module basic_1500_15000_2000_10_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_1264,In_604);
or U1 (N_1,In_531,In_496);
nand U2 (N_2,In_719,In_1020);
and U3 (N_3,In_560,In_1143);
nor U4 (N_4,In_1441,In_672);
or U5 (N_5,In_1479,In_115);
and U6 (N_6,In_415,In_1431);
or U7 (N_7,In_993,In_1254);
and U8 (N_8,In_1468,In_469);
nand U9 (N_9,In_274,In_518);
xnor U10 (N_10,In_650,In_1412);
or U11 (N_11,In_444,In_760);
and U12 (N_12,In_588,In_1274);
nand U13 (N_13,In_1373,In_543);
xor U14 (N_14,In_114,In_535);
nor U15 (N_15,In_270,In_1462);
and U16 (N_16,In_1340,In_61);
nand U17 (N_17,In_1011,In_207);
xor U18 (N_18,In_1142,In_285);
nand U19 (N_19,In_641,In_1453);
nor U20 (N_20,In_1138,In_1283);
nor U21 (N_21,In_1113,In_1115);
nand U22 (N_22,In_969,In_622);
xnor U23 (N_23,In_1211,In_554);
or U24 (N_24,In_1314,In_865);
xor U25 (N_25,In_500,In_434);
or U26 (N_26,In_1247,In_253);
xnor U27 (N_27,In_1126,In_305);
and U28 (N_28,In_1108,In_302);
nor U29 (N_29,In_1003,In_618);
xor U30 (N_30,In_1118,In_1219);
nand U31 (N_31,In_1351,In_1377);
or U32 (N_32,In_1300,In_929);
or U33 (N_33,In_1325,In_435);
xor U34 (N_34,In_866,In_325);
and U35 (N_35,In_636,In_92);
xnor U36 (N_36,In_1117,In_629);
nor U37 (N_37,In_141,In_627);
xnor U38 (N_38,In_737,In_1111);
nand U39 (N_39,In_255,In_70);
or U40 (N_40,In_833,In_1475);
and U41 (N_41,In_813,In_1469);
or U42 (N_42,In_928,In_49);
or U43 (N_43,In_1258,In_244);
nor U44 (N_44,In_35,In_726);
or U45 (N_45,In_353,In_418);
nor U46 (N_46,In_1072,In_228);
or U47 (N_47,In_177,In_212);
nand U48 (N_48,In_1225,In_220);
nand U49 (N_49,In_907,In_768);
xnor U50 (N_50,In_1363,In_473);
nor U51 (N_51,In_293,In_175);
and U52 (N_52,In_852,In_288);
xnor U53 (N_53,In_692,In_569);
nor U54 (N_54,In_861,In_989);
and U55 (N_55,In_1064,In_1365);
nor U56 (N_56,In_121,In_671);
nor U57 (N_57,In_315,In_421);
and U58 (N_58,In_1201,In_33);
nor U59 (N_59,In_593,In_830);
and U60 (N_60,In_232,In_362);
nor U61 (N_61,In_1043,In_871);
and U62 (N_62,In_1284,In_984);
and U63 (N_63,In_294,In_656);
xnor U64 (N_64,In_1311,In_669);
and U65 (N_65,In_599,In_180);
nand U66 (N_66,In_995,In_313);
or U67 (N_67,In_170,In_1195);
or U68 (N_68,In_798,In_1275);
nand U69 (N_69,In_231,In_385);
nor U70 (N_70,In_158,In_897);
and U71 (N_71,In_1161,In_1433);
nand U72 (N_72,In_1191,In_136);
nor U73 (N_73,In_783,In_1316);
xnor U74 (N_74,In_1372,In_1070);
xnor U75 (N_75,In_396,In_1477);
nor U76 (N_76,In_63,In_823);
or U77 (N_77,In_227,In_194);
and U78 (N_78,In_1151,In_475);
xnor U79 (N_79,In_748,In_499);
nor U80 (N_80,In_786,In_1063);
and U81 (N_81,In_598,In_1052);
xor U82 (N_82,In_1010,In_1327);
nand U83 (N_83,In_1307,In_159);
or U84 (N_84,In_1368,In_595);
and U85 (N_85,In_188,In_1134);
or U86 (N_86,In_246,In_1400);
nor U87 (N_87,In_279,In_1393);
and U88 (N_88,In_829,In_178);
xnor U89 (N_89,In_615,In_321);
nor U90 (N_90,In_827,In_254);
and U91 (N_91,In_1246,In_1175);
and U92 (N_92,In_44,In_163);
xor U93 (N_93,In_428,In_366);
or U94 (N_94,In_297,In_795);
nor U95 (N_95,In_1082,In_1007);
or U96 (N_96,In_195,In_624);
and U97 (N_97,In_292,In_420);
nor U98 (N_98,In_68,In_788);
nand U99 (N_99,In_1212,In_777);
nand U100 (N_100,In_1234,In_705);
nor U101 (N_101,In_509,In_12);
or U102 (N_102,In_1171,In_240);
or U103 (N_103,In_135,In_809);
and U104 (N_104,In_1374,In_609);
xnor U105 (N_105,In_432,In_34);
xnor U106 (N_106,In_26,In_967);
or U107 (N_107,In_800,In_191);
xnor U108 (N_108,In_298,In_1075);
nand U109 (N_109,In_1091,In_258);
and U110 (N_110,In_948,In_91);
xnor U111 (N_111,In_1152,In_395);
and U112 (N_112,In_520,In_525);
and U113 (N_113,In_576,In_1077);
or U114 (N_114,In_1014,In_397);
nor U115 (N_115,In_512,In_57);
or U116 (N_116,In_80,In_1490);
nor U117 (N_117,In_352,In_1170);
nor U118 (N_118,In_983,In_259);
and U119 (N_119,In_241,In_1438);
and U120 (N_120,In_284,In_1062);
or U121 (N_121,In_1001,In_822);
or U122 (N_122,In_763,In_710);
nor U123 (N_123,In_371,In_693);
or U124 (N_124,In_713,In_562);
or U125 (N_125,In_1390,In_447);
nor U126 (N_126,In_476,In_1244);
nand U127 (N_127,In_649,In_167);
nor U128 (N_128,In_433,In_660);
or U129 (N_129,In_106,In_935);
or U130 (N_130,In_832,In_899);
xor U131 (N_131,In_1147,In_1360);
nor U132 (N_132,In_387,In_470);
and U133 (N_133,In_775,In_105);
nor U134 (N_134,In_377,In_966);
xor U135 (N_135,In_938,In_1202);
and U136 (N_136,In_790,In_482);
and U137 (N_137,In_1491,In_139);
or U138 (N_138,In_1173,In_217);
xor U139 (N_139,In_320,In_900);
or U140 (N_140,In_546,In_1228);
or U141 (N_141,In_516,In_1252);
xor U142 (N_142,In_1455,In_1016);
nor U143 (N_143,In_547,In_1496);
nor U144 (N_144,In_480,In_908);
nand U145 (N_145,In_417,In_1447);
or U146 (N_146,In_683,In_128);
nor U147 (N_147,In_489,In_1405);
and U148 (N_148,In_621,In_1317);
nor U149 (N_149,In_508,In_1304);
nand U150 (N_150,In_1250,In_970);
or U151 (N_151,In_374,In_961);
nand U152 (N_152,In_1487,In_247);
xnor U153 (N_153,In_881,In_1299);
and U154 (N_154,In_787,In_1277);
and U155 (N_155,In_174,In_1087);
nand U156 (N_156,In_1124,In_424);
nand U157 (N_157,In_811,In_205);
or U158 (N_158,In_962,In_1039);
nand U159 (N_159,In_601,In_715);
and U160 (N_160,In_1426,In_917);
or U161 (N_161,In_124,In_1055);
nor U162 (N_162,In_1302,In_986);
or U163 (N_163,In_687,In_684);
and U164 (N_164,In_441,In_81);
xnor U165 (N_165,In_653,In_379);
nor U166 (N_166,In_774,In_836);
nand U167 (N_167,In_341,In_1473);
xnor U168 (N_168,In_797,In_982);
or U169 (N_169,In_407,In_514);
and U170 (N_170,In_754,In_125);
xor U171 (N_171,In_1230,In_893);
or U172 (N_172,In_219,In_1413);
xor U173 (N_173,In_197,In_1318);
nor U174 (N_174,In_1410,In_349);
nor U175 (N_175,In_152,In_161);
nor U176 (N_176,In_1189,In_607);
and U177 (N_177,In_41,In_845);
or U178 (N_178,In_766,In_1498);
or U179 (N_179,In_506,In_591);
nand U180 (N_180,In_154,In_815);
xnor U181 (N_181,In_1294,In_1125);
or U182 (N_182,In_991,In_701);
nand U183 (N_183,In_700,In_102);
xnor U184 (N_184,In_97,In_1397);
xor U185 (N_185,In_1345,In_276);
nor U186 (N_186,In_1388,In_1429);
nand U187 (N_187,In_388,In_1464);
nor U188 (N_188,In_1236,In_59);
xor U189 (N_189,In_443,In_734);
nand U190 (N_190,In_182,In_873);
nor U191 (N_191,In_1404,In_1216);
or U192 (N_192,In_582,In_1364);
nor U193 (N_193,In_1367,In_1110);
and U194 (N_194,In_585,In_877);
or U195 (N_195,In_130,In_612);
and U196 (N_196,In_1199,In_1215);
nor U197 (N_197,In_1094,In_1000);
nand U198 (N_198,In_816,In_1492);
nor U199 (N_199,In_333,In_390);
or U200 (N_200,In_1458,In_818);
or U201 (N_201,In_376,In_56);
or U202 (N_202,In_580,In_1459);
xor U203 (N_203,In_1423,In_51);
nor U204 (N_204,In_1478,In_256);
nand U205 (N_205,In_1029,In_1306);
and U206 (N_206,In_450,In_1352);
nand U207 (N_207,In_1044,In_100);
and U208 (N_208,In_1078,In_1164);
nor U209 (N_209,In_427,In_556);
nand U210 (N_210,In_488,In_453);
and U211 (N_211,In_1241,In_1023);
nor U212 (N_212,In_237,In_381);
nand U213 (N_213,In_1223,In_640);
or U214 (N_214,In_160,In_803);
or U215 (N_215,In_913,In_31);
nand U216 (N_216,In_1132,In_1406);
xor U217 (N_217,In_312,In_586);
nor U218 (N_218,In_211,In_1021);
xor U219 (N_219,In_883,In_156);
xnor U220 (N_220,In_1398,In_805);
nor U221 (N_221,In_1148,In_1452);
nor U222 (N_222,In_1030,In_120);
nor U223 (N_223,In_1386,In_72);
nor U224 (N_224,In_1081,In_1424);
xor U225 (N_225,In_630,In_1494);
and U226 (N_226,In_1349,In_226);
xnor U227 (N_227,In_817,In_215);
or U228 (N_228,In_1335,In_1288);
or U229 (N_229,In_245,In_950);
xnor U230 (N_230,In_584,In_310);
or U231 (N_231,In_3,In_625);
and U232 (N_232,In_1184,In_771);
and U233 (N_233,In_1017,In_412);
and U234 (N_234,In_1483,In_229);
nand U235 (N_235,In_1050,In_725);
or U236 (N_236,In_268,In_411);
xor U237 (N_237,In_402,In_637);
or U238 (N_238,In_1012,In_25);
nand U239 (N_239,In_372,In_394);
and U240 (N_240,In_1319,In_451);
nor U241 (N_241,In_755,In_467);
nand U242 (N_242,In_38,In_1339);
nor U243 (N_243,In_537,In_272);
or U244 (N_244,In_1235,In_351);
nand U245 (N_245,In_1322,In_1231);
or U246 (N_246,In_1,In_466);
nand U247 (N_247,In_1119,In_662);
and U248 (N_248,In_1137,In_1032);
nor U249 (N_249,In_842,In_931);
or U250 (N_250,In_958,In_848);
nor U251 (N_251,In_1221,In_721);
nand U252 (N_252,In_691,In_1217);
nand U253 (N_253,In_183,In_510);
nand U254 (N_254,In_323,In_64);
or U255 (N_255,In_730,In_1061);
nand U256 (N_256,In_670,In_126);
and U257 (N_257,In_1018,In_378);
or U258 (N_258,In_565,In_925);
nand U259 (N_259,In_736,In_1355);
nor U260 (N_260,In_990,In_934);
nor U261 (N_261,In_753,In_1303);
and U262 (N_262,In_1331,In_493);
and U263 (N_263,In_561,In_1154);
nand U264 (N_264,In_155,In_1460);
nand U265 (N_265,In_794,In_262);
nand U266 (N_266,In_487,In_1396);
xor U267 (N_267,In_1315,In_769);
and U268 (N_268,In_360,In_578);
nand U269 (N_269,In_214,In_694);
nor U270 (N_270,In_311,In_1379);
and U271 (N_271,In_146,In_511);
and U272 (N_272,In_1463,In_939);
xor U273 (N_273,In_67,In_749);
and U274 (N_274,In_923,In_895);
xnor U275 (N_275,In_812,In_551);
and U276 (N_276,In_463,In_644);
or U277 (N_277,In_633,In_46);
and U278 (N_278,In_1196,In_1414);
and U279 (N_279,In_828,In_666);
nand U280 (N_280,In_265,In_359);
xor U281 (N_281,In_416,In_5);
and U282 (N_282,In_1204,In_1287);
or U283 (N_283,In_1457,In_738);
nand U284 (N_284,In_697,In_1358);
or U285 (N_285,In_957,In_810);
nor U286 (N_286,In_223,In_614);
nor U287 (N_287,In_706,In_342);
and U288 (N_288,In_550,In_403);
and U289 (N_289,In_304,In_890);
nand U290 (N_290,In_1430,In_1272);
or U291 (N_291,In_731,In_968);
nor U292 (N_292,In_1357,In_847);
or U293 (N_293,In_233,In_1146);
and U294 (N_294,In_712,In_1408);
nor U295 (N_295,In_912,In_383);
xnor U296 (N_296,In_1178,In_885);
xor U297 (N_297,In_54,In_147);
nor U298 (N_298,In_841,In_117);
nor U299 (N_299,In_1323,In_875);
nand U300 (N_300,In_109,In_1180);
nor U301 (N_301,In_951,In_1093);
xor U302 (N_302,In_704,In_1172);
nor U303 (N_303,In_95,In_1359);
nor U304 (N_304,In_485,In_1298);
or U305 (N_305,In_679,In_430);
xor U306 (N_306,In_1454,In_856);
xor U307 (N_307,In_239,In_620);
xor U308 (N_308,In_1167,In_826);
xor U309 (N_309,In_896,In_698);
and U310 (N_310,In_477,In_490);
xnor U311 (N_311,In_1428,In_1045);
and U312 (N_312,In_186,In_1025);
nor U313 (N_313,In_198,In_558);
xor U314 (N_314,In_918,In_542);
nor U315 (N_315,In_355,In_501);
xnor U316 (N_316,In_1289,In_1107);
xnor U317 (N_317,In_752,In_727);
nand U318 (N_318,In_1290,In_1227);
nor U319 (N_319,In_527,In_1391);
nand U320 (N_320,In_122,In_502);
xor U321 (N_321,In_567,In_1467);
nand U322 (N_322,In_440,In_651);
or U323 (N_323,In_235,In_1347);
xor U324 (N_324,In_399,In_203);
or U325 (N_325,In_718,In_657);
xnor U326 (N_326,In_47,In_555);
xor U327 (N_327,In_1008,In_464);
and U328 (N_328,In_1135,In_76);
xnor U329 (N_329,In_62,In_600);
nand U330 (N_330,In_523,In_807);
and U331 (N_331,In_665,In_437);
or U332 (N_332,In_613,In_521);
or U333 (N_333,In_368,In_1471);
or U334 (N_334,In_1004,In_1472);
nand U335 (N_335,In_1425,In_872);
nor U336 (N_336,In_481,In_208);
xor U337 (N_337,In_1450,In_1165);
and U338 (N_338,In_740,In_491);
or U339 (N_339,In_677,In_932);
and U340 (N_340,In_921,In_1402);
nor U341 (N_341,In_347,In_1337);
and U342 (N_342,In_414,In_854);
and U343 (N_343,In_78,In_659);
nand U344 (N_344,In_324,In_1489);
and U345 (N_345,In_112,In_1076);
nor U346 (N_346,In_486,In_448);
nand U347 (N_347,In_619,In_953);
nor U348 (N_348,In_1185,In_1033);
xor U349 (N_349,In_111,In_1238);
nor U350 (N_350,In_894,In_1129);
nor U351 (N_351,In_1069,In_295);
nor U352 (N_352,In_18,In_1278);
nor U353 (N_353,In_1361,In_66);
or U354 (N_354,In_911,In_171);
and U355 (N_355,In_632,In_184);
nand U356 (N_356,In_90,In_709);
nand U357 (N_357,In_389,In_99);
xnor U358 (N_358,In_1401,In_1286);
or U359 (N_359,In_1149,In_1197);
xor U360 (N_360,In_446,In_597);
or U361 (N_361,In_398,In_747);
and U362 (N_362,In_83,In_1255);
and U363 (N_363,In_977,In_792);
and U364 (N_364,In_716,In_1047);
xnor U365 (N_365,In_785,In_901);
nor U366 (N_366,In_1326,In_834);
xor U367 (N_367,In_344,In_1267);
or U368 (N_368,In_548,In_201);
or U369 (N_369,In_1205,In_218);
and U370 (N_370,In_20,In_1495);
xor U371 (N_371,In_634,In_965);
nand U372 (N_372,In_994,In_1269);
nor U373 (N_373,In_1085,In_1329);
nand U374 (N_374,In_140,In_744);
or U375 (N_375,In_616,In_350);
or U376 (N_376,In_1305,In_71);
nor U377 (N_377,In_1336,In_519);
nand U378 (N_378,In_1207,In_1394);
nor U379 (N_379,In_316,In_257);
nor U380 (N_380,In_166,In_855);
nand U381 (N_381,In_1210,In_606);
nor U382 (N_382,In_639,In_1160);
nand U383 (N_383,In_438,In_1240);
nand U384 (N_384,In_1024,In_442);
and U385 (N_385,In_1169,In_789);
nor U386 (N_386,In_1259,In_686);
or U387 (N_387,In_973,In_814);
or U388 (N_388,In_552,In_234);
nand U389 (N_389,In_583,In_859);
and U390 (N_390,In_264,In_707);
nand U391 (N_391,In_1066,In_116);
or U392 (N_392,In_356,In_964);
nand U393 (N_393,In_674,In_972);
xnor U394 (N_394,In_39,In_27);
and U395 (N_395,In_676,In_858);
xor U396 (N_396,In_714,In_1439);
or U397 (N_397,In_457,In_667);
nand U398 (N_398,In_1268,In_910);
nand U399 (N_399,In_844,In_978);
or U400 (N_400,In_1470,In_592);
nand U401 (N_401,In_802,In_190);
or U402 (N_402,In_123,In_210);
nor U403 (N_403,In_340,In_162);
and U404 (N_404,In_914,In_84);
and U405 (N_405,In_24,In_127);
nor U406 (N_406,In_1333,In_1432);
or U407 (N_407,In_946,In_425);
nand U408 (N_408,In_761,In_1291);
and U409 (N_409,In_472,In_997);
nand U410 (N_410,In_53,In_6);
nor U411 (N_411,In_1101,In_98);
and U412 (N_412,In_617,In_299);
nor U413 (N_413,In_626,In_455);
nor U414 (N_414,In_436,In_1153);
and U415 (N_415,In_1209,In_678);
nor U416 (N_416,In_1266,In_87);
nor U417 (N_417,In_176,In_505);
nand U418 (N_418,In_157,In_887);
and U419 (N_419,In_974,In_1198);
xor U420 (N_420,In_750,In_43);
and U421 (N_421,In_118,In_916);
nor U422 (N_422,In_857,In_878);
nor U423 (N_423,In_48,In_263);
or U424 (N_424,In_1177,In_1086);
and U425 (N_425,In_898,In_1140);
and U426 (N_426,In_942,In_780);
nor U427 (N_427,In_1222,In_1249);
and U428 (N_428,In_1488,In_1366);
nand U429 (N_429,In_1163,In_1485);
nand U430 (N_430,In_1369,In_1395);
xor U431 (N_431,In_746,In_1059);
nand U432 (N_432,In_1418,In_365);
nand U433 (N_433,In_138,In_1451);
nand U434 (N_434,In_13,In_148);
nand U435 (N_435,In_764,In_926);
nand U436 (N_436,In_361,In_431);
xnor U437 (N_437,In_1192,In_22);
xor U438 (N_438,In_423,In_539);
and U439 (N_439,In_30,In_937);
or U440 (N_440,In_52,In_759);
and U441 (N_441,In_1200,In_963);
nor U442 (N_442,In_1054,In_1292);
nor U443 (N_443,In_658,In_1053);
nor U444 (N_444,In_602,In_1038);
nor U445 (N_445,In_1174,In_532);
xor U446 (N_446,In_196,In_849);
and U447 (N_447,In_1461,In_999);
or U448 (N_448,In_456,In_835);
xor U449 (N_449,In_346,In_9);
and U450 (N_450,In_1068,In_1090);
or U451 (N_451,In_471,In_979);
nand U452 (N_452,In_1042,In_1122);
nand U453 (N_453,In_892,In_1145);
nor U454 (N_454,In_82,In_507);
nand U455 (N_455,In_1067,In_544);
xnor U456 (N_456,In_400,In_133);
or U457 (N_457,In_1446,In_1338);
xor U458 (N_458,In_867,In_663);
xor U459 (N_459,In_93,In_1407);
nand U460 (N_460,In_296,In_648);
and U461 (N_461,In_851,In_1261);
xor U462 (N_462,In_426,In_1481);
or U463 (N_463,In_336,In_202);
or U464 (N_464,In_758,In_1098);
nor U465 (N_465,In_206,In_603);
xor U466 (N_466,In_1301,In_1420);
and U467 (N_467,In_267,In_909);
nor U468 (N_468,In_308,In_454);
xor U469 (N_469,In_661,In_149);
or U470 (N_470,In_708,In_549);
nor U471 (N_471,In_1476,In_1232);
nor U472 (N_472,In_652,In_1334);
nor U473 (N_473,In_976,In_280);
nor U474 (N_474,In_17,In_1048);
xor U475 (N_475,In_307,In_742);
nor U476 (N_476,In_1380,In_363);
and U477 (N_477,In_401,In_791);
nor U478 (N_478,In_281,In_497);
or U479 (N_479,In_1220,In_404);
xor U480 (N_480,In_1088,In_1034);
or U481 (N_481,In_86,In_209);
nand U482 (N_482,In_131,In_1436);
xnor U483 (N_483,In_940,In_1256);
nor U484 (N_484,In_225,In_992);
nor U485 (N_485,In_793,In_904);
and U486 (N_486,In_906,In_271);
and U487 (N_487,In_1448,In_696);
nand U488 (N_488,In_605,In_581);
nor U489 (N_489,In_572,In_882);
xnor U490 (N_490,In_1381,In_77);
or U491 (N_491,In_1350,In_862);
xor U492 (N_492,In_1265,In_28);
nand U493 (N_493,In_870,In_169);
or U494 (N_494,In_2,In_1005);
nand U495 (N_495,In_419,In_1348);
or U496 (N_496,In_1031,In_1282);
nor U497 (N_497,In_1409,In_1186);
xnor U498 (N_498,In_50,In_729);
nor U499 (N_499,In_413,In_1141);
and U500 (N_500,In_1058,In_1296);
xor U501 (N_501,In_335,In_492);
xnor U502 (N_502,In_1271,In_513);
xor U503 (N_503,In_494,In_949);
xnor U504 (N_504,In_981,In_1187);
or U505 (N_505,In_944,In_1466);
or U506 (N_506,In_1037,In_886);
and U507 (N_507,In_1028,In_277);
nor U508 (N_508,In_1486,In_647);
or U509 (N_509,In_724,In_1179);
xnor U510 (N_510,In_732,In_96);
xnor U511 (N_511,In_1324,In_1226);
and U512 (N_512,In_998,In_801);
or U513 (N_513,In_348,In_664);
nand U514 (N_514,In_1166,In_29);
or U515 (N_515,In_685,In_60);
or U516 (N_516,In_846,In_947);
xor U517 (N_517,In_960,In_462);
nor U518 (N_518,In_1100,In_1310);
nand U519 (N_519,In_689,In_1130);
nor U520 (N_520,In_1239,In_108);
xor U521 (N_521,In_1112,In_273);
or U522 (N_522,In_1083,In_1474);
and U523 (N_523,In_1136,In_1009);
xor U524 (N_524,In_289,In_825);
or U525 (N_525,In_319,In_461);
nor U526 (N_526,In_199,In_1121);
nand U527 (N_527,In_216,In_11);
xnor U528 (N_528,In_975,In_819);
and U529 (N_529,In_1080,In_902);
nand U530 (N_530,In_1279,In_1041);
or U531 (N_531,In_1482,In_172);
nand U532 (N_532,In_831,In_393);
xnor U533 (N_533,In_317,In_611);
xnor U534 (N_534,In_474,In_1353);
xnor U535 (N_535,In_610,In_369);
xor U536 (N_536,In_779,In_375);
or U537 (N_537,In_1293,In_339);
nand U538 (N_538,In_1362,In_32);
nor U539 (N_539,In_1057,In_309);
xor U540 (N_540,In_1084,In_460);
xnor U541 (N_541,In_1060,In_23);
nor U542 (N_542,In_132,In_1285);
xnor U543 (N_543,In_820,In_107);
nand U544 (N_544,In_517,In_524);
xor U545 (N_545,In_269,In_1444);
xor U546 (N_546,In_837,In_327);
and U547 (N_547,In_1309,In_1123);
and U548 (N_548,In_690,In_380);
nand U549 (N_549,In_903,In_1182);
or U550 (N_550,In_1168,In_688);
and U551 (N_551,In_682,In_282);
xnor U552 (N_552,In_74,In_1183);
nor U553 (N_553,In_249,In_699);
and U554 (N_554,In_422,In_367);
xnor U555 (N_555,In_996,In_557);
nand U556 (N_556,In_1208,In_589);
nor U557 (N_557,In_668,In_596);
or U558 (N_558,In_142,In_1276);
or U559 (N_559,In_943,In_1242);
and U560 (N_560,In_113,In_250);
and U561 (N_561,In_574,In_1206);
and U562 (N_562,In_876,In_1035);
nor U563 (N_563,In_1442,In_635);
xnor U564 (N_564,In_15,In_1036);
nand U565 (N_565,In_345,In_728);
nor U566 (N_566,In_631,In_338);
xor U567 (N_567,In_329,In_330);
xnor U568 (N_568,In_1027,In_0);
nand U569 (N_569,In_65,In_465);
xnor U570 (N_570,In_628,In_1181);
nor U571 (N_571,In_252,In_370);
nand U572 (N_572,In_545,In_533);
and U573 (N_573,In_781,In_743);
nor U574 (N_574,In_409,In_1421);
or U575 (N_575,In_7,In_21);
nand U576 (N_576,In_608,In_566);
xor U577 (N_577,In_1332,In_1229);
nand U578 (N_578,In_1190,In_364);
or U579 (N_579,In_1382,In_645);
nor U580 (N_580,In_880,In_1213);
nand U581 (N_581,In_1026,In_88);
nor U582 (N_582,In_1158,In_1176);
xnor U583 (N_583,In_326,In_129);
or U584 (N_584,In_868,In_1378);
or U585 (N_585,In_538,In_741);
nand U586 (N_586,In_702,In_55);
or U587 (N_587,In_1096,In_623);
or U588 (N_588,In_515,In_69);
and U589 (N_589,In_980,In_1218);
nand U590 (N_590,In_429,In_590);
nor U591 (N_591,In_843,In_382);
nand U592 (N_592,In_1243,In_1434);
or U593 (N_593,In_1341,In_1342);
nand U594 (N_594,In_1013,In_1371);
xor U595 (N_595,In_568,In_778);
xor U596 (N_596,In_230,In_1370);
nor U597 (N_597,In_776,In_1403);
nand U598 (N_598,In_577,In_571);
nor U599 (N_599,In_722,In_654);
or U600 (N_600,In_915,In_408);
or U601 (N_601,In_459,In_1480);
or U602 (N_602,In_1049,In_526);
xnor U603 (N_603,In_1437,In_36);
xnor U604 (N_604,In_1389,In_278);
nor U605 (N_605,In_1263,In_185);
and U606 (N_606,In_594,In_151);
nand U607 (N_607,In_1015,In_181);
xnor U608 (N_608,In_449,In_756);
nor U609 (N_609,In_1273,In_1109);
nor U610 (N_610,In_806,In_406);
nand U611 (N_611,In_1392,In_1074);
xnor U612 (N_612,In_1106,In_1384);
and U613 (N_613,In_1375,In_222);
xnor U614 (N_614,In_373,In_933);
xor U615 (N_615,In_522,In_19);
xor U616 (N_616,In_1104,In_75);
nand U617 (N_617,In_879,In_955);
nand U618 (N_618,In_173,In_1281);
or U619 (N_619,In_498,In_204);
nor U620 (N_620,In_804,In_103);
and U621 (N_621,In_733,In_261);
nor U622 (N_622,In_528,In_290);
and U623 (N_623,In_874,In_286);
or U624 (N_624,In_1116,In_1105);
xnor U625 (N_625,In_1399,In_1193);
xnor U626 (N_626,In_720,In_439);
or U627 (N_627,In_1155,In_1383);
or U628 (N_628,In_1046,In_1120);
nand U629 (N_629,In_717,In_936);
xor U630 (N_630,In_1065,In_808);
xnor U631 (N_631,In_8,In_642);
xnor U632 (N_632,In_1343,In_553);
or U633 (N_633,In_1295,In_905);
or U634 (N_634,In_1214,In_988);
or U635 (N_635,In_1385,In_559);
nand U636 (N_636,In_959,In_1097);
nand U637 (N_637,In_134,In_1449);
or U638 (N_638,In_314,In_1194);
nand U639 (N_639,In_985,In_248);
nor U640 (N_640,In_4,In_1328);
and U641 (N_641,In_187,In_484);
nand U642 (N_642,In_927,In_1330);
xnor U643 (N_643,In_920,In_1128);
and U644 (N_644,In_840,In_573);
or U645 (N_645,In_483,In_85);
nand U646 (N_646,In_673,In_1262);
or U647 (N_647,In_945,In_541);
or U648 (N_648,In_1422,In_655);
nand U649 (N_649,In_318,In_1144);
or U650 (N_650,In_334,In_1245);
and U651 (N_651,In_1280,In_343);
nor U652 (N_652,In_889,In_153);
xor U653 (N_653,In_735,In_579);
or U654 (N_654,In_838,In_322);
nand U655 (N_655,In_745,In_1002);
and U656 (N_656,In_530,In_79);
nor U657 (N_657,In_675,In_1440);
xnor U658 (N_658,In_332,In_110);
and U659 (N_659,In_260,In_1387);
or U660 (N_660,In_1312,In_638);
or U661 (N_661,In_1435,In_213);
and U662 (N_662,In_1260,In_445);
or U663 (N_663,In_1019,In_1376);
nor U664 (N_664,In_1416,In_479);
nor U665 (N_665,In_236,In_145);
nand U666 (N_666,In_495,In_243);
and U667 (N_667,In_919,In_410);
nor U668 (N_668,In_1257,In_405);
xor U669 (N_669,In_1308,In_824);
xor U670 (N_670,In_1443,In_238);
or U671 (N_671,In_587,In_762);
and U672 (N_672,In_799,In_189);
xor U673 (N_673,In_1248,In_89);
nand U674 (N_674,In_767,In_952);
and U675 (N_675,In_971,In_1499);
xnor U676 (N_676,In_1022,In_956);
nand U677 (N_677,In_540,In_392);
xnor U678 (N_678,In_751,In_863);
nor U679 (N_679,In_303,In_144);
nor U680 (N_680,In_821,In_357);
or U681 (N_681,In_1127,In_10);
and U682 (N_682,In_143,In_1095);
or U683 (N_683,In_1150,In_1162);
nand U684 (N_684,In_504,In_850);
nor U685 (N_685,In_1139,In_723);
nand U686 (N_686,In_1133,In_891);
and U687 (N_687,In_42,In_37);
nand U688 (N_688,In_864,In_681);
and U689 (N_689,In_1270,In_16);
nor U690 (N_690,In_137,In_1251);
nor U691 (N_691,In_168,In_853);
nand U692 (N_692,In_680,In_884);
nand U693 (N_693,In_242,In_529);
nand U694 (N_694,In_1415,In_192);
nor U695 (N_695,In_987,In_1427);
and U696 (N_696,In_458,In_924);
nand U697 (N_697,In_104,In_784);
nand U698 (N_698,In_757,In_1103);
nor U699 (N_699,In_224,In_1354);
nand U700 (N_700,In_1321,In_1411);
and U701 (N_701,In_1073,In_391);
and U702 (N_702,In_94,In_1131);
nand U703 (N_703,In_922,In_1224);
nor U704 (N_704,In_1465,In_287);
or U705 (N_705,In_283,In_1089);
xor U706 (N_706,In_1484,In_1006);
nor U707 (N_707,In_1159,In_300);
nand U708 (N_708,In_1099,In_14);
and U709 (N_709,In_101,In_468);
or U710 (N_710,In_1233,In_1493);
and U711 (N_711,In_1497,In_73);
and U712 (N_712,In_739,In_1156);
nand U713 (N_713,In_1237,In_1320);
nand U714 (N_714,In_306,In_860);
xnor U715 (N_715,In_1417,In_1040);
and U716 (N_716,In_266,In_1456);
and U717 (N_717,In_570,In_1114);
or U718 (N_718,In_888,In_1157);
and U719 (N_719,In_1313,In_954);
and U720 (N_720,In_1051,In_646);
nor U721 (N_721,In_251,In_193);
or U722 (N_722,In_1253,In_358);
or U723 (N_723,In_164,In_1445);
nand U724 (N_724,In_839,In_165);
or U725 (N_725,In_711,In_45);
nor U726 (N_726,In_575,In_119);
or U727 (N_727,In_1346,In_1188);
nand U728 (N_728,In_40,In_563);
or U729 (N_729,In_796,In_534);
xor U730 (N_730,In_695,In_930);
and U731 (N_731,In_1092,In_773);
xnor U732 (N_732,In_275,In_1356);
nand U733 (N_733,In_354,In_1297);
xnor U734 (N_734,In_782,In_150);
nor U735 (N_735,In_941,In_301);
or U736 (N_736,In_478,In_564);
and U737 (N_737,In_386,In_1419);
nand U738 (N_738,In_772,In_328);
nand U739 (N_739,In_221,In_384);
xnor U740 (N_740,In_291,In_1056);
nor U741 (N_741,In_337,In_200);
or U742 (N_742,In_536,In_452);
xor U743 (N_743,In_1203,In_1079);
or U744 (N_744,In_643,In_869);
or U745 (N_745,In_770,In_1344);
and U746 (N_746,In_703,In_331);
nand U747 (N_747,In_179,In_503);
or U748 (N_748,In_58,In_1102);
xnor U749 (N_749,In_1071,In_765);
or U750 (N_750,In_693,In_159);
or U751 (N_751,In_289,In_82);
nor U752 (N_752,In_573,In_611);
nand U753 (N_753,In_1413,In_1356);
nor U754 (N_754,In_519,In_1000);
or U755 (N_755,In_312,In_383);
xnor U756 (N_756,In_760,In_1138);
or U757 (N_757,In_1291,In_1177);
xor U758 (N_758,In_707,In_515);
nand U759 (N_759,In_221,In_202);
and U760 (N_760,In_59,In_361);
and U761 (N_761,In_1260,In_1023);
nor U762 (N_762,In_1059,In_539);
nand U763 (N_763,In_563,In_157);
xnor U764 (N_764,In_1026,In_1040);
nor U765 (N_765,In_104,In_910);
nor U766 (N_766,In_932,In_1485);
nand U767 (N_767,In_514,In_377);
xnor U768 (N_768,In_1214,In_956);
nand U769 (N_769,In_1129,In_705);
nor U770 (N_770,In_1189,In_1111);
or U771 (N_771,In_888,In_780);
xnor U772 (N_772,In_1054,In_1313);
xor U773 (N_773,In_1393,In_879);
xnor U774 (N_774,In_1380,In_1169);
or U775 (N_775,In_301,In_1149);
and U776 (N_776,In_1425,In_316);
and U777 (N_777,In_1141,In_964);
or U778 (N_778,In_139,In_11);
and U779 (N_779,In_343,In_1054);
and U780 (N_780,In_1483,In_131);
nor U781 (N_781,In_1346,In_472);
nand U782 (N_782,In_1423,In_893);
nand U783 (N_783,In_1465,In_1409);
xnor U784 (N_784,In_413,In_800);
or U785 (N_785,In_1235,In_192);
nand U786 (N_786,In_129,In_1498);
and U787 (N_787,In_1228,In_667);
and U788 (N_788,In_1295,In_827);
and U789 (N_789,In_946,In_944);
and U790 (N_790,In_564,In_88);
or U791 (N_791,In_532,In_21);
xor U792 (N_792,In_1348,In_934);
or U793 (N_793,In_588,In_416);
and U794 (N_794,In_687,In_346);
xor U795 (N_795,In_771,In_251);
nor U796 (N_796,In_918,In_1367);
nor U797 (N_797,In_1302,In_482);
nor U798 (N_798,In_67,In_295);
and U799 (N_799,In_718,In_1250);
xnor U800 (N_800,In_1108,In_139);
nand U801 (N_801,In_131,In_229);
and U802 (N_802,In_850,In_122);
xor U803 (N_803,In_1326,In_1155);
nor U804 (N_804,In_215,In_1211);
nor U805 (N_805,In_1146,In_627);
nor U806 (N_806,In_799,In_1074);
nor U807 (N_807,In_1177,In_953);
nor U808 (N_808,In_1100,In_58);
nand U809 (N_809,In_1047,In_579);
nand U810 (N_810,In_1436,In_314);
or U811 (N_811,In_1079,In_1130);
and U812 (N_812,In_140,In_587);
nor U813 (N_813,In_256,In_461);
and U814 (N_814,In_1348,In_962);
nor U815 (N_815,In_1382,In_446);
xor U816 (N_816,In_1082,In_163);
xor U817 (N_817,In_281,In_642);
xnor U818 (N_818,In_821,In_583);
nor U819 (N_819,In_524,In_591);
nor U820 (N_820,In_1051,In_766);
nand U821 (N_821,In_1100,In_975);
xnor U822 (N_822,In_184,In_1357);
or U823 (N_823,In_1125,In_1473);
and U824 (N_824,In_305,In_468);
xnor U825 (N_825,In_1276,In_1142);
or U826 (N_826,In_489,In_728);
nand U827 (N_827,In_231,In_228);
nor U828 (N_828,In_46,In_882);
xnor U829 (N_829,In_859,In_232);
nor U830 (N_830,In_256,In_695);
nand U831 (N_831,In_870,In_540);
nand U832 (N_832,In_84,In_1238);
nor U833 (N_833,In_1001,In_551);
and U834 (N_834,In_890,In_897);
or U835 (N_835,In_1031,In_566);
or U836 (N_836,In_85,In_446);
or U837 (N_837,In_887,In_715);
nand U838 (N_838,In_376,In_1012);
or U839 (N_839,In_170,In_1136);
nand U840 (N_840,In_298,In_612);
nor U841 (N_841,In_50,In_817);
nand U842 (N_842,In_800,In_634);
or U843 (N_843,In_315,In_819);
and U844 (N_844,In_531,In_1340);
and U845 (N_845,In_733,In_570);
and U846 (N_846,In_47,In_378);
or U847 (N_847,In_1453,In_1482);
or U848 (N_848,In_1158,In_1038);
nor U849 (N_849,In_1436,In_572);
and U850 (N_850,In_1160,In_525);
xnor U851 (N_851,In_755,In_856);
xnor U852 (N_852,In_948,In_1281);
or U853 (N_853,In_665,In_19);
nor U854 (N_854,In_672,In_1468);
or U855 (N_855,In_1223,In_1340);
nand U856 (N_856,In_367,In_510);
nor U857 (N_857,In_192,In_92);
xor U858 (N_858,In_1185,In_463);
nor U859 (N_859,In_1016,In_479);
nand U860 (N_860,In_1277,In_423);
or U861 (N_861,In_185,In_1486);
xor U862 (N_862,In_749,In_306);
and U863 (N_863,In_562,In_125);
or U864 (N_864,In_304,In_247);
xnor U865 (N_865,In_571,In_1346);
or U866 (N_866,In_200,In_420);
and U867 (N_867,In_215,In_1086);
nor U868 (N_868,In_947,In_949);
nand U869 (N_869,In_171,In_88);
or U870 (N_870,In_111,In_808);
nor U871 (N_871,In_601,In_1355);
and U872 (N_872,In_233,In_619);
and U873 (N_873,In_508,In_417);
nand U874 (N_874,In_279,In_37);
and U875 (N_875,In_703,In_1195);
nand U876 (N_876,In_319,In_980);
or U877 (N_877,In_464,In_385);
xnor U878 (N_878,In_345,In_803);
or U879 (N_879,In_1373,In_545);
nand U880 (N_880,In_1408,In_1030);
nor U881 (N_881,In_412,In_1);
xor U882 (N_882,In_743,In_327);
nor U883 (N_883,In_931,In_989);
xnor U884 (N_884,In_962,In_779);
nand U885 (N_885,In_1412,In_1208);
xnor U886 (N_886,In_1218,In_403);
xor U887 (N_887,In_893,In_218);
nor U888 (N_888,In_1408,In_1130);
and U889 (N_889,In_856,In_317);
and U890 (N_890,In_972,In_1067);
and U891 (N_891,In_57,In_768);
nor U892 (N_892,In_49,In_1341);
and U893 (N_893,In_372,In_106);
nand U894 (N_894,In_788,In_1032);
and U895 (N_895,In_1213,In_303);
xor U896 (N_896,In_573,In_1012);
nand U897 (N_897,In_995,In_10);
nor U898 (N_898,In_1131,In_1174);
or U899 (N_899,In_227,In_281);
nor U900 (N_900,In_93,In_673);
nand U901 (N_901,In_829,In_1493);
and U902 (N_902,In_18,In_847);
nor U903 (N_903,In_412,In_431);
and U904 (N_904,In_477,In_1182);
and U905 (N_905,In_1084,In_421);
and U906 (N_906,In_858,In_374);
or U907 (N_907,In_1083,In_1186);
xnor U908 (N_908,In_1131,In_1034);
xnor U909 (N_909,In_671,In_1436);
xor U910 (N_910,In_1247,In_905);
xor U911 (N_911,In_232,In_1467);
and U912 (N_912,In_66,In_787);
and U913 (N_913,In_1236,In_1353);
or U914 (N_914,In_350,In_1010);
and U915 (N_915,In_141,In_1250);
or U916 (N_916,In_863,In_1174);
or U917 (N_917,In_1046,In_261);
xor U918 (N_918,In_1449,In_1427);
or U919 (N_919,In_773,In_1492);
and U920 (N_920,In_1173,In_291);
nor U921 (N_921,In_762,In_1465);
and U922 (N_922,In_712,In_521);
nor U923 (N_923,In_594,In_668);
or U924 (N_924,In_1042,In_27);
nand U925 (N_925,In_280,In_816);
or U926 (N_926,In_553,In_1244);
and U927 (N_927,In_436,In_1334);
nand U928 (N_928,In_17,In_891);
xnor U929 (N_929,In_99,In_770);
nor U930 (N_930,In_1066,In_1461);
xnor U931 (N_931,In_1110,In_632);
xnor U932 (N_932,In_343,In_161);
or U933 (N_933,In_1449,In_928);
and U934 (N_934,In_1038,In_579);
nand U935 (N_935,In_262,In_1327);
nor U936 (N_936,In_1288,In_663);
and U937 (N_937,In_520,In_474);
nor U938 (N_938,In_1052,In_273);
or U939 (N_939,In_78,In_188);
nor U940 (N_940,In_220,In_1295);
nand U941 (N_941,In_69,In_1221);
nor U942 (N_942,In_946,In_985);
and U943 (N_943,In_319,In_299);
or U944 (N_944,In_1461,In_237);
xor U945 (N_945,In_1494,In_1052);
or U946 (N_946,In_729,In_1160);
nor U947 (N_947,In_881,In_780);
nor U948 (N_948,In_661,In_157);
nor U949 (N_949,In_1162,In_1307);
nor U950 (N_950,In_218,In_1029);
or U951 (N_951,In_1312,In_715);
xor U952 (N_952,In_1123,In_1287);
nand U953 (N_953,In_1317,In_198);
and U954 (N_954,In_1328,In_62);
xor U955 (N_955,In_1396,In_1108);
nand U956 (N_956,In_909,In_55);
xnor U957 (N_957,In_865,In_1464);
and U958 (N_958,In_1036,In_1065);
nand U959 (N_959,In_1180,In_415);
xnor U960 (N_960,In_1282,In_353);
nand U961 (N_961,In_499,In_862);
or U962 (N_962,In_403,In_944);
and U963 (N_963,In_912,In_882);
and U964 (N_964,In_1177,In_195);
or U965 (N_965,In_29,In_1236);
nor U966 (N_966,In_125,In_1333);
xnor U967 (N_967,In_1276,In_297);
nand U968 (N_968,In_1168,In_1452);
xnor U969 (N_969,In_1020,In_402);
nor U970 (N_970,In_1375,In_276);
nand U971 (N_971,In_271,In_803);
or U972 (N_972,In_1066,In_815);
or U973 (N_973,In_504,In_978);
xor U974 (N_974,In_902,In_114);
and U975 (N_975,In_911,In_368);
nor U976 (N_976,In_240,In_1048);
nand U977 (N_977,In_80,In_583);
and U978 (N_978,In_963,In_382);
xnor U979 (N_979,In_1462,In_1131);
xor U980 (N_980,In_937,In_843);
nand U981 (N_981,In_223,In_1108);
and U982 (N_982,In_1247,In_1477);
xor U983 (N_983,In_104,In_1091);
nand U984 (N_984,In_299,In_552);
nand U985 (N_985,In_846,In_860);
nor U986 (N_986,In_417,In_654);
nand U987 (N_987,In_193,In_1302);
xor U988 (N_988,In_571,In_1198);
or U989 (N_989,In_1065,In_778);
nor U990 (N_990,In_886,In_1226);
nand U991 (N_991,In_846,In_1419);
and U992 (N_992,In_574,In_456);
nand U993 (N_993,In_371,In_1048);
xnor U994 (N_994,In_637,In_822);
or U995 (N_995,In_597,In_655);
and U996 (N_996,In_187,In_235);
or U997 (N_997,In_389,In_868);
nor U998 (N_998,In_693,In_790);
and U999 (N_999,In_1326,In_94);
nor U1000 (N_1000,In_944,In_402);
xor U1001 (N_1001,In_620,In_1277);
xnor U1002 (N_1002,In_1324,In_979);
and U1003 (N_1003,In_1338,In_620);
nor U1004 (N_1004,In_81,In_262);
or U1005 (N_1005,In_1286,In_998);
and U1006 (N_1006,In_42,In_1358);
or U1007 (N_1007,In_310,In_405);
or U1008 (N_1008,In_1235,In_201);
nand U1009 (N_1009,In_874,In_10);
or U1010 (N_1010,In_1042,In_10);
or U1011 (N_1011,In_439,In_1026);
or U1012 (N_1012,In_493,In_881);
nor U1013 (N_1013,In_1243,In_502);
xnor U1014 (N_1014,In_159,In_1489);
or U1015 (N_1015,In_1297,In_1287);
nor U1016 (N_1016,In_403,In_1259);
and U1017 (N_1017,In_1296,In_320);
nand U1018 (N_1018,In_1103,In_823);
nand U1019 (N_1019,In_60,In_8);
nand U1020 (N_1020,In_1158,In_69);
nor U1021 (N_1021,In_583,In_1059);
or U1022 (N_1022,In_361,In_235);
and U1023 (N_1023,In_86,In_506);
or U1024 (N_1024,In_89,In_1461);
or U1025 (N_1025,In_323,In_267);
xor U1026 (N_1026,In_444,In_41);
nand U1027 (N_1027,In_683,In_486);
nor U1028 (N_1028,In_797,In_1113);
nor U1029 (N_1029,In_911,In_414);
nand U1030 (N_1030,In_1056,In_249);
and U1031 (N_1031,In_456,In_760);
nand U1032 (N_1032,In_1274,In_58);
nor U1033 (N_1033,In_540,In_322);
and U1034 (N_1034,In_229,In_718);
and U1035 (N_1035,In_1226,In_185);
xor U1036 (N_1036,In_1425,In_116);
and U1037 (N_1037,In_1033,In_324);
nor U1038 (N_1038,In_433,In_644);
and U1039 (N_1039,In_950,In_994);
and U1040 (N_1040,In_350,In_1008);
and U1041 (N_1041,In_1052,In_149);
nand U1042 (N_1042,In_1259,In_1296);
xor U1043 (N_1043,In_138,In_223);
or U1044 (N_1044,In_702,In_730);
nor U1045 (N_1045,In_164,In_1260);
nand U1046 (N_1046,In_147,In_32);
and U1047 (N_1047,In_1007,In_616);
and U1048 (N_1048,In_171,In_1021);
and U1049 (N_1049,In_973,In_354);
or U1050 (N_1050,In_74,In_1088);
xnor U1051 (N_1051,In_291,In_1101);
and U1052 (N_1052,In_696,In_170);
or U1053 (N_1053,In_236,In_1445);
and U1054 (N_1054,In_730,In_1296);
nor U1055 (N_1055,In_1275,In_1435);
and U1056 (N_1056,In_1075,In_35);
nand U1057 (N_1057,In_317,In_585);
and U1058 (N_1058,In_1177,In_125);
nand U1059 (N_1059,In_720,In_886);
or U1060 (N_1060,In_1041,In_1300);
and U1061 (N_1061,In_8,In_0);
xor U1062 (N_1062,In_615,In_995);
xnor U1063 (N_1063,In_667,In_705);
xor U1064 (N_1064,In_1118,In_983);
xnor U1065 (N_1065,In_416,In_1042);
nand U1066 (N_1066,In_83,In_158);
or U1067 (N_1067,In_91,In_972);
and U1068 (N_1068,In_683,In_787);
nand U1069 (N_1069,In_94,In_1384);
nor U1070 (N_1070,In_764,In_680);
xor U1071 (N_1071,In_855,In_1397);
or U1072 (N_1072,In_526,In_1301);
nor U1073 (N_1073,In_716,In_273);
nand U1074 (N_1074,In_733,In_818);
nor U1075 (N_1075,In_301,In_992);
nor U1076 (N_1076,In_1271,In_124);
or U1077 (N_1077,In_1279,In_132);
xor U1078 (N_1078,In_901,In_1030);
xnor U1079 (N_1079,In_1142,In_565);
nor U1080 (N_1080,In_15,In_777);
nand U1081 (N_1081,In_258,In_1274);
xnor U1082 (N_1082,In_449,In_1246);
nor U1083 (N_1083,In_816,In_711);
nand U1084 (N_1084,In_1254,In_68);
and U1085 (N_1085,In_917,In_685);
or U1086 (N_1086,In_24,In_252);
nor U1087 (N_1087,In_1028,In_689);
nand U1088 (N_1088,In_84,In_885);
xor U1089 (N_1089,In_763,In_1269);
and U1090 (N_1090,In_1010,In_56);
xnor U1091 (N_1091,In_524,In_401);
nor U1092 (N_1092,In_125,In_1166);
nor U1093 (N_1093,In_277,In_118);
and U1094 (N_1094,In_1112,In_1079);
nand U1095 (N_1095,In_1104,In_114);
and U1096 (N_1096,In_351,In_844);
or U1097 (N_1097,In_8,In_402);
nor U1098 (N_1098,In_747,In_381);
nand U1099 (N_1099,In_1222,In_648);
nand U1100 (N_1100,In_592,In_507);
nand U1101 (N_1101,In_1134,In_299);
and U1102 (N_1102,In_1477,In_799);
and U1103 (N_1103,In_1399,In_1364);
or U1104 (N_1104,In_784,In_1250);
or U1105 (N_1105,In_125,In_650);
nor U1106 (N_1106,In_502,In_268);
and U1107 (N_1107,In_652,In_160);
and U1108 (N_1108,In_1054,In_1488);
and U1109 (N_1109,In_93,In_251);
and U1110 (N_1110,In_1331,In_667);
and U1111 (N_1111,In_1377,In_271);
and U1112 (N_1112,In_1410,In_624);
xor U1113 (N_1113,In_866,In_1288);
xnor U1114 (N_1114,In_1420,In_666);
xor U1115 (N_1115,In_489,In_1389);
nor U1116 (N_1116,In_1039,In_218);
and U1117 (N_1117,In_1445,In_356);
or U1118 (N_1118,In_171,In_727);
or U1119 (N_1119,In_1365,In_1422);
nor U1120 (N_1120,In_612,In_1405);
nand U1121 (N_1121,In_1243,In_617);
nor U1122 (N_1122,In_1251,In_925);
xor U1123 (N_1123,In_1189,In_980);
nand U1124 (N_1124,In_1401,In_974);
or U1125 (N_1125,In_1347,In_1386);
and U1126 (N_1126,In_694,In_392);
and U1127 (N_1127,In_349,In_751);
or U1128 (N_1128,In_357,In_779);
and U1129 (N_1129,In_1357,In_429);
or U1130 (N_1130,In_1369,In_809);
nand U1131 (N_1131,In_1427,In_1293);
nor U1132 (N_1132,In_566,In_1330);
and U1133 (N_1133,In_388,In_589);
xnor U1134 (N_1134,In_877,In_543);
xnor U1135 (N_1135,In_584,In_152);
or U1136 (N_1136,In_86,In_678);
or U1137 (N_1137,In_953,In_734);
nand U1138 (N_1138,In_1424,In_729);
and U1139 (N_1139,In_1453,In_1448);
nand U1140 (N_1140,In_787,In_128);
xnor U1141 (N_1141,In_1416,In_1231);
nor U1142 (N_1142,In_417,In_1032);
and U1143 (N_1143,In_633,In_304);
nor U1144 (N_1144,In_988,In_345);
nand U1145 (N_1145,In_1188,In_914);
or U1146 (N_1146,In_986,In_205);
xor U1147 (N_1147,In_1242,In_1061);
and U1148 (N_1148,In_825,In_398);
or U1149 (N_1149,In_250,In_670);
or U1150 (N_1150,In_104,In_1186);
nor U1151 (N_1151,In_441,In_219);
xnor U1152 (N_1152,In_1052,In_1212);
xnor U1153 (N_1153,In_1010,In_339);
and U1154 (N_1154,In_1253,In_834);
nand U1155 (N_1155,In_1227,In_1256);
nand U1156 (N_1156,In_1452,In_490);
nand U1157 (N_1157,In_777,In_1105);
and U1158 (N_1158,In_579,In_702);
or U1159 (N_1159,In_480,In_949);
or U1160 (N_1160,In_34,In_1034);
or U1161 (N_1161,In_482,In_104);
xor U1162 (N_1162,In_1045,In_1030);
and U1163 (N_1163,In_214,In_379);
or U1164 (N_1164,In_180,In_338);
xnor U1165 (N_1165,In_81,In_1141);
or U1166 (N_1166,In_1318,In_495);
or U1167 (N_1167,In_843,In_835);
or U1168 (N_1168,In_1084,In_180);
or U1169 (N_1169,In_364,In_1365);
xor U1170 (N_1170,In_340,In_503);
nand U1171 (N_1171,In_119,In_69);
nand U1172 (N_1172,In_895,In_418);
xor U1173 (N_1173,In_1413,In_157);
xnor U1174 (N_1174,In_987,In_1291);
nor U1175 (N_1175,In_1455,In_654);
and U1176 (N_1176,In_246,In_475);
nand U1177 (N_1177,In_1223,In_173);
nand U1178 (N_1178,In_1114,In_1372);
nor U1179 (N_1179,In_830,In_1194);
and U1180 (N_1180,In_441,In_424);
and U1181 (N_1181,In_113,In_214);
nor U1182 (N_1182,In_124,In_293);
or U1183 (N_1183,In_827,In_577);
nor U1184 (N_1184,In_162,In_628);
and U1185 (N_1185,In_1287,In_1025);
nor U1186 (N_1186,In_684,In_1462);
xor U1187 (N_1187,In_1436,In_1340);
and U1188 (N_1188,In_932,In_1313);
nand U1189 (N_1189,In_1224,In_1087);
nor U1190 (N_1190,In_1401,In_1050);
nand U1191 (N_1191,In_182,In_553);
nand U1192 (N_1192,In_475,In_1017);
xnor U1193 (N_1193,In_1151,In_1274);
and U1194 (N_1194,In_528,In_526);
and U1195 (N_1195,In_1030,In_1118);
nor U1196 (N_1196,In_761,In_488);
xor U1197 (N_1197,In_1119,In_1421);
nand U1198 (N_1198,In_933,In_823);
xor U1199 (N_1199,In_590,In_749);
and U1200 (N_1200,In_38,In_451);
nor U1201 (N_1201,In_436,In_1346);
or U1202 (N_1202,In_332,In_100);
or U1203 (N_1203,In_1187,In_226);
and U1204 (N_1204,In_327,In_151);
nand U1205 (N_1205,In_1404,In_1066);
nor U1206 (N_1206,In_999,In_1312);
xnor U1207 (N_1207,In_1164,In_674);
xnor U1208 (N_1208,In_475,In_599);
and U1209 (N_1209,In_1193,In_1024);
nor U1210 (N_1210,In_1317,In_4);
nand U1211 (N_1211,In_735,In_445);
xnor U1212 (N_1212,In_776,In_1442);
and U1213 (N_1213,In_61,In_709);
and U1214 (N_1214,In_632,In_1456);
xor U1215 (N_1215,In_1222,In_867);
nand U1216 (N_1216,In_1068,In_206);
nor U1217 (N_1217,In_1082,In_974);
xor U1218 (N_1218,In_303,In_1148);
or U1219 (N_1219,In_779,In_453);
nand U1220 (N_1220,In_30,In_656);
or U1221 (N_1221,In_41,In_899);
and U1222 (N_1222,In_34,In_1398);
nand U1223 (N_1223,In_1366,In_517);
nand U1224 (N_1224,In_408,In_1485);
nand U1225 (N_1225,In_1003,In_451);
nor U1226 (N_1226,In_1405,In_856);
xor U1227 (N_1227,In_1220,In_1028);
or U1228 (N_1228,In_1214,In_785);
and U1229 (N_1229,In_1474,In_490);
xnor U1230 (N_1230,In_1235,In_1468);
and U1231 (N_1231,In_1380,In_1112);
xor U1232 (N_1232,In_235,In_1155);
or U1233 (N_1233,In_1162,In_379);
and U1234 (N_1234,In_67,In_457);
and U1235 (N_1235,In_1009,In_265);
xnor U1236 (N_1236,In_242,In_1068);
and U1237 (N_1237,In_1476,In_459);
nor U1238 (N_1238,In_675,In_690);
nor U1239 (N_1239,In_244,In_369);
xnor U1240 (N_1240,In_33,In_1235);
nor U1241 (N_1241,In_1463,In_913);
and U1242 (N_1242,In_343,In_733);
nor U1243 (N_1243,In_1463,In_1045);
or U1244 (N_1244,In_927,In_366);
nor U1245 (N_1245,In_1365,In_1041);
nor U1246 (N_1246,In_1419,In_135);
xnor U1247 (N_1247,In_1194,In_222);
xor U1248 (N_1248,In_318,In_1065);
xnor U1249 (N_1249,In_899,In_401);
and U1250 (N_1250,In_876,In_1312);
xnor U1251 (N_1251,In_624,In_852);
nand U1252 (N_1252,In_891,In_1371);
xnor U1253 (N_1253,In_820,In_257);
and U1254 (N_1254,In_226,In_1018);
nor U1255 (N_1255,In_904,In_1400);
or U1256 (N_1256,In_412,In_247);
and U1257 (N_1257,In_1017,In_858);
and U1258 (N_1258,In_1465,In_97);
nand U1259 (N_1259,In_622,In_1244);
nand U1260 (N_1260,In_1131,In_1235);
and U1261 (N_1261,In_148,In_170);
or U1262 (N_1262,In_262,In_358);
xnor U1263 (N_1263,In_171,In_476);
nand U1264 (N_1264,In_538,In_1007);
nand U1265 (N_1265,In_1244,In_1048);
nand U1266 (N_1266,In_1359,In_682);
nor U1267 (N_1267,In_356,In_1010);
or U1268 (N_1268,In_974,In_732);
nand U1269 (N_1269,In_1158,In_945);
xor U1270 (N_1270,In_1409,In_753);
and U1271 (N_1271,In_185,In_872);
or U1272 (N_1272,In_1058,In_1226);
xor U1273 (N_1273,In_287,In_846);
or U1274 (N_1274,In_1492,In_67);
xor U1275 (N_1275,In_734,In_1139);
nor U1276 (N_1276,In_396,In_618);
nand U1277 (N_1277,In_374,In_388);
and U1278 (N_1278,In_261,In_722);
or U1279 (N_1279,In_1306,In_300);
and U1280 (N_1280,In_911,In_539);
and U1281 (N_1281,In_1157,In_962);
xnor U1282 (N_1282,In_89,In_321);
nor U1283 (N_1283,In_817,In_144);
nor U1284 (N_1284,In_1474,In_592);
nor U1285 (N_1285,In_796,In_518);
and U1286 (N_1286,In_1303,In_122);
or U1287 (N_1287,In_282,In_302);
or U1288 (N_1288,In_1240,In_1390);
nand U1289 (N_1289,In_1479,In_1297);
xnor U1290 (N_1290,In_1386,In_33);
xor U1291 (N_1291,In_205,In_935);
or U1292 (N_1292,In_181,In_853);
xnor U1293 (N_1293,In_481,In_987);
and U1294 (N_1294,In_1327,In_1474);
xor U1295 (N_1295,In_544,In_1214);
xnor U1296 (N_1296,In_376,In_79);
nor U1297 (N_1297,In_380,In_1007);
nand U1298 (N_1298,In_685,In_62);
or U1299 (N_1299,In_545,In_1389);
xnor U1300 (N_1300,In_1473,In_1405);
xor U1301 (N_1301,In_1218,In_377);
xnor U1302 (N_1302,In_1055,In_1401);
and U1303 (N_1303,In_540,In_974);
and U1304 (N_1304,In_600,In_1012);
xor U1305 (N_1305,In_1400,In_430);
nand U1306 (N_1306,In_113,In_1096);
xor U1307 (N_1307,In_760,In_909);
nand U1308 (N_1308,In_1413,In_903);
nor U1309 (N_1309,In_261,In_300);
nor U1310 (N_1310,In_326,In_1322);
nand U1311 (N_1311,In_1468,In_1084);
xnor U1312 (N_1312,In_1255,In_1367);
or U1313 (N_1313,In_1222,In_608);
or U1314 (N_1314,In_799,In_37);
nand U1315 (N_1315,In_1352,In_633);
or U1316 (N_1316,In_898,In_1486);
or U1317 (N_1317,In_1112,In_380);
xnor U1318 (N_1318,In_354,In_530);
and U1319 (N_1319,In_654,In_1290);
and U1320 (N_1320,In_313,In_21);
nand U1321 (N_1321,In_624,In_310);
xnor U1322 (N_1322,In_955,In_412);
nor U1323 (N_1323,In_309,In_1166);
nor U1324 (N_1324,In_1332,In_1383);
nand U1325 (N_1325,In_419,In_30);
nand U1326 (N_1326,In_723,In_623);
and U1327 (N_1327,In_1111,In_1041);
nor U1328 (N_1328,In_61,In_90);
nor U1329 (N_1329,In_231,In_1482);
xnor U1330 (N_1330,In_724,In_942);
and U1331 (N_1331,In_1380,In_451);
nor U1332 (N_1332,In_1075,In_219);
xnor U1333 (N_1333,In_890,In_529);
xnor U1334 (N_1334,In_832,In_1125);
or U1335 (N_1335,In_1346,In_954);
nand U1336 (N_1336,In_728,In_239);
nor U1337 (N_1337,In_701,In_1437);
nor U1338 (N_1338,In_1314,In_1483);
nand U1339 (N_1339,In_1232,In_428);
nand U1340 (N_1340,In_674,In_5);
nand U1341 (N_1341,In_673,In_772);
and U1342 (N_1342,In_170,In_243);
nor U1343 (N_1343,In_530,In_535);
and U1344 (N_1344,In_511,In_1327);
or U1345 (N_1345,In_1328,In_815);
nor U1346 (N_1346,In_90,In_483);
and U1347 (N_1347,In_538,In_54);
or U1348 (N_1348,In_1127,In_268);
or U1349 (N_1349,In_1313,In_246);
nand U1350 (N_1350,In_766,In_490);
or U1351 (N_1351,In_1200,In_410);
and U1352 (N_1352,In_1157,In_885);
and U1353 (N_1353,In_250,In_302);
nand U1354 (N_1354,In_407,In_545);
nor U1355 (N_1355,In_195,In_840);
nor U1356 (N_1356,In_990,In_21);
nand U1357 (N_1357,In_1254,In_978);
nor U1358 (N_1358,In_231,In_465);
and U1359 (N_1359,In_636,In_557);
nand U1360 (N_1360,In_1267,In_839);
and U1361 (N_1361,In_1259,In_58);
and U1362 (N_1362,In_442,In_1365);
or U1363 (N_1363,In_216,In_1104);
nor U1364 (N_1364,In_1175,In_1351);
nor U1365 (N_1365,In_1289,In_1468);
or U1366 (N_1366,In_1353,In_1213);
nand U1367 (N_1367,In_1456,In_133);
nand U1368 (N_1368,In_738,In_77);
nor U1369 (N_1369,In_34,In_328);
nand U1370 (N_1370,In_214,In_513);
nand U1371 (N_1371,In_459,In_953);
nor U1372 (N_1372,In_830,In_862);
or U1373 (N_1373,In_105,In_336);
xor U1374 (N_1374,In_44,In_1370);
and U1375 (N_1375,In_651,In_426);
xor U1376 (N_1376,In_1462,In_835);
nand U1377 (N_1377,In_732,In_415);
or U1378 (N_1378,In_608,In_239);
xnor U1379 (N_1379,In_479,In_227);
or U1380 (N_1380,In_134,In_208);
and U1381 (N_1381,In_639,In_174);
xor U1382 (N_1382,In_1488,In_8);
xor U1383 (N_1383,In_124,In_13);
xor U1384 (N_1384,In_1448,In_1109);
and U1385 (N_1385,In_915,In_118);
xor U1386 (N_1386,In_114,In_1366);
nand U1387 (N_1387,In_1208,In_481);
or U1388 (N_1388,In_1122,In_1266);
nor U1389 (N_1389,In_716,In_1351);
and U1390 (N_1390,In_607,In_836);
xor U1391 (N_1391,In_15,In_587);
xor U1392 (N_1392,In_460,In_697);
nand U1393 (N_1393,In_1167,In_1038);
nand U1394 (N_1394,In_205,In_301);
nand U1395 (N_1395,In_1320,In_122);
nand U1396 (N_1396,In_305,In_179);
nand U1397 (N_1397,In_358,In_459);
nand U1398 (N_1398,In_49,In_796);
and U1399 (N_1399,In_122,In_1271);
nor U1400 (N_1400,In_265,In_1310);
or U1401 (N_1401,In_607,In_387);
nor U1402 (N_1402,In_222,In_1365);
and U1403 (N_1403,In_515,In_277);
and U1404 (N_1404,In_335,In_1364);
nand U1405 (N_1405,In_1366,In_953);
xnor U1406 (N_1406,In_900,In_168);
or U1407 (N_1407,In_1262,In_540);
and U1408 (N_1408,In_1083,In_1232);
or U1409 (N_1409,In_1277,In_1491);
nor U1410 (N_1410,In_187,In_1104);
or U1411 (N_1411,In_854,In_1211);
nand U1412 (N_1412,In_205,In_219);
nand U1413 (N_1413,In_1043,In_1416);
and U1414 (N_1414,In_1483,In_1206);
nand U1415 (N_1415,In_1183,In_1312);
or U1416 (N_1416,In_50,In_773);
nand U1417 (N_1417,In_1004,In_210);
or U1418 (N_1418,In_1118,In_738);
xor U1419 (N_1419,In_1250,In_592);
and U1420 (N_1420,In_423,In_1012);
or U1421 (N_1421,In_403,In_689);
xnor U1422 (N_1422,In_39,In_254);
nor U1423 (N_1423,In_1126,In_894);
nand U1424 (N_1424,In_1153,In_740);
and U1425 (N_1425,In_892,In_88);
or U1426 (N_1426,In_1268,In_810);
nand U1427 (N_1427,In_1438,In_701);
nand U1428 (N_1428,In_1441,In_755);
xor U1429 (N_1429,In_201,In_665);
nor U1430 (N_1430,In_1013,In_557);
or U1431 (N_1431,In_1464,In_359);
xor U1432 (N_1432,In_1078,In_1362);
xor U1433 (N_1433,In_214,In_1);
xnor U1434 (N_1434,In_297,In_56);
nor U1435 (N_1435,In_911,In_551);
xnor U1436 (N_1436,In_1406,In_362);
nand U1437 (N_1437,In_1329,In_1461);
nand U1438 (N_1438,In_1232,In_839);
nor U1439 (N_1439,In_12,In_673);
nor U1440 (N_1440,In_1302,In_478);
and U1441 (N_1441,In_164,In_293);
or U1442 (N_1442,In_910,In_1041);
nand U1443 (N_1443,In_1453,In_139);
and U1444 (N_1444,In_1255,In_852);
nor U1445 (N_1445,In_640,In_1126);
nand U1446 (N_1446,In_1380,In_259);
nor U1447 (N_1447,In_628,In_1226);
and U1448 (N_1448,In_674,In_928);
nor U1449 (N_1449,In_530,In_1193);
nor U1450 (N_1450,In_1092,In_1214);
xor U1451 (N_1451,In_1103,In_339);
and U1452 (N_1452,In_191,In_467);
or U1453 (N_1453,In_919,In_121);
nand U1454 (N_1454,In_1118,In_1111);
or U1455 (N_1455,In_756,In_1486);
xor U1456 (N_1456,In_443,In_678);
or U1457 (N_1457,In_972,In_877);
nand U1458 (N_1458,In_126,In_72);
and U1459 (N_1459,In_56,In_1035);
and U1460 (N_1460,In_615,In_8);
and U1461 (N_1461,In_1329,In_1420);
and U1462 (N_1462,In_201,In_380);
nand U1463 (N_1463,In_19,In_1289);
and U1464 (N_1464,In_1030,In_1178);
and U1465 (N_1465,In_919,In_723);
nor U1466 (N_1466,In_137,In_932);
nor U1467 (N_1467,In_657,In_655);
nand U1468 (N_1468,In_82,In_21);
xor U1469 (N_1469,In_112,In_1157);
or U1470 (N_1470,In_244,In_104);
and U1471 (N_1471,In_754,In_525);
or U1472 (N_1472,In_260,In_757);
nand U1473 (N_1473,In_1237,In_512);
and U1474 (N_1474,In_1093,In_9);
nand U1475 (N_1475,In_315,In_1068);
or U1476 (N_1476,In_1323,In_210);
or U1477 (N_1477,In_1115,In_1090);
nand U1478 (N_1478,In_455,In_1381);
nor U1479 (N_1479,In_646,In_683);
nand U1480 (N_1480,In_98,In_267);
nand U1481 (N_1481,In_236,In_596);
nand U1482 (N_1482,In_962,In_1273);
nand U1483 (N_1483,In_1460,In_394);
nor U1484 (N_1484,In_487,In_32);
nand U1485 (N_1485,In_655,In_1276);
or U1486 (N_1486,In_770,In_748);
nand U1487 (N_1487,In_1384,In_560);
nand U1488 (N_1488,In_326,In_1338);
nand U1489 (N_1489,In_1324,In_670);
and U1490 (N_1490,In_476,In_1133);
or U1491 (N_1491,In_740,In_1484);
nand U1492 (N_1492,In_442,In_708);
nor U1493 (N_1493,In_185,In_1339);
nor U1494 (N_1494,In_1419,In_1312);
or U1495 (N_1495,In_1177,In_795);
nor U1496 (N_1496,In_1295,In_268);
and U1497 (N_1497,In_1318,In_698);
or U1498 (N_1498,In_859,In_565);
xor U1499 (N_1499,In_700,In_362);
nor U1500 (N_1500,N_956,N_698);
and U1501 (N_1501,N_33,N_658);
and U1502 (N_1502,N_1209,N_1348);
nand U1503 (N_1503,N_935,N_877);
or U1504 (N_1504,N_1440,N_1396);
nor U1505 (N_1505,N_189,N_918);
nor U1506 (N_1506,N_899,N_1311);
nor U1507 (N_1507,N_1373,N_586);
and U1508 (N_1508,N_1285,N_852);
xnor U1509 (N_1509,N_591,N_1393);
nand U1510 (N_1510,N_1456,N_1163);
nand U1511 (N_1511,N_1107,N_349);
nor U1512 (N_1512,N_914,N_421);
nand U1513 (N_1513,N_1310,N_835);
nor U1514 (N_1514,N_1319,N_1390);
nand U1515 (N_1515,N_1087,N_1450);
nor U1516 (N_1516,N_729,N_197);
xor U1517 (N_1517,N_293,N_505);
nand U1518 (N_1518,N_926,N_923);
xor U1519 (N_1519,N_406,N_358);
or U1520 (N_1520,N_364,N_432);
nand U1521 (N_1521,N_982,N_1183);
xor U1522 (N_1522,N_1244,N_1300);
nor U1523 (N_1523,N_760,N_342);
nand U1524 (N_1524,N_1382,N_776);
nor U1525 (N_1525,N_1427,N_920);
or U1526 (N_1526,N_670,N_1239);
xnor U1527 (N_1527,N_105,N_1108);
xnor U1528 (N_1528,N_1461,N_1082);
nor U1529 (N_1529,N_575,N_592);
nor U1530 (N_1530,N_225,N_773);
nand U1531 (N_1531,N_114,N_113);
and U1532 (N_1532,N_1193,N_182);
nand U1533 (N_1533,N_1229,N_929);
and U1534 (N_1534,N_1175,N_1271);
nor U1535 (N_1535,N_1179,N_649);
nand U1536 (N_1536,N_1474,N_1477);
or U1537 (N_1537,N_141,N_266);
or U1538 (N_1538,N_453,N_1353);
xor U1539 (N_1539,N_73,N_862);
nand U1540 (N_1540,N_854,N_904);
nor U1541 (N_1541,N_234,N_48);
nor U1542 (N_1542,N_507,N_617);
nor U1543 (N_1543,N_526,N_1492);
nor U1544 (N_1544,N_1488,N_1008);
xnor U1545 (N_1545,N_41,N_129);
nand U1546 (N_1546,N_177,N_1035);
nor U1547 (N_1547,N_1443,N_513);
nand U1548 (N_1548,N_111,N_101);
or U1549 (N_1549,N_993,N_715);
or U1550 (N_1550,N_790,N_91);
nor U1551 (N_1551,N_1439,N_1070);
nand U1552 (N_1552,N_395,N_337);
or U1553 (N_1553,N_1326,N_539);
or U1554 (N_1554,N_860,N_520);
or U1555 (N_1555,N_1255,N_825);
nand U1556 (N_1556,N_1418,N_352);
xnor U1557 (N_1557,N_420,N_1421);
xor U1558 (N_1558,N_1487,N_1288);
nor U1559 (N_1559,N_613,N_1429);
and U1560 (N_1560,N_861,N_538);
nand U1561 (N_1561,N_147,N_878);
and U1562 (N_1562,N_599,N_456);
nor U1563 (N_1563,N_1242,N_1369);
or U1564 (N_1564,N_208,N_374);
xnor U1565 (N_1565,N_1227,N_1270);
xor U1566 (N_1566,N_487,N_36);
and U1567 (N_1567,N_1030,N_1134);
and U1568 (N_1568,N_655,N_145);
nand U1569 (N_1569,N_1447,N_1187);
and U1570 (N_1570,N_801,N_221);
nand U1571 (N_1571,N_69,N_960);
nor U1572 (N_1572,N_277,N_754);
or U1573 (N_1573,N_438,N_531);
xor U1574 (N_1574,N_637,N_1406);
or U1575 (N_1575,N_786,N_204);
xnor U1576 (N_1576,N_271,N_517);
xor U1577 (N_1577,N_1394,N_881);
and U1578 (N_1578,N_572,N_131);
or U1579 (N_1579,N_1281,N_370);
xnor U1580 (N_1580,N_1092,N_143);
or U1581 (N_1581,N_85,N_598);
xnor U1582 (N_1582,N_1269,N_594);
or U1583 (N_1583,N_1056,N_2);
or U1584 (N_1584,N_1385,N_1071);
nor U1585 (N_1585,N_1036,N_390);
xnor U1586 (N_1586,N_1253,N_1233);
xor U1587 (N_1587,N_466,N_905);
nand U1588 (N_1588,N_1155,N_723);
nand U1589 (N_1589,N_1045,N_1061);
nand U1590 (N_1590,N_1391,N_725);
or U1591 (N_1591,N_396,N_672);
nand U1592 (N_1592,N_1132,N_693);
nand U1593 (N_1593,N_200,N_40);
or U1594 (N_1594,N_1408,N_1445);
xor U1595 (N_1595,N_1154,N_311);
xnor U1596 (N_1596,N_152,N_1400);
nor U1597 (N_1597,N_694,N_1121);
nand U1598 (N_1598,N_983,N_56);
or U1599 (N_1599,N_1162,N_787);
xnor U1600 (N_1600,N_726,N_172);
nor U1601 (N_1601,N_1338,N_407);
and U1602 (N_1602,N_1117,N_44);
xnor U1603 (N_1603,N_14,N_79);
and U1604 (N_1604,N_940,N_659);
and U1605 (N_1605,N_1014,N_31);
and U1606 (N_1606,N_377,N_1322);
and U1607 (N_1607,N_485,N_46);
xor U1608 (N_1608,N_344,N_621);
xnor U1609 (N_1609,N_1276,N_1012);
or U1610 (N_1610,N_537,N_889);
or U1611 (N_1611,N_921,N_232);
or U1612 (N_1612,N_302,N_669);
nand U1613 (N_1613,N_890,N_671);
xor U1614 (N_1614,N_979,N_448);
nor U1615 (N_1615,N_124,N_1282);
and U1616 (N_1616,N_455,N_1411);
nor U1617 (N_1617,N_1223,N_560);
nor U1618 (N_1618,N_1279,N_950);
xnor U1619 (N_1619,N_30,N_1342);
and U1620 (N_1620,N_1169,N_1113);
and U1621 (N_1621,N_345,N_1063);
or U1622 (N_1622,N_1368,N_1325);
xnor U1623 (N_1623,N_1225,N_1431);
or U1624 (N_1624,N_25,N_704);
nand U1625 (N_1625,N_508,N_1389);
xnor U1626 (N_1626,N_1435,N_1337);
xor U1627 (N_1627,N_902,N_199);
xnor U1628 (N_1628,N_267,N_112);
xor U1629 (N_1629,N_815,N_1031);
nand U1630 (N_1630,N_567,N_1318);
nand U1631 (N_1631,N_1160,N_27);
or U1632 (N_1632,N_361,N_436);
and U1633 (N_1633,N_70,N_238);
and U1634 (N_1634,N_948,N_84);
nor U1635 (N_1635,N_509,N_1251);
and U1636 (N_1636,N_896,N_994);
or U1637 (N_1637,N_439,N_1123);
nor U1638 (N_1638,N_1438,N_134);
and U1639 (N_1639,N_807,N_761);
nor U1640 (N_1640,N_156,N_1415);
nor U1641 (N_1641,N_435,N_1375);
and U1642 (N_1642,N_660,N_589);
xor U1643 (N_1643,N_1230,N_176);
xor U1644 (N_1644,N_445,N_632);
xnor U1645 (N_1645,N_75,N_876);
nand U1646 (N_1646,N_1360,N_908);
nor U1647 (N_1647,N_774,N_151);
nand U1648 (N_1648,N_148,N_1497);
nand U1649 (N_1649,N_1339,N_568);
xnor U1650 (N_1650,N_251,N_405);
nand U1651 (N_1651,N_169,N_366);
and U1652 (N_1652,N_1138,N_997);
or U1653 (N_1653,N_664,N_240);
nand U1654 (N_1654,N_12,N_1034);
nand U1655 (N_1655,N_387,N_1432);
nand U1656 (N_1656,N_365,N_1041);
nor U1657 (N_1657,N_388,N_892);
nand U1658 (N_1658,N_392,N_719);
or U1659 (N_1659,N_759,N_429);
or U1660 (N_1660,N_1424,N_1218);
or U1661 (N_1661,N_1470,N_161);
and U1662 (N_1662,N_1297,N_1228);
and U1663 (N_1663,N_356,N_223);
and U1664 (N_1664,N_1452,N_1266);
or U1665 (N_1665,N_1054,N_1211);
and U1666 (N_1666,N_1112,N_848);
and U1667 (N_1667,N_1430,N_510);
and U1668 (N_1668,N_1114,N_1142);
or U1669 (N_1669,N_1321,N_1192);
and U1670 (N_1670,N_934,N_300);
nor U1671 (N_1671,N_1202,N_498);
and U1672 (N_1672,N_1245,N_357);
or U1673 (N_1673,N_532,N_1130);
nor U1674 (N_1674,N_931,N_393);
nand U1675 (N_1675,N_433,N_243);
nor U1676 (N_1676,N_434,N_990);
nor U1677 (N_1677,N_967,N_314);
nor U1678 (N_1678,N_891,N_1298);
nor U1679 (N_1679,N_823,N_491);
or U1680 (N_1680,N_400,N_813);
xnor U1681 (N_1681,N_335,N_1366);
nand U1682 (N_1682,N_951,N_62);
and U1683 (N_1683,N_77,N_551);
and U1684 (N_1684,N_1309,N_292);
and U1685 (N_1685,N_1324,N_468);
or U1686 (N_1686,N_995,N_1290);
or U1687 (N_1687,N_628,N_1482);
or U1688 (N_1688,N_409,N_1124);
nor U1689 (N_1689,N_654,N_1143);
nand U1690 (N_1690,N_1139,N_603);
xnor U1691 (N_1691,N_1101,N_484);
nor U1692 (N_1692,N_1205,N_1009);
xor U1693 (N_1693,N_925,N_1062);
and U1694 (N_1694,N_1267,N_1473);
nand U1695 (N_1695,N_987,N_697);
and U1696 (N_1696,N_705,N_958);
nand U1697 (N_1697,N_1350,N_1081);
or U1698 (N_1698,N_95,N_536);
and U1699 (N_1699,N_268,N_1174);
nor U1700 (N_1700,N_886,N_796);
and U1701 (N_1701,N_461,N_457);
nand U1702 (N_1702,N_196,N_847);
nor U1703 (N_1703,N_126,N_241);
xnor U1704 (N_1704,N_945,N_1098);
and U1705 (N_1705,N_408,N_108);
nor U1706 (N_1706,N_1133,N_888);
nand U1707 (N_1707,N_578,N_78);
and U1708 (N_1708,N_1096,N_584);
or U1709 (N_1709,N_136,N_245);
and U1710 (N_1710,N_566,N_1404);
nand U1711 (N_1711,N_724,N_735);
and U1712 (N_1712,N_690,N_884);
xor U1713 (N_1713,N_362,N_619);
and U1714 (N_1714,N_313,N_936);
and U1715 (N_1715,N_820,N_389);
and U1716 (N_1716,N_858,N_1469);
and U1717 (N_1717,N_946,N_1040);
or U1718 (N_1718,N_1046,N_1414);
or U1719 (N_1719,N_810,N_1475);
or U1720 (N_1720,N_18,N_1257);
or U1721 (N_1721,N_215,N_1376);
or U1722 (N_1722,N_1278,N_1097);
or U1723 (N_1723,N_1131,N_1027);
nor U1724 (N_1724,N_29,N_702);
xnor U1725 (N_1725,N_1274,N_919);
and U1726 (N_1726,N_1259,N_316);
nor U1727 (N_1727,N_1115,N_700);
and U1728 (N_1728,N_306,N_175);
nand U1729 (N_1729,N_1434,N_51);
xor U1730 (N_1730,N_373,N_515);
nor U1731 (N_1731,N_7,N_677);
nand U1732 (N_1732,N_116,N_679);
or U1733 (N_1733,N_359,N_764);
xor U1734 (N_1734,N_100,N_250);
nor U1735 (N_1735,N_618,N_1095);
nor U1736 (N_1736,N_88,N_473);
or U1737 (N_1737,N_418,N_1345);
or U1738 (N_1738,N_804,N_558);
nand U1739 (N_1739,N_587,N_699);
xnor U1740 (N_1740,N_1146,N_678);
or U1741 (N_1741,N_1305,N_795);
or U1742 (N_1742,N_989,N_280);
and U1743 (N_1743,N_1044,N_5);
nand U1744 (N_1744,N_1494,N_1178);
xnor U1745 (N_1745,N_1005,N_1196);
nand U1746 (N_1746,N_486,N_1354);
nor U1747 (N_1747,N_283,N_1362);
nor U1748 (N_1748,N_1053,N_1197);
or U1749 (N_1749,N_1216,N_1145);
and U1750 (N_1750,N_47,N_720);
xnor U1751 (N_1751,N_262,N_290);
nand U1752 (N_1752,N_684,N_185);
nand U1753 (N_1753,N_673,N_440);
or U1754 (N_1754,N_949,N_1377);
nor U1755 (N_1755,N_533,N_834);
or U1756 (N_1756,N_287,N_742);
xnor U1757 (N_1757,N_1428,N_163);
or U1758 (N_1758,N_1120,N_1294);
or U1759 (N_1759,N_1306,N_228);
nor U1760 (N_1760,N_135,N_981);
and U1761 (N_1761,N_1363,N_8);
and U1762 (N_1762,N_1011,N_1176);
nor U1763 (N_1763,N_713,N_1454);
xor U1764 (N_1764,N_569,N_635);
or U1765 (N_1765,N_733,N_178);
or U1766 (N_1766,N_1472,N_310);
nor U1767 (N_1767,N_231,N_1261);
nor U1768 (N_1768,N_816,N_717);
nor U1769 (N_1769,N_331,N_1457);
and U1770 (N_1770,N_1484,N_264);
nor U1771 (N_1771,N_1080,N_631);
nand U1772 (N_1772,N_401,N_552);
and U1773 (N_1773,N_1222,N_1365);
nand U1774 (N_1774,N_992,N_1103);
nand U1775 (N_1775,N_1003,N_442);
and U1776 (N_1776,N_588,N_523);
or U1777 (N_1777,N_504,N_608);
and U1778 (N_1778,N_1453,N_38);
xnor U1779 (N_1779,N_1280,N_644);
or U1780 (N_1780,N_840,N_1328);
xor U1781 (N_1781,N_346,N_755);
nand U1782 (N_1782,N_893,N_850);
and U1783 (N_1783,N_276,N_246);
nand U1784 (N_1784,N_1180,N_739);
nor U1785 (N_1785,N_1313,N_695);
or U1786 (N_1786,N_86,N_996);
and U1787 (N_1787,N_666,N_668);
nand U1788 (N_1788,N_963,N_194);
and U1789 (N_1789,N_559,N_218);
nor U1790 (N_1790,N_593,N_210);
nand U1791 (N_1791,N_601,N_917);
and U1792 (N_1792,N_187,N_1398);
or U1793 (N_1793,N_322,N_1307);
and U1794 (N_1794,N_1020,N_752);
nand U1795 (N_1795,N_939,N_90);
nor U1796 (N_1796,N_880,N_1073);
and U1797 (N_1797,N_1479,N_160);
or U1798 (N_1798,N_1286,N_428);
or U1799 (N_1799,N_502,N_158);
and U1800 (N_1800,N_64,N_355);
xnor U1801 (N_1801,N_585,N_417);
nor U1802 (N_1802,N_1182,N_610);
or U1803 (N_1803,N_506,N_1093);
and U1804 (N_1804,N_495,N_1077);
nor U1805 (N_1805,N_959,N_1249);
nor U1806 (N_1806,N_63,N_696);
nand U1807 (N_1807,N_897,N_1);
nand U1808 (N_1808,N_1372,N_1153);
nor U1809 (N_1809,N_159,N_192);
nor U1810 (N_1810,N_125,N_636);
nor U1811 (N_1811,N_1426,N_1204);
and U1812 (N_1812,N_765,N_1171);
xnor U1813 (N_1813,N_1068,N_1268);
nor U1814 (N_1814,N_579,N_872);
and U1815 (N_1815,N_132,N_595);
or U1816 (N_1816,N_1442,N_818);
nor U1817 (N_1817,N_916,N_330);
nor U1818 (N_1818,N_1361,N_437);
nor U1819 (N_1819,N_778,N_34);
nor U1820 (N_1820,N_550,N_379);
nor U1821 (N_1821,N_146,N_667);
nor U1822 (N_1822,N_371,N_1149);
or U1823 (N_1823,N_1015,N_710);
xnor U1824 (N_1824,N_216,N_827);
nand U1825 (N_1825,N_273,N_309);
nand U1826 (N_1826,N_315,N_22);
or U1827 (N_1827,N_1055,N_519);
and U1828 (N_1828,N_912,N_770);
nand U1829 (N_1829,N_1224,N_1065);
and U1830 (N_1830,N_831,N_1240);
and U1831 (N_1831,N_122,N_806);
nand U1832 (N_1832,N_333,N_783);
and U1833 (N_1833,N_746,N_201);
nor U1834 (N_1834,N_328,N_811);
nor U1835 (N_1835,N_350,N_1207);
xnor U1836 (N_1836,N_757,N_573);
and U1837 (N_1837,N_730,N_625);
xor U1838 (N_1838,N_1156,N_1386);
nor U1839 (N_1839,N_1191,N_492);
xor U1840 (N_1840,N_42,N_1147);
or U1841 (N_1841,N_450,N_184);
nor U1842 (N_1842,N_1201,N_1302);
or U1843 (N_1843,N_985,N_846);
and U1844 (N_1844,N_270,N_446);
xnor U1845 (N_1845,N_1275,N_65);
or U1846 (N_1846,N_142,N_867);
and U1847 (N_1847,N_419,N_797);
or U1848 (N_1848,N_1258,N_477);
xnor U1849 (N_1849,N_173,N_590);
nand U1850 (N_1850,N_999,N_525);
or U1851 (N_1851,N_1448,N_1116);
xnor U1852 (N_1852,N_954,N_235);
nand U1853 (N_1853,N_1181,N_383);
xnor U1854 (N_1854,N_1140,N_839);
or U1855 (N_1855,N_381,N_1273);
or U1856 (N_1856,N_728,N_883);
xnor U1857 (N_1857,N_565,N_1059);
or U1858 (N_1858,N_616,N_1118);
or U1859 (N_1859,N_1330,N_1425);
nand U1860 (N_1860,N_829,N_1066);
and U1861 (N_1861,N_1122,N_736);
nor U1862 (N_1862,N_1496,N_1157);
nand U1863 (N_1863,N_866,N_53);
nor U1864 (N_1864,N_1481,N_1141);
nand U1865 (N_1865,N_1247,N_1293);
nand U1866 (N_1866,N_641,N_1329);
or U1867 (N_1867,N_853,N_812);
nand U1868 (N_1868,N_67,N_303);
nand U1869 (N_1869,N_743,N_1170);
and U1870 (N_1870,N_582,N_1126);
xor U1871 (N_1871,N_869,N_363);
nor U1872 (N_1872,N_1190,N_441);
xor U1873 (N_1873,N_794,N_288);
nand U1874 (N_1874,N_1371,N_1332);
or U1875 (N_1875,N_991,N_895);
nor U1876 (N_1876,N_727,N_943);
nand U1877 (N_1877,N_545,N_222);
or U1878 (N_1878,N_1079,N_685);
nand U1879 (N_1879,N_256,N_1189);
and U1880 (N_1880,N_416,N_646);
xnor U1881 (N_1881,N_263,N_427);
xnor U1882 (N_1882,N_1083,N_59);
or U1883 (N_1883,N_1076,N_43);
xor U1884 (N_1884,N_229,N_1099);
or U1885 (N_1885,N_885,N_1359);
or U1886 (N_1886,N_324,N_443);
and U1887 (N_1887,N_179,N_879);
nand U1888 (N_1888,N_1048,N_50);
or U1889 (N_1889,N_398,N_581);
and U1890 (N_1890,N_535,N_1219);
and U1891 (N_1891,N_1001,N_255);
xnor U1892 (N_1892,N_482,N_875);
or U1893 (N_1893,N_1004,N_1032);
or U1894 (N_1894,N_932,N_1084);
xor U1895 (N_1895,N_556,N_788);
xor U1896 (N_1896,N_1463,N_107);
or U1897 (N_1897,N_154,N_771);
nand U1898 (N_1898,N_777,N_252);
nor U1899 (N_1899,N_1416,N_1033);
nor U1900 (N_1900,N_832,N_460);
or U1901 (N_1901,N_1347,N_1422);
and U1902 (N_1902,N_580,N_411);
nor U1903 (N_1903,N_476,N_630);
or U1904 (N_1904,N_1026,N_609);
nand U1905 (N_1905,N_612,N_496);
nand U1906 (N_1906,N_785,N_1395);
nand U1907 (N_1907,N_549,N_737);
nand U1908 (N_1908,N_109,N_97);
or U1909 (N_1909,N_745,N_195);
nor U1910 (N_1910,N_574,N_213);
nor U1911 (N_1911,N_425,N_1106);
xor U1912 (N_1912,N_412,N_464);
and U1913 (N_1913,N_657,N_947);
and U1914 (N_1914,N_296,N_89);
and U1915 (N_1915,N_23,N_1308);
and U1916 (N_1916,N_563,N_348);
and U1917 (N_1917,N_808,N_965);
xnor U1918 (N_1918,N_817,N_650);
xor U1919 (N_1919,N_170,N_928);
nor U1920 (N_1920,N_843,N_499);
xor U1921 (N_1921,N_1254,N_244);
nor U1922 (N_1922,N_1444,N_1127);
and U1923 (N_1923,N_1017,N_1128);
nor U1924 (N_1924,N_1291,N_938);
nand U1925 (N_1925,N_712,N_611);
nor U1926 (N_1926,N_680,N_369);
nand U1927 (N_1927,N_894,N_92);
nor U1928 (N_1928,N_211,N_226);
nand U1929 (N_1929,N_826,N_756);
and U1930 (N_1930,N_561,N_749);
xnor U1931 (N_1931,N_127,N_1064);
xnor U1932 (N_1932,N_318,N_72);
or U1933 (N_1933,N_207,N_500);
or U1934 (N_1934,N_55,N_1407);
nor U1935 (N_1935,N_1417,N_741);
xor U1936 (N_1936,N_71,N_1016);
nand U1937 (N_1937,N_1025,N_740);
or U1938 (N_1938,N_451,N_171);
or U1939 (N_1939,N_326,N_1057);
xnor U1940 (N_1940,N_1217,N_1344);
nor U1941 (N_1941,N_1480,N_1058);
nor U1942 (N_1942,N_553,N_115);
nor U1943 (N_1943,N_304,N_1090);
xor U1944 (N_1944,N_1029,N_530);
and U1945 (N_1945,N_721,N_110);
nand U1946 (N_1946,N_1349,N_254);
nor U1947 (N_1947,N_909,N_1383);
xnor U1948 (N_1948,N_528,N_518);
and U1949 (N_1949,N_868,N_1265);
xor U1950 (N_1950,N_769,N_1413);
xor U1951 (N_1951,N_286,N_1185);
or U1952 (N_1952,N_1334,N_1381);
nor U1953 (N_1953,N_351,N_1161);
xor U1954 (N_1954,N_144,N_1210);
nor U1955 (N_1955,N_970,N_1323);
xnor U1956 (N_1956,N_384,N_782);
and U1957 (N_1957,N_793,N_1088);
and U1958 (N_1958,N_953,N_1264);
nor U1959 (N_1959,N_360,N_842);
and U1960 (N_1960,N_661,N_1314);
and U1961 (N_1961,N_962,N_763);
nand U1962 (N_1962,N_157,N_340);
and U1963 (N_1963,N_291,N_620);
or U1964 (N_1964,N_1006,N_1167);
nand U1965 (N_1965,N_1295,N_738);
or U1966 (N_1966,N_1260,N_1110);
nand U1967 (N_1967,N_1412,N_856);
and U1968 (N_1968,N_798,N_527);
nand U1969 (N_1969,N_0,N_1214);
nand U1970 (N_1970,N_480,N_955);
or U1971 (N_1971,N_423,N_1013);
or U1972 (N_1972,N_233,N_767);
or U1973 (N_1973,N_404,N_82);
xor U1974 (N_1974,N_1405,N_859);
xnor U1975 (N_1975,N_1485,N_230);
and U1976 (N_1976,N_103,N_1246);
nand U1977 (N_1977,N_1464,N_426);
nor U1978 (N_1978,N_924,N_39);
xnor U1979 (N_1979,N_541,N_1403);
and U1980 (N_1980,N_49,N_751);
and U1981 (N_1981,N_4,N_1067);
and U1982 (N_1982,N_343,N_653);
and U1983 (N_1983,N_833,N_1441);
or U1984 (N_1984,N_489,N_472);
and U1985 (N_1985,N_915,N_516);
nor U1986 (N_1986,N_220,N_863);
nand U1987 (N_1987,N_1490,N_647);
nor U1988 (N_1988,N_494,N_120);
or U1989 (N_1989,N_1198,N_471);
nand U1990 (N_1990,N_1150,N_968);
xor U1991 (N_1991,N_284,N_139);
and U1992 (N_1992,N_174,N_1378);
xor U1993 (N_1993,N_855,N_583);
xnor U1994 (N_1994,N_307,N_781);
and U1995 (N_1995,N_155,N_1256);
and U1996 (N_1996,N_957,N_372);
and U1997 (N_1997,N_805,N_1331);
nand U1998 (N_1998,N_544,N_1236);
nand U1999 (N_1999,N_984,N_87);
nor U2000 (N_2000,N_1272,N_775);
nand U2001 (N_2001,N_1397,N_1007);
or U2002 (N_2002,N_903,N_214);
xnor U2003 (N_2003,N_629,N_1213);
or U2004 (N_2004,N_1215,N_714);
nand U2005 (N_2005,N_60,N_1250);
or U2006 (N_2006,N_399,N_910);
and U2007 (N_2007,N_1235,N_1460);
nor U2008 (N_2008,N_153,N_164);
and U2009 (N_2009,N_639,N_627);
xnor U2010 (N_2010,N_289,N_140);
nor U2011 (N_2011,N_998,N_422);
or U2012 (N_2012,N_253,N_841);
and U2013 (N_2013,N_1462,N_534);
nand U2014 (N_2014,N_665,N_138);
nor U2015 (N_2015,N_1320,N_922);
or U2016 (N_2016,N_298,N_1410);
nand U2017 (N_2017,N_341,N_1458);
or U2018 (N_2018,N_260,N_317);
or U2019 (N_2019,N_701,N_378);
or U2020 (N_2020,N_864,N_1125);
xor U2021 (N_2021,N_1491,N_941);
nor U2022 (N_2022,N_1263,N_332);
nand U2023 (N_2023,N_488,N_319);
or U2024 (N_2024,N_54,N_1471);
nand U2025 (N_2025,N_278,N_236);
nor U2026 (N_2026,N_548,N_16);
xnor U2027 (N_2027,N_614,N_975);
and U2028 (N_2028,N_1042,N_424);
xnor U2029 (N_2029,N_1296,N_716);
xor U2030 (N_2030,N_1148,N_543);
or U2031 (N_2031,N_966,N_1238);
nand U2032 (N_2032,N_339,N_104);
or U2033 (N_2033,N_604,N_606);
nor U2034 (N_2034,N_1287,N_1078);
and U2035 (N_2035,N_1104,N_198);
nand U2036 (N_2036,N_600,N_1144);
and U2037 (N_2037,N_96,N_822);
nand U2038 (N_2038,N_1340,N_1437);
xnor U2039 (N_2039,N_607,N_1237);
and U2040 (N_2040,N_1241,N_837);
nor U2041 (N_2041,N_479,N_1039);
xnor U2042 (N_2042,N_809,N_465);
and U2043 (N_2043,N_933,N_206);
nand U2044 (N_2044,N_708,N_675);
nand U2045 (N_2045,N_1177,N_1050);
xor U2046 (N_2046,N_15,N_1168);
and U2047 (N_2047,N_217,N_1399);
nand U2048 (N_2048,N_988,N_663);
nand U2049 (N_2049,N_643,N_547);
nand U2050 (N_2050,N_1493,N_301);
or U2051 (N_2051,N_571,N_1102);
or U2052 (N_2052,N_1446,N_1166);
xor U2053 (N_2053,N_1423,N_753);
or U2054 (N_2054,N_784,N_626);
or U2055 (N_2055,N_58,N_83);
xor U2056 (N_2056,N_380,N_542);
and U2057 (N_2057,N_119,N_37);
nor U2058 (N_2058,N_1208,N_942);
or U2059 (N_2059,N_1129,N_166);
or U2060 (N_2060,N_676,N_1449);
or U2061 (N_2061,N_265,N_1387);
xor U2062 (N_2062,N_961,N_927);
nor U2063 (N_2063,N_1333,N_475);
xnor U2064 (N_2064,N_193,N_281);
nand U2065 (N_2065,N_258,N_98);
nor U2066 (N_2066,N_431,N_454);
nor U2067 (N_2067,N_1234,N_1364);
and U2068 (N_2068,N_106,N_368);
or U2069 (N_2069,N_824,N_282);
nor U2070 (N_2070,N_1220,N_849);
or U2071 (N_2071,N_1024,N_493);
or U2072 (N_2072,N_467,N_1038);
nor U2073 (N_2073,N_972,N_1047);
and U2074 (N_2074,N_602,N_239);
or U2075 (N_2075,N_779,N_376);
or U2076 (N_2076,N_687,N_353);
and U2077 (N_2077,N_622,N_978);
xnor U2078 (N_2078,N_52,N_944);
nand U2079 (N_2079,N_1151,N_205);
and U2080 (N_2080,N_1135,N_681);
nor U2081 (N_2081,N_1074,N_80);
or U2082 (N_2082,N_1119,N_1010);
nor U2083 (N_2083,N_68,N_1303);
and U2084 (N_2084,N_74,N_1352);
nand U2085 (N_2085,N_1409,N_873);
or U2086 (N_2086,N_887,N_648);
and U2087 (N_2087,N_121,N_367);
or U2088 (N_2088,N_1419,N_973);
nor U2089 (N_2089,N_165,N_130);
xor U2090 (N_2090,N_911,N_734);
nand U2091 (N_2091,N_181,N_462);
nor U2092 (N_2092,N_1243,N_1022);
and U2093 (N_2093,N_249,N_913);
xor U2094 (N_2094,N_882,N_907);
or U2095 (N_2095,N_413,N_19);
nor U2096 (N_2096,N_709,N_35);
or U2097 (N_2097,N_686,N_633);
xor U2098 (N_2098,N_562,N_186);
nor U2099 (N_2099,N_1292,N_1343);
or U2100 (N_2100,N_118,N_1498);
nand U2101 (N_2101,N_772,N_792);
or U2102 (N_2102,N_1226,N_1358);
or U2103 (N_2103,N_10,N_605);
and U2104 (N_2104,N_906,N_1341);
nor U2105 (N_2105,N_403,N_452);
nand U2106 (N_2106,N_93,N_683);
and U2107 (N_2107,N_149,N_1200);
xor U2108 (N_2108,N_748,N_789);
nor U2109 (N_2109,N_766,N_1433);
nor U2110 (N_2110,N_449,N_1356);
and U2111 (N_2111,N_1199,N_651);
or U2112 (N_2112,N_722,N_969);
xnor U2113 (N_2113,N_1052,N_937);
xor U2114 (N_2114,N_747,N_1051);
xnor U2115 (N_2115,N_168,N_1203);
nand U2116 (N_2116,N_845,N_1137);
nand U2117 (N_2117,N_976,N_656);
nand U2118 (N_2118,N_227,N_638);
or U2119 (N_2119,N_800,N_279);
nor U2120 (N_2120,N_870,N_1312);
and U2121 (N_2121,N_930,N_325);
nor U2122 (N_2122,N_6,N_259);
nor U2123 (N_2123,N_410,N_799);
and U2124 (N_2124,N_688,N_295);
nor U2125 (N_2125,N_323,N_1468);
nand U2126 (N_2126,N_964,N_576);
or U2127 (N_2127,N_123,N_497);
and U2128 (N_2128,N_1194,N_117);
and U2129 (N_2129,N_1315,N_731);
or U2130 (N_2130,N_338,N_386);
or U2131 (N_2131,N_819,N_1019);
nor U2132 (N_2132,N_1489,N_478);
and U2133 (N_2133,N_1476,N_1184);
or U2134 (N_2134,N_718,N_26);
nand U2135 (N_2135,N_1100,N_385);
and U2136 (N_2136,N_1478,N_470);
or U2137 (N_2137,N_242,N_312);
nand U2138 (N_2138,N_137,N_1165);
or U2139 (N_2139,N_692,N_447);
xor U2140 (N_2140,N_1188,N_9);
nor U2141 (N_2141,N_1304,N_980);
nor U2142 (N_2142,N_1086,N_320);
nor U2143 (N_2143,N_857,N_1317);
or U2144 (N_2144,N_645,N_750);
xnor U2145 (N_2145,N_1152,N_802);
nor U2146 (N_2146,N_1158,N_257);
or U2147 (N_2147,N_202,N_546);
or U2148 (N_2148,N_1327,N_564);
and U2149 (N_2149,N_1388,N_382);
and U2150 (N_2150,N_61,N_971);
or U2151 (N_2151,N_615,N_521);
and U2152 (N_2152,N_624,N_1284);
xor U2153 (N_2153,N_188,N_596);
nand U2154 (N_2154,N_483,N_768);
and U2155 (N_2155,N_1173,N_662);
or U2156 (N_2156,N_3,N_512);
nor U2157 (N_2157,N_444,N_1420);
and U2158 (N_2158,N_1085,N_1459);
xor U2159 (N_2159,N_524,N_102);
and U2160 (N_2160,N_133,N_1186);
nor U2161 (N_2161,N_623,N_1195);
xnor U2162 (N_2162,N_1486,N_1466);
xor U2163 (N_2163,N_1091,N_838);
nor U2164 (N_2164,N_458,N_481);
xor U2165 (N_2165,N_209,N_522);
nor U2166 (N_2166,N_1379,N_514);
nor U2167 (N_2167,N_1021,N_1402);
and U2168 (N_2168,N_459,N_305);
nand U2169 (N_2169,N_1367,N_871);
and U2170 (N_2170,N_952,N_1111);
or U2171 (N_2171,N_1465,N_652);
or U2172 (N_2172,N_1451,N_1384);
and U2173 (N_2173,N_732,N_1301);
nand U2174 (N_2174,N_554,N_901);
and U2175 (N_2175,N_1043,N_299);
or U2176 (N_2176,N_490,N_1357);
and U2177 (N_2177,N_1232,N_830);
or U2178 (N_2178,N_269,N_851);
and U2179 (N_2179,N_1436,N_66);
xor U2180 (N_2180,N_555,N_874);
nand U2181 (N_2181,N_285,N_1380);
and U2182 (N_2182,N_844,N_224);
xor U2183 (N_2183,N_691,N_248);
and U2184 (N_2184,N_203,N_791);
or U2185 (N_2185,N_1037,N_1023);
nand U2186 (N_2186,N_28,N_1002);
or U2187 (N_2187,N_463,N_327);
xor U2188 (N_2188,N_1075,N_1018);
nand U2189 (N_2189,N_674,N_167);
or U2190 (N_2190,N_1069,N_334);
xnor U2191 (N_2191,N_758,N_1136);
and U2192 (N_2192,N_900,N_329);
nand U2193 (N_2193,N_1028,N_32);
nand U2194 (N_2194,N_308,N_294);
nand U2195 (N_2195,N_744,N_1370);
nor U2196 (N_2196,N_375,N_13);
nor U2197 (N_2197,N_1467,N_1283);
xor U2198 (N_2198,N_212,N_898);
xor U2199 (N_2199,N_190,N_1351);
or U2200 (N_2200,N_17,N_577);
nand U2201 (N_2201,N_1455,N_836);
nor U2202 (N_2202,N_57,N_501);
nor U2203 (N_2203,N_336,N_977);
nand U2204 (N_2204,N_1499,N_703);
and U2205 (N_2205,N_642,N_706);
xor U2206 (N_2206,N_1072,N_762);
nor U2207 (N_2207,N_45,N_321);
or U2208 (N_2208,N_183,N_1105);
nor U2209 (N_2209,N_1089,N_191);
and U2210 (N_2210,N_414,N_1164);
xnor U2211 (N_2211,N_1049,N_237);
and U2212 (N_2212,N_430,N_1277);
xor U2213 (N_2213,N_1252,N_24);
and U2214 (N_2214,N_1355,N_689);
or U2215 (N_2215,N_821,N_597);
nand U2216 (N_2216,N_1060,N_1299);
and U2217 (N_2217,N_1206,N_803);
xor U2218 (N_2218,N_1483,N_540);
or U2219 (N_2219,N_1231,N_274);
or U2220 (N_2220,N_272,N_707);
and U2221 (N_2221,N_11,N_1495);
and U2222 (N_2222,N_1094,N_828);
nand U2223 (N_2223,N_99,N_865);
or U2224 (N_2224,N_974,N_275);
or U2225 (N_2225,N_1401,N_1335);
or U2226 (N_2226,N_354,N_128);
and U2227 (N_2227,N_347,N_503);
and U2228 (N_2228,N_94,N_219);
and U2229 (N_2229,N_415,N_1248);
or U2230 (N_2230,N_1172,N_1374);
or U2231 (N_2231,N_261,N_1316);
nor U2232 (N_2232,N_180,N_391);
nand U2233 (N_2233,N_711,N_511);
nand U2234 (N_2234,N_150,N_1346);
nand U2235 (N_2235,N_529,N_682);
and U2236 (N_2236,N_1212,N_1336);
nor U2237 (N_2237,N_634,N_297);
nor U2238 (N_2238,N_1159,N_780);
nor U2239 (N_2239,N_986,N_397);
nor U2240 (N_2240,N_469,N_247);
nor U2241 (N_2241,N_1392,N_557);
nand U2242 (N_2242,N_474,N_21);
and U2243 (N_2243,N_570,N_1221);
and U2244 (N_2244,N_814,N_402);
nor U2245 (N_2245,N_394,N_1000);
nor U2246 (N_2246,N_81,N_1262);
xnor U2247 (N_2247,N_1109,N_162);
nand U2248 (N_2248,N_1289,N_640);
or U2249 (N_2249,N_76,N_20);
and U2250 (N_2250,N_405,N_659);
or U2251 (N_2251,N_1179,N_1081);
nor U2252 (N_2252,N_1037,N_326);
nand U2253 (N_2253,N_288,N_1491);
or U2254 (N_2254,N_322,N_1084);
nand U2255 (N_2255,N_386,N_704);
nand U2256 (N_2256,N_716,N_669);
nor U2257 (N_2257,N_1136,N_494);
or U2258 (N_2258,N_813,N_310);
nor U2259 (N_2259,N_272,N_1094);
and U2260 (N_2260,N_841,N_425);
or U2261 (N_2261,N_1446,N_636);
nand U2262 (N_2262,N_863,N_1424);
and U2263 (N_2263,N_339,N_496);
nand U2264 (N_2264,N_422,N_1238);
nor U2265 (N_2265,N_1007,N_1142);
nand U2266 (N_2266,N_68,N_1308);
or U2267 (N_2267,N_834,N_607);
nor U2268 (N_2268,N_956,N_284);
nor U2269 (N_2269,N_413,N_747);
and U2270 (N_2270,N_1000,N_14);
nand U2271 (N_2271,N_969,N_711);
or U2272 (N_2272,N_881,N_695);
nor U2273 (N_2273,N_649,N_815);
xnor U2274 (N_2274,N_1027,N_1118);
nand U2275 (N_2275,N_605,N_989);
or U2276 (N_2276,N_313,N_287);
or U2277 (N_2277,N_1387,N_674);
xor U2278 (N_2278,N_1327,N_1051);
nor U2279 (N_2279,N_462,N_1001);
and U2280 (N_2280,N_750,N_52);
nor U2281 (N_2281,N_299,N_727);
nand U2282 (N_2282,N_1152,N_863);
and U2283 (N_2283,N_267,N_787);
nand U2284 (N_2284,N_495,N_676);
nor U2285 (N_2285,N_555,N_428);
nand U2286 (N_2286,N_214,N_492);
and U2287 (N_2287,N_1073,N_570);
or U2288 (N_2288,N_723,N_392);
xnor U2289 (N_2289,N_638,N_1386);
nor U2290 (N_2290,N_892,N_0);
nor U2291 (N_2291,N_34,N_451);
or U2292 (N_2292,N_1074,N_31);
and U2293 (N_2293,N_1428,N_815);
nand U2294 (N_2294,N_1421,N_1182);
nor U2295 (N_2295,N_452,N_1483);
nor U2296 (N_2296,N_763,N_1263);
nor U2297 (N_2297,N_1340,N_298);
nand U2298 (N_2298,N_905,N_480);
nand U2299 (N_2299,N_466,N_303);
nor U2300 (N_2300,N_1146,N_939);
xor U2301 (N_2301,N_905,N_81);
and U2302 (N_2302,N_398,N_659);
nor U2303 (N_2303,N_169,N_1171);
nand U2304 (N_2304,N_692,N_790);
nor U2305 (N_2305,N_673,N_1247);
xnor U2306 (N_2306,N_643,N_688);
xnor U2307 (N_2307,N_1287,N_473);
nor U2308 (N_2308,N_722,N_237);
and U2309 (N_2309,N_953,N_1005);
or U2310 (N_2310,N_1476,N_32);
and U2311 (N_2311,N_835,N_485);
xor U2312 (N_2312,N_1039,N_311);
or U2313 (N_2313,N_1139,N_10);
and U2314 (N_2314,N_299,N_989);
or U2315 (N_2315,N_484,N_1124);
xnor U2316 (N_2316,N_111,N_517);
and U2317 (N_2317,N_1083,N_665);
and U2318 (N_2318,N_866,N_1227);
or U2319 (N_2319,N_138,N_1068);
or U2320 (N_2320,N_1239,N_817);
or U2321 (N_2321,N_499,N_190);
and U2322 (N_2322,N_784,N_520);
nand U2323 (N_2323,N_276,N_155);
or U2324 (N_2324,N_1045,N_696);
nor U2325 (N_2325,N_375,N_1484);
nand U2326 (N_2326,N_474,N_130);
or U2327 (N_2327,N_1102,N_1222);
xnor U2328 (N_2328,N_1024,N_583);
or U2329 (N_2329,N_317,N_1228);
nor U2330 (N_2330,N_60,N_1060);
and U2331 (N_2331,N_376,N_1347);
nor U2332 (N_2332,N_437,N_954);
xnor U2333 (N_2333,N_382,N_1425);
nor U2334 (N_2334,N_714,N_297);
nor U2335 (N_2335,N_320,N_847);
xor U2336 (N_2336,N_725,N_294);
nor U2337 (N_2337,N_209,N_265);
nand U2338 (N_2338,N_164,N_341);
nand U2339 (N_2339,N_926,N_617);
xor U2340 (N_2340,N_5,N_1496);
xnor U2341 (N_2341,N_1061,N_1482);
or U2342 (N_2342,N_507,N_1182);
nand U2343 (N_2343,N_1145,N_700);
xnor U2344 (N_2344,N_1442,N_944);
and U2345 (N_2345,N_80,N_750);
nor U2346 (N_2346,N_567,N_1161);
nand U2347 (N_2347,N_679,N_1373);
and U2348 (N_2348,N_914,N_1309);
or U2349 (N_2349,N_1437,N_27);
xor U2350 (N_2350,N_1201,N_1458);
or U2351 (N_2351,N_96,N_335);
or U2352 (N_2352,N_636,N_659);
or U2353 (N_2353,N_587,N_1096);
nand U2354 (N_2354,N_211,N_428);
or U2355 (N_2355,N_1304,N_1122);
or U2356 (N_2356,N_511,N_177);
nor U2357 (N_2357,N_1342,N_693);
or U2358 (N_2358,N_1157,N_346);
and U2359 (N_2359,N_1496,N_292);
nand U2360 (N_2360,N_568,N_1355);
or U2361 (N_2361,N_512,N_747);
or U2362 (N_2362,N_1072,N_161);
xor U2363 (N_2363,N_1408,N_360);
or U2364 (N_2364,N_1107,N_1077);
nand U2365 (N_2365,N_1211,N_1062);
or U2366 (N_2366,N_248,N_398);
nor U2367 (N_2367,N_592,N_654);
nor U2368 (N_2368,N_644,N_754);
nor U2369 (N_2369,N_602,N_559);
nand U2370 (N_2370,N_1036,N_1336);
or U2371 (N_2371,N_156,N_1405);
nand U2372 (N_2372,N_236,N_259);
and U2373 (N_2373,N_1403,N_806);
nand U2374 (N_2374,N_1332,N_1084);
or U2375 (N_2375,N_1070,N_42);
or U2376 (N_2376,N_1118,N_407);
or U2377 (N_2377,N_1287,N_1188);
nand U2378 (N_2378,N_1195,N_580);
nor U2379 (N_2379,N_1460,N_849);
or U2380 (N_2380,N_177,N_752);
or U2381 (N_2381,N_1321,N_1072);
nand U2382 (N_2382,N_1106,N_1187);
or U2383 (N_2383,N_437,N_919);
nand U2384 (N_2384,N_666,N_1033);
nand U2385 (N_2385,N_938,N_444);
nand U2386 (N_2386,N_217,N_1382);
and U2387 (N_2387,N_954,N_446);
nand U2388 (N_2388,N_1262,N_954);
nand U2389 (N_2389,N_1420,N_205);
and U2390 (N_2390,N_198,N_1430);
nor U2391 (N_2391,N_578,N_127);
and U2392 (N_2392,N_1372,N_1367);
and U2393 (N_2393,N_945,N_408);
and U2394 (N_2394,N_40,N_386);
xor U2395 (N_2395,N_1045,N_501);
nand U2396 (N_2396,N_186,N_626);
and U2397 (N_2397,N_1480,N_664);
nand U2398 (N_2398,N_365,N_931);
or U2399 (N_2399,N_1119,N_156);
xor U2400 (N_2400,N_1305,N_1266);
or U2401 (N_2401,N_805,N_951);
and U2402 (N_2402,N_434,N_696);
xor U2403 (N_2403,N_947,N_703);
nand U2404 (N_2404,N_745,N_1416);
nand U2405 (N_2405,N_1393,N_1154);
or U2406 (N_2406,N_1335,N_1168);
and U2407 (N_2407,N_374,N_25);
and U2408 (N_2408,N_1374,N_845);
and U2409 (N_2409,N_340,N_1301);
xnor U2410 (N_2410,N_1009,N_800);
and U2411 (N_2411,N_1240,N_1473);
xnor U2412 (N_2412,N_1105,N_757);
nor U2413 (N_2413,N_75,N_861);
nand U2414 (N_2414,N_1250,N_394);
nand U2415 (N_2415,N_902,N_854);
xor U2416 (N_2416,N_844,N_1334);
nand U2417 (N_2417,N_1088,N_1319);
nor U2418 (N_2418,N_321,N_1475);
or U2419 (N_2419,N_1051,N_548);
xnor U2420 (N_2420,N_868,N_821);
nand U2421 (N_2421,N_743,N_328);
and U2422 (N_2422,N_1248,N_643);
xnor U2423 (N_2423,N_882,N_754);
or U2424 (N_2424,N_1428,N_17);
nand U2425 (N_2425,N_944,N_21);
nor U2426 (N_2426,N_932,N_1113);
nor U2427 (N_2427,N_580,N_475);
and U2428 (N_2428,N_1038,N_1286);
and U2429 (N_2429,N_1492,N_65);
nor U2430 (N_2430,N_1353,N_86);
nand U2431 (N_2431,N_968,N_1182);
nand U2432 (N_2432,N_888,N_1042);
or U2433 (N_2433,N_478,N_1266);
or U2434 (N_2434,N_1487,N_1377);
xnor U2435 (N_2435,N_1252,N_1359);
xor U2436 (N_2436,N_1369,N_1010);
nand U2437 (N_2437,N_424,N_346);
or U2438 (N_2438,N_1300,N_400);
xor U2439 (N_2439,N_347,N_590);
nor U2440 (N_2440,N_903,N_1229);
xnor U2441 (N_2441,N_861,N_13);
nand U2442 (N_2442,N_1415,N_1222);
xnor U2443 (N_2443,N_1246,N_1195);
nor U2444 (N_2444,N_525,N_425);
and U2445 (N_2445,N_371,N_1435);
and U2446 (N_2446,N_548,N_1030);
or U2447 (N_2447,N_1270,N_309);
or U2448 (N_2448,N_301,N_855);
nor U2449 (N_2449,N_585,N_851);
xor U2450 (N_2450,N_904,N_584);
nand U2451 (N_2451,N_634,N_1248);
and U2452 (N_2452,N_76,N_1367);
or U2453 (N_2453,N_836,N_586);
xnor U2454 (N_2454,N_364,N_1012);
xor U2455 (N_2455,N_499,N_469);
or U2456 (N_2456,N_693,N_1323);
or U2457 (N_2457,N_1178,N_172);
xnor U2458 (N_2458,N_1417,N_339);
and U2459 (N_2459,N_723,N_194);
nor U2460 (N_2460,N_1120,N_326);
or U2461 (N_2461,N_1451,N_1302);
nor U2462 (N_2462,N_1085,N_283);
and U2463 (N_2463,N_838,N_1153);
nor U2464 (N_2464,N_951,N_709);
nor U2465 (N_2465,N_259,N_17);
xnor U2466 (N_2466,N_1108,N_1170);
nand U2467 (N_2467,N_331,N_839);
and U2468 (N_2468,N_894,N_161);
nor U2469 (N_2469,N_1355,N_1379);
xnor U2470 (N_2470,N_845,N_273);
or U2471 (N_2471,N_465,N_1203);
xor U2472 (N_2472,N_1489,N_750);
and U2473 (N_2473,N_581,N_781);
nor U2474 (N_2474,N_1193,N_459);
and U2475 (N_2475,N_300,N_1311);
nor U2476 (N_2476,N_12,N_617);
and U2477 (N_2477,N_951,N_53);
nand U2478 (N_2478,N_724,N_595);
nand U2479 (N_2479,N_1346,N_427);
xor U2480 (N_2480,N_1434,N_909);
nand U2481 (N_2481,N_920,N_17);
xnor U2482 (N_2482,N_1210,N_873);
xor U2483 (N_2483,N_334,N_288);
nor U2484 (N_2484,N_1232,N_231);
xor U2485 (N_2485,N_86,N_5);
nand U2486 (N_2486,N_1329,N_901);
or U2487 (N_2487,N_457,N_33);
xnor U2488 (N_2488,N_427,N_591);
xor U2489 (N_2489,N_1051,N_1052);
nor U2490 (N_2490,N_348,N_474);
and U2491 (N_2491,N_1340,N_556);
nand U2492 (N_2492,N_653,N_1191);
nand U2493 (N_2493,N_1325,N_189);
and U2494 (N_2494,N_978,N_30);
nor U2495 (N_2495,N_115,N_303);
nand U2496 (N_2496,N_1168,N_247);
xnor U2497 (N_2497,N_1273,N_1415);
nand U2498 (N_2498,N_1121,N_919);
or U2499 (N_2499,N_1262,N_602);
and U2500 (N_2500,N_1221,N_662);
xor U2501 (N_2501,N_1485,N_535);
nor U2502 (N_2502,N_182,N_822);
nand U2503 (N_2503,N_1243,N_793);
nor U2504 (N_2504,N_910,N_1225);
nand U2505 (N_2505,N_363,N_42);
or U2506 (N_2506,N_563,N_1005);
xnor U2507 (N_2507,N_1173,N_1455);
nor U2508 (N_2508,N_411,N_1255);
nor U2509 (N_2509,N_1366,N_397);
nor U2510 (N_2510,N_1017,N_1322);
nand U2511 (N_2511,N_561,N_870);
nand U2512 (N_2512,N_367,N_801);
and U2513 (N_2513,N_722,N_1116);
or U2514 (N_2514,N_1173,N_1058);
xor U2515 (N_2515,N_1043,N_164);
nor U2516 (N_2516,N_1213,N_1490);
or U2517 (N_2517,N_753,N_914);
nand U2518 (N_2518,N_296,N_1084);
nand U2519 (N_2519,N_5,N_1031);
xor U2520 (N_2520,N_188,N_583);
or U2521 (N_2521,N_197,N_191);
nand U2522 (N_2522,N_900,N_1089);
or U2523 (N_2523,N_1269,N_336);
nor U2524 (N_2524,N_764,N_1083);
xnor U2525 (N_2525,N_549,N_479);
or U2526 (N_2526,N_647,N_399);
and U2527 (N_2527,N_1057,N_1464);
and U2528 (N_2528,N_491,N_275);
nor U2529 (N_2529,N_778,N_1248);
nand U2530 (N_2530,N_780,N_1452);
or U2531 (N_2531,N_1490,N_184);
or U2532 (N_2532,N_251,N_707);
or U2533 (N_2533,N_168,N_501);
or U2534 (N_2534,N_1075,N_724);
or U2535 (N_2535,N_1440,N_489);
nand U2536 (N_2536,N_453,N_966);
nor U2537 (N_2537,N_1069,N_1415);
nor U2538 (N_2538,N_1364,N_9);
or U2539 (N_2539,N_1086,N_968);
nand U2540 (N_2540,N_591,N_1177);
and U2541 (N_2541,N_1188,N_24);
or U2542 (N_2542,N_968,N_881);
nor U2543 (N_2543,N_1148,N_1029);
nand U2544 (N_2544,N_1303,N_182);
xor U2545 (N_2545,N_493,N_418);
and U2546 (N_2546,N_1117,N_569);
nor U2547 (N_2547,N_269,N_1408);
and U2548 (N_2548,N_251,N_1309);
nand U2549 (N_2549,N_1392,N_1211);
and U2550 (N_2550,N_77,N_660);
or U2551 (N_2551,N_78,N_1380);
or U2552 (N_2552,N_1399,N_1486);
and U2553 (N_2553,N_245,N_613);
xnor U2554 (N_2554,N_1422,N_693);
nor U2555 (N_2555,N_566,N_1175);
xnor U2556 (N_2556,N_1069,N_1397);
or U2557 (N_2557,N_274,N_437);
xnor U2558 (N_2558,N_1161,N_233);
or U2559 (N_2559,N_143,N_414);
nand U2560 (N_2560,N_740,N_144);
nand U2561 (N_2561,N_907,N_26);
nand U2562 (N_2562,N_1323,N_1276);
xnor U2563 (N_2563,N_880,N_1260);
and U2564 (N_2564,N_430,N_698);
and U2565 (N_2565,N_933,N_1375);
and U2566 (N_2566,N_828,N_1499);
or U2567 (N_2567,N_721,N_1478);
nor U2568 (N_2568,N_461,N_799);
xor U2569 (N_2569,N_83,N_305);
nand U2570 (N_2570,N_241,N_460);
nor U2571 (N_2571,N_1101,N_672);
or U2572 (N_2572,N_841,N_508);
nor U2573 (N_2573,N_830,N_333);
xnor U2574 (N_2574,N_977,N_1380);
and U2575 (N_2575,N_2,N_925);
xor U2576 (N_2576,N_701,N_1473);
nand U2577 (N_2577,N_491,N_1116);
xor U2578 (N_2578,N_1141,N_700);
xor U2579 (N_2579,N_1055,N_1143);
nand U2580 (N_2580,N_183,N_1069);
nand U2581 (N_2581,N_692,N_1088);
nand U2582 (N_2582,N_492,N_1399);
xor U2583 (N_2583,N_1359,N_1377);
nand U2584 (N_2584,N_758,N_281);
and U2585 (N_2585,N_1306,N_323);
nor U2586 (N_2586,N_1295,N_972);
xor U2587 (N_2587,N_1400,N_281);
or U2588 (N_2588,N_324,N_1046);
nor U2589 (N_2589,N_1094,N_636);
xnor U2590 (N_2590,N_889,N_379);
and U2591 (N_2591,N_182,N_59);
nand U2592 (N_2592,N_462,N_1475);
nand U2593 (N_2593,N_36,N_1061);
or U2594 (N_2594,N_246,N_729);
and U2595 (N_2595,N_484,N_798);
or U2596 (N_2596,N_771,N_100);
or U2597 (N_2597,N_738,N_1020);
nand U2598 (N_2598,N_886,N_828);
nor U2599 (N_2599,N_782,N_889);
and U2600 (N_2600,N_717,N_1272);
and U2601 (N_2601,N_1178,N_1056);
and U2602 (N_2602,N_636,N_375);
and U2603 (N_2603,N_44,N_1064);
xor U2604 (N_2604,N_984,N_707);
nor U2605 (N_2605,N_375,N_587);
and U2606 (N_2606,N_414,N_739);
nor U2607 (N_2607,N_102,N_1397);
xnor U2608 (N_2608,N_851,N_1162);
nand U2609 (N_2609,N_150,N_1162);
or U2610 (N_2610,N_126,N_302);
and U2611 (N_2611,N_247,N_19);
and U2612 (N_2612,N_260,N_1052);
or U2613 (N_2613,N_861,N_347);
or U2614 (N_2614,N_901,N_1441);
nand U2615 (N_2615,N_111,N_1103);
nor U2616 (N_2616,N_345,N_697);
and U2617 (N_2617,N_309,N_367);
nor U2618 (N_2618,N_273,N_1159);
or U2619 (N_2619,N_256,N_1246);
or U2620 (N_2620,N_727,N_231);
xnor U2621 (N_2621,N_88,N_42);
nand U2622 (N_2622,N_117,N_286);
and U2623 (N_2623,N_300,N_279);
nor U2624 (N_2624,N_357,N_120);
nor U2625 (N_2625,N_782,N_716);
and U2626 (N_2626,N_1434,N_882);
xor U2627 (N_2627,N_63,N_409);
xnor U2628 (N_2628,N_353,N_1370);
and U2629 (N_2629,N_1416,N_447);
nor U2630 (N_2630,N_204,N_406);
nand U2631 (N_2631,N_219,N_456);
and U2632 (N_2632,N_274,N_693);
xor U2633 (N_2633,N_374,N_741);
and U2634 (N_2634,N_1035,N_935);
xnor U2635 (N_2635,N_46,N_591);
and U2636 (N_2636,N_625,N_430);
xor U2637 (N_2637,N_1189,N_813);
nand U2638 (N_2638,N_986,N_1236);
or U2639 (N_2639,N_152,N_1212);
xor U2640 (N_2640,N_814,N_1240);
nor U2641 (N_2641,N_807,N_535);
or U2642 (N_2642,N_105,N_1329);
and U2643 (N_2643,N_1400,N_946);
or U2644 (N_2644,N_190,N_1030);
nor U2645 (N_2645,N_976,N_1379);
xnor U2646 (N_2646,N_447,N_1305);
or U2647 (N_2647,N_526,N_963);
nand U2648 (N_2648,N_1196,N_1406);
or U2649 (N_2649,N_951,N_863);
nand U2650 (N_2650,N_817,N_813);
nor U2651 (N_2651,N_127,N_428);
nor U2652 (N_2652,N_449,N_503);
xor U2653 (N_2653,N_1087,N_1405);
xor U2654 (N_2654,N_982,N_846);
or U2655 (N_2655,N_1364,N_204);
and U2656 (N_2656,N_646,N_1338);
xor U2657 (N_2657,N_290,N_193);
xor U2658 (N_2658,N_553,N_1379);
nand U2659 (N_2659,N_1443,N_454);
or U2660 (N_2660,N_710,N_50);
or U2661 (N_2661,N_76,N_115);
and U2662 (N_2662,N_208,N_1383);
or U2663 (N_2663,N_504,N_554);
or U2664 (N_2664,N_1009,N_911);
and U2665 (N_2665,N_1113,N_1254);
and U2666 (N_2666,N_378,N_505);
nand U2667 (N_2667,N_937,N_1021);
xor U2668 (N_2668,N_516,N_1115);
nor U2669 (N_2669,N_657,N_1138);
xnor U2670 (N_2670,N_1481,N_1257);
or U2671 (N_2671,N_435,N_1283);
xor U2672 (N_2672,N_61,N_693);
or U2673 (N_2673,N_866,N_194);
and U2674 (N_2674,N_608,N_1271);
or U2675 (N_2675,N_377,N_572);
and U2676 (N_2676,N_910,N_1138);
xor U2677 (N_2677,N_950,N_958);
xnor U2678 (N_2678,N_790,N_187);
nand U2679 (N_2679,N_621,N_544);
nor U2680 (N_2680,N_1381,N_105);
xor U2681 (N_2681,N_1356,N_275);
nand U2682 (N_2682,N_594,N_525);
xor U2683 (N_2683,N_667,N_746);
xor U2684 (N_2684,N_1476,N_1468);
nor U2685 (N_2685,N_149,N_9);
nor U2686 (N_2686,N_1412,N_826);
xor U2687 (N_2687,N_887,N_192);
nand U2688 (N_2688,N_448,N_807);
nand U2689 (N_2689,N_156,N_1386);
xnor U2690 (N_2690,N_542,N_1244);
nor U2691 (N_2691,N_162,N_985);
xnor U2692 (N_2692,N_833,N_257);
xor U2693 (N_2693,N_207,N_243);
and U2694 (N_2694,N_747,N_859);
xor U2695 (N_2695,N_564,N_789);
nor U2696 (N_2696,N_24,N_1003);
nand U2697 (N_2697,N_253,N_1431);
nor U2698 (N_2698,N_63,N_314);
xnor U2699 (N_2699,N_867,N_329);
and U2700 (N_2700,N_301,N_1277);
xnor U2701 (N_2701,N_1052,N_1258);
and U2702 (N_2702,N_1402,N_30);
and U2703 (N_2703,N_913,N_533);
or U2704 (N_2704,N_577,N_1154);
and U2705 (N_2705,N_1466,N_66);
and U2706 (N_2706,N_939,N_1087);
and U2707 (N_2707,N_251,N_1314);
nor U2708 (N_2708,N_168,N_444);
nor U2709 (N_2709,N_228,N_267);
and U2710 (N_2710,N_913,N_1046);
and U2711 (N_2711,N_1069,N_1416);
or U2712 (N_2712,N_1172,N_88);
or U2713 (N_2713,N_897,N_543);
xor U2714 (N_2714,N_14,N_1332);
nand U2715 (N_2715,N_628,N_366);
nor U2716 (N_2716,N_0,N_725);
nor U2717 (N_2717,N_682,N_1090);
nand U2718 (N_2718,N_700,N_1316);
nand U2719 (N_2719,N_1042,N_1128);
or U2720 (N_2720,N_177,N_146);
nand U2721 (N_2721,N_1369,N_657);
nand U2722 (N_2722,N_1065,N_790);
and U2723 (N_2723,N_707,N_1107);
nor U2724 (N_2724,N_320,N_338);
nor U2725 (N_2725,N_626,N_896);
or U2726 (N_2726,N_683,N_1374);
nand U2727 (N_2727,N_622,N_1032);
or U2728 (N_2728,N_80,N_1081);
and U2729 (N_2729,N_214,N_1209);
or U2730 (N_2730,N_1317,N_974);
nor U2731 (N_2731,N_141,N_554);
and U2732 (N_2732,N_1211,N_462);
or U2733 (N_2733,N_269,N_677);
nand U2734 (N_2734,N_423,N_706);
nor U2735 (N_2735,N_1404,N_950);
or U2736 (N_2736,N_821,N_609);
xor U2737 (N_2737,N_1278,N_792);
or U2738 (N_2738,N_1024,N_537);
nor U2739 (N_2739,N_927,N_17);
or U2740 (N_2740,N_552,N_1172);
nor U2741 (N_2741,N_1437,N_993);
xor U2742 (N_2742,N_277,N_119);
nand U2743 (N_2743,N_1289,N_531);
or U2744 (N_2744,N_519,N_1010);
and U2745 (N_2745,N_20,N_414);
nor U2746 (N_2746,N_741,N_995);
nand U2747 (N_2747,N_696,N_601);
and U2748 (N_2748,N_1040,N_169);
nand U2749 (N_2749,N_734,N_1467);
and U2750 (N_2750,N_1117,N_683);
and U2751 (N_2751,N_526,N_430);
or U2752 (N_2752,N_401,N_810);
or U2753 (N_2753,N_27,N_888);
or U2754 (N_2754,N_134,N_233);
and U2755 (N_2755,N_148,N_763);
nor U2756 (N_2756,N_273,N_638);
and U2757 (N_2757,N_689,N_590);
or U2758 (N_2758,N_1276,N_651);
nor U2759 (N_2759,N_174,N_1100);
xnor U2760 (N_2760,N_1026,N_316);
and U2761 (N_2761,N_1306,N_72);
xor U2762 (N_2762,N_372,N_1252);
nand U2763 (N_2763,N_501,N_933);
and U2764 (N_2764,N_1099,N_244);
nand U2765 (N_2765,N_1118,N_505);
nor U2766 (N_2766,N_900,N_30);
nand U2767 (N_2767,N_1427,N_978);
xor U2768 (N_2768,N_329,N_150);
and U2769 (N_2769,N_1363,N_264);
and U2770 (N_2770,N_1345,N_193);
and U2771 (N_2771,N_98,N_625);
or U2772 (N_2772,N_495,N_283);
xor U2773 (N_2773,N_699,N_435);
nand U2774 (N_2774,N_956,N_324);
xnor U2775 (N_2775,N_888,N_1355);
nand U2776 (N_2776,N_643,N_291);
or U2777 (N_2777,N_788,N_167);
nand U2778 (N_2778,N_778,N_465);
nand U2779 (N_2779,N_663,N_391);
nor U2780 (N_2780,N_1195,N_607);
or U2781 (N_2781,N_598,N_424);
nor U2782 (N_2782,N_1170,N_1029);
nand U2783 (N_2783,N_602,N_413);
nor U2784 (N_2784,N_233,N_421);
nand U2785 (N_2785,N_1389,N_1192);
xnor U2786 (N_2786,N_1380,N_140);
or U2787 (N_2787,N_1285,N_900);
nor U2788 (N_2788,N_888,N_627);
and U2789 (N_2789,N_36,N_315);
xor U2790 (N_2790,N_267,N_117);
nand U2791 (N_2791,N_653,N_457);
and U2792 (N_2792,N_1028,N_705);
nor U2793 (N_2793,N_1302,N_371);
xnor U2794 (N_2794,N_903,N_1415);
and U2795 (N_2795,N_1056,N_862);
nor U2796 (N_2796,N_312,N_1491);
and U2797 (N_2797,N_1470,N_1302);
xnor U2798 (N_2798,N_830,N_1312);
nor U2799 (N_2799,N_1137,N_415);
nand U2800 (N_2800,N_325,N_751);
nand U2801 (N_2801,N_1458,N_1195);
nor U2802 (N_2802,N_117,N_11);
xor U2803 (N_2803,N_1045,N_802);
nor U2804 (N_2804,N_1108,N_792);
or U2805 (N_2805,N_244,N_780);
or U2806 (N_2806,N_527,N_1428);
nand U2807 (N_2807,N_298,N_623);
and U2808 (N_2808,N_125,N_713);
and U2809 (N_2809,N_673,N_1346);
nand U2810 (N_2810,N_1403,N_1329);
or U2811 (N_2811,N_820,N_1190);
xnor U2812 (N_2812,N_259,N_841);
xnor U2813 (N_2813,N_385,N_1051);
nand U2814 (N_2814,N_1319,N_731);
and U2815 (N_2815,N_859,N_656);
nand U2816 (N_2816,N_1125,N_941);
nor U2817 (N_2817,N_1011,N_684);
nand U2818 (N_2818,N_1016,N_858);
nand U2819 (N_2819,N_1449,N_1225);
xnor U2820 (N_2820,N_806,N_1264);
and U2821 (N_2821,N_1368,N_1195);
nor U2822 (N_2822,N_940,N_330);
or U2823 (N_2823,N_1112,N_923);
xor U2824 (N_2824,N_945,N_525);
nand U2825 (N_2825,N_254,N_1090);
nand U2826 (N_2826,N_921,N_721);
xor U2827 (N_2827,N_738,N_348);
nor U2828 (N_2828,N_740,N_19);
or U2829 (N_2829,N_574,N_1285);
nor U2830 (N_2830,N_539,N_152);
or U2831 (N_2831,N_1310,N_1116);
or U2832 (N_2832,N_522,N_1485);
or U2833 (N_2833,N_1390,N_64);
nand U2834 (N_2834,N_1434,N_1352);
nand U2835 (N_2835,N_173,N_206);
nand U2836 (N_2836,N_765,N_495);
and U2837 (N_2837,N_1067,N_609);
xnor U2838 (N_2838,N_786,N_1191);
nand U2839 (N_2839,N_597,N_33);
nand U2840 (N_2840,N_364,N_354);
or U2841 (N_2841,N_254,N_465);
and U2842 (N_2842,N_584,N_198);
or U2843 (N_2843,N_1370,N_1310);
xor U2844 (N_2844,N_777,N_1123);
nor U2845 (N_2845,N_1145,N_9);
nand U2846 (N_2846,N_1486,N_433);
or U2847 (N_2847,N_1167,N_344);
or U2848 (N_2848,N_350,N_647);
xnor U2849 (N_2849,N_51,N_1133);
nor U2850 (N_2850,N_1071,N_1377);
or U2851 (N_2851,N_224,N_1351);
or U2852 (N_2852,N_1015,N_632);
nor U2853 (N_2853,N_1297,N_86);
xor U2854 (N_2854,N_1147,N_727);
or U2855 (N_2855,N_865,N_603);
and U2856 (N_2856,N_606,N_985);
xor U2857 (N_2857,N_570,N_709);
xnor U2858 (N_2858,N_1296,N_909);
or U2859 (N_2859,N_589,N_321);
or U2860 (N_2860,N_315,N_288);
nor U2861 (N_2861,N_1129,N_754);
or U2862 (N_2862,N_262,N_789);
or U2863 (N_2863,N_572,N_508);
and U2864 (N_2864,N_720,N_160);
or U2865 (N_2865,N_631,N_817);
and U2866 (N_2866,N_1265,N_1384);
or U2867 (N_2867,N_78,N_388);
nand U2868 (N_2868,N_1121,N_830);
xor U2869 (N_2869,N_1113,N_751);
and U2870 (N_2870,N_863,N_491);
xnor U2871 (N_2871,N_1450,N_354);
and U2872 (N_2872,N_1354,N_877);
nor U2873 (N_2873,N_490,N_104);
nand U2874 (N_2874,N_211,N_194);
or U2875 (N_2875,N_692,N_681);
xnor U2876 (N_2876,N_276,N_779);
nand U2877 (N_2877,N_333,N_1018);
nand U2878 (N_2878,N_950,N_185);
and U2879 (N_2879,N_76,N_711);
nand U2880 (N_2880,N_100,N_1314);
xnor U2881 (N_2881,N_1140,N_1316);
nand U2882 (N_2882,N_1044,N_617);
and U2883 (N_2883,N_723,N_671);
nor U2884 (N_2884,N_154,N_1388);
or U2885 (N_2885,N_401,N_580);
nand U2886 (N_2886,N_712,N_682);
and U2887 (N_2887,N_333,N_514);
nor U2888 (N_2888,N_111,N_144);
nand U2889 (N_2889,N_579,N_1392);
xnor U2890 (N_2890,N_169,N_312);
and U2891 (N_2891,N_1020,N_1344);
nand U2892 (N_2892,N_1027,N_203);
nor U2893 (N_2893,N_249,N_1075);
and U2894 (N_2894,N_733,N_535);
xor U2895 (N_2895,N_1180,N_158);
nor U2896 (N_2896,N_223,N_938);
nor U2897 (N_2897,N_308,N_1288);
xor U2898 (N_2898,N_49,N_970);
nor U2899 (N_2899,N_648,N_729);
nand U2900 (N_2900,N_547,N_785);
nor U2901 (N_2901,N_995,N_417);
and U2902 (N_2902,N_1407,N_318);
or U2903 (N_2903,N_59,N_447);
xnor U2904 (N_2904,N_1185,N_139);
and U2905 (N_2905,N_568,N_1199);
and U2906 (N_2906,N_81,N_1363);
or U2907 (N_2907,N_500,N_1441);
and U2908 (N_2908,N_153,N_1163);
nor U2909 (N_2909,N_92,N_614);
and U2910 (N_2910,N_86,N_1348);
or U2911 (N_2911,N_266,N_301);
nor U2912 (N_2912,N_632,N_1277);
or U2913 (N_2913,N_486,N_545);
or U2914 (N_2914,N_8,N_486);
nor U2915 (N_2915,N_551,N_246);
or U2916 (N_2916,N_166,N_400);
or U2917 (N_2917,N_1116,N_1055);
nor U2918 (N_2918,N_1436,N_1281);
and U2919 (N_2919,N_253,N_804);
xor U2920 (N_2920,N_960,N_408);
or U2921 (N_2921,N_210,N_1084);
and U2922 (N_2922,N_1496,N_22);
and U2923 (N_2923,N_309,N_1125);
xnor U2924 (N_2924,N_92,N_599);
or U2925 (N_2925,N_976,N_1289);
and U2926 (N_2926,N_1029,N_1238);
nor U2927 (N_2927,N_1372,N_1279);
xnor U2928 (N_2928,N_634,N_1079);
xor U2929 (N_2929,N_1096,N_1065);
nor U2930 (N_2930,N_402,N_887);
or U2931 (N_2931,N_1485,N_1279);
or U2932 (N_2932,N_658,N_1078);
or U2933 (N_2933,N_488,N_1267);
nand U2934 (N_2934,N_252,N_797);
and U2935 (N_2935,N_277,N_791);
and U2936 (N_2936,N_406,N_873);
nand U2937 (N_2937,N_169,N_797);
nor U2938 (N_2938,N_549,N_1009);
xor U2939 (N_2939,N_892,N_531);
or U2940 (N_2940,N_129,N_497);
xor U2941 (N_2941,N_1188,N_696);
xnor U2942 (N_2942,N_15,N_665);
or U2943 (N_2943,N_1223,N_305);
xnor U2944 (N_2944,N_1189,N_219);
nor U2945 (N_2945,N_625,N_542);
xor U2946 (N_2946,N_240,N_1163);
nand U2947 (N_2947,N_927,N_255);
nor U2948 (N_2948,N_1271,N_676);
xnor U2949 (N_2949,N_471,N_1488);
nor U2950 (N_2950,N_200,N_654);
and U2951 (N_2951,N_1468,N_1187);
xnor U2952 (N_2952,N_412,N_1064);
and U2953 (N_2953,N_987,N_688);
nor U2954 (N_2954,N_1348,N_453);
or U2955 (N_2955,N_822,N_849);
and U2956 (N_2956,N_389,N_559);
nand U2957 (N_2957,N_309,N_258);
nor U2958 (N_2958,N_275,N_1087);
nor U2959 (N_2959,N_1206,N_1073);
or U2960 (N_2960,N_683,N_1414);
nand U2961 (N_2961,N_515,N_234);
nor U2962 (N_2962,N_1333,N_594);
or U2963 (N_2963,N_1485,N_545);
nand U2964 (N_2964,N_834,N_1139);
and U2965 (N_2965,N_1380,N_245);
and U2966 (N_2966,N_859,N_39);
or U2967 (N_2967,N_1432,N_970);
or U2968 (N_2968,N_105,N_284);
and U2969 (N_2969,N_826,N_751);
and U2970 (N_2970,N_1241,N_900);
or U2971 (N_2971,N_388,N_775);
nand U2972 (N_2972,N_1336,N_924);
and U2973 (N_2973,N_68,N_167);
or U2974 (N_2974,N_643,N_1026);
and U2975 (N_2975,N_1209,N_1334);
xor U2976 (N_2976,N_386,N_632);
nor U2977 (N_2977,N_717,N_944);
nand U2978 (N_2978,N_682,N_1132);
xnor U2979 (N_2979,N_446,N_677);
nor U2980 (N_2980,N_1339,N_1313);
nand U2981 (N_2981,N_602,N_978);
nor U2982 (N_2982,N_473,N_232);
or U2983 (N_2983,N_1131,N_1013);
nand U2984 (N_2984,N_1412,N_851);
nand U2985 (N_2985,N_421,N_230);
nor U2986 (N_2986,N_1053,N_1239);
nand U2987 (N_2987,N_102,N_1375);
nor U2988 (N_2988,N_739,N_1402);
nand U2989 (N_2989,N_1414,N_210);
xnor U2990 (N_2990,N_132,N_641);
or U2991 (N_2991,N_1231,N_1137);
or U2992 (N_2992,N_209,N_1458);
xnor U2993 (N_2993,N_379,N_1450);
or U2994 (N_2994,N_515,N_64);
or U2995 (N_2995,N_568,N_1387);
xor U2996 (N_2996,N_70,N_1290);
nor U2997 (N_2997,N_1087,N_931);
xor U2998 (N_2998,N_271,N_1326);
nor U2999 (N_2999,N_515,N_317);
xor U3000 (N_3000,N_2437,N_2912);
nand U3001 (N_3001,N_1821,N_1747);
nand U3002 (N_3002,N_2257,N_2462);
nand U3003 (N_3003,N_2501,N_2846);
xor U3004 (N_3004,N_2148,N_2538);
xor U3005 (N_3005,N_2705,N_2228);
or U3006 (N_3006,N_2533,N_2315);
xor U3007 (N_3007,N_2758,N_2837);
nor U3008 (N_3008,N_2702,N_2855);
xor U3009 (N_3009,N_2962,N_1594);
xnor U3010 (N_3010,N_2728,N_1520);
nor U3011 (N_3011,N_2102,N_2623);
xor U3012 (N_3012,N_1973,N_1970);
and U3013 (N_3013,N_2770,N_2339);
xor U3014 (N_3014,N_2067,N_1631);
xnor U3015 (N_3015,N_2982,N_2337);
xnor U3016 (N_3016,N_2262,N_1515);
nor U3017 (N_3017,N_2667,N_1602);
nor U3018 (N_3018,N_1660,N_2204);
xnor U3019 (N_3019,N_1711,N_2365);
nand U3020 (N_3020,N_2905,N_2447);
xnor U3021 (N_3021,N_2466,N_1591);
and U3022 (N_3022,N_2469,N_2787);
nor U3023 (N_3023,N_2924,N_1561);
xnor U3024 (N_3024,N_1829,N_2321);
nand U3025 (N_3025,N_2009,N_2738);
nor U3026 (N_3026,N_2778,N_2868);
xor U3027 (N_3027,N_2373,N_2986);
or U3028 (N_3028,N_2499,N_2866);
or U3029 (N_3029,N_2376,N_2381);
xor U3030 (N_3030,N_2159,N_2163);
or U3031 (N_3031,N_2045,N_2990);
nor U3032 (N_3032,N_2472,N_2700);
nand U3033 (N_3033,N_2757,N_2768);
or U3034 (N_3034,N_2856,N_2825);
nor U3035 (N_3035,N_2370,N_1518);
xnor U3036 (N_3036,N_2046,N_2545);
nor U3037 (N_3037,N_2920,N_1567);
or U3038 (N_3038,N_1869,N_2968);
or U3039 (N_3039,N_2195,N_2618);
or U3040 (N_3040,N_2998,N_2411);
nor U3041 (N_3041,N_2323,N_2526);
or U3042 (N_3042,N_2449,N_1578);
nand U3043 (N_3043,N_2566,N_1511);
nor U3044 (N_3044,N_2989,N_2026);
nand U3045 (N_3045,N_1742,N_2694);
or U3046 (N_3046,N_2767,N_2173);
xnor U3047 (N_3047,N_2823,N_2596);
and U3048 (N_3048,N_2620,N_2015);
and U3049 (N_3049,N_2053,N_1697);
nand U3050 (N_3050,N_1632,N_2624);
and U3051 (N_3051,N_2695,N_1813);
and U3052 (N_3052,N_1500,N_1663);
xnor U3053 (N_3053,N_2463,N_2429);
nor U3054 (N_3054,N_2632,N_2604);
nor U3055 (N_3055,N_2249,N_2049);
nand U3056 (N_3056,N_2030,N_1886);
nor U3057 (N_3057,N_1975,N_1887);
nand U3058 (N_3058,N_2608,N_2379);
xor U3059 (N_3059,N_1992,N_1895);
nor U3060 (N_3060,N_2369,N_2577);
xnor U3061 (N_3061,N_1956,N_2503);
and U3062 (N_3062,N_2210,N_1530);
or U3063 (N_3063,N_2719,N_2234);
nor U3064 (N_3064,N_2607,N_1665);
xnor U3065 (N_3065,N_2089,N_1864);
or U3066 (N_3066,N_2384,N_2000);
and U3067 (N_3067,N_2415,N_2602);
nand U3068 (N_3068,N_2351,N_2523);
xnor U3069 (N_3069,N_2723,N_2683);
xnor U3070 (N_3070,N_2881,N_2814);
xnor U3071 (N_3071,N_2569,N_2413);
or U3072 (N_3072,N_1966,N_2421);
nand U3073 (N_3073,N_1873,N_1731);
nand U3074 (N_3074,N_2199,N_1793);
or U3075 (N_3075,N_1795,N_2600);
xnor U3076 (N_3076,N_1652,N_2169);
and U3077 (N_3077,N_2042,N_2091);
xor U3078 (N_3078,N_1807,N_2231);
nor U3079 (N_3079,N_1535,N_2997);
xnor U3080 (N_3080,N_2594,N_2528);
nor U3081 (N_3081,N_2753,N_1944);
nor U3082 (N_3082,N_1764,N_1983);
and U3083 (N_3083,N_2886,N_1712);
nand U3084 (N_3084,N_2966,N_2641);
xor U3085 (N_3085,N_2051,N_2489);
nand U3086 (N_3086,N_2140,N_1695);
nand U3087 (N_3087,N_1510,N_2542);
and U3088 (N_3088,N_2281,N_2587);
nand U3089 (N_3089,N_1748,N_2802);
xnor U3090 (N_3090,N_2827,N_2790);
xor U3091 (N_3091,N_1626,N_2335);
and U3092 (N_3092,N_2852,N_2108);
or U3093 (N_3093,N_2649,N_2079);
and U3094 (N_3094,N_2690,N_1693);
nor U3095 (N_3095,N_1884,N_2164);
or U3096 (N_3096,N_1949,N_1633);
nor U3097 (N_3097,N_2155,N_1568);
or U3098 (N_3098,N_2844,N_2237);
and U3099 (N_3099,N_1881,N_2522);
nand U3100 (N_3100,N_1553,N_1720);
and U3101 (N_3101,N_1902,N_2121);
nor U3102 (N_3102,N_2474,N_2166);
and U3103 (N_3103,N_1629,N_2959);
and U3104 (N_3104,N_1899,N_2047);
nand U3105 (N_3105,N_1668,N_2784);
and U3106 (N_3106,N_2263,N_2268);
or U3107 (N_3107,N_2675,N_1845);
nor U3108 (N_3108,N_2709,N_2934);
xor U3109 (N_3109,N_2652,N_1962);
and U3110 (N_3110,N_1686,N_2232);
and U3111 (N_3111,N_1732,N_1552);
and U3112 (N_3112,N_2725,N_1604);
or U3113 (N_3113,N_1984,N_2205);
nand U3114 (N_3114,N_2562,N_1737);
xor U3115 (N_3115,N_2185,N_2443);
and U3116 (N_3116,N_1818,N_2621);
nor U3117 (N_3117,N_2112,N_2253);
or U3118 (N_3118,N_1673,N_1825);
nand U3119 (N_3119,N_2760,N_2354);
or U3120 (N_3120,N_1539,N_2191);
or U3121 (N_3121,N_1613,N_2895);
nor U3122 (N_3122,N_2737,N_2378);
and U3123 (N_3123,N_2151,N_2282);
and U3124 (N_3124,N_2307,N_1601);
xnor U3125 (N_3125,N_1947,N_2961);
or U3126 (N_3126,N_1595,N_2084);
xor U3127 (N_3127,N_2459,N_2277);
nand U3128 (N_3128,N_2433,N_2888);
xnor U3129 (N_3129,N_1774,N_1565);
or U3130 (N_3130,N_2498,N_2976);
nand U3131 (N_3131,N_2104,N_2831);
nor U3132 (N_3132,N_2603,N_1506);
nand U3133 (N_3133,N_2028,N_2689);
nor U3134 (N_3134,N_2116,N_1932);
and U3135 (N_3135,N_2534,N_2175);
or U3136 (N_3136,N_2007,N_1819);
nor U3137 (N_3137,N_2039,N_2094);
and U3138 (N_3138,N_2201,N_2891);
nor U3139 (N_3139,N_2330,N_2877);
and U3140 (N_3140,N_2795,N_1637);
and U3141 (N_3141,N_2867,N_2525);
xor U3142 (N_3142,N_2983,N_2746);
xnor U3143 (N_3143,N_1855,N_1559);
nor U3144 (N_3144,N_2300,N_1541);
nor U3145 (N_3145,N_2589,N_1725);
and U3146 (N_3146,N_2898,N_1581);
nand U3147 (N_3147,N_1875,N_2082);
and U3148 (N_3148,N_2847,N_1779);
or U3149 (N_3149,N_2801,N_1710);
and U3150 (N_3150,N_1861,N_1880);
and U3151 (N_3151,N_2544,N_2254);
xnor U3152 (N_3152,N_2261,N_1741);
nand U3153 (N_3153,N_2014,N_2456);
and U3154 (N_3154,N_1790,N_1653);
xor U3155 (N_3155,N_1582,N_2060);
nor U3156 (N_3156,N_2440,N_2488);
or U3157 (N_3157,N_1909,N_1815);
nand U3158 (N_3158,N_2987,N_2633);
nand U3159 (N_3159,N_2763,N_1908);
and U3160 (N_3160,N_2657,N_2843);
xnor U3161 (N_3161,N_2154,N_2269);
and U3162 (N_3162,N_2988,N_1550);
nand U3163 (N_3163,N_1868,N_2054);
xor U3164 (N_3164,N_2111,N_1882);
nand U3165 (N_3165,N_1929,N_1726);
xnor U3166 (N_3166,N_2579,N_2804);
or U3167 (N_3167,N_1827,N_2884);
nand U3168 (N_3168,N_2017,N_1672);
and U3169 (N_3169,N_1914,N_1560);
or U3170 (N_3170,N_2333,N_2356);
xnor U3171 (N_3171,N_1941,N_1751);
xor U3172 (N_3172,N_2302,N_2118);
or U3173 (N_3173,N_1615,N_2643);
nand U3174 (N_3174,N_2996,N_2357);
and U3175 (N_3175,N_2640,N_2402);
and U3176 (N_3176,N_1920,N_2883);
nor U3177 (N_3177,N_2914,N_2259);
nand U3178 (N_3178,N_2434,N_2027);
nand U3179 (N_3179,N_2862,N_2087);
and U3180 (N_3180,N_2059,N_2001);
and U3181 (N_3181,N_1623,N_2043);
xnor U3182 (N_3182,N_1925,N_2771);
xnor U3183 (N_3183,N_2712,N_1658);
and U3184 (N_3184,N_1636,N_2214);
nor U3185 (N_3185,N_2114,N_2010);
xnor U3186 (N_3186,N_2482,N_2783);
nand U3187 (N_3187,N_1965,N_2793);
nor U3188 (N_3188,N_1799,N_2653);
nor U3189 (N_3189,N_2124,N_2960);
and U3190 (N_3190,N_2431,N_2505);
nor U3191 (N_3191,N_1507,N_2578);
xor U3192 (N_3192,N_2518,N_1856);
nor U3193 (N_3193,N_2865,N_1842);
xnor U3194 (N_3194,N_2872,N_2698);
or U3195 (N_3195,N_1716,N_2475);
xor U3196 (N_3196,N_2664,N_1577);
or U3197 (N_3197,N_1824,N_1890);
or U3198 (N_3198,N_1832,N_2050);
xor U3199 (N_3199,N_2860,N_2317);
nor U3200 (N_3200,N_2754,N_1717);
and U3201 (N_3201,N_2605,N_2575);
or U3202 (N_3202,N_2732,N_1900);
nand U3203 (N_3203,N_1554,N_2530);
or U3204 (N_3204,N_1876,N_1657);
xnor U3205 (N_3205,N_2994,N_2078);
or U3206 (N_3206,N_2404,N_2226);
and U3207 (N_3207,N_2264,N_2716);
and U3208 (N_3208,N_2452,N_2791);
and U3209 (N_3209,N_2899,N_1648);
nor U3210 (N_3210,N_1586,N_2340);
or U3211 (N_3211,N_2490,N_1617);
or U3212 (N_3212,N_2494,N_2985);
xor U3213 (N_3213,N_2517,N_1980);
or U3214 (N_3214,N_2828,N_2915);
and U3215 (N_3215,N_2752,N_2585);
and U3216 (N_3216,N_2182,N_2890);
xor U3217 (N_3217,N_2360,N_2703);
nor U3218 (N_3218,N_2341,N_2947);
nor U3219 (N_3219,N_2773,N_1974);
and U3220 (N_3220,N_2473,N_2691);
nand U3221 (N_3221,N_1706,N_2731);
or U3222 (N_3222,N_2240,N_2220);
and U3223 (N_3223,N_2152,N_2736);
and U3224 (N_3224,N_2869,N_2906);
nand U3225 (N_3225,N_1893,N_2808);
or U3226 (N_3226,N_2162,N_2919);
xor U3227 (N_3227,N_1757,N_2138);
xor U3228 (N_3228,N_2965,N_2574);
nand U3229 (N_3229,N_2838,N_1978);
xor U3230 (N_3230,N_1729,N_2171);
nand U3231 (N_3231,N_2468,N_1750);
and U3232 (N_3232,N_2077,N_2167);
xnor U3233 (N_3233,N_2244,N_2005);
or U3234 (N_3234,N_1718,N_1857);
or U3235 (N_3235,N_1698,N_1787);
xnor U3236 (N_3236,N_2227,N_2031);
xor U3237 (N_3237,N_2665,N_2021);
nand U3238 (N_3238,N_1843,N_2146);
or U3239 (N_3239,N_1620,N_2555);
xnor U3240 (N_3240,N_1847,N_1573);
nor U3241 (N_3241,N_2993,N_2943);
or U3242 (N_3242,N_2325,N_2180);
nand U3243 (N_3243,N_1874,N_1896);
nand U3244 (N_3244,N_2412,N_1838);
xnor U3245 (N_3245,N_1614,N_2071);
xor U3246 (N_3246,N_2597,N_2755);
or U3247 (N_3247,N_2615,N_2981);
or U3248 (N_3248,N_2418,N_2999);
xnor U3249 (N_3249,N_2647,N_2696);
nor U3250 (N_3250,N_2674,N_2887);
and U3251 (N_3251,N_1745,N_2399);
and U3252 (N_3252,N_2813,N_1570);
or U3253 (N_3253,N_2964,N_2502);
or U3254 (N_3254,N_2941,N_1923);
or U3255 (N_3255,N_2967,N_2876);
and U3256 (N_3256,N_1639,N_1796);
xor U3257 (N_3257,N_2038,N_2628);
or U3258 (N_3258,N_1894,N_1943);
or U3259 (N_3259,N_1773,N_1800);
nand U3260 (N_3260,N_2798,N_1946);
nor U3261 (N_3261,N_1728,N_1534);
nand U3262 (N_3262,N_1702,N_1866);
and U3263 (N_3263,N_2655,N_2076);
and U3264 (N_3264,N_1593,N_2511);
nor U3265 (N_3265,N_2003,N_2247);
and U3266 (N_3266,N_2439,N_1644);
nor U3267 (N_3267,N_2119,N_1624);
nand U3268 (N_3268,N_2559,N_2130);
nor U3269 (N_3269,N_1715,N_1719);
nor U3270 (N_3270,N_2455,N_1883);
or U3271 (N_3271,N_2225,N_1640);
xnor U3272 (N_3272,N_1903,N_1642);
xnor U3273 (N_3273,N_2396,N_1517);
or U3274 (N_3274,N_2699,N_2103);
or U3275 (N_3275,N_2184,N_2273);
nor U3276 (N_3276,N_2467,N_2894);
or U3277 (N_3277,N_1810,N_2721);
nand U3278 (N_3278,N_1853,N_2142);
xor U3279 (N_3279,N_1816,N_2539);
or U3280 (N_3280,N_2896,N_1905);
nor U3281 (N_3281,N_2265,N_2626);
xnor U3282 (N_3282,N_2974,N_1618);
and U3283 (N_3283,N_2342,N_2565);
xor U3284 (N_3284,N_1961,N_2697);
nand U3285 (N_3285,N_2345,N_2178);
and U3286 (N_3286,N_2931,N_2921);
xor U3287 (N_3287,N_2688,N_2979);
nor U3288 (N_3288,N_1580,N_2405);
nand U3289 (N_3289,N_2940,N_1722);
nor U3290 (N_3290,N_2367,N_1542);
or U3291 (N_3291,N_1912,N_2717);
nand U3292 (N_3292,N_2073,N_2368);
nor U3293 (N_3293,N_2854,N_2113);
nor U3294 (N_3294,N_2666,N_2900);
nor U3295 (N_3295,N_2739,N_2971);
or U3296 (N_3296,N_1931,N_2349);
and U3297 (N_3297,N_1860,N_2842);
and U3298 (N_3298,N_1901,N_2242);
nand U3299 (N_3299,N_2945,N_1736);
xor U3300 (N_3300,N_2025,N_2617);
or U3301 (N_3301,N_2892,N_1607);
nand U3302 (N_3302,N_2445,N_1851);
nand U3303 (N_3303,N_2532,N_1945);
nor U3304 (N_3304,N_2882,N_1989);
nand U3305 (N_3305,N_1681,N_2390);
nand U3306 (N_3306,N_1948,N_2950);
or U3307 (N_3307,N_1678,N_2656);
nand U3308 (N_3308,N_1817,N_1667);
nor U3309 (N_3309,N_1916,N_1994);
nor U3310 (N_3310,N_2549,N_2391);
and U3311 (N_3311,N_2070,N_2548);
nor U3312 (N_3312,N_1625,N_2871);
nand U3313 (N_3313,N_1926,N_2352);
xnor U3314 (N_3314,N_2098,N_2213);
nor U3315 (N_3315,N_2088,N_2245);
or U3316 (N_3316,N_1870,N_2540);
nand U3317 (N_3317,N_1572,N_2923);
or U3318 (N_3318,N_2794,N_2595);
nor U3319 (N_3319,N_2221,N_2660);
and U3320 (N_3320,N_1778,N_2806);
xnor U3321 (N_3321,N_1981,N_1684);
nor U3322 (N_3322,N_2181,N_2324);
or U3323 (N_3323,N_1659,N_2880);
nand U3324 (N_3324,N_1999,N_2925);
and U3325 (N_3325,N_2218,N_2074);
nand U3326 (N_3326,N_2516,N_1584);
and U3327 (N_3327,N_1872,N_2298);
nand U3328 (N_3328,N_2710,N_2645);
and U3329 (N_3329,N_1611,N_2805);
and U3330 (N_3330,N_2397,N_1608);
or U3331 (N_3331,N_2963,N_2730);
xnor U3332 (N_3332,N_1919,N_1503);
xor U3333 (N_3333,N_2110,N_2765);
nand U3334 (N_3334,N_1982,N_2011);
nor U3335 (N_3335,N_2122,N_1964);
nor U3336 (N_3336,N_2718,N_2156);
and U3337 (N_3337,N_1897,N_2822);
and U3338 (N_3338,N_2668,N_2408);
nand U3339 (N_3339,N_1533,N_1852);
nor U3340 (N_3340,N_2913,N_1524);
nor U3341 (N_3341,N_2441,N_1734);
or U3342 (N_3342,N_1791,N_2750);
xnor U3343 (N_3343,N_1752,N_2951);
xor U3344 (N_3344,N_1647,N_1933);
nand U3345 (N_3345,N_1833,N_2157);
xnor U3346 (N_3346,N_2953,N_2500);
or U3347 (N_3347,N_2029,N_1599);
nand U3348 (N_3348,N_2285,N_2648);
nand U3349 (N_3349,N_2470,N_1804);
nand U3350 (N_3350,N_1566,N_2942);
and U3351 (N_3351,N_2125,N_1739);
nand U3352 (N_3352,N_1609,N_2223);
or U3353 (N_3353,N_2601,N_2897);
nor U3354 (N_3354,N_1656,N_1598);
nor U3355 (N_3355,N_2436,N_1634);
or U3356 (N_3356,N_2090,N_2291);
and U3357 (N_3357,N_1985,N_2267);
xor U3358 (N_3358,N_2727,N_1501);
nor U3359 (N_3359,N_2677,N_2206);
nand U3360 (N_3360,N_2487,N_2616);
nand U3361 (N_3361,N_2744,N_2687);
xnor U3362 (N_3362,N_2938,N_2478);
nor U3363 (N_3363,N_1525,N_1587);
or U3364 (N_3364,N_1551,N_2188);
or U3365 (N_3365,N_1675,N_1679);
and U3366 (N_3366,N_1709,N_1844);
nand U3367 (N_3367,N_2586,N_2671);
and U3368 (N_3368,N_1676,N_2168);
and U3369 (N_3369,N_1921,N_2514);
nor U3370 (N_3370,N_1777,N_2386);
and U3371 (N_3371,N_2123,N_2400);
nor U3372 (N_3372,N_1557,N_2761);
or U3373 (N_3373,N_1808,N_2274);
nand U3374 (N_3374,N_2911,N_1723);
xor U3375 (N_3375,N_2874,N_1708);
and U3376 (N_3376,N_2450,N_2975);
nor U3377 (N_3377,N_2958,N_2251);
nor U3378 (N_3378,N_1865,N_2105);
or U3379 (N_3379,N_2055,N_2686);
xnor U3380 (N_3380,N_1990,N_1603);
xor U3381 (N_3381,N_1516,N_1937);
or U3382 (N_3382,N_1987,N_1664);
nor U3383 (N_3383,N_2510,N_2776);
nand U3384 (N_3384,N_2927,N_2592);
nand U3385 (N_3385,N_2327,N_1960);
or U3386 (N_3386,N_2093,N_2040);
nor U3387 (N_3387,N_1888,N_2442);
xor U3388 (N_3388,N_1606,N_2464);
or U3389 (N_3389,N_1913,N_1502);
xor U3390 (N_3390,N_2493,N_2928);
xor U3391 (N_3391,N_1871,N_2380);
nand U3392 (N_3392,N_2069,N_1836);
xor U3393 (N_3393,N_2537,N_2809);
or U3394 (N_3394,N_2134,N_2313);
or U3395 (N_3395,N_2629,N_1789);
xnor U3396 (N_3396,N_2132,N_1924);
nand U3397 (N_3397,N_2203,N_2200);
xnor U3398 (N_3398,N_2733,N_2304);
and U3399 (N_3399,N_2453,N_2917);
xor U3400 (N_3400,N_2451,N_2576);
nand U3401 (N_3401,N_1867,N_1877);
and U3402 (N_3402,N_2048,N_1743);
nand U3403 (N_3403,N_2086,N_2358);
and U3404 (N_3404,N_2708,N_1571);
nor U3405 (N_3405,N_2332,N_2572);
xor U3406 (N_3406,N_1548,N_2800);
nor U3407 (N_3407,N_1509,N_2187);
nor U3408 (N_3408,N_1967,N_2711);
or U3409 (N_3409,N_2144,N_1558);
nor U3410 (N_3410,N_2815,N_2957);
and U3411 (N_3411,N_2949,N_2829);
and U3412 (N_3412,N_2295,N_2266);
xor U3413 (N_3413,N_2012,N_2052);
or U3414 (N_3414,N_2248,N_2432);
nor U3415 (N_3415,N_2639,N_1645);
nand U3416 (N_3416,N_2995,N_2759);
or U3417 (N_3417,N_2062,N_2955);
xnor U3418 (N_3418,N_1628,N_2935);
nand U3419 (N_3419,N_2147,N_2546);
and U3420 (N_3420,N_2507,N_1674);
and U3421 (N_3421,N_2359,N_2419);
or U3422 (N_3422,N_2301,N_2588);
or U3423 (N_3423,N_2006,N_2819);
nand U3424 (N_3424,N_2347,N_2496);
nor U3425 (N_3425,N_2394,N_2406);
or U3426 (N_3426,N_2622,N_2280);
and U3427 (N_3427,N_2826,N_1878);
xor U3428 (N_3428,N_2969,N_2497);
xor U3429 (N_3429,N_1755,N_2531);
or U3430 (N_3430,N_2584,N_2484);
or U3431 (N_3431,N_1689,N_2194);
xnor U3432 (N_3432,N_2599,N_1555);
or U3433 (N_3433,N_2348,N_1532);
and U3434 (N_3434,N_1995,N_2387);
or U3435 (N_3435,N_2535,N_2659);
and U3436 (N_3436,N_1556,N_2509);
and U3437 (N_3437,N_2638,N_2246);
xnor U3438 (N_3438,N_2075,N_1928);
and U3439 (N_3439,N_1879,N_1850);
or U3440 (N_3440,N_1797,N_2520);
or U3441 (N_3441,N_1809,N_2864);
or U3442 (N_3442,N_1685,N_2019);
and U3443 (N_3443,N_2344,N_1760);
nor U3444 (N_3444,N_2065,N_2832);
and U3445 (N_3445,N_2136,N_2422);
or U3446 (N_3446,N_2977,N_2663);
nor U3447 (N_3447,N_2614,N_2676);
xor U3448 (N_3448,N_2127,N_2556);
and U3449 (N_3449,N_2799,N_1670);
and U3450 (N_3450,N_2504,N_1537);
nand U3451 (N_3451,N_2631,N_1754);
nor U3452 (N_3452,N_2457,N_1846);
or U3453 (N_3453,N_2662,N_1610);
or U3454 (N_3454,N_2817,N_1840);
and U3455 (N_3455,N_2590,N_2850);
and U3456 (N_3456,N_2980,N_2293);
or U3457 (N_3457,N_2311,N_2033);
or U3458 (N_3458,N_2642,N_1918);
nor U3459 (N_3459,N_1834,N_2145);
nor U3460 (N_3460,N_2780,N_2284);
or U3461 (N_3461,N_2329,N_2849);
nand U3462 (N_3462,N_2377,N_1662);
and U3463 (N_3463,N_2848,N_2785);
nand U3464 (N_3464,N_2286,N_2465);
or U3465 (N_3465,N_2841,N_1911);
or U3466 (N_3466,N_2424,N_2477);
nor U3467 (N_3467,N_1692,N_2403);
nand U3468 (N_3468,N_1848,N_2946);
xor U3469 (N_3469,N_1781,N_2287);
or U3470 (N_3470,N_2296,N_2044);
xor U3471 (N_3471,N_1683,N_2908);
nor U3472 (N_3472,N_2609,N_2715);
nor U3473 (N_3473,N_2742,N_1522);
and U3474 (N_3474,N_2834,N_2350);
nand U3475 (N_3475,N_2260,N_2080);
nor U3476 (N_3476,N_2322,N_1972);
xor U3477 (N_3477,N_1801,N_1997);
nor U3478 (N_3478,N_2083,N_2448);
xor U3479 (N_3479,N_2207,N_2192);
or U3480 (N_3480,N_2416,N_1727);
or U3481 (N_3481,N_2564,N_2561);
or U3482 (N_3482,N_1655,N_2479);
nor U3483 (N_3483,N_2581,N_1526);
nand U3484 (N_3484,N_1991,N_2833);
nand U3485 (N_3485,N_2681,N_2929);
nor U3486 (N_3486,N_2512,N_2056);
nor U3487 (N_3487,N_2508,N_1701);
and U3488 (N_3488,N_2312,N_2627);
xnor U3489 (N_3489,N_1564,N_2619);
nor U3490 (N_3490,N_2036,N_2984);
nor U3491 (N_3491,N_2936,N_1993);
nand U3492 (N_3492,N_1612,N_2909);
and U3493 (N_3493,N_1596,N_1600);
or U3494 (N_3494,N_2547,N_2004);
and U3495 (N_3495,N_2318,N_2382);
nor U3496 (N_3496,N_1730,N_2930);
and U3497 (N_3497,N_2978,N_1831);
nor U3498 (N_3498,N_1630,N_2918);
nand U3499 (N_3499,N_2423,N_2374);
nand U3500 (N_3500,N_2797,N_1771);
xnor U3501 (N_3501,N_1854,N_2414);
xnor U3502 (N_3502,N_1910,N_2870);
nor U3503 (N_3503,N_1765,N_2637);
or U3504 (N_3504,N_1696,N_2521);
nor U3505 (N_3505,N_2910,N_1976);
or U3506 (N_3506,N_2435,N_2611);
nand U3507 (N_3507,N_1744,N_2081);
and U3508 (N_3508,N_2735,N_1784);
and U3509 (N_3509,N_1538,N_2636);
nand U3510 (N_3510,N_1794,N_1759);
xnor U3511 (N_3511,N_2726,N_1576);
or U3512 (N_3512,N_2294,N_2395);
nor U3513 (N_3513,N_1849,N_2109);
nor U3514 (N_3514,N_1592,N_2672);
nor U3515 (N_3515,N_1583,N_2693);
and U3516 (N_3516,N_2022,N_2174);
or U3517 (N_3517,N_2680,N_1547);
nor U3518 (N_3518,N_2720,N_2063);
nor U3519 (N_3519,N_2551,N_1619);
xor U3520 (N_3520,N_1549,N_2289);
xnor U3521 (N_3521,N_2258,N_1651);
xnor U3522 (N_3522,N_2279,N_2131);
and U3523 (N_3523,N_2991,N_2278);
xor U3524 (N_3524,N_1805,N_2446);
or U3525 (N_3525,N_2483,N_1540);
xor U3526 (N_3526,N_2212,N_2290);
or U3527 (N_3527,N_1753,N_1776);
nand U3528 (N_3528,N_2722,N_1688);
xnor U3529 (N_3529,N_2873,N_2008);
nor U3530 (N_3530,N_1998,N_1691);
or U3531 (N_3531,N_2058,N_1977);
and U3532 (N_3532,N_2550,N_1605);
nor U3533 (N_3533,N_2034,N_2740);
xor U3534 (N_3534,N_2129,N_1767);
and U3535 (N_3535,N_2256,N_2766);
nand U3536 (N_3536,N_2309,N_2625);
or U3537 (N_3537,N_2222,N_1646);
nor U3538 (N_3538,N_1904,N_2972);
xor U3539 (N_3539,N_2346,N_2401);
or U3540 (N_3540,N_1687,N_2682);
nand U3541 (N_3541,N_1957,N_2398);
nand U3542 (N_3542,N_2491,N_2427);
and U3543 (N_3543,N_1590,N_2692);
and U3544 (N_3544,N_2480,N_2096);
nand U3545 (N_3545,N_2646,N_1758);
nand U3546 (N_3546,N_2420,N_1802);
xnor U3547 (N_3547,N_1505,N_1963);
nor U3548 (N_3548,N_2355,N_2190);
xor U3549 (N_3549,N_1814,N_2255);
xor U3550 (N_3550,N_1837,N_2684);
nand U3551 (N_3551,N_1588,N_2202);
and U3552 (N_3552,N_2219,N_2701);
xnor U3553 (N_3553,N_2685,N_2707);
nand U3554 (N_3554,N_1780,N_2743);
or U3555 (N_3555,N_2583,N_2013);
nor U3556 (N_3556,N_2383,N_2902);
or U3557 (N_3557,N_1671,N_2879);
nand U3558 (N_3558,N_1959,N_2392);
xor U3559 (N_3559,N_2336,N_1968);
nand U3560 (N_3560,N_1714,N_2948);
and U3561 (N_3561,N_1661,N_1669);
or U3562 (N_3562,N_1988,N_2495);
nand U3563 (N_3563,N_1782,N_2644);
xor U3564 (N_3564,N_2172,N_2820);
nand U3565 (N_3565,N_1812,N_1756);
nand U3566 (N_3566,N_2198,N_2305);
nand U3567 (N_3567,N_2292,N_2032);
and U3568 (N_3568,N_2916,N_2283);
nand U3569 (N_3569,N_2326,N_2101);
nand U3570 (N_3570,N_1922,N_2476);
or U3571 (N_3571,N_2177,N_1519);
nor U3572 (N_3572,N_2385,N_2553);
nor U3573 (N_3573,N_2937,N_2215);
and U3574 (N_3574,N_2541,N_1955);
xnor U3575 (N_3575,N_1746,N_2216);
nor U3576 (N_3576,N_1951,N_2779);
or U3577 (N_3577,N_2230,N_1531);
nor U3578 (N_3578,N_1763,N_2444);
or U3579 (N_3579,N_1677,N_1546);
xnor U3580 (N_3580,N_2922,N_1942);
nand U3581 (N_3581,N_2904,N_2824);
nor U3582 (N_3582,N_2460,N_2328);
and U3583 (N_3583,N_2756,N_2729);
and U3584 (N_3584,N_1749,N_1724);
and U3585 (N_3585,N_1579,N_2954);
or U3586 (N_3586,N_2807,N_2724);
nor U3587 (N_3587,N_2830,N_2428);
and U3588 (N_3588,N_1858,N_1512);
xnor U3589 (N_3589,N_2751,N_2769);
xnor U3590 (N_3590,N_1892,N_2189);
and U3591 (N_3591,N_2276,N_1798);
xor U3592 (N_3592,N_1699,N_2235);
or U3593 (N_3593,N_2243,N_1811);
nor U3594 (N_3594,N_2650,N_1528);
xnor U3595 (N_3595,N_2774,N_2582);
nor U3596 (N_3596,N_2563,N_2670);
xor U3597 (N_3597,N_1954,N_2066);
nand U3598 (N_3598,N_2092,N_2170);
and U3599 (N_3599,N_2658,N_2903);
nand U3600 (N_3600,N_2366,N_1694);
xor U3601 (N_3601,N_1935,N_2217);
xnor U3602 (N_3602,N_2775,N_1996);
or U3603 (N_3603,N_1545,N_2973);
nand U3604 (N_3604,N_2272,N_2035);
nand U3605 (N_3605,N_1806,N_1707);
or U3606 (N_3606,N_2120,N_1622);
nand U3607 (N_3607,N_2747,N_2580);
nor U3608 (N_3608,N_1690,N_1953);
or U3609 (N_3609,N_2372,N_2858);
nand U3610 (N_3610,N_1979,N_2430);
xor U3611 (N_3611,N_2297,N_2106);
xnor U3612 (N_3612,N_2893,N_1917);
nand U3613 (N_3613,N_1898,N_2851);
xor U3614 (N_3614,N_1906,N_1927);
and U3615 (N_3615,N_2186,N_2634);
nand U3616 (N_3616,N_2100,N_1971);
and U3617 (N_3617,N_2023,N_1930);
and U3618 (N_3618,N_1649,N_2679);
nand U3619 (N_3619,N_1735,N_2115);
and U3620 (N_3620,N_2362,N_1508);
or U3621 (N_3621,N_2789,N_2150);
or U3622 (N_3622,N_2812,N_2196);
nand U3623 (N_3623,N_2673,N_1828);
nand U3624 (N_3624,N_2363,N_2803);
nand U3625 (N_3625,N_2956,N_2788);
xor U3626 (N_3626,N_1915,N_2375);
nand U3627 (N_3627,N_2543,N_2209);
nor U3628 (N_3628,N_2160,N_2407);
xor U3629 (N_3629,N_2486,N_1830);
or U3630 (N_3630,N_2836,N_2792);
or U3631 (N_3631,N_2932,N_2107);
nand U3632 (N_3632,N_2593,N_1934);
xor U3633 (N_3633,N_2630,N_2529);
nand U3634 (N_3634,N_1792,N_2410);
nand U3635 (N_3635,N_2288,N_2821);
nand U3636 (N_3636,N_1841,N_2361);
xor U3637 (N_3637,N_1839,N_2425);
or U3638 (N_3638,N_2371,N_2515);
xor U3639 (N_3639,N_1863,N_2133);
and U3640 (N_3640,N_2840,N_2149);
or U3641 (N_3641,N_1523,N_2270);
or U3642 (N_3642,N_2236,N_2853);
or U3643 (N_3643,N_2485,N_2461);
nand U3644 (N_3644,N_1889,N_1733);
nor U3645 (N_3645,N_2117,N_1820);
nor U3646 (N_3646,N_2669,N_2952);
nor U3647 (N_3647,N_1638,N_2567);
and U3648 (N_3648,N_1761,N_2818);
xnor U3649 (N_3649,N_1939,N_1514);
nor U3650 (N_3650,N_1969,N_2741);
nor U3651 (N_3651,N_1521,N_2598);
or U3652 (N_3652,N_2275,N_2020);
nor U3653 (N_3653,N_2334,N_1738);
xor U3654 (N_3654,N_2128,N_2610);
xor U3655 (N_3655,N_2713,N_1713);
or U3656 (N_3656,N_2560,N_2863);
nor U3657 (N_3657,N_1835,N_2748);
or U3658 (N_3658,N_2179,N_2454);
xnor U3659 (N_3659,N_2153,N_2875);
and U3660 (N_3660,N_2211,N_2839);
nand U3661 (N_3661,N_1627,N_2506);
nand U3662 (N_3662,N_1589,N_2252);
nand U3663 (N_3663,N_2271,N_1958);
and U3664 (N_3664,N_2933,N_2513);
nand U3665 (N_3665,N_1527,N_2810);
nand U3666 (N_3666,N_2859,N_2857);
nor U3667 (N_3667,N_1822,N_2907);
and U3668 (N_3668,N_1513,N_2704);
nand U3669 (N_3669,N_2343,N_1543);
nor U3670 (N_3670,N_2238,N_1650);
xor U3671 (N_3671,N_1769,N_2458);
and U3672 (N_3672,N_2552,N_2016);
or U3673 (N_3673,N_1826,N_2471);
or U3674 (N_3674,N_2714,N_2678);
xnor U3675 (N_3675,N_2143,N_1597);
xnor U3676 (N_3676,N_2885,N_2338);
xor U3677 (N_3677,N_1544,N_2353);
and U3678 (N_3678,N_2161,N_2926);
xnor U3679 (N_3679,N_2310,N_2786);
xor U3680 (N_3680,N_1775,N_2811);
and U3681 (N_3681,N_2068,N_2331);
or U3682 (N_3682,N_2706,N_1859);
and U3683 (N_3683,N_2426,N_2364);
nor U3684 (N_3684,N_1666,N_2816);
nor U3685 (N_3685,N_1936,N_2064);
nand U3686 (N_3686,N_1504,N_1740);
and U3687 (N_3687,N_1643,N_1823);
and U3688 (N_3688,N_2135,N_2772);
xor U3689 (N_3689,N_1940,N_2176);
nor U3690 (N_3690,N_2762,N_1574);
and U3691 (N_3691,N_1891,N_2651);
and U3692 (N_3692,N_1529,N_2241);
or U3693 (N_3693,N_1682,N_1907);
nor U3694 (N_3694,N_1862,N_2037);
and U3695 (N_3695,N_2612,N_2197);
or U3696 (N_3696,N_2749,N_2845);
and U3697 (N_3697,N_2158,N_2320);
nand U3698 (N_3698,N_2388,N_2306);
nand U3699 (N_3699,N_2901,N_1772);
nor U3700 (N_3700,N_2183,N_2591);
and U3701 (N_3701,N_2299,N_1569);
nand U3702 (N_3702,N_2024,N_2796);
and U3703 (N_3703,N_2018,N_2208);
xor U3704 (N_3704,N_2613,N_2057);
nand U3705 (N_3705,N_2554,N_2568);
nor U3706 (N_3706,N_2409,N_2570);
nor U3707 (N_3707,N_1641,N_2126);
nor U3708 (N_3708,N_2571,N_2233);
nand U3709 (N_3709,N_2224,N_2654);
nor U3710 (N_3710,N_1986,N_2606);
nand U3711 (N_3711,N_2764,N_2835);
nor U3712 (N_3712,N_2250,N_1785);
nand U3713 (N_3713,N_1950,N_2097);
nand U3714 (N_3714,N_2165,N_1783);
nand U3715 (N_3715,N_1635,N_1952);
nand U3716 (N_3716,N_1654,N_2944);
nand U3717 (N_3717,N_1621,N_2002);
nand U3718 (N_3718,N_2099,N_2303);
nand U3719 (N_3719,N_2229,N_1768);
nand U3720 (N_3720,N_2314,N_2095);
or U3721 (N_3721,N_1536,N_2939);
nand U3722 (N_3722,N_2041,N_2782);
nor U3723 (N_3723,N_1704,N_1770);
nand U3724 (N_3724,N_2417,N_1788);
xnor U3725 (N_3725,N_2558,N_2527);
and U3726 (N_3726,N_1700,N_2777);
nand U3727 (N_3727,N_2519,N_1938);
and U3728 (N_3728,N_2878,N_2061);
xor U3729 (N_3729,N_2239,N_1762);
and U3730 (N_3730,N_2745,N_2661);
xnor U3731 (N_3731,N_2137,N_2316);
nor U3732 (N_3732,N_1680,N_2308);
or U3733 (N_3733,N_2393,N_1562);
xnor U3734 (N_3734,N_2992,N_2557);
nand U3735 (N_3735,N_2734,N_2573);
xor U3736 (N_3736,N_1803,N_2481);
nand U3737 (N_3737,N_1885,N_1766);
and U3738 (N_3738,N_2389,N_2193);
and U3739 (N_3739,N_2139,N_2970);
nand U3740 (N_3740,N_1616,N_2438);
nor U3741 (N_3741,N_1703,N_1575);
xor U3742 (N_3742,N_2524,N_1786);
or U3743 (N_3743,N_2861,N_2536);
and U3744 (N_3744,N_1705,N_2085);
nor U3745 (N_3745,N_1563,N_2781);
and U3746 (N_3746,N_2889,N_1585);
xor U3747 (N_3747,N_2635,N_2141);
nor U3748 (N_3748,N_1721,N_2492);
xnor U3749 (N_3749,N_2072,N_2319);
nand U3750 (N_3750,N_2343,N_2592);
xor U3751 (N_3751,N_2453,N_1887);
or U3752 (N_3752,N_2306,N_1938);
or U3753 (N_3753,N_2955,N_1605);
or U3754 (N_3754,N_2313,N_2776);
and U3755 (N_3755,N_2840,N_2922);
and U3756 (N_3756,N_2823,N_2016);
or U3757 (N_3757,N_2601,N_2171);
xor U3758 (N_3758,N_2193,N_1690);
xnor U3759 (N_3759,N_1676,N_2833);
nor U3760 (N_3760,N_2581,N_1957);
and U3761 (N_3761,N_1765,N_1788);
and U3762 (N_3762,N_2181,N_1805);
nand U3763 (N_3763,N_2809,N_2850);
and U3764 (N_3764,N_2100,N_2696);
or U3765 (N_3765,N_1979,N_2529);
or U3766 (N_3766,N_2392,N_1917);
xnor U3767 (N_3767,N_1789,N_2862);
or U3768 (N_3768,N_1704,N_2860);
nor U3769 (N_3769,N_2372,N_2714);
xor U3770 (N_3770,N_1911,N_1867);
and U3771 (N_3771,N_2170,N_2357);
or U3772 (N_3772,N_2605,N_2805);
and U3773 (N_3773,N_1560,N_2182);
and U3774 (N_3774,N_1926,N_2144);
nand U3775 (N_3775,N_2225,N_2822);
or U3776 (N_3776,N_2107,N_1686);
and U3777 (N_3777,N_1793,N_1548);
xnor U3778 (N_3778,N_2548,N_2750);
nand U3779 (N_3779,N_2713,N_1972);
nand U3780 (N_3780,N_2881,N_2984);
and U3781 (N_3781,N_1678,N_2567);
nand U3782 (N_3782,N_1666,N_2085);
nand U3783 (N_3783,N_2146,N_2516);
and U3784 (N_3784,N_1606,N_2998);
and U3785 (N_3785,N_2413,N_1649);
nand U3786 (N_3786,N_2119,N_1941);
nand U3787 (N_3787,N_2154,N_2910);
and U3788 (N_3788,N_1921,N_2973);
or U3789 (N_3789,N_2513,N_1989);
or U3790 (N_3790,N_1519,N_1824);
xnor U3791 (N_3791,N_2991,N_2514);
or U3792 (N_3792,N_2673,N_2359);
xor U3793 (N_3793,N_1860,N_2569);
and U3794 (N_3794,N_2892,N_2354);
xnor U3795 (N_3795,N_2046,N_1599);
nor U3796 (N_3796,N_1844,N_2095);
and U3797 (N_3797,N_2081,N_2548);
nor U3798 (N_3798,N_2201,N_2066);
nor U3799 (N_3799,N_2847,N_2536);
or U3800 (N_3800,N_1980,N_2466);
or U3801 (N_3801,N_1678,N_1773);
nand U3802 (N_3802,N_2208,N_2140);
and U3803 (N_3803,N_2827,N_1585);
and U3804 (N_3804,N_1646,N_2795);
and U3805 (N_3805,N_1582,N_2760);
nor U3806 (N_3806,N_2298,N_2563);
or U3807 (N_3807,N_1754,N_1833);
and U3808 (N_3808,N_2951,N_1785);
xnor U3809 (N_3809,N_1964,N_2618);
xnor U3810 (N_3810,N_2709,N_1910);
and U3811 (N_3811,N_2797,N_2312);
nand U3812 (N_3812,N_2053,N_2046);
or U3813 (N_3813,N_2062,N_2234);
and U3814 (N_3814,N_2966,N_2150);
and U3815 (N_3815,N_1717,N_1557);
nor U3816 (N_3816,N_1635,N_1790);
and U3817 (N_3817,N_2664,N_2752);
and U3818 (N_3818,N_2829,N_2176);
xnor U3819 (N_3819,N_2628,N_2275);
xnor U3820 (N_3820,N_2744,N_1565);
nand U3821 (N_3821,N_2612,N_2619);
nand U3822 (N_3822,N_2504,N_2539);
or U3823 (N_3823,N_2176,N_2377);
and U3824 (N_3824,N_1703,N_1878);
nor U3825 (N_3825,N_2943,N_2420);
and U3826 (N_3826,N_2757,N_2297);
nor U3827 (N_3827,N_2827,N_1991);
nor U3828 (N_3828,N_2082,N_1914);
nor U3829 (N_3829,N_1789,N_1676);
nor U3830 (N_3830,N_2237,N_2144);
nor U3831 (N_3831,N_2169,N_2898);
nand U3832 (N_3832,N_2041,N_1636);
nor U3833 (N_3833,N_1801,N_2787);
and U3834 (N_3834,N_1501,N_2796);
or U3835 (N_3835,N_1853,N_1842);
or U3836 (N_3836,N_2702,N_2653);
xnor U3837 (N_3837,N_1505,N_2710);
xor U3838 (N_3838,N_2490,N_2778);
and U3839 (N_3839,N_2059,N_2946);
nor U3840 (N_3840,N_1712,N_2546);
nand U3841 (N_3841,N_2762,N_2938);
or U3842 (N_3842,N_2731,N_1917);
nor U3843 (N_3843,N_2988,N_2961);
and U3844 (N_3844,N_1884,N_2538);
xor U3845 (N_3845,N_2567,N_2241);
nand U3846 (N_3846,N_2864,N_2734);
nor U3847 (N_3847,N_1884,N_2065);
nand U3848 (N_3848,N_1699,N_1612);
nand U3849 (N_3849,N_1618,N_1612);
or U3850 (N_3850,N_2282,N_2792);
nand U3851 (N_3851,N_2733,N_2751);
nand U3852 (N_3852,N_2376,N_1547);
and U3853 (N_3853,N_2749,N_1965);
and U3854 (N_3854,N_2691,N_1707);
nor U3855 (N_3855,N_2688,N_1949);
nand U3856 (N_3856,N_2682,N_2177);
nor U3857 (N_3857,N_1567,N_2218);
nand U3858 (N_3858,N_2838,N_1930);
xor U3859 (N_3859,N_2224,N_1987);
and U3860 (N_3860,N_2555,N_2341);
xnor U3861 (N_3861,N_2404,N_2927);
nor U3862 (N_3862,N_2018,N_1816);
or U3863 (N_3863,N_1937,N_1597);
nor U3864 (N_3864,N_2291,N_1580);
nor U3865 (N_3865,N_2035,N_2888);
nand U3866 (N_3866,N_2300,N_1838);
or U3867 (N_3867,N_2670,N_2807);
or U3868 (N_3868,N_2127,N_1795);
xnor U3869 (N_3869,N_2260,N_2801);
xnor U3870 (N_3870,N_2724,N_2191);
or U3871 (N_3871,N_2951,N_1527);
or U3872 (N_3872,N_2084,N_1661);
nand U3873 (N_3873,N_1940,N_2407);
nand U3874 (N_3874,N_1843,N_2724);
and U3875 (N_3875,N_2444,N_2871);
nor U3876 (N_3876,N_1879,N_1643);
and U3877 (N_3877,N_1910,N_2959);
nand U3878 (N_3878,N_2601,N_1852);
and U3879 (N_3879,N_2912,N_1553);
or U3880 (N_3880,N_2319,N_2050);
xnor U3881 (N_3881,N_1647,N_2246);
xnor U3882 (N_3882,N_2732,N_1531);
nor U3883 (N_3883,N_1785,N_2971);
and U3884 (N_3884,N_2681,N_2304);
and U3885 (N_3885,N_2736,N_2885);
and U3886 (N_3886,N_2274,N_2261);
xnor U3887 (N_3887,N_2013,N_2363);
or U3888 (N_3888,N_2973,N_1615);
and U3889 (N_3889,N_2891,N_1749);
xor U3890 (N_3890,N_2637,N_1864);
nand U3891 (N_3891,N_2384,N_2393);
nor U3892 (N_3892,N_2190,N_2873);
xor U3893 (N_3893,N_2319,N_2647);
nand U3894 (N_3894,N_2133,N_1545);
or U3895 (N_3895,N_2761,N_2754);
nand U3896 (N_3896,N_2611,N_1816);
nand U3897 (N_3897,N_2731,N_2128);
and U3898 (N_3898,N_2280,N_2227);
or U3899 (N_3899,N_2829,N_2246);
xor U3900 (N_3900,N_1793,N_2777);
nand U3901 (N_3901,N_2165,N_1807);
xnor U3902 (N_3902,N_1767,N_2756);
nand U3903 (N_3903,N_2561,N_2997);
nor U3904 (N_3904,N_1746,N_2251);
or U3905 (N_3905,N_2110,N_1908);
nor U3906 (N_3906,N_2596,N_1984);
and U3907 (N_3907,N_1672,N_2380);
nor U3908 (N_3908,N_2811,N_1912);
or U3909 (N_3909,N_1973,N_1658);
or U3910 (N_3910,N_2038,N_2335);
nand U3911 (N_3911,N_2770,N_2552);
and U3912 (N_3912,N_2934,N_1790);
or U3913 (N_3913,N_2576,N_2144);
or U3914 (N_3914,N_1638,N_1747);
and U3915 (N_3915,N_2413,N_2516);
nand U3916 (N_3916,N_2405,N_2289);
nand U3917 (N_3917,N_2165,N_2226);
or U3918 (N_3918,N_2476,N_2143);
xor U3919 (N_3919,N_2549,N_2268);
nand U3920 (N_3920,N_2925,N_2713);
or U3921 (N_3921,N_2977,N_2259);
and U3922 (N_3922,N_1975,N_2073);
or U3923 (N_3923,N_1699,N_2336);
nor U3924 (N_3924,N_1750,N_2891);
and U3925 (N_3925,N_2853,N_2558);
and U3926 (N_3926,N_2598,N_2278);
nand U3927 (N_3927,N_2584,N_2803);
nand U3928 (N_3928,N_1922,N_1966);
nor U3929 (N_3929,N_1982,N_2271);
xnor U3930 (N_3930,N_2724,N_1610);
nand U3931 (N_3931,N_1784,N_1729);
xor U3932 (N_3932,N_1866,N_2509);
xor U3933 (N_3933,N_1911,N_2509);
nor U3934 (N_3934,N_1939,N_2653);
and U3935 (N_3935,N_1800,N_1869);
nor U3936 (N_3936,N_1642,N_1879);
nor U3937 (N_3937,N_1526,N_2161);
xnor U3938 (N_3938,N_2741,N_2165);
xor U3939 (N_3939,N_1513,N_2235);
xor U3940 (N_3940,N_1969,N_2000);
and U3941 (N_3941,N_2667,N_2216);
and U3942 (N_3942,N_1754,N_1823);
xnor U3943 (N_3943,N_2478,N_2791);
nor U3944 (N_3944,N_2371,N_1917);
xor U3945 (N_3945,N_2864,N_2917);
and U3946 (N_3946,N_2729,N_1634);
xor U3947 (N_3947,N_2298,N_2703);
or U3948 (N_3948,N_1550,N_2892);
nor U3949 (N_3949,N_2947,N_2465);
and U3950 (N_3950,N_2130,N_1516);
and U3951 (N_3951,N_2462,N_1862);
nor U3952 (N_3952,N_1500,N_1626);
xnor U3953 (N_3953,N_2274,N_1896);
or U3954 (N_3954,N_2634,N_2098);
xor U3955 (N_3955,N_2738,N_1813);
nand U3956 (N_3956,N_2736,N_1765);
or U3957 (N_3957,N_1769,N_1640);
and U3958 (N_3958,N_2195,N_1614);
nor U3959 (N_3959,N_2879,N_1987);
or U3960 (N_3960,N_2441,N_1931);
and U3961 (N_3961,N_1571,N_2865);
nand U3962 (N_3962,N_2576,N_2777);
or U3963 (N_3963,N_2233,N_1841);
or U3964 (N_3964,N_1994,N_1866);
xnor U3965 (N_3965,N_2423,N_2601);
nand U3966 (N_3966,N_1757,N_1777);
and U3967 (N_3967,N_2522,N_1769);
nor U3968 (N_3968,N_2053,N_2542);
nor U3969 (N_3969,N_2872,N_1907);
nand U3970 (N_3970,N_2765,N_1950);
xnor U3971 (N_3971,N_1713,N_2041);
or U3972 (N_3972,N_2828,N_1758);
and U3973 (N_3973,N_2678,N_2924);
or U3974 (N_3974,N_1842,N_2298);
or U3975 (N_3975,N_1729,N_2287);
nand U3976 (N_3976,N_1900,N_2894);
nand U3977 (N_3977,N_1629,N_2890);
and U3978 (N_3978,N_1643,N_2325);
nand U3979 (N_3979,N_1777,N_2623);
and U3980 (N_3980,N_2611,N_1674);
nor U3981 (N_3981,N_2030,N_1891);
nor U3982 (N_3982,N_2583,N_2666);
nor U3983 (N_3983,N_1736,N_1942);
or U3984 (N_3984,N_2745,N_2801);
xnor U3985 (N_3985,N_1776,N_1692);
or U3986 (N_3986,N_2403,N_2060);
nand U3987 (N_3987,N_1692,N_2096);
xor U3988 (N_3988,N_1582,N_1557);
xnor U3989 (N_3989,N_1839,N_1596);
nor U3990 (N_3990,N_2067,N_2994);
and U3991 (N_3991,N_2551,N_2380);
or U3992 (N_3992,N_1708,N_2835);
nand U3993 (N_3993,N_2230,N_1932);
xor U3994 (N_3994,N_2594,N_1672);
nor U3995 (N_3995,N_2978,N_2557);
nand U3996 (N_3996,N_1901,N_1611);
or U3997 (N_3997,N_2151,N_2614);
nand U3998 (N_3998,N_1887,N_1673);
nor U3999 (N_3999,N_1599,N_1975);
or U4000 (N_4000,N_1527,N_2287);
xnor U4001 (N_4001,N_2189,N_2740);
and U4002 (N_4002,N_2072,N_2111);
xor U4003 (N_4003,N_1525,N_2415);
nand U4004 (N_4004,N_2084,N_2992);
and U4005 (N_4005,N_1849,N_2041);
nand U4006 (N_4006,N_1868,N_2745);
nand U4007 (N_4007,N_1607,N_1927);
and U4008 (N_4008,N_1973,N_2963);
xor U4009 (N_4009,N_2037,N_1542);
or U4010 (N_4010,N_2678,N_2155);
xor U4011 (N_4011,N_1656,N_2560);
xor U4012 (N_4012,N_2105,N_1501);
nand U4013 (N_4013,N_2641,N_2302);
xnor U4014 (N_4014,N_1926,N_2174);
xor U4015 (N_4015,N_2294,N_2732);
or U4016 (N_4016,N_2609,N_2358);
nor U4017 (N_4017,N_2831,N_1543);
and U4018 (N_4018,N_2446,N_2473);
or U4019 (N_4019,N_2430,N_1992);
nor U4020 (N_4020,N_2135,N_1529);
or U4021 (N_4021,N_2346,N_2470);
nor U4022 (N_4022,N_2311,N_2404);
or U4023 (N_4023,N_2070,N_2263);
nand U4024 (N_4024,N_1566,N_2632);
xor U4025 (N_4025,N_2876,N_2373);
nor U4026 (N_4026,N_1725,N_2332);
and U4027 (N_4027,N_2410,N_1591);
and U4028 (N_4028,N_2234,N_2283);
nor U4029 (N_4029,N_1583,N_1900);
nand U4030 (N_4030,N_2107,N_2645);
nand U4031 (N_4031,N_2784,N_2996);
nor U4032 (N_4032,N_2370,N_2755);
nand U4033 (N_4033,N_2413,N_1885);
nor U4034 (N_4034,N_2179,N_2877);
nor U4035 (N_4035,N_2867,N_2759);
nor U4036 (N_4036,N_2649,N_2322);
nor U4037 (N_4037,N_2302,N_2794);
and U4038 (N_4038,N_1514,N_2715);
xnor U4039 (N_4039,N_1853,N_1728);
or U4040 (N_4040,N_2874,N_1739);
nand U4041 (N_4041,N_1768,N_2122);
and U4042 (N_4042,N_2845,N_1572);
or U4043 (N_4043,N_2786,N_1700);
and U4044 (N_4044,N_2571,N_2741);
nand U4045 (N_4045,N_2636,N_2996);
or U4046 (N_4046,N_2362,N_2347);
nand U4047 (N_4047,N_2680,N_2603);
and U4048 (N_4048,N_1942,N_2597);
nand U4049 (N_4049,N_1620,N_2649);
or U4050 (N_4050,N_2382,N_2961);
and U4051 (N_4051,N_2740,N_2432);
nand U4052 (N_4052,N_2911,N_1925);
or U4053 (N_4053,N_2244,N_1590);
or U4054 (N_4054,N_2885,N_2149);
nor U4055 (N_4055,N_1776,N_2385);
xor U4056 (N_4056,N_2791,N_2134);
xnor U4057 (N_4057,N_2468,N_2980);
xor U4058 (N_4058,N_1510,N_2239);
and U4059 (N_4059,N_1611,N_1792);
nand U4060 (N_4060,N_2489,N_1802);
nand U4061 (N_4061,N_1511,N_2417);
and U4062 (N_4062,N_2742,N_2196);
nand U4063 (N_4063,N_2603,N_2377);
or U4064 (N_4064,N_1530,N_2692);
xor U4065 (N_4065,N_1745,N_2977);
and U4066 (N_4066,N_2091,N_1793);
nor U4067 (N_4067,N_1955,N_2354);
nor U4068 (N_4068,N_2378,N_2051);
xor U4069 (N_4069,N_2827,N_2024);
nand U4070 (N_4070,N_1599,N_2400);
or U4071 (N_4071,N_2223,N_2031);
nor U4072 (N_4072,N_2757,N_2414);
nor U4073 (N_4073,N_2922,N_2173);
nor U4074 (N_4074,N_2403,N_1515);
nand U4075 (N_4075,N_1801,N_2601);
and U4076 (N_4076,N_2629,N_2824);
nand U4077 (N_4077,N_1741,N_2315);
or U4078 (N_4078,N_2854,N_1752);
nand U4079 (N_4079,N_2839,N_2869);
xor U4080 (N_4080,N_1904,N_1913);
xnor U4081 (N_4081,N_2912,N_1520);
xnor U4082 (N_4082,N_2523,N_2082);
nand U4083 (N_4083,N_2323,N_2433);
and U4084 (N_4084,N_2181,N_2708);
xor U4085 (N_4085,N_2427,N_2951);
or U4086 (N_4086,N_1836,N_2665);
xor U4087 (N_4087,N_2866,N_2587);
or U4088 (N_4088,N_1969,N_1807);
nor U4089 (N_4089,N_1823,N_2274);
or U4090 (N_4090,N_2234,N_1525);
nand U4091 (N_4091,N_1746,N_2084);
nand U4092 (N_4092,N_2342,N_2205);
nor U4093 (N_4093,N_1682,N_2667);
nand U4094 (N_4094,N_2278,N_2657);
nand U4095 (N_4095,N_1844,N_2376);
nor U4096 (N_4096,N_2927,N_2575);
or U4097 (N_4097,N_1565,N_1799);
nand U4098 (N_4098,N_1600,N_2628);
nand U4099 (N_4099,N_1959,N_2870);
xnor U4100 (N_4100,N_2690,N_2392);
xor U4101 (N_4101,N_2145,N_1711);
xnor U4102 (N_4102,N_2241,N_1662);
nand U4103 (N_4103,N_2985,N_2922);
xor U4104 (N_4104,N_2879,N_2482);
nor U4105 (N_4105,N_1943,N_1651);
or U4106 (N_4106,N_2881,N_1904);
nor U4107 (N_4107,N_2738,N_1522);
nor U4108 (N_4108,N_1671,N_1844);
or U4109 (N_4109,N_2576,N_2711);
and U4110 (N_4110,N_1978,N_2836);
nor U4111 (N_4111,N_2415,N_2759);
and U4112 (N_4112,N_1674,N_1858);
or U4113 (N_4113,N_1640,N_2418);
and U4114 (N_4114,N_2742,N_2461);
or U4115 (N_4115,N_2818,N_2153);
nor U4116 (N_4116,N_1622,N_2083);
or U4117 (N_4117,N_1650,N_1523);
nand U4118 (N_4118,N_2128,N_1888);
or U4119 (N_4119,N_2543,N_2729);
nand U4120 (N_4120,N_1772,N_1922);
and U4121 (N_4121,N_1983,N_2588);
xnor U4122 (N_4122,N_1885,N_2522);
and U4123 (N_4123,N_2470,N_2763);
nor U4124 (N_4124,N_2784,N_2666);
and U4125 (N_4125,N_1820,N_2649);
nor U4126 (N_4126,N_2513,N_1829);
xor U4127 (N_4127,N_2812,N_2833);
xor U4128 (N_4128,N_2327,N_2634);
xnor U4129 (N_4129,N_2210,N_2202);
and U4130 (N_4130,N_2959,N_1948);
and U4131 (N_4131,N_1565,N_2680);
nor U4132 (N_4132,N_2702,N_1873);
nand U4133 (N_4133,N_2651,N_2711);
nand U4134 (N_4134,N_1821,N_1700);
nand U4135 (N_4135,N_1534,N_2749);
nor U4136 (N_4136,N_1714,N_1676);
xor U4137 (N_4137,N_2873,N_1805);
nor U4138 (N_4138,N_2123,N_1779);
and U4139 (N_4139,N_1839,N_1586);
and U4140 (N_4140,N_2229,N_1979);
and U4141 (N_4141,N_1873,N_2648);
and U4142 (N_4142,N_1910,N_1525);
xnor U4143 (N_4143,N_1530,N_2224);
nand U4144 (N_4144,N_2557,N_2556);
xnor U4145 (N_4145,N_2469,N_2286);
xor U4146 (N_4146,N_2158,N_2985);
xnor U4147 (N_4147,N_1881,N_2520);
nor U4148 (N_4148,N_2521,N_2835);
xor U4149 (N_4149,N_2442,N_2160);
or U4150 (N_4150,N_2457,N_1902);
or U4151 (N_4151,N_2911,N_2890);
nor U4152 (N_4152,N_1971,N_2924);
or U4153 (N_4153,N_2481,N_2187);
nand U4154 (N_4154,N_2617,N_1555);
nor U4155 (N_4155,N_2240,N_2328);
nor U4156 (N_4156,N_2842,N_2093);
or U4157 (N_4157,N_2379,N_2099);
xor U4158 (N_4158,N_2358,N_2497);
and U4159 (N_4159,N_2601,N_2348);
nor U4160 (N_4160,N_2297,N_2199);
or U4161 (N_4161,N_2613,N_2794);
xor U4162 (N_4162,N_1818,N_2300);
xor U4163 (N_4163,N_2485,N_2658);
nand U4164 (N_4164,N_2483,N_2929);
nor U4165 (N_4165,N_2409,N_2544);
or U4166 (N_4166,N_1760,N_1606);
xor U4167 (N_4167,N_1689,N_2503);
and U4168 (N_4168,N_2178,N_1538);
nor U4169 (N_4169,N_2578,N_1571);
and U4170 (N_4170,N_1873,N_2520);
and U4171 (N_4171,N_2055,N_2414);
and U4172 (N_4172,N_2079,N_1673);
nand U4173 (N_4173,N_1759,N_1737);
or U4174 (N_4174,N_1629,N_2771);
or U4175 (N_4175,N_1717,N_2584);
and U4176 (N_4176,N_2233,N_2121);
nand U4177 (N_4177,N_1962,N_2109);
xnor U4178 (N_4178,N_1682,N_1728);
and U4179 (N_4179,N_2808,N_2256);
nand U4180 (N_4180,N_2057,N_2285);
or U4181 (N_4181,N_2826,N_1686);
or U4182 (N_4182,N_2042,N_2752);
and U4183 (N_4183,N_1873,N_2856);
nor U4184 (N_4184,N_1885,N_1775);
xor U4185 (N_4185,N_1909,N_2363);
and U4186 (N_4186,N_2341,N_2385);
nand U4187 (N_4187,N_1663,N_2373);
xor U4188 (N_4188,N_2488,N_2179);
and U4189 (N_4189,N_1751,N_2141);
xnor U4190 (N_4190,N_2098,N_2185);
nor U4191 (N_4191,N_2774,N_2923);
or U4192 (N_4192,N_1688,N_1772);
or U4193 (N_4193,N_1654,N_1951);
and U4194 (N_4194,N_2251,N_2735);
or U4195 (N_4195,N_2287,N_2246);
and U4196 (N_4196,N_1826,N_2061);
nor U4197 (N_4197,N_2061,N_2392);
nand U4198 (N_4198,N_2686,N_2345);
nand U4199 (N_4199,N_1559,N_2779);
nor U4200 (N_4200,N_1804,N_2734);
xnor U4201 (N_4201,N_1763,N_1902);
nand U4202 (N_4202,N_2979,N_2273);
nand U4203 (N_4203,N_1772,N_2185);
xnor U4204 (N_4204,N_2934,N_2219);
and U4205 (N_4205,N_1994,N_1908);
nand U4206 (N_4206,N_2790,N_2188);
nand U4207 (N_4207,N_1809,N_1507);
and U4208 (N_4208,N_2403,N_2043);
nor U4209 (N_4209,N_1713,N_2687);
nand U4210 (N_4210,N_2629,N_1981);
xor U4211 (N_4211,N_2976,N_1774);
xor U4212 (N_4212,N_1623,N_2546);
xor U4213 (N_4213,N_2075,N_2368);
nand U4214 (N_4214,N_2322,N_2451);
and U4215 (N_4215,N_1544,N_2430);
xor U4216 (N_4216,N_2921,N_1708);
or U4217 (N_4217,N_2562,N_1632);
and U4218 (N_4218,N_2548,N_2833);
nor U4219 (N_4219,N_2778,N_1938);
nand U4220 (N_4220,N_2562,N_2354);
or U4221 (N_4221,N_2575,N_2825);
nand U4222 (N_4222,N_2148,N_2055);
xor U4223 (N_4223,N_2302,N_2638);
nor U4224 (N_4224,N_2173,N_2135);
and U4225 (N_4225,N_2157,N_1581);
or U4226 (N_4226,N_1936,N_1946);
or U4227 (N_4227,N_2900,N_1962);
nand U4228 (N_4228,N_1834,N_2172);
or U4229 (N_4229,N_2246,N_2121);
and U4230 (N_4230,N_2967,N_2910);
and U4231 (N_4231,N_2539,N_1776);
and U4232 (N_4232,N_1695,N_1765);
or U4233 (N_4233,N_1731,N_1525);
nand U4234 (N_4234,N_2707,N_1561);
nor U4235 (N_4235,N_1518,N_1577);
xor U4236 (N_4236,N_2921,N_2313);
and U4237 (N_4237,N_2458,N_2437);
nand U4238 (N_4238,N_2460,N_1886);
or U4239 (N_4239,N_2491,N_2419);
nand U4240 (N_4240,N_2620,N_1750);
xnor U4241 (N_4241,N_2716,N_2517);
or U4242 (N_4242,N_2734,N_1863);
and U4243 (N_4243,N_1840,N_2214);
xor U4244 (N_4244,N_2627,N_2645);
nand U4245 (N_4245,N_2367,N_2911);
and U4246 (N_4246,N_2164,N_1676);
xnor U4247 (N_4247,N_1634,N_2125);
and U4248 (N_4248,N_2428,N_2660);
and U4249 (N_4249,N_2679,N_2560);
and U4250 (N_4250,N_1720,N_1637);
or U4251 (N_4251,N_2277,N_2660);
xnor U4252 (N_4252,N_2442,N_2547);
or U4253 (N_4253,N_2421,N_2612);
nand U4254 (N_4254,N_1714,N_2910);
xnor U4255 (N_4255,N_2355,N_1684);
nand U4256 (N_4256,N_2197,N_2287);
nand U4257 (N_4257,N_2173,N_1980);
or U4258 (N_4258,N_1586,N_1577);
xor U4259 (N_4259,N_2642,N_2793);
xor U4260 (N_4260,N_1780,N_1637);
and U4261 (N_4261,N_1799,N_2742);
xor U4262 (N_4262,N_1804,N_1761);
nand U4263 (N_4263,N_1809,N_2581);
nor U4264 (N_4264,N_2157,N_2702);
and U4265 (N_4265,N_2109,N_1704);
or U4266 (N_4266,N_2040,N_2920);
xnor U4267 (N_4267,N_2064,N_2765);
xnor U4268 (N_4268,N_1840,N_1849);
xor U4269 (N_4269,N_2917,N_2086);
and U4270 (N_4270,N_1646,N_1616);
nor U4271 (N_4271,N_2389,N_2375);
xor U4272 (N_4272,N_1907,N_1982);
and U4273 (N_4273,N_1677,N_2420);
xor U4274 (N_4274,N_2883,N_2256);
nand U4275 (N_4275,N_2214,N_2817);
xor U4276 (N_4276,N_2917,N_2994);
xnor U4277 (N_4277,N_1595,N_1982);
nand U4278 (N_4278,N_2521,N_2439);
xor U4279 (N_4279,N_2631,N_2522);
nand U4280 (N_4280,N_1914,N_2051);
and U4281 (N_4281,N_2334,N_2231);
or U4282 (N_4282,N_2103,N_2982);
nand U4283 (N_4283,N_2708,N_2704);
nand U4284 (N_4284,N_2491,N_1878);
and U4285 (N_4285,N_1621,N_2865);
and U4286 (N_4286,N_1888,N_2016);
or U4287 (N_4287,N_2919,N_2308);
nand U4288 (N_4288,N_1863,N_1619);
nor U4289 (N_4289,N_2614,N_1951);
xor U4290 (N_4290,N_1901,N_2632);
nor U4291 (N_4291,N_2903,N_2698);
or U4292 (N_4292,N_2384,N_2813);
and U4293 (N_4293,N_2584,N_1789);
xnor U4294 (N_4294,N_2355,N_1947);
or U4295 (N_4295,N_1865,N_2691);
and U4296 (N_4296,N_2229,N_2002);
and U4297 (N_4297,N_2172,N_2220);
or U4298 (N_4298,N_2541,N_2828);
nand U4299 (N_4299,N_1980,N_2498);
or U4300 (N_4300,N_1631,N_1582);
and U4301 (N_4301,N_1539,N_2368);
and U4302 (N_4302,N_2337,N_1816);
nor U4303 (N_4303,N_2070,N_2386);
xor U4304 (N_4304,N_2315,N_1704);
xor U4305 (N_4305,N_2946,N_1841);
nand U4306 (N_4306,N_2258,N_2766);
nor U4307 (N_4307,N_2909,N_2416);
nor U4308 (N_4308,N_2894,N_2832);
or U4309 (N_4309,N_1909,N_2057);
xnor U4310 (N_4310,N_1504,N_1762);
or U4311 (N_4311,N_2940,N_1602);
and U4312 (N_4312,N_1806,N_1556);
and U4313 (N_4313,N_2393,N_2566);
nor U4314 (N_4314,N_1827,N_2889);
nand U4315 (N_4315,N_2213,N_2048);
nand U4316 (N_4316,N_2085,N_2023);
nor U4317 (N_4317,N_1933,N_2500);
xor U4318 (N_4318,N_1783,N_2826);
nand U4319 (N_4319,N_2935,N_2941);
nand U4320 (N_4320,N_2370,N_2045);
or U4321 (N_4321,N_1920,N_1626);
xnor U4322 (N_4322,N_2937,N_2314);
xor U4323 (N_4323,N_2704,N_2049);
and U4324 (N_4324,N_1975,N_1822);
nor U4325 (N_4325,N_2796,N_2897);
xnor U4326 (N_4326,N_2364,N_2301);
xor U4327 (N_4327,N_1947,N_2044);
and U4328 (N_4328,N_2129,N_1810);
nand U4329 (N_4329,N_2416,N_1613);
nand U4330 (N_4330,N_1913,N_2370);
or U4331 (N_4331,N_2928,N_2700);
nor U4332 (N_4332,N_2672,N_1831);
xnor U4333 (N_4333,N_2027,N_1933);
or U4334 (N_4334,N_2029,N_2692);
nand U4335 (N_4335,N_2066,N_2470);
xnor U4336 (N_4336,N_1919,N_2889);
or U4337 (N_4337,N_1987,N_2252);
and U4338 (N_4338,N_1611,N_2736);
nand U4339 (N_4339,N_1957,N_2014);
and U4340 (N_4340,N_2750,N_2835);
nor U4341 (N_4341,N_2313,N_1737);
nor U4342 (N_4342,N_1880,N_2237);
nor U4343 (N_4343,N_1660,N_2747);
or U4344 (N_4344,N_1513,N_2259);
nand U4345 (N_4345,N_1734,N_1601);
and U4346 (N_4346,N_1682,N_2164);
or U4347 (N_4347,N_2442,N_2349);
or U4348 (N_4348,N_2605,N_1632);
and U4349 (N_4349,N_1852,N_2177);
xor U4350 (N_4350,N_2558,N_1860);
nand U4351 (N_4351,N_2969,N_1910);
xnor U4352 (N_4352,N_2034,N_1758);
nand U4353 (N_4353,N_2051,N_2375);
or U4354 (N_4354,N_2234,N_1918);
nor U4355 (N_4355,N_1652,N_2825);
or U4356 (N_4356,N_1602,N_1832);
and U4357 (N_4357,N_2086,N_1591);
nand U4358 (N_4358,N_2221,N_2589);
and U4359 (N_4359,N_2028,N_1729);
nor U4360 (N_4360,N_2868,N_1574);
or U4361 (N_4361,N_2591,N_2182);
xnor U4362 (N_4362,N_2033,N_2070);
or U4363 (N_4363,N_1748,N_2902);
or U4364 (N_4364,N_1691,N_2248);
nor U4365 (N_4365,N_2119,N_2084);
or U4366 (N_4366,N_1654,N_2425);
nor U4367 (N_4367,N_2435,N_2524);
nand U4368 (N_4368,N_2044,N_2992);
nor U4369 (N_4369,N_1683,N_1673);
or U4370 (N_4370,N_2497,N_1983);
nand U4371 (N_4371,N_1608,N_2187);
nor U4372 (N_4372,N_2482,N_2826);
xnor U4373 (N_4373,N_2099,N_2162);
xor U4374 (N_4374,N_2845,N_2596);
or U4375 (N_4375,N_2791,N_2201);
nor U4376 (N_4376,N_1786,N_2989);
and U4377 (N_4377,N_1575,N_2448);
nor U4378 (N_4378,N_2338,N_2908);
or U4379 (N_4379,N_2876,N_2984);
or U4380 (N_4380,N_2002,N_1751);
xnor U4381 (N_4381,N_1799,N_1623);
xor U4382 (N_4382,N_2038,N_2692);
and U4383 (N_4383,N_1900,N_1523);
xnor U4384 (N_4384,N_2090,N_2020);
xnor U4385 (N_4385,N_2818,N_2834);
nand U4386 (N_4386,N_2433,N_2495);
and U4387 (N_4387,N_1688,N_1565);
nor U4388 (N_4388,N_2818,N_2054);
and U4389 (N_4389,N_1823,N_2195);
nor U4390 (N_4390,N_2716,N_1657);
or U4391 (N_4391,N_2551,N_2899);
and U4392 (N_4392,N_1662,N_2673);
or U4393 (N_4393,N_2400,N_2777);
and U4394 (N_4394,N_2174,N_1524);
and U4395 (N_4395,N_2818,N_2001);
and U4396 (N_4396,N_2791,N_2977);
or U4397 (N_4397,N_2844,N_2875);
or U4398 (N_4398,N_2805,N_2986);
and U4399 (N_4399,N_2576,N_2810);
nor U4400 (N_4400,N_2354,N_2269);
or U4401 (N_4401,N_2462,N_2347);
or U4402 (N_4402,N_1640,N_2576);
nand U4403 (N_4403,N_2040,N_1558);
and U4404 (N_4404,N_1619,N_2198);
xor U4405 (N_4405,N_1829,N_2546);
xnor U4406 (N_4406,N_2619,N_2159);
xor U4407 (N_4407,N_2765,N_2108);
xnor U4408 (N_4408,N_1900,N_2892);
nand U4409 (N_4409,N_2506,N_2811);
or U4410 (N_4410,N_2780,N_1770);
or U4411 (N_4411,N_1695,N_1506);
nand U4412 (N_4412,N_1850,N_2043);
nor U4413 (N_4413,N_2346,N_2740);
nor U4414 (N_4414,N_2316,N_2593);
nor U4415 (N_4415,N_1690,N_2283);
and U4416 (N_4416,N_1916,N_2117);
or U4417 (N_4417,N_1944,N_2354);
nand U4418 (N_4418,N_1588,N_1740);
and U4419 (N_4419,N_2466,N_1815);
xor U4420 (N_4420,N_2810,N_2361);
xor U4421 (N_4421,N_1802,N_2027);
nand U4422 (N_4422,N_1635,N_2015);
and U4423 (N_4423,N_2758,N_1510);
or U4424 (N_4424,N_2597,N_2831);
or U4425 (N_4425,N_2815,N_2184);
nor U4426 (N_4426,N_2303,N_2701);
nand U4427 (N_4427,N_2715,N_2679);
nand U4428 (N_4428,N_1995,N_1796);
nand U4429 (N_4429,N_2180,N_2272);
nand U4430 (N_4430,N_1704,N_1839);
xor U4431 (N_4431,N_2215,N_1621);
xnor U4432 (N_4432,N_2829,N_2885);
nor U4433 (N_4433,N_1958,N_2917);
and U4434 (N_4434,N_2888,N_2492);
and U4435 (N_4435,N_2879,N_1980);
and U4436 (N_4436,N_1737,N_2342);
or U4437 (N_4437,N_1878,N_2923);
and U4438 (N_4438,N_2173,N_2358);
and U4439 (N_4439,N_2177,N_2208);
or U4440 (N_4440,N_2031,N_2971);
nand U4441 (N_4441,N_1810,N_2326);
xor U4442 (N_4442,N_1914,N_2472);
xor U4443 (N_4443,N_1903,N_2819);
and U4444 (N_4444,N_1555,N_1505);
xor U4445 (N_4445,N_2595,N_1502);
and U4446 (N_4446,N_2757,N_1923);
and U4447 (N_4447,N_1678,N_2911);
nand U4448 (N_4448,N_2038,N_2394);
nand U4449 (N_4449,N_2647,N_1645);
nor U4450 (N_4450,N_1630,N_2141);
or U4451 (N_4451,N_2737,N_2298);
xnor U4452 (N_4452,N_1847,N_2697);
nor U4453 (N_4453,N_1507,N_2570);
nand U4454 (N_4454,N_1917,N_2551);
nor U4455 (N_4455,N_2434,N_1797);
nor U4456 (N_4456,N_2898,N_2224);
nor U4457 (N_4457,N_2502,N_2293);
or U4458 (N_4458,N_2013,N_2119);
or U4459 (N_4459,N_1910,N_1783);
nor U4460 (N_4460,N_2521,N_2327);
nor U4461 (N_4461,N_2187,N_1618);
or U4462 (N_4462,N_1717,N_2352);
and U4463 (N_4463,N_1778,N_2235);
and U4464 (N_4464,N_1955,N_2118);
or U4465 (N_4465,N_1909,N_2923);
or U4466 (N_4466,N_2032,N_2355);
nand U4467 (N_4467,N_2629,N_1909);
and U4468 (N_4468,N_1772,N_2153);
nand U4469 (N_4469,N_1980,N_2026);
xnor U4470 (N_4470,N_2810,N_2353);
xor U4471 (N_4471,N_2357,N_2462);
or U4472 (N_4472,N_2544,N_2013);
nor U4473 (N_4473,N_2149,N_2573);
xor U4474 (N_4474,N_2423,N_2951);
nand U4475 (N_4475,N_1851,N_2365);
and U4476 (N_4476,N_1692,N_2055);
nor U4477 (N_4477,N_2934,N_2861);
nor U4478 (N_4478,N_2963,N_2254);
nand U4479 (N_4479,N_1858,N_1564);
nor U4480 (N_4480,N_2877,N_2743);
or U4481 (N_4481,N_2898,N_1620);
and U4482 (N_4482,N_1689,N_2059);
and U4483 (N_4483,N_2555,N_2677);
xor U4484 (N_4484,N_2712,N_2541);
nand U4485 (N_4485,N_2939,N_1735);
and U4486 (N_4486,N_1666,N_2489);
or U4487 (N_4487,N_2721,N_1911);
nor U4488 (N_4488,N_2046,N_1696);
xor U4489 (N_4489,N_1850,N_2269);
and U4490 (N_4490,N_2394,N_1709);
xor U4491 (N_4491,N_2918,N_2440);
nor U4492 (N_4492,N_2927,N_2632);
nor U4493 (N_4493,N_1752,N_2319);
or U4494 (N_4494,N_1749,N_2326);
nand U4495 (N_4495,N_2893,N_1908);
nand U4496 (N_4496,N_1911,N_2181);
xor U4497 (N_4497,N_1881,N_2901);
and U4498 (N_4498,N_2847,N_2800);
or U4499 (N_4499,N_2011,N_2740);
xnor U4500 (N_4500,N_3182,N_3586);
and U4501 (N_4501,N_4126,N_3839);
or U4502 (N_4502,N_4197,N_3192);
xnor U4503 (N_4503,N_3255,N_3505);
xor U4504 (N_4504,N_4073,N_4405);
or U4505 (N_4505,N_3357,N_3821);
and U4506 (N_4506,N_3576,N_3570);
nor U4507 (N_4507,N_4082,N_4050);
xor U4508 (N_4508,N_4267,N_4212);
nand U4509 (N_4509,N_3427,N_3828);
nor U4510 (N_4510,N_3591,N_3201);
or U4511 (N_4511,N_4366,N_4016);
xnor U4512 (N_4512,N_3419,N_3414);
or U4513 (N_4513,N_3812,N_3254);
and U4514 (N_4514,N_3196,N_3230);
nand U4515 (N_4515,N_3481,N_4314);
nor U4516 (N_4516,N_4176,N_4344);
nor U4517 (N_4517,N_3952,N_3112);
nand U4518 (N_4518,N_4364,N_3897);
nand U4519 (N_4519,N_3014,N_3880);
and U4520 (N_4520,N_3019,N_4084);
and U4521 (N_4521,N_3767,N_4068);
or U4522 (N_4522,N_3550,N_3150);
nand U4523 (N_4523,N_3604,N_3284);
and U4524 (N_4524,N_3883,N_3363);
xnor U4525 (N_4525,N_3486,N_3455);
xnor U4526 (N_4526,N_4418,N_3408);
nor U4527 (N_4527,N_3000,N_3130);
nand U4528 (N_4528,N_4341,N_3643);
or U4529 (N_4529,N_3453,N_3690);
and U4530 (N_4530,N_4386,N_3248);
xnor U4531 (N_4531,N_4428,N_4420);
nor U4532 (N_4532,N_3823,N_4227);
xnor U4533 (N_4533,N_4419,N_4247);
nor U4534 (N_4534,N_3713,N_3556);
or U4535 (N_4535,N_3833,N_3282);
nor U4536 (N_4536,N_4063,N_4069);
and U4537 (N_4537,N_4178,N_3057);
and U4538 (N_4538,N_4289,N_4061);
and U4539 (N_4539,N_3647,N_3631);
nand U4540 (N_4540,N_4125,N_3772);
and U4541 (N_4541,N_4146,N_4306);
or U4542 (N_4542,N_3675,N_3422);
nand U4543 (N_4543,N_4020,N_3537);
and U4544 (N_4544,N_4170,N_3781);
or U4545 (N_4545,N_4464,N_4269);
nand U4546 (N_4546,N_4083,N_3306);
xor U4547 (N_4547,N_4433,N_3773);
and U4548 (N_4548,N_3857,N_3371);
or U4549 (N_4549,N_3696,N_3871);
xnor U4550 (N_4550,N_3080,N_3754);
nor U4551 (N_4551,N_3267,N_3409);
and U4552 (N_4552,N_4272,N_3385);
and U4553 (N_4553,N_3558,N_4488);
nor U4554 (N_4554,N_3769,N_4116);
nor U4555 (N_4555,N_3168,N_3918);
xor U4556 (N_4556,N_3935,N_4240);
or U4557 (N_4557,N_3499,N_3161);
nor U4558 (N_4558,N_3341,N_3129);
nor U4559 (N_4559,N_3652,N_4299);
and U4560 (N_4560,N_3036,N_3110);
xnor U4561 (N_4561,N_3940,N_3572);
xnor U4562 (N_4562,N_4079,N_4128);
nand U4563 (N_4563,N_3712,N_3032);
or U4564 (N_4564,N_4097,N_4393);
nor U4565 (N_4565,N_3734,N_3686);
and U4566 (N_4566,N_3579,N_3017);
and U4567 (N_4567,N_3983,N_3293);
nor U4568 (N_4568,N_4437,N_4111);
xor U4569 (N_4569,N_3756,N_3273);
and U4570 (N_4570,N_3523,N_3753);
xor U4571 (N_4571,N_4431,N_3829);
nor U4572 (N_4572,N_4179,N_3216);
nand U4573 (N_4573,N_3418,N_4296);
nor U4574 (N_4574,N_3082,N_3491);
or U4575 (N_4575,N_4301,N_3529);
nand U4576 (N_4576,N_3008,N_3394);
or U4577 (N_4577,N_4481,N_4319);
or U4578 (N_4578,N_3976,N_4077);
or U4579 (N_4579,N_4101,N_3866);
and U4580 (N_4580,N_4136,N_3600);
nor U4581 (N_4581,N_3506,N_4000);
xor U4582 (N_4582,N_4311,N_3382);
and U4583 (N_4583,N_4307,N_4354);
and U4584 (N_4584,N_3636,N_4155);
and U4585 (N_4585,N_3396,N_4066);
xnor U4586 (N_4586,N_4279,N_3795);
xor U4587 (N_4587,N_3645,N_4138);
or U4588 (N_4588,N_3185,N_4490);
nor U4589 (N_4589,N_3628,N_4198);
nor U4590 (N_4590,N_4193,N_4142);
nor U4591 (N_4591,N_3512,N_4292);
and U4592 (N_4592,N_4495,N_4394);
nor U4593 (N_4593,N_3778,N_3266);
xor U4594 (N_4594,N_3722,N_4435);
nand U4595 (N_4595,N_4389,N_3961);
and U4596 (N_4596,N_4172,N_4003);
and U4597 (N_4597,N_3583,N_4338);
nor U4598 (N_4598,N_4283,N_3519);
and U4599 (N_4599,N_4022,N_4373);
and U4600 (N_4600,N_3531,N_3748);
nor U4601 (N_4601,N_3659,N_3485);
nor U4602 (N_4602,N_3641,N_4447);
xnor U4603 (N_4603,N_4166,N_3687);
and U4604 (N_4604,N_3058,N_3165);
nand U4605 (N_4605,N_3830,N_4105);
nand U4606 (N_4606,N_3252,N_3937);
and U4607 (N_4607,N_3740,N_4315);
and U4608 (N_4608,N_3808,N_3428);
nand U4609 (N_4609,N_4165,N_4270);
nand U4610 (N_4610,N_3494,N_3752);
or U4611 (N_4611,N_4233,N_3179);
or U4612 (N_4612,N_3791,N_4032);
nor U4613 (N_4613,N_3120,N_4297);
nand U4614 (N_4614,N_3336,N_3692);
xnor U4615 (N_4615,N_3048,N_3475);
xor U4616 (N_4616,N_3009,N_3038);
nor U4617 (N_4617,N_3896,N_4329);
and U4618 (N_4618,N_3184,N_3815);
or U4619 (N_4619,N_3317,N_3814);
and U4620 (N_4620,N_3356,N_3303);
and U4621 (N_4621,N_3542,N_4019);
xor U4622 (N_4622,N_4305,N_3551);
xor U4623 (N_4623,N_3202,N_3318);
nor U4624 (N_4624,N_3820,N_3606);
or U4625 (N_4625,N_3931,N_3194);
or U4626 (N_4626,N_4472,N_3043);
or U4627 (N_4627,N_3545,N_4245);
nor U4628 (N_4628,N_4205,N_3077);
xor U4629 (N_4629,N_3089,N_4446);
nand U4630 (N_4630,N_3471,N_3510);
or U4631 (N_4631,N_3214,N_4324);
and U4632 (N_4632,N_3169,N_4187);
or U4633 (N_4633,N_3580,N_4340);
or U4634 (N_4634,N_3941,N_3978);
xnor U4635 (N_4635,N_4429,N_4293);
nand U4636 (N_4636,N_3390,N_3372);
nor U4637 (N_4637,N_3642,N_4453);
nand U4638 (N_4638,N_3307,N_4094);
and U4639 (N_4639,N_3650,N_3905);
and U4640 (N_4640,N_3800,N_3953);
or U4641 (N_4641,N_3707,N_3904);
or U4642 (N_4642,N_4281,N_4460);
or U4643 (N_4643,N_4201,N_3208);
xnor U4644 (N_4644,N_3850,N_4027);
or U4645 (N_4645,N_3780,N_3508);
xor U4646 (N_4646,N_3251,N_3527);
xor U4647 (N_4647,N_3682,N_3386);
nand U4648 (N_4648,N_4448,N_3714);
nor U4649 (N_4649,N_4371,N_3725);
xnor U4650 (N_4650,N_4377,N_4457);
nand U4651 (N_4651,N_4333,N_3775);
or U4652 (N_4652,N_3015,N_3536);
xnor U4653 (N_4653,N_4362,N_3233);
or U4654 (N_4654,N_3012,N_3835);
nor U4655 (N_4655,N_3105,N_3916);
and U4656 (N_4656,N_3278,N_4452);
and U4657 (N_4657,N_3805,N_3242);
nand U4658 (N_4658,N_3374,N_3164);
nand U4659 (N_4659,N_3802,N_3296);
xnor U4660 (N_4660,N_3400,N_3421);
xnor U4661 (N_4661,N_3993,N_3539);
or U4662 (N_4662,N_4347,N_3315);
or U4663 (N_4663,N_3730,N_3083);
or U4664 (N_4664,N_4028,N_3991);
nand U4665 (N_4665,N_4328,N_3220);
xor U4666 (N_4666,N_4018,N_3430);
and U4667 (N_4667,N_3774,N_3660);
nand U4668 (N_4668,N_4114,N_4023);
and U4669 (N_4669,N_3885,N_3362);
and U4670 (N_4670,N_3697,N_3259);
xor U4671 (N_4671,N_3724,N_3788);
or U4672 (N_4672,N_4339,N_3140);
xnor U4673 (N_4673,N_3138,N_3644);
nor U4674 (N_4674,N_3555,N_3424);
nor U4675 (N_4675,N_3465,N_4007);
nand U4676 (N_4676,N_4242,N_4103);
nor U4677 (N_4677,N_4130,N_3117);
nand U4678 (N_4678,N_3030,N_4234);
xor U4679 (N_4679,N_3187,N_3440);
nand U4680 (N_4680,N_3244,N_4057);
nor U4681 (N_4681,N_3258,N_4288);
and U4682 (N_4682,N_3005,N_3035);
nor U4683 (N_4683,N_3776,N_3342);
and U4684 (N_4684,N_4291,N_3658);
nand U4685 (N_4685,N_3560,N_4383);
nor U4686 (N_4686,N_3403,N_3627);
or U4687 (N_4687,N_3156,N_3909);
nor U4688 (N_4688,N_4218,N_4332);
nand U4689 (N_4689,N_4026,N_3344);
nand U4690 (N_4690,N_4033,N_3526);
nor U4691 (N_4691,N_4115,N_3862);
and U4692 (N_4692,N_3297,N_4408);
nor U4693 (N_4693,N_3898,N_3167);
xnor U4694 (N_4694,N_4056,N_3437);
or U4695 (N_4695,N_4425,N_3314);
and U4696 (N_4696,N_3966,N_4204);
and U4697 (N_4697,N_3972,N_3786);
or U4698 (N_4698,N_3176,N_3792);
or U4699 (N_4699,N_4403,N_4396);
and U4700 (N_4700,N_4238,N_4298);
nor U4701 (N_4701,N_4127,N_3115);
xor U4702 (N_4702,N_3877,N_3137);
nand U4703 (N_4703,N_3420,N_4439);
nand U4704 (N_4704,N_3118,N_4098);
nor U4705 (N_4705,N_4192,N_4219);
xnor U4706 (N_4706,N_3231,N_3521);
nor U4707 (N_4707,N_3163,N_3973);
nor U4708 (N_4708,N_3949,N_4322);
or U4709 (N_4709,N_3013,N_3124);
and U4710 (N_4710,N_3106,N_4134);
nand U4711 (N_4711,N_4042,N_4398);
and U4712 (N_4712,N_3869,N_4356);
or U4713 (N_4713,N_3655,N_4417);
or U4714 (N_4714,N_4411,N_3899);
and U4715 (N_4715,N_4380,N_3876);
xnor U4716 (N_4716,N_3148,N_3022);
or U4717 (N_4717,N_3698,N_4232);
xor U4718 (N_4718,N_3771,N_4183);
and U4719 (N_4719,N_3737,N_3376);
or U4720 (N_4720,N_3107,N_4294);
xor U4721 (N_4721,N_3407,N_4335);
and U4722 (N_4722,N_4214,N_3287);
nand U4723 (N_4723,N_4081,N_3971);
xnor U4724 (N_4724,N_3728,N_3186);
nand U4725 (N_4725,N_3480,N_4017);
or U4726 (N_4726,N_3253,N_3703);
and U4727 (N_4727,N_3274,N_3392);
nor U4728 (N_4728,N_3665,N_4467);
and U4729 (N_4729,N_3018,N_3159);
or U4730 (N_4730,N_3195,N_3676);
nor U4731 (N_4731,N_3964,N_3663);
nor U4732 (N_4732,N_3654,N_4392);
xnor U4733 (N_4733,N_3436,N_4002);
and U4734 (N_4734,N_3601,N_3152);
and U4735 (N_4735,N_3908,N_3640);
nor U4736 (N_4736,N_3339,N_3878);
and U4737 (N_4737,N_3711,N_4226);
and U4738 (N_4738,N_4323,N_4388);
xnor U4739 (N_4739,N_3181,N_3178);
and U4740 (N_4740,N_3467,N_3744);
nand U4741 (N_4741,N_4475,N_3996);
and U4742 (N_4742,N_3548,N_4235);
xor U4743 (N_4743,N_4090,N_4038);
nor U4744 (N_4744,N_3229,N_4182);
xor U4745 (N_4745,N_3567,N_3649);
and U4746 (N_4746,N_4053,N_3813);
nand U4747 (N_4747,N_4132,N_3189);
nor U4748 (N_4748,N_3096,N_3388);
nor U4749 (N_4749,N_3350,N_4361);
or U4750 (N_4750,N_3810,N_4015);
or U4751 (N_4751,N_3262,N_3701);
nand U4752 (N_4752,N_3476,N_3693);
xor U4753 (N_4753,N_3981,N_3349);
xor U4754 (N_4754,N_4367,N_3629);
or U4755 (N_4755,N_4195,N_3352);
nor U4756 (N_4756,N_3291,N_4256);
or U4757 (N_4757,N_3323,N_3716);
nor U4758 (N_4758,N_4345,N_3568);
or U4759 (N_4759,N_4159,N_3530);
and U4760 (N_4760,N_4313,N_3651);
or U4761 (N_4761,N_3429,N_3538);
xnor U4762 (N_4762,N_3582,N_3474);
xnor U4763 (N_4763,N_4241,N_3546);
xnor U4764 (N_4764,N_4284,N_3102);
nand U4765 (N_4765,N_3395,N_4080);
xor U4766 (N_4766,N_3068,N_3482);
xor U4767 (N_4767,N_3171,N_3369);
nor U4768 (N_4768,N_4499,N_3779);
or U4769 (N_4769,N_3127,N_3797);
xnor U4770 (N_4770,N_4440,N_3843);
and U4771 (N_4771,N_3033,N_3842);
nor U4772 (N_4772,N_4237,N_4060);
nor U4773 (N_4773,N_3379,N_3915);
nor U4774 (N_4774,N_3328,N_3515);
xor U4775 (N_4775,N_4492,N_4331);
or U4776 (N_4776,N_3360,N_3459);
nand U4777 (N_4777,N_3045,N_3708);
nand U4778 (N_4778,N_3348,N_3272);
nand U4779 (N_4779,N_4211,N_4058);
nor U4780 (N_4780,N_4102,N_3219);
or U4781 (N_4781,N_4310,N_3340);
and U4782 (N_4782,N_4484,N_3925);
nand U4783 (N_4783,N_3922,N_4352);
xnor U4784 (N_4784,N_3544,N_3321);
and U4785 (N_4785,N_4265,N_3479);
xor U4786 (N_4786,N_4251,N_4466);
nand U4787 (N_4787,N_3415,N_4434);
or U4788 (N_4788,N_3046,N_3276);
xor U4789 (N_4789,N_3330,N_4175);
or U4790 (N_4790,N_3581,N_3919);
or U4791 (N_4791,N_3602,N_4399);
nand U4792 (N_4792,N_4229,N_4140);
xnor U4793 (N_4793,N_3329,N_3007);
xor U4794 (N_4794,N_3126,N_4406);
and U4795 (N_4795,N_3086,N_3028);
or U4796 (N_4796,N_4282,N_4054);
or U4797 (N_4797,N_3836,N_3451);
and U4798 (N_4798,N_3589,N_3888);
nor U4799 (N_4799,N_3818,N_4275);
or U4800 (N_4800,N_4099,N_4423);
xnor U4801 (N_4801,N_3367,N_3784);
xnor U4802 (N_4802,N_3950,N_4171);
or U4803 (N_4803,N_3070,N_4008);
xor U4804 (N_4804,N_3621,N_4494);
nor U4805 (N_4805,N_3995,N_3504);
nor U4806 (N_4806,N_3166,N_4030);
and U4807 (N_4807,N_3975,N_3280);
nand U4808 (N_4808,N_3794,N_4308);
nand U4809 (N_4809,N_3074,N_4223);
nand U4810 (N_4810,N_3705,N_4150);
xnor U4811 (N_4811,N_3378,N_3782);
nand U4812 (N_4812,N_3986,N_3003);
nor U4813 (N_4813,N_3912,N_3084);
or U4814 (N_4814,N_3518,N_4257);
and U4815 (N_4815,N_4129,N_4470);
nand U4816 (N_4816,N_4185,N_3669);
xnor U4817 (N_4817,N_4104,N_3689);
and U4818 (N_4818,N_3943,N_3623);
and U4819 (N_4819,N_3135,N_4385);
and U4820 (N_4820,N_4342,N_4372);
nor U4821 (N_4821,N_3337,N_3345);
nor U4822 (N_4822,N_3099,N_3806);
nor U4823 (N_4823,N_3222,N_3399);
or U4824 (N_4824,N_3463,N_4100);
nand U4825 (N_4825,N_4153,N_3569);
nand U4826 (N_4826,N_3932,N_3445);
or U4827 (N_4827,N_3155,N_3006);
nor U4828 (N_4828,N_4285,N_4106);
xnor U4829 (N_4829,N_3679,N_3511);
and U4830 (N_4830,N_4424,N_4262);
nor U4831 (N_4831,N_4365,N_4215);
or U4832 (N_4832,N_3218,N_3997);
nand U4833 (N_4833,N_4149,N_3809);
nand U4834 (N_4834,N_3639,N_3980);
nand U4835 (N_4835,N_3144,N_3071);
or U4836 (N_4836,N_3522,N_4255);
and U4837 (N_4837,N_3861,N_3439);
nor U4838 (N_4838,N_3011,N_4051);
nor U4839 (N_4839,N_3726,N_3232);
nor U4840 (N_4840,N_3078,N_3358);
nor U4841 (N_4841,N_4259,N_3989);
nor U4842 (N_4842,N_3840,N_4407);
nand U4843 (N_4843,N_4133,N_3999);
nand U4844 (N_4844,N_3260,N_4184);
xnor U4845 (N_4845,N_3204,N_4312);
and U4846 (N_4846,N_3607,N_3928);
or U4847 (N_4847,N_3132,N_3936);
nor U4848 (N_4848,N_3867,N_3653);
nand U4849 (N_4849,N_3370,N_4163);
and U4850 (N_4850,N_3816,N_4065);
nor U4851 (N_4851,N_3079,N_3023);
and U4852 (N_4852,N_3533,N_3624);
or U4853 (N_4853,N_3359,N_3844);
or U4854 (N_4854,N_4387,N_3063);
and U4855 (N_4855,N_3532,N_4210);
nand U4856 (N_4856,N_3865,N_4239);
and U4857 (N_4857,N_3826,N_3552);
and U4858 (N_4858,N_3121,N_3547);
nand U4859 (N_4859,N_3327,N_3295);
and U4860 (N_4860,N_3270,N_4276);
nor U4861 (N_4861,N_3747,N_3947);
nand U4862 (N_4862,N_3487,N_3309);
xor U4863 (N_4863,N_3501,N_3709);
xor U4864 (N_4864,N_3462,N_4055);
and U4865 (N_4865,N_4248,N_3031);
xnor U4866 (N_4866,N_3587,N_3488);
nand U4867 (N_4867,N_3847,N_3852);
nand U4868 (N_4868,N_4360,N_4326);
nor U4869 (N_4869,N_4085,N_4161);
xnor U4870 (N_4870,N_3900,N_3901);
xnor U4871 (N_4871,N_3319,N_3930);
xor U4872 (N_4872,N_3346,N_3226);
or U4873 (N_4873,N_3069,N_3749);
nor U4874 (N_4874,N_3332,N_3870);
xnor U4875 (N_4875,N_4112,N_3768);
nand U4876 (N_4876,N_3425,N_3442);
xor U4877 (N_4877,N_4209,N_3605);
nor U4878 (N_4878,N_3597,N_3745);
xnor U4879 (N_4879,N_3434,N_3312);
xnor U4880 (N_4880,N_3147,N_3405);
and U4881 (N_4881,N_3097,N_3055);
xnor U4882 (N_4882,N_3819,N_3020);
xnor U4883 (N_4883,N_3757,N_4225);
nor U4884 (N_4884,N_4432,N_3913);
or U4885 (N_4885,N_3109,N_4334);
nor U4886 (N_4886,N_3059,N_3391);
and U4887 (N_4887,N_3128,N_4445);
and U4888 (N_4888,N_3695,N_4273);
and U4889 (N_4889,N_3305,N_4011);
and U4890 (N_4890,N_3796,N_4089);
or U4891 (N_4891,N_3064,N_4468);
or U4892 (N_4892,N_4369,N_3541);
xor U4893 (N_4893,N_3879,N_4391);
xnor U4894 (N_4894,N_4188,N_4124);
xnor U4895 (N_4895,N_4181,N_4249);
nor U4896 (N_4896,N_3777,N_3114);
xnor U4897 (N_4897,N_4477,N_3962);
nor U4898 (N_4898,N_4168,N_3100);
and U4899 (N_4899,N_4045,N_3793);
xnor U4900 (N_4900,N_3268,N_3575);
nand U4901 (N_4901,N_3603,N_3497);
or U4902 (N_4902,N_4064,N_4160);
nand U4903 (N_4903,N_3368,N_3264);
and U4904 (N_4904,N_3613,N_4337);
xor U4905 (N_4905,N_3402,N_3618);
and U4906 (N_4906,N_3619,N_3383);
nand U4907 (N_4907,N_4286,N_4031);
or U4908 (N_4908,N_3225,N_4461);
nor U4909 (N_4909,N_3503,N_3113);
and U4910 (N_4910,N_3743,N_4449);
or U4911 (N_4911,N_4156,N_3746);
and U4912 (N_4912,N_3566,N_3721);
nand U4913 (N_4913,N_3308,N_3448);
nor U4914 (N_4914,N_3066,N_4379);
or U4915 (N_4915,N_3733,N_3052);
xor U4916 (N_4916,N_3131,N_3310);
xnor U4917 (N_4917,N_3191,N_3210);
or U4918 (N_4918,N_4200,N_3955);
nor U4919 (N_4919,N_3617,N_4421);
or U4920 (N_4920,N_3719,N_4295);
nor U4921 (N_4921,N_3633,N_4122);
xor U4922 (N_4922,N_4052,N_3817);
nand U4923 (N_4923,N_4402,N_4462);
nor U4924 (N_4924,N_3119,N_3635);
nor U4925 (N_4925,N_3732,N_3584);
xnor U4926 (N_4926,N_3288,N_4154);
or U4927 (N_4927,N_3944,N_3670);
and U4928 (N_4928,N_3979,N_4436);
xnor U4929 (N_4929,N_3237,N_3688);
or U4930 (N_4930,N_3081,N_3304);
or U4931 (N_4931,N_3513,N_3271);
or U4932 (N_4932,N_4095,N_3520);
xnor U4933 (N_4933,N_3827,N_3894);
nand U4934 (N_4934,N_3458,N_3466);
and U4935 (N_4935,N_3302,N_4415);
nor U4936 (N_4936,N_3456,N_3141);
xor U4937 (N_4937,N_4118,N_4479);
xor U4938 (N_4938,N_3946,N_3404);
and U4939 (N_4939,N_3438,N_3984);
xnor U4940 (N_4940,N_3939,N_4152);
or U4941 (N_4941,N_4368,N_3927);
xnor U4942 (N_4942,N_3384,N_3433);
and U4943 (N_4943,N_3460,N_3449);
xnor U4944 (N_4944,N_4316,N_3143);
xor U4945 (N_4945,N_3873,N_3236);
and U4946 (N_4946,N_3149,N_4348);
nand U4947 (N_4947,N_3042,N_3238);
nor U4948 (N_4948,N_4086,N_3301);
nand U4949 (N_4949,N_4498,N_3763);
or U4950 (N_4950,N_3553,N_4280);
or U4951 (N_4951,N_3316,N_3626);
nand U4952 (N_4952,N_4001,N_3470);
or U4953 (N_4953,N_4137,N_3087);
or U4954 (N_4954,N_3412,N_4474);
and U4955 (N_4955,N_4072,N_4148);
and U4956 (N_4956,N_3257,N_3333);
or U4957 (N_4957,N_3249,N_4497);
and U4958 (N_4958,N_3738,N_3090);
xnor U4959 (N_4959,N_3095,N_4190);
or U4960 (N_4960,N_3637,N_3889);
nor U4961 (N_4961,N_3672,N_3596);
nand U4962 (N_4962,N_4287,N_3625);
nand U4963 (N_4963,N_4422,N_4317);
xnor U4964 (N_4964,N_4351,N_4370);
and U4965 (N_4965,N_3413,N_4049);
xor U4966 (N_4966,N_4143,N_3807);
and U4967 (N_4967,N_3571,N_4131);
nor U4968 (N_4968,N_4455,N_3516);
and U4969 (N_4969,N_3588,N_4300);
nor U4970 (N_4970,N_4220,N_4350);
nand U4971 (N_4971,N_4107,N_4169);
or U4972 (N_4972,N_3798,N_3620);
or U4973 (N_4973,N_4109,N_3938);
nor U4974 (N_4974,N_3982,N_3366);
xor U4975 (N_4975,N_3911,N_3211);
nor U4976 (N_4976,N_4006,N_4443);
nand U4977 (N_4977,N_4009,N_4302);
or U4978 (N_4978,N_3426,N_4473);
nor U4979 (N_4979,N_4246,N_3585);
nand U4980 (N_4980,N_3561,N_3162);
xnor U4981 (N_4981,N_4147,N_4349);
or U4982 (N_4982,N_4194,N_4024);
xnor U4983 (N_4983,N_3294,N_4378);
and U4984 (N_4984,N_3235,N_3334);
nand U4985 (N_4985,N_3801,N_3103);
nor U4986 (N_4986,N_3261,N_4224);
nor U4987 (N_4987,N_3373,N_4034);
nor U4988 (N_4988,N_3313,N_4208);
or U4989 (N_4989,N_4117,N_3454);
nor U4990 (N_4990,N_4384,N_3859);
xor U4991 (N_4991,N_3563,N_3024);
nor U4992 (N_4992,N_3151,N_3578);
nand U4993 (N_4993,N_3755,N_3331);
and U4994 (N_4994,N_3338,N_3172);
xor U4995 (N_4995,N_3684,N_3656);
nand U4996 (N_4996,N_3864,N_3298);
xor U4997 (N_4997,N_3706,N_3785);
and U4998 (N_4998,N_3612,N_3401);
xnor U4999 (N_4999,N_3849,N_3397);
nor U5000 (N_5000,N_3729,N_3514);
or U5001 (N_5001,N_3224,N_3142);
and U5002 (N_5002,N_3246,N_3489);
and U5003 (N_5003,N_3205,N_3892);
xor U5004 (N_5004,N_3175,N_3203);
or U5005 (N_5005,N_4320,N_4043);
nand U5006 (N_5006,N_3256,N_3634);
nor U5007 (N_5007,N_3929,N_3848);
or U5008 (N_5008,N_3450,N_3493);
nand U5009 (N_5009,N_3914,N_3906);
xnor U5010 (N_5010,N_3838,N_3067);
and U5011 (N_5011,N_3177,N_3920);
xor U5012 (N_5012,N_3760,N_3787);
or U5013 (N_5013,N_3039,N_4353);
or U5014 (N_5014,N_4206,N_3863);
xor U5015 (N_5015,N_3431,N_4139);
and U5016 (N_5016,N_4463,N_3389);
xnor U5017 (N_5017,N_3281,N_3685);
nand U5018 (N_5018,N_3361,N_3406);
xor U5019 (N_5019,N_3674,N_3285);
or U5020 (N_5020,N_4014,N_3882);
nand U5021 (N_5021,N_4013,N_3783);
or U5022 (N_5022,N_3299,N_4254);
xnor U5023 (N_5023,N_3959,N_4021);
or U5024 (N_5024,N_3803,N_4277);
or U5025 (N_5025,N_3180,N_4216);
and U5026 (N_5026,N_3207,N_4359);
nor U5027 (N_5027,N_3154,N_4046);
nand U5028 (N_5028,N_4071,N_4450);
nor U5029 (N_5029,N_3292,N_3498);
nor U5030 (N_5030,N_3985,N_3846);
xnor U5031 (N_5031,N_4469,N_3234);
nor U5032 (N_5032,N_3410,N_3353);
or U5033 (N_5033,N_3874,N_3855);
xnor U5034 (N_5034,N_3790,N_3764);
xnor U5035 (N_5035,N_4096,N_4157);
nor U5036 (N_5036,N_4363,N_4180);
and U5037 (N_5037,N_3001,N_4113);
nor U5038 (N_5038,N_3034,N_3193);
xnor U5039 (N_5039,N_4035,N_3146);
xor U5040 (N_5040,N_3960,N_3824);
xnor U5041 (N_5041,N_4203,N_4491);
nand U5042 (N_5042,N_4230,N_3300);
nand U5043 (N_5043,N_3076,N_3461);
or U5044 (N_5044,N_4309,N_3263);
xor U5045 (N_5045,N_3432,N_3666);
and U5046 (N_5046,N_3592,N_3765);
and U5047 (N_5047,N_4228,N_3170);
nand U5048 (N_5048,N_3887,N_3444);
xor U5049 (N_5049,N_3988,N_3040);
nand U5050 (N_5050,N_3073,N_3072);
nand U5051 (N_5051,N_3477,N_3221);
nor U5052 (N_5052,N_4213,N_4401);
xnor U5053 (N_5053,N_3832,N_3265);
xor U5054 (N_5054,N_3942,N_3464);
or U5055 (N_5055,N_4123,N_3535);
and U5056 (N_5056,N_3381,N_3411);
or U5057 (N_5057,N_3029,N_4303);
nor U5058 (N_5058,N_3926,N_4036);
nor U5059 (N_5059,N_3239,N_4357);
nand U5060 (N_5060,N_4266,N_4162);
and U5061 (N_5061,N_3183,N_4478);
or U5062 (N_5062,N_4135,N_3277);
nand U5063 (N_5063,N_3923,N_3473);
nor U5064 (N_5064,N_3851,N_3500);
and U5065 (N_5065,N_3965,N_3021);
or U5066 (N_5066,N_3608,N_4075);
or U5067 (N_5067,N_3967,N_3026);
or U5068 (N_5068,N_4260,N_3990);
or U5069 (N_5069,N_3718,N_3243);
xor U5070 (N_5070,N_3104,N_3134);
xor U5071 (N_5071,N_3101,N_3227);
xnor U5072 (N_5072,N_3811,N_4252);
nand U5073 (N_5073,N_4236,N_3657);
and U5074 (N_5074,N_4087,N_3215);
xnor U5075 (N_5075,N_4158,N_4395);
xnor U5076 (N_5076,N_3699,N_3858);
xnor U5077 (N_5077,N_3691,N_3921);
xnor U5078 (N_5078,N_3452,N_3700);
and U5079 (N_5079,N_3630,N_3398);
or U5080 (N_5080,N_4390,N_4410);
nand U5081 (N_5081,N_3375,N_3133);
and U5082 (N_5082,N_4037,N_3974);
xnor U5083 (N_5083,N_3895,N_4325);
or U5084 (N_5084,N_3153,N_4253);
and U5085 (N_5085,N_4186,N_4261);
nor U5086 (N_5086,N_3056,N_4145);
xnor U5087 (N_5087,N_3478,N_3320);
xnor U5088 (N_5088,N_4151,N_4059);
or U5089 (N_5089,N_4327,N_3213);
nand U5090 (N_5090,N_4321,N_3594);
and U5091 (N_5091,N_3393,N_3751);
nor U5092 (N_5092,N_4438,N_3116);
xnor U5093 (N_5093,N_3188,N_3173);
and U5094 (N_5094,N_4271,N_3540);
or U5095 (N_5095,N_3881,N_3441);
and U5096 (N_5096,N_3492,N_4480);
or U5097 (N_5097,N_3994,N_3355);
and U5098 (N_5098,N_3903,N_3275);
or U5099 (N_5099,N_3041,N_3250);
or U5100 (N_5100,N_3595,N_4416);
or U5101 (N_5101,N_3593,N_3661);
xnor U5102 (N_5102,N_3562,N_3956);
and U5103 (N_5103,N_3365,N_3190);
xnor U5104 (N_5104,N_3094,N_4164);
or U5105 (N_5105,N_3992,N_3948);
xnor U5106 (N_5106,N_3435,N_3525);
and U5107 (N_5107,N_3158,N_4442);
or U5108 (N_5108,N_3934,N_4485);
or U5109 (N_5109,N_3742,N_3615);
or U5110 (N_5110,N_4191,N_3758);
xnor U5111 (N_5111,N_3343,N_3247);
xor U5112 (N_5112,N_4404,N_4048);
nand U5113 (N_5113,N_3469,N_4088);
nor U5114 (N_5114,N_3060,N_4041);
nor U5115 (N_5115,N_3609,N_4119);
and U5116 (N_5116,N_3891,N_3610);
xor U5117 (N_5117,N_3240,N_3710);
or U5118 (N_5118,N_3958,N_3098);
xnor U5119 (N_5119,N_3598,N_4091);
and U5120 (N_5120,N_3085,N_3969);
nand U5121 (N_5121,N_4482,N_3614);
or U5122 (N_5122,N_3681,N_4346);
nor U5123 (N_5123,N_3717,N_4231);
nand U5124 (N_5124,N_3590,N_4496);
or U5125 (N_5125,N_3577,N_3831);
and U5126 (N_5126,N_3311,N_3423);
nor U5127 (N_5127,N_4381,N_4264);
nor U5128 (N_5128,N_3047,N_4070);
nor U5129 (N_5129,N_4465,N_3622);
nor U5130 (N_5130,N_3907,N_3053);
nor U5131 (N_5131,N_4141,N_3054);
or U5132 (N_5132,N_3322,N_4413);
or U5133 (N_5133,N_3416,N_3198);
and U5134 (N_5134,N_4476,N_3557);
nor U5135 (N_5135,N_3902,N_3223);
nor U5136 (N_5136,N_3289,N_3049);
nor U5137 (N_5137,N_3123,N_3025);
nor U5138 (N_5138,N_3139,N_3092);
nand U5139 (N_5139,N_3977,N_3761);
or U5140 (N_5140,N_4062,N_4039);
nand U5141 (N_5141,N_3088,N_3667);
nor U5142 (N_5142,N_3125,N_4044);
nor U5143 (N_5143,N_4202,N_3573);
nand U5144 (N_5144,N_3484,N_3122);
xnor U5145 (N_5145,N_3616,N_3822);
nand U5146 (N_5146,N_4221,N_3443);
or U5147 (N_5147,N_3269,N_3668);
xor U5148 (N_5148,N_4196,N_3770);
nand U5149 (N_5149,N_4409,N_3002);
nor U5150 (N_5150,N_4397,N_3945);
or U5151 (N_5151,N_4426,N_3495);
xnor U5152 (N_5152,N_3678,N_3010);
and U5153 (N_5153,N_4040,N_4374);
xnor U5154 (N_5154,N_3741,N_4274);
nor U5155 (N_5155,N_3091,N_4244);
nand U5156 (N_5156,N_3559,N_3283);
and U5157 (N_5157,N_3174,N_3004);
or U5158 (N_5158,N_3789,N_4382);
nor U5159 (N_5159,N_3739,N_3854);
and U5160 (N_5160,N_3825,N_3868);
xnor U5161 (N_5161,N_4120,N_4414);
xor U5162 (N_5162,N_3554,N_3662);
nor U5163 (N_5163,N_3680,N_3093);
xor U5164 (N_5164,N_3549,N_4268);
or U5165 (N_5165,N_4029,N_4189);
nand U5166 (N_5166,N_4441,N_4444);
xor U5167 (N_5167,N_3910,N_3447);
and U5168 (N_5168,N_4217,N_3720);
nor U5169 (N_5169,N_4173,N_4471);
nand U5170 (N_5170,N_3446,N_3351);
nor U5171 (N_5171,N_3957,N_4330);
or U5172 (N_5172,N_3543,N_4355);
xnor U5173 (N_5173,N_4093,N_3286);
and U5174 (N_5174,N_3347,N_4010);
and U5175 (N_5175,N_4486,N_3884);
and U5176 (N_5176,N_3970,N_3694);
nor U5177 (N_5177,N_4483,N_3217);
nand U5178 (N_5178,N_4487,N_3924);
xor U5179 (N_5179,N_3646,N_3565);
nor U5180 (N_5180,N_3241,N_3417);
nor U5181 (N_5181,N_3528,N_3704);
or U5182 (N_5182,N_3325,N_3037);
nand U5183 (N_5183,N_3853,N_3468);
or U5184 (N_5184,N_4174,N_3987);
nor U5185 (N_5185,N_3648,N_4343);
or U5186 (N_5186,N_3380,N_3611);
nand U5187 (N_5187,N_3564,N_3136);
xnor U5188 (N_5188,N_3364,N_3496);
nor U5189 (N_5189,N_3723,N_3715);
xor U5190 (N_5190,N_3893,N_3875);
nor U5191 (N_5191,N_3759,N_3050);
and U5192 (N_5192,N_3841,N_3856);
nor U5193 (N_5193,N_4451,N_4110);
and U5194 (N_5194,N_4290,N_3677);
and U5195 (N_5195,N_4222,N_3804);
or U5196 (N_5196,N_3075,N_3963);
xor U5197 (N_5197,N_4376,N_3354);
nor U5198 (N_5198,N_3890,N_3279);
nand U5199 (N_5199,N_4400,N_3998);
xor U5200 (N_5200,N_3324,N_4358);
nand U5201 (N_5201,N_3731,N_3387);
or U5202 (N_5202,N_3727,N_4263);
xnor U5203 (N_5203,N_3483,N_4005);
and U5204 (N_5204,N_3200,N_3917);
xnor U5205 (N_5205,N_3206,N_3762);
or U5206 (N_5206,N_3157,N_4459);
nor U5207 (N_5207,N_3245,N_3599);
and U5208 (N_5208,N_3016,N_3472);
nand U5209 (N_5209,N_4304,N_3671);
or U5210 (N_5210,N_4318,N_4207);
xor U5211 (N_5211,N_4427,N_3502);
nor U5212 (N_5212,N_4278,N_3160);
nor U5213 (N_5213,N_3933,N_4092);
nor U5214 (N_5214,N_4025,N_3750);
and U5215 (N_5215,N_4456,N_3673);
nor U5216 (N_5216,N_4121,N_3664);
xor U5217 (N_5217,N_4144,N_3517);
or U5218 (N_5218,N_3377,N_3702);
nor U5219 (N_5219,N_3534,N_3199);
or U5220 (N_5220,N_3632,N_3051);
nand U5221 (N_5221,N_4004,N_4258);
nor U5222 (N_5222,N_3108,N_4177);
xnor U5223 (N_5223,N_3111,N_3574);
nand U5224 (N_5224,N_3145,N_3683);
and U5225 (N_5225,N_3290,N_3065);
nand U5226 (N_5226,N_4199,N_3209);
and U5227 (N_5227,N_4012,N_3228);
nor U5228 (N_5228,N_4375,N_3062);
or U5229 (N_5229,N_4047,N_3212);
or U5230 (N_5230,N_3197,N_3735);
nor U5231 (N_5231,N_4336,N_3027);
nand U5232 (N_5232,N_3951,N_3509);
and U5233 (N_5233,N_4454,N_4458);
nand U5234 (N_5234,N_4074,N_3335);
nor U5235 (N_5235,N_3834,N_4078);
or U5236 (N_5236,N_3061,N_3845);
and U5237 (N_5237,N_4243,N_3860);
and U5238 (N_5238,N_3524,N_4489);
and U5239 (N_5239,N_3507,N_4250);
xor U5240 (N_5240,N_3638,N_4412);
nor U5241 (N_5241,N_3872,N_3837);
or U5242 (N_5242,N_4167,N_3044);
xor U5243 (N_5243,N_3954,N_3736);
or U5244 (N_5244,N_4430,N_3766);
or U5245 (N_5245,N_4493,N_3326);
xor U5246 (N_5246,N_4067,N_3968);
nand U5247 (N_5247,N_4108,N_3490);
and U5248 (N_5248,N_3886,N_3799);
and U5249 (N_5249,N_4076,N_3457);
nor U5250 (N_5250,N_3990,N_3364);
nand U5251 (N_5251,N_3125,N_4269);
or U5252 (N_5252,N_3597,N_3054);
or U5253 (N_5253,N_3799,N_3395);
and U5254 (N_5254,N_4407,N_3288);
nand U5255 (N_5255,N_3103,N_3517);
nand U5256 (N_5256,N_3837,N_3282);
nor U5257 (N_5257,N_3467,N_3842);
xnor U5258 (N_5258,N_4107,N_3021);
xor U5259 (N_5259,N_3545,N_3846);
nand U5260 (N_5260,N_3474,N_3716);
or U5261 (N_5261,N_3432,N_3046);
nand U5262 (N_5262,N_3007,N_3142);
nor U5263 (N_5263,N_3571,N_3741);
or U5264 (N_5264,N_4251,N_3167);
xnor U5265 (N_5265,N_3653,N_3250);
and U5266 (N_5266,N_3537,N_3351);
nor U5267 (N_5267,N_4079,N_4289);
nor U5268 (N_5268,N_3901,N_3333);
or U5269 (N_5269,N_3139,N_3494);
nor U5270 (N_5270,N_3900,N_3115);
nor U5271 (N_5271,N_4112,N_3716);
xor U5272 (N_5272,N_3170,N_3036);
nand U5273 (N_5273,N_3017,N_3407);
and U5274 (N_5274,N_3199,N_4204);
or U5275 (N_5275,N_3088,N_3490);
nand U5276 (N_5276,N_3146,N_3982);
and U5277 (N_5277,N_3325,N_4469);
nand U5278 (N_5278,N_4482,N_3961);
or U5279 (N_5279,N_3197,N_3377);
xnor U5280 (N_5280,N_3592,N_4027);
nand U5281 (N_5281,N_4116,N_4222);
nand U5282 (N_5282,N_4335,N_3086);
nand U5283 (N_5283,N_4055,N_4249);
xnor U5284 (N_5284,N_4086,N_4395);
nand U5285 (N_5285,N_3547,N_3564);
xor U5286 (N_5286,N_3768,N_4009);
nor U5287 (N_5287,N_3842,N_3885);
nand U5288 (N_5288,N_3781,N_3700);
nor U5289 (N_5289,N_4317,N_3847);
and U5290 (N_5290,N_3675,N_3440);
or U5291 (N_5291,N_4279,N_3573);
nand U5292 (N_5292,N_4064,N_3026);
and U5293 (N_5293,N_3255,N_3762);
or U5294 (N_5294,N_3757,N_3906);
or U5295 (N_5295,N_3117,N_3630);
or U5296 (N_5296,N_4196,N_3440);
or U5297 (N_5297,N_3155,N_3870);
or U5298 (N_5298,N_3851,N_3037);
nand U5299 (N_5299,N_3175,N_3320);
nand U5300 (N_5300,N_4011,N_3042);
nand U5301 (N_5301,N_3802,N_3877);
xnor U5302 (N_5302,N_3368,N_3520);
nand U5303 (N_5303,N_3805,N_3493);
xnor U5304 (N_5304,N_3117,N_3200);
nor U5305 (N_5305,N_3175,N_3946);
xor U5306 (N_5306,N_3677,N_3797);
nor U5307 (N_5307,N_3277,N_3076);
or U5308 (N_5308,N_3925,N_3924);
and U5309 (N_5309,N_4394,N_4200);
nor U5310 (N_5310,N_3096,N_4383);
nor U5311 (N_5311,N_4016,N_4092);
nor U5312 (N_5312,N_4287,N_4389);
nor U5313 (N_5313,N_3980,N_3033);
xnor U5314 (N_5314,N_3454,N_4090);
nor U5315 (N_5315,N_3130,N_4499);
or U5316 (N_5316,N_4291,N_3708);
and U5317 (N_5317,N_4301,N_3311);
or U5318 (N_5318,N_4098,N_3154);
nor U5319 (N_5319,N_3406,N_3950);
or U5320 (N_5320,N_3597,N_3561);
and U5321 (N_5321,N_3207,N_3139);
nor U5322 (N_5322,N_4374,N_4321);
nor U5323 (N_5323,N_3875,N_3722);
or U5324 (N_5324,N_3383,N_3847);
or U5325 (N_5325,N_4188,N_3795);
and U5326 (N_5326,N_3839,N_4282);
and U5327 (N_5327,N_3902,N_3818);
xnor U5328 (N_5328,N_3622,N_3370);
xnor U5329 (N_5329,N_3154,N_4121);
and U5330 (N_5330,N_3614,N_3516);
nor U5331 (N_5331,N_3816,N_4319);
or U5332 (N_5332,N_4118,N_3721);
nand U5333 (N_5333,N_4442,N_3986);
nor U5334 (N_5334,N_3574,N_3611);
nor U5335 (N_5335,N_3324,N_3158);
nor U5336 (N_5336,N_3964,N_3505);
xor U5337 (N_5337,N_4312,N_4258);
or U5338 (N_5338,N_4309,N_4117);
xnor U5339 (N_5339,N_3482,N_4159);
nor U5340 (N_5340,N_4393,N_4439);
or U5341 (N_5341,N_4096,N_3778);
or U5342 (N_5342,N_3699,N_3564);
nor U5343 (N_5343,N_4292,N_3888);
or U5344 (N_5344,N_4391,N_4469);
and U5345 (N_5345,N_3961,N_3439);
and U5346 (N_5346,N_4038,N_3086);
nor U5347 (N_5347,N_4007,N_4059);
or U5348 (N_5348,N_4449,N_4280);
nor U5349 (N_5349,N_3923,N_3050);
nor U5350 (N_5350,N_3528,N_4469);
and U5351 (N_5351,N_3377,N_3743);
or U5352 (N_5352,N_3420,N_3248);
xnor U5353 (N_5353,N_3407,N_4293);
nand U5354 (N_5354,N_4094,N_3777);
xnor U5355 (N_5355,N_3393,N_4406);
xnor U5356 (N_5356,N_3960,N_3972);
and U5357 (N_5357,N_4111,N_3196);
nand U5358 (N_5358,N_3553,N_3325);
nand U5359 (N_5359,N_4279,N_4301);
nor U5360 (N_5360,N_3662,N_3139);
nand U5361 (N_5361,N_4306,N_3796);
nor U5362 (N_5362,N_3503,N_4050);
nor U5363 (N_5363,N_3155,N_4143);
nand U5364 (N_5364,N_3778,N_3971);
nor U5365 (N_5365,N_3698,N_3927);
nor U5366 (N_5366,N_4242,N_4000);
or U5367 (N_5367,N_4203,N_3331);
or U5368 (N_5368,N_3074,N_4258);
nor U5369 (N_5369,N_4234,N_3367);
and U5370 (N_5370,N_3639,N_3010);
and U5371 (N_5371,N_3491,N_4100);
or U5372 (N_5372,N_3692,N_3641);
nor U5373 (N_5373,N_3722,N_4193);
nor U5374 (N_5374,N_3864,N_4447);
nor U5375 (N_5375,N_3588,N_4167);
or U5376 (N_5376,N_3060,N_4423);
xnor U5377 (N_5377,N_3324,N_3297);
nor U5378 (N_5378,N_3589,N_3310);
xnor U5379 (N_5379,N_3942,N_3018);
or U5380 (N_5380,N_3973,N_3750);
nor U5381 (N_5381,N_3154,N_3377);
and U5382 (N_5382,N_3522,N_3814);
nor U5383 (N_5383,N_4380,N_3684);
and U5384 (N_5384,N_3367,N_3075);
xnor U5385 (N_5385,N_3383,N_4224);
nor U5386 (N_5386,N_4357,N_4093);
or U5387 (N_5387,N_3162,N_3687);
or U5388 (N_5388,N_3002,N_4345);
or U5389 (N_5389,N_3979,N_3706);
or U5390 (N_5390,N_4063,N_3259);
xor U5391 (N_5391,N_4142,N_3022);
xnor U5392 (N_5392,N_3646,N_3692);
xnor U5393 (N_5393,N_3807,N_3563);
or U5394 (N_5394,N_3354,N_3276);
and U5395 (N_5395,N_3850,N_4129);
nor U5396 (N_5396,N_3653,N_3707);
and U5397 (N_5397,N_3647,N_3954);
or U5398 (N_5398,N_4085,N_4038);
and U5399 (N_5399,N_3438,N_3618);
or U5400 (N_5400,N_3515,N_4296);
nand U5401 (N_5401,N_4495,N_3931);
and U5402 (N_5402,N_4107,N_3579);
nand U5403 (N_5403,N_4419,N_3576);
nor U5404 (N_5404,N_4135,N_4497);
nand U5405 (N_5405,N_4333,N_3769);
and U5406 (N_5406,N_3967,N_3555);
or U5407 (N_5407,N_3154,N_4017);
or U5408 (N_5408,N_4400,N_3327);
nor U5409 (N_5409,N_3290,N_3792);
or U5410 (N_5410,N_3052,N_3811);
nor U5411 (N_5411,N_3038,N_3066);
xor U5412 (N_5412,N_3971,N_4215);
xor U5413 (N_5413,N_3770,N_4214);
nor U5414 (N_5414,N_3403,N_4088);
or U5415 (N_5415,N_3951,N_3381);
or U5416 (N_5416,N_4471,N_3608);
nor U5417 (N_5417,N_3911,N_4225);
nand U5418 (N_5418,N_3382,N_3026);
and U5419 (N_5419,N_4099,N_3018);
or U5420 (N_5420,N_3927,N_3253);
xnor U5421 (N_5421,N_3413,N_3472);
nor U5422 (N_5422,N_3487,N_3424);
and U5423 (N_5423,N_3991,N_3952);
or U5424 (N_5424,N_3675,N_4051);
xnor U5425 (N_5425,N_3595,N_3411);
and U5426 (N_5426,N_3076,N_3175);
xnor U5427 (N_5427,N_4208,N_4417);
xor U5428 (N_5428,N_3826,N_3474);
nor U5429 (N_5429,N_4000,N_4385);
and U5430 (N_5430,N_4376,N_3453);
nand U5431 (N_5431,N_3966,N_4470);
or U5432 (N_5432,N_4149,N_4411);
xnor U5433 (N_5433,N_3970,N_4233);
and U5434 (N_5434,N_4486,N_4410);
nand U5435 (N_5435,N_3328,N_4286);
xor U5436 (N_5436,N_3631,N_3749);
and U5437 (N_5437,N_4299,N_3476);
and U5438 (N_5438,N_4364,N_3483);
and U5439 (N_5439,N_4049,N_4342);
or U5440 (N_5440,N_3825,N_4331);
nand U5441 (N_5441,N_4096,N_4464);
or U5442 (N_5442,N_4116,N_3865);
nand U5443 (N_5443,N_4495,N_3981);
and U5444 (N_5444,N_3610,N_3187);
and U5445 (N_5445,N_3316,N_3810);
and U5446 (N_5446,N_4164,N_4484);
xnor U5447 (N_5447,N_3373,N_4050);
nand U5448 (N_5448,N_3922,N_4277);
and U5449 (N_5449,N_3053,N_4263);
nor U5450 (N_5450,N_4267,N_4451);
or U5451 (N_5451,N_3817,N_3710);
nor U5452 (N_5452,N_4052,N_4496);
nor U5453 (N_5453,N_4253,N_3024);
xor U5454 (N_5454,N_4133,N_3264);
and U5455 (N_5455,N_4059,N_4004);
xnor U5456 (N_5456,N_3180,N_4346);
or U5457 (N_5457,N_4322,N_4423);
xnor U5458 (N_5458,N_3416,N_3955);
or U5459 (N_5459,N_3059,N_3216);
xor U5460 (N_5460,N_3807,N_3532);
and U5461 (N_5461,N_4049,N_3075);
nand U5462 (N_5462,N_3499,N_3710);
xor U5463 (N_5463,N_3049,N_3217);
nand U5464 (N_5464,N_3206,N_3536);
xnor U5465 (N_5465,N_4465,N_3806);
nand U5466 (N_5466,N_3258,N_4270);
or U5467 (N_5467,N_3969,N_4295);
xor U5468 (N_5468,N_3609,N_3794);
xor U5469 (N_5469,N_3777,N_3980);
or U5470 (N_5470,N_3876,N_3731);
and U5471 (N_5471,N_3996,N_3485);
and U5472 (N_5472,N_3957,N_3333);
and U5473 (N_5473,N_3230,N_3689);
or U5474 (N_5474,N_4059,N_3211);
or U5475 (N_5475,N_3078,N_3559);
xnor U5476 (N_5476,N_4322,N_3754);
and U5477 (N_5477,N_4276,N_3079);
xnor U5478 (N_5478,N_3200,N_3208);
or U5479 (N_5479,N_4286,N_4497);
nor U5480 (N_5480,N_3712,N_3963);
nand U5481 (N_5481,N_3107,N_3197);
and U5482 (N_5482,N_3833,N_3503);
nor U5483 (N_5483,N_3162,N_3200);
nand U5484 (N_5484,N_3006,N_3009);
nor U5485 (N_5485,N_3169,N_3487);
nand U5486 (N_5486,N_3958,N_3562);
and U5487 (N_5487,N_4205,N_3125);
nor U5488 (N_5488,N_3914,N_4308);
and U5489 (N_5489,N_4195,N_4242);
nand U5490 (N_5490,N_4431,N_3043);
xnor U5491 (N_5491,N_3050,N_3597);
or U5492 (N_5492,N_4253,N_3146);
nor U5493 (N_5493,N_4374,N_3787);
or U5494 (N_5494,N_3123,N_4179);
and U5495 (N_5495,N_4093,N_4212);
xor U5496 (N_5496,N_3614,N_4030);
nand U5497 (N_5497,N_4142,N_4410);
nor U5498 (N_5498,N_3538,N_3248);
or U5499 (N_5499,N_3631,N_3500);
xor U5500 (N_5500,N_4231,N_3030);
and U5501 (N_5501,N_3415,N_4003);
nand U5502 (N_5502,N_4206,N_4225);
or U5503 (N_5503,N_4000,N_3356);
and U5504 (N_5504,N_3746,N_4219);
nand U5505 (N_5505,N_3006,N_3277);
xor U5506 (N_5506,N_3414,N_3299);
or U5507 (N_5507,N_3079,N_3605);
nor U5508 (N_5508,N_4103,N_4374);
and U5509 (N_5509,N_3856,N_3835);
nand U5510 (N_5510,N_3906,N_3466);
xor U5511 (N_5511,N_3171,N_4112);
and U5512 (N_5512,N_4077,N_3657);
and U5513 (N_5513,N_3598,N_4278);
nand U5514 (N_5514,N_3703,N_3760);
xor U5515 (N_5515,N_4475,N_3912);
xnor U5516 (N_5516,N_3653,N_3992);
nand U5517 (N_5517,N_4305,N_3505);
and U5518 (N_5518,N_3904,N_3750);
or U5519 (N_5519,N_3564,N_3437);
and U5520 (N_5520,N_3892,N_4006);
and U5521 (N_5521,N_3275,N_4034);
or U5522 (N_5522,N_4423,N_4012);
and U5523 (N_5523,N_3685,N_3471);
and U5524 (N_5524,N_3047,N_3016);
nor U5525 (N_5525,N_4404,N_3449);
nand U5526 (N_5526,N_3011,N_3019);
or U5527 (N_5527,N_3324,N_3591);
xor U5528 (N_5528,N_4044,N_3161);
and U5529 (N_5529,N_4499,N_3932);
and U5530 (N_5530,N_3270,N_3429);
xor U5531 (N_5531,N_3534,N_3437);
nand U5532 (N_5532,N_4353,N_3884);
xor U5533 (N_5533,N_3724,N_3739);
nor U5534 (N_5534,N_3162,N_4194);
nand U5535 (N_5535,N_3504,N_3301);
or U5536 (N_5536,N_3758,N_4342);
and U5537 (N_5537,N_3121,N_3395);
nor U5538 (N_5538,N_4353,N_4381);
or U5539 (N_5539,N_3502,N_3941);
or U5540 (N_5540,N_3979,N_3976);
and U5541 (N_5541,N_3126,N_3295);
xnor U5542 (N_5542,N_3461,N_3225);
xor U5543 (N_5543,N_4334,N_4050);
or U5544 (N_5544,N_4246,N_3593);
nand U5545 (N_5545,N_4057,N_4147);
xor U5546 (N_5546,N_3221,N_3569);
or U5547 (N_5547,N_4177,N_3779);
nor U5548 (N_5548,N_3092,N_4320);
and U5549 (N_5549,N_3622,N_3118);
and U5550 (N_5550,N_4440,N_3760);
nor U5551 (N_5551,N_4042,N_3250);
nor U5552 (N_5552,N_3595,N_4170);
and U5553 (N_5553,N_3250,N_3737);
or U5554 (N_5554,N_3823,N_3448);
and U5555 (N_5555,N_3630,N_3171);
or U5556 (N_5556,N_3726,N_3883);
nor U5557 (N_5557,N_4008,N_4416);
xor U5558 (N_5558,N_3890,N_3389);
nand U5559 (N_5559,N_3285,N_4345);
or U5560 (N_5560,N_3490,N_3894);
nand U5561 (N_5561,N_4480,N_3373);
nand U5562 (N_5562,N_4268,N_3468);
nor U5563 (N_5563,N_4332,N_3242);
and U5564 (N_5564,N_3734,N_4017);
nand U5565 (N_5565,N_4447,N_3344);
nand U5566 (N_5566,N_3228,N_4401);
nand U5567 (N_5567,N_4231,N_3887);
nor U5568 (N_5568,N_4408,N_3471);
nand U5569 (N_5569,N_3396,N_3180);
or U5570 (N_5570,N_4385,N_3921);
and U5571 (N_5571,N_3273,N_3175);
nand U5572 (N_5572,N_3661,N_4447);
and U5573 (N_5573,N_3686,N_3131);
xor U5574 (N_5574,N_4199,N_3686);
or U5575 (N_5575,N_4402,N_4127);
or U5576 (N_5576,N_3277,N_3784);
nand U5577 (N_5577,N_3502,N_3736);
nand U5578 (N_5578,N_4369,N_3795);
nor U5579 (N_5579,N_4127,N_4173);
or U5580 (N_5580,N_3667,N_3414);
nand U5581 (N_5581,N_3032,N_4467);
nor U5582 (N_5582,N_3737,N_4438);
or U5583 (N_5583,N_3159,N_3725);
nand U5584 (N_5584,N_4256,N_3050);
and U5585 (N_5585,N_3295,N_4412);
xor U5586 (N_5586,N_3325,N_3022);
xor U5587 (N_5587,N_3288,N_3665);
nand U5588 (N_5588,N_3445,N_3087);
or U5589 (N_5589,N_3723,N_4405);
or U5590 (N_5590,N_3300,N_4396);
nand U5591 (N_5591,N_3796,N_3503);
or U5592 (N_5592,N_4434,N_4220);
and U5593 (N_5593,N_3999,N_3274);
or U5594 (N_5594,N_3567,N_3371);
and U5595 (N_5595,N_3675,N_3876);
nor U5596 (N_5596,N_3590,N_4259);
xnor U5597 (N_5597,N_3340,N_3062);
nand U5598 (N_5598,N_3478,N_3108);
nand U5599 (N_5599,N_4490,N_3147);
nor U5600 (N_5600,N_3358,N_4426);
nor U5601 (N_5601,N_4160,N_4251);
nor U5602 (N_5602,N_3695,N_3684);
xor U5603 (N_5603,N_3758,N_3837);
nand U5604 (N_5604,N_3028,N_4058);
and U5605 (N_5605,N_3185,N_4335);
xor U5606 (N_5606,N_4065,N_4240);
and U5607 (N_5607,N_3695,N_3624);
xor U5608 (N_5608,N_3854,N_4096);
and U5609 (N_5609,N_4219,N_3522);
and U5610 (N_5610,N_3225,N_3958);
nor U5611 (N_5611,N_4420,N_3363);
nand U5612 (N_5612,N_3989,N_4123);
xnor U5613 (N_5613,N_3812,N_3005);
or U5614 (N_5614,N_3425,N_3550);
xor U5615 (N_5615,N_3276,N_3093);
xor U5616 (N_5616,N_4342,N_4126);
nand U5617 (N_5617,N_4155,N_4091);
or U5618 (N_5618,N_3422,N_3629);
xor U5619 (N_5619,N_3130,N_3358);
and U5620 (N_5620,N_3734,N_3322);
xor U5621 (N_5621,N_3226,N_4449);
nand U5622 (N_5622,N_4132,N_4418);
or U5623 (N_5623,N_3057,N_4411);
or U5624 (N_5624,N_3175,N_3197);
nand U5625 (N_5625,N_3541,N_3386);
nand U5626 (N_5626,N_3917,N_3723);
nand U5627 (N_5627,N_3966,N_3147);
and U5628 (N_5628,N_3222,N_3999);
xor U5629 (N_5629,N_3749,N_3998);
xor U5630 (N_5630,N_3726,N_3506);
nand U5631 (N_5631,N_4223,N_3473);
xnor U5632 (N_5632,N_4435,N_3540);
xnor U5633 (N_5633,N_4035,N_3022);
or U5634 (N_5634,N_4299,N_4144);
xnor U5635 (N_5635,N_3258,N_4020);
and U5636 (N_5636,N_3859,N_3052);
xor U5637 (N_5637,N_3385,N_4191);
and U5638 (N_5638,N_3912,N_4481);
or U5639 (N_5639,N_3333,N_4364);
nand U5640 (N_5640,N_3430,N_3337);
or U5641 (N_5641,N_3418,N_3629);
xor U5642 (N_5642,N_3158,N_3351);
xnor U5643 (N_5643,N_4294,N_3119);
nand U5644 (N_5644,N_3345,N_3910);
nor U5645 (N_5645,N_3074,N_3416);
nor U5646 (N_5646,N_3841,N_4039);
nand U5647 (N_5647,N_3668,N_3253);
nor U5648 (N_5648,N_3031,N_3140);
xnor U5649 (N_5649,N_4243,N_3076);
or U5650 (N_5650,N_3021,N_3527);
or U5651 (N_5651,N_3605,N_3889);
nor U5652 (N_5652,N_4396,N_3860);
xnor U5653 (N_5653,N_3230,N_3374);
or U5654 (N_5654,N_3285,N_4057);
nand U5655 (N_5655,N_3126,N_3562);
and U5656 (N_5656,N_3500,N_3184);
xnor U5657 (N_5657,N_3391,N_3978);
nor U5658 (N_5658,N_3226,N_3299);
nand U5659 (N_5659,N_3181,N_4306);
or U5660 (N_5660,N_3641,N_4460);
xnor U5661 (N_5661,N_3053,N_4285);
xor U5662 (N_5662,N_4296,N_4096);
or U5663 (N_5663,N_4425,N_3847);
and U5664 (N_5664,N_3665,N_3681);
or U5665 (N_5665,N_3552,N_3565);
and U5666 (N_5666,N_3444,N_3593);
nand U5667 (N_5667,N_3950,N_3410);
and U5668 (N_5668,N_4480,N_4222);
or U5669 (N_5669,N_3254,N_3940);
nand U5670 (N_5670,N_3963,N_4311);
nand U5671 (N_5671,N_4203,N_3302);
nand U5672 (N_5672,N_3957,N_3928);
nor U5673 (N_5673,N_3866,N_3222);
and U5674 (N_5674,N_3462,N_4434);
nand U5675 (N_5675,N_4215,N_3516);
nor U5676 (N_5676,N_3915,N_3880);
and U5677 (N_5677,N_3228,N_3114);
nor U5678 (N_5678,N_3408,N_3625);
and U5679 (N_5679,N_3944,N_3454);
or U5680 (N_5680,N_3776,N_3274);
and U5681 (N_5681,N_4498,N_4055);
or U5682 (N_5682,N_3053,N_4406);
nand U5683 (N_5683,N_3592,N_3746);
nor U5684 (N_5684,N_4215,N_3051);
xor U5685 (N_5685,N_3477,N_3581);
xor U5686 (N_5686,N_4034,N_3987);
and U5687 (N_5687,N_3288,N_3338);
nand U5688 (N_5688,N_4018,N_3147);
nor U5689 (N_5689,N_3022,N_3651);
xnor U5690 (N_5690,N_3611,N_3552);
xor U5691 (N_5691,N_3053,N_3898);
and U5692 (N_5692,N_4304,N_4102);
xor U5693 (N_5693,N_3865,N_4337);
nand U5694 (N_5694,N_4439,N_3604);
nand U5695 (N_5695,N_3443,N_3397);
and U5696 (N_5696,N_4317,N_4148);
xnor U5697 (N_5697,N_3332,N_4179);
nor U5698 (N_5698,N_3168,N_3529);
nor U5699 (N_5699,N_4454,N_3716);
xor U5700 (N_5700,N_4181,N_4272);
nor U5701 (N_5701,N_3906,N_3281);
xnor U5702 (N_5702,N_4376,N_3156);
nor U5703 (N_5703,N_3627,N_3237);
nand U5704 (N_5704,N_3379,N_4194);
nand U5705 (N_5705,N_3835,N_3421);
nand U5706 (N_5706,N_4154,N_4178);
nand U5707 (N_5707,N_3433,N_4313);
nor U5708 (N_5708,N_4297,N_3783);
nand U5709 (N_5709,N_4429,N_3171);
nand U5710 (N_5710,N_3830,N_3380);
nand U5711 (N_5711,N_3184,N_4080);
nor U5712 (N_5712,N_4324,N_4373);
nor U5713 (N_5713,N_4104,N_4280);
and U5714 (N_5714,N_3189,N_3251);
or U5715 (N_5715,N_4298,N_3539);
nand U5716 (N_5716,N_3633,N_4321);
or U5717 (N_5717,N_3780,N_4257);
nand U5718 (N_5718,N_3780,N_3337);
nand U5719 (N_5719,N_4007,N_3387);
and U5720 (N_5720,N_4253,N_3777);
xnor U5721 (N_5721,N_3112,N_3835);
nand U5722 (N_5722,N_3409,N_3939);
or U5723 (N_5723,N_3267,N_3634);
or U5724 (N_5724,N_3413,N_3079);
nand U5725 (N_5725,N_4196,N_3238);
or U5726 (N_5726,N_4403,N_3841);
and U5727 (N_5727,N_3107,N_3997);
xnor U5728 (N_5728,N_3989,N_3535);
xnor U5729 (N_5729,N_3825,N_3055);
xor U5730 (N_5730,N_3991,N_3677);
and U5731 (N_5731,N_3460,N_3082);
xnor U5732 (N_5732,N_4270,N_3924);
or U5733 (N_5733,N_3238,N_3867);
xor U5734 (N_5734,N_3768,N_4457);
nand U5735 (N_5735,N_4389,N_4132);
nand U5736 (N_5736,N_4292,N_3454);
nor U5737 (N_5737,N_3380,N_3117);
xor U5738 (N_5738,N_3809,N_3095);
xnor U5739 (N_5739,N_4060,N_3837);
xnor U5740 (N_5740,N_3786,N_3080);
nand U5741 (N_5741,N_4125,N_3838);
xnor U5742 (N_5742,N_3156,N_3341);
nand U5743 (N_5743,N_3916,N_3666);
or U5744 (N_5744,N_4102,N_3447);
nor U5745 (N_5745,N_3322,N_3024);
or U5746 (N_5746,N_4203,N_3004);
nand U5747 (N_5747,N_3155,N_3395);
xnor U5748 (N_5748,N_4096,N_3868);
and U5749 (N_5749,N_3447,N_4304);
nand U5750 (N_5750,N_3233,N_4458);
or U5751 (N_5751,N_4121,N_3096);
nor U5752 (N_5752,N_3118,N_4446);
nand U5753 (N_5753,N_4070,N_3747);
nor U5754 (N_5754,N_4112,N_3444);
or U5755 (N_5755,N_3996,N_3805);
xor U5756 (N_5756,N_4074,N_4395);
nor U5757 (N_5757,N_3540,N_4143);
nor U5758 (N_5758,N_4018,N_3977);
and U5759 (N_5759,N_4164,N_4017);
nor U5760 (N_5760,N_3582,N_3872);
nand U5761 (N_5761,N_3772,N_3531);
xor U5762 (N_5762,N_3366,N_4481);
or U5763 (N_5763,N_4365,N_4174);
nand U5764 (N_5764,N_3389,N_3241);
nand U5765 (N_5765,N_4331,N_3568);
or U5766 (N_5766,N_3366,N_3802);
xor U5767 (N_5767,N_3111,N_3092);
or U5768 (N_5768,N_3798,N_3519);
or U5769 (N_5769,N_3932,N_4434);
and U5770 (N_5770,N_3988,N_3668);
xnor U5771 (N_5771,N_3721,N_3929);
nand U5772 (N_5772,N_4300,N_3984);
and U5773 (N_5773,N_3234,N_4060);
nand U5774 (N_5774,N_3180,N_3635);
nand U5775 (N_5775,N_3689,N_3493);
nand U5776 (N_5776,N_4145,N_3381);
nand U5777 (N_5777,N_3105,N_4040);
nor U5778 (N_5778,N_4352,N_3424);
nand U5779 (N_5779,N_4094,N_3377);
and U5780 (N_5780,N_3167,N_3939);
xor U5781 (N_5781,N_3283,N_3196);
xor U5782 (N_5782,N_3005,N_3496);
nand U5783 (N_5783,N_3136,N_4406);
or U5784 (N_5784,N_3137,N_3985);
xor U5785 (N_5785,N_4489,N_3111);
nor U5786 (N_5786,N_3755,N_3630);
nor U5787 (N_5787,N_3987,N_3823);
xnor U5788 (N_5788,N_4294,N_3190);
nor U5789 (N_5789,N_4309,N_3610);
and U5790 (N_5790,N_4342,N_3084);
nor U5791 (N_5791,N_4141,N_3057);
xnor U5792 (N_5792,N_3173,N_4097);
nor U5793 (N_5793,N_3958,N_4376);
or U5794 (N_5794,N_3864,N_3649);
nand U5795 (N_5795,N_3594,N_4220);
xnor U5796 (N_5796,N_3492,N_4245);
nand U5797 (N_5797,N_4371,N_4428);
or U5798 (N_5798,N_4269,N_3637);
nor U5799 (N_5799,N_4298,N_3989);
nand U5800 (N_5800,N_3663,N_4294);
or U5801 (N_5801,N_3036,N_3715);
and U5802 (N_5802,N_3053,N_4299);
or U5803 (N_5803,N_3927,N_3215);
xor U5804 (N_5804,N_3999,N_4316);
xor U5805 (N_5805,N_3315,N_4116);
and U5806 (N_5806,N_3952,N_3436);
and U5807 (N_5807,N_3915,N_3309);
and U5808 (N_5808,N_3004,N_4206);
xnor U5809 (N_5809,N_4074,N_4133);
nor U5810 (N_5810,N_3744,N_3101);
and U5811 (N_5811,N_3437,N_4107);
and U5812 (N_5812,N_4437,N_3738);
nand U5813 (N_5813,N_4228,N_3609);
xnor U5814 (N_5814,N_4074,N_3918);
or U5815 (N_5815,N_3615,N_4042);
nand U5816 (N_5816,N_4308,N_3874);
nand U5817 (N_5817,N_4479,N_3837);
nand U5818 (N_5818,N_3967,N_4062);
xor U5819 (N_5819,N_3467,N_3623);
nor U5820 (N_5820,N_4128,N_3480);
nor U5821 (N_5821,N_3252,N_3901);
and U5822 (N_5822,N_3008,N_4416);
and U5823 (N_5823,N_4261,N_3962);
nand U5824 (N_5824,N_3687,N_4241);
nand U5825 (N_5825,N_3057,N_3565);
and U5826 (N_5826,N_3163,N_3856);
and U5827 (N_5827,N_4157,N_3130);
or U5828 (N_5828,N_3133,N_3982);
nor U5829 (N_5829,N_3251,N_3604);
and U5830 (N_5830,N_3888,N_3926);
nand U5831 (N_5831,N_4423,N_3371);
nor U5832 (N_5832,N_3180,N_3100);
nand U5833 (N_5833,N_4399,N_4306);
and U5834 (N_5834,N_3066,N_4218);
and U5835 (N_5835,N_3216,N_3101);
nor U5836 (N_5836,N_4251,N_3835);
or U5837 (N_5837,N_3778,N_4264);
nor U5838 (N_5838,N_3899,N_3619);
or U5839 (N_5839,N_3057,N_3242);
nand U5840 (N_5840,N_3186,N_3093);
or U5841 (N_5841,N_3795,N_3715);
xnor U5842 (N_5842,N_4359,N_4027);
or U5843 (N_5843,N_3426,N_4277);
or U5844 (N_5844,N_4149,N_3231);
nor U5845 (N_5845,N_3274,N_4362);
xor U5846 (N_5846,N_3632,N_3946);
or U5847 (N_5847,N_3548,N_4343);
or U5848 (N_5848,N_3122,N_4055);
nand U5849 (N_5849,N_3438,N_3624);
and U5850 (N_5850,N_3737,N_4174);
nand U5851 (N_5851,N_3716,N_4041);
xor U5852 (N_5852,N_4037,N_3715);
nor U5853 (N_5853,N_3015,N_3292);
nor U5854 (N_5854,N_3022,N_3645);
nand U5855 (N_5855,N_3135,N_4008);
nor U5856 (N_5856,N_3429,N_3024);
nor U5857 (N_5857,N_3514,N_4417);
xor U5858 (N_5858,N_3410,N_3615);
nand U5859 (N_5859,N_4099,N_3283);
nor U5860 (N_5860,N_4400,N_3003);
or U5861 (N_5861,N_3160,N_4312);
or U5862 (N_5862,N_4362,N_3868);
nand U5863 (N_5863,N_4408,N_3725);
nor U5864 (N_5864,N_3536,N_3025);
and U5865 (N_5865,N_4000,N_3976);
xnor U5866 (N_5866,N_3458,N_3852);
or U5867 (N_5867,N_4480,N_4498);
nor U5868 (N_5868,N_3466,N_3233);
nor U5869 (N_5869,N_4426,N_3576);
nor U5870 (N_5870,N_3626,N_4426);
or U5871 (N_5871,N_4421,N_3014);
nand U5872 (N_5872,N_3199,N_4186);
nor U5873 (N_5873,N_4487,N_3874);
and U5874 (N_5874,N_3149,N_4226);
xnor U5875 (N_5875,N_4180,N_3632);
xor U5876 (N_5876,N_4066,N_4491);
nand U5877 (N_5877,N_3755,N_3895);
nor U5878 (N_5878,N_3912,N_3997);
and U5879 (N_5879,N_4325,N_3677);
and U5880 (N_5880,N_4177,N_3398);
nor U5881 (N_5881,N_3302,N_3988);
xnor U5882 (N_5882,N_3130,N_3225);
or U5883 (N_5883,N_3716,N_3503);
nor U5884 (N_5884,N_3337,N_3530);
nor U5885 (N_5885,N_3297,N_3873);
nor U5886 (N_5886,N_3707,N_3127);
xor U5887 (N_5887,N_3643,N_4136);
and U5888 (N_5888,N_3997,N_4289);
xnor U5889 (N_5889,N_3063,N_3942);
and U5890 (N_5890,N_3972,N_3210);
or U5891 (N_5891,N_4011,N_3289);
nor U5892 (N_5892,N_4364,N_3840);
nor U5893 (N_5893,N_3082,N_4298);
and U5894 (N_5894,N_3799,N_3057);
nor U5895 (N_5895,N_4386,N_3807);
or U5896 (N_5896,N_4148,N_3841);
nand U5897 (N_5897,N_3520,N_4297);
nand U5898 (N_5898,N_3387,N_3155);
nand U5899 (N_5899,N_3233,N_3804);
nand U5900 (N_5900,N_3832,N_3998);
nand U5901 (N_5901,N_3439,N_3846);
xnor U5902 (N_5902,N_4421,N_3839);
xor U5903 (N_5903,N_3834,N_3976);
and U5904 (N_5904,N_4382,N_3566);
xnor U5905 (N_5905,N_4294,N_3049);
and U5906 (N_5906,N_3859,N_3365);
or U5907 (N_5907,N_3729,N_4155);
or U5908 (N_5908,N_3071,N_4136);
nand U5909 (N_5909,N_3691,N_3965);
nand U5910 (N_5910,N_4008,N_3454);
nor U5911 (N_5911,N_3582,N_3659);
and U5912 (N_5912,N_3943,N_3651);
xnor U5913 (N_5913,N_3682,N_4386);
nor U5914 (N_5914,N_3131,N_3543);
or U5915 (N_5915,N_4107,N_3317);
nand U5916 (N_5916,N_3544,N_4491);
xnor U5917 (N_5917,N_3960,N_3998);
nor U5918 (N_5918,N_3182,N_4494);
nand U5919 (N_5919,N_4028,N_4352);
nor U5920 (N_5920,N_3566,N_3104);
nor U5921 (N_5921,N_4406,N_3992);
nor U5922 (N_5922,N_3350,N_3092);
nand U5923 (N_5923,N_4447,N_4411);
nor U5924 (N_5924,N_4105,N_3945);
nor U5925 (N_5925,N_3867,N_3321);
nand U5926 (N_5926,N_4013,N_3775);
or U5927 (N_5927,N_3860,N_3698);
nand U5928 (N_5928,N_3546,N_3816);
nor U5929 (N_5929,N_3456,N_4240);
nor U5930 (N_5930,N_4397,N_3456);
nor U5931 (N_5931,N_3701,N_3762);
xor U5932 (N_5932,N_3039,N_3553);
nor U5933 (N_5933,N_3772,N_4229);
nor U5934 (N_5934,N_4375,N_3147);
and U5935 (N_5935,N_3157,N_3323);
xnor U5936 (N_5936,N_4214,N_4378);
nand U5937 (N_5937,N_3364,N_3224);
xor U5938 (N_5938,N_3049,N_3426);
nand U5939 (N_5939,N_3174,N_3227);
and U5940 (N_5940,N_3275,N_3345);
nand U5941 (N_5941,N_3769,N_3587);
nor U5942 (N_5942,N_4307,N_3548);
nor U5943 (N_5943,N_4088,N_4412);
xor U5944 (N_5944,N_3319,N_4005);
and U5945 (N_5945,N_3877,N_3183);
nor U5946 (N_5946,N_3984,N_3460);
or U5947 (N_5947,N_3143,N_3222);
or U5948 (N_5948,N_3408,N_3330);
or U5949 (N_5949,N_3426,N_3164);
and U5950 (N_5950,N_3547,N_4018);
or U5951 (N_5951,N_3288,N_3227);
or U5952 (N_5952,N_3285,N_4058);
nor U5953 (N_5953,N_3117,N_3944);
and U5954 (N_5954,N_3094,N_3353);
or U5955 (N_5955,N_3953,N_4299);
or U5956 (N_5956,N_4210,N_3881);
xnor U5957 (N_5957,N_3948,N_3063);
nor U5958 (N_5958,N_4441,N_3903);
xnor U5959 (N_5959,N_4142,N_4158);
xnor U5960 (N_5960,N_3681,N_3659);
nand U5961 (N_5961,N_4400,N_3829);
xnor U5962 (N_5962,N_3850,N_4013);
and U5963 (N_5963,N_4064,N_3083);
nor U5964 (N_5964,N_3565,N_3622);
xor U5965 (N_5965,N_3560,N_4452);
nor U5966 (N_5966,N_4486,N_4104);
or U5967 (N_5967,N_3738,N_4475);
nor U5968 (N_5968,N_3940,N_3676);
or U5969 (N_5969,N_4394,N_4451);
and U5970 (N_5970,N_4354,N_3295);
or U5971 (N_5971,N_3420,N_3718);
nor U5972 (N_5972,N_3560,N_3734);
and U5973 (N_5973,N_3409,N_4342);
and U5974 (N_5974,N_4451,N_3713);
nor U5975 (N_5975,N_3805,N_3332);
or U5976 (N_5976,N_3823,N_4222);
and U5977 (N_5977,N_3800,N_3494);
xnor U5978 (N_5978,N_3329,N_3898);
or U5979 (N_5979,N_3389,N_4242);
and U5980 (N_5980,N_3001,N_3003);
xor U5981 (N_5981,N_4215,N_3526);
or U5982 (N_5982,N_3690,N_4099);
nand U5983 (N_5983,N_3354,N_3812);
nand U5984 (N_5984,N_3232,N_3228);
or U5985 (N_5985,N_4086,N_3876);
or U5986 (N_5986,N_3889,N_3226);
or U5987 (N_5987,N_3369,N_4241);
and U5988 (N_5988,N_3085,N_3754);
xnor U5989 (N_5989,N_4309,N_4064);
xnor U5990 (N_5990,N_4344,N_4221);
nand U5991 (N_5991,N_3364,N_3674);
and U5992 (N_5992,N_3820,N_4388);
and U5993 (N_5993,N_3884,N_3212);
xnor U5994 (N_5994,N_3350,N_4177);
xor U5995 (N_5995,N_4466,N_4080);
nor U5996 (N_5996,N_3542,N_3565);
or U5997 (N_5997,N_4362,N_3736);
and U5998 (N_5998,N_4076,N_3268);
nor U5999 (N_5999,N_3206,N_3800);
and U6000 (N_6000,N_5615,N_5460);
nand U6001 (N_6001,N_5556,N_5516);
nand U6002 (N_6002,N_5465,N_5273);
or U6003 (N_6003,N_5474,N_4758);
or U6004 (N_6004,N_4593,N_5950);
nor U6005 (N_6005,N_5498,N_5094);
xnor U6006 (N_6006,N_5937,N_4917);
xor U6007 (N_6007,N_4509,N_5590);
nand U6008 (N_6008,N_5877,N_4609);
and U6009 (N_6009,N_5960,N_5352);
or U6010 (N_6010,N_5632,N_5593);
nand U6011 (N_6011,N_5411,N_5421);
xor U6012 (N_6012,N_4994,N_5437);
xnor U6013 (N_6013,N_4781,N_4576);
nor U6014 (N_6014,N_5161,N_5467);
xor U6015 (N_6015,N_5767,N_4881);
nand U6016 (N_6016,N_4908,N_4885);
or U6017 (N_6017,N_4860,N_5799);
nand U6018 (N_6018,N_5662,N_5745);
or U6019 (N_6019,N_5637,N_4633);
and U6020 (N_6020,N_5609,N_5842);
nor U6021 (N_6021,N_5654,N_4963);
and U6022 (N_6022,N_5359,N_5093);
nor U6023 (N_6023,N_4699,N_5688);
or U6024 (N_6024,N_5521,N_5869);
nor U6025 (N_6025,N_5451,N_5680);
nand U6026 (N_6026,N_4500,N_4669);
nand U6027 (N_6027,N_4537,N_4899);
or U6028 (N_6028,N_5969,N_5202);
xor U6029 (N_6029,N_4681,N_4978);
nand U6030 (N_6030,N_5364,N_5413);
xor U6031 (N_6031,N_5630,N_5362);
nor U6032 (N_6032,N_5208,N_5019);
nor U6033 (N_6033,N_5222,N_5007);
or U6034 (N_6034,N_5552,N_5509);
xor U6035 (N_6035,N_5901,N_4897);
nand U6036 (N_6036,N_5756,N_4754);
or U6037 (N_6037,N_5572,N_4878);
xor U6038 (N_6038,N_5712,N_5714);
xor U6039 (N_6039,N_5732,N_5984);
nand U6040 (N_6040,N_5097,N_5720);
and U6041 (N_6041,N_4722,N_4560);
and U6042 (N_6042,N_5043,N_5887);
nand U6043 (N_6043,N_5049,N_5929);
and U6044 (N_6044,N_5059,N_4698);
and U6045 (N_6045,N_5039,N_4735);
nor U6046 (N_6046,N_5428,N_5271);
or U6047 (N_6047,N_5782,N_5321);
nand U6048 (N_6048,N_5484,N_4588);
and U6049 (N_6049,N_5227,N_5213);
nand U6050 (N_6050,N_5963,N_4931);
xnor U6051 (N_6051,N_4721,N_5753);
nand U6052 (N_6052,N_5416,N_4896);
and U6053 (N_6053,N_4850,N_4581);
xnor U6054 (N_6054,N_5348,N_5382);
xor U6055 (N_6055,N_5709,N_5517);
xnor U6056 (N_6056,N_4523,N_5829);
nand U6057 (N_6057,N_5330,N_4515);
nor U6058 (N_6058,N_5957,N_5543);
nor U6059 (N_6059,N_5511,N_5849);
nand U6060 (N_6060,N_4997,N_5353);
xor U6061 (N_6061,N_4594,N_5973);
nor U6062 (N_6062,N_5979,N_5080);
xnor U6063 (N_6063,N_5163,N_4985);
or U6064 (N_6064,N_5325,N_5812);
nor U6065 (N_6065,N_5017,N_5880);
xor U6066 (N_6066,N_4554,N_5100);
nor U6067 (N_6067,N_5985,N_5311);
nand U6068 (N_6068,N_4519,N_5703);
nand U6069 (N_6069,N_4864,N_5324);
nor U6070 (N_6070,N_5997,N_5713);
or U6071 (N_6071,N_5586,N_4914);
and U6072 (N_6072,N_5711,N_4742);
or U6073 (N_6073,N_4779,N_5394);
nand U6074 (N_6074,N_5559,N_5351);
or U6075 (N_6075,N_5898,N_5840);
and U6076 (N_6076,N_5641,N_4506);
and U6077 (N_6077,N_4961,N_5149);
nor U6078 (N_6078,N_5810,N_5990);
or U6079 (N_6079,N_5975,N_4550);
nand U6080 (N_6080,N_5537,N_5333);
and U6081 (N_6081,N_5788,N_5482);
nor U6082 (N_6082,N_5403,N_5150);
and U6083 (N_6083,N_5101,N_4818);
or U6084 (N_6084,N_5457,N_5237);
xnor U6085 (N_6085,N_5006,N_4636);
and U6086 (N_6086,N_5073,N_5248);
and U6087 (N_6087,N_5494,N_5790);
nor U6088 (N_6088,N_4525,N_5770);
or U6089 (N_6089,N_5485,N_5759);
or U6090 (N_6090,N_5279,N_4763);
nor U6091 (N_6091,N_4549,N_4545);
or U6092 (N_6092,N_5122,N_4946);
or U6093 (N_6093,N_5553,N_5504);
nand U6094 (N_6094,N_5337,N_4949);
and U6095 (N_6095,N_4565,N_5747);
xnor U6096 (N_6096,N_5169,N_4535);
nor U6097 (N_6097,N_5156,N_5454);
xor U6098 (N_6098,N_5340,N_5468);
or U6099 (N_6099,N_5211,N_5220);
nand U6100 (N_6100,N_5653,N_5057);
nor U6101 (N_6101,N_5078,N_5589);
or U6102 (N_6102,N_4906,N_4952);
xnor U6103 (N_6103,N_5105,N_5439);
xnor U6104 (N_6104,N_5347,N_5534);
xnor U6105 (N_6105,N_5346,N_4888);
nand U6106 (N_6106,N_5107,N_5938);
or U6107 (N_6107,N_4745,N_4691);
and U6108 (N_6108,N_5328,N_4770);
nand U6109 (N_6109,N_5786,N_4579);
nand U6110 (N_6110,N_5806,N_5585);
nor U6111 (N_6111,N_5805,N_4816);
and U6112 (N_6112,N_4842,N_4834);
nor U6113 (N_6113,N_4924,N_4883);
and U6114 (N_6114,N_5447,N_4585);
xor U6115 (N_6115,N_4548,N_4959);
nand U6116 (N_6116,N_5339,N_4514);
nand U6117 (N_6117,N_4948,N_4647);
nand U6118 (N_6118,N_5133,N_5409);
and U6119 (N_6119,N_5168,N_5631);
and U6120 (N_6120,N_5299,N_5327);
nand U6121 (N_6121,N_5573,N_5594);
or U6122 (N_6122,N_5084,N_5081);
and U6123 (N_6123,N_4709,N_5866);
or U6124 (N_6124,N_5233,N_4562);
nand U6125 (N_6125,N_4760,N_5578);
or U6126 (N_6126,N_5261,N_5003);
nor U6127 (N_6127,N_5129,N_4720);
nand U6128 (N_6128,N_4811,N_5683);
nand U6129 (N_6129,N_5378,N_4992);
xnor U6130 (N_6130,N_5022,N_4582);
and U6131 (N_6131,N_5209,N_4668);
or U6132 (N_6132,N_4522,N_5913);
nand U6133 (N_6133,N_4701,N_4993);
nor U6134 (N_6134,N_5800,N_4889);
xnor U6135 (N_6135,N_4958,N_5964);
nor U6136 (N_6136,N_4655,N_5200);
nor U6137 (N_6137,N_4680,N_4704);
nand U6138 (N_6138,N_5920,N_5966);
nand U6139 (N_6139,N_5453,N_5999);
and U6140 (N_6140,N_5036,N_5496);
nor U6141 (N_6141,N_5427,N_4871);
and U6142 (N_6142,N_5157,N_5557);
nand U6143 (N_6143,N_5729,N_5981);
nand U6144 (N_6144,N_4879,N_4696);
xor U6145 (N_6145,N_5462,N_5260);
nor U6146 (N_6146,N_5531,N_4910);
nand U6147 (N_6147,N_4546,N_4640);
nor U6148 (N_6148,N_5808,N_5216);
nand U6149 (N_6149,N_4858,N_5250);
xnor U6150 (N_6150,N_5648,N_4711);
nand U6151 (N_6151,N_4945,N_5188);
nand U6152 (N_6152,N_4607,N_5197);
nand U6153 (N_6153,N_5768,N_5616);
xor U6154 (N_6154,N_5332,N_5254);
nand U6155 (N_6155,N_5180,N_5923);
nand U6156 (N_6156,N_5833,N_5655);
or U6157 (N_6157,N_4956,N_5758);
nor U6158 (N_6158,N_4942,N_5315);
xor U6159 (N_6159,N_5915,N_4969);
nor U6160 (N_6160,N_4521,N_4559);
nor U6161 (N_6161,N_5367,N_5523);
and U6162 (N_6162,N_5848,N_5158);
nor U6163 (N_6163,N_5099,N_5571);
nor U6164 (N_6164,N_5414,N_5947);
nor U6165 (N_6165,N_5604,N_5210);
and U6166 (N_6166,N_5313,N_4644);
or U6167 (N_6167,N_4915,N_4999);
xor U6168 (N_6168,N_5395,N_4977);
nand U6169 (N_6169,N_5141,N_4991);
xor U6170 (N_6170,N_4815,N_5448);
and U6171 (N_6171,N_5090,N_5173);
nor U6172 (N_6172,N_5623,N_4873);
nand U6173 (N_6173,N_5748,N_5676);
and U6174 (N_6174,N_5539,N_5846);
or U6175 (N_6175,N_5673,N_5934);
nand U6176 (N_6176,N_5961,N_5410);
nand U6177 (N_6177,N_4671,N_4557);
nand U6178 (N_6178,N_5851,N_4510);
and U6179 (N_6179,N_5251,N_5493);
or U6180 (N_6180,N_5828,N_5355);
nor U6181 (N_6181,N_4829,N_5859);
nor U6182 (N_6182,N_4662,N_4567);
and U6183 (N_6183,N_5306,N_4518);
xnor U6184 (N_6184,N_5283,N_5816);
xor U6185 (N_6185,N_5420,N_5894);
nor U6186 (N_6186,N_4789,N_5684);
or U6187 (N_6187,N_5032,N_5154);
and U6188 (N_6188,N_5567,N_5266);
nor U6189 (N_6189,N_5706,N_4836);
or U6190 (N_6190,N_4808,N_4533);
or U6191 (N_6191,N_5265,N_5948);
or U6192 (N_6192,N_4667,N_5102);
nor U6193 (N_6193,N_5137,N_4928);
and U6194 (N_6194,N_5638,N_4813);
or U6195 (N_6195,N_5582,N_4964);
nand U6196 (N_6196,N_4773,N_5972);
or U6197 (N_6197,N_5243,N_4578);
nor U6198 (N_6198,N_4654,N_5164);
nand U6199 (N_6199,N_5231,N_4979);
xor U6200 (N_6200,N_4855,N_4632);
and U6201 (N_6201,N_5384,N_5933);
and U6202 (N_6202,N_4685,N_5576);
xnor U6203 (N_6203,N_4706,N_5388);
xor U6204 (N_6204,N_4649,N_5825);
or U6205 (N_6205,N_5206,N_4817);
and U6206 (N_6206,N_4859,N_4646);
xnor U6207 (N_6207,N_5379,N_5269);
xor U6208 (N_6208,N_5000,N_5489);
or U6209 (N_6209,N_5435,N_4725);
or U6210 (N_6210,N_5693,N_5704);
or U6211 (N_6211,N_5242,N_4972);
or U6212 (N_6212,N_4622,N_5912);
or U6213 (N_6213,N_5469,N_5924);
and U6214 (N_6214,N_4987,N_4971);
xor U6215 (N_6215,N_4894,N_5148);
and U6216 (N_6216,N_5440,N_4812);
and U6217 (N_6217,N_4869,N_5323);
nand U6218 (N_6218,N_4531,N_5830);
and U6219 (N_6219,N_4672,N_4650);
or U6220 (N_6220,N_5921,N_4827);
or U6221 (N_6221,N_5766,N_5811);
or U6222 (N_6222,N_5177,N_4935);
xor U6223 (N_6223,N_4980,N_4947);
nand U6224 (N_6224,N_5499,N_4976);
and U6225 (N_6225,N_4708,N_5218);
or U6226 (N_6226,N_4785,N_5635);
nor U6227 (N_6227,N_5142,N_4605);
or U6228 (N_6228,N_4930,N_5867);
nor U6229 (N_6229,N_4762,N_4595);
or U6230 (N_6230,N_5185,N_5116);
or U6231 (N_6231,N_4503,N_5245);
nor U6232 (N_6232,N_5292,N_5500);
nor U6233 (N_6233,N_4695,N_4511);
or U6234 (N_6234,N_4921,N_5858);
and U6235 (N_6235,N_5807,N_5434);
nor U6236 (N_6236,N_4868,N_4823);
and U6237 (N_6237,N_5375,N_4538);
and U6238 (N_6238,N_5610,N_4527);
nor U6239 (N_6239,N_5138,N_5108);
nand U6240 (N_6240,N_5377,N_5383);
and U6241 (N_6241,N_5885,N_4505);
xor U6242 (N_6242,N_4625,N_5834);
or U6243 (N_6243,N_5935,N_5731);
nand U6244 (N_6244,N_4558,N_5695);
or U6245 (N_6245,N_5952,N_5796);
and U6246 (N_6246,N_5455,N_5905);
xnor U6247 (N_6247,N_5986,N_5497);
nand U6248 (N_6248,N_4875,N_5404);
nand U6249 (N_6249,N_5492,N_5502);
and U6250 (N_6250,N_5749,N_4715);
or U6251 (N_6251,N_5661,N_5183);
xnor U6252 (N_6252,N_5679,N_5244);
nand U6253 (N_6253,N_5374,N_5086);
or U6254 (N_6254,N_5916,N_4748);
xnor U6255 (N_6255,N_5646,N_5599);
xnor U6256 (N_6256,N_5575,N_4596);
and U6257 (N_6257,N_5287,N_5879);
or U6258 (N_6258,N_4601,N_5838);
nand U6259 (N_6259,N_5195,N_4995);
xor U6260 (N_6260,N_5071,N_4920);
and U6261 (N_6261,N_4670,N_4744);
xor U6262 (N_6262,N_4981,N_5368);
nor U6263 (N_6263,N_5707,N_4919);
and U6264 (N_6264,N_5182,N_4610);
nor U6265 (N_6265,N_5855,N_5886);
and U6266 (N_6266,N_4577,N_5918);
and U6267 (N_6267,N_5075,N_5344);
nand U6268 (N_6268,N_4989,N_5087);
or U6269 (N_6269,N_4792,N_5996);
nand U6270 (N_6270,N_5692,N_5350);
nand U6271 (N_6271,N_5162,N_5776);
and U6272 (N_6272,N_4737,N_4675);
and U6273 (N_6273,N_5736,N_4877);
or U6274 (N_6274,N_4790,N_5818);
nand U6275 (N_6275,N_5284,N_4966);
nor U6276 (N_6276,N_5988,N_4597);
and U6277 (N_6277,N_4892,N_5705);
nor U6278 (N_6278,N_4730,N_5878);
xor U6279 (N_6279,N_5288,N_5666);
xor U6280 (N_6280,N_5338,N_4743);
nor U6281 (N_6281,N_5167,N_5300);
and U6282 (N_6282,N_5088,N_5238);
or U6283 (N_6283,N_5798,N_4656);
xnor U6284 (N_6284,N_5402,N_5291);
and U6285 (N_6285,N_5433,N_5987);
and U6286 (N_6286,N_4922,N_5971);
xor U6287 (N_6287,N_5940,N_5405);
xor U6288 (N_6288,N_5698,N_4723);
or U6289 (N_6289,N_4974,N_4973);
nor U6290 (N_6290,N_5779,N_4824);
nand U6291 (N_6291,N_4810,N_4843);
nand U6292 (N_6292,N_4512,N_5746);
nand U6293 (N_6293,N_4738,N_5488);
and U6294 (N_6294,N_4544,N_5871);
nand U6295 (N_6295,N_5479,N_5762);
or U6296 (N_6296,N_5053,N_5664);
nor U6297 (N_6297,N_5121,N_4913);
and U6298 (N_6298,N_5184,N_5235);
or U6299 (N_6299,N_5246,N_5120);
xor U6300 (N_6300,N_5381,N_5717);
nor U6301 (N_6301,N_5312,N_5503);
or U6302 (N_6302,N_4530,N_4716);
and U6303 (N_6303,N_5289,N_5004);
nor U6304 (N_6304,N_5471,N_5780);
xor U6305 (N_6305,N_5522,N_5893);
or U6306 (N_6306,N_5742,N_5942);
nand U6307 (N_6307,N_4782,N_4587);
and U6308 (N_6308,N_4658,N_4940);
or U6309 (N_6309,N_5526,N_5970);
and U6310 (N_6310,N_4923,N_4882);
nand U6311 (N_6311,N_4733,N_5002);
and U6312 (N_6312,N_4757,N_4838);
nand U6313 (N_6313,N_5794,N_5056);
nand U6314 (N_6314,N_5380,N_5951);
nor U6315 (N_6315,N_4905,N_4661);
xor U6316 (N_6316,N_5845,N_5070);
nand U6317 (N_6317,N_4543,N_5670);
nor U6318 (N_6318,N_5547,N_4589);
and U6319 (N_6319,N_4697,N_5760);
xnor U6320 (N_6320,N_5741,N_5645);
nand U6321 (N_6321,N_4957,N_5595);
xor U6322 (N_6322,N_5215,N_5614);
nand U6323 (N_6323,N_4804,N_4944);
nand U6324 (N_6324,N_5217,N_4586);
and U6325 (N_6325,N_4682,N_4614);
nand U6326 (N_6326,N_5239,N_5761);
or U6327 (N_6327,N_5360,N_5956);
nand U6328 (N_6328,N_4890,N_5777);
and U6329 (N_6329,N_4805,N_4592);
and U6330 (N_6330,N_5995,N_5696);
xor U6331 (N_6331,N_5847,N_4844);
nor U6332 (N_6332,N_5134,N_5658);
nor U6333 (N_6333,N_5596,N_5194);
nor U6334 (N_6334,N_5681,N_5976);
or U6335 (N_6335,N_5257,N_5429);
xnor U6336 (N_6336,N_5914,N_5165);
nor U6337 (N_6337,N_5307,N_4620);
nand U6338 (N_6338,N_5015,N_5669);
nor U6339 (N_6339,N_5663,N_5345);
or U6340 (N_6340,N_5558,N_5201);
and U6341 (N_6341,N_5769,N_4541);
xnor U6342 (N_6342,N_4840,N_5065);
and U6343 (N_6343,N_5945,N_5293);
nand U6344 (N_6344,N_4955,N_5754);
and U6345 (N_6345,N_5813,N_5038);
nand U6346 (N_6346,N_4569,N_5387);
nor U6347 (N_6347,N_5560,N_5740);
or U6348 (N_6348,N_4852,N_5856);
and U6349 (N_6349,N_4604,N_5587);
nor U6350 (N_6350,N_5372,N_4925);
and U6351 (N_6351,N_4851,N_5025);
or U6352 (N_6352,N_5225,N_5668);
and U6353 (N_6353,N_4665,N_5258);
or U6354 (N_6354,N_5532,N_4561);
nand U6355 (N_6355,N_4643,N_5843);
xor U6356 (N_6356,N_4727,N_4623);
xnor U6357 (N_6357,N_5919,N_5481);
or U6358 (N_6358,N_5936,N_4825);
nor U6359 (N_6359,N_5170,N_5068);
or U6360 (N_6360,N_5054,N_4573);
xnor U6361 (N_6361,N_5487,N_4849);
nand U6362 (N_6362,N_4707,N_4756);
nor U6363 (N_6363,N_4787,N_4542);
or U6364 (N_6364,N_5702,N_4659);
or U6365 (N_6365,N_5820,N_5385);
nor U6366 (N_6366,N_4839,N_5665);
nor U6367 (N_6367,N_5308,N_5889);
nor U6368 (N_6368,N_5906,N_5675);
nor U6369 (N_6369,N_5581,N_5104);
nand U6370 (N_6370,N_5275,N_5644);
nand U6371 (N_6371,N_5021,N_4719);
xor U6372 (N_6372,N_5115,N_4903);
nor U6373 (N_6373,N_5392,N_4854);
xor U6374 (N_6374,N_4831,N_5892);
xnor U6375 (N_6375,N_5331,N_4996);
and U6376 (N_6376,N_4806,N_4602);
nand U6377 (N_6377,N_5771,N_4528);
xnor U6378 (N_6378,N_5930,N_5602);
nand U6379 (N_6379,N_4613,N_4874);
xnor U6380 (N_6380,N_5822,N_5109);
and U6381 (N_6381,N_4982,N_5114);
xor U6382 (N_6382,N_5095,N_5890);
xor U6383 (N_6383,N_5529,N_4606);
xnor U6384 (N_6384,N_5844,N_5626);
nand U6385 (N_6385,N_5044,N_5047);
or U6386 (N_6386,N_5365,N_5011);
nand U6387 (N_6387,N_4657,N_4703);
nor U6388 (N_6388,N_5309,N_5295);
nand U6389 (N_6389,N_4876,N_5391);
nand U6390 (N_6390,N_5026,N_5236);
xor U6391 (N_6391,N_5297,N_4953);
nand U6392 (N_6392,N_5659,N_4688);
or U6393 (N_6393,N_4867,N_5819);
nor U6394 (N_6394,N_5939,N_4861);
nand U6395 (N_6395,N_4778,N_5001);
or U6396 (N_6396,N_5791,N_5865);
nand U6397 (N_6397,N_5091,N_5787);
xor U6398 (N_6398,N_4962,N_5136);
and U6399 (N_6399,N_5230,N_5153);
xor U6400 (N_6400,N_5809,N_4872);
or U6401 (N_6401,N_4771,N_5320);
and U6402 (N_6402,N_4863,N_5750);
nor U6403 (N_6403,N_5601,N_4652);
xor U6404 (N_6404,N_5778,N_5296);
or U6405 (N_6405,N_5793,N_5135);
nand U6406 (N_6406,N_5827,N_4536);
and U6407 (N_6407,N_5196,N_5998);
or U6408 (N_6408,N_5821,N_5259);
xor U6409 (N_6409,N_4794,N_4988);
nor U6410 (N_6410,N_5881,N_5274);
and U6411 (N_6411,N_5256,N_5624);
nor U6412 (N_6412,N_5922,N_5804);
nand U6413 (N_6413,N_5145,N_4651);
xor U6414 (N_6414,N_5181,N_5608);
xnor U6415 (N_6415,N_4516,N_5119);
nor U6416 (N_6416,N_5398,N_5528);
or U6417 (N_6417,N_5917,N_5160);
nor U6418 (N_6418,N_4761,N_5221);
or U6419 (N_6419,N_4700,N_4570);
or U6420 (N_6420,N_5048,N_5396);
xor U6421 (N_6421,N_5249,N_5466);
and U6422 (N_6422,N_5179,N_5190);
and U6423 (N_6423,N_4630,N_5700);
and U6424 (N_6424,N_4960,N_4801);
and U6425 (N_6425,N_4753,N_5204);
and U6426 (N_6426,N_5735,N_5132);
and U6427 (N_6427,N_4786,N_5724);
and U6428 (N_6428,N_5792,N_5613);
nor U6429 (N_6429,N_5326,N_5533);
xor U6430 (N_6430,N_5408,N_4887);
xnor U6431 (N_6431,N_5035,N_5737);
nor U6432 (N_6432,N_4551,N_5450);
and U6433 (N_6433,N_5187,N_5214);
or U6434 (N_6434,N_4866,N_5010);
nand U6435 (N_6435,N_5473,N_5899);
and U6436 (N_6436,N_5322,N_5801);
nand U6437 (N_6437,N_5699,N_5861);
or U6438 (N_6438,N_4751,N_5130);
or U6439 (N_6439,N_4619,N_4783);
nor U6440 (N_6440,N_4769,N_4608);
and U6441 (N_6441,N_5728,N_5329);
nor U6442 (N_6442,N_5802,N_4970);
and U6443 (N_6443,N_4990,N_4954);
nor U6444 (N_6444,N_5535,N_4777);
xor U6445 (N_6445,N_4566,N_4984);
and U6446 (N_6446,N_5579,N_5541);
nor U6447 (N_6447,N_5076,N_4814);
and U6448 (N_6448,N_5874,N_5862);
and U6449 (N_6449,N_5824,N_5727);
nor U6450 (N_6450,N_5127,N_4616);
xnor U6451 (N_6451,N_4739,N_5667);
nand U6452 (N_6452,N_5992,N_4631);
and U6453 (N_6453,N_5089,N_5316);
or U6454 (N_6454,N_4835,N_4713);
nand U6455 (N_6455,N_5977,N_5551);
nor U6456 (N_6456,N_5954,N_5524);
and U6457 (N_6457,N_5159,N_5123);
nor U6458 (N_6458,N_4639,N_5682);
xor U6459 (N_6459,N_4927,N_5690);
or U6460 (N_6460,N_5106,N_5495);
xnor U6461 (N_6461,N_4684,N_5171);
nand U6462 (N_6462,N_5519,N_5252);
nand U6463 (N_6463,N_5478,N_5198);
or U6464 (N_6464,N_5009,N_5476);
nor U6465 (N_6465,N_5536,N_5725);
nand U6466 (N_6466,N_5041,N_5369);
or U6467 (N_6467,N_5826,N_4615);
xor U6468 (N_6468,N_5240,N_5456);
xor U6469 (N_6469,N_4621,N_4918);
nand U6470 (N_6470,N_5775,N_4502);
xor U6471 (N_6471,N_5928,N_4642);
nand U6472 (N_6472,N_5708,N_5030);
nand U6473 (N_6473,N_5949,N_5738);
and U6474 (N_6474,N_5510,N_5540);
or U6475 (N_6475,N_4853,N_5925);
or U6476 (N_6476,N_4555,N_5286);
or U6477 (N_6477,N_5904,N_5545);
nand U6478 (N_6478,N_5739,N_5464);
nor U6479 (N_6479,N_4793,N_5013);
nor U6480 (N_6480,N_4628,N_4912);
nand U6481 (N_6481,N_5390,N_4694);
and U6482 (N_6482,N_5968,N_5040);
xor U6483 (N_6483,N_5441,N_5946);
or U6484 (N_6484,N_5525,N_5219);
xor U6485 (N_6485,N_4617,N_5491);
and U6486 (N_6486,N_4513,N_5797);
or U6487 (N_6487,N_4845,N_5733);
xnor U6488 (N_6488,N_4848,N_5354);
nor U6489 (N_6489,N_4936,N_4575);
and U6490 (N_6490,N_4690,N_5263);
xnor U6491 (N_6491,N_5612,N_5103);
xnor U6492 (N_6492,N_5371,N_4774);
nor U6493 (N_6493,N_5554,N_4600);
xor U6494 (N_6494,N_5247,N_5520);
xnor U6495 (N_6495,N_5577,N_5016);
nand U6496 (N_6496,N_5883,N_4710);
nand U6497 (N_6497,N_5926,N_5125);
xnor U6498 (N_6498,N_5023,N_5508);
nand U6499 (N_6499,N_5152,N_4911);
xnor U6500 (N_6500,N_5505,N_5373);
nor U6501 (N_6501,N_5189,N_5565);
xnor U6502 (N_6502,N_5908,N_4798);
and U6503 (N_6503,N_5897,N_5051);
and U6504 (N_6504,N_5991,N_5486);
xor U6505 (N_6505,N_4939,N_5515);
nor U6506 (N_6506,N_5475,N_4676);
or U6507 (N_6507,N_4776,N_4599);
nand U6508 (N_6508,N_4534,N_5784);
or U6509 (N_6509,N_5343,N_4687);
nand U6510 (N_6510,N_4508,N_5853);
xor U6511 (N_6511,N_5282,N_4532);
or U6512 (N_6512,N_5803,N_5438);
nor U6513 (N_6513,N_4791,N_5876);
nor U6514 (N_6514,N_5423,N_5174);
nand U6515 (N_6515,N_4702,N_5012);
nor U6516 (N_6516,N_4833,N_5472);
or U6517 (N_6517,N_5882,N_5752);
xor U6518 (N_6518,N_5270,N_4752);
and U6519 (N_6519,N_5018,N_5600);
nor U6520 (N_6520,N_5671,N_5642);
and U6521 (N_6521,N_5294,N_5077);
and U6522 (N_6522,N_5191,N_5873);
nor U6523 (N_6523,N_5628,N_5927);
and U6524 (N_6524,N_4712,N_5817);
or U6525 (N_6525,N_4856,N_4635);
nor U6526 (N_6526,N_5605,N_4683);
or U6527 (N_6527,N_5814,N_5785);
nand U6528 (N_6528,N_4517,N_4664);
xnor U6529 (N_6529,N_4880,N_4590);
nand U6530 (N_6530,N_4618,N_4564);
nand U6531 (N_6531,N_5166,N_5518);
or U6532 (N_6532,N_5841,N_4893);
and U6533 (N_6533,N_5363,N_4747);
or U6534 (N_6534,N_5255,N_5226);
or U6535 (N_6535,N_5203,N_4504);
and U6536 (N_6536,N_5060,N_5562);
nand U6537 (N_6537,N_5446,N_5098);
and U6538 (N_6538,N_5079,N_5501);
xor U6539 (N_6539,N_4692,N_5978);
nand U6540 (N_6540,N_4571,N_5967);
nand U6541 (N_6541,N_5431,N_4714);
or U6542 (N_6542,N_5461,N_5241);
and U6543 (N_6543,N_5634,N_5649);
or U6544 (N_6544,N_5028,N_5512);
xnor U6545 (N_6545,N_5932,N_4634);
and U6546 (N_6546,N_4539,N_5417);
or U6547 (N_6547,N_5863,N_5193);
xnor U6548 (N_6548,N_4741,N_4629);
and U6549 (N_6549,N_4898,N_5490);
and U6550 (N_6550,N_4965,N_5783);
xor U6551 (N_6551,N_5111,N_5764);
nand U6552 (N_6552,N_4645,N_4820);
nand U6553 (N_6553,N_5620,N_5621);
nand U6554 (N_6554,N_5005,N_4520);
and U6555 (N_6555,N_5870,N_5744);
xor U6556 (N_6556,N_5564,N_5430);
and U6557 (N_6557,N_5640,N_5570);
nor U6558 (N_6558,N_5058,N_5192);
and U6559 (N_6559,N_4580,N_4932);
or U6560 (N_6560,N_5598,N_5272);
and U6561 (N_6561,N_4736,N_4967);
xor U6562 (N_6562,N_5267,N_5548);
and U6563 (N_6563,N_5302,N_5400);
or U6564 (N_6564,N_5857,N_5633);
or U6565 (N_6565,N_5832,N_4563);
and U6566 (N_6566,N_4746,N_5151);
xnor U6567 (N_6567,N_5895,N_5931);
and U6568 (N_6568,N_4626,N_5902);
and U6569 (N_6569,N_4677,N_5580);
or U6570 (N_6570,N_4950,N_5305);
xor U6571 (N_6571,N_5424,N_5530);
nor U6572 (N_6572,N_4729,N_5280);
xor U6573 (N_6573,N_4679,N_4938);
and U6574 (N_6574,N_5442,N_4900);
xnor U6575 (N_6575,N_4916,N_5831);
xnor U6576 (N_6576,N_5872,N_5607);
nand U6577 (N_6577,N_5650,N_4891);
nor U6578 (N_6578,N_5356,N_4807);
nor U6579 (N_6579,N_5253,N_5689);
xnor U6580 (N_6580,N_5389,N_4902);
nor U6581 (N_6581,N_4686,N_5033);
nor U6582 (N_6582,N_5232,N_4884);
and U6583 (N_6583,N_4627,N_5186);
nand U6584 (N_6584,N_5701,N_4526);
nand U6585 (N_6585,N_5278,N_5144);
or U6586 (N_6586,N_5124,N_4830);
xnor U6587 (N_6587,N_5452,N_4857);
nor U6588 (N_6588,N_4611,N_4780);
xor U6589 (N_6589,N_5426,N_5835);
nand U6590 (N_6590,N_5636,N_5603);
nor U6591 (N_6591,N_4572,N_4766);
or U6592 (N_6592,N_5854,N_4837);
nand U6593 (N_6593,N_4724,N_4772);
and U6594 (N_6594,N_5781,N_5436);
nand U6595 (N_6595,N_5643,N_4666);
xor U6596 (N_6596,N_5082,N_4809);
nand U6597 (N_6597,N_4904,N_5314);
nand U6598 (N_6598,N_5941,N_5147);
xor U6599 (N_6599,N_5763,N_4507);
nor U6600 (N_6600,N_5349,N_5031);
and U6601 (N_6601,N_5341,N_4529);
nand U6602 (N_6602,N_5674,N_5024);
xor U6603 (N_6603,N_5677,N_5422);
xnor U6604 (N_6604,N_4583,N_5691);
or U6605 (N_6605,N_5176,N_4862);
or U6606 (N_6606,N_5357,N_4553);
or U6607 (N_6607,N_5860,N_5974);
and U6608 (N_6608,N_5140,N_5298);
nand U6609 (N_6609,N_5419,N_5660);
nor U6610 (N_6610,N_4660,N_5625);
or U6611 (N_6611,N_5721,N_4802);
nor U6612 (N_6612,N_4983,N_4740);
nand U6613 (N_6613,N_5281,N_4726);
nor U6614 (N_6614,N_4673,N_5730);
or U6615 (N_6615,N_4886,N_5953);
or U6616 (N_6616,N_4797,N_5506);
and U6617 (N_6617,N_4765,N_5980);
nor U6618 (N_6618,N_5958,N_4552);
or U6619 (N_6619,N_5418,N_5561);
xor U6620 (N_6620,N_5896,N_5029);
and U6621 (N_6621,N_5710,N_4847);
or U6622 (N_6622,N_5483,N_4788);
nand U6623 (N_6623,N_5067,N_5318);
and U6624 (N_6624,N_4822,N_5425);
xnor U6625 (N_6625,N_4540,N_4775);
xor U6626 (N_6626,N_5366,N_5606);
xor U6627 (N_6627,N_5463,N_5480);
xnor U6628 (N_6628,N_4937,N_5020);
and U6629 (N_6629,N_4584,N_4933);
xnor U6630 (N_6630,N_5982,N_5722);
xnor U6631 (N_6631,N_5074,N_5647);
nand U6632 (N_6632,N_4568,N_5837);
or U6633 (N_6633,N_5139,N_5205);
nor U6634 (N_6634,N_5128,N_5584);
nor U6635 (N_6635,N_5627,N_5443);
and U6636 (N_6636,N_4556,N_5795);
and U6637 (N_6637,N_4718,N_5629);
or U6638 (N_6638,N_5055,N_5401);
nand U6639 (N_6639,N_4731,N_4907);
or U6640 (N_6640,N_5397,N_5126);
and U6641 (N_6641,N_5765,N_4734);
or U6642 (N_6642,N_4998,N_5588);
and U6643 (N_6643,N_5268,N_5891);
xnor U6644 (N_6644,N_5212,N_4767);
nand U6645 (N_6645,N_5262,N_4846);
nand U6646 (N_6646,N_4895,N_4574);
xnor U6647 (N_6647,N_5583,N_5112);
nand U6648 (N_6648,N_5888,N_5045);
nand U6649 (N_6649,N_5955,N_5507);
xor U6650 (N_6650,N_5118,N_5301);
and U6651 (N_6651,N_5037,N_5989);
xnor U6652 (N_6652,N_5096,N_5072);
or U6653 (N_6653,N_5983,N_5694);
nand U6654 (N_6654,N_5772,N_4909);
or U6655 (N_6655,N_5566,N_4768);
xnor U6656 (N_6656,N_5046,N_5449);
or U6657 (N_6657,N_5303,N_4943);
nor U6658 (N_6658,N_4764,N_5358);
or U6659 (N_6659,N_5868,N_5757);
and U6660 (N_6660,N_5718,N_5064);
nand U6661 (N_6661,N_5550,N_5789);
or U6662 (N_6662,N_5597,N_5228);
nand U6663 (N_6663,N_5994,N_5574);
xnor U6664 (N_6664,N_4750,N_5276);
and U6665 (N_6665,N_5207,N_5907);
and U6666 (N_6666,N_4784,N_4803);
and U6667 (N_6667,N_5386,N_4828);
nor U6668 (N_6668,N_5069,N_5317);
and U6669 (N_6669,N_5066,N_4501);
nand U6670 (N_6670,N_5052,N_5407);
nand U6671 (N_6671,N_4821,N_4598);
nor U6672 (N_6672,N_4749,N_4796);
and U6673 (N_6673,N_4648,N_5361);
xnor U6674 (N_6674,N_5672,N_5117);
xor U6675 (N_6675,N_5113,N_4826);
or U6676 (N_6676,N_5083,N_5014);
or U6677 (N_6677,N_5569,N_5546);
nor U6678 (N_6678,N_4795,N_4653);
and U6679 (N_6679,N_4603,N_4926);
nor U6680 (N_6680,N_5458,N_5290);
nand U6681 (N_6681,N_5155,N_5370);
xor U6682 (N_6682,N_4612,N_4799);
nor U6683 (N_6683,N_5959,N_4624);
xnor U6684 (N_6684,N_5042,N_4929);
or U6685 (N_6685,N_5944,N_5734);
xnor U6686 (N_6686,N_5131,N_5697);
nor U6687 (N_6687,N_5110,N_5823);
and U6688 (N_6688,N_5027,N_5773);
and U6689 (N_6689,N_5061,N_4865);
or U6690 (N_6690,N_5143,N_5617);
and U6691 (N_6691,N_5993,N_4941);
and U6692 (N_6692,N_5903,N_5568);
xnor U6693 (N_6693,N_5336,N_5836);
or U6694 (N_6694,N_5611,N_4901);
or U6695 (N_6695,N_5549,N_5459);
nor U6696 (N_6696,N_5678,N_5900);
nor U6697 (N_6697,N_5618,N_4591);
xor U6698 (N_6698,N_4819,N_5726);
nor U6699 (N_6699,N_5444,N_4975);
nand U6700 (N_6700,N_4637,N_5393);
nand U6701 (N_6701,N_5911,N_4841);
and U6702 (N_6702,N_5774,N_5687);
xor U6703 (N_6703,N_5514,N_4951);
nor U6704 (N_6704,N_5264,N_4663);
nand U6705 (N_6705,N_5146,N_5652);
and U6706 (N_6706,N_5234,N_5875);
nor U6707 (N_6707,N_5008,N_4759);
or U6708 (N_6708,N_5555,N_5864);
nand U6709 (N_6709,N_5965,N_4732);
nand U6710 (N_6710,N_5591,N_5304);
xor U6711 (N_6711,N_5224,N_4641);
or U6712 (N_6712,N_5910,N_5723);
or U6713 (N_6713,N_4689,N_5909);
nand U6714 (N_6714,N_5432,N_4934);
nand U6715 (N_6715,N_5544,N_5406);
or U6716 (N_6716,N_4728,N_4678);
or U6717 (N_6717,N_5743,N_5715);
and U6718 (N_6718,N_4717,N_5719);
nor U6719 (N_6719,N_5656,N_4638);
nand U6720 (N_6720,N_4968,N_5399);
and U6721 (N_6721,N_5538,N_5050);
nand U6722 (N_6722,N_4693,N_5716);
xor U6723 (N_6723,N_5852,N_5651);
or U6724 (N_6724,N_5839,N_5085);
and U6725 (N_6725,N_5172,N_5685);
or U6726 (N_6726,N_5415,N_5175);
xor U6727 (N_6727,N_5884,N_5062);
or U6728 (N_6728,N_5622,N_4986);
nor U6729 (N_6729,N_5542,N_5285);
or U6730 (N_6730,N_5412,N_5686);
or U6731 (N_6731,N_5850,N_5034);
and U6732 (N_6732,N_5639,N_5470);
nor U6733 (N_6733,N_5277,N_5751);
xor U6734 (N_6734,N_5199,N_5229);
and U6735 (N_6735,N_4705,N_5223);
xnor U6736 (N_6736,N_5943,N_5342);
and U6737 (N_6737,N_5755,N_5513);
nor U6738 (N_6738,N_5445,N_5962);
nor U6739 (N_6739,N_5563,N_5319);
and U6740 (N_6740,N_5310,N_4870);
or U6741 (N_6741,N_4832,N_4755);
and U6742 (N_6742,N_5063,N_4524);
nand U6743 (N_6743,N_5657,N_5092);
xnor U6744 (N_6744,N_5376,N_5815);
nand U6745 (N_6745,N_5334,N_5335);
nand U6746 (N_6746,N_4674,N_5477);
xor U6747 (N_6747,N_5527,N_5178);
or U6748 (N_6748,N_4800,N_4547);
nand U6749 (N_6749,N_5619,N_5592);
nor U6750 (N_6750,N_5123,N_5731);
and U6751 (N_6751,N_5745,N_5910);
xor U6752 (N_6752,N_5135,N_5171);
nand U6753 (N_6753,N_5781,N_5548);
and U6754 (N_6754,N_5626,N_4980);
or U6755 (N_6755,N_4821,N_5764);
and U6756 (N_6756,N_5794,N_5557);
nor U6757 (N_6757,N_4551,N_5535);
nor U6758 (N_6758,N_5978,N_5370);
xor U6759 (N_6759,N_5642,N_5296);
or U6760 (N_6760,N_5910,N_5621);
or U6761 (N_6761,N_5352,N_5092);
nor U6762 (N_6762,N_5838,N_5149);
and U6763 (N_6763,N_5695,N_5663);
or U6764 (N_6764,N_5770,N_4854);
and U6765 (N_6765,N_5568,N_4522);
and U6766 (N_6766,N_5612,N_4933);
xnor U6767 (N_6767,N_5566,N_5800);
or U6768 (N_6768,N_5909,N_5152);
or U6769 (N_6769,N_4709,N_4558);
and U6770 (N_6770,N_5377,N_5754);
and U6771 (N_6771,N_5555,N_4610);
or U6772 (N_6772,N_4960,N_5826);
nor U6773 (N_6773,N_5992,N_5141);
nand U6774 (N_6774,N_5253,N_4887);
nand U6775 (N_6775,N_4723,N_4778);
and U6776 (N_6776,N_5828,N_5743);
nor U6777 (N_6777,N_5275,N_5694);
xnor U6778 (N_6778,N_5999,N_4806);
or U6779 (N_6779,N_5952,N_4915);
and U6780 (N_6780,N_5825,N_4859);
nor U6781 (N_6781,N_5351,N_5813);
xor U6782 (N_6782,N_5894,N_4892);
nand U6783 (N_6783,N_5612,N_5458);
xnor U6784 (N_6784,N_5205,N_5610);
or U6785 (N_6785,N_5097,N_5294);
and U6786 (N_6786,N_4734,N_4839);
xnor U6787 (N_6787,N_5960,N_4541);
or U6788 (N_6788,N_5766,N_4728);
nand U6789 (N_6789,N_4715,N_5214);
xnor U6790 (N_6790,N_5429,N_5190);
xor U6791 (N_6791,N_5612,N_4739);
or U6792 (N_6792,N_5261,N_4944);
or U6793 (N_6793,N_5222,N_5822);
nor U6794 (N_6794,N_5610,N_5824);
nand U6795 (N_6795,N_4607,N_5823);
xor U6796 (N_6796,N_5509,N_5448);
or U6797 (N_6797,N_5850,N_4787);
nand U6798 (N_6798,N_5023,N_5467);
nor U6799 (N_6799,N_5097,N_4993);
or U6800 (N_6800,N_5837,N_5659);
or U6801 (N_6801,N_5892,N_5573);
and U6802 (N_6802,N_5313,N_5871);
xor U6803 (N_6803,N_5137,N_5918);
and U6804 (N_6804,N_5219,N_5041);
nand U6805 (N_6805,N_4822,N_4769);
xor U6806 (N_6806,N_4501,N_5211);
and U6807 (N_6807,N_5310,N_5854);
nor U6808 (N_6808,N_5025,N_5377);
nand U6809 (N_6809,N_5088,N_4778);
nand U6810 (N_6810,N_4825,N_5647);
xor U6811 (N_6811,N_5014,N_5375);
or U6812 (N_6812,N_5435,N_4539);
xor U6813 (N_6813,N_5213,N_5415);
and U6814 (N_6814,N_4843,N_4858);
or U6815 (N_6815,N_5579,N_4694);
xor U6816 (N_6816,N_5393,N_5070);
xnor U6817 (N_6817,N_4520,N_5978);
xnor U6818 (N_6818,N_4822,N_5327);
and U6819 (N_6819,N_4658,N_4807);
nand U6820 (N_6820,N_5638,N_4824);
and U6821 (N_6821,N_5550,N_4670);
nand U6822 (N_6822,N_5346,N_5605);
nand U6823 (N_6823,N_4824,N_5415);
or U6824 (N_6824,N_4814,N_5726);
nand U6825 (N_6825,N_4568,N_5096);
xor U6826 (N_6826,N_4761,N_4946);
xor U6827 (N_6827,N_5284,N_5301);
nand U6828 (N_6828,N_5428,N_5139);
xnor U6829 (N_6829,N_4506,N_5773);
nor U6830 (N_6830,N_4724,N_4615);
nand U6831 (N_6831,N_4693,N_5681);
and U6832 (N_6832,N_5192,N_5320);
or U6833 (N_6833,N_4786,N_5361);
nand U6834 (N_6834,N_5388,N_5940);
nand U6835 (N_6835,N_5536,N_5075);
nor U6836 (N_6836,N_5689,N_5935);
and U6837 (N_6837,N_5764,N_4958);
or U6838 (N_6838,N_5359,N_5959);
nand U6839 (N_6839,N_5547,N_4549);
and U6840 (N_6840,N_4898,N_5860);
or U6841 (N_6841,N_5587,N_4529);
or U6842 (N_6842,N_5832,N_5586);
or U6843 (N_6843,N_5480,N_4561);
nand U6844 (N_6844,N_5495,N_5960);
nand U6845 (N_6845,N_4640,N_4792);
nand U6846 (N_6846,N_5398,N_5285);
or U6847 (N_6847,N_5036,N_5615);
nand U6848 (N_6848,N_5020,N_5077);
or U6849 (N_6849,N_4844,N_5725);
or U6850 (N_6850,N_5954,N_5966);
or U6851 (N_6851,N_5162,N_5974);
or U6852 (N_6852,N_5758,N_4756);
nand U6853 (N_6853,N_4872,N_4825);
nand U6854 (N_6854,N_4971,N_5937);
and U6855 (N_6855,N_4715,N_4914);
xnor U6856 (N_6856,N_5795,N_5433);
nand U6857 (N_6857,N_5983,N_5890);
and U6858 (N_6858,N_5245,N_5080);
nor U6859 (N_6859,N_5293,N_4906);
and U6860 (N_6860,N_5105,N_5359);
xnor U6861 (N_6861,N_5279,N_5631);
nor U6862 (N_6862,N_4780,N_4514);
nand U6863 (N_6863,N_5306,N_4623);
xnor U6864 (N_6864,N_4640,N_5344);
or U6865 (N_6865,N_4816,N_5526);
nor U6866 (N_6866,N_5082,N_4511);
or U6867 (N_6867,N_5595,N_5900);
nor U6868 (N_6868,N_5215,N_4640);
xor U6869 (N_6869,N_5416,N_5774);
and U6870 (N_6870,N_5153,N_5511);
nand U6871 (N_6871,N_5439,N_5909);
xor U6872 (N_6872,N_4662,N_4754);
xnor U6873 (N_6873,N_5519,N_5895);
or U6874 (N_6874,N_4689,N_5152);
or U6875 (N_6875,N_4832,N_4775);
nor U6876 (N_6876,N_4702,N_5068);
and U6877 (N_6877,N_4958,N_5469);
xor U6878 (N_6878,N_5123,N_4944);
or U6879 (N_6879,N_5185,N_4728);
and U6880 (N_6880,N_4956,N_5899);
nor U6881 (N_6881,N_5688,N_4991);
and U6882 (N_6882,N_5945,N_5895);
xor U6883 (N_6883,N_5350,N_4946);
xnor U6884 (N_6884,N_4508,N_4657);
or U6885 (N_6885,N_5287,N_5421);
nand U6886 (N_6886,N_5151,N_5031);
and U6887 (N_6887,N_4584,N_4683);
nor U6888 (N_6888,N_4595,N_4530);
nor U6889 (N_6889,N_5356,N_4504);
nor U6890 (N_6890,N_4929,N_4979);
nor U6891 (N_6891,N_5756,N_5206);
nand U6892 (N_6892,N_5568,N_4666);
xnor U6893 (N_6893,N_5687,N_4810);
xor U6894 (N_6894,N_5459,N_5002);
and U6895 (N_6895,N_5347,N_4572);
nand U6896 (N_6896,N_5366,N_4526);
and U6897 (N_6897,N_5970,N_5716);
nand U6898 (N_6898,N_5241,N_5994);
and U6899 (N_6899,N_5275,N_5681);
and U6900 (N_6900,N_5409,N_5922);
or U6901 (N_6901,N_5542,N_5517);
nor U6902 (N_6902,N_5203,N_4846);
or U6903 (N_6903,N_5284,N_4946);
xor U6904 (N_6904,N_5229,N_4956);
nand U6905 (N_6905,N_5365,N_5806);
or U6906 (N_6906,N_5485,N_5285);
xnor U6907 (N_6907,N_4566,N_5414);
nor U6908 (N_6908,N_4915,N_5190);
or U6909 (N_6909,N_5049,N_5640);
and U6910 (N_6910,N_4686,N_5071);
nand U6911 (N_6911,N_5440,N_4738);
nor U6912 (N_6912,N_5096,N_4519);
xor U6913 (N_6913,N_5657,N_4851);
and U6914 (N_6914,N_4542,N_4755);
nand U6915 (N_6915,N_5888,N_5784);
xnor U6916 (N_6916,N_5837,N_5101);
xor U6917 (N_6917,N_5270,N_5159);
xor U6918 (N_6918,N_4985,N_5854);
xor U6919 (N_6919,N_4916,N_4913);
nand U6920 (N_6920,N_5792,N_4792);
xnor U6921 (N_6921,N_5964,N_5832);
nor U6922 (N_6922,N_4805,N_5293);
xnor U6923 (N_6923,N_4830,N_5256);
and U6924 (N_6924,N_4724,N_5057);
xnor U6925 (N_6925,N_5773,N_4704);
xor U6926 (N_6926,N_5476,N_5739);
nand U6927 (N_6927,N_5770,N_4613);
nor U6928 (N_6928,N_4733,N_5077);
or U6929 (N_6929,N_4898,N_5520);
and U6930 (N_6930,N_5512,N_4523);
nor U6931 (N_6931,N_4966,N_4944);
xnor U6932 (N_6932,N_4989,N_4914);
or U6933 (N_6933,N_5895,N_5942);
and U6934 (N_6934,N_5903,N_4608);
and U6935 (N_6935,N_4857,N_5831);
xor U6936 (N_6936,N_4719,N_4989);
and U6937 (N_6937,N_5248,N_5346);
and U6938 (N_6938,N_5816,N_5437);
and U6939 (N_6939,N_4579,N_5599);
nand U6940 (N_6940,N_5659,N_4894);
xnor U6941 (N_6941,N_4591,N_4939);
or U6942 (N_6942,N_5929,N_4535);
xor U6943 (N_6943,N_4845,N_5471);
xnor U6944 (N_6944,N_5016,N_5427);
nor U6945 (N_6945,N_5932,N_5354);
nor U6946 (N_6946,N_5100,N_4643);
xnor U6947 (N_6947,N_5350,N_5277);
or U6948 (N_6948,N_5819,N_5880);
xnor U6949 (N_6949,N_5336,N_4927);
nor U6950 (N_6950,N_4540,N_5570);
and U6951 (N_6951,N_4544,N_5286);
or U6952 (N_6952,N_5173,N_4722);
or U6953 (N_6953,N_5075,N_5513);
nand U6954 (N_6954,N_5875,N_5501);
xor U6955 (N_6955,N_5634,N_5358);
xor U6956 (N_6956,N_5458,N_4720);
and U6957 (N_6957,N_5204,N_5310);
nor U6958 (N_6958,N_5373,N_5310);
xnor U6959 (N_6959,N_4611,N_5402);
or U6960 (N_6960,N_5976,N_4567);
and U6961 (N_6961,N_5729,N_5696);
nand U6962 (N_6962,N_5666,N_5315);
nand U6963 (N_6963,N_4711,N_5485);
nor U6964 (N_6964,N_5680,N_5944);
and U6965 (N_6965,N_5443,N_5196);
xor U6966 (N_6966,N_5153,N_5971);
nand U6967 (N_6967,N_5006,N_5360);
nor U6968 (N_6968,N_5623,N_4643);
xnor U6969 (N_6969,N_5885,N_5206);
nor U6970 (N_6970,N_4579,N_5444);
or U6971 (N_6971,N_5809,N_4648);
xnor U6972 (N_6972,N_5959,N_5551);
or U6973 (N_6973,N_5055,N_5067);
or U6974 (N_6974,N_5429,N_5828);
and U6975 (N_6975,N_4797,N_5050);
xnor U6976 (N_6976,N_4528,N_4598);
nand U6977 (N_6977,N_5381,N_4793);
nor U6978 (N_6978,N_4816,N_5540);
or U6979 (N_6979,N_5965,N_4887);
nand U6980 (N_6980,N_5415,N_5044);
nor U6981 (N_6981,N_5617,N_5790);
nor U6982 (N_6982,N_4981,N_5276);
or U6983 (N_6983,N_5756,N_5003);
xor U6984 (N_6984,N_5784,N_5892);
nor U6985 (N_6985,N_5471,N_4679);
nand U6986 (N_6986,N_5944,N_4725);
or U6987 (N_6987,N_4598,N_5115);
nor U6988 (N_6988,N_5831,N_4718);
and U6989 (N_6989,N_4666,N_4869);
nor U6990 (N_6990,N_5745,N_4766);
nand U6991 (N_6991,N_4644,N_5235);
or U6992 (N_6992,N_4800,N_5890);
xor U6993 (N_6993,N_5123,N_5935);
and U6994 (N_6994,N_4840,N_5833);
or U6995 (N_6995,N_4833,N_4926);
and U6996 (N_6996,N_5525,N_4869);
nand U6997 (N_6997,N_5540,N_5901);
or U6998 (N_6998,N_4790,N_5150);
nor U6999 (N_6999,N_5312,N_5071);
xnor U7000 (N_7000,N_5269,N_5693);
nand U7001 (N_7001,N_4857,N_4674);
xnor U7002 (N_7002,N_5397,N_5437);
or U7003 (N_7003,N_4661,N_5719);
xnor U7004 (N_7004,N_5764,N_4864);
nand U7005 (N_7005,N_5676,N_4715);
xor U7006 (N_7006,N_4603,N_4743);
nor U7007 (N_7007,N_5061,N_4591);
or U7008 (N_7008,N_5184,N_4577);
nand U7009 (N_7009,N_5441,N_5006);
xor U7010 (N_7010,N_5235,N_5323);
nand U7011 (N_7011,N_5413,N_5401);
nor U7012 (N_7012,N_4881,N_5029);
nand U7013 (N_7013,N_5754,N_5511);
and U7014 (N_7014,N_4724,N_5015);
or U7015 (N_7015,N_5149,N_5842);
xor U7016 (N_7016,N_5198,N_4506);
nor U7017 (N_7017,N_5124,N_4747);
xnor U7018 (N_7018,N_4920,N_4714);
nor U7019 (N_7019,N_5951,N_5674);
or U7020 (N_7020,N_5919,N_4868);
xnor U7021 (N_7021,N_4636,N_5857);
xnor U7022 (N_7022,N_4764,N_5278);
nor U7023 (N_7023,N_5295,N_4654);
xnor U7024 (N_7024,N_5418,N_5153);
and U7025 (N_7025,N_5430,N_4774);
nand U7026 (N_7026,N_5912,N_4914);
nand U7027 (N_7027,N_5356,N_4763);
nand U7028 (N_7028,N_5770,N_5781);
nor U7029 (N_7029,N_4845,N_5960);
nand U7030 (N_7030,N_5534,N_5124);
nor U7031 (N_7031,N_5663,N_4820);
and U7032 (N_7032,N_4996,N_5161);
or U7033 (N_7033,N_5193,N_5384);
and U7034 (N_7034,N_4983,N_5763);
xor U7035 (N_7035,N_4659,N_5736);
or U7036 (N_7036,N_4788,N_5086);
nor U7037 (N_7037,N_5532,N_5790);
nand U7038 (N_7038,N_4573,N_4587);
and U7039 (N_7039,N_5408,N_4670);
or U7040 (N_7040,N_4544,N_4965);
nand U7041 (N_7041,N_5321,N_5803);
or U7042 (N_7042,N_5202,N_4877);
and U7043 (N_7043,N_5815,N_5614);
nor U7044 (N_7044,N_5322,N_4955);
and U7045 (N_7045,N_5556,N_4742);
nand U7046 (N_7046,N_5872,N_4656);
and U7047 (N_7047,N_5140,N_4785);
nor U7048 (N_7048,N_4863,N_4538);
nand U7049 (N_7049,N_4943,N_5801);
nand U7050 (N_7050,N_4703,N_5936);
nand U7051 (N_7051,N_5632,N_5884);
and U7052 (N_7052,N_4879,N_4920);
nand U7053 (N_7053,N_4687,N_4616);
and U7054 (N_7054,N_5280,N_4579);
nand U7055 (N_7055,N_4640,N_5362);
and U7056 (N_7056,N_5382,N_4679);
nor U7057 (N_7057,N_5877,N_5664);
and U7058 (N_7058,N_5904,N_5124);
or U7059 (N_7059,N_5655,N_5422);
xor U7060 (N_7060,N_5582,N_4924);
and U7061 (N_7061,N_5961,N_4910);
or U7062 (N_7062,N_5669,N_4655);
nor U7063 (N_7063,N_5596,N_5929);
nand U7064 (N_7064,N_4759,N_5575);
or U7065 (N_7065,N_5216,N_5702);
xor U7066 (N_7066,N_5746,N_5052);
nor U7067 (N_7067,N_5361,N_4610);
or U7068 (N_7068,N_5033,N_4895);
and U7069 (N_7069,N_5787,N_5621);
and U7070 (N_7070,N_5483,N_5627);
nand U7071 (N_7071,N_5772,N_4707);
and U7072 (N_7072,N_5941,N_4858);
or U7073 (N_7073,N_5064,N_5131);
or U7074 (N_7074,N_4941,N_4636);
nand U7075 (N_7075,N_5970,N_5249);
and U7076 (N_7076,N_5876,N_5460);
nand U7077 (N_7077,N_4856,N_5641);
nand U7078 (N_7078,N_4876,N_5883);
or U7079 (N_7079,N_4706,N_5138);
xnor U7080 (N_7080,N_5042,N_4678);
nor U7081 (N_7081,N_5166,N_5515);
and U7082 (N_7082,N_4549,N_4994);
nand U7083 (N_7083,N_4517,N_5485);
or U7084 (N_7084,N_4876,N_4979);
xor U7085 (N_7085,N_4561,N_5840);
nor U7086 (N_7086,N_5992,N_4651);
xor U7087 (N_7087,N_5789,N_5037);
nor U7088 (N_7088,N_5522,N_5751);
or U7089 (N_7089,N_5219,N_5947);
or U7090 (N_7090,N_5893,N_4521);
or U7091 (N_7091,N_5201,N_5987);
xnor U7092 (N_7092,N_5551,N_4703);
and U7093 (N_7093,N_4817,N_5645);
nor U7094 (N_7094,N_5436,N_5027);
nor U7095 (N_7095,N_5961,N_4954);
nand U7096 (N_7096,N_5786,N_4762);
or U7097 (N_7097,N_5656,N_5842);
or U7098 (N_7098,N_5981,N_5365);
nand U7099 (N_7099,N_4911,N_5644);
or U7100 (N_7100,N_4854,N_5565);
nand U7101 (N_7101,N_4653,N_4836);
xnor U7102 (N_7102,N_5758,N_4989);
nor U7103 (N_7103,N_5067,N_5627);
xor U7104 (N_7104,N_4515,N_5756);
nand U7105 (N_7105,N_5998,N_4972);
nand U7106 (N_7106,N_4502,N_4989);
or U7107 (N_7107,N_5798,N_5382);
and U7108 (N_7108,N_5008,N_5890);
nand U7109 (N_7109,N_4846,N_4606);
nor U7110 (N_7110,N_4606,N_5161);
nand U7111 (N_7111,N_5005,N_4751);
and U7112 (N_7112,N_5888,N_5669);
nor U7113 (N_7113,N_4550,N_5029);
or U7114 (N_7114,N_5757,N_5247);
or U7115 (N_7115,N_4717,N_5058);
nand U7116 (N_7116,N_5886,N_4818);
nor U7117 (N_7117,N_4682,N_5512);
and U7118 (N_7118,N_5564,N_5831);
nor U7119 (N_7119,N_5391,N_4905);
or U7120 (N_7120,N_5990,N_5042);
or U7121 (N_7121,N_4530,N_4834);
and U7122 (N_7122,N_4765,N_5630);
xnor U7123 (N_7123,N_4608,N_5418);
or U7124 (N_7124,N_4924,N_5010);
and U7125 (N_7125,N_5948,N_4848);
nor U7126 (N_7126,N_5786,N_5919);
xor U7127 (N_7127,N_4637,N_4731);
nor U7128 (N_7128,N_4599,N_4924);
nor U7129 (N_7129,N_4552,N_4525);
xnor U7130 (N_7130,N_5818,N_4879);
or U7131 (N_7131,N_5257,N_5340);
nand U7132 (N_7132,N_5938,N_4867);
or U7133 (N_7133,N_5521,N_5244);
nand U7134 (N_7134,N_5400,N_5683);
or U7135 (N_7135,N_5844,N_5448);
and U7136 (N_7136,N_5371,N_4760);
nand U7137 (N_7137,N_5058,N_4697);
xnor U7138 (N_7138,N_4543,N_5064);
xor U7139 (N_7139,N_5459,N_5347);
xnor U7140 (N_7140,N_5175,N_5076);
or U7141 (N_7141,N_4914,N_5528);
and U7142 (N_7142,N_5743,N_5806);
nor U7143 (N_7143,N_4751,N_5742);
nor U7144 (N_7144,N_4990,N_5591);
xor U7145 (N_7145,N_5699,N_5865);
or U7146 (N_7146,N_5648,N_5653);
xnor U7147 (N_7147,N_4659,N_4652);
or U7148 (N_7148,N_4671,N_5975);
nor U7149 (N_7149,N_5634,N_4769);
xor U7150 (N_7150,N_5739,N_5778);
or U7151 (N_7151,N_4743,N_5922);
nand U7152 (N_7152,N_5430,N_4642);
and U7153 (N_7153,N_4791,N_4614);
nor U7154 (N_7154,N_5619,N_5444);
and U7155 (N_7155,N_5977,N_5254);
and U7156 (N_7156,N_5841,N_5133);
nand U7157 (N_7157,N_5954,N_5122);
xnor U7158 (N_7158,N_5787,N_5976);
and U7159 (N_7159,N_5960,N_4515);
xnor U7160 (N_7160,N_5220,N_4623);
xnor U7161 (N_7161,N_5837,N_5572);
nor U7162 (N_7162,N_5047,N_4863);
nor U7163 (N_7163,N_5219,N_4590);
nand U7164 (N_7164,N_5807,N_5913);
nor U7165 (N_7165,N_5973,N_5328);
and U7166 (N_7166,N_5671,N_5152);
xor U7167 (N_7167,N_5560,N_4966);
xnor U7168 (N_7168,N_4792,N_4820);
nor U7169 (N_7169,N_5702,N_5763);
nor U7170 (N_7170,N_5829,N_4732);
nand U7171 (N_7171,N_5026,N_5441);
or U7172 (N_7172,N_5408,N_5603);
or U7173 (N_7173,N_5325,N_4987);
nor U7174 (N_7174,N_5163,N_4995);
xor U7175 (N_7175,N_4782,N_5765);
xnor U7176 (N_7176,N_4787,N_5705);
xor U7177 (N_7177,N_5579,N_5050);
nor U7178 (N_7178,N_4919,N_4856);
and U7179 (N_7179,N_4904,N_4581);
nor U7180 (N_7180,N_4679,N_5840);
xor U7181 (N_7181,N_5675,N_5622);
nand U7182 (N_7182,N_4626,N_5113);
xnor U7183 (N_7183,N_5624,N_5670);
and U7184 (N_7184,N_5297,N_4618);
and U7185 (N_7185,N_5652,N_5412);
nand U7186 (N_7186,N_4843,N_5729);
or U7187 (N_7187,N_5818,N_4854);
nand U7188 (N_7188,N_4971,N_4901);
or U7189 (N_7189,N_5277,N_5412);
nor U7190 (N_7190,N_4658,N_5430);
and U7191 (N_7191,N_4544,N_5105);
nor U7192 (N_7192,N_5239,N_4672);
or U7193 (N_7193,N_4773,N_4993);
nor U7194 (N_7194,N_5677,N_5563);
xnor U7195 (N_7195,N_5389,N_4984);
nand U7196 (N_7196,N_5781,N_5939);
nand U7197 (N_7197,N_4673,N_4534);
nor U7198 (N_7198,N_4934,N_4887);
and U7199 (N_7199,N_5118,N_4889);
nor U7200 (N_7200,N_5652,N_5382);
nand U7201 (N_7201,N_5943,N_5222);
or U7202 (N_7202,N_5146,N_5383);
nand U7203 (N_7203,N_5469,N_5584);
or U7204 (N_7204,N_4503,N_4673);
nor U7205 (N_7205,N_5930,N_5517);
or U7206 (N_7206,N_5203,N_5719);
or U7207 (N_7207,N_5204,N_5552);
and U7208 (N_7208,N_5078,N_4771);
nand U7209 (N_7209,N_5507,N_5247);
or U7210 (N_7210,N_5688,N_4703);
or U7211 (N_7211,N_5300,N_5773);
xor U7212 (N_7212,N_5283,N_4661);
nand U7213 (N_7213,N_5710,N_5456);
nor U7214 (N_7214,N_4836,N_5740);
or U7215 (N_7215,N_4593,N_5559);
nor U7216 (N_7216,N_5256,N_5919);
nand U7217 (N_7217,N_5195,N_4679);
nand U7218 (N_7218,N_5548,N_5519);
xnor U7219 (N_7219,N_5715,N_5498);
nand U7220 (N_7220,N_5618,N_5798);
nand U7221 (N_7221,N_4509,N_4948);
or U7222 (N_7222,N_5595,N_5386);
nand U7223 (N_7223,N_5276,N_4550);
nand U7224 (N_7224,N_4514,N_5642);
nor U7225 (N_7225,N_5970,N_5812);
or U7226 (N_7226,N_4665,N_5606);
nor U7227 (N_7227,N_5869,N_5707);
nor U7228 (N_7228,N_5292,N_5156);
xnor U7229 (N_7229,N_5341,N_5716);
xor U7230 (N_7230,N_5671,N_4958);
xor U7231 (N_7231,N_4528,N_4676);
and U7232 (N_7232,N_5624,N_5044);
xor U7233 (N_7233,N_5176,N_5233);
nor U7234 (N_7234,N_4806,N_5452);
or U7235 (N_7235,N_4658,N_4619);
or U7236 (N_7236,N_5146,N_5668);
nand U7237 (N_7237,N_5864,N_5700);
nand U7238 (N_7238,N_4502,N_5527);
xor U7239 (N_7239,N_4672,N_5936);
nor U7240 (N_7240,N_5043,N_5653);
xor U7241 (N_7241,N_5624,N_4995);
nor U7242 (N_7242,N_5393,N_5006);
xnor U7243 (N_7243,N_4625,N_5462);
xor U7244 (N_7244,N_5339,N_4691);
nor U7245 (N_7245,N_4899,N_5982);
nand U7246 (N_7246,N_5517,N_5787);
or U7247 (N_7247,N_5156,N_5273);
and U7248 (N_7248,N_5874,N_4592);
and U7249 (N_7249,N_5579,N_5392);
xnor U7250 (N_7250,N_5855,N_5643);
xor U7251 (N_7251,N_5528,N_5502);
and U7252 (N_7252,N_4923,N_5174);
xor U7253 (N_7253,N_5856,N_5270);
or U7254 (N_7254,N_5613,N_4602);
nand U7255 (N_7255,N_4501,N_5157);
xnor U7256 (N_7256,N_5669,N_4908);
nor U7257 (N_7257,N_5284,N_5072);
nand U7258 (N_7258,N_5266,N_5656);
and U7259 (N_7259,N_5339,N_5414);
nand U7260 (N_7260,N_4980,N_4678);
or U7261 (N_7261,N_4925,N_4876);
or U7262 (N_7262,N_4977,N_5382);
nor U7263 (N_7263,N_5398,N_4711);
and U7264 (N_7264,N_5852,N_4665);
nor U7265 (N_7265,N_5049,N_5421);
nand U7266 (N_7266,N_5512,N_4620);
and U7267 (N_7267,N_4955,N_5865);
nor U7268 (N_7268,N_4859,N_5878);
xnor U7269 (N_7269,N_5590,N_5246);
xnor U7270 (N_7270,N_5951,N_4638);
and U7271 (N_7271,N_4819,N_4710);
and U7272 (N_7272,N_5884,N_5938);
nor U7273 (N_7273,N_5124,N_5354);
nand U7274 (N_7274,N_5712,N_4762);
nand U7275 (N_7275,N_4702,N_4621);
or U7276 (N_7276,N_5158,N_5644);
nand U7277 (N_7277,N_4922,N_5796);
or U7278 (N_7278,N_5970,N_5631);
or U7279 (N_7279,N_4966,N_5380);
or U7280 (N_7280,N_5779,N_5373);
nand U7281 (N_7281,N_5661,N_5674);
or U7282 (N_7282,N_4972,N_5159);
nand U7283 (N_7283,N_5458,N_5946);
or U7284 (N_7284,N_5013,N_5980);
xor U7285 (N_7285,N_5888,N_5731);
nand U7286 (N_7286,N_5380,N_5516);
xnor U7287 (N_7287,N_4807,N_4599);
nor U7288 (N_7288,N_4671,N_4822);
nand U7289 (N_7289,N_5652,N_5938);
xor U7290 (N_7290,N_4764,N_5265);
or U7291 (N_7291,N_5016,N_5314);
nor U7292 (N_7292,N_5755,N_4599);
xor U7293 (N_7293,N_4779,N_5356);
nand U7294 (N_7294,N_4678,N_4956);
and U7295 (N_7295,N_4893,N_4632);
nand U7296 (N_7296,N_5794,N_4959);
and U7297 (N_7297,N_4515,N_5605);
nor U7298 (N_7298,N_5690,N_4918);
nand U7299 (N_7299,N_5884,N_5542);
xor U7300 (N_7300,N_5910,N_5311);
nand U7301 (N_7301,N_5294,N_5407);
or U7302 (N_7302,N_5489,N_4733);
nand U7303 (N_7303,N_4541,N_5617);
or U7304 (N_7304,N_5038,N_4732);
or U7305 (N_7305,N_5175,N_5836);
xnor U7306 (N_7306,N_4850,N_5543);
and U7307 (N_7307,N_5753,N_4755);
xnor U7308 (N_7308,N_5048,N_5509);
nor U7309 (N_7309,N_5475,N_4818);
and U7310 (N_7310,N_5055,N_4891);
and U7311 (N_7311,N_5317,N_5086);
xnor U7312 (N_7312,N_5789,N_5475);
nand U7313 (N_7313,N_4945,N_5596);
or U7314 (N_7314,N_5896,N_5440);
nand U7315 (N_7315,N_5152,N_5940);
and U7316 (N_7316,N_5877,N_5694);
nand U7317 (N_7317,N_5460,N_5913);
nand U7318 (N_7318,N_5329,N_5667);
or U7319 (N_7319,N_4811,N_4749);
or U7320 (N_7320,N_5221,N_4941);
or U7321 (N_7321,N_4932,N_5599);
and U7322 (N_7322,N_5835,N_5586);
and U7323 (N_7323,N_4528,N_5220);
and U7324 (N_7324,N_4895,N_5678);
and U7325 (N_7325,N_4930,N_4588);
xor U7326 (N_7326,N_5737,N_5532);
or U7327 (N_7327,N_5322,N_4741);
nor U7328 (N_7328,N_5548,N_5348);
or U7329 (N_7329,N_5219,N_5310);
nor U7330 (N_7330,N_5145,N_5197);
and U7331 (N_7331,N_4931,N_5907);
nor U7332 (N_7332,N_4507,N_5488);
or U7333 (N_7333,N_5865,N_4913);
and U7334 (N_7334,N_5559,N_5849);
and U7335 (N_7335,N_4702,N_5894);
nand U7336 (N_7336,N_5277,N_5181);
nor U7337 (N_7337,N_5994,N_4741);
nand U7338 (N_7338,N_5539,N_5910);
or U7339 (N_7339,N_4560,N_5199);
nand U7340 (N_7340,N_5291,N_4816);
xor U7341 (N_7341,N_4611,N_5598);
xor U7342 (N_7342,N_5725,N_4672);
or U7343 (N_7343,N_5729,N_4544);
or U7344 (N_7344,N_4543,N_5675);
nor U7345 (N_7345,N_5133,N_5495);
xnor U7346 (N_7346,N_5078,N_4513);
or U7347 (N_7347,N_5066,N_4746);
and U7348 (N_7348,N_4510,N_5656);
nand U7349 (N_7349,N_5987,N_4595);
nor U7350 (N_7350,N_4953,N_5117);
xnor U7351 (N_7351,N_4619,N_5057);
nand U7352 (N_7352,N_5123,N_5312);
or U7353 (N_7353,N_5198,N_5231);
nand U7354 (N_7354,N_5021,N_4795);
xnor U7355 (N_7355,N_4960,N_4552);
xor U7356 (N_7356,N_4591,N_5763);
nand U7357 (N_7357,N_4928,N_5450);
nand U7358 (N_7358,N_4955,N_5047);
nor U7359 (N_7359,N_5891,N_4703);
or U7360 (N_7360,N_5250,N_4816);
nor U7361 (N_7361,N_4699,N_5357);
or U7362 (N_7362,N_4719,N_5753);
nor U7363 (N_7363,N_5604,N_5389);
and U7364 (N_7364,N_5259,N_5225);
nand U7365 (N_7365,N_5764,N_5828);
nand U7366 (N_7366,N_5353,N_5557);
and U7367 (N_7367,N_5590,N_4684);
nand U7368 (N_7368,N_5168,N_5248);
xor U7369 (N_7369,N_5989,N_4902);
nand U7370 (N_7370,N_5785,N_4540);
nand U7371 (N_7371,N_5634,N_4889);
xor U7372 (N_7372,N_5389,N_5275);
xor U7373 (N_7373,N_5582,N_5718);
nor U7374 (N_7374,N_4893,N_5047);
xnor U7375 (N_7375,N_5443,N_5087);
xnor U7376 (N_7376,N_5210,N_4605);
xor U7377 (N_7377,N_5579,N_4627);
or U7378 (N_7378,N_5105,N_4665);
and U7379 (N_7379,N_4852,N_4670);
nand U7380 (N_7380,N_5703,N_5607);
and U7381 (N_7381,N_5986,N_5173);
nor U7382 (N_7382,N_5481,N_5835);
xor U7383 (N_7383,N_5525,N_4601);
nand U7384 (N_7384,N_4610,N_4730);
and U7385 (N_7385,N_5019,N_5433);
or U7386 (N_7386,N_5831,N_5945);
xor U7387 (N_7387,N_5680,N_4657);
and U7388 (N_7388,N_4676,N_5568);
and U7389 (N_7389,N_4733,N_4866);
and U7390 (N_7390,N_5612,N_4600);
nand U7391 (N_7391,N_4553,N_5450);
nand U7392 (N_7392,N_4802,N_4827);
nor U7393 (N_7393,N_5908,N_5126);
xnor U7394 (N_7394,N_5547,N_5113);
nor U7395 (N_7395,N_4612,N_4571);
xor U7396 (N_7396,N_5302,N_4634);
or U7397 (N_7397,N_5107,N_5341);
xor U7398 (N_7398,N_5448,N_5507);
or U7399 (N_7399,N_5466,N_5518);
or U7400 (N_7400,N_5907,N_5340);
xor U7401 (N_7401,N_5715,N_5352);
nand U7402 (N_7402,N_4777,N_5692);
and U7403 (N_7403,N_5335,N_5064);
nor U7404 (N_7404,N_4886,N_4890);
or U7405 (N_7405,N_5176,N_5748);
and U7406 (N_7406,N_5740,N_5673);
nor U7407 (N_7407,N_4663,N_4778);
nor U7408 (N_7408,N_5499,N_5227);
and U7409 (N_7409,N_5408,N_5727);
xnor U7410 (N_7410,N_5502,N_5388);
nand U7411 (N_7411,N_5333,N_5054);
xnor U7412 (N_7412,N_4885,N_5200);
and U7413 (N_7413,N_5101,N_5716);
or U7414 (N_7414,N_5774,N_4647);
xor U7415 (N_7415,N_5268,N_5282);
or U7416 (N_7416,N_4909,N_5371);
or U7417 (N_7417,N_5712,N_5890);
or U7418 (N_7418,N_4590,N_5147);
xor U7419 (N_7419,N_5362,N_5766);
xor U7420 (N_7420,N_4523,N_4994);
or U7421 (N_7421,N_5151,N_5299);
xor U7422 (N_7422,N_4659,N_5450);
xnor U7423 (N_7423,N_5075,N_5523);
xor U7424 (N_7424,N_5888,N_4586);
and U7425 (N_7425,N_5978,N_5882);
nand U7426 (N_7426,N_4901,N_5314);
nand U7427 (N_7427,N_5617,N_4750);
and U7428 (N_7428,N_4579,N_5637);
nor U7429 (N_7429,N_4752,N_5809);
or U7430 (N_7430,N_5413,N_5028);
xnor U7431 (N_7431,N_5896,N_4705);
xnor U7432 (N_7432,N_5224,N_5703);
xor U7433 (N_7433,N_5565,N_5029);
nor U7434 (N_7434,N_5589,N_5654);
nor U7435 (N_7435,N_4919,N_4748);
and U7436 (N_7436,N_4525,N_5348);
or U7437 (N_7437,N_5612,N_5653);
nor U7438 (N_7438,N_4665,N_4569);
nand U7439 (N_7439,N_5562,N_5471);
nand U7440 (N_7440,N_5852,N_5971);
and U7441 (N_7441,N_5677,N_4541);
or U7442 (N_7442,N_5155,N_5968);
xnor U7443 (N_7443,N_4533,N_5500);
nand U7444 (N_7444,N_5225,N_5639);
nor U7445 (N_7445,N_4878,N_5134);
and U7446 (N_7446,N_4975,N_4510);
or U7447 (N_7447,N_5421,N_4975);
or U7448 (N_7448,N_5657,N_5153);
xnor U7449 (N_7449,N_5300,N_5796);
nand U7450 (N_7450,N_5164,N_4599);
nand U7451 (N_7451,N_5511,N_5666);
nand U7452 (N_7452,N_5145,N_5807);
and U7453 (N_7453,N_5017,N_4774);
nand U7454 (N_7454,N_5268,N_5777);
or U7455 (N_7455,N_5637,N_5948);
or U7456 (N_7456,N_4997,N_5414);
nor U7457 (N_7457,N_4830,N_5539);
or U7458 (N_7458,N_4998,N_5294);
and U7459 (N_7459,N_5289,N_5065);
nand U7460 (N_7460,N_5142,N_5771);
xor U7461 (N_7461,N_5489,N_5803);
nor U7462 (N_7462,N_4642,N_4919);
nor U7463 (N_7463,N_5598,N_5299);
nor U7464 (N_7464,N_5289,N_4846);
nor U7465 (N_7465,N_5989,N_5494);
nand U7466 (N_7466,N_5360,N_5020);
and U7467 (N_7467,N_4693,N_4726);
nand U7468 (N_7468,N_5086,N_5115);
and U7469 (N_7469,N_5610,N_5395);
xor U7470 (N_7470,N_4896,N_4531);
xor U7471 (N_7471,N_5869,N_5674);
and U7472 (N_7472,N_5972,N_5557);
xnor U7473 (N_7473,N_4783,N_4501);
xor U7474 (N_7474,N_5928,N_4962);
or U7475 (N_7475,N_5941,N_5145);
nor U7476 (N_7476,N_4827,N_5092);
nand U7477 (N_7477,N_4751,N_5183);
and U7478 (N_7478,N_5814,N_5881);
nor U7479 (N_7479,N_5797,N_5528);
nand U7480 (N_7480,N_4997,N_4655);
xnor U7481 (N_7481,N_5183,N_5806);
nor U7482 (N_7482,N_4744,N_4707);
nor U7483 (N_7483,N_4632,N_5930);
xor U7484 (N_7484,N_5401,N_5347);
nand U7485 (N_7485,N_5307,N_5849);
nand U7486 (N_7486,N_4808,N_5158);
and U7487 (N_7487,N_4643,N_5112);
xnor U7488 (N_7488,N_5177,N_5928);
or U7489 (N_7489,N_5173,N_5803);
or U7490 (N_7490,N_4753,N_5781);
nand U7491 (N_7491,N_5410,N_4805);
and U7492 (N_7492,N_5588,N_4976);
or U7493 (N_7493,N_4802,N_5461);
and U7494 (N_7494,N_4698,N_4754);
nand U7495 (N_7495,N_5762,N_5672);
nor U7496 (N_7496,N_4641,N_5467);
nand U7497 (N_7497,N_5578,N_4837);
nor U7498 (N_7498,N_5125,N_5809);
nor U7499 (N_7499,N_5704,N_5092);
or U7500 (N_7500,N_6120,N_7013);
nand U7501 (N_7501,N_6160,N_6572);
nand U7502 (N_7502,N_7320,N_6916);
xnor U7503 (N_7503,N_7299,N_7348);
nand U7504 (N_7504,N_7489,N_6668);
and U7505 (N_7505,N_6837,N_7370);
and U7506 (N_7506,N_7279,N_7168);
or U7507 (N_7507,N_6569,N_6355);
xnor U7508 (N_7508,N_6672,N_6301);
nor U7509 (N_7509,N_6548,N_6481);
xor U7510 (N_7510,N_6789,N_6619);
and U7511 (N_7511,N_6831,N_7425);
or U7512 (N_7512,N_6998,N_6248);
nand U7513 (N_7513,N_7100,N_7077);
nand U7514 (N_7514,N_6103,N_7030);
nand U7515 (N_7515,N_7126,N_6943);
nor U7516 (N_7516,N_6760,N_7475);
xor U7517 (N_7517,N_6568,N_6071);
nand U7518 (N_7518,N_7387,N_7223);
nor U7519 (N_7519,N_6231,N_7288);
nor U7520 (N_7520,N_6935,N_6762);
and U7521 (N_7521,N_7280,N_6714);
or U7522 (N_7522,N_7461,N_6726);
nor U7523 (N_7523,N_6681,N_7448);
nor U7524 (N_7524,N_6022,N_6890);
nor U7525 (N_7525,N_6529,N_6086);
xor U7526 (N_7526,N_7263,N_7353);
xor U7527 (N_7527,N_7290,N_6305);
xor U7528 (N_7528,N_6869,N_6618);
and U7529 (N_7529,N_7397,N_6209);
nor U7530 (N_7530,N_6132,N_6982);
xor U7531 (N_7531,N_7275,N_6267);
xnor U7532 (N_7532,N_6639,N_6731);
nand U7533 (N_7533,N_6912,N_6069);
or U7534 (N_7534,N_6676,N_6922);
nand U7535 (N_7535,N_6490,N_6908);
or U7536 (N_7536,N_6854,N_6117);
nand U7537 (N_7537,N_6409,N_6506);
or U7538 (N_7538,N_6723,N_6663);
and U7539 (N_7539,N_7464,N_7486);
nand U7540 (N_7540,N_6246,N_6748);
or U7541 (N_7541,N_6265,N_7191);
xnor U7542 (N_7542,N_6390,N_7453);
and U7543 (N_7543,N_6292,N_6673);
nand U7544 (N_7544,N_7006,N_7333);
nor U7545 (N_7545,N_6695,N_6424);
nand U7546 (N_7546,N_6995,N_6735);
and U7547 (N_7547,N_6013,N_6553);
and U7548 (N_7548,N_6923,N_7197);
or U7549 (N_7549,N_6338,N_6549);
xnor U7550 (N_7550,N_6483,N_7094);
nor U7551 (N_7551,N_7061,N_6072);
nor U7552 (N_7552,N_7154,N_6719);
and U7553 (N_7553,N_6880,N_6848);
xnor U7554 (N_7554,N_6858,N_6394);
or U7555 (N_7555,N_6530,N_6039);
nor U7556 (N_7556,N_6196,N_6147);
nor U7557 (N_7557,N_7024,N_7106);
xnor U7558 (N_7558,N_7091,N_6818);
nand U7559 (N_7559,N_6946,N_6996);
nand U7560 (N_7560,N_6223,N_6392);
xnor U7561 (N_7561,N_6194,N_7241);
and U7562 (N_7562,N_6368,N_6769);
nor U7563 (N_7563,N_7225,N_7146);
xnor U7564 (N_7564,N_6260,N_7322);
or U7565 (N_7565,N_6929,N_6070);
and U7566 (N_7566,N_6232,N_6359);
nor U7567 (N_7567,N_7351,N_6036);
nand U7568 (N_7568,N_6646,N_6849);
nand U7569 (N_7569,N_7075,N_6791);
or U7570 (N_7570,N_7407,N_6757);
and U7571 (N_7571,N_7008,N_6430);
nor U7572 (N_7572,N_7483,N_6012);
nor U7573 (N_7573,N_6520,N_7233);
nand U7574 (N_7574,N_7287,N_6892);
and U7575 (N_7575,N_6893,N_6855);
and U7576 (N_7576,N_6993,N_6488);
nand U7577 (N_7577,N_6289,N_7041);
or U7578 (N_7578,N_7457,N_6614);
and U7579 (N_7579,N_7189,N_7498);
nand U7580 (N_7580,N_6786,N_6242);
nand U7581 (N_7581,N_7270,N_6198);
nor U7582 (N_7582,N_7214,N_6158);
or U7583 (N_7583,N_7449,N_7166);
nor U7584 (N_7584,N_6307,N_7059);
or U7585 (N_7585,N_6253,N_7246);
xnor U7586 (N_7586,N_7156,N_6006);
nor U7587 (N_7587,N_7203,N_7266);
nand U7588 (N_7588,N_6032,N_6244);
and U7589 (N_7589,N_6073,N_6886);
xor U7590 (N_7590,N_6367,N_6299);
nand U7591 (N_7591,N_6050,N_7173);
and U7592 (N_7592,N_6501,N_6959);
xor U7593 (N_7593,N_6396,N_6097);
nand U7594 (N_7594,N_6913,N_6110);
xnor U7595 (N_7595,N_6341,N_7467);
xnor U7596 (N_7596,N_6712,N_6556);
and U7597 (N_7597,N_6397,N_7400);
nor U7598 (N_7598,N_6797,N_6832);
or U7599 (N_7599,N_6531,N_6709);
nor U7600 (N_7600,N_6990,N_6443);
xnor U7601 (N_7601,N_6817,N_7021);
xnor U7602 (N_7602,N_6108,N_6107);
nand U7603 (N_7603,N_7226,N_6128);
nand U7604 (N_7604,N_6985,N_6122);
or U7605 (N_7605,N_7178,N_7128);
or U7606 (N_7606,N_6274,N_7140);
or U7607 (N_7607,N_6452,N_6186);
or U7608 (N_7608,N_6241,N_7070);
or U7609 (N_7609,N_7375,N_6114);
nor U7610 (N_7610,N_7384,N_7155);
and U7611 (N_7611,N_6235,N_6782);
and U7612 (N_7612,N_7216,N_6677);
xor U7613 (N_7613,N_6351,N_6466);
xnor U7614 (N_7614,N_6015,N_7343);
and U7615 (N_7615,N_6846,N_6577);
or U7616 (N_7616,N_6717,N_6251);
xor U7617 (N_7617,N_6428,N_7151);
or U7618 (N_7618,N_6376,N_6016);
and U7619 (N_7619,N_7079,N_7119);
or U7620 (N_7620,N_6809,N_6536);
or U7621 (N_7621,N_6420,N_7081);
xor U7622 (N_7622,N_6062,N_6933);
nand U7623 (N_7623,N_6322,N_7358);
or U7624 (N_7624,N_7098,N_7201);
nor U7625 (N_7625,N_6977,N_7244);
nand U7626 (N_7626,N_6219,N_6736);
nor U7627 (N_7627,N_6840,N_7235);
and U7628 (N_7628,N_6302,N_7002);
nand U7629 (N_7629,N_7108,N_6539);
nand U7630 (N_7630,N_6711,N_7010);
and U7631 (N_7631,N_6578,N_7285);
xnor U7632 (N_7632,N_6391,N_6361);
xor U7633 (N_7633,N_6965,N_6513);
and U7634 (N_7634,N_6872,N_6927);
nor U7635 (N_7635,N_6662,N_6247);
xor U7636 (N_7636,N_6624,N_6090);
nor U7637 (N_7637,N_6727,N_7272);
and U7638 (N_7638,N_6279,N_7310);
or U7639 (N_7639,N_7423,N_7097);
xnor U7640 (N_7640,N_6542,N_6085);
xor U7641 (N_7641,N_6089,N_6528);
xnor U7642 (N_7642,N_6565,N_6525);
nand U7643 (N_7643,N_7090,N_6027);
nand U7644 (N_7644,N_7043,N_6875);
or U7645 (N_7645,N_6199,N_6417);
nor U7646 (N_7646,N_7137,N_7136);
nand U7647 (N_7647,N_7200,N_6824);
and U7648 (N_7648,N_6608,N_6991);
and U7649 (N_7649,N_6213,N_6562);
and U7650 (N_7650,N_6821,N_6802);
and U7651 (N_7651,N_6951,N_7102);
nand U7652 (N_7652,N_7176,N_6534);
and U7653 (N_7653,N_6137,N_7009);
nor U7654 (N_7654,N_6353,N_7324);
nor U7655 (N_7655,N_6220,N_7406);
and U7656 (N_7656,N_6820,N_7293);
nor U7657 (N_7657,N_7190,N_7332);
or U7658 (N_7658,N_7175,N_6187);
and U7659 (N_7659,N_7346,N_6115);
xnor U7660 (N_7660,N_6093,N_6519);
and U7661 (N_7661,N_6078,N_6526);
xor U7662 (N_7662,N_6839,N_6243);
and U7663 (N_7663,N_6871,N_6787);
or U7664 (N_7664,N_6499,N_6701);
nand U7665 (N_7665,N_6370,N_6543);
and U7666 (N_7666,N_6680,N_6540);
and U7667 (N_7667,N_6647,N_6412);
and U7668 (N_7668,N_6945,N_7242);
nand U7669 (N_7669,N_6266,N_6202);
nor U7670 (N_7670,N_6557,N_7307);
and U7671 (N_7671,N_7344,N_6642);
and U7672 (N_7672,N_6868,N_6329);
or U7673 (N_7673,N_7000,N_6617);
nand U7674 (N_7674,N_7488,N_6395);
and U7675 (N_7675,N_7222,N_7305);
or U7676 (N_7676,N_6659,N_7133);
xor U7677 (N_7677,N_6878,N_6947);
nor U7678 (N_7678,N_7085,N_7089);
or U7679 (N_7679,N_6920,N_6427);
xnor U7680 (N_7680,N_6785,N_7491);
nor U7681 (N_7681,N_7329,N_7122);
xnor U7682 (N_7682,N_7007,N_6747);
and U7683 (N_7683,N_7159,N_6864);
nand U7684 (N_7684,N_6522,N_7205);
nor U7685 (N_7685,N_6865,N_7107);
nor U7686 (N_7686,N_6829,N_6643);
xnor U7687 (N_7687,N_6034,N_6626);
nand U7688 (N_7688,N_7112,N_6573);
nor U7689 (N_7689,N_7063,N_6176);
xor U7690 (N_7690,N_6467,N_6105);
nand U7691 (N_7691,N_6127,N_6239);
xor U7692 (N_7692,N_6773,N_6583);
or U7693 (N_7693,N_7012,N_6783);
and U7694 (N_7694,N_6683,N_7217);
and U7695 (N_7695,N_6234,N_6862);
xor U7696 (N_7696,N_6410,N_6560);
or U7697 (N_7697,N_7416,N_7308);
xnor U7698 (N_7698,N_6589,N_6250);
nand U7699 (N_7699,N_6303,N_6166);
and U7700 (N_7700,N_6909,N_7476);
nor U7701 (N_7701,N_6599,N_7269);
nor U7702 (N_7702,N_6502,N_7141);
nand U7703 (N_7703,N_7474,N_7148);
and U7704 (N_7704,N_7158,N_6331);
xnor U7705 (N_7705,N_6371,N_7034);
nor U7706 (N_7706,N_6435,N_6588);
or U7707 (N_7707,N_6358,N_7295);
nor U7708 (N_7708,N_6559,N_6374);
or U7709 (N_7709,N_7150,N_6771);
or U7710 (N_7710,N_6928,N_6067);
and U7711 (N_7711,N_6660,N_6884);
nand U7712 (N_7712,N_6159,N_6124);
xor U7713 (N_7713,N_6068,N_7327);
nand U7714 (N_7714,N_6554,N_6587);
or U7715 (N_7715,N_7111,N_6134);
nand U7716 (N_7716,N_7212,N_6170);
xnor U7717 (N_7717,N_6805,N_6810);
xnor U7718 (N_7718,N_6604,N_6458);
or U7719 (N_7719,N_7183,N_7444);
nand U7720 (N_7720,N_6964,N_6739);
nand U7721 (N_7721,N_6295,N_6171);
and U7722 (N_7722,N_6637,N_6255);
or U7723 (N_7723,N_7447,N_7105);
nand U7724 (N_7724,N_6563,N_6429);
and U7725 (N_7725,N_6294,N_6915);
or U7726 (N_7726,N_6636,N_7347);
or U7727 (N_7727,N_7033,N_6883);
and U7728 (N_7728,N_6335,N_6401);
xnor U7729 (N_7729,N_6230,N_6441);
xor U7730 (N_7730,N_6907,N_6957);
or U7731 (N_7731,N_7236,N_6455);
and U7732 (N_7732,N_7497,N_6189);
and U7733 (N_7733,N_6183,N_6980);
or U7734 (N_7734,N_6896,N_7338);
nand U7735 (N_7735,N_7314,N_6765);
or U7736 (N_7736,N_6753,N_6332);
and U7737 (N_7737,N_6140,N_6104);
nor U7738 (N_7738,N_6261,N_6641);
nand U7739 (N_7739,N_7181,N_6776);
nand U7740 (N_7740,N_6203,N_7393);
and U7741 (N_7741,N_6382,N_6386);
or U7742 (N_7742,N_6009,N_6629);
and U7743 (N_7743,N_6537,N_6208);
and U7744 (N_7744,N_6487,N_6345);
or U7745 (N_7745,N_6888,N_6106);
and U7746 (N_7746,N_6149,N_7401);
and U7747 (N_7747,N_6168,N_7382);
nor U7748 (N_7748,N_7363,N_6432);
nor U7749 (N_7749,N_6779,N_7029);
or U7750 (N_7750,N_7131,N_6986);
nand U7751 (N_7751,N_6906,N_6421);
or U7752 (N_7752,N_6738,N_6635);
nand U7753 (N_7753,N_7139,N_7256);
or U7754 (N_7754,N_7127,N_6764);
nand U7755 (N_7755,N_6602,N_7248);
nor U7756 (N_7756,N_7252,N_6754);
and U7757 (N_7757,N_6669,N_6612);
or U7758 (N_7758,N_7202,N_6477);
and U7759 (N_7759,N_7080,N_6287);
nand U7760 (N_7760,N_6362,N_7328);
xor U7761 (N_7761,N_7035,N_6857);
nor U7762 (N_7762,N_6877,N_6080);
nand U7763 (N_7763,N_6627,N_7428);
xor U7764 (N_7764,N_6347,N_7377);
xnor U7765 (N_7765,N_6224,N_6767);
nor U7766 (N_7766,N_6770,N_6205);
and U7767 (N_7767,N_7392,N_7073);
or U7768 (N_7768,N_7121,N_7462);
nor U7769 (N_7769,N_6121,N_6442);
or U7770 (N_7770,N_6508,N_6277);
xnor U7771 (N_7771,N_6592,N_6378);
nor U7772 (N_7772,N_6237,N_7004);
nor U7773 (N_7773,N_6112,N_6030);
or U7774 (N_7774,N_6807,N_6879);
or U7775 (N_7775,N_6111,N_7083);
nor U7776 (N_7776,N_7240,N_6190);
and U7777 (N_7777,N_7101,N_6413);
and U7778 (N_7778,N_6418,N_6628);
nand U7779 (N_7779,N_7317,N_6609);
nor U7780 (N_7780,N_6590,N_6567);
nor U7781 (N_7781,N_6264,N_6968);
and U7782 (N_7782,N_7412,N_7039);
nor U7783 (N_7783,N_6450,N_7326);
nor U7784 (N_7784,N_6285,N_6297);
nand U7785 (N_7785,N_6507,N_6552);
and U7786 (N_7786,N_6276,N_6052);
and U7787 (N_7787,N_7169,N_7262);
nor U7788 (N_7788,N_6698,N_7231);
nor U7789 (N_7789,N_6010,N_6280);
nor U7790 (N_7790,N_6055,N_7422);
and U7791 (N_7791,N_6473,N_6720);
xnor U7792 (N_7792,N_6970,N_6045);
nand U7793 (N_7793,N_6486,N_6262);
xnor U7794 (N_7794,N_7334,N_7078);
or U7795 (N_7795,N_6218,N_7493);
xor U7796 (N_7796,N_7067,N_6252);
and U7797 (N_7797,N_6570,N_6504);
nor U7798 (N_7798,N_6925,N_6227);
or U7799 (N_7799,N_7250,N_6752);
nor U7800 (N_7800,N_7345,N_7357);
nand U7801 (N_7801,N_6891,N_7415);
xnor U7802 (N_7802,N_6425,N_7389);
or U7803 (N_7803,N_7204,N_7304);
or U7804 (N_7804,N_6611,N_6154);
and U7805 (N_7805,N_7220,N_6269);
nor U7806 (N_7806,N_6622,N_7051);
and U7807 (N_7807,N_6705,N_7047);
nor U7808 (N_7808,N_6257,N_6216);
or U7809 (N_7809,N_7315,N_6703);
or U7810 (N_7810,N_6532,N_6087);
nor U7811 (N_7811,N_6324,N_6256);
xnor U7812 (N_7812,N_7038,N_6098);
nand U7813 (N_7813,N_6650,N_6161);
nor U7814 (N_7814,N_7103,N_6037);
nand U7815 (N_7815,N_7247,N_6966);
or U7816 (N_7816,N_6498,N_6685);
nand U7817 (N_7817,N_7048,N_7277);
and U7818 (N_7818,N_6902,N_6060);
nor U7819 (N_7819,N_7452,N_6517);
nand U7820 (N_7820,N_6480,N_6434);
xnor U7821 (N_7821,N_6623,N_6291);
nor U7822 (N_7822,N_7441,N_7433);
nor U7823 (N_7823,N_6873,N_6400);
nor U7824 (N_7824,N_6874,N_6372);
nand U7825 (N_7825,N_6679,N_7074);
and U7826 (N_7826,N_6579,N_6591);
xor U7827 (N_7827,N_6828,N_7227);
xor U7828 (N_7828,N_7254,N_6638);
xor U7829 (N_7829,N_6598,N_6984);
and U7830 (N_7830,N_7228,N_6162);
or U7831 (N_7831,N_6926,N_7469);
or U7832 (N_7832,N_6066,N_7022);
or U7833 (N_7833,N_6939,N_6387);
or U7834 (N_7834,N_6919,N_6942);
or U7835 (N_7835,N_7463,N_6155);
nand U7836 (N_7836,N_7300,N_6388);
or U7837 (N_7837,N_6349,N_6475);
nand U7838 (N_7838,N_6179,N_6706);
or U7839 (N_7839,N_6164,N_6142);
or U7840 (N_7840,N_6309,N_6950);
nand U7841 (N_7841,N_7352,N_6798);
or U7842 (N_7842,N_6803,N_7005);
nor U7843 (N_7843,N_6393,N_6687);
nand U7844 (N_7844,N_6585,N_6233);
nand U7845 (N_7845,N_7420,N_6304);
or U7846 (N_7846,N_6897,N_7208);
or U7847 (N_7847,N_7411,N_6894);
nand U7848 (N_7848,N_6917,N_6887);
and U7849 (N_7849,N_7219,N_6236);
and U7850 (N_7850,N_7003,N_6594);
nand U7851 (N_7851,N_7198,N_7120);
xor U7852 (N_7852,N_7062,N_7257);
or U7853 (N_7853,N_6876,N_7193);
or U7854 (N_7854,N_7330,N_6664);
nand U7855 (N_7855,N_7323,N_6937);
and U7856 (N_7856,N_6094,N_7454);
xnor U7857 (N_7857,N_7408,N_6206);
or U7858 (N_7858,N_7028,N_6621);
nand U7859 (N_7859,N_6713,N_7138);
nor U7860 (N_7860,N_7117,N_6652);
xnor U7861 (N_7861,N_6651,N_6983);
and U7862 (N_7862,N_6582,N_7395);
or U7863 (N_7863,N_7276,N_6457);
or U7864 (N_7864,N_7410,N_6981);
or U7865 (N_7865,N_6956,N_6180);
nor U7866 (N_7866,N_7068,N_7490);
nand U7867 (N_7867,N_6328,N_6509);
nand U7868 (N_7868,N_7360,N_6742);
nor U7869 (N_7869,N_7368,N_6576);
or U7870 (N_7870,N_6156,N_7229);
and U7871 (N_7871,N_6047,N_6150);
nand U7872 (N_7872,N_6924,N_7273);
and U7873 (N_7873,N_6023,N_6340);
and U7874 (N_7874,N_6722,N_7499);
xor U7875 (N_7875,N_7109,N_7292);
nand U7876 (N_7876,N_6750,N_6082);
nand U7877 (N_7877,N_6700,N_6385);
nor U7878 (N_7878,N_7278,N_6311);
and U7879 (N_7879,N_7088,N_6973);
nand U7880 (N_7880,N_7485,N_6172);
or U7881 (N_7881,N_7232,N_7113);
or U7882 (N_7882,N_6408,N_6586);
and U7883 (N_7883,N_7355,N_7342);
xor U7884 (N_7884,N_6002,N_6157);
xnor U7885 (N_7885,N_6325,N_6661);
nor U7886 (N_7886,N_6333,N_6063);
or U7887 (N_7887,N_6476,N_6535);
and U7888 (N_7888,N_7437,N_6138);
xor U7889 (N_7889,N_6046,N_6356);
nor U7890 (N_7890,N_7291,N_6384);
and U7891 (N_7891,N_6497,N_6028);
nand U7892 (N_7892,N_7398,N_7157);
nand U7893 (N_7893,N_7045,N_7367);
or U7894 (N_7894,N_7152,N_6263);
and U7895 (N_7895,N_6215,N_6270);
and U7896 (N_7896,N_6479,N_6018);
xnor U7897 (N_7897,N_7218,N_6383);
or U7898 (N_7898,N_6744,N_6492);
nand U7899 (N_7899,N_6035,N_6099);
xor U7900 (N_7900,N_7414,N_6249);
nand U7901 (N_7901,N_6694,N_6667);
or U7902 (N_7902,N_7302,N_7224);
or U7903 (N_7903,N_6029,N_6976);
nand U7904 (N_7904,N_6640,N_6228);
or U7905 (N_7905,N_6240,N_6584);
or U7906 (N_7906,N_6468,N_6905);
or U7907 (N_7907,N_7480,N_7471);
and U7908 (N_7908,N_6702,N_6881);
xnor U7909 (N_7909,N_6348,N_6343);
xnor U7910 (N_7910,N_6987,N_6900);
xnor U7911 (N_7911,N_7267,N_7056);
xor U7912 (N_7912,N_6008,N_6489);
nand U7913 (N_7913,N_6403,N_6146);
or U7914 (N_7914,N_7478,N_7366);
and U7915 (N_7915,N_7016,N_6399);
xor U7916 (N_7916,N_6955,N_6523);
xor U7917 (N_7917,N_7147,N_7296);
nand U7918 (N_7918,N_7430,N_7477);
and U7919 (N_7919,N_6139,N_6564);
nand U7920 (N_7920,N_7429,N_7072);
nor U7921 (N_7921,N_7192,N_7130);
nand U7922 (N_7922,N_6377,N_7372);
nor U7923 (N_7923,N_7361,N_6775);
nor U7924 (N_7924,N_6281,N_7115);
and U7925 (N_7925,N_6931,N_6648);
or U7926 (N_7926,N_6566,N_7238);
nor U7927 (N_7927,N_7135,N_7015);
nand U7928 (N_7928,N_6729,N_6684);
xor U7929 (N_7929,N_6019,N_6152);
nor U7930 (N_7930,N_6516,N_6954);
xor U7931 (N_7931,N_7470,N_7268);
nor U7932 (N_7932,N_6630,N_7417);
and U7933 (N_7933,N_6352,N_6431);
nand U7934 (N_7934,N_6949,N_6484);
nor U7935 (N_7935,N_6439,N_6366);
nand U7936 (N_7936,N_6318,N_6320);
or U7937 (N_7937,N_6800,N_6766);
xnor U7938 (N_7938,N_6632,N_6173);
nand U7939 (N_7939,N_6426,N_6469);
and U7940 (N_7940,N_7456,N_6795);
or U7941 (N_7941,N_6058,N_6064);
and U7942 (N_7942,N_6859,N_6153);
or U7943 (N_7943,N_6181,N_7055);
and U7944 (N_7944,N_6020,N_7496);
nor U7945 (N_7945,N_6436,N_6689);
nand U7946 (N_7946,N_7259,N_6823);
or U7947 (N_7947,N_6607,N_6021);
or U7948 (N_7948,N_6169,N_6781);
nor U7949 (N_7949,N_6038,N_7298);
nand U7950 (N_7950,N_6518,N_6671);
nand U7951 (N_7951,N_7084,N_6414);
and U7952 (N_7952,N_6645,N_7432);
xnor U7953 (N_7953,N_6379,N_6844);
and U7954 (N_7954,N_6461,N_7142);
or U7955 (N_7955,N_7185,N_7132);
nand U7956 (N_7956,N_7032,N_6616);
nand U7957 (N_7957,N_7284,N_6811);
or U7958 (N_7958,N_7439,N_7093);
nand U7959 (N_7959,N_6545,N_6211);
nand U7960 (N_7960,N_6521,N_6992);
and U7961 (N_7961,N_6938,N_7435);
nand U7962 (N_7962,N_7162,N_6524);
nand U7963 (N_7963,N_6188,N_7194);
and U7964 (N_7964,N_6195,N_6282);
nand U7965 (N_7965,N_7446,N_6278);
or U7966 (N_7966,N_6596,N_7466);
xor U7967 (N_7967,N_6048,N_6245);
xnor U7968 (N_7968,N_6288,N_6081);
xor U7969 (N_7969,N_6315,N_6551);
nor U7970 (N_7970,N_6088,N_6936);
nor U7971 (N_7971,N_6808,N_6631);
nand U7972 (N_7972,N_7170,N_6836);
nand U7973 (N_7973,N_7260,N_7354);
xor U7974 (N_7974,N_6686,N_7057);
nor U7975 (N_7975,N_6095,N_6710);
xor U7976 (N_7976,N_6784,N_7378);
nor U7977 (N_7977,N_7054,N_6972);
xor U7978 (N_7978,N_6960,N_6313);
and U7979 (N_7979,N_6999,N_7206);
nor U7980 (N_7980,N_7396,N_6963);
nand U7981 (N_7981,N_7442,N_7438);
nor U7982 (N_7982,N_6734,N_6512);
nand U7983 (N_7983,N_6474,N_6838);
xnor U7984 (N_7984,N_6365,N_6699);
nor U7985 (N_7985,N_7014,N_7369);
nand U7986 (N_7986,N_6024,N_6268);
nand U7987 (N_7987,N_6780,N_6889);
nand U7988 (N_7988,N_7019,N_6944);
xor U7989 (N_7989,N_6721,N_7373);
and U7990 (N_7990,N_6674,N_6969);
nand U7991 (N_7991,N_7379,N_7443);
nand U7992 (N_7992,N_7405,N_6449);
nand U7993 (N_7993,N_7243,N_7472);
and U7994 (N_7994,N_6841,N_6197);
or U7995 (N_7995,N_7311,N_7011);
and U7996 (N_7996,N_7149,N_6415);
and U7997 (N_7997,N_7195,N_6581);
or U7998 (N_7998,N_6059,N_6751);
nand U7999 (N_7999,N_6774,N_6077);
nor U8000 (N_8000,N_7281,N_6192);
nand U8001 (N_8001,N_6496,N_6126);
xnor U8002 (N_8002,N_7318,N_7255);
nor U8003 (N_8003,N_6763,N_6193);
nor U8004 (N_8004,N_7086,N_7163);
or U8005 (N_8005,N_6514,N_6541);
or U8006 (N_8006,N_6593,N_7445);
nand U8007 (N_8007,N_6041,N_7371);
nor U8008 (N_8008,N_6327,N_7099);
nor U8009 (N_8009,N_6463,N_6113);
and U8010 (N_8010,N_6678,N_6207);
nand U8011 (N_8011,N_7264,N_6571);
xnor U8012 (N_8012,N_6918,N_6438);
or U8013 (N_8013,N_6042,N_6603);
nand U8014 (N_8014,N_6538,N_6655);
nand U8015 (N_8015,N_6454,N_7309);
nand U8016 (N_8016,N_7376,N_6422);
and U8017 (N_8017,N_6336,N_6580);
nor U8018 (N_8018,N_6478,N_7071);
or U8019 (N_8019,N_6238,N_6011);
xor U8020 (N_8020,N_7110,N_6494);
nor U8021 (N_8021,N_6119,N_6357);
or U8022 (N_8022,N_7144,N_7118);
nand U8023 (N_8023,N_7313,N_6561);
xnor U8024 (N_8024,N_7383,N_6404);
xor U8025 (N_8025,N_6411,N_6437);
or U8026 (N_8026,N_6856,N_7385);
nor U8027 (N_8027,N_6952,N_7306);
and U8028 (N_8028,N_7286,N_6101);
or U8029 (N_8029,N_6204,N_6056);
nand U8030 (N_8030,N_6555,N_6283);
xor U8031 (N_8031,N_7335,N_7044);
and U8032 (N_8032,N_7455,N_7481);
xor U8033 (N_8033,N_6445,N_7321);
nor U8034 (N_8034,N_7040,N_6813);
nand U8035 (N_8035,N_6574,N_6904);
nand U8036 (N_8036,N_6932,N_7271);
and U8037 (N_8037,N_6495,N_6953);
and U8038 (N_8038,N_7245,N_6974);
nor U8039 (N_8039,N_6148,N_6812);
nand U8040 (N_8040,N_6544,N_6174);
and U8041 (N_8041,N_6842,N_7188);
or U8042 (N_8042,N_6527,N_6910);
nor U8043 (N_8043,N_6003,N_6930);
and U8044 (N_8044,N_6136,N_6749);
xor U8045 (N_8045,N_7312,N_6040);
nand U8046 (N_8046,N_6471,N_7125);
and U8047 (N_8047,N_7403,N_6100);
nor U8048 (N_8048,N_6547,N_6860);
nand U8049 (N_8049,N_7082,N_6914);
xnor U8050 (N_8050,N_6716,N_6321);
or U8051 (N_8051,N_6360,N_6272);
nand U8052 (N_8052,N_7186,N_7164);
or U8053 (N_8053,N_6462,N_6123);
xnor U8054 (N_8054,N_6053,N_6882);
xnor U8055 (N_8055,N_7213,N_6354);
and U8056 (N_8056,N_7134,N_6004);
nand U8057 (N_8057,N_7046,N_6144);
or U8058 (N_8058,N_6696,N_6819);
or U8059 (N_8059,N_6482,N_7209);
nand U8060 (N_8060,N_6001,N_6755);
xor U8061 (N_8061,N_6334,N_7116);
and U8062 (N_8062,N_6296,N_6778);
xor U8063 (N_8063,N_7171,N_6866);
nor U8064 (N_8064,N_6133,N_7399);
xor U8065 (N_8065,N_7258,N_6118);
xnor U8066 (N_8066,N_6286,N_7095);
and U8067 (N_8067,N_7386,N_7388);
nor U8068 (N_8068,N_7440,N_7274);
nor U8069 (N_8069,N_6440,N_6310);
and U8070 (N_8070,N_7418,N_6342);
xor U8071 (N_8071,N_6201,N_6725);
or U8072 (N_8072,N_6323,N_6373);
xnor U8073 (N_8073,N_6448,N_6826);
and U8074 (N_8074,N_7283,N_6690);
nor U8075 (N_8075,N_7282,N_7336);
or U8076 (N_8076,N_7374,N_6693);
xnor U8077 (N_8077,N_6258,N_6708);
xor U8078 (N_8078,N_6314,N_6625);
nor U8079 (N_8079,N_6834,N_6790);
nand U8080 (N_8080,N_7025,N_6273);
or U8081 (N_8081,N_7460,N_6740);
nor U8082 (N_8082,N_7380,N_7172);
and U8083 (N_8083,N_7349,N_6326);
xor U8084 (N_8084,N_6804,N_6758);
and U8085 (N_8085,N_7419,N_6899);
and U8086 (N_8086,N_6948,N_6165);
xnor U8087 (N_8087,N_7319,N_6337);
nand U8088 (N_8088,N_7161,N_6033);
nand U8089 (N_8089,N_7356,N_7421);
or U8090 (N_8090,N_6178,N_6306);
and U8091 (N_8091,N_7426,N_6691);
nor U8092 (N_8092,N_6670,N_7087);
and U8093 (N_8093,N_7187,N_6962);
xor U8094 (N_8094,N_6026,N_7468);
or U8095 (N_8095,N_7301,N_6167);
nor U8096 (N_8096,N_6654,N_7066);
and U8097 (N_8097,N_6911,N_6298);
nor U8098 (N_8098,N_6191,N_6921);
or U8099 (N_8099,N_7482,N_6835);
xor U8100 (N_8100,N_7114,N_7065);
nand U8101 (N_8101,N_6460,N_6444);
and U8102 (N_8102,N_6605,N_6316);
nand U8103 (N_8103,N_6451,N_7221);
xor U8104 (N_8104,N_7069,N_7153);
or U8105 (N_8105,N_7325,N_7196);
nand U8106 (N_8106,N_6017,N_6402);
or U8107 (N_8107,N_6092,N_6845);
xor U8108 (N_8108,N_7123,N_6433);
nor U8109 (N_8109,N_6346,N_7215);
nand U8110 (N_8110,N_6275,N_6746);
and U8111 (N_8111,N_7341,N_6515);
nor U8112 (N_8112,N_6657,N_7331);
and U8113 (N_8113,N_6788,N_7167);
nor U8114 (N_8114,N_6792,N_6000);
nand U8115 (N_8115,N_7340,N_6822);
xor U8116 (N_8116,N_6453,N_7492);
xor U8117 (N_8117,N_6682,N_7207);
nor U8118 (N_8118,N_7424,N_7145);
and U8119 (N_8119,N_6885,N_6732);
nand U8120 (N_8120,N_6730,N_6075);
and U8121 (N_8121,N_6109,N_6049);
nand U8122 (N_8122,N_7018,N_6491);
xnor U8123 (N_8123,N_6472,N_7049);
xnor U8124 (N_8124,N_6743,N_6794);
or U8125 (N_8125,N_6610,N_6125);
nand U8126 (N_8126,N_6074,N_6850);
nand U8127 (N_8127,N_7359,N_6533);
or U8128 (N_8128,N_6141,N_6419);
nor U8129 (N_8129,N_6503,N_7316);
nand U8130 (N_8130,N_6416,N_6459);
and U8131 (N_8131,N_6129,N_6423);
nand U8132 (N_8132,N_6546,N_6044);
and U8133 (N_8133,N_6656,N_6130);
or U8134 (N_8134,N_6284,N_6761);
nand U8135 (N_8135,N_6505,N_7391);
xor U8136 (N_8136,N_6575,N_6665);
nand U8137 (N_8137,N_7265,N_6606);
nor U8138 (N_8138,N_6025,N_6200);
or U8139 (N_8139,N_6851,N_7165);
or U8140 (N_8140,N_7184,N_6697);
and U8141 (N_8141,N_6806,N_6903);
or U8142 (N_8142,N_6330,N_6317);
or U8143 (N_8143,N_7365,N_6259);
xnor U8144 (N_8144,N_6975,N_6979);
or U8145 (N_8145,N_7473,N_7031);
nand U8146 (N_8146,N_6091,N_6600);
and U8147 (N_8147,N_7042,N_6051);
and U8148 (N_8148,N_6380,N_6843);
or U8149 (N_8149,N_7199,N_6210);
or U8150 (N_8150,N_6465,N_6801);
nand U8151 (N_8151,N_6633,N_7494);
nand U8152 (N_8152,N_7058,N_6079);
nor U8153 (N_8153,N_6217,N_6369);
or U8154 (N_8154,N_6500,N_7253);
nand U8155 (N_8155,N_6151,N_6407);
or U8156 (N_8156,N_7210,N_6978);
nand U8157 (N_8157,N_7020,N_6116);
and U8158 (N_8158,N_6212,N_6221);
or U8159 (N_8159,N_7237,N_6300);
or U8160 (N_8160,N_6398,N_6961);
nor U8161 (N_8161,N_7053,N_6934);
and U8162 (N_8162,N_6061,N_6861);
xnor U8163 (N_8163,N_6737,N_6350);
nor U8164 (N_8164,N_6901,N_6102);
or U8165 (N_8165,N_6759,N_6005);
nor U8166 (N_8166,N_6615,N_6014);
and U8167 (N_8167,N_6595,N_6756);
nand U8168 (N_8168,N_7458,N_7180);
xor U8169 (N_8169,N_6704,N_6406);
xnor U8170 (N_8170,N_6511,N_6988);
and U8171 (N_8171,N_6816,N_6863);
or U8172 (N_8172,N_6815,N_6793);
nor U8173 (N_8173,N_6895,N_6644);
and U8174 (N_8174,N_7023,N_6182);
nand U8175 (N_8175,N_7001,N_7431);
nor U8176 (N_8176,N_6226,N_6363);
and U8177 (N_8177,N_7394,N_7350);
and U8178 (N_8178,N_6084,N_6364);
or U8179 (N_8179,N_7402,N_7104);
xor U8180 (N_8180,N_7434,N_6043);
nor U8181 (N_8181,N_6688,N_6825);
xor U8182 (N_8182,N_6225,N_6745);
nand U8183 (N_8183,N_6558,N_7230);
nor U8184 (N_8184,N_6796,N_6707);
or U8185 (N_8185,N_6852,N_6184);
nor U8186 (N_8186,N_6971,N_6007);
nand U8187 (N_8187,N_6083,N_7465);
nand U8188 (N_8188,N_6613,N_6339);
and U8189 (N_8189,N_7037,N_7249);
and U8190 (N_8190,N_6456,N_7427);
nand U8191 (N_8191,N_7177,N_6131);
nand U8192 (N_8192,N_7436,N_6649);
nor U8193 (N_8193,N_6675,N_6389);
nand U8194 (N_8194,N_6847,N_7182);
or U8195 (N_8195,N_6493,N_6741);
nand U8196 (N_8196,N_7495,N_7027);
and U8197 (N_8197,N_6344,N_6620);
or U8198 (N_8198,N_6692,N_6728);
nand U8199 (N_8199,N_7036,N_7381);
and U8200 (N_8200,N_6446,N_7064);
or U8201 (N_8201,N_6031,N_6941);
and U8202 (N_8202,N_7294,N_6733);
xor U8203 (N_8203,N_7450,N_7017);
nor U8204 (N_8204,N_6485,N_6799);
nor U8205 (N_8205,N_6827,N_7076);
or U8206 (N_8206,N_6177,N_6989);
nand U8207 (N_8207,N_7390,N_7129);
xor U8208 (N_8208,N_6054,N_6653);
and U8209 (N_8209,N_7261,N_7096);
nand U8210 (N_8210,N_6163,N_6814);
xnor U8211 (N_8211,N_6229,N_7362);
xor U8212 (N_8212,N_6853,N_7337);
and U8213 (N_8213,N_7234,N_6293);
or U8214 (N_8214,N_6958,N_6254);
nor U8215 (N_8215,N_6464,N_7179);
and U8216 (N_8216,N_6308,N_6870);
xnor U8217 (N_8217,N_7409,N_6867);
xnor U8218 (N_8218,N_7339,N_7289);
and U8219 (N_8219,N_7459,N_6718);
nand U8220 (N_8220,N_7404,N_6076);
nand U8221 (N_8221,N_6214,N_6375);
xor U8222 (N_8222,N_7297,N_7124);
xor U8223 (N_8223,N_7487,N_6724);
or U8224 (N_8224,N_6601,N_6222);
or U8225 (N_8225,N_7451,N_6175);
and U8226 (N_8226,N_7303,N_6997);
or U8227 (N_8227,N_6768,N_6994);
nor U8228 (N_8228,N_6597,N_6898);
and U8229 (N_8229,N_6830,N_6470);
xor U8230 (N_8230,N_7143,N_7052);
xnor U8231 (N_8231,N_7092,N_6312);
or U8232 (N_8232,N_6290,N_6143);
xor U8233 (N_8233,N_6065,N_7160);
nand U8234 (N_8234,N_6271,N_6772);
xnor U8235 (N_8235,N_6185,N_7050);
or U8236 (N_8236,N_6096,N_6634);
nor U8237 (N_8237,N_6381,N_6940);
nor U8238 (N_8238,N_6666,N_6658);
nor U8239 (N_8239,N_7251,N_6510);
or U8240 (N_8240,N_7239,N_6447);
or U8241 (N_8241,N_6135,N_6057);
nor U8242 (N_8242,N_7479,N_6319);
nand U8243 (N_8243,N_6777,N_6967);
xnor U8244 (N_8244,N_6405,N_7174);
and U8245 (N_8245,N_7060,N_6833);
and U8246 (N_8246,N_7484,N_6715);
nor U8247 (N_8247,N_7211,N_7364);
or U8248 (N_8248,N_7413,N_7026);
nand U8249 (N_8249,N_6550,N_6145);
nor U8250 (N_8250,N_7224,N_7380);
xnor U8251 (N_8251,N_7050,N_6335);
nor U8252 (N_8252,N_6658,N_6803);
xor U8253 (N_8253,N_7297,N_6592);
xnor U8254 (N_8254,N_6557,N_6812);
xor U8255 (N_8255,N_6725,N_6551);
nor U8256 (N_8256,N_7192,N_6760);
xor U8257 (N_8257,N_6576,N_7375);
or U8258 (N_8258,N_6943,N_7127);
nand U8259 (N_8259,N_6866,N_6153);
nand U8260 (N_8260,N_6915,N_6140);
and U8261 (N_8261,N_7239,N_6018);
nor U8262 (N_8262,N_7390,N_6854);
xor U8263 (N_8263,N_6060,N_6887);
nand U8264 (N_8264,N_6183,N_6015);
and U8265 (N_8265,N_7040,N_7157);
and U8266 (N_8266,N_6754,N_7240);
xnor U8267 (N_8267,N_6298,N_7089);
nand U8268 (N_8268,N_7309,N_7220);
nor U8269 (N_8269,N_6975,N_7399);
and U8270 (N_8270,N_6511,N_6186);
or U8271 (N_8271,N_7044,N_6699);
or U8272 (N_8272,N_7194,N_6474);
or U8273 (N_8273,N_6560,N_7062);
nand U8274 (N_8274,N_7277,N_6454);
and U8275 (N_8275,N_6410,N_7013);
or U8276 (N_8276,N_6888,N_6493);
nor U8277 (N_8277,N_6441,N_6450);
and U8278 (N_8278,N_7373,N_7232);
or U8279 (N_8279,N_6971,N_7342);
or U8280 (N_8280,N_6585,N_7326);
nor U8281 (N_8281,N_6368,N_6445);
and U8282 (N_8282,N_6312,N_6870);
or U8283 (N_8283,N_6935,N_7180);
or U8284 (N_8284,N_6269,N_6473);
nand U8285 (N_8285,N_7475,N_6548);
nor U8286 (N_8286,N_7269,N_7036);
nor U8287 (N_8287,N_7419,N_7354);
xor U8288 (N_8288,N_6637,N_6951);
xor U8289 (N_8289,N_6816,N_6554);
or U8290 (N_8290,N_6947,N_7408);
or U8291 (N_8291,N_7075,N_6602);
nor U8292 (N_8292,N_6920,N_6353);
or U8293 (N_8293,N_6474,N_7023);
xor U8294 (N_8294,N_6936,N_6338);
or U8295 (N_8295,N_6320,N_6076);
and U8296 (N_8296,N_6451,N_6742);
nand U8297 (N_8297,N_7473,N_7248);
xor U8298 (N_8298,N_6870,N_7360);
and U8299 (N_8299,N_7493,N_7222);
nand U8300 (N_8300,N_6854,N_6874);
xor U8301 (N_8301,N_6021,N_6871);
or U8302 (N_8302,N_6084,N_6915);
or U8303 (N_8303,N_6203,N_7168);
nand U8304 (N_8304,N_7102,N_6557);
nand U8305 (N_8305,N_6832,N_6177);
nand U8306 (N_8306,N_6506,N_7222);
nor U8307 (N_8307,N_6821,N_6330);
nor U8308 (N_8308,N_7111,N_7077);
and U8309 (N_8309,N_6317,N_6218);
xnor U8310 (N_8310,N_6594,N_6866);
and U8311 (N_8311,N_6944,N_6209);
nor U8312 (N_8312,N_7442,N_6283);
and U8313 (N_8313,N_6869,N_6450);
or U8314 (N_8314,N_6574,N_7462);
nor U8315 (N_8315,N_6409,N_7330);
nor U8316 (N_8316,N_6598,N_6968);
nor U8317 (N_8317,N_6102,N_6376);
nand U8318 (N_8318,N_6175,N_6484);
or U8319 (N_8319,N_7122,N_7478);
xor U8320 (N_8320,N_6823,N_6485);
nor U8321 (N_8321,N_6469,N_6763);
nor U8322 (N_8322,N_6090,N_7245);
nor U8323 (N_8323,N_6049,N_6812);
and U8324 (N_8324,N_6532,N_7361);
nand U8325 (N_8325,N_6646,N_6902);
nand U8326 (N_8326,N_7134,N_6267);
or U8327 (N_8327,N_7102,N_6496);
nand U8328 (N_8328,N_7186,N_7031);
nand U8329 (N_8329,N_6274,N_6438);
nand U8330 (N_8330,N_6056,N_6275);
xor U8331 (N_8331,N_6779,N_6053);
nand U8332 (N_8332,N_7488,N_6659);
or U8333 (N_8333,N_7244,N_6712);
and U8334 (N_8334,N_6820,N_7273);
xnor U8335 (N_8335,N_7411,N_7319);
and U8336 (N_8336,N_7169,N_7214);
or U8337 (N_8337,N_7066,N_6672);
nor U8338 (N_8338,N_6732,N_6241);
nand U8339 (N_8339,N_6269,N_7178);
xnor U8340 (N_8340,N_6636,N_7070);
or U8341 (N_8341,N_6335,N_6470);
xnor U8342 (N_8342,N_6809,N_6434);
nor U8343 (N_8343,N_7199,N_7473);
and U8344 (N_8344,N_6261,N_6554);
nand U8345 (N_8345,N_6735,N_6856);
nor U8346 (N_8346,N_7496,N_7261);
xnor U8347 (N_8347,N_6183,N_7010);
nand U8348 (N_8348,N_7447,N_6033);
xor U8349 (N_8349,N_7400,N_7119);
or U8350 (N_8350,N_6742,N_6190);
xor U8351 (N_8351,N_6596,N_6946);
nor U8352 (N_8352,N_6521,N_6774);
and U8353 (N_8353,N_6750,N_6316);
or U8354 (N_8354,N_7275,N_7114);
nand U8355 (N_8355,N_6189,N_7222);
xor U8356 (N_8356,N_6595,N_6777);
and U8357 (N_8357,N_6717,N_6004);
xor U8358 (N_8358,N_7044,N_6698);
xor U8359 (N_8359,N_6713,N_7238);
nand U8360 (N_8360,N_7440,N_7388);
xnor U8361 (N_8361,N_7270,N_7264);
xnor U8362 (N_8362,N_7094,N_6137);
xnor U8363 (N_8363,N_6636,N_6615);
nand U8364 (N_8364,N_7201,N_6913);
nor U8365 (N_8365,N_6485,N_7430);
nand U8366 (N_8366,N_7019,N_7298);
nand U8367 (N_8367,N_7165,N_6501);
and U8368 (N_8368,N_6796,N_6649);
and U8369 (N_8369,N_6559,N_6522);
nand U8370 (N_8370,N_7092,N_6702);
nor U8371 (N_8371,N_7427,N_7053);
xnor U8372 (N_8372,N_6390,N_6762);
and U8373 (N_8373,N_6865,N_7163);
nand U8374 (N_8374,N_6004,N_6411);
nand U8375 (N_8375,N_6161,N_7083);
and U8376 (N_8376,N_6837,N_6102);
nor U8377 (N_8377,N_7187,N_7432);
nand U8378 (N_8378,N_6991,N_6961);
nor U8379 (N_8379,N_6858,N_7095);
nand U8380 (N_8380,N_7020,N_7136);
xnor U8381 (N_8381,N_6212,N_7358);
nand U8382 (N_8382,N_6902,N_6876);
or U8383 (N_8383,N_7005,N_6530);
nor U8384 (N_8384,N_6128,N_6114);
nand U8385 (N_8385,N_6490,N_6287);
nor U8386 (N_8386,N_7078,N_7138);
nor U8387 (N_8387,N_6429,N_6097);
and U8388 (N_8388,N_6331,N_7024);
xnor U8389 (N_8389,N_7313,N_6632);
or U8390 (N_8390,N_6408,N_7185);
nor U8391 (N_8391,N_6146,N_6514);
nor U8392 (N_8392,N_6951,N_7252);
nand U8393 (N_8393,N_6125,N_6114);
or U8394 (N_8394,N_6232,N_6592);
nand U8395 (N_8395,N_6119,N_6362);
and U8396 (N_8396,N_7157,N_7384);
nand U8397 (N_8397,N_6182,N_6711);
nand U8398 (N_8398,N_6346,N_7354);
and U8399 (N_8399,N_7229,N_7343);
nor U8400 (N_8400,N_6346,N_7330);
and U8401 (N_8401,N_6811,N_6378);
nor U8402 (N_8402,N_6924,N_6389);
or U8403 (N_8403,N_6264,N_7010);
nand U8404 (N_8404,N_6570,N_7278);
and U8405 (N_8405,N_6293,N_6823);
or U8406 (N_8406,N_6435,N_7078);
and U8407 (N_8407,N_6844,N_6306);
nand U8408 (N_8408,N_6529,N_6778);
nor U8409 (N_8409,N_7128,N_6037);
and U8410 (N_8410,N_6751,N_6319);
and U8411 (N_8411,N_6139,N_6472);
nand U8412 (N_8412,N_6201,N_6318);
or U8413 (N_8413,N_6725,N_6226);
nor U8414 (N_8414,N_6619,N_7113);
nand U8415 (N_8415,N_6597,N_7343);
nor U8416 (N_8416,N_6454,N_6638);
nand U8417 (N_8417,N_6695,N_7155);
xnor U8418 (N_8418,N_6005,N_6764);
nor U8419 (N_8419,N_7438,N_7407);
xnor U8420 (N_8420,N_6513,N_6698);
and U8421 (N_8421,N_6951,N_7372);
nand U8422 (N_8422,N_7126,N_6809);
nor U8423 (N_8423,N_6836,N_7472);
or U8424 (N_8424,N_7310,N_6536);
xor U8425 (N_8425,N_6817,N_7423);
nor U8426 (N_8426,N_6214,N_6355);
nand U8427 (N_8427,N_6021,N_6249);
or U8428 (N_8428,N_7267,N_6357);
and U8429 (N_8429,N_7426,N_6010);
xnor U8430 (N_8430,N_7407,N_6383);
nor U8431 (N_8431,N_6530,N_6535);
xnor U8432 (N_8432,N_6090,N_6470);
and U8433 (N_8433,N_6568,N_6610);
xor U8434 (N_8434,N_7189,N_6378);
or U8435 (N_8435,N_7094,N_7057);
or U8436 (N_8436,N_6617,N_7180);
nand U8437 (N_8437,N_7298,N_6953);
or U8438 (N_8438,N_6842,N_7362);
and U8439 (N_8439,N_7462,N_6570);
and U8440 (N_8440,N_6436,N_6005);
and U8441 (N_8441,N_6056,N_6306);
nand U8442 (N_8442,N_6986,N_6288);
nor U8443 (N_8443,N_6186,N_6183);
or U8444 (N_8444,N_7267,N_6496);
or U8445 (N_8445,N_6078,N_6245);
or U8446 (N_8446,N_6763,N_7233);
and U8447 (N_8447,N_6573,N_6289);
and U8448 (N_8448,N_6021,N_7379);
xor U8449 (N_8449,N_7269,N_7374);
xor U8450 (N_8450,N_6533,N_7143);
xor U8451 (N_8451,N_7046,N_6989);
nand U8452 (N_8452,N_7098,N_6718);
nand U8453 (N_8453,N_6708,N_6959);
xor U8454 (N_8454,N_7398,N_6312);
nor U8455 (N_8455,N_7125,N_6048);
xnor U8456 (N_8456,N_6654,N_6642);
xnor U8457 (N_8457,N_6186,N_7339);
nand U8458 (N_8458,N_6861,N_6378);
nor U8459 (N_8459,N_6545,N_6523);
and U8460 (N_8460,N_7120,N_7387);
nor U8461 (N_8461,N_6646,N_6650);
and U8462 (N_8462,N_6505,N_6579);
nand U8463 (N_8463,N_6962,N_6670);
nand U8464 (N_8464,N_7081,N_7198);
nor U8465 (N_8465,N_6285,N_6612);
or U8466 (N_8466,N_6771,N_6919);
xnor U8467 (N_8467,N_7298,N_6036);
nor U8468 (N_8468,N_6267,N_6628);
or U8469 (N_8469,N_6857,N_6402);
nor U8470 (N_8470,N_6216,N_6029);
and U8471 (N_8471,N_6770,N_6915);
and U8472 (N_8472,N_7156,N_6020);
and U8473 (N_8473,N_6991,N_6228);
or U8474 (N_8474,N_7094,N_6024);
xnor U8475 (N_8475,N_6074,N_6020);
or U8476 (N_8476,N_6670,N_6748);
or U8477 (N_8477,N_6154,N_7294);
xor U8478 (N_8478,N_6424,N_7180);
nor U8479 (N_8479,N_6885,N_7315);
nand U8480 (N_8480,N_7186,N_6400);
nand U8481 (N_8481,N_7470,N_7284);
or U8482 (N_8482,N_6805,N_7455);
nand U8483 (N_8483,N_6822,N_7028);
or U8484 (N_8484,N_7398,N_6734);
nand U8485 (N_8485,N_6321,N_6587);
nand U8486 (N_8486,N_6214,N_6766);
xor U8487 (N_8487,N_6521,N_6653);
and U8488 (N_8488,N_6945,N_7359);
or U8489 (N_8489,N_7071,N_6247);
nand U8490 (N_8490,N_6911,N_6368);
nor U8491 (N_8491,N_7474,N_6679);
nand U8492 (N_8492,N_7412,N_7094);
xnor U8493 (N_8493,N_6025,N_7297);
and U8494 (N_8494,N_6373,N_6629);
or U8495 (N_8495,N_6763,N_6769);
or U8496 (N_8496,N_6097,N_7209);
xnor U8497 (N_8497,N_6871,N_7456);
and U8498 (N_8498,N_6387,N_7395);
nor U8499 (N_8499,N_7194,N_6459);
or U8500 (N_8500,N_6543,N_6936);
xnor U8501 (N_8501,N_6167,N_7008);
nand U8502 (N_8502,N_6449,N_7219);
xnor U8503 (N_8503,N_7341,N_7397);
and U8504 (N_8504,N_7294,N_7039);
or U8505 (N_8505,N_6916,N_6020);
nor U8506 (N_8506,N_7486,N_6395);
nor U8507 (N_8507,N_6580,N_6786);
nand U8508 (N_8508,N_6301,N_6822);
nand U8509 (N_8509,N_6268,N_6475);
and U8510 (N_8510,N_6354,N_7194);
nand U8511 (N_8511,N_7408,N_6247);
or U8512 (N_8512,N_7352,N_6659);
and U8513 (N_8513,N_7022,N_6426);
nor U8514 (N_8514,N_7329,N_6724);
or U8515 (N_8515,N_6732,N_6273);
xnor U8516 (N_8516,N_6656,N_6412);
nand U8517 (N_8517,N_6804,N_6219);
nand U8518 (N_8518,N_7414,N_6685);
or U8519 (N_8519,N_6731,N_7328);
nand U8520 (N_8520,N_7415,N_6118);
and U8521 (N_8521,N_7219,N_6523);
xor U8522 (N_8522,N_6612,N_6078);
xor U8523 (N_8523,N_6941,N_6339);
or U8524 (N_8524,N_6850,N_6866);
nor U8525 (N_8525,N_6787,N_6427);
xnor U8526 (N_8526,N_6412,N_6788);
and U8527 (N_8527,N_6664,N_6824);
or U8528 (N_8528,N_6944,N_6304);
nor U8529 (N_8529,N_6376,N_7262);
xnor U8530 (N_8530,N_6277,N_6823);
xnor U8531 (N_8531,N_7171,N_6593);
nand U8532 (N_8532,N_7031,N_6221);
xor U8533 (N_8533,N_7075,N_7271);
and U8534 (N_8534,N_6683,N_6692);
or U8535 (N_8535,N_7066,N_6692);
nor U8536 (N_8536,N_6886,N_7211);
nor U8537 (N_8537,N_6296,N_7262);
or U8538 (N_8538,N_6871,N_7023);
nor U8539 (N_8539,N_6712,N_6386);
nand U8540 (N_8540,N_6199,N_6685);
xnor U8541 (N_8541,N_6078,N_6485);
nor U8542 (N_8542,N_6153,N_6207);
or U8543 (N_8543,N_7481,N_6920);
xor U8544 (N_8544,N_6477,N_6612);
nand U8545 (N_8545,N_6596,N_6349);
nand U8546 (N_8546,N_6467,N_6740);
xnor U8547 (N_8547,N_6884,N_7482);
or U8548 (N_8548,N_7456,N_6135);
nand U8549 (N_8549,N_6645,N_6013);
nand U8550 (N_8550,N_6620,N_7435);
nand U8551 (N_8551,N_6996,N_6875);
nor U8552 (N_8552,N_6200,N_7190);
and U8553 (N_8553,N_6865,N_6747);
and U8554 (N_8554,N_6414,N_6506);
nor U8555 (N_8555,N_6144,N_6021);
and U8556 (N_8556,N_6869,N_7430);
xor U8557 (N_8557,N_6462,N_6945);
nor U8558 (N_8558,N_6280,N_6453);
or U8559 (N_8559,N_6682,N_6736);
nor U8560 (N_8560,N_7360,N_6279);
or U8561 (N_8561,N_6248,N_7008);
and U8562 (N_8562,N_6097,N_6459);
xnor U8563 (N_8563,N_7348,N_6239);
or U8564 (N_8564,N_6045,N_6618);
xnor U8565 (N_8565,N_6427,N_6629);
xor U8566 (N_8566,N_7378,N_7260);
nor U8567 (N_8567,N_6971,N_7409);
xnor U8568 (N_8568,N_7015,N_6132);
nor U8569 (N_8569,N_7339,N_7468);
xnor U8570 (N_8570,N_6734,N_7090);
xnor U8571 (N_8571,N_6148,N_6723);
and U8572 (N_8572,N_6452,N_7367);
xnor U8573 (N_8573,N_6236,N_6110);
nor U8574 (N_8574,N_7413,N_7221);
and U8575 (N_8575,N_6850,N_6951);
and U8576 (N_8576,N_6131,N_7297);
and U8577 (N_8577,N_6570,N_6212);
xnor U8578 (N_8578,N_6117,N_7436);
nand U8579 (N_8579,N_7283,N_6340);
nand U8580 (N_8580,N_6251,N_7443);
and U8581 (N_8581,N_7464,N_6525);
or U8582 (N_8582,N_6044,N_7448);
nand U8583 (N_8583,N_6557,N_6352);
xnor U8584 (N_8584,N_7388,N_7381);
and U8585 (N_8585,N_7301,N_6870);
nand U8586 (N_8586,N_6537,N_6889);
and U8587 (N_8587,N_7075,N_6595);
nand U8588 (N_8588,N_6993,N_6639);
or U8589 (N_8589,N_6544,N_7088);
nor U8590 (N_8590,N_6583,N_6559);
nor U8591 (N_8591,N_7068,N_6165);
or U8592 (N_8592,N_6850,N_6013);
nand U8593 (N_8593,N_6840,N_6043);
and U8594 (N_8594,N_6497,N_7319);
and U8595 (N_8595,N_6677,N_7277);
nand U8596 (N_8596,N_6713,N_6555);
xor U8597 (N_8597,N_6367,N_6844);
or U8598 (N_8598,N_6200,N_6604);
or U8599 (N_8599,N_6209,N_6930);
and U8600 (N_8600,N_6670,N_6486);
xor U8601 (N_8601,N_6403,N_6617);
and U8602 (N_8602,N_6535,N_6938);
nand U8603 (N_8603,N_6695,N_7316);
nor U8604 (N_8604,N_7111,N_6700);
xnor U8605 (N_8605,N_6030,N_6591);
nor U8606 (N_8606,N_6417,N_7041);
nor U8607 (N_8607,N_6336,N_7372);
and U8608 (N_8608,N_6499,N_7320);
xnor U8609 (N_8609,N_6232,N_6450);
or U8610 (N_8610,N_7466,N_6670);
xor U8611 (N_8611,N_7294,N_7385);
nand U8612 (N_8612,N_6145,N_6134);
or U8613 (N_8613,N_6462,N_7001);
nor U8614 (N_8614,N_6042,N_6607);
nor U8615 (N_8615,N_6034,N_7441);
nor U8616 (N_8616,N_6214,N_6123);
and U8617 (N_8617,N_6465,N_6057);
nand U8618 (N_8618,N_6842,N_7034);
nor U8619 (N_8619,N_6048,N_6560);
nand U8620 (N_8620,N_6072,N_6463);
and U8621 (N_8621,N_6602,N_6594);
nor U8622 (N_8622,N_7061,N_6324);
or U8623 (N_8623,N_6482,N_6649);
xnor U8624 (N_8624,N_6317,N_7050);
and U8625 (N_8625,N_6953,N_6380);
nand U8626 (N_8626,N_6099,N_6344);
and U8627 (N_8627,N_6114,N_6386);
nor U8628 (N_8628,N_7189,N_6485);
nand U8629 (N_8629,N_6572,N_6538);
nor U8630 (N_8630,N_6569,N_6283);
and U8631 (N_8631,N_6387,N_6307);
xor U8632 (N_8632,N_6685,N_6837);
and U8633 (N_8633,N_7127,N_6639);
or U8634 (N_8634,N_6985,N_6662);
nor U8635 (N_8635,N_6225,N_7298);
nand U8636 (N_8636,N_6868,N_6452);
or U8637 (N_8637,N_7164,N_6239);
nor U8638 (N_8638,N_6970,N_7349);
xor U8639 (N_8639,N_6219,N_6404);
xnor U8640 (N_8640,N_6731,N_6361);
or U8641 (N_8641,N_6340,N_7373);
or U8642 (N_8642,N_6417,N_6498);
or U8643 (N_8643,N_7485,N_7154);
xnor U8644 (N_8644,N_7124,N_7375);
and U8645 (N_8645,N_6062,N_6837);
nor U8646 (N_8646,N_7040,N_6201);
nand U8647 (N_8647,N_6551,N_7420);
nor U8648 (N_8648,N_7294,N_6692);
and U8649 (N_8649,N_6373,N_7428);
nand U8650 (N_8650,N_7195,N_6637);
nor U8651 (N_8651,N_7433,N_6314);
or U8652 (N_8652,N_6048,N_7124);
nor U8653 (N_8653,N_6099,N_6985);
or U8654 (N_8654,N_6630,N_6307);
nor U8655 (N_8655,N_6525,N_7257);
nand U8656 (N_8656,N_6767,N_6828);
nor U8657 (N_8657,N_6264,N_7064);
or U8658 (N_8658,N_6572,N_6523);
and U8659 (N_8659,N_6390,N_6763);
nor U8660 (N_8660,N_7446,N_6737);
nand U8661 (N_8661,N_6152,N_6315);
or U8662 (N_8662,N_6037,N_6124);
and U8663 (N_8663,N_6957,N_6354);
or U8664 (N_8664,N_6737,N_7084);
or U8665 (N_8665,N_7301,N_7453);
xor U8666 (N_8666,N_6652,N_6529);
and U8667 (N_8667,N_6287,N_6607);
nand U8668 (N_8668,N_6096,N_6940);
and U8669 (N_8669,N_6987,N_6874);
xnor U8670 (N_8670,N_6570,N_7410);
or U8671 (N_8671,N_6954,N_6348);
nor U8672 (N_8672,N_7393,N_7042);
or U8673 (N_8673,N_7177,N_7029);
nand U8674 (N_8674,N_6773,N_6660);
xor U8675 (N_8675,N_6284,N_6749);
xnor U8676 (N_8676,N_6450,N_6569);
nor U8677 (N_8677,N_6798,N_7329);
nor U8678 (N_8678,N_6322,N_6881);
nand U8679 (N_8679,N_6462,N_6259);
or U8680 (N_8680,N_6522,N_7317);
or U8681 (N_8681,N_6174,N_6805);
or U8682 (N_8682,N_6448,N_6360);
and U8683 (N_8683,N_7154,N_6829);
nor U8684 (N_8684,N_7113,N_7391);
and U8685 (N_8685,N_6564,N_7358);
and U8686 (N_8686,N_6790,N_6229);
nand U8687 (N_8687,N_6128,N_6297);
xor U8688 (N_8688,N_6136,N_6569);
nand U8689 (N_8689,N_6215,N_7448);
nor U8690 (N_8690,N_6431,N_7455);
or U8691 (N_8691,N_7227,N_6557);
nand U8692 (N_8692,N_6776,N_6765);
and U8693 (N_8693,N_6546,N_6199);
or U8694 (N_8694,N_7369,N_6298);
xnor U8695 (N_8695,N_7388,N_6241);
nand U8696 (N_8696,N_6819,N_6496);
or U8697 (N_8697,N_6398,N_6876);
nand U8698 (N_8698,N_7059,N_7255);
nor U8699 (N_8699,N_6611,N_6841);
xnor U8700 (N_8700,N_6808,N_6716);
or U8701 (N_8701,N_7219,N_7237);
xor U8702 (N_8702,N_6074,N_6149);
or U8703 (N_8703,N_6843,N_6721);
nor U8704 (N_8704,N_6409,N_7372);
or U8705 (N_8705,N_6235,N_6887);
nand U8706 (N_8706,N_6718,N_7007);
nand U8707 (N_8707,N_7328,N_6855);
and U8708 (N_8708,N_7080,N_7050);
and U8709 (N_8709,N_6162,N_7092);
and U8710 (N_8710,N_6957,N_6147);
xnor U8711 (N_8711,N_6477,N_6569);
xnor U8712 (N_8712,N_6408,N_6136);
and U8713 (N_8713,N_7167,N_6187);
nor U8714 (N_8714,N_6958,N_6421);
nand U8715 (N_8715,N_6857,N_6388);
nor U8716 (N_8716,N_7234,N_7114);
and U8717 (N_8717,N_7412,N_6577);
and U8718 (N_8718,N_7049,N_6697);
and U8719 (N_8719,N_6436,N_6674);
and U8720 (N_8720,N_6482,N_6030);
xnor U8721 (N_8721,N_6488,N_7014);
or U8722 (N_8722,N_6322,N_6733);
nor U8723 (N_8723,N_7400,N_6384);
or U8724 (N_8724,N_7102,N_6296);
nand U8725 (N_8725,N_6044,N_6262);
nor U8726 (N_8726,N_7350,N_6861);
or U8727 (N_8727,N_6721,N_6716);
and U8728 (N_8728,N_7470,N_6684);
nand U8729 (N_8729,N_6067,N_6276);
and U8730 (N_8730,N_6575,N_6324);
nand U8731 (N_8731,N_6449,N_7173);
nand U8732 (N_8732,N_7003,N_6765);
nand U8733 (N_8733,N_6585,N_6334);
nor U8734 (N_8734,N_7114,N_7092);
nor U8735 (N_8735,N_7289,N_7260);
nor U8736 (N_8736,N_6324,N_7212);
nand U8737 (N_8737,N_6493,N_6583);
and U8738 (N_8738,N_7288,N_6634);
nand U8739 (N_8739,N_7035,N_7063);
or U8740 (N_8740,N_7427,N_6686);
and U8741 (N_8741,N_6987,N_7282);
and U8742 (N_8742,N_6053,N_6639);
and U8743 (N_8743,N_7384,N_7374);
and U8744 (N_8744,N_6969,N_7496);
xor U8745 (N_8745,N_7113,N_6351);
or U8746 (N_8746,N_6295,N_6431);
nand U8747 (N_8747,N_6140,N_7092);
nor U8748 (N_8748,N_6429,N_6233);
nand U8749 (N_8749,N_6211,N_6473);
and U8750 (N_8750,N_7175,N_7148);
xnor U8751 (N_8751,N_7063,N_6598);
xnor U8752 (N_8752,N_6900,N_7453);
or U8753 (N_8753,N_6847,N_6206);
xnor U8754 (N_8754,N_6665,N_7124);
and U8755 (N_8755,N_6989,N_7408);
nor U8756 (N_8756,N_6765,N_6599);
xnor U8757 (N_8757,N_6625,N_6049);
and U8758 (N_8758,N_6092,N_6286);
and U8759 (N_8759,N_7412,N_6638);
or U8760 (N_8760,N_6654,N_6303);
nand U8761 (N_8761,N_7246,N_6447);
nand U8762 (N_8762,N_7308,N_6192);
or U8763 (N_8763,N_6564,N_6258);
nor U8764 (N_8764,N_6255,N_6749);
nor U8765 (N_8765,N_6005,N_6389);
nor U8766 (N_8766,N_7341,N_6065);
xor U8767 (N_8767,N_6795,N_6209);
xnor U8768 (N_8768,N_6841,N_6982);
and U8769 (N_8769,N_6396,N_7256);
and U8770 (N_8770,N_7099,N_7272);
nor U8771 (N_8771,N_7392,N_6215);
and U8772 (N_8772,N_7475,N_7222);
and U8773 (N_8773,N_7120,N_6180);
and U8774 (N_8774,N_6377,N_6056);
nand U8775 (N_8775,N_6921,N_7009);
nand U8776 (N_8776,N_6286,N_7047);
xnor U8777 (N_8777,N_6403,N_6401);
nand U8778 (N_8778,N_6534,N_6436);
xor U8779 (N_8779,N_7027,N_7360);
or U8780 (N_8780,N_6600,N_6262);
nor U8781 (N_8781,N_7362,N_6092);
nor U8782 (N_8782,N_6691,N_6234);
xor U8783 (N_8783,N_6234,N_7461);
nor U8784 (N_8784,N_6310,N_6895);
nand U8785 (N_8785,N_6609,N_7116);
or U8786 (N_8786,N_6401,N_7371);
or U8787 (N_8787,N_7200,N_6808);
nor U8788 (N_8788,N_7475,N_6037);
or U8789 (N_8789,N_7320,N_7271);
nand U8790 (N_8790,N_6945,N_6967);
and U8791 (N_8791,N_6276,N_6723);
nor U8792 (N_8792,N_7252,N_6041);
nand U8793 (N_8793,N_6457,N_6228);
nand U8794 (N_8794,N_7188,N_6591);
or U8795 (N_8795,N_6972,N_6801);
nor U8796 (N_8796,N_7226,N_6631);
nand U8797 (N_8797,N_6556,N_6258);
or U8798 (N_8798,N_6525,N_6106);
nor U8799 (N_8799,N_6698,N_6298);
and U8800 (N_8800,N_7371,N_6538);
nor U8801 (N_8801,N_7401,N_6338);
and U8802 (N_8802,N_7181,N_6715);
or U8803 (N_8803,N_6643,N_6261);
nor U8804 (N_8804,N_6520,N_6997);
nor U8805 (N_8805,N_6045,N_6674);
or U8806 (N_8806,N_6775,N_6366);
nor U8807 (N_8807,N_6602,N_6352);
and U8808 (N_8808,N_6192,N_7067);
xnor U8809 (N_8809,N_6123,N_7080);
or U8810 (N_8810,N_6378,N_6045);
or U8811 (N_8811,N_6529,N_7198);
xnor U8812 (N_8812,N_7421,N_7408);
and U8813 (N_8813,N_7105,N_6420);
nor U8814 (N_8814,N_6842,N_6819);
nor U8815 (N_8815,N_6437,N_6050);
and U8816 (N_8816,N_6022,N_6812);
nand U8817 (N_8817,N_6453,N_6018);
or U8818 (N_8818,N_6797,N_6518);
and U8819 (N_8819,N_7401,N_6966);
or U8820 (N_8820,N_6303,N_6905);
nor U8821 (N_8821,N_6551,N_7398);
nand U8822 (N_8822,N_6449,N_6502);
xnor U8823 (N_8823,N_7475,N_6749);
or U8824 (N_8824,N_6309,N_6957);
nor U8825 (N_8825,N_6116,N_6437);
and U8826 (N_8826,N_7027,N_6239);
nand U8827 (N_8827,N_7445,N_7247);
xor U8828 (N_8828,N_6582,N_7184);
nor U8829 (N_8829,N_7444,N_6532);
nand U8830 (N_8830,N_7450,N_6677);
nor U8831 (N_8831,N_6615,N_6972);
nand U8832 (N_8832,N_7002,N_7109);
or U8833 (N_8833,N_6929,N_6861);
or U8834 (N_8834,N_6939,N_6180);
and U8835 (N_8835,N_6650,N_6747);
nand U8836 (N_8836,N_7343,N_6185);
nor U8837 (N_8837,N_7097,N_6747);
or U8838 (N_8838,N_7401,N_7115);
and U8839 (N_8839,N_6788,N_6304);
or U8840 (N_8840,N_6259,N_6330);
xor U8841 (N_8841,N_7480,N_6930);
xor U8842 (N_8842,N_6333,N_6224);
nand U8843 (N_8843,N_6464,N_7266);
nand U8844 (N_8844,N_6772,N_6818);
xnor U8845 (N_8845,N_7100,N_6990);
and U8846 (N_8846,N_7156,N_6068);
xor U8847 (N_8847,N_6352,N_7453);
or U8848 (N_8848,N_6327,N_7025);
and U8849 (N_8849,N_6315,N_6188);
and U8850 (N_8850,N_7224,N_6002);
nor U8851 (N_8851,N_6620,N_7384);
xnor U8852 (N_8852,N_6961,N_6227);
and U8853 (N_8853,N_6637,N_6510);
or U8854 (N_8854,N_6184,N_7403);
or U8855 (N_8855,N_7094,N_6663);
xnor U8856 (N_8856,N_6083,N_7152);
or U8857 (N_8857,N_6404,N_6003);
nor U8858 (N_8858,N_6268,N_6307);
or U8859 (N_8859,N_7240,N_7321);
xnor U8860 (N_8860,N_6264,N_6411);
and U8861 (N_8861,N_6770,N_6731);
or U8862 (N_8862,N_6702,N_6634);
xnor U8863 (N_8863,N_6929,N_7058);
nand U8864 (N_8864,N_6220,N_7228);
nand U8865 (N_8865,N_7368,N_6135);
or U8866 (N_8866,N_7164,N_7463);
nor U8867 (N_8867,N_6035,N_6572);
nand U8868 (N_8868,N_6796,N_6518);
and U8869 (N_8869,N_6042,N_6489);
or U8870 (N_8870,N_7288,N_6171);
nor U8871 (N_8871,N_7488,N_6809);
xor U8872 (N_8872,N_6583,N_6042);
and U8873 (N_8873,N_7309,N_6332);
nand U8874 (N_8874,N_6060,N_6197);
xnor U8875 (N_8875,N_6161,N_6199);
or U8876 (N_8876,N_6089,N_6399);
nor U8877 (N_8877,N_6920,N_6077);
or U8878 (N_8878,N_6929,N_6732);
xnor U8879 (N_8879,N_7140,N_6560);
xor U8880 (N_8880,N_7293,N_7046);
nor U8881 (N_8881,N_6162,N_7052);
nor U8882 (N_8882,N_7345,N_6254);
nor U8883 (N_8883,N_7175,N_6434);
or U8884 (N_8884,N_7191,N_6576);
nor U8885 (N_8885,N_7215,N_7092);
and U8886 (N_8886,N_6404,N_6208);
nor U8887 (N_8887,N_6238,N_7496);
xor U8888 (N_8888,N_6996,N_6575);
xnor U8889 (N_8889,N_6757,N_7229);
nand U8890 (N_8890,N_6506,N_7160);
nand U8891 (N_8891,N_7005,N_6563);
nand U8892 (N_8892,N_6998,N_7370);
and U8893 (N_8893,N_7343,N_6362);
xor U8894 (N_8894,N_6659,N_6737);
or U8895 (N_8895,N_7120,N_6984);
or U8896 (N_8896,N_7395,N_6186);
and U8897 (N_8897,N_6107,N_6902);
or U8898 (N_8898,N_6854,N_6445);
xnor U8899 (N_8899,N_6475,N_6266);
nand U8900 (N_8900,N_7474,N_6060);
and U8901 (N_8901,N_7066,N_7356);
and U8902 (N_8902,N_6091,N_7315);
xor U8903 (N_8903,N_6786,N_6599);
xnor U8904 (N_8904,N_7166,N_6471);
or U8905 (N_8905,N_6263,N_6685);
xor U8906 (N_8906,N_6635,N_7308);
or U8907 (N_8907,N_7172,N_6967);
and U8908 (N_8908,N_6855,N_6351);
and U8909 (N_8909,N_6476,N_6090);
nand U8910 (N_8910,N_7427,N_6889);
nand U8911 (N_8911,N_7047,N_6214);
nor U8912 (N_8912,N_6921,N_6070);
xnor U8913 (N_8913,N_7256,N_7429);
nand U8914 (N_8914,N_6348,N_7395);
or U8915 (N_8915,N_6643,N_6801);
nand U8916 (N_8916,N_6892,N_6466);
or U8917 (N_8917,N_6162,N_7182);
and U8918 (N_8918,N_6434,N_6878);
nand U8919 (N_8919,N_6788,N_6229);
and U8920 (N_8920,N_6206,N_6175);
nand U8921 (N_8921,N_6570,N_7371);
xnor U8922 (N_8922,N_6894,N_6785);
nor U8923 (N_8923,N_6616,N_7281);
nand U8924 (N_8924,N_6074,N_6814);
or U8925 (N_8925,N_6940,N_6479);
or U8926 (N_8926,N_6811,N_6809);
or U8927 (N_8927,N_6413,N_6336);
and U8928 (N_8928,N_7305,N_6551);
xnor U8929 (N_8929,N_7148,N_6958);
xnor U8930 (N_8930,N_7093,N_6318);
xor U8931 (N_8931,N_6479,N_7174);
xnor U8932 (N_8932,N_7370,N_7037);
nor U8933 (N_8933,N_7476,N_7475);
or U8934 (N_8934,N_7180,N_7200);
or U8935 (N_8935,N_6407,N_6216);
nor U8936 (N_8936,N_6454,N_6449);
or U8937 (N_8937,N_6434,N_7467);
nor U8938 (N_8938,N_6444,N_7438);
nand U8939 (N_8939,N_7109,N_6225);
or U8940 (N_8940,N_7281,N_7228);
xor U8941 (N_8941,N_6392,N_7249);
nor U8942 (N_8942,N_7423,N_6006);
nor U8943 (N_8943,N_6410,N_6652);
or U8944 (N_8944,N_6413,N_6468);
xor U8945 (N_8945,N_7486,N_6216);
or U8946 (N_8946,N_7227,N_6551);
xnor U8947 (N_8947,N_7420,N_6822);
or U8948 (N_8948,N_7333,N_6938);
xnor U8949 (N_8949,N_7014,N_7389);
nand U8950 (N_8950,N_7129,N_7327);
and U8951 (N_8951,N_6700,N_7214);
xor U8952 (N_8952,N_6897,N_6216);
and U8953 (N_8953,N_6348,N_7074);
and U8954 (N_8954,N_6870,N_7165);
xor U8955 (N_8955,N_7200,N_6624);
and U8956 (N_8956,N_6334,N_6446);
xor U8957 (N_8957,N_7231,N_6749);
or U8958 (N_8958,N_6417,N_7491);
nor U8959 (N_8959,N_6077,N_6820);
and U8960 (N_8960,N_6981,N_6466);
xor U8961 (N_8961,N_6757,N_6349);
or U8962 (N_8962,N_7312,N_6685);
xor U8963 (N_8963,N_6349,N_6137);
or U8964 (N_8964,N_6062,N_7181);
xnor U8965 (N_8965,N_6793,N_6554);
nor U8966 (N_8966,N_6890,N_6459);
nand U8967 (N_8967,N_6954,N_6037);
or U8968 (N_8968,N_6167,N_6807);
or U8969 (N_8969,N_6508,N_6142);
nand U8970 (N_8970,N_7228,N_7381);
or U8971 (N_8971,N_6837,N_6652);
nor U8972 (N_8972,N_7411,N_6500);
or U8973 (N_8973,N_7127,N_7105);
xnor U8974 (N_8974,N_6247,N_6725);
and U8975 (N_8975,N_6959,N_7098);
nand U8976 (N_8976,N_7115,N_6144);
and U8977 (N_8977,N_6186,N_6397);
or U8978 (N_8978,N_6080,N_6467);
or U8979 (N_8979,N_7137,N_6248);
and U8980 (N_8980,N_6750,N_6946);
and U8981 (N_8981,N_6273,N_6280);
nor U8982 (N_8982,N_6207,N_7224);
or U8983 (N_8983,N_7486,N_7481);
nor U8984 (N_8984,N_6293,N_6059);
and U8985 (N_8985,N_6115,N_6231);
and U8986 (N_8986,N_7097,N_6828);
and U8987 (N_8987,N_7049,N_6033);
and U8988 (N_8988,N_6128,N_6046);
nand U8989 (N_8989,N_6118,N_7058);
or U8990 (N_8990,N_7014,N_6950);
nand U8991 (N_8991,N_7404,N_6221);
xor U8992 (N_8992,N_7156,N_6359);
xor U8993 (N_8993,N_6157,N_6979);
or U8994 (N_8994,N_6560,N_7182);
or U8995 (N_8995,N_7191,N_7450);
or U8996 (N_8996,N_6896,N_6377);
and U8997 (N_8997,N_6646,N_7459);
and U8998 (N_8998,N_6454,N_6300);
and U8999 (N_8999,N_6186,N_6706);
xnor U9000 (N_9000,N_8184,N_8301);
nand U9001 (N_9001,N_8501,N_8669);
nand U9002 (N_9002,N_8633,N_7653);
nand U9003 (N_9003,N_8744,N_8917);
or U9004 (N_9004,N_7582,N_7883);
or U9005 (N_9005,N_8262,N_8174);
and U9006 (N_9006,N_7696,N_8728);
nor U9007 (N_9007,N_7766,N_8791);
nor U9008 (N_9008,N_7570,N_8990);
xnor U9009 (N_9009,N_8467,N_8764);
nor U9010 (N_9010,N_8115,N_8182);
xnor U9011 (N_9011,N_8930,N_8891);
nand U9012 (N_9012,N_7658,N_7809);
nor U9013 (N_9013,N_8879,N_8040);
xnor U9014 (N_9014,N_8581,N_7567);
nand U9015 (N_9015,N_8660,N_8529);
or U9016 (N_9016,N_8640,N_8574);
or U9017 (N_9017,N_7907,N_8083);
xor U9018 (N_9018,N_7845,N_8114);
and U9019 (N_9019,N_8927,N_7690);
and U9020 (N_9020,N_7751,N_7675);
nand U9021 (N_9021,N_8779,N_8484);
xnor U9022 (N_9022,N_8796,N_8761);
nor U9023 (N_9023,N_7948,N_8307);
and U9024 (N_9024,N_7531,N_7600);
nand U9025 (N_9025,N_7754,N_8429);
nor U9026 (N_9026,N_8547,N_7572);
or U9027 (N_9027,N_8552,N_8940);
nand U9028 (N_9028,N_8588,N_8492);
and U9029 (N_9029,N_8831,N_7862);
nor U9030 (N_9030,N_8934,N_7958);
xnor U9031 (N_9031,N_8306,N_8226);
nor U9032 (N_9032,N_8131,N_8849);
and U9033 (N_9033,N_8192,N_8625);
xnor U9034 (N_9034,N_8185,N_8896);
xnor U9035 (N_9035,N_8228,N_7872);
or U9036 (N_9036,N_7668,N_8903);
xor U9037 (N_9037,N_7821,N_7681);
nand U9038 (N_9038,N_7991,N_7786);
and U9039 (N_9039,N_8460,N_8388);
nand U9040 (N_9040,N_8027,N_8159);
and U9041 (N_9041,N_8942,N_8936);
nand U9042 (N_9042,N_7526,N_8980);
and U9043 (N_9043,N_7566,N_8537);
nor U9044 (N_9044,N_8026,N_8736);
and U9045 (N_9045,N_7993,N_8399);
or U9046 (N_9046,N_8546,N_7753);
nand U9047 (N_9047,N_7741,N_8740);
nand U9048 (N_9048,N_8878,N_8496);
and U9049 (N_9049,N_8289,N_8005);
nand U9050 (N_9050,N_7599,N_8441);
or U9051 (N_9051,N_7995,N_8569);
or U9052 (N_9052,N_8583,N_8048);
nand U9053 (N_9053,N_7825,N_8682);
xnor U9054 (N_9054,N_7933,N_7711);
xor U9055 (N_9055,N_8366,N_7530);
xor U9056 (N_9056,N_7693,N_8885);
nor U9057 (N_9057,N_8287,N_7647);
nand U9058 (N_9058,N_7501,N_8834);
nor U9059 (N_9059,N_8420,N_8915);
xnor U9060 (N_9060,N_8679,N_8476);
or U9061 (N_9061,N_8424,N_8756);
nor U9062 (N_9062,N_8911,N_7971);
nor U9063 (N_9063,N_7774,N_8607);
nor U9064 (N_9064,N_7619,N_8926);
xor U9065 (N_9065,N_7922,N_7866);
or U9066 (N_9066,N_7554,N_7822);
and U9067 (N_9067,N_8909,N_8272);
and U9068 (N_9068,N_8076,N_8527);
nand U9069 (N_9069,N_8630,N_8737);
xnor U9070 (N_9070,N_8579,N_8517);
or U9071 (N_9071,N_7855,N_8385);
nor U9072 (N_9072,N_8555,N_8269);
nand U9073 (N_9073,N_8983,N_7801);
xnor U9074 (N_9074,N_8683,N_8402);
xor U9075 (N_9075,N_7630,N_8644);
or U9076 (N_9076,N_8642,N_8599);
nor U9077 (N_9077,N_8187,N_8266);
and U9078 (N_9078,N_8075,N_8271);
and U9079 (N_9079,N_8726,N_8818);
xor U9080 (N_9080,N_8895,N_8912);
nor U9081 (N_9081,N_8168,N_8037);
xor U9082 (N_9082,N_8098,N_8541);
xor U9083 (N_9083,N_8512,N_7757);
nor U9084 (N_9084,N_8299,N_8322);
or U9085 (N_9085,N_8809,N_8015);
and U9086 (N_9086,N_7574,N_8246);
xor U9087 (N_9087,N_8994,N_8274);
xor U9088 (N_9088,N_8065,N_7882);
and U9089 (N_9089,N_7601,N_8982);
nor U9090 (N_9090,N_7939,N_7556);
or U9091 (N_9091,N_7695,N_7520);
or U9092 (N_9092,N_7587,N_8802);
or U9093 (N_9093,N_7729,N_7833);
and U9094 (N_9094,N_7738,N_8386);
xor U9095 (N_9095,N_8584,N_7789);
xor U9096 (N_9096,N_8924,N_8945);
and U9097 (N_9097,N_7942,N_7542);
nor U9098 (N_9098,N_8444,N_7854);
and U9099 (N_9099,N_7873,N_7655);
or U9100 (N_9100,N_7674,N_7981);
nor U9101 (N_9101,N_8550,N_8433);
nand U9102 (N_9102,N_7899,N_8178);
nand U9103 (N_9103,N_7591,N_7876);
and U9104 (N_9104,N_7955,N_7585);
xnor U9105 (N_9105,N_8752,N_8066);
nor U9106 (N_9106,N_8361,N_7692);
nand U9107 (N_9107,N_8454,N_8795);
or U9108 (N_9108,N_8353,N_8523);
and U9109 (N_9109,N_8247,N_7747);
or U9110 (N_9110,N_8920,N_8419);
nand U9111 (N_9111,N_8524,N_8698);
xnor U9112 (N_9112,N_7590,N_8916);
and U9113 (N_9113,N_8975,N_8499);
or U9114 (N_9114,N_7843,N_8296);
xnor U9115 (N_9115,N_8031,N_8163);
xor U9116 (N_9116,N_8145,N_7549);
xnor U9117 (N_9117,N_7637,N_8064);
nand U9118 (N_9118,N_8594,N_8350);
or U9119 (N_9119,N_8151,N_8913);
nor U9120 (N_9120,N_8807,N_7671);
nor U9121 (N_9121,N_7588,N_8827);
nor U9122 (N_9122,N_7764,N_8876);
or U9123 (N_9123,N_8459,N_7778);
and U9124 (N_9124,N_7967,N_8883);
nand U9125 (N_9125,N_8097,N_8355);
xnor U9126 (N_9126,N_8403,N_8021);
nand U9127 (N_9127,N_8149,N_8691);
xnor U9128 (N_9128,N_8381,N_8848);
and U9129 (N_9129,N_8465,N_8073);
nor U9130 (N_9130,N_7553,N_7635);
nor U9131 (N_9131,N_8582,N_8139);
xnor U9132 (N_9132,N_8856,N_7787);
or U9133 (N_9133,N_7578,N_7652);
nor U9134 (N_9134,N_8252,N_8566);
or U9135 (N_9135,N_8999,N_8578);
and U9136 (N_9136,N_8238,N_8536);
xnor U9137 (N_9137,N_8970,N_8223);
nor U9138 (N_9138,N_8641,N_7663);
or U9139 (N_9139,N_8820,N_8201);
and U9140 (N_9140,N_8119,N_8839);
and U9141 (N_9141,N_8088,N_8416);
nor U9142 (N_9142,N_7612,N_8789);
xnor U9143 (N_9143,N_8199,N_7594);
xor U9144 (N_9144,N_7800,N_7932);
xor U9145 (N_9145,N_8910,N_7505);
nor U9146 (N_9146,N_8870,N_8564);
xnor U9147 (N_9147,N_7592,N_8525);
and U9148 (N_9148,N_7765,N_8413);
nor U9149 (N_9149,N_7889,N_7654);
nor U9150 (N_9150,N_7563,N_8535);
nand U9151 (N_9151,N_7888,N_7506);
or U9152 (N_9152,N_8998,N_7768);
or U9153 (N_9153,N_7545,N_7557);
nand U9154 (N_9154,N_8367,N_7755);
nor U9155 (N_9155,N_7529,N_8814);
and U9156 (N_9156,N_8610,N_8605);
nand U9157 (N_9157,N_8471,N_8260);
or U9158 (N_9158,N_8346,N_7909);
or U9159 (N_9159,N_8613,N_8464);
xnor U9160 (N_9160,N_8935,N_7519);
xnor U9161 (N_9161,N_7508,N_8632);
nor U9162 (N_9162,N_8696,N_8657);
xnor U9163 (N_9163,N_8225,N_7734);
nor U9164 (N_9164,N_8030,N_7963);
or U9165 (N_9165,N_8276,N_8964);
nand U9166 (N_9166,N_8977,N_7914);
and U9167 (N_9167,N_8906,N_8662);
xnor U9168 (N_9168,N_8611,N_7871);
and U9169 (N_9169,N_7807,N_8699);
xor U9170 (N_9170,N_8538,N_8019);
and U9171 (N_9171,N_8677,N_8823);
or U9172 (N_9172,N_8253,N_7941);
nor U9173 (N_9173,N_8079,N_7790);
nor U9174 (N_9174,N_8622,N_8943);
xnor U9175 (N_9175,N_8111,N_7752);
nor U9176 (N_9176,N_8825,N_8816);
nor U9177 (N_9177,N_7987,N_7636);
xor U9178 (N_9178,N_8035,N_8741);
or U9179 (N_9179,N_8319,N_8714);
or U9180 (N_9180,N_8323,N_8109);
nand U9181 (N_9181,N_8860,N_7742);
xnor U9182 (N_9182,N_7921,N_8635);
nor U9183 (N_9183,N_8077,N_8855);
and U9184 (N_9184,N_8370,N_8798);
nand U9185 (N_9185,N_7935,N_8559);
and U9186 (N_9186,N_7705,N_8297);
or U9187 (N_9187,N_8093,N_8136);
xnor U9188 (N_9188,N_8422,N_8781);
nand U9189 (N_9189,N_7965,N_7975);
nand U9190 (N_9190,N_7723,N_8347);
and U9191 (N_9191,N_7969,N_8655);
or U9192 (N_9192,N_8376,N_8001);
xor U9193 (N_9193,N_8283,N_7950);
or U9194 (N_9194,N_7890,N_8576);
nor U9195 (N_9195,N_8522,N_8689);
nand U9196 (N_9196,N_7504,N_8939);
xnor U9197 (N_9197,N_8750,N_8061);
nand U9198 (N_9198,N_8869,N_8428);
or U9199 (N_9199,N_7885,N_8058);
xnor U9200 (N_9200,N_7928,N_8591);
nand U9201 (N_9201,N_7806,N_8830);
and U9202 (N_9202,N_8208,N_8009);
xor U9203 (N_9203,N_8013,N_7606);
and U9204 (N_9204,N_8749,N_8585);
nor U9205 (N_9205,N_8776,N_7595);
nand U9206 (N_9206,N_7852,N_8273);
xnor U9207 (N_9207,N_8162,N_8688);
nor U9208 (N_9208,N_8971,N_7829);
xnor U9209 (N_9209,N_7886,N_8380);
and U9210 (N_9210,N_8294,N_7811);
and U9211 (N_9211,N_8447,N_8084);
nor U9212 (N_9212,N_8236,N_7929);
and U9213 (N_9213,N_7988,N_8561);
xnor U9214 (N_9214,N_8440,N_8286);
nand U9215 (N_9215,N_8356,N_8684);
nor U9216 (N_9216,N_8067,N_8049);
and U9217 (N_9217,N_8745,N_8120);
or U9218 (N_9218,N_8601,N_7500);
and U9219 (N_9219,N_8117,N_7547);
or U9220 (N_9220,N_7716,N_8325);
and U9221 (N_9221,N_8494,N_8375);
xor U9222 (N_9222,N_8626,N_8722);
nor U9223 (N_9223,N_8110,N_8743);
and U9224 (N_9224,N_7713,N_8693);
xnor U9225 (N_9225,N_8104,N_8063);
xnor U9226 (N_9226,N_7569,N_8106);
nand U9227 (N_9227,N_8957,N_7731);
and U9228 (N_9228,N_7999,N_7536);
and U9229 (N_9229,N_8121,N_8933);
or U9230 (N_9230,N_7736,N_8025);
nor U9231 (N_9231,N_8897,N_8706);
and U9232 (N_9232,N_8553,N_8060);
xor U9233 (N_9233,N_7634,N_8557);
nor U9234 (N_9234,N_7979,N_8062);
nor U9235 (N_9235,N_8974,N_8202);
xor U9236 (N_9236,N_8495,N_8995);
nor U9237 (N_9237,N_8604,N_7552);
xor U9238 (N_9238,N_8071,N_7620);
xnor U9239 (N_9239,N_8087,N_8290);
or U9240 (N_9240,N_8560,N_8503);
xnor U9241 (N_9241,N_8739,N_7511);
nor U9242 (N_9242,N_8291,N_8214);
nand U9243 (N_9243,N_7537,N_7830);
and U9244 (N_9244,N_8854,N_7947);
and U9245 (N_9245,N_7703,N_8141);
nor U9246 (N_9246,N_7953,N_8100);
xnor U9247 (N_9247,N_8360,N_8784);
or U9248 (N_9248,N_8221,N_8890);
nor U9249 (N_9249,N_7515,N_8603);
nand U9250 (N_9250,N_8409,N_7605);
xor U9251 (N_9251,N_8227,N_7761);
nand U9252 (N_9252,N_7678,N_8313);
or U9253 (N_9253,N_8300,N_8142);
and U9254 (N_9254,N_8656,N_7997);
nand U9255 (N_9255,N_8379,N_8080);
and U9256 (N_9256,N_8263,N_7721);
xnor U9257 (N_9257,N_8690,N_8183);
or U9258 (N_9258,N_8785,N_8858);
xnor U9259 (N_9259,N_8309,N_7616);
or U9260 (N_9260,N_8195,N_8851);
nor U9261 (N_9261,N_7524,N_7859);
nand U9262 (N_9262,N_7722,N_8445);
nor U9263 (N_9263,N_8256,N_8593);
nand U9264 (N_9264,N_7666,N_8123);
and U9265 (N_9265,N_8947,N_7824);
nand U9266 (N_9266,N_8658,N_7911);
xnor U9267 (N_9267,N_7715,N_7805);
or U9268 (N_9268,N_8480,N_7593);
nand U9269 (N_9269,N_7684,N_7804);
nor U9270 (N_9270,N_7864,N_7784);
or U9271 (N_9271,N_7608,N_8542);
xor U9272 (N_9272,N_7986,N_8664);
and U9273 (N_9273,N_8042,N_7857);
xor U9274 (N_9274,N_7930,N_7974);
or U9275 (N_9275,N_8623,N_8292);
and U9276 (N_9276,N_8639,N_7669);
nand U9277 (N_9277,N_8137,N_8008);
nand U9278 (N_9278,N_7740,N_7733);
xnor U9279 (N_9279,N_8710,N_8144);
or U9280 (N_9280,N_7743,N_7904);
xor U9281 (N_9281,N_7571,N_8616);
nand U9282 (N_9282,N_8963,N_8861);
and U9283 (N_9283,N_8932,N_8918);
or U9284 (N_9284,N_7628,N_8993);
xor U9285 (N_9285,N_8410,N_8996);
xor U9286 (N_9286,N_7580,N_8806);
nand U9287 (N_9287,N_8819,N_8308);
nor U9288 (N_9288,N_8986,N_7642);
and U9289 (N_9289,N_8738,N_8218);
xor U9290 (N_9290,N_8505,N_7699);
nand U9291 (N_9291,N_8427,N_7522);
nor U9292 (N_9292,N_8426,N_7614);
xnor U9293 (N_9293,N_8176,N_7584);
nand U9294 (N_9294,N_8485,N_8598);
nor U9295 (N_9295,N_8384,N_8050);
xor U9296 (N_9296,N_8398,N_7903);
or U9297 (N_9297,N_8654,N_7532);
or U9298 (N_9298,N_7686,N_7577);
nor U9299 (N_9299,N_8340,N_8196);
nor U9300 (N_9300,N_7788,N_8395);
xor U9301 (N_9301,N_8705,N_7610);
xnor U9302 (N_9302,N_8295,N_8328);
nand U9303 (N_9303,N_7701,N_8965);
xnor U9304 (N_9304,N_7648,N_7561);
xnor U9305 (N_9305,N_8742,N_8334);
xor U9306 (N_9306,N_7662,N_8242);
or U9307 (N_9307,N_8091,N_8374);
and U9308 (N_9308,N_8908,N_8258);
nand U9309 (N_9309,N_8359,N_8181);
nor U9310 (N_9310,N_8602,N_7836);
nor U9311 (N_9311,N_8280,N_7962);
or U9312 (N_9312,N_8680,N_8431);
xnor U9313 (N_9313,N_8217,N_8961);
nand U9314 (N_9314,N_7613,N_8797);
nor U9315 (N_9315,N_7850,N_7513);
nor U9316 (N_9316,N_7808,N_7989);
nand U9317 (N_9317,N_8003,N_7867);
and U9318 (N_9318,N_8674,N_8694);
nor U9319 (N_9319,N_8345,N_7672);
and U9320 (N_9320,N_8462,N_7860);
or U9321 (N_9321,N_8650,N_8069);
nand U9322 (N_9322,N_8944,N_8315);
nor U9323 (N_9323,N_8695,N_8866);
xor U9324 (N_9324,N_7603,N_8392);
or U9325 (N_9325,N_7920,N_8390);
or U9326 (N_9326,N_8824,N_8024);
xnor U9327 (N_9327,N_7802,N_8434);
nand U9328 (N_9328,N_8596,N_8755);
xnor U9329 (N_9329,N_8298,N_8383);
nand U9330 (N_9330,N_8777,N_7810);
xor U9331 (N_9331,N_7990,N_8249);
xnor U9332 (N_9332,N_7823,N_7937);
nand U9333 (N_9333,N_8277,N_8127);
or U9334 (N_9334,N_8634,N_7992);
xor U9335 (N_9335,N_7688,N_8767);
nand U9336 (N_9336,N_7670,N_7881);
nand U9337 (N_9337,N_8166,N_8719);
nor U9338 (N_9338,N_8748,N_8829);
nand U9339 (N_9339,N_7626,N_8017);
or U9340 (N_9340,N_8177,N_8082);
and U9341 (N_9341,N_7949,N_7803);
nand U9342 (N_9342,N_7739,N_7994);
xnor U9343 (N_9343,N_8946,N_7797);
nor U9344 (N_9344,N_7792,N_8889);
nand U9345 (N_9345,N_7523,N_8125);
nor U9346 (N_9346,N_8488,N_8438);
xnor U9347 (N_9347,N_8518,N_7762);
and U9348 (N_9348,N_7714,N_8101);
and U9349 (N_9349,N_8081,N_8222);
and U9350 (N_9350,N_7970,N_7581);
nand U9351 (N_9351,N_8700,N_7780);
nor U9352 (N_9352,N_8959,N_8255);
and U9353 (N_9353,N_7615,N_8051);
xor U9354 (N_9354,N_7717,N_8801);
nor U9355 (N_9355,N_7785,N_7913);
and U9356 (N_9356,N_8198,N_8880);
nor U9357 (N_9357,N_8257,N_8096);
nor U9358 (N_9358,N_8960,N_8703);
and U9359 (N_9359,N_8224,N_8620);
nor U9360 (N_9360,N_8671,N_8905);
nor U9361 (N_9361,N_8155,N_8780);
nand U9362 (N_9362,N_7848,N_8270);
nand U9363 (N_9363,N_8717,N_8378);
and U9364 (N_9364,N_8812,N_8165);
nand U9365 (N_9365,N_7502,N_7891);
nand U9366 (N_9366,N_8105,N_8868);
and U9367 (N_9367,N_8989,N_8790);
nand U9368 (N_9368,N_7934,N_7517);
xnor U9369 (N_9369,N_8676,N_8118);
xnor U9370 (N_9370,N_7812,N_8152);
and U9371 (N_9371,N_8489,N_7618);
nor U9372 (N_9372,N_8126,N_8898);
nand U9373 (N_9373,N_8483,N_7507);
nand U9374 (N_9374,N_7617,N_8925);
and U9375 (N_9375,N_7772,N_8955);
and U9376 (N_9376,N_8430,N_7641);
nand U9377 (N_9377,N_7957,N_8772);
xnor U9378 (N_9378,N_7781,N_8029);
and U9379 (N_9379,N_8432,N_8991);
or U9380 (N_9380,N_8043,N_7951);
or U9381 (N_9381,N_7814,N_8763);
xor U9382 (N_9382,N_8461,N_8245);
or U9383 (N_9383,N_8808,N_8609);
or U9384 (N_9384,N_7640,N_7827);
or U9385 (N_9385,N_8507,N_8044);
nor U9386 (N_9386,N_8330,N_8016);
and U9387 (N_9387,N_8000,N_8826);
xor U9388 (N_9388,N_8953,N_7573);
nor U9389 (N_9389,N_8979,N_8156);
nor U9390 (N_9390,N_8941,N_8759);
nor U9391 (N_9391,N_8362,N_8702);
xor U9392 (N_9392,N_8615,N_7707);
and U9393 (N_9393,N_7737,N_7777);
xor U9394 (N_9394,N_8161,N_7842);
and U9395 (N_9395,N_7983,N_8648);
xnor U9396 (N_9396,N_8614,N_8393);
nand U9397 (N_9397,N_8397,N_7835);
and U9398 (N_9398,N_7694,N_7844);
xnor U9399 (N_9399,N_8766,N_8194);
nand U9400 (N_9400,N_7831,N_7708);
nand U9401 (N_9401,N_8180,N_8968);
or U9402 (N_9402,N_8568,N_8173);
or U9403 (N_9403,N_8978,N_7858);
xor U9404 (N_9404,N_8544,N_7847);
nand U9405 (N_9405,N_7589,N_8608);
nor U9406 (N_9406,N_7576,N_8985);
xor U9407 (N_9407,N_8382,N_8701);
nand U9408 (N_9408,N_8768,N_8859);
nor U9409 (N_9409,N_8130,N_8487);
and U9410 (N_9410,N_8357,N_7894);
and U9411 (N_9411,N_8086,N_8264);
nor U9412 (N_9412,N_8665,N_8239);
and U9413 (N_9413,N_7541,N_8175);
or U9414 (N_9414,N_7925,N_8251);
and U9415 (N_9415,N_7945,N_8436);
nand U9416 (N_9416,N_7624,N_8725);
xnor U9417 (N_9417,N_8220,N_7575);
and U9418 (N_9418,N_8765,N_8113);
and U9419 (N_9419,N_7946,N_8365);
nand U9420 (N_9420,N_8022,N_7849);
or U9421 (N_9421,N_8753,N_8606);
nor U9422 (N_9422,N_8449,N_7880);
nand U9423 (N_9423,N_8627,N_8841);
nor U9424 (N_9424,N_8881,N_8311);
nand U9425 (N_9425,N_8129,N_7720);
or U9426 (N_9426,N_8810,N_7817);
xor U9427 (N_9427,N_7915,N_8046);
xor U9428 (N_9428,N_8059,N_7732);
nor U9429 (N_9429,N_7869,N_8099);
xor U9430 (N_9430,N_7689,N_8846);
and U9431 (N_9431,N_8884,N_8842);
or U9432 (N_9432,N_7667,N_8203);
xor U9433 (N_9433,N_8592,N_8519);
nand U9434 (N_9434,N_8533,N_7525);
nand U9435 (N_9435,N_8708,N_8850);
and U9436 (N_9436,N_8647,N_8036);
and U9437 (N_9437,N_7851,N_8548);
xnor U9438 (N_9438,N_7996,N_8888);
xnor U9439 (N_9439,N_7856,N_8733);
nand U9440 (N_9440,N_8754,N_7796);
and U9441 (N_9441,N_8976,N_8510);
nor U9442 (N_9442,N_8054,N_8469);
xor U9443 (N_9443,N_8646,N_8302);
xnor U9444 (N_9444,N_7902,N_8774);
and U9445 (N_9445,N_8233,N_8670);
nand U9446 (N_9446,N_7841,N_8709);
and U9447 (N_9447,N_8329,N_8278);
xor U9448 (N_9448,N_8805,N_8707);
and U9449 (N_9449,N_8659,N_8844);
and U9450 (N_9450,N_8211,N_7896);
and U9451 (N_9451,N_7727,N_7514);
xnor U9452 (N_9452,N_8692,N_7795);
or U9453 (N_9453,N_7656,N_8565);
or U9454 (N_9454,N_8443,N_7712);
and U9455 (N_9455,N_8800,N_7799);
nor U9456 (N_9456,N_8477,N_7709);
or U9457 (N_9457,N_8624,N_7539);
nand U9458 (N_9458,N_7770,N_7650);
or U9459 (N_9459,N_7638,N_8490);
nor U9460 (N_9460,N_8284,N_7621);
xor U9461 (N_9461,N_7535,N_8778);
xor U9462 (N_9462,N_8351,N_8103);
and U9463 (N_9463,N_7918,N_7968);
or U9464 (N_9464,N_7980,N_7878);
xnor U9465 (N_9465,N_8637,N_7657);
xor U9466 (N_9466,N_8268,N_8303);
nand U9467 (N_9467,N_8358,N_8919);
and U9468 (N_9468,N_8147,N_8992);
nor U9469 (N_9469,N_7917,N_8265);
or U9470 (N_9470,N_7730,N_8415);
and U9471 (N_9471,N_7927,N_8751);
and U9472 (N_9472,N_8951,N_8335);
and U9473 (N_9473,N_7728,N_7559);
xnor U9474 (N_9474,N_8463,N_7905);
and U9475 (N_9475,N_8852,N_8092);
nor U9476 (N_9476,N_8138,N_8718);
nand U9477 (N_9477,N_8108,N_8468);
xnor U9478 (N_9478,N_7673,N_7661);
or U9479 (N_9479,N_8562,N_8840);
nor U9480 (N_9480,N_7597,N_7565);
and U9481 (N_9481,N_8007,N_8275);
nor U9482 (N_9482,N_7538,N_8773);
and U9483 (N_9483,N_8716,N_8803);
nand U9484 (N_9484,N_7750,N_8686);
and U9485 (N_9485,N_7516,N_8572);
nor U9486 (N_9486,N_8972,N_8843);
xor U9487 (N_9487,N_8727,N_8526);
or U9488 (N_9488,N_7960,N_8886);
or U9489 (N_9489,N_8327,N_7697);
nor U9490 (N_9490,N_8954,N_8762);
xnor U9491 (N_9491,N_8681,N_8758);
or U9492 (N_9492,N_8244,N_8871);
and U9493 (N_9493,N_8653,N_8668);
nor U9494 (N_9494,N_8857,N_8377);
nor U9495 (N_9495,N_7875,N_7512);
nand U9496 (N_9496,N_7926,N_7916);
and U9497 (N_9497,N_7870,N_8023);
nand U9498 (N_9498,N_8206,N_8401);
and U9499 (N_9499,N_8408,N_8085);
and U9500 (N_9500,N_7791,N_8847);
nor U9501 (N_9501,N_8337,N_7893);
or U9502 (N_9502,N_8056,N_7644);
or U9503 (N_9503,N_7745,N_8451);
nor U9504 (N_9504,N_8645,N_8651);
or U9505 (N_9505,N_8528,N_8169);
nand U9506 (N_9506,N_7629,N_8811);
nor U9507 (N_9507,N_8874,N_8041);
or U9508 (N_9508,N_7651,N_8193);
nand U9509 (N_9509,N_7868,N_8864);
or U9510 (N_9510,N_8838,N_8473);
or U9511 (N_9511,N_8997,N_8216);
and U9512 (N_9512,N_8458,N_8219);
or U9513 (N_9513,N_8344,N_8332);
xor U9514 (N_9514,N_8070,N_8212);
nor U9515 (N_9515,N_8575,N_8534);
nor U9516 (N_9516,N_8405,N_8600);
xor U9517 (N_9517,N_8732,N_8783);
xor U9518 (N_9518,N_8312,N_7706);
nor U9519 (N_9519,N_8389,N_8835);
xnor U9520 (N_9520,N_8675,N_7956);
and U9521 (N_9521,N_7702,N_8729);
nor U9522 (N_9522,N_8241,N_8962);
nor U9523 (N_9523,N_8039,N_8958);
nor U9524 (N_9524,N_8179,N_8902);
and U9525 (N_9525,N_7982,N_7749);
nand U9526 (N_9526,N_8074,N_8837);
nor U9527 (N_9527,N_8904,N_8146);
xor U9528 (N_9528,N_8425,N_7865);
nor U9529 (N_9529,N_8190,N_8240);
or U9530 (N_9530,N_8414,N_7685);
and U9531 (N_9531,N_8004,N_7944);
xor U9532 (N_9532,N_8047,N_7704);
or U9533 (N_9533,N_8938,N_7892);
xor U9534 (N_9534,N_7551,N_8734);
nor U9535 (N_9535,N_7846,N_7767);
and U9536 (N_9536,N_8372,N_8229);
nand U9537 (N_9537,N_7639,N_7998);
and U9538 (N_9538,N_8304,N_8318);
nor U9539 (N_9539,N_7659,N_8479);
xnor U9540 (N_9540,N_8002,N_8186);
and U9541 (N_9541,N_8338,N_8988);
nand U9542 (N_9542,N_8140,N_7895);
nor U9543 (N_9543,N_7839,N_8636);
or U9544 (N_9544,N_8124,N_8164);
or U9545 (N_9545,N_8279,N_7583);
or U9546 (N_9546,N_8587,N_8929);
nand U9547 (N_9547,N_7884,N_7735);
xnor U9548 (N_9548,N_8072,N_8288);
nor U9549 (N_9549,N_8010,N_8466);
or U9550 (N_9550,N_7775,N_8987);
xnor U9551 (N_9551,N_7625,N_7609);
or U9552 (N_9552,N_8687,N_8554);
nor U9553 (N_9553,N_8478,N_7510);
nor U9554 (N_9554,N_8931,N_8508);
and U9555 (N_9555,N_8053,N_8981);
xor U9556 (N_9556,N_7645,N_8590);
or U9557 (N_9557,N_8793,N_7649);
nand U9558 (N_9558,N_8411,N_8713);
nor U9559 (N_9559,N_7973,N_8786);
xor U9560 (N_9560,N_8540,N_8556);
or U9561 (N_9561,N_8724,N_7923);
or U9562 (N_9562,N_8794,N_8769);
and U9563 (N_9563,N_8107,N_8364);
and U9564 (N_9564,N_8712,N_8324);
xor U9565 (N_9565,N_7760,N_8412);
and U9566 (N_9566,N_7664,N_8720);
and U9567 (N_9567,N_8207,N_8404);
and U9568 (N_9568,N_7840,N_8455);
xnor U9569 (N_9569,N_7598,N_8439);
xor U9570 (N_9570,N_8267,N_8899);
and U9571 (N_9571,N_8316,N_7794);
and U9572 (N_9572,N_7503,N_7548);
xor U9573 (N_9573,N_8135,N_8612);
nand U9574 (N_9574,N_8310,N_8493);
nand U9575 (N_9575,N_8617,N_8914);
or U9576 (N_9576,N_8514,N_8928);
nand U9577 (N_9577,N_7646,N_7748);
or U9578 (N_9578,N_8619,N_8014);
xor U9579 (N_9579,N_7682,N_7940);
xor U9580 (N_9580,N_7756,N_8573);
and U9581 (N_9581,N_8423,N_8200);
xor U9582 (N_9582,N_8937,N_8012);
xor U9583 (N_9583,N_7863,N_7725);
nor U9584 (N_9584,N_8354,N_8577);
xor U9585 (N_9585,N_8032,N_8813);
or U9586 (N_9586,N_7985,N_8667);
xor U9587 (N_9587,N_8452,N_7665);
nand U9588 (N_9588,N_7633,N_7710);
nand U9589 (N_9589,N_8363,N_8336);
and U9590 (N_9590,N_7769,N_7746);
or U9591 (N_9591,N_8775,N_7631);
nor U9592 (N_9592,N_7954,N_8629);
nand U9593 (N_9593,N_7680,N_7783);
nand U9594 (N_9594,N_8134,N_8730);
and U9595 (N_9595,N_8853,N_7782);
and U9596 (N_9596,N_8254,N_8396);
nor U9597 (N_9597,N_7562,N_8006);
or U9598 (N_9598,N_8470,N_8089);
xnor U9599 (N_9599,N_7518,N_8901);
xor U9600 (N_9600,N_8011,N_8250);
xor U9601 (N_9601,N_8923,N_8417);
xnor U9602 (N_9602,N_8631,N_7719);
nor U9603 (N_9603,N_7700,N_8597);
or U9604 (N_9604,N_7533,N_7877);
and U9605 (N_9605,N_8095,N_7611);
nand U9606 (N_9606,N_8333,N_8731);
and U9607 (N_9607,N_8833,N_8661);
nor U9608 (N_9608,N_8567,N_8394);
xor U9609 (N_9609,N_8232,N_8872);
and U9610 (N_9610,N_8132,N_7602);
nor U9611 (N_9611,N_7586,N_8018);
nand U9612 (N_9612,N_7726,N_7977);
and U9613 (N_9613,N_8893,N_8320);
nand U9614 (N_9614,N_8956,N_8618);
nor U9615 (N_9615,N_8666,N_8317);
nor U9616 (N_9616,N_7832,N_8143);
nor U9617 (N_9617,N_8188,N_8516);
and U9618 (N_9618,N_7879,N_8685);
nand U9619 (N_9619,N_7908,N_8442);
xor U9620 (N_9620,N_8760,N_8907);
or U9621 (N_9621,N_8170,N_8502);
nand U9622 (N_9622,N_8715,N_7959);
nor U9623 (N_9623,N_8352,N_8894);
nand U9624 (N_9624,N_7874,N_7820);
nor U9625 (N_9625,N_8877,N_7919);
nand U9626 (N_9626,N_8532,N_7677);
nand U9627 (N_9627,N_8673,N_8133);
or U9628 (N_9628,N_7509,N_8509);
nor U9629 (N_9629,N_7972,N_8342);
or U9630 (N_9630,N_8248,N_7931);
nor U9631 (N_9631,N_7816,N_8530);
or U9632 (N_9632,N_8034,N_7984);
nor U9633 (N_9633,N_8078,N_7952);
nand U9634 (N_9634,N_7826,N_8305);
nand U9635 (N_9635,N_7528,N_8543);
xor U9636 (N_9636,N_8406,N_8373);
or U9637 (N_9637,N_7596,N_7819);
and U9638 (N_9638,N_7676,N_7861);
or U9639 (N_9639,N_7758,N_8314);
nand U9640 (N_9640,N_8511,N_7815);
xor U9641 (N_9641,N_8865,N_7924);
nand U9642 (N_9642,N_8628,N_8922);
xor U9643 (N_9643,N_8504,N_8475);
and U9644 (N_9644,N_8817,N_8875);
nor U9645 (N_9645,N_7938,N_8435);
and U9646 (N_9646,N_8321,N_8497);
nor U9647 (N_9647,N_8821,N_7779);
nand U9648 (N_9648,N_8259,N_8038);
nor U9649 (N_9649,N_8204,N_8952);
nor U9650 (N_9650,N_8457,N_7687);
xnor U9651 (N_9651,N_7698,N_7691);
and U9652 (N_9652,N_8832,N_8652);
or U9653 (N_9653,N_8506,N_8400);
or U9654 (N_9654,N_7546,N_8157);
and U9655 (N_9655,N_8348,N_7901);
xnor U9656 (N_9656,N_7744,N_8235);
nand U9657 (N_9657,N_8437,N_7521);
nor U9658 (N_9658,N_8391,N_8234);
or U9659 (N_9659,N_7759,N_8326);
or U9660 (N_9660,N_8873,N_8033);
and U9661 (N_9661,N_8486,N_8158);
nand U9662 (N_9662,N_8747,N_7718);
xnor U9663 (N_9663,N_8237,N_7887);
nand U9664 (N_9664,N_7900,N_8282);
nand U9665 (N_9665,N_8735,N_8515);
nand U9666 (N_9666,N_8862,N_7623);
or U9667 (N_9667,N_8189,N_8453);
or U9668 (N_9668,N_8293,N_8150);
nor U9669 (N_9669,N_7763,N_8672);
xnor U9670 (N_9670,N_8160,N_8531);
nor U9671 (N_9671,N_7912,N_8815);
xnor U9672 (N_9672,N_8407,N_7776);
xnor U9673 (N_9673,N_7568,N_8052);
or U9674 (N_9674,N_8697,N_8570);
and U9675 (N_9675,N_8967,N_7906);
nor U9676 (N_9676,N_8481,N_7853);
xor U9677 (N_9677,N_7898,N_8521);
or U9678 (N_9678,N_8057,N_8210);
nor U9679 (N_9679,N_8828,N_8549);
and U9680 (N_9680,N_8649,N_7643);
nand U9681 (N_9681,N_8921,N_8172);
nand U9682 (N_9682,N_8723,N_8867);
and U9683 (N_9683,N_7943,N_7632);
nand U9684 (N_9684,N_8571,N_8787);
nand U9685 (N_9685,N_8369,N_8094);
and U9686 (N_9686,N_7961,N_7604);
or U9687 (N_9687,N_8563,N_7798);
nand U9688 (N_9688,N_8836,N_8586);
and U9689 (N_9689,N_8205,N_8331);
nand U9690 (N_9690,N_8595,N_7813);
and U9691 (N_9691,N_8213,N_8128);
xor U9692 (N_9692,N_8513,N_8055);
nor U9693 (N_9693,N_8678,N_7544);
nor U9694 (N_9694,N_8882,N_8782);
nand U9695 (N_9695,N_8545,N_7834);
or U9696 (N_9696,N_8704,N_8045);
nor U9697 (N_9697,N_8450,N_7543);
and U9698 (N_9698,N_8491,N_8231);
nor U9699 (N_9699,N_7936,N_8498);
xnor U9700 (N_9700,N_7793,N_8863);
and U9701 (N_9701,N_8757,N_7910);
nand U9702 (N_9702,N_8020,N_7607);
nor U9703 (N_9703,N_8822,N_8446);
or U9704 (N_9704,N_8171,N_8950);
xnor U9705 (N_9705,N_7966,N_8112);
or U9706 (N_9706,N_8520,N_8799);
nor U9707 (N_9707,N_8102,N_8230);
or U9708 (N_9708,N_7679,N_8191);
nor U9709 (N_9709,N_8474,N_8421);
nand U9710 (N_9710,N_7627,N_8638);
and U9711 (N_9711,N_8285,N_8771);
nand U9712 (N_9712,N_7771,N_8090);
nand U9713 (N_9713,N_8792,N_8243);
nor U9714 (N_9714,N_8456,N_7837);
or U9715 (N_9715,N_8973,N_7540);
and U9716 (N_9716,N_7564,N_8122);
nand U9717 (N_9717,N_7976,N_8900);
nor U9718 (N_9718,N_8663,N_8215);
xor U9719 (N_9719,N_8589,N_8551);
or U9720 (N_9720,N_8558,N_7555);
or U9721 (N_9721,N_7818,N_8371);
and U9722 (N_9722,N_8068,N_7622);
nor U9723 (N_9723,N_8154,N_8948);
nor U9724 (N_9724,N_7558,N_8621);
and U9725 (N_9725,N_8804,N_7527);
xnor U9726 (N_9726,N_8845,N_8643);
nor U9727 (N_9727,N_7724,N_7683);
xor U9728 (N_9728,N_8349,N_8580);
or U9729 (N_9729,N_8788,N_8969);
xor U9730 (N_9730,N_8418,N_8148);
or U9731 (N_9731,N_8341,N_7560);
and U9732 (N_9732,N_7964,N_8387);
nor U9733 (N_9733,N_8281,N_7660);
xor U9734 (N_9734,N_7897,N_8343);
nor U9735 (N_9735,N_8028,N_8746);
nand U9736 (N_9736,N_8153,N_8770);
nor U9737 (N_9737,N_8711,N_7978);
nand U9738 (N_9738,N_7828,N_8539);
nor U9739 (N_9739,N_8984,N_8482);
or U9740 (N_9740,N_8116,N_8167);
and U9741 (N_9741,N_8261,N_8721);
xor U9742 (N_9742,N_8887,N_7534);
nor U9743 (N_9743,N_8197,N_7550);
xnor U9744 (N_9744,N_8966,N_7773);
nand U9745 (N_9745,N_8892,N_8339);
xor U9746 (N_9746,N_8949,N_8500);
nand U9747 (N_9747,N_8472,N_8209);
and U9748 (N_9748,N_8448,N_8368);
nand U9749 (N_9749,N_7838,N_7579);
nand U9750 (N_9750,N_8165,N_8288);
nor U9751 (N_9751,N_8346,N_8285);
or U9752 (N_9752,N_7661,N_7513);
xor U9753 (N_9753,N_8686,N_8942);
and U9754 (N_9754,N_8507,N_7535);
nand U9755 (N_9755,N_8511,N_7990);
xnor U9756 (N_9756,N_7702,N_8323);
or U9757 (N_9757,N_8314,N_8370);
and U9758 (N_9758,N_8970,N_8174);
nand U9759 (N_9759,N_7503,N_7836);
nand U9760 (N_9760,N_7981,N_7817);
nand U9761 (N_9761,N_8093,N_7763);
nor U9762 (N_9762,N_7543,N_8050);
xor U9763 (N_9763,N_8452,N_7838);
nor U9764 (N_9764,N_8183,N_8981);
and U9765 (N_9765,N_8500,N_7766);
nor U9766 (N_9766,N_8654,N_8576);
nand U9767 (N_9767,N_8794,N_7777);
and U9768 (N_9768,N_8585,N_8086);
and U9769 (N_9769,N_7519,N_8140);
xnor U9770 (N_9770,N_7595,N_8891);
nand U9771 (N_9771,N_7718,N_7633);
or U9772 (N_9772,N_7547,N_8202);
xnor U9773 (N_9773,N_8353,N_7804);
xnor U9774 (N_9774,N_8928,N_7966);
nor U9775 (N_9775,N_7955,N_8854);
nor U9776 (N_9776,N_8724,N_8948);
nor U9777 (N_9777,N_8102,N_8035);
nor U9778 (N_9778,N_8610,N_8485);
xor U9779 (N_9779,N_8398,N_8892);
or U9780 (N_9780,N_8923,N_8852);
xnor U9781 (N_9781,N_8507,N_8215);
xor U9782 (N_9782,N_7721,N_8093);
or U9783 (N_9783,N_8117,N_8901);
nor U9784 (N_9784,N_8635,N_7754);
or U9785 (N_9785,N_8623,N_7609);
and U9786 (N_9786,N_8230,N_8384);
nor U9787 (N_9787,N_7536,N_8114);
xnor U9788 (N_9788,N_8817,N_7991);
nor U9789 (N_9789,N_8234,N_8383);
nand U9790 (N_9790,N_8630,N_8368);
or U9791 (N_9791,N_8248,N_8679);
or U9792 (N_9792,N_7606,N_8138);
and U9793 (N_9793,N_7842,N_8939);
nor U9794 (N_9794,N_8755,N_7759);
nand U9795 (N_9795,N_7510,N_8927);
nand U9796 (N_9796,N_8632,N_8646);
or U9797 (N_9797,N_7781,N_7900);
or U9798 (N_9798,N_8228,N_7519);
and U9799 (N_9799,N_8726,N_7796);
nor U9800 (N_9800,N_7635,N_7646);
xnor U9801 (N_9801,N_8888,N_7959);
nor U9802 (N_9802,N_8484,N_7739);
nand U9803 (N_9803,N_8714,N_8636);
or U9804 (N_9804,N_8612,N_7967);
or U9805 (N_9805,N_8807,N_8840);
and U9806 (N_9806,N_8956,N_7504);
and U9807 (N_9807,N_7505,N_8499);
nand U9808 (N_9808,N_8216,N_8594);
xnor U9809 (N_9809,N_7755,N_7641);
xnor U9810 (N_9810,N_7940,N_7504);
or U9811 (N_9811,N_8219,N_7604);
xor U9812 (N_9812,N_8778,N_8601);
xor U9813 (N_9813,N_8554,N_8099);
or U9814 (N_9814,N_8160,N_8208);
and U9815 (N_9815,N_7844,N_7771);
and U9816 (N_9816,N_7815,N_8907);
nor U9817 (N_9817,N_8848,N_7804);
and U9818 (N_9818,N_8017,N_7781);
xor U9819 (N_9819,N_7626,N_8987);
or U9820 (N_9820,N_8375,N_8854);
and U9821 (N_9821,N_8749,N_7901);
nor U9822 (N_9822,N_8293,N_8639);
and U9823 (N_9823,N_8267,N_8178);
xnor U9824 (N_9824,N_8639,N_7986);
nor U9825 (N_9825,N_7617,N_8914);
and U9826 (N_9826,N_8879,N_8300);
and U9827 (N_9827,N_8980,N_7881);
nor U9828 (N_9828,N_7942,N_7589);
nand U9829 (N_9829,N_7510,N_8135);
nor U9830 (N_9830,N_8115,N_8063);
or U9831 (N_9831,N_8703,N_8979);
or U9832 (N_9832,N_7857,N_8989);
nand U9833 (N_9833,N_8433,N_7624);
nand U9834 (N_9834,N_8930,N_8834);
nor U9835 (N_9835,N_8620,N_8790);
nor U9836 (N_9836,N_8850,N_8262);
xnor U9837 (N_9837,N_7547,N_8513);
xor U9838 (N_9838,N_8038,N_7970);
xnor U9839 (N_9839,N_8367,N_8907);
or U9840 (N_9840,N_7690,N_7879);
nor U9841 (N_9841,N_8907,N_8292);
nand U9842 (N_9842,N_8943,N_7810);
or U9843 (N_9843,N_8732,N_8139);
nor U9844 (N_9844,N_7574,N_8077);
nor U9845 (N_9845,N_7570,N_8442);
nor U9846 (N_9846,N_8743,N_7759);
xnor U9847 (N_9847,N_8759,N_8652);
nand U9848 (N_9848,N_8056,N_8935);
nand U9849 (N_9849,N_8952,N_8496);
nand U9850 (N_9850,N_8484,N_8700);
xnor U9851 (N_9851,N_8483,N_8764);
nand U9852 (N_9852,N_8891,N_8770);
nand U9853 (N_9853,N_7998,N_8661);
and U9854 (N_9854,N_8065,N_8745);
nand U9855 (N_9855,N_8512,N_8081);
or U9856 (N_9856,N_8601,N_8570);
or U9857 (N_9857,N_8664,N_8216);
or U9858 (N_9858,N_8806,N_8587);
and U9859 (N_9859,N_8743,N_7889);
and U9860 (N_9860,N_8499,N_8303);
xnor U9861 (N_9861,N_8445,N_7891);
and U9862 (N_9862,N_8980,N_7892);
nor U9863 (N_9863,N_8891,N_8429);
nand U9864 (N_9864,N_7744,N_8438);
and U9865 (N_9865,N_8494,N_8803);
xor U9866 (N_9866,N_7631,N_8933);
xor U9867 (N_9867,N_8957,N_7578);
xnor U9868 (N_9868,N_7792,N_7732);
nor U9869 (N_9869,N_8616,N_7623);
or U9870 (N_9870,N_7682,N_8676);
nand U9871 (N_9871,N_7568,N_8735);
nor U9872 (N_9872,N_8457,N_8244);
xnor U9873 (N_9873,N_8911,N_8250);
xnor U9874 (N_9874,N_7841,N_7894);
xor U9875 (N_9875,N_8803,N_8720);
or U9876 (N_9876,N_8966,N_8311);
xor U9877 (N_9877,N_7908,N_7777);
or U9878 (N_9878,N_8334,N_7529);
and U9879 (N_9879,N_8606,N_8804);
nor U9880 (N_9880,N_8785,N_7803);
or U9881 (N_9881,N_7659,N_8947);
nand U9882 (N_9882,N_8562,N_7602);
nor U9883 (N_9883,N_8019,N_8456);
nand U9884 (N_9884,N_8981,N_8119);
nor U9885 (N_9885,N_8067,N_8531);
nand U9886 (N_9886,N_7746,N_8423);
xnor U9887 (N_9887,N_8626,N_8010);
nand U9888 (N_9888,N_8115,N_8944);
xor U9889 (N_9889,N_8961,N_8257);
and U9890 (N_9890,N_7586,N_7699);
nand U9891 (N_9891,N_7884,N_8324);
nor U9892 (N_9892,N_7530,N_8661);
nand U9893 (N_9893,N_8038,N_7793);
nand U9894 (N_9894,N_8237,N_8492);
or U9895 (N_9895,N_7722,N_8982);
and U9896 (N_9896,N_8561,N_7932);
xnor U9897 (N_9897,N_7571,N_7659);
or U9898 (N_9898,N_7553,N_8762);
nor U9899 (N_9899,N_7565,N_7637);
or U9900 (N_9900,N_8724,N_7557);
and U9901 (N_9901,N_8322,N_8164);
or U9902 (N_9902,N_8088,N_8446);
and U9903 (N_9903,N_8445,N_8841);
and U9904 (N_9904,N_8388,N_8851);
xor U9905 (N_9905,N_8465,N_8269);
xor U9906 (N_9906,N_8343,N_8656);
and U9907 (N_9907,N_8186,N_8428);
xnor U9908 (N_9908,N_8525,N_7831);
nor U9909 (N_9909,N_8780,N_7800);
xnor U9910 (N_9910,N_7870,N_7576);
nand U9911 (N_9911,N_8489,N_7937);
nor U9912 (N_9912,N_8149,N_8234);
and U9913 (N_9913,N_8827,N_8789);
and U9914 (N_9914,N_8724,N_8337);
nand U9915 (N_9915,N_8042,N_8875);
and U9916 (N_9916,N_7557,N_7760);
and U9917 (N_9917,N_7875,N_8062);
and U9918 (N_9918,N_8550,N_8085);
or U9919 (N_9919,N_8929,N_7991);
and U9920 (N_9920,N_8506,N_8952);
nand U9921 (N_9921,N_8556,N_8203);
and U9922 (N_9922,N_8402,N_7556);
or U9923 (N_9923,N_7812,N_7819);
nand U9924 (N_9924,N_7725,N_8174);
nand U9925 (N_9925,N_8169,N_8223);
xor U9926 (N_9926,N_7916,N_7985);
nor U9927 (N_9927,N_8436,N_7943);
xor U9928 (N_9928,N_8127,N_7981);
nor U9929 (N_9929,N_8947,N_7870);
and U9930 (N_9930,N_8922,N_8611);
xnor U9931 (N_9931,N_7687,N_8984);
xor U9932 (N_9932,N_8337,N_7699);
and U9933 (N_9933,N_7918,N_7647);
or U9934 (N_9934,N_7562,N_8695);
or U9935 (N_9935,N_7672,N_8632);
xnor U9936 (N_9936,N_8065,N_8188);
and U9937 (N_9937,N_8084,N_8818);
xnor U9938 (N_9938,N_8666,N_8882);
xor U9939 (N_9939,N_8724,N_8102);
xnor U9940 (N_9940,N_8734,N_7528);
nor U9941 (N_9941,N_8135,N_8618);
nor U9942 (N_9942,N_8121,N_8954);
nand U9943 (N_9943,N_8431,N_8055);
and U9944 (N_9944,N_8670,N_8487);
nor U9945 (N_9945,N_8413,N_8539);
and U9946 (N_9946,N_8161,N_8229);
or U9947 (N_9947,N_8582,N_8558);
nor U9948 (N_9948,N_8917,N_8809);
nor U9949 (N_9949,N_8623,N_8793);
or U9950 (N_9950,N_8502,N_7545);
xor U9951 (N_9951,N_8670,N_8819);
nand U9952 (N_9952,N_8353,N_8544);
xor U9953 (N_9953,N_8731,N_8555);
nand U9954 (N_9954,N_8893,N_7649);
or U9955 (N_9955,N_8173,N_8012);
or U9956 (N_9956,N_7877,N_7945);
nand U9957 (N_9957,N_8539,N_8400);
and U9958 (N_9958,N_8454,N_8692);
nand U9959 (N_9959,N_8170,N_8627);
nand U9960 (N_9960,N_7502,N_8705);
and U9961 (N_9961,N_8107,N_8188);
nor U9962 (N_9962,N_7926,N_8355);
or U9963 (N_9963,N_8429,N_7886);
nor U9964 (N_9964,N_8491,N_8866);
nor U9965 (N_9965,N_8263,N_7795);
or U9966 (N_9966,N_8968,N_8238);
and U9967 (N_9967,N_8966,N_8394);
or U9968 (N_9968,N_8490,N_7819);
nor U9969 (N_9969,N_7903,N_8797);
and U9970 (N_9970,N_8985,N_8387);
nand U9971 (N_9971,N_8569,N_8356);
nor U9972 (N_9972,N_8360,N_8147);
or U9973 (N_9973,N_7901,N_7868);
nor U9974 (N_9974,N_8403,N_7996);
nand U9975 (N_9975,N_8979,N_8824);
or U9976 (N_9976,N_8123,N_7696);
nand U9977 (N_9977,N_8257,N_8662);
xor U9978 (N_9978,N_8011,N_8827);
and U9979 (N_9979,N_7980,N_7958);
nand U9980 (N_9980,N_8307,N_7771);
and U9981 (N_9981,N_7664,N_7696);
or U9982 (N_9982,N_8396,N_8058);
xor U9983 (N_9983,N_8687,N_7614);
nand U9984 (N_9984,N_8950,N_8843);
nand U9985 (N_9985,N_7651,N_7803);
xnor U9986 (N_9986,N_7825,N_7755);
nand U9987 (N_9987,N_8848,N_7995);
nor U9988 (N_9988,N_8238,N_8911);
nand U9989 (N_9989,N_8288,N_8162);
nand U9990 (N_9990,N_8695,N_8659);
nor U9991 (N_9991,N_7682,N_8649);
nand U9992 (N_9992,N_8752,N_8445);
and U9993 (N_9993,N_8284,N_8875);
and U9994 (N_9994,N_8200,N_8838);
and U9995 (N_9995,N_8941,N_8356);
and U9996 (N_9996,N_7816,N_8001);
and U9997 (N_9997,N_8839,N_8825);
and U9998 (N_9998,N_8490,N_7843);
or U9999 (N_9999,N_8565,N_8189);
nor U10000 (N_10000,N_8351,N_8763);
or U10001 (N_10001,N_8531,N_7936);
or U10002 (N_10002,N_8395,N_8733);
and U10003 (N_10003,N_7628,N_8589);
xnor U10004 (N_10004,N_8337,N_8022);
nor U10005 (N_10005,N_8597,N_8586);
or U10006 (N_10006,N_8152,N_8485);
and U10007 (N_10007,N_8931,N_7618);
and U10008 (N_10008,N_8456,N_8078);
or U10009 (N_10009,N_8038,N_8769);
xor U10010 (N_10010,N_8328,N_7910);
nor U10011 (N_10011,N_8981,N_7829);
nand U10012 (N_10012,N_8285,N_8615);
or U10013 (N_10013,N_8291,N_7545);
and U10014 (N_10014,N_8203,N_8423);
nand U10015 (N_10015,N_7992,N_8348);
and U10016 (N_10016,N_7683,N_7786);
nand U10017 (N_10017,N_8767,N_8355);
or U10018 (N_10018,N_8956,N_7752);
or U10019 (N_10019,N_8200,N_8722);
and U10020 (N_10020,N_8626,N_8794);
xor U10021 (N_10021,N_8391,N_7506);
xnor U10022 (N_10022,N_8760,N_7917);
xor U10023 (N_10023,N_8252,N_8165);
and U10024 (N_10024,N_8557,N_8948);
nor U10025 (N_10025,N_7836,N_8522);
or U10026 (N_10026,N_8734,N_7902);
and U10027 (N_10027,N_8900,N_8952);
and U10028 (N_10028,N_8537,N_8037);
nand U10029 (N_10029,N_7734,N_7912);
or U10030 (N_10030,N_7726,N_8991);
nand U10031 (N_10031,N_8695,N_8210);
xnor U10032 (N_10032,N_8597,N_8269);
nor U10033 (N_10033,N_7534,N_8994);
or U10034 (N_10034,N_8628,N_8003);
xnor U10035 (N_10035,N_8581,N_8970);
or U10036 (N_10036,N_8705,N_8786);
nor U10037 (N_10037,N_7652,N_7557);
or U10038 (N_10038,N_8944,N_8471);
or U10039 (N_10039,N_8062,N_7654);
nor U10040 (N_10040,N_8647,N_8362);
xor U10041 (N_10041,N_8254,N_7805);
xnor U10042 (N_10042,N_7639,N_7962);
nand U10043 (N_10043,N_7546,N_8747);
nand U10044 (N_10044,N_8124,N_8630);
nand U10045 (N_10045,N_7607,N_8041);
nand U10046 (N_10046,N_8075,N_7901);
nand U10047 (N_10047,N_8104,N_7973);
nor U10048 (N_10048,N_8816,N_7940);
nand U10049 (N_10049,N_7765,N_8500);
xor U10050 (N_10050,N_8474,N_7785);
nand U10051 (N_10051,N_8458,N_8738);
xnor U10052 (N_10052,N_7828,N_8540);
or U10053 (N_10053,N_8472,N_8297);
nor U10054 (N_10054,N_8511,N_8878);
nor U10055 (N_10055,N_8051,N_7586);
and U10056 (N_10056,N_8853,N_8843);
or U10057 (N_10057,N_8684,N_7754);
xnor U10058 (N_10058,N_7509,N_8329);
xnor U10059 (N_10059,N_8174,N_8506);
nand U10060 (N_10060,N_8813,N_8155);
xor U10061 (N_10061,N_8105,N_7622);
and U10062 (N_10062,N_8215,N_8202);
xnor U10063 (N_10063,N_8286,N_8993);
or U10064 (N_10064,N_8081,N_7841);
nand U10065 (N_10065,N_8206,N_8791);
nor U10066 (N_10066,N_8730,N_7732);
xor U10067 (N_10067,N_8095,N_7593);
nor U10068 (N_10068,N_7715,N_7584);
and U10069 (N_10069,N_8743,N_8324);
and U10070 (N_10070,N_8739,N_8922);
nand U10071 (N_10071,N_7999,N_7995);
and U10072 (N_10072,N_8484,N_7833);
nand U10073 (N_10073,N_8496,N_8863);
and U10074 (N_10074,N_8106,N_8748);
or U10075 (N_10075,N_8943,N_8031);
nand U10076 (N_10076,N_7881,N_8665);
xor U10077 (N_10077,N_8061,N_7670);
and U10078 (N_10078,N_8081,N_8554);
nand U10079 (N_10079,N_7590,N_8182);
nor U10080 (N_10080,N_8683,N_7608);
and U10081 (N_10081,N_8925,N_7956);
and U10082 (N_10082,N_8157,N_7726);
and U10083 (N_10083,N_8828,N_7654);
nand U10084 (N_10084,N_8913,N_7938);
nor U10085 (N_10085,N_8415,N_8872);
nand U10086 (N_10086,N_8875,N_8133);
nand U10087 (N_10087,N_8934,N_8874);
xnor U10088 (N_10088,N_7974,N_8811);
nor U10089 (N_10089,N_7747,N_8762);
and U10090 (N_10090,N_8270,N_7832);
or U10091 (N_10091,N_8063,N_8472);
nand U10092 (N_10092,N_8117,N_8319);
nor U10093 (N_10093,N_7825,N_8951);
and U10094 (N_10094,N_7731,N_7924);
nand U10095 (N_10095,N_7677,N_8471);
nor U10096 (N_10096,N_8710,N_7508);
nand U10097 (N_10097,N_8337,N_8647);
nor U10098 (N_10098,N_8272,N_7739);
xnor U10099 (N_10099,N_7888,N_8238);
or U10100 (N_10100,N_8721,N_8211);
nand U10101 (N_10101,N_8910,N_8307);
or U10102 (N_10102,N_8749,N_8799);
and U10103 (N_10103,N_8189,N_8147);
xor U10104 (N_10104,N_8048,N_8445);
and U10105 (N_10105,N_8279,N_8968);
or U10106 (N_10106,N_7872,N_7946);
or U10107 (N_10107,N_7807,N_7961);
nor U10108 (N_10108,N_7780,N_7576);
nand U10109 (N_10109,N_8776,N_8504);
or U10110 (N_10110,N_7851,N_7707);
xnor U10111 (N_10111,N_8214,N_7732);
and U10112 (N_10112,N_7545,N_8182);
xnor U10113 (N_10113,N_8011,N_7833);
nor U10114 (N_10114,N_8429,N_8922);
nor U10115 (N_10115,N_8248,N_8224);
nor U10116 (N_10116,N_8642,N_7761);
xnor U10117 (N_10117,N_8266,N_8685);
nor U10118 (N_10118,N_8374,N_7910);
nand U10119 (N_10119,N_8342,N_8914);
and U10120 (N_10120,N_8416,N_8768);
and U10121 (N_10121,N_8497,N_7611);
nor U10122 (N_10122,N_8752,N_8285);
nand U10123 (N_10123,N_8953,N_7706);
nand U10124 (N_10124,N_8823,N_7541);
nor U10125 (N_10125,N_7717,N_8725);
xnor U10126 (N_10126,N_8758,N_7702);
and U10127 (N_10127,N_8720,N_8267);
or U10128 (N_10128,N_7601,N_7523);
nand U10129 (N_10129,N_7811,N_8415);
or U10130 (N_10130,N_7590,N_8899);
or U10131 (N_10131,N_8310,N_7846);
or U10132 (N_10132,N_8210,N_8083);
nor U10133 (N_10133,N_7717,N_8858);
xor U10134 (N_10134,N_8102,N_7646);
and U10135 (N_10135,N_8901,N_8268);
or U10136 (N_10136,N_8874,N_8836);
or U10137 (N_10137,N_8464,N_8777);
xnor U10138 (N_10138,N_8373,N_7691);
and U10139 (N_10139,N_8470,N_8195);
nor U10140 (N_10140,N_8127,N_8785);
or U10141 (N_10141,N_8687,N_8507);
or U10142 (N_10142,N_8760,N_8597);
or U10143 (N_10143,N_8344,N_8411);
nand U10144 (N_10144,N_7708,N_8234);
nand U10145 (N_10145,N_8206,N_7791);
or U10146 (N_10146,N_8926,N_7919);
or U10147 (N_10147,N_7536,N_7809);
nand U10148 (N_10148,N_8795,N_7906);
nand U10149 (N_10149,N_8797,N_7599);
and U10150 (N_10150,N_7873,N_8713);
and U10151 (N_10151,N_8053,N_8959);
nor U10152 (N_10152,N_7703,N_7945);
and U10153 (N_10153,N_8876,N_7924);
and U10154 (N_10154,N_8787,N_7598);
or U10155 (N_10155,N_8272,N_8858);
nand U10156 (N_10156,N_8605,N_7709);
or U10157 (N_10157,N_8368,N_8758);
xnor U10158 (N_10158,N_8970,N_8850);
and U10159 (N_10159,N_8504,N_8057);
and U10160 (N_10160,N_7779,N_7657);
or U10161 (N_10161,N_7872,N_8715);
nand U10162 (N_10162,N_8147,N_8608);
xor U10163 (N_10163,N_8544,N_8642);
and U10164 (N_10164,N_8211,N_8876);
or U10165 (N_10165,N_7892,N_8107);
and U10166 (N_10166,N_8770,N_7933);
and U10167 (N_10167,N_8360,N_8699);
nor U10168 (N_10168,N_8720,N_7675);
nand U10169 (N_10169,N_8066,N_7519);
nand U10170 (N_10170,N_8111,N_8547);
xnor U10171 (N_10171,N_8606,N_8731);
or U10172 (N_10172,N_7714,N_8422);
xor U10173 (N_10173,N_8317,N_8376);
and U10174 (N_10174,N_7790,N_7702);
or U10175 (N_10175,N_7650,N_8494);
nor U10176 (N_10176,N_8835,N_8681);
nand U10177 (N_10177,N_8110,N_8585);
nor U10178 (N_10178,N_7891,N_8710);
and U10179 (N_10179,N_8190,N_8070);
and U10180 (N_10180,N_8609,N_8521);
nor U10181 (N_10181,N_8263,N_8758);
and U10182 (N_10182,N_8931,N_7672);
and U10183 (N_10183,N_8299,N_8262);
and U10184 (N_10184,N_7781,N_8171);
or U10185 (N_10185,N_8749,N_8180);
xnor U10186 (N_10186,N_7696,N_7669);
xor U10187 (N_10187,N_8763,N_7540);
nand U10188 (N_10188,N_7746,N_8794);
nand U10189 (N_10189,N_7509,N_8393);
nand U10190 (N_10190,N_8713,N_8758);
and U10191 (N_10191,N_7998,N_8159);
nand U10192 (N_10192,N_8677,N_8612);
or U10193 (N_10193,N_7826,N_8442);
xnor U10194 (N_10194,N_8573,N_8461);
and U10195 (N_10195,N_7603,N_7519);
and U10196 (N_10196,N_8864,N_8238);
nand U10197 (N_10197,N_7626,N_7664);
nor U10198 (N_10198,N_8882,N_8063);
nor U10199 (N_10199,N_8461,N_7780);
nand U10200 (N_10200,N_8015,N_7729);
and U10201 (N_10201,N_7604,N_8577);
nand U10202 (N_10202,N_8874,N_8955);
nand U10203 (N_10203,N_7555,N_7989);
xor U10204 (N_10204,N_7895,N_7767);
or U10205 (N_10205,N_8426,N_7889);
and U10206 (N_10206,N_8066,N_7752);
or U10207 (N_10207,N_8021,N_7653);
nand U10208 (N_10208,N_8729,N_8973);
nand U10209 (N_10209,N_8234,N_8463);
nand U10210 (N_10210,N_7512,N_8864);
nand U10211 (N_10211,N_7579,N_8332);
or U10212 (N_10212,N_8190,N_8495);
xnor U10213 (N_10213,N_8684,N_8376);
and U10214 (N_10214,N_7733,N_8538);
and U10215 (N_10215,N_8380,N_8112);
nand U10216 (N_10216,N_8726,N_7518);
or U10217 (N_10217,N_7677,N_8108);
and U10218 (N_10218,N_8168,N_7589);
nand U10219 (N_10219,N_7585,N_7758);
and U10220 (N_10220,N_8994,N_8194);
nand U10221 (N_10221,N_8790,N_7723);
nor U10222 (N_10222,N_7747,N_8689);
nor U10223 (N_10223,N_7500,N_8580);
and U10224 (N_10224,N_8154,N_8188);
nand U10225 (N_10225,N_8440,N_8496);
nor U10226 (N_10226,N_8518,N_8204);
nor U10227 (N_10227,N_7910,N_8398);
xor U10228 (N_10228,N_8786,N_8531);
xnor U10229 (N_10229,N_8726,N_7653);
and U10230 (N_10230,N_7964,N_7778);
or U10231 (N_10231,N_8562,N_8171);
nand U10232 (N_10232,N_8960,N_7659);
nand U10233 (N_10233,N_7886,N_7513);
xor U10234 (N_10234,N_7538,N_8292);
nor U10235 (N_10235,N_7881,N_8400);
nor U10236 (N_10236,N_7982,N_7734);
or U10237 (N_10237,N_8208,N_7794);
nand U10238 (N_10238,N_8797,N_7582);
nor U10239 (N_10239,N_8966,N_7884);
nor U10240 (N_10240,N_8632,N_7764);
nor U10241 (N_10241,N_8519,N_7665);
or U10242 (N_10242,N_7677,N_8586);
xnor U10243 (N_10243,N_8712,N_7560);
nand U10244 (N_10244,N_8771,N_8996);
nor U10245 (N_10245,N_7657,N_7987);
or U10246 (N_10246,N_8621,N_7593);
nand U10247 (N_10247,N_7844,N_8521);
or U10248 (N_10248,N_7534,N_7921);
xor U10249 (N_10249,N_8235,N_8787);
xor U10250 (N_10250,N_8643,N_7554);
or U10251 (N_10251,N_8865,N_8511);
nand U10252 (N_10252,N_8282,N_8169);
nand U10253 (N_10253,N_8969,N_8236);
nand U10254 (N_10254,N_7892,N_8852);
or U10255 (N_10255,N_8673,N_8816);
nand U10256 (N_10256,N_8833,N_8914);
and U10257 (N_10257,N_8624,N_7969);
xor U10258 (N_10258,N_7815,N_7806);
nand U10259 (N_10259,N_8674,N_7657);
nor U10260 (N_10260,N_8967,N_8237);
nand U10261 (N_10261,N_7677,N_8744);
or U10262 (N_10262,N_8420,N_8761);
and U10263 (N_10263,N_7637,N_7729);
nand U10264 (N_10264,N_8742,N_8956);
xnor U10265 (N_10265,N_8360,N_8477);
nor U10266 (N_10266,N_8363,N_8220);
nand U10267 (N_10267,N_8344,N_8376);
xor U10268 (N_10268,N_8554,N_7659);
nor U10269 (N_10269,N_7543,N_7723);
and U10270 (N_10270,N_8988,N_8210);
nand U10271 (N_10271,N_8186,N_8823);
xnor U10272 (N_10272,N_8065,N_7807);
nor U10273 (N_10273,N_7613,N_8169);
xor U10274 (N_10274,N_8064,N_8760);
nand U10275 (N_10275,N_7703,N_8169);
nor U10276 (N_10276,N_7960,N_7792);
or U10277 (N_10277,N_7838,N_7780);
nand U10278 (N_10278,N_7796,N_8653);
and U10279 (N_10279,N_8517,N_8625);
nor U10280 (N_10280,N_7816,N_8458);
xnor U10281 (N_10281,N_8870,N_8352);
xnor U10282 (N_10282,N_7862,N_8513);
nor U10283 (N_10283,N_8121,N_8071);
and U10284 (N_10284,N_8792,N_7876);
xor U10285 (N_10285,N_8197,N_8934);
nand U10286 (N_10286,N_7962,N_8966);
and U10287 (N_10287,N_8990,N_8617);
or U10288 (N_10288,N_8555,N_7714);
or U10289 (N_10289,N_8888,N_7737);
or U10290 (N_10290,N_8104,N_8810);
nor U10291 (N_10291,N_7579,N_8696);
xor U10292 (N_10292,N_8915,N_7599);
nor U10293 (N_10293,N_8302,N_8218);
xnor U10294 (N_10294,N_8430,N_8579);
or U10295 (N_10295,N_8908,N_8197);
and U10296 (N_10296,N_8244,N_8134);
or U10297 (N_10297,N_8673,N_8792);
and U10298 (N_10298,N_8915,N_8921);
nand U10299 (N_10299,N_8730,N_7523);
xnor U10300 (N_10300,N_8334,N_7992);
nor U10301 (N_10301,N_8552,N_8396);
xor U10302 (N_10302,N_8220,N_8445);
nor U10303 (N_10303,N_8274,N_8876);
and U10304 (N_10304,N_7817,N_8497);
nand U10305 (N_10305,N_8761,N_8327);
or U10306 (N_10306,N_7956,N_8640);
or U10307 (N_10307,N_8858,N_8010);
and U10308 (N_10308,N_8138,N_8100);
or U10309 (N_10309,N_8081,N_8682);
nand U10310 (N_10310,N_8295,N_7930);
and U10311 (N_10311,N_8121,N_7657);
nand U10312 (N_10312,N_7588,N_8759);
nand U10313 (N_10313,N_8447,N_8295);
or U10314 (N_10314,N_7749,N_8858);
nand U10315 (N_10315,N_8518,N_8147);
nand U10316 (N_10316,N_7905,N_8115);
and U10317 (N_10317,N_8530,N_8410);
or U10318 (N_10318,N_8281,N_7506);
xor U10319 (N_10319,N_8565,N_8731);
and U10320 (N_10320,N_7648,N_8214);
and U10321 (N_10321,N_7549,N_7668);
nand U10322 (N_10322,N_8442,N_8822);
xnor U10323 (N_10323,N_8251,N_8665);
and U10324 (N_10324,N_7564,N_8353);
nor U10325 (N_10325,N_7766,N_8602);
nor U10326 (N_10326,N_8480,N_8924);
nand U10327 (N_10327,N_7665,N_7850);
nand U10328 (N_10328,N_7820,N_8770);
or U10329 (N_10329,N_8100,N_7509);
and U10330 (N_10330,N_7789,N_8598);
xnor U10331 (N_10331,N_8738,N_8510);
nor U10332 (N_10332,N_8368,N_7543);
and U10333 (N_10333,N_8907,N_8908);
and U10334 (N_10334,N_8265,N_8546);
nor U10335 (N_10335,N_8640,N_7613);
xor U10336 (N_10336,N_8700,N_8398);
nand U10337 (N_10337,N_7740,N_8847);
nor U10338 (N_10338,N_7977,N_7782);
and U10339 (N_10339,N_8698,N_7831);
nor U10340 (N_10340,N_7991,N_8536);
xnor U10341 (N_10341,N_8421,N_7653);
nor U10342 (N_10342,N_8958,N_7819);
xor U10343 (N_10343,N_8570,N_8289);
xnor U10344 (N_10344,N_7843,N_7859);
or U10345 (N_10345,N_8663,N_8596);
or U10346 (N_10346,N_7500,N_8711);
or U10347 (N_10347,N_8465,N_8514);
nor U10348 (N_10348,N_7908,N_7720);
nor U10349 (N_10349,N_8473,N_8118);
or U10350 (N_10350,N_7528,N_7780);
or U10351 (N_10351,N_7508,N_8096);
nand U10352 (N_10352,N_8120,N_8716);
and U10353 (N_10353,N_8602,N_7786);
or U10354 (N_10354,N_8297,N_7511);
xor U10355 (N_10355,N_7542,N_8474);
nand U10356 (N_10356,N_8909,N_7749);
xnor U10357 (N_10357,N_8955,N_8490);
xor U10358 (N_10358,N_8492,N_7752);
and U10359 (N_10359,N_8512,N_8781);
nor U10360 (N_10360,N_8244,N_8329);
and U10361 (N_10361,N_7994,N_8988);
nor U10362 (N_10362,N_8522,N_8005);
nand U10363 (N_10363,N_8097,N_8257);
nand U10364 (N_10364,N_8849,N_8983);
nand U10365 (N_10365,N_8871,N_8944);
xor U10366 (N_10366,N_7971,N_8654);
nor U10367 (N_10367,N_8391,N_8003);
nand U10368 (N_10368,N_7524,N_8430);
and U10369 (N_10369,N_7533,N_7950);
and U10370 (N_10370,N_7814,N_7530);
and U10371 (N_10371,N_7956,N_8691);
xor U10372 (N_10372,N_8648,N_7637);
nand U10373 (N_10373,N_8827,N_8654);
and U10374 (N_10374,N_8393,N_8712);
xnor U10375 (N_10375,N_7706,N_7858);
nand U10376 (N_10376,N_8113,N_8025);
or U10377 (N_10377,N_7988,N_8873);
xor U10378 (N_10378,N_7725,N_7578);
and U10379 (N_10379,N_8558,N_8130);
or U10380 (N_10380,N_8151,N_8418);
and U10381 (N_10381,N_8932,N_7830);
and U10382 (N_10382,N_7718,N_8159);
nor U10383 (N_10383,N_8153,N_8238);
or U10384 (N_10384,N_7859,N_7985);
and U10385 (N_10385,N_8367,N_7723);
or U10386 (N_10386,N_8714,N_8602);
and U10387 (N_10387,N_8045,N_8009);
or U10388 (N_10388,N_8006,N_8895);
and U10389 (N_10389,N_8026,N_7745);
or U10390 (N_10390,N_7549,N_8919);
nand U10391 (N_10391,N_8949,N_7543);
and U10392 (N_10392,N_8268,N_8715);
nand U10393 (N_10393,N_8264,N_8500);
or U10394 (N_10394,N_8941,N_8765);
nor U10395 (N_10395,N_8633,N_7990);
xnor U10396 (N_10396,N_8650,N_8566);
nand U10397 (N_10397,N_8804,N_8406);
and U10398 (N_10398,N_8185,N_8461);
or U10399 (N_10399,N_8359,N_8783);
and U10400 (N_10400,N_8851,N_8566);
nor U10401 (N_10401,N_7975,N_8868);
nor U10402 (N_10402,N_7682,N_8351);
nor U10403 (N_10403,N_8775,N_8708);
nor U10404 (N_10404,N_8765,N_8743);
nor U10405 (N_10405,N_8812,N_7547);
or U10406 (N_10406,N_8492,N_8506);
or U10407 (N_10407,N_8127,N_8927);
xor U10408 (N_10408,N_8463,N_7749);
or U10409 (N_10409,N_7852,N_8510);
xnor U10410 (N_10410,N_8972,N_8166);
xor U10411 (N_10411,N_7794,N_8393);
and U10412 (N_10412,N_7521,N_8620);
xor U10413 (N_10413,N_8756,N_8069);
and U10414 (N_10414,N_8719,N_8459);
or U10415 (N_10415,N_8729,N_8126);
xnor U10416 (N_10416,N_8416,N_8810);
and U10417 (N_10417,N_7803,N_7714);
nand U10418 (N_10418,N_8594,N_8769);
or U10419 (N_10419,N_8922,N_8740);
and U10420 (N_10420,N_8097,N_8481);
or U10421 (N_10421,N_8664,N_8313);
or U10422 (N_10422,N_8580,N_8457);
nand U10423 (N_10423,N_8120,N_8972);
xor U10424 (N_10424,N_8085,N_7842);
and U10425 (N_10425,N_7905,N_8228);
and U10426 (N_10426,N_8998,N_7822);
nand U10427 (N_10427,N_8859,N_7608);
and U10428 (N_10428,N_8132,N_8080);
or U10429 (N_10429,N_8811,N_8646);
and U10430 (N_10430,N_7680,N_8751);
nand U10431 (N_10431,N_8449,N_7547);
nor U10432 (N_10432,N_8329,N_7724);
and U10433 (N_10433,N_8939,N_8726);
and U10434 (N_10434,N_8821,N_7915);
nor U10435 (N_10435,N_8817,N_8025);
nand U10436 (N_10436,N_8236,N_8634);
xnor U10437 (N_10437,N_8615,N_8112);
nor U10438 (N_10438,N_8121,N_8547);
xor U10439 (N_10439,N_8099,N_8081);
or U10440 (N_10440,N_7605,N_8973);
or U10441 (N_10441,N_7739,N_7719);
or U10442 (N_10442,N_8865,N_7944);
nor U10443 (N_10443,N_8910,N_7645);
xor U10444 (N_10444,N_7763,N_8706);
or U10445 (N_10445,N_8127,N_8405);
nor U10446 (N_10446,N_8694,N_8438);
nor U10447 (N_10447,N_7872,N_7940);
nor U10448 (N_10448,N_8770,N_8646);
nor U10449 (N_10449,N_8976,N_8787);
and U10450 (N_10450,N_8528,N_8558);
nor U10451 (N_10451,N_7540,N_8626);
nand U10452 (N_10452,N_8223,N_7613);
and U10453 (N_10453,N_8674,N_8637);
nor U10454 (N_10454,N_8324,N_8425);
nor U10455 (N_10455,N_8384,N_7670);
and U10456 (N_10456,N_7748,N_8252);
xnor U10457 (N_10457,N_8068,N_8854);
nand U10458 (N_10458,N_7737,N_8617);
or U10459 (N_10459,N_8836,N_8041);
and U10460 (N_10460,N_8101,N_7867);
nor U10461 (N_10461,N_7991,N_7580);
nand U10462 (N_10462,N_8324,N_8438);
nand U10463 (N_10463,N_8584,N_7681);
and U10464 (N_10464,N_7885,N_8373);
xor U10465 (N_10465,N_8078,N_7702);
nand U10466 (N_10466,N_8874,N_7934);
nand U10467 (N_10467,N_7865,N_8723);
nand U10468 (N_10468,N_7929,N_7902);
or U10469 (N_10469,N_8673,N_8729);
xnor U10470 (N_10470,N_7871,N_8601);
or U10471 (N_10471,N_8282,N_8952);
and U10472 (N_10472,N_8079,N_7888);
or U10473 (N_10473,N_7788,N_8806);
xnor U10474 (N_10474,N_8281,N_7601);
nor U10475 (N_10475,N_7580,N_8850);
nand U10476 (N_10476,N_7671,N_8014);
nor U10477 (N_10477,N_8781,N_8458);
xnor U10478 (N_10478,N_7677,N_7737);
xor U10479 (N_10479,N_8705,N_8726);
xor U10480 (N_10480,N_8693,N_8045);
and U10481 (N_10481,N_8956,N_7965);
nand U10482 (N_10482,N_7786,N_7720);
xnor U10483 (N_10483,N_7898,N_7836);
or U10484 (N_10484,N_7618,N_8446);
nand U10485 (N_10485,N_7780,N_8801);
nand U10486 (N_10486,N_8158,N_8273);
nor U10487 (N_10487,N_8809,N_7858);
nor U10488 (N_10488,N_8113,N_8989);
xnor U10489 (N_10489,N_7774,N_8300);
or U10490 (N_10490,N_8596,N_8443);
nand U10491 (N_10491,N_8719,N_8153);
or U10492 (N_10492,N_8369,N_8013);
xnor U10493 (N_10493,N_8201,N_8588);
and U10494 (N_10494,N_8353,N_7723);
nand U10495 (N_10495,N_8824,N_8686);
nand U10496 (N_10496,N_8762,N_8558);
nor U10497 (N_10497,N_8833,N_8525);
nand U10498 (N_10498,N_8720,N_7979);
and U10499 (N_10499,N_8501,N_7740);
xor U10500 (N_10500,N_10207,N_9245);
nand U10501 (N_10501,N_9046,N_9005);
nor U10502 (N_10502,N_9431,N_10410);
xor U10503 (N_10503,N_9669,N_9800);
or U10504 (N_10504,N_9704,N_10067);
or U10505 (N_10505,N_9138,N_9938);
or U10506 (N_10506,N_10461,N_9838);
and U10507 (N_10507,N_9296,N_10448);
nand U10508 (N_10508,N_9775,N_10333);
nand U10509 (N_10509,N_9678,N_10418);
nand U10510 (N_10510,N_9128,N_10476);
and U10511 (N_10511,N_10271,N_10364);
nand U10512 (N_10512,N_10016,N_9489);
xnor U10513 (N_10513,N_9780,N_9386);
xor U10514 (N_10514,N_9546,N_9663);
nand U10515 (N_10515,N_9793,N_10171);
xor U10516 (N_10516,N_9873,N_10345);
or U10517 (N_10517,N_10199,N_9496);
nor U10518 (N_10518,N_10085,N_9284);
xnor U10519 (N_10519,N_9575,N_10146);
xnor U10520 (N_10520,N_10111,N_9200);
xor U10521 (N_10521,N_9139,N_10323);
and U10522 (N_10522,N_10373,N_10482);
and U10523 (N_10523,N_9685,N_9957);
xnor U10524 (N_10524,N_9734,N_9751);
xor U10525 (N_10525,N_9494,N_10175);
nor U10526 (N_10526,N_9184,N_9833);
or U10527 (N_10527,N_10159,N_10494);
xor U10528 (N_10528,N_9151,N_9823);
nor U10529 (N_10529,N_9287,N_10102);
and U10530 (N_10530,N_10413,N_9075);
and U10531 (N_10531,N_10001,N_10121);
nand U10532 (N_10532,N_9047,N_10213);
or U10533 (N_10533,N_9541,N_9760);
nor U10534 (N_10534,N_10335,N_9480);
nand U10535 (N_10535,N_9478,N_10267);
or U10536 (N_10536,N_9518,N_9629);
or U10537 (N_10537,N_10491,N_9658);
or U10538 (N_10538,N_9469,N_10361);
nor U10539 (N_10539,N_10412,N_9730);
and U10540 (N_10540,N_9032,N_9285);
and U10541 (N_10541,N_9656,N_9363);
nor U10542 (N_10542,N_9746,N_10354);
nor U10543 (N_10543,N_9310,N_10210);
nand U10544 (N_10544,N_10318,N_9269);
nor U10545 (N_10545,N_9053,N_9410);
xnor U10546 (N_10546,N_9272,N_9871);
and U10547 (N_10547,N_9670,N_9112);
or U10548 (N_10548,N_10157,N_10309);
xor U10549 (N_10549,N_10201,N_9655);
xor U10550 (N_10550,N_9812,N_9198);
xor U10551 (N_10551,N_10303,N_9117);
nor U10552 (N_10552,N_10208,N_10156);
or U10553 (N_10553,N_9065,N_10088);
and U10554 (N_10554,N_9179,N_9796);
and U10555 (N_10555,N_9896,N_10368);
or U10556 (N_10556,N_10116,N_10093);
nand U10557 (N_10557,N_10423,N_10465);
and U10558 (N_10558,N_9461,N_9076);
xnor U10559 (N_10559,N_9440,N_9766);
and U10560 (N_10560,N_9512,N_9609);
nor U10561 (N_10561,N_9264,N_9343);
nand U10562 (N_10562,N_10438,N_9149);
nor U10563 (N_10563,N_9853,N_10339);
xor U10564 (N_10564,N_10139,N_10185);
or U10565 (N_10565,N_9974,N_10141);
nor U10566 (N_10566,N_10252,N_9216);
xor U10567 (N_10567,N_9167,N_9523);
xor U10568 (N_10568,N_10084,N_9289);
nor U10569 (N_10569,N_9391,N_9166);
and U10570 (N_10570,N_9207,N_9246);
nor U10571 (N_10571,N_9733,N_9722);
nor U10572 (N_10572,N_9868,N_9037);
and U10573 (N_10573,N_10394,N_9735);
and U10574 (N_10574,N_9606,N_10051);
nand U10575 (N_10575,N_9031,N_10120);
nor U10576 (N_10576,N_10038,N_10444);
and U10577 (N_10577,N_9615,N_9499);
xor U10578 (N_10578,N_9181,N_9333);
nand U10579 (N_10579,N_9651,N_10115);
nor U10580 (N_10580,N_10162,N_9732);
nor U10581 (N_10581,N_9068,N_10399);
xor U10582 (N_10582,N_9716,N_10452);
and U10583 (N_10583,N_9306,N_9807);
or U10584 (N_10584,N_9073,N_9249);
or U10585 (N_10585,N_10459,N_9015);
xnor U10586 (N_10586,N_9404,N_9254);
nor U10587 (N_10587,N_9842,N_9966);
nand U10588 (N_10588,N_10401,N_10429);
and U10589 (N_10589,N_9094,N_9026);
and U10590 (N_10590,N_9729,N_9811);
nor U10591 (N_10591,N_9994,N_10225);
nand U10592 (N_10592,N_10166,N_9418);
nor U10593 (N_10593,N_9758,N_9805);
and U10594 (N_10594,N_9750,N_10173);
or U10595 (N_10595,N_9185,N_9761);
nor U10596 (N_10596,N_9215,N_10384);
xnor U10597 (N_10597,N_9486,N_10163);
or U10598 (N_10598,N_9498,N_10081);
nand U10599 (N_10599,N_9755,N_9612);
nand U10600 (N_10600,N_9454,N_10238);
nand U10601 (N_10601,N_10376,N_9959);
nand U10602 (N_10602,N_9382,N_9532);
nor U10603 (N_10603,N_10348,N_10018);
nor U10604 (N_10604,N_9859,N_9262);
nand U10605 (N_10605,N_9998,N_9725);
nor U10606 (N_10606,N_9432,N_9781);
and U10607 (N_10607,N_10231,N_9282);
xnor U10608 (N_10608,N_9594,N_9338);
or U10609 (N_10609,N_10234,N_9302);
or U10610 (N_10610,N_9401,N_9061);
and U10611 (N_10611,N_9243,N_9949);
xnor U10612 (N_10612,N_10206,N_9370);
nor U10613 (N_10613,N_10239,N_9411);
nand U10614 (N_10614,N_10241,N_9836);
xor U10615 (N_10615,N_10181,N_10420);
xnor U10616 (N_10616,N_10196,N_9280);
nand U10617 (N_10617,N_9014,N_10472);
or U10618 (N_10618,N_9535,N_9027);
and U10619 (N_10619,N_9011,N_9673);
xnor U10620 (N_10620,N_9964,N_9039);
and U10621 (N_10621,N_9196,N_9968);
and U10622 (N_10622,N_9118,N_10408);
and U10623 (N_10623,N_9267,N_10477);
xor U10624 (N_10624,N_9681,N_9520);
and U10625 (N_10625,N_9174,N_10300);
xor U10626 (N_10626,N_9795,N_10349);
and U10627 (N_10627,N_9709,N_10086);
nand U10628 (N_10628,N_10402,N_9617);
nand U10629 (N_10629,N_9036,N_10365);
xor U10630 (N_10630,N_9855,N_9740);
nand U10631 (N_10631,N_9915,N_9721);
xnor U10632 (N_10632,N_10106,N_10329);
nand U10633 (N_10633,N_10257,N_9345);
nor U10634 (N_10634,N_9893,N_9872);
xnor U10635 (N_10635,N_10277,N_9955);
nand U10636 (N_10636,N_9195,N_10460);
and U10637 (N_10637,N_9506,N_10062);
or U10638 (N_10638,N_10489,N_10462);
or U10639 (N_10639,N_9259,N_9038);
and U10640 (N_10640,N_9420,N_9258);
xor U10641 (N_10641,N_10190,N_9281);
xnor U10642 (N_10642,N_9274,N_10114);
and U10643 (N_10643,N_9419,N_9475);
or U10644 (N_10644,N_9500,N_10385);
or U10645 (N_10645,N_9328,N_9144);
nand U10646 (N_10646,N_9143,N_9637);
nor U10647 (N_10647,N_9803,N_9407);
nand U10648 (N_10648,N_10336,N_9979);
nor U10649 (N_10649,N_10055,N_9801);
xor U10650 (N_10650,N_9388,N_9712);
nor U10651 (N_10651,N_9764,N_9205);
nor U10652 (N_10652,N_9771,N_9313);
nor U10653 (N_10653,N_10097,N_10312);
xor U10654 (N_10654,N_9720,N_10321);
nor U10655 (N_10655,N_9577,N_9986);
or U10656 (N_10656,N_9164,N_10050);
or U10657 (N_10657,N_10296,N_9778);
nand U10658 (N_10658,N_10355,N_9409);
nand U10659 (N_10659,N_9349,N_9161);
nand U10660 (N_10660,N_9028,N_9643);
and U10661 (N_10661,N_9129,N_10029);
nor U10662 (N_10662,N_9747,N_9408);
nand U10663 (N_10663,N_9157,N_9318);
and U10664 (N_10664,N_9277,N_9589);
nor U10665 (N_10665,N_9371,N_10442);
or U10666 (N_10666,N_9443,N_10005);
xnor U10667 (N_10667,N_9999,N_10256);
nor U10668 (N_10668,N_9621,N_9858);
or U10669 (N_10669,N_10367,N_9237);
xnor U10670 (N_10670,N_10428,N_9692);
nor U10671 (N_10671,N_9828,N_10202);
nand U10672 (N_10672,N_10306,N_9946);
nand U10673 (N_10673,N_9743,N_9696);
or U10674 (N_10674,N_10127,N_10248);
nor U10675 (N_10675,N_10052,N_10200);
nor U10676 (N_10676,N_9360,N_10073);
and U10677 (N_10677,N_10470,N_9152);
xnor U10678 (N_10678,N_10466,N_9070);
nand U10679 (N_10679,N_9001,N_9742);
and U10680 (N_10680,N_10311,N_9002);
and U10681 (N_10681,N_9922,N_9201);
nand U10682 (N_10682,N_9912,N_9482);
nand U10683 (N_10683,N_9741,N_10341);
nor U10684 (N_10684,N_10059,N_10144);
and U10685 (N_10685,N_9556,N_9422);
xor U10686 (N_10686,N_9774,N_10104);
xor U10687 (N_10687,N_9885,N_10135);
nor U10688 (N_10688,N_10362,N_10356);
nor U10689 (N_10689,N_9104,N_9517);
nor U10690 (N_10690,N_10289,N_10165);
nor U10691 (N_10691,N_9794,N_9162);
xor U10692 (N_10692,N_9081,N_10358);
xnor U10693 (N_10693,N_9314,N_9867);
and U10694 (N_10694,N_9942,N_10126);
nor U10695 (N_10695,N_10150,N_9777);
and U10696 (N_10696,N_9640,N_9448);
and U10697 (N_10697,N_9791,N_9403);
and U10698 (N_10698,N_9592,N_9693);
or U10699 (N_10699,N_10471,N_9736);
or U10700 (N_10700,N_9159,N_10077);
nand U10701 (N_10701,N_9114,N_9189);
xnor U10702 (N_10702,N_9103,N_9472);
xor U10703 (N_10703,N_9372,N_9940);
xor U10704 (N_10704,N_9210,N_9717);
and U10705 (N_10705,N_9286,N_9560);
or U10706 (N_10706,N_10147,N_9579);
and U10707 (N_10707,N_9214,N_9610);
xnor U10708 (N_10708,N_9158,N_10069);
xor U10709 (N_10709,N_10468,N_9248);
nor U10710 (N_10710,N_9533,N_10021);
and U10711 (N_10711,N_9822,N_10158);
and U10712 (N_10712,N_9485,N_9906);
nor U10713 (N_10713,N_10193,N_9133);
nor U10714 (N_10714,N_9030,N_10002);
nand U10715 (N_10715,N_10030,N_9645);
nand U10716 (N_10716,N_10124,N_10281);
and U10717 (N_10717,N_9559,N_9996);
nor U10718 (N_10718,N_9083,N_10143);
nor U10719 (N_10719,N_9902,N_10488);
nand U10720 (N_10720,N_9169,N_9235);
or U10721 (N_10721,N_9728,N_10273);
or U10722 (N_10722,N_9635,N_9653);
nand U10723 (N_10723,N_9695,N_9434);
nor U10724 (N_10724,N_9102,N_9706);
and U10725 (N_10725,N_10390,N_9035);
or U10726 (N_10726,N_9305,N_9564);
nand U10727 (N_10727,N_9659,N_10142);
or U10728 (N_10728,N_9087,N_10017);
or U10729 (N_10729,N_9462,N_9319);
nand U10730 (N_10730,N_10386,N_9298);
xnor U10731 (N_10731,N_10000,N_9897);
or U10732 (N_10732,N_10270,N_9111);
and U10733 (N_10733,N_10089,N_10262);
nand U10734 (N_10734,N_9191,N_9973);
nor U10735 (N_10735,N_10416,N_10109);
xor U10736 (N_10736,N_10222,N_9334);
and U10737 (N_10737,N_9194,N_9596);
nand U10738 (N_10738,N_9519,N_9850);
and U10739 (N_10739,N_9347,N_10314);
nor U10740 (N_10740,N_9051,N_10205);
nand U10741 (N_10741,N_9991,N_9576);
or U10742 (N_10742,N_9505,N_9845);
or U10743 (N_10743,N_9782,N_10041);
nor U10744 (N_10744,N_10454,N_9753);
or U10745 (N_10745,N_10266,N_9240);
nand U10746 (N_10746,N_9394,N_9359);
xnor U10747 (N_10747,N_9012,N_9299);
nor U10748 (N_10748,N_9251,N_9187);
or U10749 (N_10749,N_9528,N_10083);
nor U10750 (N_10750,N_9808,N_9137);
xor U10751 (N_10751,N_9348,N_10176);
nor U10752 (N_10752,N_9894,N_9545);
and U10753 (N_10753,N_9447,N_9982);
nor U10754 (N_10754,N_9745,N_10149);
nor U10755 (N_10755,N_10337,N_9779);
xnor U10756 (N_10756,N_9424,N_9935);
or U10757 (N_10757,N_9204,N_9852);
or U10758 (N_10758,N_10322,N_10170);
or U10759 (N_10759,N_10483,N_10406);
or U10760 (N_10760,N_10285,N_9683);
nand U10761 (N_10761,N_9978,N_9837);
nand U10762 (N_10762,N_10422,N_9352);
nor U10763 (N_10763,N_9341,N_10112);
xnor U10764 (N_10764,N_10027,N_10434);
xor U10765 (N_10765,N_9713,N_10183);
or U10766 (N_10766,N_10148,N_9303);
xnor U10767 (N_10767,N_10046,N_9092);
nor U10768 (N_10768,N_9123,N_9444);
nor U10769 (N_10769,N_10226,N_9238);
and U10770 (N_10770,N_9355,N_9049);
nand U10771 (N_10771,N_9088,N_9947);
nor U10772 (N_10772,N_10079,N_10486);
nor U10773 (N_10773,N_9600,N_9776);
xnor U10774 (N_10774,N_9866,N_9358);
nor U10775 (N_10775,N_9936,N_9555);
or U10776 (N_10776,N_9367,N_9266);
or U10777 (N_10777,N_9402,N_10012);
or U10778 (N_10778,N_9430,N_10383);
nor U10779 (N_10779,N_9309,N_10229);
nand U10780 (N_10780,N_10119,N_9405);
nand U10781 (N_10781,N_9731,N_9628);
or U10782 (N_10782,N_9710,N_9748);
nand U10783 (N_10783,N_9458,N_9183);
or U10784 (N_10784,N_9043,N_9186);
or U10785 (N_10785,N_10048,N_9242);
or U10786 (N_10786,N_10179,N_9826);
xor U10787 (N_10787,N_10375,N_10198);
xor U10788 (N_10788,N_9718,N_9160);
and U10789 (N_10789,N_10265,N_9105);
nand U10790 (N_10790,N_9626,N_9881);
xor U10791 (N_10791,N_9672,N_9539);
nor U10792 (N_10792,N_10094,N_9311);
xor U10793 (N_10793,N_9300,N_9086);
or U10794 (N_10794,N_9236,N_9326);
nor U10795 (N_10795,N_9346,N_9876);
or U10796 (N_10796,N_9260,N_10223);
nor U10797 (N_10797,N_9737,N_9513);
or U10798 (N_10798,N_9292,N_10426);
nor U10799 (N_10799,N_9377,N_9271);
or U10800 (N_10800,N_9297,N_9965);
and U10801 (N_10801,N_9985,N_9983);
or U10802 (N_10802,N_10324,N_10437);
or U10803 (N_10803,N_10327,N_9707);
or U10804 (N_10804,N_9381,N_9180);
xnor U10805 (N_10805,N_9754,N_10007);
and U10806 (N_10806,N_10319,N_9090);
nor U10807 (N_10807,N_9213,N_9414);
and U10808 (N_10808,N_10174,N_10122);
nor U10809 (N_10809,N_9903,N_9016);
xnor U10810 (N_10810,N_9079,N_9464);
nor U10811 (N_10811,N_9784,N_10317);
nand U10812 (N_10812,N_10431,N_10009);
nand U10813 (N_10813,N_9182,N_9572);
xor U10814 (N_10814,N_9724,N_9665);
xnor U10815 (N_10815,N_9193,N_9082);
and U10816 (N_10816,N_9085,N_9293);
nor U10817 (N_10817,N_9586,N_9602);
nand U10818 (N_10818,N_10216,N_9603);
or U10819 (N_10819,N_9723,N_9132);
nand U10820 (N_10820,N_10136,N_10090);
xnor U10821 (N_10821,N_9768,N_9497);
or U10822 (N_10822,N_10182,N_9757);
nor U10823 (N_10823,N_10308,N_9374);
nand U10824 (N_10824,N_9142,N_9060);
nor U10825 (N_10825,N_10405,N_9883);
and U10826 (N_10826,N_9316,N_10260);
or U10827 (N_10827,N_10215,N_9763);
and U10828 (N_10828,N_10293,N_9294);
nor U10829 (N_10829,N_9887,N_9041);
xnor U10830 (N_10830,N_9437,N_9633);
or U10831 (N_10831,N_9146,N_9176);
or U10832 (N_10832,N_9054,N_9932);
nand U10833 (N_10833,N_9997,N_9165);
nor U10834 (N_10834,N_9385,N_10425);
xnor U10835 (N_10835,N_9702,N_9990);
nor U10836 (N_10836,N_9632,N_9923);
xnor U10837 (N_10837,N_9574,N_9003);
or U10838 (N_10838,N_9767,N_10279);
nand U10839 (N_10839,N_9429,N_9045);
nor U10840 (N_10840,N_9916,N_10137);
and U10841 (N_10841,N_9765,N_9098);
or U10842 (N_10842,N_9809,N_9154);
nor U10843 (N_10843,N_9066,N_9379);
or U10844 (N_10844,N_9905,N_9749);
or U10845 (N_10845,N_9770,N_9023);
nand U10846 (N_10846,N_9125,N_9178);
or U10847 (N_10847,N_9821,N_9911);
and U10848 (N_10848,N_10160,N_10499);
and U10849 (N_10849,N_10230,N_9329);
xor U10850 (N_10850,N_9988,N_9890);
nor U10851 (N_10851,N_9846,N_10212);
and U10852 (N_10852,N_9554,N_9368);
nand U10853 (N_10853,N_9017,N_9703);
nand U10854 (N_10854,N_10228,N_9566);
nor U10855 (N_10855,N_9400,N_9477);
xnor U10856 (N_10856,N_10435,N_9057);
nand U10857 (N_10857,N_9799,N_10024);
or U10858 (N_10858,N_9342,N_9854);
nor U10859 (N_10859,N_10350,N_9558);
and U10860 (N_10860,N_9416,N_10474);
or U10861 (N_10861,N_10473,N_10129);
and U10862 (N_10862,N_9279,N_10363);
and U10863 (N_10863,N_9206,N_9727);
xor U10864 (N_10864,N_9050,N_10071);
and U10865 (N_10865,N_9843,N_9888);
or U10866 (N_10866,N_10145,N_10113);
and U10867 (N_10867,N_10269,N_10334);
nor U10868 (N_10868,N_9536,N_10065);
xor U10869 (N_10869,N_9177,N_9530);
nor U10870 (N_10870,N_9217,N_10186);
nor U10871 (N_10871,N_9642,N_9276);
nand U10872 (N_10872,N_9832,N_10332);
and U10873 (N_10873,N_9492,N_10161);
nor U10874 (N_10874,N_9413,N_10152);
and U10875 (N_10875,N_9317,N_9992);
nand U10876 (N_10876,N_9627,N_9790);
nor U10877 (N_10877,N_9202,N_9056);
or U10878 (N_10878,N_9892,N_10495);
and U10879 (N_10879,N_9582,N_10404);
nor U10880 (N_10880,N_9759,N_9847);
nand U10881 (N_10881,N_9229,N_10484);
or U10882 (N_10882,N_9361,N_9662);
or U10883 (N_10883,N_10338,N_9397);
nor U10884 (N_10884,N_10302,N_9975);
xnor U10885 (N_10885,N_10087,N_10091);
and U10886 (N_10886,N_9101,N_10283);
nor U10887 (N_10887,N_9290,N_9726);
nor U10888 (N_10888,N_10249,N_10344);
nor U10889 (N_10889,N_9212,N_9584);
nand U10890 (N_10890,N_9926,N_9463);
nand U10891 (N_10891,N_9813,N_9525);
xnor U10892 (N_10892,N_10037,N_9667);
or U10893 (N_10893,N_10400,N_9884);
and U10894 (N_10894,N_10110,N_9072);
nor U10895 (N_10895,N_10360,N_9147);
or U10896 (N_10896,N_9719,N_9550);
nand U10897 (N_10897,N_10315,N_9288);
nor U10898 (N_10898,N_9354,N_9442);
and U10899 (N_10899,N_9487,N_9918);
or U10900 (N_10900,N_9421,N_9451);
nor U10901 (N_10901,N_9583,N_9022);
nor U10902 (N_10902,N_10020,N_9715);
nand U10903 (N_10903,N_9131,N_9963);
or U10904 (N_10904,N_9452,N_10282);
xnor U10905 (N_10905,N_9450,N_9508);
xor U10906 (N_10906,N_9886,N_9007);
nand U10907 (N_10907,N_10330,N_9543);
or U10908 (N_10908,N_9917,N_9676);
and U10909 (N_10909,N_10347,N_10264);
and U10910 (N_10910,N_9699,N_9537);
and U10911 (N_10911,N_10047,N_9484);
xor U10912 (N_10912,N_10388,N_9531);
and U10913 (N_10913,N_9616,N_10236);
nor U10914 (N_10914,N_9898,N_9362);
nor U10915 (N_10915,N_9364,N_9563);
xnor U10916 (N_10916,N_10105,N_9869);
xnor U10917 (N_10917,N_9106,N_9226);
nor U10918 (N_10918,N_9369,N_10025);
xnor U10919 (N_10919,N_10439,N_9383);
nor U10920 (N_10920,N_9124,N_9814);
or U10921 (N_10921,N_10353,N_9829);
nand U10922 (N_10922,N_9199,N_10251);
and U10923 (N_10923,N_9456,N_10214);
or U10924 (N_10924,N_10481,N_10006);
nand U10925 (N_10925,N_10301,N_9009);
nor U10926 (N_10926,N_9446,N_9396);
and U10927 (N_10927,N_9470,N_9445);
nor U10928 (N_10928,N_9690,N_9646);
and U10929 (N_10929,N_9827,N_9067);
nand U10930 (N_10930,N_9504,N_10023);
xnor U10931 (N_10931,N_9211,N_10427);
and U10932 (N_10932,N_10445,N_9581);
nand U10933 (N_10933,N_9514,N_9618);
or U10934 (N_10934,N_9415,N_9995);
or U10935 (N_10935,N_9700,N_9173);
xnor U10936 (N_10936,N_9686,N_9126);
nor U10937 (N_10937,N_10053,N_9654);
nor U10938 (N_10938,N_9588,N_10366);
and U10939 (N_10939,N_9590,N_9561);
xnor U10940 (N_10940,N_10022,N_9671);
nor U10941 (N_10941,N_10204,N_9772);
and U10942 (N_10942,N_9527,N_9320);
and U10943 (N_10943,N_9605,N_9516);
nor U10944 (N_10944,N_9325,N_9952);
or U10945 (N_10945,N_9900,N_9789);
nor U10946 (N_10946,N_9029,N_9473);
and U10947 (N_10947,N_9908,N_10187);
or U10948 (N_10948,N_9096,N_10192);
or U10949 (N_10949,N_9380,N_9426);
xnor U10950 (N_10950,N_9077,N_9939);
and U10951 (N_10951,N_10058,N_9384);
nand U10952 (N_10952,N_10443,N_10057);
nand U10953 (N_10953,N_10235,N_9153);
xor U10954 (N_10954,N_9666,N_9944);
or U10955 (N_10955,N_10064,N_9816);
and U10956 (N_10956,N_9870,N_9353);
or U10957 (N_10957,N_10132,N_9471);
or U10958 (N_10958,N_9636,N_9684);
and U10959 (N_10959,N_9930,N_10253);
and U10960 (N_10960,N_10151,N_9878);
nand U10961 (N_10961,N_10272,N_10209);
or U10962 (N_10962,N_9503,N_9481);
nand U10963 (N_10963,N_9427,N_9483);
or U10964 (N_10964,N_9048,N_10294);
nor U10965 (N_10965,N_9108,N_9175);
nand U10966 (N_10966,N_9967,N_9792);
or U10967 (N_10967,N_9257,N_10032);
nor U10968 (N_10968,N_9951,N_9308);
nor U10969 (N_10969,N_9324,N_10117);
and U10970 (N_10970,N_9219,N_10259);
nand U10971 (N_10971,N_9171,N_9406);
nor U10972 (N_10972,N_10374,N_9899);
nor U10973 (N_10973,N_10220,N_10343);
and U10974 (N_10974,N_9568,N_9679);
and U10975 (N_10975,N_9107,N_9232);
nor U10976 (N_10976,N_9392,N_9798);
and U10977 (N_10977,N_9378,N_10453);
xnor U10978 (N_10978,N_9804,N_10458);
or U10979 (N_10979,N_9802,N_9552);
and U10980 (N_10980,N_9649,N_9844);
and U10981 (N_10981,N_9501,N_9291);
and U10982 (N_10982,N_9275,N_10130);
and U10983 (N_10983,N_9895,N_9093);
nor U10984 (N_10984,N_10060,N_9019);
nand U10985 (N_10985,N_9247,N_9344);
or U10986 (N_10986,N_10154,N_9241);
and U10987 (N_10987,N_10153,N_9920);
nand U10988 (N_10988,N_10138,N_9190);
xor U10989 (N_10989,N_9295,N_10232);
or U10990 (N_10990,N_9479,N_10436);
nand U10991 (N_10991,N_10298,N_9981);
nor U10992 (N_10992,N_10326,N_9648);
nand U10993 (N_10993,N_10372,N_9849);
or U10994 (N_10994,N_9987,N_9033);
and U10995 (N_10995,N_9502,N_9835);
nor U10996 (N_10996,N_9860,N_9739);
nand U10997 (N_10997,N_9569,N_10242);
nand U10998 (N_10998,N_9925,N_9490);
xor U10999 (N_10999,N_10393,N_9954);
or U11000 (N_11000,N_9010,N_10134);
or U11001 (N_11001,N_9909,N_9650);
xnor U11002 (N_11002,N_9110,N_10325);
or U11003 (N_11003,N_9270,N_9071);
xnor U11004 (N_11004,N_10101,N_9620);
or U11005 (N_11005,N_9544,N_9021);
nor U11006 (N_11006,N_9425,N_10455);
xor U11007 (N_11007,N_9390,N_9253);
or U11008 (N_11008,N_10492,N_9675);
or U11009 (N_11009,N_9366,N_9595);
xnor U11010 (N_11010,N_10480,N_9914);
nor U11011 (N_11011,N_9064,N_10305);
xnor U11012 (N_11012,N_9668,N_9977);
nor U11013 (N_11013,N_10100,N_9697);
and U11014 (N_11014,N_9332,N_9208);
nor U11015 (N_11015,N_9433,N_9524);
or U11016 (N_11016,N_9453,N_10218);
nand U11017 (N_11017,N_9565,N_10240);
nand U11018 (N_11018,N_9788,N_9435);
nor U11019 (N_11019,N_10033,N_10098);
and U11020 (N_11020,N_10074,N_10003);
or U11021 (N_11021,N_9170,N_9080);
nand U11022 (N_11022,N_10013,N_9928);
nand U11023 (N_11023,N_10382,N_9412);
or U11024 (N_11024,N_10417,N_9542);
nor U11025 (N_11025,N_9488,N_9907);
or U11026 (N_11026,N_10040,N_9340);
nor U11027 (N_11027,N_9441,N_10340);
and U11028 (N_11028,N_9115,N_10221);
nand U11029 (N_11029,N_10072,N_9913);
or U11030 (N_11030,N_10015,N_9660);
and U11031 (N_11031,N_10061,N_9074);
nand U11032 (N_11032,N_10316,N_9336);
nand U11033 (N_11033,N_9958,N_9493);
and U11034 (N_11034,N_9323,N_9943);
xor U11035 (N_11035,N_10261,N_10432);
xor U11036 (N_11036,N_9356,N_10424);
nor U11037 (N_11037,N_9578,N_9910);
nand U11038 (N_11038,N_9580,N_10346);
nor U11039 (N_11039,N_9436,N_9919);
nand U11040 (N_11040,N_10082,N_9815);
nand U11041 (N_11041,N_9069,N_9273);
xnor U11042 (N_11042,N_9006,N_9122);
xor U11043 (N_11043,N_9607,N_10398);
nand U11044 (N_11044,N_9571,N_10133);
nand U11045 (N_11045,N_9634,N_9465);
or U11046 (N_11046,N_9630,N_10010);
nor U11047 (N_11047,N_9882,N_9817);
and U11048 (N_11048,N_9825,N_9099);
xor U11049 (N_11049,N_9034,N_9466);
and U11050 (N_11050,N_9593,N_9806);
or U11051 (N_11051,N_10463,N_9495);
and U11052 (N_11052,N_9130,N_10469);
nor U11053 (N_11053,N_9491,N_9962);
nand U11054 (N_11054,N_10457,N_9562);
xnor U11055 (N_11055,N_9841,N_9052);
nand U11056 (N_11056,N_9976,N_9283);
and U11057 (N_11057,N_9614,N_10189);
or U11058 (N_11058,N_9304,N_9155);
nand U11059 (N_11059,N_10419,N_9119);
nand U11060 (N_11060,N_9399,N_9971);
or U11061 (N_11061,N_9197,N_9769);
xor U11062 (N_11062,N_10286,N_9188);
or U11063 (N_11063,N_10044,N_10250);
nor U11064 (N_11064,N_9339,N_9682);
and U11065 (N_11065,N_9510,N_9192);
nand U11066 (N_11066,N_9134,N_10275);
xnor U11067 (N_11067,N_9989,N_10255);
nor U11068 (N_11068,N_9387,N_9861);
and U11069 (N_11069,N_9234,N_9687);
nand U11070 (N_11070,N_9570,N_9953);
or U11071 (N_11071,N_10245,N_10403);
and U11072 (N_11072,N_9058,N_10172);
xor U11073 (N_11073,N_10194,N_10219);
or U11074 (N_11074,N_10396,N_9830);
xnor U11075 (N_11075,N_9708,N_9148);
xor U11076 (N_11076,N_9127,N_9145);
or U11077 (N_11077,N_9889,N_9222);
nand U11078 (N_11078,N_9831,N_9095);
nand U11079 (N_11079,N_9820,N_9711);
or U11080 (N_11080,N_10369,N_9141);
nand U11081 (N_11081,N_10080,N_9877);
and U11082 (N_11082,N_9457,N_9657);
xor U11083 (N_11083,N_9549,N_9529);
or U11084 (N_11084,N_9927,N_10357);
nor U11085 (N_11085,N_9857,N_9714);
nand U11086 (N_11086,N_10066,N_9762);
and U11087 (N_11087,N_10167,N_9376);
nor U11088 (N_11088,N_10421,N_9455);
xnor U11089 (N_11089,N_10411,N_9331);
xor U11090 (N_11090,N_10395,N_10407);
xnor U11091 (N_11091,N_9389,N_10378);
or U11092 (N_11092,N_9970,N_9357);
nand U11093 (N_11093,N_9140,N_9934);
nor U11094 (N_11094,N_10274,N_9203);
nor U11095 (N_11095,N_10034,N_10475);
nand U11096 (N_11096,N_9515,N_10075);
and U11097 (N_11097,N_9335,N_10031);
and U11098 (N_11098,N_10042,N_9945);
or U11099 (N_11099,N_10479,N_9078);
nor U11100 (N_11100,N_10244,N_9921);
nor U11101 (N_11101,N_10379,N_9937);
nor U11102 (N_11102,N_9252,N_9221);
nor U11103 (N_11103,N_10451,N_9459);
nand U11104 (N_11104,N_9862,N_9268);
nand U11105 (N_11105,N_9557,N_10096);
nand U11106 (N_11106,N_10370,N_10387);
and U11107 (N_11107,N_9752,N_9109);
or U11108 (N_11108,N_10180,N_10276);
xnor U11109 (N_11109,N_9611,N_9661);
nand U11110 (N_11110,N_9423,N_10039);
or U11111 (N_11111,N_9100,N_10237);
nor U11112 (N_11112,N_9929,N_9691);
nand U11113 (N_11113,N_9865,N_9969);
nand U11114 (N_11114,N_9063,N_9008);
nand U11115 (N_11115,N_10191,N_9786);
xor U11116 (N_11116,N_9321,N_9522);
and U11117 (N_11117,N_9688,N_10246);
nor U11118 (N_11118,N_9467,N_9624);
xnor U11119 (N_11119,N_9756,N_10076);
xor U11120 (N_11120,N_10140,N_9819);
and U11121 (N_11121,N_9136,N_10043);
nor U11122 (N_11122,N_9228,N_10128);
xor U11123 (N_11123,N_9623,N_9567);
nor U11124 (N_11124,N_10278,N_9025);
and U11125 (N_11125,N_9834,N_9664);
and U11126 (N_11126,N_9880,N_9224);
nor U11127 (N_11127,N_10496,N_9024);
and U11128 (N_11128,N_9647,N_9573);
and U11129 (N_11129,N_9044,N_9091);
and U11130 (N_11130,N_10184,N_9225);
nor U11131 (N_11131,N_9449,N_10415);
and U11132 (N_11132,N_10054,N_10299);
xnor U11133 (N_11133,N_9172,N_10280);
xnor U11134 (N_11134,N_9000,N_10290);
nand U11135 (N_11135,N_10485,N_9652);
nand U11136 (N_11136,N_9972,N_9476);
or U11137 (N_11137,N_10168,N_9312);
and U11138 (N_11138,N_9585,N_9738);
or U11139 (N_11139,N_9840,N_9534);
nor U11140 (N_11140,N_9393,N_9587);
or U11141 (N_11141,N_9120,N_10493);
xor U11142 (N_11142,N_9698,N_9601);
or U11143 (N_11143,N_9511,N_9322);
nor U11144 (N_11144,N_9810,N_9933);
nand U11145 (N_11145,N_9604,N_10011);
or U11146 (N_11146,N_9507,N_9255);
nor U11147 (N_11147,N_9961,N_10320);
xnor U11148 (N_11148,N_10447,N_10092);
nor U11149 (N_11149,N_9680,N_10095);
xor U11150 (N_11150,N_10103,N_9265);
nand U11151 (N_11151,N_9055,N_9641);
nor U11152 (N_11152,N_9327,N_9230);
nand U11153 (N_11153,N_9597,N_9787);
and U11154 (N_11154,N_10233,N_10389);
xor U11155 (N_11155,N_9851,N_9350);
nor U11156 (N_11156,N_10307,N_9218);
nand U11157 (N_11157,N_9818,N_9622);
nand U11158 (N_11158,N_9980,N_9156);
or U11159 (N_11159,N_9315,N_10391);
and U11160 (N_11160,N_10108,N_10328);
xnor U11161 (N_11161,N_10178,N_10440);
nand U11162 (N_11162,N_10441,N_9398);
nor U11163 (N_11163,N_9956,N_10297);
xnor U11164 (N_11164,N_10211,N_10292);
nor U11165 (N_11165,N_9783,N_9864);
and U11166 (N_11166,N_9931,N_10456);
nor U11167 (N_11167,N_9301,N_9365);
and U11168 (N_11168,N_9891,N_10263);
and U11169 (N_11169,N_9018,N_9163);
nor U11170 (N_11170,N_9351,N_10414);
nand U11171 (N_11171,N_9839,N_10028);
nand U11172 (N_11172,N_10310,N_9705);
and U11173 (N_11173,N_10291,N_10392);
xnor U11174 (N_11174,N_9089,N_10254);
and U11175 (N_11175,N_9209,N_9644);
nand U11176 (N_11176,N_10304,N_9875);
xnor U11177 (N_11177,N_9548,N_9428);
nand U11178 (N_11178,N_9168,N_9468);
xnor U11179 (N_11179,N_10351,N_10014);
nand U11180 (N_11180,N_10243,N_9042);
xor U11181 (N_11181,N_9040,N_9261);
xnor U11182 (N_11182,N_10331,N_10131);
nor U11183 (N_11183,N_9677,N_9744);
nand U11184 (N_11184,N_10478,N_10026);
and U11185 (N_11185,N_10045,N_9638);
nor U11186 (N_11186,N_9256,N_9941);
xor U11187 (N_11187,N_9375,N_10450);
xnor U11188 (N_11188,N_9509,N_9135);
nand U11189 (N_11189,N_10446,N_9223);
and U11190 (N_11190,N_9474,N_10078);
nand U11191 (N_11191,N_10188,N_9395);
xor U11192 (N_11192,N_10004,N_10224);
nor U11193 (N_11193,N_10008,N_9113);
nand U11194 (N_11194,N_10380,N_10123);
nand U11195 (N_11195,N_10464,N_10498);
nand U11196 (N_11196,N_9121,N_9984);
xnor U11197 (N_11197,N_9797,N_10371);
and U11198 (N_11198,N_10227,N_9020);
xor U11199 (N_11199,N_9639,N_9417);
nor U11200 (N_11200,N_10107,N_9373);
nor U11201 (N_11201,N_9608,N_10247);
nor U11202 (N_11202,N_9538,N_9553);
nor U11203 (N_11203,N_9619,N_9591);
nand U11204 (N_11204,N_9521,N_10433);
nand U11205 (N_11205,N_10099,N_10467);
xor U11206 (N_11206,N_9701,N_9250);
xnor U11207 (N_11207,N_9337,N_9773);
nor U11208 (N_11208,N_9960,N_9674);
xor U11209 (N_11209,N_10352,N_9863);
nor U11210 (N_11210,N_9239,N_9278);
xnor U11211 (N_11211,N_9004,N_9785);
or U11212 (N_11212,N_9244,N_10258);
and U11213 (N_11213,N_9948,N_10049);
or U11214 (N_11214,N_9150,N_10164);
nand U11215 (N_11215,N_9848,N_9220);
or U11216 (N_11216,N_9059,N_9526);
and U11217 (N_11217,N_9824,N_9993);
and U11218 (N_11218,N_9547,N_10155);
xnor U11219 (N_11219,N_9540,N_9013);
nor U11220 (N_11220,N_9233,N_9307);
or U11221 (N_11221,N_10490,N_10169);
nor U11222 (N_11222,N_10035,N_10056);
and U11223 (N_11223,N_9263,N_10359);
xor U11224 (N_11224,N_10203,N_10036);
nor U11225 (N_11225,N_10068,N_9116);
xnor U11226 (N_11226,N_10288,N_9694);
nor U11227 (N_11227,N_10118,N_10295);
or U11228 (N_11228,N_9613,N_10287);
or U11229 (N_11229,N_10197,N_9625);
nand U11230 (N_11230,N_10449,N_10487);
xor U11231 (N_11231,N_10377,N_10430);
xnor U11232 (N_11232,N_9438,N_9062);
nand U11233 (N_11233,N_9330,N_9460);
nand U11234 (N_11234,N_10019,N_10342);
or U11235 (N_11235,N_10268,N_10195);
or U11236 (N_11236,N_10409,N_9689);
nor U11237 (N_11237,N_9551,N_9950);
xnor U11238 (N_11238,N_9856,N_9598);
nor U11239 (N_11239,N_9904,N_9924);
nor U11240 (N_11240,N_9901,N_9439);
nor U11241 (N_11241,N_10177,N_10397);
or U11242 (N_11242,N_10313,N_9874);
xor U11243 (N_11243,N_10063,N_9227);
nor U11244 (N_11244,N_9879,N_9631);
and U11245 (N_11245,N_10125,N_10284);
nand U11246 (N_11246,N_9599,N_10381);
nand U11247 (N_11247,N_10070,N_9084);
nor U11248 (N_11248,N_9097,N_10497);
xor U11249 (N_11249,N_10217,N_9231);
xor U11250 (N_11250,N_10374,N_9837);
nor U11251 (N_11251,N_9941,N_10289);
and U11252 (N_11252,N_9203,N_9550);
or U11253 (N_11253,N_9924,N_9524);
and U11254 (N_11254,N_10299,N_9695);
nor U11255 (N_11255,N_10000,N_9379);
nor U11256 (N_11256,N_10085,N_10491);
or U11257 (N_11257,N_9214,N_9868);
and U11258 (N_11258,N_10066,N_10113);
xnor U11259 (N_11259,N_10035,N_9485);
xnor U11260 (N_11260,N_9791,N_9341);
and U11261 (N_11261,N_9694,N_10376);
nor U11262 (N_11262,N_10282,N_9799);
and U11263 (N_11263,N_9320,N_9966);
and U11264 (N_11264,N_10290,N_9370);
xor U11265 (N_11265,N_9879,N_9277);
nor U11266 (N_11266,N_9733,N_9486);
nand U11267 (N_11267,N_9557,N_9212);
and U11268 (N_11268,N_9659,N_10407);
or U11269 (N_11269,N_10124,N_9980);
nand U11270 (N_11270,N_10456,N_9077);
xnor U11271 (N_11271,N_9060,N_10021);
nor U11272 (N_11272,N_10154,N_9897);
nand U11273 (N_11273,N_10455,N_9341);
and U11274 (N_11274,N_10097,N_9673);
and U11275 (N_11275,N_9162,N_10121);
nor U11276 (N_11276,N_9937,N_9091);
or U11277 (N_11277,N_9449,N_9535);
nand U11278 (N_11278,N_9948,N_9494);
nor U11279 (N_11279,N_10088,N_9823);
nand U11280 (N_11280,N_10063,N_10202);
nand U11281 (N_11281,N_9534,N_9166);
nor U11282 (N_11282,N_9828,N_10168);
nor U11283 (N_11283,N_10201,N_9061);
nor U11284 (N_11284,N_9711,N_9456);
xor U11285 (N_11285,N_10033,N_9672);
and U11286 (N_11286,N_10038,N_10006);
xor U11287 (N_11287,N_9669,N_9618);
or U11288 (N_11288,N_9604,N_9374);
nand U11289 (N_11289,N_9663,N_10383);
or U11290 (N_11290,N_10160,N_10266);
nand U11291 (N_11291,N_10020,N_9312);
nor U11292 (N_11292,N_9169,N_9878);
nor U11293 (N_11293,N_10279,N_9088);
and U11294 (N_11294,N_10117,N_9561);
xor U11295 (N_11295,N_9356,N_9047);
nand U11296 (N_11296,N_9042,N_10030);
nand U11297 (N_11297,N_10238,N_9410);
nor U11298 (N_11298,N_10430,N_9451);
xnor U11299 (N_11299,N_9199,N_10404);
xor U11300 (N_11300,N_10431,N_9367);
or U11301 (N_11301,N_9321,N_9593);
or U11302 (N_11302,N_10421,N_9594);
nor U11303 (N_11303,N_9929,N_9888);
and U11304 (N_11304,N_9010,N_9717);
nor U11305 (N_11305,N_9036,N_9359);
nor U11306 (N_11306,N_9168,N_9633);
and U11307 (N_11307,N_9392,N_9241);
and U11308 (N_11308,N_9912,N_10327);
nor U11309 (N_11309,N_9898,N_9640);
xor U11310 (N_11310,N_10178,N_10080);
and U11311 (N_11311,N_9059,N_9238);
nor U11312 (N_11312,N_9912,N_9693);
and U11313 (N_11313,N_9222,N_9304);
and U11314 (N_11314,N_9156,N_10338);
nor U11315 (N_11315,N_9514,N_9360);
or U11316 (N_11316,N_10036,N_9646);
nand U11317 (N_11317,N_9123,N_9622);
xor U11318 (N_11318,N_10144,N_9017);
nor U11319 (N_11319,N_9717,N_9471);
nand U11320 (N_11320,N_9556,N_9365);
nor U11321 (N_11321,N_9009,N_9019);
nor U11322 (N_11322,N_9245,N_9393);
and U11323 (N_11323,N_9814,N_10407);
or U11324 (N_11324,N_9925,N_10294);
nand U11325 (N_11325,N_9619,N_9718);
nor U11326 (N_11326,N_9662,N_10089);
and U11327 (N_11327,N_9826,N_10095);
nand U11328 (N_11328,N_9113,N_9851);
xnor U11329 (N_11329,N_9268,N_9508);
nor U11330 (N_11330,N_9283,N_9117);
nor U11331 (N_11331,N_9583,N_9590);
and U11332 (N_11332,N_9338,N_10064);
and U11333 (N_11333,N_10233,N_9486);
nand U11334 (N_11334,N_9167,N_10292);
nand U11335 (N_11335,N_9825,N_9601);
xnor U11336 (N_11336,N_9563,N_9085);
and U11337 (N_11337,N_10114,N_10079);
nor U11338 (N_11338,N_9721,N_9396);
nor U11339 (N_11339,N_9837,N_9542);
and U11340 (N_11340,N_9190,N_10120);
nand U11341 (N_11341,N_9583,N_9175);
xnor U11342 (N_11342,N_10103,N_9499);
or U11343 (N_11343,N_9417,N_9452);
xnor U11344 (N_11344,N_10275,N_9635);
xor U11345 (N_11345,N_10442,N_10048);
nand U11346 (N_11346,N_9454,N_9238);
and U11347 (N_11347,N_9888,N_9477);
nor U11348 (N_11348,N_9662,N_9329);
or U11349 (N_11349,N_9836,N_10361);
or U11350 (N_11350,N_10211,N_9153);
xor U11351 (N_11351,N_10147,N_10361);
xnor U11352 (N_11352,N_9736,N_10307);
nand U11353 (N_11353,N_10043,N_9919);
or U11354 (N_11354,N_9689,N_10204);
or U11355 (N_11355,N_9663,N_9672);
nor U11356 (N_11356,N_10029,N_9972);
and U11357 (N_11357,N_9298,N_9290);
or U11358 (N_11358,N_9149,N_9074);
and U11359 (N_11359,N_10224,N_9982);
nor U11360 (N_11360,N_9057,N_9258);
nand U11361 (N_11361,N_10364,N_9588);
xor U11362 (N_11362,N_10133,N_9742);
and U11363 (N_11363,N_9180,N_9799);
xnor U11364 (N_11364,N_9520,N_9355);
or U11365 (N_11365,N_9567,N_9741);
and U11366 (N_11366,N_10425,N_10455);
xnor U11367 (N_11367,N_9169,N_10120);
xnor U11368 (N_11368,N_10059,N_9768);
nand U11369 (N_11369,N_9108,N_10008);
or U11370 (N_11370,N_10491,N_9442);
xor U11371 (N_11371,N_9560,N_9284);
or U11372 (N_11372,N_9748,N_9811);
nor U11373 (N_11373,N_10451,N_9896);
nor U11374 (N_11374,N_9238,N_10263);
nor U11375 (N_11375,N_9614,N_9393);
xor U11376 (N_11376,N_9767,N_10175);
nor U11377 (N_11377,N_9475,N_9942);
nor U11378 (N_11378,N_9769,N_9882);
and U11379 (N_11379,N_9242,N_9638);
nand U11380 (N_11380,N_9892,N_10253);
and U11381 (N_11381,N_10475,N_9998);
nand U11382 (N_11382,N_10349,N_9815);
or U11383 (N_11383,N_9929,N_9487);
nand U11384 (N_11384,N_9601,N_10253);
and U11385 (N_11385,N_10242,N_9603);
xor U11386 (N_11386,N_9621,N_9109);
nand U11387 (N_11387,N_9005,N_10051);
xnor U11388 (N_11388,N_9825,N_9261);
and U11389 (N_11389,N_9375,N_10045);
and U11390 (N_11390,N_9728,N_10306);
xor U11391 (N_11391,N_9116,N_9288);
or U11392 (N_11392,N_10246,N_10117);
nor U11393 (N_11393,N_9942,N_9883);
nand U11394 (N_11394,N_9392,N_9409);
nor U11395 (N_11395,N_10353,N_9161);
and U11396 (N_11396,N_10093,N_9048);
nand U11397 (N_11397,N_9184,N_9342);
nand U11398 (N_11398,N_9970,N_10337);
or U11399 (N_11399,N_10304,N_9237);
nor U11400 (N_11400,N_10258,N_10010);
and U11401 (N_11401,N_9115,N_10348);
or U11402 (N_11402,N_9068,N_9002);
xnor U11403 (N_11403,N_10305,N_9268);
xnor U11404 (N_11404,N_9483,N_9648);
xnor U11405 (N_11405,N_10382,N_9818);
or U11406 (N_11406,N_9958,N_9988);
nand U11407 (N_11407,N_9132,N_9615);
nand U11408 (N_11408,N_9452,N_9600);
nor U11409 (N_11409,N_10312,N_9249);
xnor U11410 (N_11410,N_9272,N_9768);
and U11411 (N_11411,N_9734,N_9041);
and U11412 (N_11412,N_9267,N_9833);
or U11413 (N_11413,N_10433,N_9301);
or U11414 (N_11414,N_9435,N_9776);
and U11415 (N_11415,N_10029,N_9506);
xor U11416 (N_11416,N_10311,N_10431);
or U11417 (N_11417,N_10296,N_9145);
nand U11418 (N_11418,N_9534,N_9038);
xnor U11419 (N_11419,N_10235,N_9640);
xnor U11420 (N_11420,N_9248,N_9638);
and U11421 (N_11421,N_10389,N_9864);
xnor U11422 (N_11422,N_9966,N_10249);
nor U11423 (N_11423,N_9027,N_10074);
xnor U11424 (N_11424,N_9705,N_10313);
and U11425 (N_11425,N_10474,N_10485);
xnor U11426 (N_11426,N_9656,N_10464);
nand U11427 (N_11427,N_9185,N_9123);
nand U11428 (N_11428,N_10278,N_10207);
and U11429 (N_11429,N_9076,N_9551);
nand U11430 (N_11430,N_9002,N_10329);
nand U11431 (N_11431,N_9099,N_9272);
nand U11432 (N_11432,N_9267,N_9484);
and U11433 (N_11433,N_9019,N_9817);
and U11434 (N_11434,N_10295,N_9270);
or U11435 (N_11435,N_9715,N_9018);
nor U11436 (N_11436,N_9160,N_9565);
xnor U11437 (N_11437,N_9250,N_9799);
and U11438 (N_11438,N_10417,N_9265);
nand U11439 (N_11439,N_9855,N_10360);
and U11440 (N_11440,N_10396,N_9964);
or U11441 (N_11441,N_10059,N_9704);
or U11442 (N_11442,N_9600,N_10090);
xnor U11443 (N_11443,N_9079,N_9223);
nor U11444 (N_11444,N_9781,N_10476);
nand U11445 (N_11445,N_9734,N_9694);
xor U11446 (N_11446,N_9154,N_9867);
xnor U11447 (N_11447,N_9763,N_9026);
and U11448 (N_11448,N_9424,N_9136);
nand U11449 (N_11449,N_9694,N_9312);
or U11450 (N_11450,N_9970,N_10359);
and U11451 (N_11451,N_9998,N_10268);
nand U11452 (N_11452,N_9872,N_10298);
nand U11453 (N_11453,N_10481,N_9454);
nand U11454 (N_11454,N_10387,N_9732);
nor U11455 (N_11455,N_10353,N_10107);
nand U11456 (N_11456,N_9073,N_9931);
or U11457 (N_11457,N_9255,N_9010);
xor U11458 (N_11458,N_10240,N_9726);
xnor U11459 (N_11459,N_10243,N_10396);
xor U11460 (N_11460,N_10474,N_9239);
nand U11461 (N_11461,N_9908,N_9019);
xor U11462 (N_11462,N_10142,N_9678);
and U11463 (N_11463,N_10308,N_10249);
nand U11464 (N_11464,N_9873,N_9750);
nor U11465 (N_11465,N_9973,N_9977);
nor U11466 (N_11466,N_9816,N_9975);
and U11467 (N_11467,N_9572,N_10464);
and U11468 (N_11468,N_9904,N_9536);
and U11469 (N_11469,N_10012,N_9399);
and U11470 (N_11470,N_9473,N_9016);
and U11471 (N_11471,N_9483,N_10469);
nand U11472 (N_11472,N_9424,N_9266);
xnor U11473 (N_11473,N_10045,N_9683);
nor U11474 (N_11474,N_9127,N_9979);
or U11475 (N_11475,N_9691,N_10403);
xnor U11476 (N_11476,N_10196,N_9191);
or U11477 (N_11477,N_9952,N_9434);
xor U11478 (N_11478,N_10369,N_9018);
xor U11479 (N_11479,N_9271,N_9574);
nand U11480 (N_11480,N_9709,N_9448);
or U11481 (N_11481,N_10025,N_9148);
xor U11482 (N_11482,N_10005,N_10414);
nor U11483 (N_11483,N_10045,N_9757);
nand U11484 (N_11484,N_9224,N_9217);
nand U11485 (N_11485,N_10395,N_9851);
xor U11486 (N_11486,N_9277,N_10099);
or U11487 (N_11487,N_9832,N_9272);
xnor U11488 (N_11488,N_10352,N_10158);
nand U11489 (N_11489,N_9005,N_10065);
nand U11490 (N_11490,N_9933,N_9518);
xnor U11491 (N_11491,N_9283,N_9602);
or U11492 (N_11492,N_10048,N_9282);
or U11493 (N_11493,N_9534,N_10413);
and U11494 (N_11494,N_9479,N_10155);
or U11495 (N_11495,N_10181,N_9088);
xnor U11496 (N_11496,N_10137,N_10405);
xnor U11497 (N_11497,N_9408,N_9122);
xnor U11498 (N_11498,N_9251,N_9573);
xor U11499 (N_11499,N_9673,N_9094);
nor U11500 (N_11500,N_9020,N_9233);
nor U11501 (N_11501,N_10013,N_9013);
nand U11502 (N_11502,N_9895,N_9974);
and U11503 (N_11503,N_9263,N_10308);
nand U11504 (N_11504,N_9127,N_9112);
nand U11505 (N_11505,N_9067,N_9682);
and U11506 (N_11506,N_9011,N_9543);
xor U11507 (N_11507,N_9453,N_9999);
nand U11508 (N_11508,N_9171,N_10416);
nand U11509 (N_11509,N_9799,N_9096);
nor U11510 (N_11510,N_9468,N_9815);
nor U11511 (N_11511,N_9394,N_9763);
xor U11512 (N_11512,N_9616,N_9467);
or U11513 (N_11513,N_10491,N_10088);
xor U11514 (N_11514,N_9664,N_9382);
or U11515 (N_11515,N_10493,N_9416);
and U11516 (N_11516,N_9383,N_10499);
nor U11517 (N_11517,N_9899,N_9596);
and U11518 (N_11518,N_10450,N_9422);
nor U11519 (N_11519,N_10017,N_9362);
xor U11520 (N_11520,N_10092,N_9372);
nor U11521 (N_11521,N_10436,N_10325);
and U11522 (N_11522,N_10433,N_10149);
or U11523 (N_11523,N_9337,N_10437);
or U11524 (N_11524,N_10220,N_9444);
or U11525 (N_11525,N_9779,N_9758);
and U11526 (N_11526,N_9378,N_9229);
xor U11527 (N_11527,N_9702,N_10336);
nor U11528 (N_11528,N_9187,N_9221);
nor U11529 (N_11529,N_9353,N_9999);
nor U11530 (N_11530,N_9474,N_9172);
xor U11531 (N_11531,N_9678,N_9451);
nand U11532 (N_11532,N_9947,N_9957);
nand U11533 (N_11533,N_9487,N_10042);
and U11534 (N_11534,N_9772,N_9563);
and U11535 (N_11535,N_9034,N_9667);
nand U11536 (N_11536,N_9209,N_9302);
nand U11537 (N_11537,N_9714,N_9630);
xor U11538 (N_11538,N_10125,N_9627);
xnor U11539 (N_11539,N_9089,N_9967);
and U11540 (N_11540,N_9369,N_9147);
nand U11541 (N_11541,N_9367,N_9858);
or U11542 (N_11542,N_9296,N_9731);
and U11543 (N_11543,N_9880,N_10146);
nor U11544 (N_11544,N_9020,N_10023);
and U11545 (N_11545,N_10316,N_9102);
nor U11546 (N_11546,N_10365,N_10165);
and U11547 (N_11547,N_10297,N_10374);
or U11548 (N_11548,N_9189,N_9210);
nand U11549 (N_11549,N_9921,N_9298);
xnor U11550 (N_11550,N_9578,N_10107);
nand U11551 (N_11551,N_9270,N_10264);
or U11552 (N_11552,N_9485,N_10235);
nor U11553 (N_11553,N_9419,N_9182);
xor U11554 (N_11554,N_10401,N_10113);
nand U11555 (N_11555,N_9757,N_9436);
nor U11556 (N_11556,N_9812,N_9808);
or U11557 (N_11557,N_10021,N_9077);
and U11558 (N_11558,N_9600,N_9932);
and U11559 (N_11559,N_10454,N_9052);
nand U11560 (N_11560,N_10064,N_9975);
and U11561 (N_11561,N_9552,N_9081);
nor U11562 (N_11562,N_9888,N_9283);
and U11563 (N_11563,N_9827,N_10032);
nand U11564 (N_11564,N_10223,N_9828);
and U11565 (N_11565,N_9738,N_9056);
nor U11566 (N_11566,N_9835,N_10132);
nor U11567 (N_11567,N_9331,N_9865);
nor U11568 (N_11568,N_10195,N_9209);
or U11569 (N_11569,N_10425,N_9777);
nor U11570 (N_11570,N_9389,N_10290);
xnor U11571 (N_11571,N_9612,N_9332);
and U11572 (N_11572,N_9493,N_9853);
and U11573 (N_11573,N_10404,N_9251);
and U11574 (N_11574,N_9279,N_9155);
xor U11575 (N_11575,N_9270,N_10301);
or U11576 (N_11576,N_9805,N_9505);
nor U11577 (N_11577,N_9814,N_9630);
and U11578 (N_11578,N_9763,N_9102);
or U11579 (N_11579,N_9533,N_9065);
or U11580 (N_11580,N_9416,N_9570);
or U11581 (N_11581,N_9606,N_9790);
nand U11582 (N_11582,N_10229,N_10493);
or U11583 (N_11583,N_10463,N_10070);
nand U11584 (N_11584,N_10391,N_9133);
nand U11585 (N_11585,N_9641,N_10407);
xnor U11586 (N_11586,N_9775,N_10447);
nor U11587 (N_11587,N_9489,N_9595);
and U11588 (N_11588,N_9070,N_9108);
nor U11589 (N_11589,N_9338,N_9238);
xnor U11590 (N_11590,N_10450,N_9250);
nand U11591 (N_11591,N_9017,N_9714);
xor U11592 (N_11592,N_10130,N_10168);
or U11593 (N_11593,N_10248,N_10499);
or U11594 (N_11594,N_10101,N_9842);
or U11595 (N_11595,N_10494,N_9449);
and U11596 (N_11596,N_9932,N_9466);
nand U11597 (N_11597,N_10022,N_10195);
nand U11598 (N_11598,N_10432,N_9940);
xnor U11599 (N_11599,N_10090,N_9469);
or U11600 (N_11600,N_9925,N_9730);
and U11601 (N_11601,N_9461,N_9411);
and U11602 (N_11602,N_10102,N_9274);
nand U11603 (N_11603,N_9030,N_9555);
or U11604 (N_11604,N_9765,N_9288);
xor U11605 (N_11605,N_9428,N_9349);
or U11606 (N_11606,N_9327,N_9681);
nand U11607 (N_11607,N_9784,N_9532);
nor U11608 (N_11608,N_10292,N_9806);
and U11609 (N_11609,N_9444,N_9361);
nand U11610 (N_11610,N_9104,N_9912);
nor U11611 (N_11611,N_9880,N_9039);
or U11612 (N_11612,N_9524,N_9428);
xnor U11613 (N_11613,N_10078,N_9264);
and U11614 (N_11614,N_9668,N_9594);
nor U11615 (N_11615,N_9658,N_9833);
or U11616 (N_11616,N_9120,N_9643);
or U11617 (N_11617,N_10415,N_10065);
nor U11618 (N_11618,N_9214,N_10370);
and U11619 (N_11619,N_9634,N_10257);
xor U11620 (N_11620,N_9639,N_10433);
and U11621 (N_11621,N_9388,N_9892);
and U11622 (N_11622,N_9059,N_9601);
nor U11623 (N_11623,N_9534,N_9772);
and U11624 (N_11624,N_9648,N_9993);
or U11625 (N_11625,N_9556,N_9066);
xnor U11626 (N_11626,N_9631,N_10194);
and U11627 (N_11627,N_9578,N_9949);
nor U11628 (N_11628,N_9807,N_10356);
nor U11629 (N_11629,N_9816,N_9897);
and U11630 (N_11630,N_10098,N_9891);
or U11631 (N_11631,N_9732,N_10380);
xor U11632 (N_11632,N_9263,N_10338);
nand U11633 (N_11633,N_9302,N_9944);
nor U11634 (N_11634,N_9382,N_9157);
nor U11635 (N_11635,N_9448,N_9741);
nand U11636 (N_11636,N_9889,N_9208);
nand U11637 (N_11637,N_9301,N_10081);
nor U11638 (N_11638,N_9678,N_10417);
and U11639 (N_11639,N_10192,N_9027);
and U11640 (N_11640,N_9097,N_9704);
xor U11641 (N_11641,N_9120,N_10278);
nor U11642 (N_11642,N_9142,N_10311);
or U11643 (N_11643,N_10253,N_10415);
or U11644 (N_11644,N_9522,N_9646);
nand U11645 (N_11645,N_9686,N_9000);
nor U11646 (N_11646,N_9154,N_9637);
nand U11647 (N_11647,N_10033,N_10242);
or U11648 (N_11648,N_10260,N_9206);
xnor U11649 (N_11649,N_10045,N_9323);
nor U11650 (N_11650,N_9464,N_9368);
or U11651 (N_11651,N_9284,N_9739);
or U11652 (N_11652,N_9034,N_9613);
and U11653 (N_11653,N_9169,N_9552);
and U11654 (N_11654,N_10088,N_9084);
xnor U11655 (N_11655,N_10135,N_9072);
and U11656 (N_11656,N_9740,N_9198);
and U11657 (N_11657,N_9694,N_9443);
xor U11658 (N_11658,N_9943,N_10481);
and U11659 (N_11659,N_9645,N_9889);
nor U11660 (N_11660,N_10353,N_10278);
xor U11661 (N_11661,N_10166,N_10159);
xor U11662 (N_11662,N_9895,N_9562);
xnor U11663 (N_11663,N_9658,N_9562);
nand U11664 (N_11664,N_9477,N_9644);
xnor U11665 (N_11665,N_9016,N_9837);
nand U11666 (N_11666,N_9112,N_9093);
nand U11667 (N_11667,N_10086,N_9297);
nor U11668 (N_11668,N_10414,N_9966);
xor U11669 (N_11669,N_9489,N_10401);
or U11670 (N_11670,N_9385,N_10039);
xor U11671 (N_11671,N_9955,N_9776);
and U11672 (N_11672,N_9149,N_9874);
nor U11673 (N_11673,N_9382,N_10358);
nand U11674 (N_11674,N_9410,N_9482);
nand U11675 (N_11675,N_9166,N_9036);
and U11676 (N_11676,N_9330,N_9987);
xor U11677 (N_11677,N_10440,N_9851);
nor U11678 (N_11678,N_10057,N_9238);
nor U11679 (N_11679,N_10155,N_10356);
xnor U11680 (N_11680,N_10050,N_10025);
nand U11681 (N_11681,N_10262,N_9406);
nand U11682 (N_11682,N_9105,N_10336);
nor U11683 (N_11683,N_10352,N_10243);
xnor U11684 (N_11684,N_9778,N_9726);
or U11685 (N_11685,N_10396,N_9838);
nor U11686 (N_11686,N_9419,N_9300);
nor U11687 (N_11687,N_9161,N_9995);
or U11688 (N_11688,N_9928,N_9639);
or U11689 (N_11689,N_9132,N_9151);
nor U11690 (N_11690,N_9942,N_9990);
or U11691 (N_11691,N_9738,N_10405);
and U11692 (N_11692,N_10256,N_9524);
and U11693 (N_11693,N_10090,N_9995);
xnor U11694 (N_11694,N_9127,N_9097);
and U11695 (N_11695,N_9584,N_10116);
nor U11696 (N_11696,N_9103,N_9904);
xor U11697 (N_11697,N_9626,N_9249);
nor U11698 (N_11698,N_9119,N_9441);
and U11699 (N_11699,N_9230,N_9459);
xnor U11700 (N_11700,N_9145,N_9702);
xnor U11701 (N_11701,N_10113,N_9309);
xor U11702 (N_11702,N_9033,N_9131);
nor U11703 (N_11703,N_10160,N_10372);
nor U11704 (N_11704,N_9953,N_9450);
or U11705 (N_11705,N_9934,N_9539);
nand U11706 (N_11706,N_10166,N_9347);
nand U11707 (N_11707,N_9117,N_10345);
nand U11708 (N_11708,N_10088,N_9410);
and U11709 (N_11709,N_10091,N_9945);
nand U11710 (N_11710,N_9581,N_10242);
nor U11711 (N_11711,N_9893,N_10100);
nand U11712 (N_11712,N_10344,N_9565);
xnor U11713 (N_11713,N_9044,N_10453);
nor U11714 (N_11714,N_9112,N_9634);
nand U11715 (N_11715,N_9793,N_9796);
xnor U11716 (N_11716,N_9709,N_10078);
xor U11717 (N_11717,N_9290,N_9765);
or U11718 (N_11718,N_9070,N_9134);
xnor U11719 (N_11719,N_10048,N_10054);
nand U11720 (N_11720,N_9334,N_10022);
and U11721 (N_11721,N_10058,N_9301);
or U11722 (N_11722,N_9047,N_9323);
or U11723 (N_11723,N_9076,N_10226);
xor U11724 (N_11724,N_9158,N_10005);
xor U11725 (N_11725,N_10067,N_10311);
nor U11726 (N_11726,N_9627,N_9541);
xnor U11727 (N_11727,N_10422,N_10442);
nor U11728 (N_11728,N_9957,N_9870);
xor U11729 (N_11729,N_9049,N_9280);
and U11730 (N_11730,N_9050,N_10169);
nand U11731 (N_11731,N_10255,N_10314);
nor U11732 (N_11732,N_9695,N_10126);
or U11733 (N_11733,N_9239,N_9217);
xor U11734 (N_11734,N_10161,N_9094);
or U11735 (N_11735,N_9460,N_9366);
xor U11736 (N_11736,N_9789,N_10356);
or U11737 (N_11737,N_9004,N_9973);
nor U11738 (N_11738,N_9903,N_9219);
xor U11739 (N_11739,N_9140,N_9628);
or U11740 (N_11740,N_9831,N_9102);
nand U11741 (N_11741,N_9427,N_9957);
nor U11742 (N_11742,N_9519,N_9724);
or U11743 (N_11743,N_10260,N_9744);
nor U11744 (N_11744,N_10469,N_9644);
nor U11745 (N_11745,N_9037,N_10259);
and U11746 (N_11746,N_10125,N_9402);
xnor U11747 (N_11747,N_9366,N_9517);
nand U11748 (N_11748,N_10203,N_9069);
xor U11749 (N_11749,N_9631,N_10095);
xnor U11750 (N_11750,N_9492,N_9769);
or U11751 (N_11751,N_9823,N_10487);
or U11752 (N_11752,N_10249,N_9850);
xor U11753 (N_11753,N_10048,N_9722);
nand U11754 (N_11754,N_9352,N_9143);
and U11755 (N_11755,N_9362,N_9954);
nor U11756 (N_11756,N_10456,N_10336);
or U11757 (N_11757,N_9165,N_9160);
xor U11758 (N_11758,N_9859,N_9802);
nand U11759 (N_11759,N_9235,N_9894);
xnor U11760 (N_11760,N_10355,N_9850);
nand U11761 (N_11761,N_9469,N_9085);
nand U11762 (N_11762,N_10011,N_10302);
or U11763 (N_11763,N_9941,N_9479);
or U11764 (N_11764,N_9725,N_9891);
and U11765 (N_11765,N_9193,N_9558);
nor U11766 (N_11766,N_9204,N_10138);
nor U11767 (N_11767,N_9949,N_9846);
nand U11768 (N_11768,N_10375,N_9654);
or U11769 (N_11769,N_9335,N_9806);
or U11770 (N_11770,N_9128,N_10312);
nand U11771 (N_11771,N_9525,N_9273);
and U11772 (N_11772,N_9044,N_9726);
nand U11773 (N_11773,N_9969,N_9601);
xor U11774 (N_11774,N_9974,N_9722);
or U11775 (N_11775,N_9179,N_9362);
nor U11776 (N_11776,N_9339,N_10233);
xor U11777 (N_11777,N_9208,N_9872);
xor U11778 (N_11778,N_9453,N_9807);
xor U11779 (N_11779,N_9308,N_9526);
or U11780 (N_11780,N_10358,N_10257);
and U11781 (N_11781,N_10235,N_9441);
or U11782 (N_11782,N_9150,N_10222);
xnor U11783 (N_11783,N_10499,N_10485);
xor U11784 (N_11784,N_10295,N_10090);
and U11785 (N_11785,N_9793,N_10325);
xor U11786 (N_11786,N_9853,N_9288);
and U11787 (N_11787,N_9711,N_9307);
nand U11788 (N_11788,N_10242,N_10176);
or U11789 (N_11789,N_9406,N_9307);
xnor U11790 (N_11790,N_9741,N_9487);
or U11791 (N_11791,N_9749,N_9050);
xnor U11792 (N_11792,N_10046,N_10462);
and U11793 (N_11793,N_9349,N_9385);
nor U11794 (N_11794,N_9629,N_9285);
xnor U11795 (N_11795,N_9877,N_9143);
or U11796 (N_11796,N_9845,N_9285);
nand U11797 (N_11797,N_9363,N_9719);
nand U11798 (N_11798,N_9934,N_10295);
nand U11799 (N_11799,N_9126,N_9622);
nand U11800 (N_11800,N_9865,N_9778);
or U11801 (N_11801,N_10196,N_9426);
or U11802 (N_11802,N_9002,N_10270);
or U11803 (N_11803,N_9014,N_9991);
nor U11804 (N_11804,N_9754,N_9144);
and U11805 (N_11805,N_10222,N_9088);
nor U11806 (N_11806,N_10143,N_10057);
xor U11807 (N_11807,N_9727,N_9910);
nor U11808 (N_11808,N_9950,N_9578);
xor U11809 (N_11809,N_9079,N_9413);
or U11810 (N_11810,N_9592,N_9130);
and U11811 (N_11811,N_9218,N_9906);
and U11812 (N_11812,N_10245,N_9905);
or U11813 (N_11813,N_9607,N_9065);
or U11814 (N_11814,N_10142,N_9629);
xor U11815 (N_11815,N_10426,N_9834);
nor U11816 (N_11816,N_9194,N_10370);
or U11817 (N_11817,N_9800,N_9634);
nor U11818 (N_11818,N_10065,N_9344);
and U11819 (N_11819,N_9709,N_9387);
nand U11820 (N_11820,N_9487,N_9356);
nor U11821 (N_11821,N_9750,N_9058);
or U11822 (N_11822,N_9245,N_10120);
and U11823 (N_11823,N_10473,N_9307);
xnor U11824 (N_11824,N_10423,N_10072);
xnor U11825 (N_11825,N_10499,N_9526);
and U11826 (N_11826,N_9505,N_9421);
nand U11827 (N_11827,N_10305,N_9822);
nor U11828 (N_11828,N_9865,N_10296);
nand U11829 (N_11829,N_10202,N_9592);
or U11830 (N_11830,N_9152,N_9229);
nand U11831 (N_11831,N_9777,N_9850);
and U11832 (N_11832,N_9672,N_10266);
xor U11833 (N_11833,N_10148,N_10479);
or U11834 (N_11834,N_10024,N_10159);
nor U11835 (N_11835,N_9432,N_9231);
xnor U11836 (N_11836,N_10336,N_9917);
nand U11837 (N_11837,N_9157,N_9187);
and U11838 (N_11838,N_10000,N_10244);
nor U11839 (N_11839,N_9036,N_9111);
nor U11840 (N_11840,N_9988,N_9541);
or U11841 (N_11841,N_10296,N_9873);
xnor U11842 (N_11842,N_10067,N_9844);
or U11843 (N_11843,N_9250,N_10252);
or U11844 (N_11844,N_9456,N_9186);
and U11845 (N_11845,N_9967,N_9854);
xor U11846 (N_11846,N_9332,N_10478);
nand U11847 (N_11847,N_9029,N_9400);
and U11848 (N_11848,N_9053,N_9923);
nor U11849 (N_11849,N_9274,N_9142);
and U11850 (N_11850,N_9695,N_9711);
nand U11851 (N_11851,N_9340,N_9384);
xnor U11852 (N_11852,N_9438,N_9730);
nand U11853 (N_11853,N_9416,N_9397);
nand U11854 (N_11854,N_10088,N_9875);
and U11855 (N_11855,N_10449,N_10210);
nor U11856 (N_11856,N_9083,N_9383);
nor U11857 (N_11857,N_9773,N_9726);
nor U11858 (N_11858,N_10151,N_10427);
and U11859 (N_11859,N_9740,N_10433);
nor U11860 (N_11860,N_9281,N_10468);
nand U11861 (N_11861,N_9970,N_10294);
nand U11862 (N_11862,N_9638,N_9093);
xnor U11863 (N_11863,N_9613,N_9295);
or U11864 (N_11864,N_10410,N_9820);
or U11865 (N_11865,N_10232,N_9247);
nor U11866 (N_11866,N_10279,N_9981);
nand U11867 (N_11867,N_9966,N_10050);
nand U11868 (N_11868,N_9785,N_9300);
nor U11869 (N_11869,N_10040,N_9001);
and U11870 (N_11870,N_10426,N_9230);
nor U11871 (N_11871,N_9298,N_9627);
xnor U11872 (N_11872,N_9571,N_9615);
or U11873 (N_11873,N_10367,N_9886);
nand U11874 (N_11874,N_9066,N_9509);
and U11875 (N_11875,N_9948,N_9068);
xnor U11876 (N_11876,N_9252,N_9320);
and U11877 (N_11877,N_10265,N_9035);
nor U11878 (N_11878,N_9525,N_9852);
nor U11879 (N_11879,N_9842,N_10145);
or U11880 (N_11880,N_9644,N_9578);
xor U11881 (N_11881,N_9346,N_9388);
nand U11882 (N_11882,N_10055,N_10261);
and U11883 (N_11883,N_10084,N_10442);
and U11884 (N_11884,N_10016,N_9409);
nor U11885 (N_11885,N_10088,N_9821);
nand U11886 (N_11886,N_10058,N_9764);
xnor U11887 (N_11887,N_9901,N_9848);
or U11888 (N_11888,N_9135,N_9946);
and U11889 (N_11889,N_9210,N_9595);
and U11890 (N_11890,N_9890,N_10147);
nand U11891 (N_11891,N_10036,N_10237);
nor U11892 (N_11892,N_9172,N_9096);
and U11893 (N_11893,N_9358,N_9177);
nand U11894 (N_11894,N_9874,N_9542);
xor U11895 (N_11895,N_9678,N_10085);
and U11896 (N_11896,N_9646,N_9903);
nand U11897 (N_11897,N_9414,N_9715);
and U11898 (N_11898,N_9777,N_9395);
or U11899 (N_11899,N_10458,N_9571);
nand U11900 (N_11900,N_9255,N_10099);
nor U11901 (N_11901,N_9182,N_9672);
and U11902 (N_11902,N_9366,N_9949);
xnor U11903 (N_11903,N_10411,N_9221);
nor U11904 (N_11904,N_10189,N_9596);
xor U11905 (N_11905,N_9644,N_9949);
nor U11906 (N_11906,N_9486,N_9423);
nor U11907 (N_11907,N_9260,N_10417);
or U11908 (N_11908,N_9923,N_9222);
xor U11909 (N_11909,N_10357,N_9475);
and U11910 (N_11910,N_9595,N_9258);
nand U11911 (N_11911,N_10232,N_9577);
xnor U11912 (N_11912,N_10138,N_9208);
nor U11913 (N_11913,N_9302,N_10017);
nand U11914 (N_11914,N_9782,N_10478);
or U11915 (N_11915,N_10150,N_9041);
xor U11916 (N_11916,N_10474,N_9617);
xor U11917 (N_11917,N_10420,N_9728);
xor U11918 (N_11918,N_9030,N_9230);
nand U11919 (N_11919,N_9094,N_9713);
xnor U11920 (N_11920,N_9193,N_10308);
nor U11921 (N_11921,N_10441,N_9897);
nand U11922 (N_11922,N_9512,N_10204);
or U11923 (N_11923,N_9264,N_10245);
xnor U11924 (N_11924,N_9175,N_10171);
nor U11925 (N_11925,N_9563,N_10424);
nor U11926 (N_11926,N_10103,N_9562);
and U11927 (N_11927,N_9812,N_9468);
xor U11928 (N_11928,N_9090,N_10345);
and U11929 (N_11929,N_9192,N_9952);
and U11930 (N_11930,N_9993,N_9927);
and U11931 (N_11931,N_9393,N_10202);
and U11932 (N_11932,N_10226,N_9555);
or U11933 (N_11933,N_9873,N_9624);
xor U11934 (N_11934,N_10451,N_10293);
and U11935 (N_11935,N_10040,N_9448);
or U11936 (N_11936,N_9488,N_10309);
or U11937 (N_11937,N_9050,N_9580);
xnor U11938 (N_11938,N_9053,N_10206);
and U11939 (N_11939,N_9264,N_9779);
and U11940 (N_11940,N_9425,N_9574);
nor U11941 (N_11941,N_10463,N_9770);
or U11942 (N_11942,N_9444,N_9170);
xor U11943 (N_11943,N_10165,N_9091);
nor U11944 (N_11944,N_9595,N_9584);
nand U11945 (N_11945,N_10362,N_10200);
nand U11946 (N_11946,N_9641,N_10465);
xor U11947 (N_11947,N_9813,N_10426);
or U11948 (N_11948,N_9568,N_10348);
nor U11949 (N_11949,N_9918,N_9482);
nand U11950 (N_11950,N_10131,N_10312);
xnor U11951 (N_11951,N_10360,N_10351);
and U11952 (N_11952,N_10085,N_9862);
nor U11953 (N_11953,N_9929,N_9181);
or U11954 (N_11954,N_9756,N_9512);
and U11955 (N_11955,N_9700,N_9224);
or U11956 (N_11956,N_9918,N_9885);
nor U11957 (N_11957,N_9798,N_9231);
xnor U11958 (N_11958,N_10025,N_9195);
nand U11959 (N_11959,N_9117,N_10301);
or U11960 (N_11960,N_9143,N_10165);
nand U11961 (N_11961,N_10281,N_10255);
nor U11962 (N_11962,N_10111,N_10036);
and U11963 (N_11963,N_10104,N_10423);
xnor U11964 (N_11964,N_9309,N_9977);
nor U11965 (N_11965,N_9310,N_10415);
xor U11966 (N_11966,N_9955,N_9787);
and U11967 (N_11967,N_9746,N_9534);
nor U11968 (N_11968,N_9771,N_9836);
nand U11969 (N_11969,N_9127,N_9778);
nand U11970 (N_11970,N_9323,N_9487);
nor U11971 (N_11971,N_9984,N_9358);
nor U11972 (N_11972,N_10097,N_10141);
or U11973 (N_11973,N_10002,N_10342);
xnor U11974 (N_11974,N_9005,N_10325);
or U11975 (N_11975,N_9322,N_10272);
xnor U11976 (N_11976,N_9824,N_9316);
nor U11977 (N_11977,N_10059,N_10174);
and U11978 (N_11978,N_10407,N_10386);
xor U11979 (N_11979,N_9819,N_9901);
xor U11980 (N_11980,N_10105,N_9711);
nor U11981 (N_11981,N_9754,N_9038);
nand U11982 (N_11982,N_9570,N_9167);
xor U11983 (N_11983,N_10494,N_10437);
xnor U11984 (N_11984,N_9756,N_9433);
nor U11985 (N_11985,N_9188,N_9550);
nor U11986 (N_11986,N_10229,N_10132);
or U11987 (N_11987,N_10002,N_10339);
nand U11988 (N_11988,N_9165,N_9368);
nand U11989 (N_11989,N_9391,N_9806);
or U11990 (N_11990,N_10211,N_9049);
xor U11991 (N_11991,N_9756,N_9590);
xor U11992 (N_11992,N_9043,N_9235);
and U11993 (N_11993,N_10145,N_9757);
nand U11994 (N_11994,N_10077,N_9783);
nand U11995 (N_11995,N_9412,N_10132);
nand U11996 (N_11996,N_10004,N_10062);
nand U11997 (N_11997,N_10008,N_9175);
nand U11998 (N_11998,N_9169,N_10451);
xnor U11999 (N_11999,N_9125,N_9854);
or U12000 (N_12000,N_11706,N_11265);
nand U12001 (N_12001,N_11449,N_10598);
or U12002 (N_12002,N_11747,N_11285);
nand U12003 (N_12003,N_11567,N_11239);
and U12004 (N_12004,N_11486,N_10567);
or U12005 (N_12005,N_11614,N_11073);
and U12006 (N_12006,N_10924,N_11993);
nor U12007 (N_12007,N_11731,N_11446);
and U12008 (N_12008,N_11734,N_11912);
or U12009 (N_12009,N_11241,N_10688);
xnor U12010 (N_12010,N_10736,N_11115);
and U12011 (N_12011,N_10712,N_10915);
and U12012 (N_12012,N_11774,N_11742);
xnor U12013 (N_12013,N_11832,N_10600);
nand U12014 (N_12014,N_11368,N_11652);
xnor U12015 (N_12015,N_11735,N_11992);
nand U12016 (N_12016,N_11246,N_10585);
nor U12017 (N_12017,N_11506,N_10895);
and U12018 (N_12018,N_10738,N_11006);
and U12019 (N_12019,N_11269,N_10641);
and U12020 (N_12020,N_10979,N_10954);
nand U12021 (N_12021,N_10861,N_11540);
xnor U12022 (N_12022,N_11337,N_11383);
nand U12023 (N_12023,N_11234,N_11692);
xor U12024 (N_12024,N_10591,N_11112);
nor U12025 (N_12025,N_11494,N_11635);
xor U12026 (N_12026,N_10938,N_11661);
xnor U12027 (N_12027,N_10507,N_11932);
nand U12028 (N_12028,N_11447,N_10742);
nand U12029 (N_12029,N_11012,N_11913);
xnor U12030 (N_12030,N_10822,N_10682);
nor U12031 (N_12031,N_11210,N_11878);
and U12032 (N_12032,N_11238,N_10616);
nand U12033 (N_12033,N_10811,N_11429);
nand U12034 (N_12034,N_10680,N_11862);
xnor U12035 (N_12035,N_11184,N_10662);
xnor U12036 (N_12036,N_11709,N_11031);
nand U12037 (N_12037,N_10885,N_11746);
nand U12038 (N_12038,N_10597,N_11434);
nor U12039 (N_12039,N_11532,N_11122);
xor U12040 (N_12040,N_10946,N_11025);
nor U12041 (N_12041,N_11630,N_11398);
nand U12042 (N_12042,N_10886,N_10615);
or U12043 (N_12043,N_11631,N_10750);
and U12044 (N_12044,N_10685,N_11615);
and U12045 (N_12045,N_11471,N_11312);
and U12046 (N_12046,N_10543,N_10710);
and U12047 (N_12047,N_11625,N_11147);
xor U12048 (N_12048,N_10996,N_11588);
nor U12049 (N_12049,N_11552,N_11215);
xnor U12050 (N_12050,N_10699,N_11657);
or U12051 (N_12051,N_10661,N_11839);
nand U12052 (N_12052,N_11099,N_11185);
and U12053 (N_12053,N_11335,N_11771);
nor U12054 (N_12054,N_10723,N_10834);
xor U12055 (N_12055,N_10559,N_10576);
nor U12056 (N_12056,N_11008,N_11310);
nand U12057 (N_12057,N_10744,N_11138);
nor U12058 (N_12058,N_11518,N_11050);
or U12059 (N_12059,N_11790,N_10858);
xnor U12060 (N_12060,N_10583,N_11564);
and U12061 (N_12061,N_11780,N_11290);
nor U12062 (N_12062,N_11703,N_11413);
xnor U12063 (N_12063,N_10827,N_11578);
and U12064 (N_12064,N_11690,N_11497);
or U12065 (N_12065,N_10883,N_11281);
nand U12066 (N_12066,N_11872,N_11928);
or U12067 (N_12067,N_11792,N_11204);
and U12068 (N_12068,N_11075,N_11755);
and U12069 (N_12069,N_11880,N_10521);
and U12070 (N_12070,N_11427,N_10893);
nor U12071 (N_12071,N_11618,N_11745);
nor U12072 (N_12072,N_10823,N_11390);
nand U12073 (N_12073,N_10629,N_11814);
xnor U12074 (N_12074,N_10556,N_11410);
xnor U12075 (N_12075,N_11543,N_10577);
and U12076 (N_12076,N_11266,N_11760);
xnor U12077 (N_12077,N_11612,N_10604);
or U12078 (N_12078,N_10876,N_10651);
xnor U12079 (N_12079,N_11693,N_11385);
and U12080 (N_12080,N_10809,N_11902);
xor U12081 (N_12081,N_11177,N_11178);
nand U12082 (N_12082,N_11049,N_11289);
or U12083 (N_12083,N_11923,N_11977);
xor U12084 (N_12084,N_11864,N_11000);
xor U12085 (N_12085,N_10913,N_11757);
and U12086 (N_12086,N_10960,N_10584);
nand U12087 (N_12087,N_11549,N_11988);
nand U12088 (N_12088,N_10792,N_11871);
nor U12089 (N_12089,N_10855,N_10638);
xnor U12090 (N_12090,N_11304,N_11996);
nor U12091 (N_12091,N_10956,N_11991);
xor U12092 (N_12092,N_11605,N_10833);
or U12093 (N_12093,N_11736,N_11081);
or U12094 (N_12094,N_11901,N_11906);
xor U12095 (N_12095,N_11953,N_11607);
xnor U12096 (N_12096,N_11647,N_10509);
xnor U12097 (N_12097,N_10803,N_10944);
xor U12098 (N_12098,N_11576,N_11551);
nor U12099 (N_12099,N_11949,N_11950);
and U12100 (N_12100,N_10967,N_11525);
nand U12101 (N_12101,N_11719,N_11749);
xnor U12102 (N_12102,N_10733,N_11341);
or U12103 (N_12103,N_10801,N_11989);
xnor U12104 (N_12104,N_11331,N_10660);
and U12105 (N_12105,N_11009,N_10757);
nand U12106 (N_12106,N_11909,N_11581);
xor U12107 (N_12107,N_11198,N_11788);
xnor U12108 (N_12108,N_10903,N_11557);
nor U12109 (N_12109,N_11333,N_11085);
and U12110 (N_12110,N_11628,N_11051);
nand U12111 (N_12111,N_11848,N_10961);
xor U12112 (N_12112,N_11058,N_10725);
nand U12113 (N_12113,N_11979,N_11695);
nor U12114 (N_12114,N_10706,N_10802);
or U12115 (N_12115,N_10872,N_11641);
nand U12116 (N_12116,N_10874,N_11765);
nor U12117 (N_12117,N_10531,N_10845);
nor U12118 (N_12118,N_11712,N_11392);
nor U12119 (N_12119,N_11538,N_11599);
and U12120 (N_12120,N_11272,N_11109);
nor U12121 (N_12121,N_11029,N_10752);
xnor U12122 (N_12122,N_11119,N_10994);
or U12123 (N_12123,N_11512,N_11523);
and U12124 (N_12124,N_11343,N_11741);
or U12125 (N_12125,N_11639,N_11918);
and U12126 (N_12126,N_11257,N_10523);
and U12127 (N_12127,N_10628,N_10675);
and U12128 (N_12128,N_10578,N_11980);
nand U12129 (N_12129,N_11035,N_11033);
nor U12130 (N_12130,N_11587,N_10730);
nand U12131 (N_12131,N_11271,N_10739);
xnor U12132 (N_12132,N_11597,N_11422);
and U12133 (N_12133,N_11252,N_11221);
nor U12134 (N_12134,N_11188,N_11968);
and U12135 (N_12135,N_11855,N_11573);
nand U12136 (N_12136,N_10678,N_11300);
nor U12137 (N_12137,N_11710,N_11898);
and U12138 (N_12138,N_11211,N_11786);
nor U12139 (N_12139,N_10784,N_11516);
and U12140 (N_12140,N_10995,N_10653);
xnor U12141 (N_12141,N_11847,N_11756);
nor U12142 (N_12142,N_11773,N_10973);
nor U12143 (N_12143,N_10511,N_10982);
nor U12144 (N_12144,N_11379,N_10761);
nand U12145 (N_12145,N_11854,N_11268);
nor U12146 (N_12146,N_11232,N_11260);
nand U12147 (N_12147,N_11811,N_11259);
xor U12148 (N_12148,N_11451,N_11620);
nand U12149 (N_12149,N_11859,N_10663);
nor U12150 (N_12150,N_10846,N_10852);
nand U12151 (N_12151,N_11280,N_11226);
nand U12152 (N_12152,N_11632,N_11127);
or U12153 (N_12153,N_11342,N_11868);
and U12154 (N_12154,N_10613,N_10520);
nor U12155 (N_12155,N_11126,N_11024);
xor U12156 (N_12156,N_10970,N_11296);
nor U12157 (N_12157,N_10546,N_11469);
nor U12158 (N_12158,N_10514,N_11155);
nand U12159 (N_12159,N_11242,N_10878);
nand U12160 (N_12160,N_11524,N_10525);
nand U12161 (N_12161,N_11262,N_10528);
or U12162 (N_12162,N_10650,N_11815);
nor U12163 (N_12163,N_11776,N_11003);
xor U12164 (N_12164,N_11930,N_11542);
or U12165 (N_12165,N_11857,N_10606);
or U12166 (N_12166,N_10636,N_10605);
nand U12167 (N_12167,N_11403,N_11806);
xnor U12168 (N_12168,N_11227,N_11802);
and U12169 (N_12169,N_10542,N_11481);
xnor U12170 (N_12170,N_11955,N_10909);
xnor U12171 (N_12171,N_11927,N_11345);
xnor U12172 (N_12172,N_11584,N_11400);
nand U12173 (N_12173,N_11782,N_11145);
xor U12174 (N_12174,N_11648,N_11546);
nor U12175 (N_12175,N_10880,N_10934);
nand U12176 (N_12176,N_11526,N_10700);
xnor U12177 (N_12177,N_11603,N_11062);
or U12178 (N_12178,N_11640,N_11201);
and U12179 (N_12179,N_11521,N_11350);
and U12180 (N_12180,N_11078,N_10748);
nor U12181 (N_12181,N_10781,N_10544);
and U12182 (N_12182,N_11946,N_10697);
xor U12183 (N_12183,N_10670,N_11353);
and U12184 (N_12184,N_11154,N_11541);
or U12185 (N_12185,N_11087,N_10592);
nand U12186 (N_12186,N_10873,N_11495);
nor U12187 (N_12187,N_10571,N_10950);
and U12188 (N_12188,N_10690,N_11807);
nor U12189 (N_12189,N_11298,N_10770);
xnor U12190 (N_12190,N_11669,N_11517);
nand U12191 (N_12191,N_11671,N_10758);
xor U12192 (N_12192,N_11863,N_10947);
or U12193 (N_12193,N_10842,N_10987);
nor U12194 (N_12194,N_11384,N_10639);
and U12195 (N_12195,N_10993,N_11600);
and U12196 (N_12196,N_10821,N_11254);
and U12197 (N_12197,N_11483,N_11327);
and U12198 (N_12198,N_11818,N_11834);
nand U12199 (N_12199,N_10743,N_11228);
nand U12200 (N_12200,N_11100,N_10790);
nand U12201 (N_12201,N_11504,N_11954);
nand U12202 (N_12202,N_11365,N_10922);
nor U12203 (N_12203,N_10704,N_10702);
xnor U12204 (N_12204,N_11501,N_11047);
and U12205 (N_12205,N_11091,N_10930);
xor U12206 (N_12206,N_11108,N_11409);
and U12207 (N_12207,N_10839,N_11467);
xor U12208 (N_12208,N_11424,N_11173);
nand U12209 (N_12209,N_10687,N_11443);
nand U12210 (N_12210,N_10870,N_10911);
or U12211 (N_12211,N_11642,N_10515);
nor U12212 (N_12212,N_11161,N_11206);
or U12213 (N_12213,N_11374,N_11137);
nor U12214 (N_12214,N_11141,N_11924);
nand U12215 (N_12215,N_10527,N_10575);
xor U12216 (N_12216,N_11027,N_10889);
xor U12217 (N_12217,N_10554,N_11513);
nor U12218 (N_12218,N_11558,N_11478);
xor U12219 (N_12219,N_11083,N_11613);
nand U12220 (N_12220,N_11480,N_11767);
nor U12221 (N_12221,N_11611,N_11225);
nor U12222 (N_12222,N_11382,N_11836);
nand U12223 (N_12223,N_11900,N_11948);
or U12224 (N_12224,N_11363,N_10588);
nor U12225 (N_12225,N_11438,N_11925);
or U12226 (N_12226,N_11275,N_10611);
or U12227 (N_12227,N_11415,N_10727);
nand U12228 (N_12228,N_11196,N_11684);
nand U12229 (N_12229,N_10871,N_10853);
or U12230 (N_12230,N_10539,N_11701);
nor U12231 (N_12231,N_10709,N_11897);
nand U12232 (N_12232,N_11231,N_11441);
nor U12233 (N_12233,N_10829,N_11287);
or U12234 (N_12234,N_11510,N_10789);
nand U12235 (N_12235,N_11922,N_11514);
xnor U12236 (N_12236,N_11825,N_11740);
nor U12237 (N_12237,N_11136,N_10879);
nor U12238 (N_12238,N_10620,N_11633);
or U12239 (N_12239,N_11837,N_11941);
nand U12240 (N_12240,N_11355,N_10732);
nor U12241 (N_12241,N_10847,N_11426);
xnor U12242 (N_12242,N_11937,N_11842);
nor U12243 (N_12243,N_10892,N_11969);
xor U12244 (N_12244,N_11961,N_10512);
nor U12245 (N_12245,N_11899,N_11216);
xor U12246 (N_12246,N_11399,N_11308);
nand U12247 (N_12247,N_11299,N_11655);
and U12248 (N_12248,N_11841,N_10537);
xnor U12249 (N_12249,N_10652,N_11131);
nor U12250 (N_12250,N_11015,N_11676);
nor U12251 (N_12251,N_11255,N_11369);
nor U12252 (N_12252,N_10898,N_10551);
nand U12253 (N_12253,N_11174,N_10608);
nand U12254 (N_12254,N_10983,N_11354);
or U12255 (N_12255,N_10658,N_11130);
or U12256 (N_12256,N_10817,N_11711);
or U12257 (N_12257,N_11240,N_11649);
nand U12258 (N_12258,N_10881,N_11063);
and U12259 (N_12259,N_10557,N_11235);
and U12260 (N_12260,N_11678,N_11534);
or U12261 (N_12261,N_11812,N_11737);
and U12262 (N_12262,N_11450,N_11966);
nand U12263 (N_12263,N_11219,N_11046);
and U12264 (N_12264,N_11598,N_11001);
and U12265 (N_12265,N_10560,N_11143);
nand U12266 (N_12266,N_11865,N_11785);
or U12267 (N_12267,N_11978,N_11391);
nand U12268 (N_12268,N_10558,N_10500);
and U12269 (N_12269,N_11082,N_11650);
nor U12270 (N_12270,N_11997,N_11402);
or U12271 (N_12271,N_10582,N_11042);
nor U12272 (N_12272,N_11116,N_10785);
and U12273 (N_12273,N_10989,N_10717);
nor U12274 (N_12274,N_11853,N_11183);
or U12275 (N_12275,N_11778,N_10957);
or U12276 (N_12276,N_11401,N_10856);
or U12277 (N_12277,N_10698,N_11846);
xnor U12278 (N_12278,N_10695,N_11707);
or U12279 (N_12279,N_10741,N_11781);
and U12280 (N_12280,N_11258,N_10780);
or U12281 (N_12281,N_11187,N_11653);
or U12282 (N_12282,N_11039,N_11585);
xnor U12283 (N_12283,N_11437,N_11609);
xnor U12284 (N_12284,N_11835,N_11140);
and U12285 (N_12285,N_11456,N_11366);
and U12286 (N_12286,N_10634,N_10580);
or U12287 (N_12287,N_11784,N_11995);
nand U12288 (N_12288,N_11586,N_11889);
or U12289 (N_12289,N_11887,N_10666);
or U12290 (N_12290,N_11626,N_11861);
xnor U12291 (N_12291,N_10971,N_10664);
nor U12292 (N_12292,N_10796,N_10617);
nand U12293 (N_12293,N_11654,N_11247);
xnor U12294 (N_12294,N_11824,N_11651);
nor U12295 (N_12295,N_10986,N_11111);
xor U12296 (N_12296,N_11459,N_11153);
nor U12297 (N_12297,N_10831,N_11761);
xor U12298 (N_12298,N_11321,N_11945);
or U12299 (N_12299,N_11687,N_10923);
nand U12300 (N_12300,N_10693,N_10503);
nor U12301 (N_12301,N_10948,N_11556);
xnor U12302 (N_12302,N_10774,N_10549);
xor U12303 (N_12303,N_11002,N_11301);
or U12304 (N_12304,N_11851,N_11207);
xnor U12305 (N_12305,N_11214,N_11903);
and U12306 (N_12306,N_10935,N_11984);
nand U12307 (N_12307,N_10762,N_10804);
nand U12308 (N_12308,N_11224,N_11146);
nor U12309 (N_12309,N_11487,N_11306);
or U12310 (N_12310,N_10825,N_11502);
and U12311 (N_12311,N_11565,N_10731);
or U12312 (N_12312,N_11055,N_11753);
nor U12313 (N_12313,N_11118,N_11931);
or U12314 (N_12314,N_10978,N_11570);
nand U12315 (N_12315,N_10764,N_11005);
xor U12316 (N_12316,N_10838,N_11559);
nand U12317 (N_12317,N_10850,N_10621);
nor U12318 (N_12318,N_11358,N_11579);
xor U12319 (N_12319,N_11905,N_11831);
or U12320 (N_12320,N_10716,N_11357);
xor U12321 (N_12321,N_11370,N_11139);
xnor U12322 (N_12322,N_11274,N_11129);
nand U12323 (N_12323,N_11939,N_11417);
nand U12324 (N_12324,N_11103,N_10976);
or U12325 (N_12325,N_10635,N_11772);
or U12326 (N_12326,N_11970,N_11577);
xor U12327 (N_12327,N_11376,N_11372);
or U12328 (N_12328,N_11346,N_10925);
and U12329 (N_12329,N_11168,N_11076);
xor U12330 (N_12330,N_11074,N_11465);
or U12331 (N_12331,N_10800,N_11072);
or U12332 (N_12332,N_11016,N_10953);
nand U12333 (N_12333,N_11974,N_11233);
or U12334 (N_12334,N_10767,N_10656);
nor U12335 (N_12335,N_11535,N_10713);
xor U12336 (N_12336,N_10619,N_11022);
xor U12337 (N_12337,N_10965,N_11533);
and U12338 (N_12338,N_11389,N_11037);
xnor U12339 (N_12339,N_10633,N_10808);
nor U12340 (N_12340,N_10771,N_11220);
nand U12341 (N_12341,N_10673,N_11762);
nor U12342 (N_12342,N_10566,N_11263);
nor U12343 (N_12343,N_10955,N_11998);
or U12344 (N_12344,N_11328,N_11721);
nand U12345 (N_12345,N_11591,N_10734);
xnor U12346 (N_12346,N_10769,N_11412);
nor U12347 (N_12347,N_10642,N_10927);
nor U12348 (N_12348,N_10863,N_10990);
or U12349 (N_12349,N_11810,N_11248);
or U12350 (N_12350,N_10644,N_10533);
xnor U12351 (N_12351,N_10541,N_11169);
nand U12352 (N_12352,N_10759,N_11805);
and U12353 (N_12353,N_11895,N_11869);
or U12354 (N_12354,N_10504,N_11470);
nand U12355 (N_12355,N_11666,N_10648);
nand U12356 (N_12356,N_10686,N_11550);
nor U12357 (N_12357,N_11890,N_10910);
nor U12358 (N_12358,N_11102,N_10798);
xnor U12359 (N_12359,N_11416,N_11826);
nand U12360 (N_12360,N_10937,N_10772);
nand U12361 (N_12361,N_10791,N_11303);
nor U12362 (N_12362,N_10696,N_11194);
and U12363 (N_12363,N_10522,N_11688);
xnor U12364 (N_12364,N_11957,N_10779);
nand U12365 (N_12365,N_11791,N_11420);
or U12366 (N_12366,N_11052,N_10508);
or U12367 (N_12367,N_11999,N_10787);
and U12368 (N_12368,N_11423,N_10891);
nand U12369 (N_12369,N_10875,N_11668);
xnor U12370 (N_12370,N_11849,N_11894);
nor U12371 (N_12371,N_11729,N_11987);
nor U12372 (N_12372,N_11044,N_11014);
nor U12373 (N_12373,N_11041,N_11457);
and U12374 (N_12374,N_10538,N_10835);
or U12375 (N_12375,N_10722,N_11681);
and U12376 (N_12376,N_11689,N_11458);
or U12377 (N_12377,N_11844,N_10988);
xor U12378 (N_12378,N_11870,N_10939);
nand U12379 (N_12379,N_11404,N_11876);
and U12380 (N_12380,N_10540,N_11562);
and U12381 (N_12381,N_11574,N_10864);
nor U12382 (N_12382,N_11503,N_11720);
xor U12383 (N_12383,N_11770,N_10669);
and U12384 (N_12384,N_10799,N_11627);
nand U12385 (N_12385,N_11691,N_11004);
xor U12386 (N_12386,N_11309,N_11679);
xor U12387 (N_12387,N_11482,N_10899);
nor U12388 (N_12388,N_11943,N_11388);
xor U12389 (N_12389,N_11172,N_11123);
and U12390 (N_12390,N_11209,N_10806);
nand U12391 (N_12391,N_11594,N_11873);
nor U12392 (N_12392,N_11572,N_11125);
xnor U12393 (N_12393,N_11332,N_11951);
or U12394 (N_12394,N_10506,N_10708);
xor U12395 (N_12395,N_11536,N_10768);
nor U12396 (N_12396,N_11833,N_11933);
or U12397 (N_12397,N_11601,N_11011);
and U12398 (N_12398,N_11674,N_11317);
xnor U12399 (N_12399,N_11697,N_11580);
nand U12400 (N_12400,N_10820,N_11251);
or U12401 (N_12401,N_11699,N_11499);
or U12402 (N_12402,N_11132,N_11726);
nor U12403 (N_12403,N_11708,N_11982);
nor U12404 (N_12404,N_10602,N_11843);
or U12405 (N_12405,N_10705,N_10726);
nand U12406 (N_12406,N_11973,N_10920);
xor U12407 (N_12407,N_11208,N_10857);
nor U12408 (N_12408,N_11783,N_10623);
nand U12409 (N_12409,N_10677,N_10918);
or U12410 (N_12410,N_10794,N_10607);
or U12411 (N_12411,N_10921,N_11881);
xor U12412 (N_12412,N_10884,N_10581);
and U12413 (N_12413,N_10958,N_11714);
or U12414 (N_12414,N_10562,N_11329);
nor U12415 (N_12415,N_11728,N_10715);
nor U12416 (N_12416,N_11067,N_11944);
nor U12417 (N_12417,N_11798,N_11057);
and U12418 (N_12418,N_11971,N_11682);
nor U12419 (N_12419,N_10659,N_11098);
and U12420 (N_12420,N_11644,N_11466);
xor U12421 (N_12421,N_11463,N_11356);
xnor U12422 (N_12422,N_11882,N_11079);
xor U12423 (N_12423,N_11432,N_11670);
nor U12424 (N_12424,N_11621,N_10904);
and U12425 (N_12425,N_11326,N_11938);
and U12426 (N_12426,N_10691,N_11789);
nand U12427 (N_12427,N_11318,N_11320);
and U12428 (N_12428,N_10718,N_11694);
or U12429 (N_12429,N_11981,N_11484);
xnor U12430 (N_12430,N_11637,N_11917);
xnor U12431 (N_12431,N_10951,N_10745);
and U12432 (N_12432,N_11967,N_11730);
or U12433 (N_12433,N_10991,N_11157);
or U12434 (N_12434,N_10962,N_11645);
nor U12435 (N_12435,N_11270,N_10964);
and U12436 (N_12436,N_10902,N_11519);
nand U12437 (N_12437,N_10724,N_10977);
xnor U12438 (N_12438,N_11330,N_10843);
and U12439 (N_12439,N_11860,N_11439);
or U12440 (N_12440,N_11566,N_11821);
nand U12441 (N_12441,N_11407,N_11380);
nor U12442 (N_12442,N_10997,N_11489);
xnor U12443 (N_12443,N_10689,N_10755);
nand U12444 (N_12444,N_10740,N_10665);
and U12445 (N_12445,N_11793,N_10912);
and U12446 (N_12446,N_10753,N_11646);
nor U12447 (N_12447,N_10942,N_10729);
xnor U12448 (N_12448,N_11243,N_10778);
nor U12449 (N_12449,N_11779,N_11539);
nand U12450 (N_12450,N_11959,N_11673);
nand U12451 (N_12451,N_10711,N_10654);
or U12452 (N_12452,N_10795,N_11505);
nor U12453 (N_12453,N_11582,N_10535);
xnor U12454 (N_12454,N_11277,N_11528);
and U12455 (N_12455,N_11947,N_11752);
nand U12456 (N_12456,N_10919,N_11222);
or U12457 (N_12457,N_11093,N_11910);
nor U12458 (N_12458,N_11186,N_10945);
nand U12459 (N_12459,N_10933,N_10932);
nor U12460 (N_12460,N_11908,N_11479);
and U12461 (N_12461,N_11795,N_11364);
nand U12462 (N_12462,N_11769,N_11934);
and U12463 (N_12463,N_11144,N_11829);
nor U12464 (N_12464,N_10818,N_11715);
xnor U12465 (N_12465,N_11373,N_11452);
xor U12466 (N_12466,N_10815,N_11511);
xnor U12467 (N_12467,N_10568,N_10980);
nor U12468 (N_12468,N_11395,N_11856);
or U12469 (N_12469,N_11267,N_10972);
or U12470 (N_12470,N_11718,N_11474);
and U12471 (N_12471,N_10837,N_10579);
and U12472 (N_12472,N_11593,N_11347);
nand U12473 (N_12473,N_10649,N_11583);
nand U12474 (N_12474,N_11629,N_11095);
xnor U12475 (N_12475,N_11292,N_11460);
nor U12476 (N_12476,N_10630,N_11230);
nand U12477 (N_12477,N_10936,N_11663);
nor U12478 (N_12478,N_11751,N_11283);
nand U12479 (N_12479,N_11801,N_10545);
nand U12480 (N_12480,N_11827,N_10844);
or U12481 (N_12481,N_11743,N_11020);
or U12482 (N_12482,N_11884,N_11563);
xnor U12483 (N_12483,N_11101,N_11375);
and U12484 (N_12484,N_10805,N_11929);
and U12485 (N_12485,N_11171,N_11685);
nor U12486 (N_12486,N_10631,N_11069);
nand U12487 (N_12487,N_11371,N_11492);
nand U12488 (N_12488,N_11602,N_11104);
and U12489 (N_12489,N_10728,N_10657);
xnor U12490 (N_12490,N_10679,N_10694);
nor U12491 (N_12491,N_11148,N_11433);
xor U12492 (N_12492,N_11253,N_10550);
and U12493 (N_12493,N_11808,N_11819);
or U12494 (N_12494,N_11162,N_11038);
xnor U12495 (N_12495,N_11976,N_11092);
xor U12496 (N_12496,N_11664,N_11121);
nor U12497 (N_12497,N_10572,N_11084);
nand U12498 (N_12498,N_11282,N_11921);
or U12499 (N_12499,N_11595,N_10783);
or U12500 (N_12500,N_11396,N_10941);
xor U12501 (N_12501,N_11295,N_11656);
xor U12502 (N_12502,N_11799,N_10684);
nand U12503 (N_12503,N_11455,N_11936);
nand U12504 (N_12504,N_11545,N_11472);
or U12505 (N_12505,N_11017,N_10756);
nor U12506 (N_12506,N_11096,N_10836);
and U12507 (N_12507,N_11182,N_11094);
xnor U12508 (N_12508,N_11175,N_11893);
xnor U12509 (N_12509,N_10564,N_11569);
nor U12510 (N_12510,N_10599,N_11705);
xor U12511 (N_12511,N_11361,N_10985);
nor U12512 (N_12512,N_11750,N_10793);
xor U12513 (N_12513,N_11181,N_10992);
and U12514 (N_12514,N_10981,N_11286);
nand U12515 (N_12515,N_10614,N_11940);
xnor U12516 (N_12516,N_11325,N_11405);
nand U12517 (N_12517,N_11097,N_10529);
nand U12518 (N_12518,N_11278,N_10943);
nor U12519 (N_12519,N_11962,N_11419);
xnor U12520 (N_12520,N_11874,N_11675);
or U12521 (N_12521,N_11804,N_11313);
nor U12522 (N_12522,N_11488,N_10974);
xnor U12523 (N_12523,N_10646,N_11195);
nor U12524 (N_12524,N_11911,N_11021);
and U12525 (N_12525,N_10609,N_10782);
nor U12526 (N_12526,N_11527,N_10624);
or U12527 (N_12527,N_10612,N_11284);
or U12528 (N_12528,N_11800,N_11026);
or U12529 (N_12529,N_10553,N_11250);
xor U12530 (N_12530,N_11748,N_11764);
nand U12531 (N_12531,N_11828,N_10854);
xor U12532 (N_12532,N_10890,N_10574);
nand U12533 (N_12533,N_10622,N_11034);
or U12534 (N_12534,N_11066,N_11152);
or U12535 (N_12535,N_10907,N_10812);
nand U12536 (N_12536,N_11134,N_11244);
nor U12537 (N_12537,N_11133,N_11975);
or U12538 (N_12538,N_11952,N_11787);
xor U12539 (N_12539,N_10868,N_11387);
or U12540 (N_12540,N_10916,N_11496);
xor U12541 (N_12541,N_10751,N_11964);
or U12542 (N_12542,N_10832,N_10952);
and U12543 (N_12543,N_10593,N_11202);
and U12544 (N_12544,N_11520,N_11490);
or U12545 (N_12545,N_11411,N_11218);
xor U12546 (N_12546,N_10703,N_11150);
and U12547 (N_12547,N_11686,N_11324);
or U12548 (N_12548,N_11491,N_11575);
and U12549 (N_12549,N_10999,N_11273);
and U12550 (N_12550,N_10849,N_11340);
and U12551 (N_12551,N_11667,N_11942);
xor U12552 (N_12552,N_10766,N_11189);
and U12553 (N_12553,N_10555,N_11725);
xnor U12554 (N_12554,N_10869,N_11165);
nand U12555 (N_12555,N_11885,N_11845);
nor U12556 (N_12556,N_11858,N_11500);
and U12557 (N_12557,N_10510,N_11142);
xnor U12558 (N_12558,N_11775,N_10735);
xor U12559 (N_12559,N_10749,N_10747);
or U12560 (N_12560,N_11030,N_11907);
or U12561 (N_12561,N_10610,N_10518);
or U12562 (N_12562,N_10968,N_11604);
xnor U12563 (N_12563,N_11394,N_11840);
nor U12564 (N_12564,N_11048,N_11696);
nand U12565 (N_12565,N_10618,N_11023);
and U12566 (N_12566,N_10645,N_11156);
xnor U12567 (N_12567,N_11896,N_11193);
or U12568 (N_12568,N_11716,N_11891);
xor U12569 (N_12569,N_10901,N_11170);
and U12570 (N_12570,N_11315,N_10859);
and U12571 (N_12571,N_11803,N_11237);
or U12572 (N_12572,N_11068,N_11105);
nand U12573 (N_12573,N_10626,N_11823);
and U12574 (N_12574,N_10776,N_10721);
or U12575 (N_12575,N_11418,N_10627);
or U12576 (N_12576,N_10536,N_11212);
nor U12577 (N_12577,N_10914,N_11179);
or U12578 (N_12578,N_11249,N_10746);
and U12579 (N_12579,N_11061,N_11191);
or U12580 (N_12580,N_11117,N_11445);
nand U12581 (N_12581,N_11739,N_10865);
or U12582 (N_12582,N_10840,N_11311);
nor U12583 (N_12583,N_11816,N_11149);
and U12584 (N_12584,N_10773,N_10683);
nand U12585 (N_12585,N_10841,N_10570);
and U12586 (N_12586,N_11531,N_11128);
and U12587 (N_12587,N_11813,N_11197);
nor U12588 (N_12588,N_11658,N_11972);
and U12589 (N_12589,N_11636,N_11809);
and U12590 (N_12590,N_10707,N_11256);
xor U12591 (N_12591,N_10900,N_11983);
and U12592 (N_12592,N_11158,N_10819);
or U12593 (N_12593,N_11548,N_10851);
and U12594 (N_12594,N_11617,N_11677);
nand U12595 (N_12595,N_11817,N_10788);
and U12596 (N_12596,N_11028,N_10826);
nor U12597 (N_12597,N_10969,N_11744);
xnor U12598 (N_12598,N_11431,N_11683);
xor U12599 (N_12599,N_11421,N_11838);
xor U12600 (N_12600,N_11381,N_11349);
nor U12601 (N_12601,N_11086,N_11107);
or U12602 (N_12602,N_11279,N_10984);
and U12603 (N_12603,N_11018,N_11956);
nor U12604 (N_12604,N_11203,N_11344);
nor U12605 (N_12605,N_11223,N_11754);
nand U12606 (N_12606,N_11920,N_11397);
nand U12607 (N_12607,N_10647,N_11619);
nor U12608 (N_12608,N_10807,N_11454);
xor U12609 (N_12609,N_10813,N_10681);
nor U12610 (N_12610,N_10797,N_11090);
or U12611 (N_12611,N_11060,N_11164);
xnor U12612 (N_12612,N_10587,N_11070);
or U12613 (N_12613,N_10882,N_10905);
nor U12614 (N_12614,N_10765,N_10877);
and U12615 (N_12615,N_10502,N_11190);
nor U12616 (N_12616,N_10519,N_11622);
xor U12617 (N_12617,N_11554,N_11036);
nand U12618 (N_12618,N_11430,N_11704);
nand U12619 (N_12619,N_11713,N_11360);
or U12620 (N_12620,N_10517,N_11444);
and U12621 (N_12621,N_11336,N_10906);
and U12622 (N_12622,N_10632,N_10828);
nand U12623 (N_12623,N_11406,N_11334);
and U12624 (N_12624,N_11378,N_10860);
nor U12625 (N_12625,N_10940,N_11352);
nor U12626 (N_12626,N_11013,N_10866);
or U12627 (N_12627,N_11643,N_11555);
xor U12628 (N_12628,N_11960,N_10547);
nor U12629 (N_12629,N_11166,N_11916);
nand U12630 (N_12630,N_11509,N_10625);
xnor U12631 (N_12631,N_10637,N_11077);
xor U12632 (N_12632,N_11294,N_10929);
nand U12633 (N_12633,N_10532,N_11114);
and U12634 (N_12634,N_11485,N_11377);
nand U12635 (N_12635,N_10565,N_11348);
nand U12636 (N_12636,N_11990,N_10586);
nand U12637 (N_12637,N_11477,N_11733);
nor U12638 (N_12638,N_11359,N_10719);
nor U12639 (N_12639,N_11537,N_11180);
nor U12640 (N_12640,N_11297,N_11732);
and U12641 (N_12641,N_10959,N_11425);
and U12642 (N_12642,N_11610,N_11698);
or U12643 (N_12643,N_11229,N_11866);
or U12644 (N_12644,N_11568,N_10786);
xnor U12645 (N_12645,N_11043,N_10552);
nand U12646 (N_12646,N_10998,N_11010);
nor U12647 (N_12647,N_10501,N_11493);
nor U12648 (N_12648,N_11738,N_11071);
and U12649 (N_12649,N_10513,N_11056);
xnor U12650 (N_12650,N_11159,N_10596);
nor U12651 (N_12651,N_11797,N_11634);
and U12652 (N_12652,N_11766,N_10516);
nor U12653 (N_12653,N_11507,N_11888);
and U12654 (N_12654,N_11919,N_11120);
xor U12655 (N_12655,N_11963,N_11850);
nor U12656 (N_12656,N_10763,N_11462);
or U12657 (N_12657,N_11291,N_11768);
or U12658 (N_12658,N_11089,N_10810);
nand U12659 (N_12659,N_11822,N_10963);
and U12660 (N_12660,N_11763,N_11616);
and U12661 (N_12661,N_11464,N_10917);
and U12662 (N_12662,N_11199,N_11498);
and U12663 (N_12663,N_11886,N_10824);
and U12664 (N_12664,N_11515,N_10569);
nand U12665 (N_12665,N_11316,N_10714);
nand U12666 (N_12666,N_11830,N_11151);
or U12667 (N_12667,N_11007,N_11442);
nand U12668 (N_12668,N_10601,N_11717);
or U12669 (N_12669,N_11724,N_11160);
xor U12670 (N_12670,N_11700,N_11264);
nand U12671 (N_12671,N_11665,N_11059);
nand U12672 (N_12672,N_11985,N_10894);
nand U12673 (N_12673,N_10862,N_11624);
nor U12674 (N_12674,N_11288,N_11436);
xnor U12675 (N_12675,N_11307,N_11702);
or U12676 (N_12676,N_11414,N_11040);
xor U12677 (N_12677,N_11547,N_11560);
nor U12678 (N_12678,N_11883,N_11820);
or U12679 (N_12679,N_11638,N_11875);
nor U12680 (N_12680,N_11124,N_11386);
and U12681 (N_12681,N_10589,N_11261);
and U12682 (N_12682,N_10676,N_11200);
nor U12683 (N_12683,N_11428,N_11054);
nand U12684 (N_12684,N_10603,N_10674);
nand U12685 (N_12685,N_11508,N_10926);
nand U12686 (N_12686,N_11553,N_10830);
or U12687 (N_12687,N_10867,N_10530);
and U12688 (N_12688,N_10777,N_11672);
xor U12689 (N_12689,N_10975,N_11217);
or U12690 (N_12690,N_10897,N_11879);
nor U12691 (N_12691,N_11660,N_11522);
and U12692 (N_12692,N_11914,N_11045);
xor U12693 (N_12693,N_11338,N_11623);
or U12694 (N_12694,N_11777,N_11926);
and U12695 (N_12695,N_10573,N_11935);
nand U12696 (N_12696,N_11892,N_11994);
nand U12697 (N_12697,N_11192,N_10966);
xor U12698 (N_12698,N_11019,N_11276);
or U12699 (N_12699,N_11796,N_11176);
nor U12700 (N_12700,N_11245,N_11727);
and U12701 (N_12701,N_10548,N_11167);
xor U12702 (N_12702,N_11461,N_10848);
or U12703 (N_12703,N_11608,N_11759);
or U12704 (N_12704,N_10754,N_10667);
nand U12705 (N_12705,N_11590,N_11440);
xor U12706 (N_12706,N_11064,N_11236);
nand U12707 (N_12707,N_10668,N_10524);
nor U12708 (N_12708,N_11293,N_11877);
nor U12709 (N_12709,N_11722,N_10534);
xnor U12710 (N_12710,N_10737,N_11794);
xor U12711 (N_12711,N_11659,N_11596);
xor U12712 (N_12712,N_10760,N_10505);
nand U12713 (N_12713,N_11723,N_11110);
xor U12714 (N_12714,N_11606,N_11986);
and U12715 (N_12715,N_11032,N_10561);
or U12716 (N_12716,N_11468,N_11476);
or U12717 (N_12717,N_10928,N_11323);
or U12718 (N_12718,N_10692,N_10595);
and U12719 (N_12719,N_11367,N_11662);
and U12720 (N_12720,N_11351,N_11589);
nor U12721 (N_12721,N_10816,N_11113);
nand U12722 (N_12722,N_11362,N_10526);
and U12723 (N_12723,N_11213,N_10655);
and U12724 (N_12724,N_11393,N_10814);
xor U12725 (N_12725,N_11561,N_11339);
or U12726 (N_12726,N_10563,N_11302);
nor U12727 (N_12727,N_11205,N_11305);
nor U12728 (N_12728,N_10671,N_11915);
nor U12729 (N_12729,N_10775,N_11106);
and U12730 (N_12730,N_10590,N_11904);
nand U12731 (N_12731,N_11314,N_11867);
and U12732 (N_12732,N_11758,N_10640);
nand U12733 (N_12733,N_10887,N_10896);
and U12734 (N_12734,N_11448,N_10672);
or U12735 (N_12735,N_10908,N_10594);
nand U12736 (N_12736,N_11053,N_11965);
nor U12737 (N_12737,N_11529,N_11544);
and U12738 (N_12738,N_11135,N_10888);
or U12739 (N_12739,N_11319,N_11163);
or U12740 (N_12740,N_11080,N_10931);
nor U12741 (N_12741,N_11592,N_11408);
xnor U12742 (N_12742,N_10701,N_11088);
nand U12743 (N_12743,N_11435,N_11852);
nor U12744 (N_12744,N_11453,N_11473);
nor U12745 (N_12745,N_11475,N_11680);
nand U12746 (N_12746,N_10949,N_11065);
nor U12747 (N_12747,N_10643,N_10720);
nand U12748 (N_12748,N_11958,N_11530);
nor U12749 (N_12749,N_11322,N_11571);
xor U12750 (N_12750,N_11491,N_11606);
xnor U12751 (N_12751,N_10512,N_10983);
xnor U12752 (N_12752,N_10955,N_10672);
nor U12753 (N_12753,N_10815,N_11313);
and U12754 (N_12754,N_11030,N_10595);
or U12755 (N_12755,N_11695,N_11698);
nand U12756 (N_12756,N_11743,N_11360);
xnor U12757 (N_12757,N_10961,N_10653);
and U12758 (N_12758,N_10645,N_11449);
and U12759 (N_12759,N_11160,N_11239);
or U12760 (N_12760,N_11577,N_10544);
or U12761 (N_12761,N_10897,N_10637);
and U12762 (N_12762,N_11302,N_11685);
xor U12763 (N_12763,N_11862,N_11916);
or U12764 (N_12764,N_11620,N_10545);
or U12765 (N_12765,N_10608,N_11550);
and U12766 (N_12766,N_10781,N_10652);
nor U12767 (N_12767,N_11166,N_11389);
nand U12768 (N_12768,N_11035,N_11698);
and U12769 (N_12769,N_11335,N_11035);
or U12770 (N_12770,N_11494,N_11701);
and U12771 (N_12771,N_11145,N_11245);
nand U12772 (N_12772,N_10889,N_11092);
and U12773 (N_12773,N_11517,N_10536);
and U12774 (N_12774,N_11250,N_11764);
or U12775 (N_12775,N_11307,N_10820);
and U12776 (N_12776,N_11252,N_11541);
nand U12777 (N_12777,N_10733,N_11304);
nor U12778 (N_12778,N_10527,N_11028);
xor U12779 (N_12779,N_11275,N_11690);
or U12780 (N_12780,N_10866,N_11687);
xor U12781 (N_12781,N_11907,N_11467);
or U12782 (N_12782,N_10507,N_11612);
xnor U12783 (N_12783,N_10788,N_10719);
and U12784 (N_12784,N_10812,N_10824);
xor U12785 (N_12785,N_10910,N_11358);
nand U12786 (N_12786,N_10835,N_11097);
and U12787 (N_12787,N_11829,N_11517);
or U12788 (N_12788,N_10542,N_11819);
xor U12789 (N_12789,N_11038,N_10565);
and U12790 (N_12790,N_11125,N_11518);
or U12791 (N_12791,N_11369,N_10806);
and U12792 (N_12792,N_10869,N_11780);
nor U12793 (N_12793,N_10967,N_10703);
or U12794 (N_12794,N_11557,N_11606);
nand U12795 (N_12795,N_11024,N_11210);
and U12796 (N_12796,N_11107,N_11119);
xnor U12797 (N_12797,N_11932,N_10990);
xnor U12798 (N_12798,N_10525,N_10941);
nor U12799 (N_12799,N_10578,N_10590);
nor U12800 (N_12800,N_10600,N_10843);
nand U12801 (N_12801,N_11770,N_11182);
nand U12802 (N_12802,N_11945,N_11871);
or U12803 (N_12803,N_11343,N_11835);
or U12804 (N_12804,N_11674,N_10543);
or U12805 (N_12805,N_11537,N_10989);
nor U12806 (N_12806,N_10737,N_11132);
and U12807 (N_12807,N_11464,N_11294);
nor U12808 (N_12808,N_11263,N_11512);
and U12809 (N_12809,N_10970,N_10898);
xor U12810 (N_12810,N_11430,N_11533);
nor U12811 (N_12811,N_11648,N_10539);
and U12812 (N_12812,N_11922,N_11180);
nor U12813 (N_12813,N_11767,N_10593);
xor U12814 (N_12814,N_11010,N_11395);
xnor U12815 (N_12815,N_10562,N_11569);
nand U12816 (N_12816,N_11055,N_11533);
xor U12817 (N_12817,N_11870,N_11808);
or U12818 (N_12818,N_10707,N_11258);
xnor U12819 (N_12819,N_11229,N_11280);
nand U12820 (N_12820,N_11486,N_11440);
or U12821 (N_12821,N_11793,N_11719);
and U12822 (N_12822,N_10989,N_11521);
or U12823 (N_12823,N_10656,N_10855);
and U12824 (N_12824,N_11698,N_11770);
nand U12825 (N_12825,N_11355,N_11963);
xor U12826 (N_12826,N_11843,N_11062);
xor U12827 (N_12827,N_10787,N_11457);
nor U12828 (N_12828,N_11379,N_11623);
nor U12829 (N_12829,N_11941,N_10997);
nand U12830 (N_12830,N_11273,N_11525);
or U12831 (N_12831,N_11209,N_11174);
or U12832 (N_12832,N_10769,N_11798);
nand U12833 (N_12833,N_11948,N_11677);
and U12834 (N_12834,N_11504,N_10996);
and U12835 (N_12835,N_11089,N_11043);
nand U12836 (N_12836,N_11952,N_11820);
and U12837 (N_12837,N_10530,N_11243);
xor U12838 (N_12838,N_10547,N_10751);
and U12839 (N_12839,N_10582,N_11420);
nand U12840 (N_12840,N_10991,N_11861);
nand U12841 (N_12841,N_10654,N_11937);
nand U12842 (N_12842,N_10829,N_10503);
nor U12843 (N_12843,N_11840,N_11740);
nor U12844 (N_12844,N_11728,N_11853);
or U12845 (N_12845,N_11477,N_11678);
nor U12846 (N_12846,N_11461,N_10829);
nor U12847 (N_12847,N_10926,N_10905);
nor U12848 (N_12848,N_10572,N_11189);
nor U12849 (N_12849,N_11721,N_11731);
or U12850 (N_12850,N_10991,N_11314);
nor U12851 (N_12851,N_10748,N_11048);
or U12852 (N_12852,N_10882,N_11899);
or U12853 (N_12853,N_11433,N_11664);
nand U12854 (N_12854,N_11883,N_11009);
nand U12855 (N_12855,N_10630,N_11848);
nand U12856 (N_12856,N_11642,N_11382);
nand U12857 (N_12857,N_11378,N_11198);
xor U12858 (N_12858,N_11958,N_11382);
nor U12859 (N_12859,N_11173,N_11401);
nand U12860 (N_12860,N_10548,N_10514);
nor U12861 (N_12861,N_10712,N_11396);
nor U12862 (N_12862,N_10915,N_11436);
xnor U12863 (N_12863,N_10616,N_10853);
nand U12864 (N_12864,N_10831,N_11470);
nand U12865 (N_12865,N_11597,N_11366);
or U12866 (N_12866,N_11110,N_10736);
or U12867 (N_12867,N_10745,N_10701);
nand U12868 (N_12868,N_10741,N_10670);
and U12869 (N_12869,N_11775,N_10918);
nor U12870 (N_12870,N_11978,N_11995);
and U12871 (N_12871,N_11904,N_11482);
or U12872 (N_12872,N_11039,N_11527);
and U12873 (N_12873,N_11662,N_11272);
nand U12874 (N_12874,N_11633,N_10578);
nor U12875 (N_12875,N_11100,N_10980);
xor U12876 (N_12876,N_11482,N_11193);
and U12877 (N_12877,N_11155,N_11029);
and U12878 (N_12878,N_10981,N_10889);
nor U12879 (N_12879,N_11491,N_10862);
nor U12880 (N_12880,N_11289,N_11038);
and U12881 (N_12881,N_11228,N_11853);
or U12882 (N_12882,N_10943,N_11893);
xor U12883 (N_12883,N_11354,N_10867);
and U12884 (N_12884,N_11630,N_10729);
nor U12885 (N_12885,N_11605,N_10802);
nor U12886 (N_12886,N_10910,N_11666);
and U12887 (N_12887,N_11293,N_11999);
nor U12888 (N_12888,N_11158,N_10845);
nor U12889 (N_12889,N_10634,N_11637);
nor U12890 (N_12890,N_10781,N_11236);
xnor U12891 (N_12891,N_11007,N_11956);
xor U12892 (N_12892,N_11700,N_10815);
and U12893 (N_12893,N_10555,N_11611);
nand U12894 (N_12894,N_11612,N_11253);
nor U12895 (N_12895,N_10653,N_11874);
xor U12896 (N_12896,N_10950,N_11390);
xor U12897 (N_12897,N_11008,N_10665);
xor U12898 (N_12898,N_11821,N_11005);
xor U12899 (N_12899,N_11974,N_11322);
nor U12900 (N_12900,N_10978,N_10727);
xnor U12901 (N_12901,N_10804,N_10922);
nor U12902 (N_12902,N_11321,N_10551);
or U12903 (N_12903,N_11454,N_10819);
nand U12904 (N_12904,N_11351,N_10706);
xnor U12905 (N_12905,N_11264,N_11361);
nor U12906 (N_12906,N_11196,N_11586);
nor U12907 (N_12907,N_11425,N_11210);
nand U12908 (N_12908,N_11498,N_11426);
xnor U12909 (N_12909,N_11240,N_10606);
nor U12910 (N_12910,N_10679,N_11427);
or U12911 (N_12911,N_11250,N_11067);
nor U12912 (N_12912,N_11895,N_11344);
nor U12913 (N_12913,N_11846,N_11856);
xnor U12914 (N_12914,N_11291,N_11784);
xor U12915 (N_12915,N_11135,N_11713);
xor U12916 (N_12916,N_10529,N_11997);
nand U12917 (N_12917,N_10783,N_11831);
xnor U12918 (N_12918,N_11999,N_11540);
nor U12919 (N_12919,N_10551,N_11006);
and U12920 (N_12920,N_11325,N_11859);
and U12921 (N_12921,N_10570,N_11375);
or U12922 (N_12922,N_11551,N_10735);
or U12923 (N_12923,N_10716,N_11272);
and U12924 (N_12924,N_11928,N_10698);
xnor U12925 (N_12925,N_11400,N_10585);
or U12926 (N_12926,N_11616,N_10581);
and U12927 (N_12927,N_10910,N_10877);
and U12928 (N_12928,N_11789,N_11701);
or U12929 (N_12929,N_10520,N_11758);
and U12930 (N_12930,N_11505,N_11399);
nand U12931 (N_12931,N_11056,N_11495);
xor U12932 (N_12932,N_11003,N_11745);
nor U12933 (N_12933,N_11515,N_11706);
nand U12934 (N_12934,N_11887,N_11855);
nand U12935 (N_12935,N_10922,N_10821);
and U12936 (N_12936,N_11686,N_10518);
nor U12937 (N_12937,N_11770,N_11132);
xnor U12938 (N_12938,N_10758,N_11368);
or U12939 (N_12939,N_11481,N_10871);
nand U12940 (N_12940,N_11939,N_11515);
xnor U12941 (N_12941,N_11357,N_11253);
nor U12942 (N_12942,N_11881,N_10549);
and U12943 (N_12943,N_11273,N_11014);
xor U12944 (N_12944,N_10629,N_10673);
xnor U12945 (N_12945,N_11828,N_11861);
or U12946 (N_12946,N_10936,N_10895);
nor U12947 (N_12947,N_11264,N_10924);
or U12948 (N_12948,N_11978,N_11464);
xnor U12949 (N_12949,N_10704,N_10799);
nand U12950 (N_12950,N_11963,N_11887);
nand U12951 (N_12951,N_11496,N_11069);
and U12952 (N_12952,N_10998,N_11400);
xor U12953 (N_12953,N_10740,N_10966);
xor U12954 (N_12954,N_10962,N_10980);
and U12955 (N_12955,N_11902,N_10556);
and U12956 (N_12956,N_11004,N_11628);
nand U12957 (N_12957,N_11419,N_11541);
nor U12958 (N_12958,N_11571,N_11303);
xnor U12959 (N_12959,N_11873,N_10689);
xnor U12960 (N_12960,N_10791,N_11162);
xnor U12961 (N_12961,N_10824,N_11467);
nor U12962 (N_12962,N_10832,N_11078);
nand U12963 (N_12963,N_10729,N_11956);
xor U12964 (N_12964,N_11165,N_11543);
or U12965 (N_12965,N_10536,N_11714);
and U12966 (N_12966,N_11232,N_10923);
xnor U12967 (N_12967,N_10811,N_11319);
nand U12968 (N_12968,N_11289,N_11302);
nor U12969 (N_12969,N_11845,N_10753);
nor U12970 (N_12970,N_11881,N_11942);
nand U12971 (N_12971,N_10743,N_11628);
and U12972 (N_12972,N_10986,N_11869);
nand U12973 (N_12973,N_11383,N_11667);
xor U12974 (N_12974,N_10927,N_11850);
nand U12975 (N_12975,N_10986,N_11083);
nand U12976 (N_12976,N_10994,N_11985);
and U12977 (N_12977,N_11748,N_10840);
or U12978 (N_12978,N_10531,N_10952);
xnor U12979 (N_12979,N_11515,N_11506);
nand U12980 (N_12980,N_10713,N_11643);
nand U12981 (N_12981,N_10531,N_10695);
nand U12982 (N_12982,N_10827,N_11152);
nor U12983 (N_12983,N_11975,N_11539);
nand U12984 (N_12984,N_11734,N_11314);
and U12985 (N_12985,N_11044,N_10553);
nor U12986 (N_12986,N_11391,N_11945);
and U12987 (N_12987,N_11500,N_10980);
and U12988 (N_12988,N_10711,N_11379);
or U12989 (N_12989,N_11881,N_10572);
nand U12990 (N_12990,N_11773,N_10923);
or U12991 (N_12991,N_11450,N_11272);
nor U12992 (N_12992,N_11836,N_10513);
nor U12993 (N_12993,N_10920,N_11463);
or U12994 (N_12994,N_11436,N_11088);
nor U12995 (N_12995,N_11055,N_10713);
xnor U12996 (N_12996,N_11451,N_11632);
xnor U12997 (N_12997,N_11123,N_10783);
xnor U12998 (N_12998,N_11470,N_10629);
and U12999 (N_12999,N_11192,N_11784);
xnor U13000 (N_13000,N_11771,N_10549);
nor U13001 (N_13001,N_11950,N_11022);
xnor U13002 (N_13002,N_11769,N_11372);
nand U13003 (N_13003,N_11995,N_11596);
xor U13004 (N_13004,N_10892,N_10857);
and U13005 (N_13005,N_10910,N_11436);
or U13006 (N_13006,N_10669,N_11962);
and U13007 (N_13007,N_11132,N_10597);
or U13008 (N_13008,N_10853,N_11566);
or U13009 (N_13009,N_10927,N_11125);
xnor U13010 (N_13010,N_10690,N_11982);
or U13011 (N_13011,N_11450,N_11689);
nand U13012 (N_13012,N_10790,N_11522);
or U13013 (N_13013,N_10740,N_11927);
xnor U13014 (N_13014,N_11623,N_10521);
and U13015 (N_13015,N_11039,N_11075);
nor U13016 (N_13016,N_11330,N_11966);
nand U13017 (N_13017,N_11643,N_11705);
nand U13018 (N_13018,N_11483,N_11276);
nor U13019 (N_13019,N_10923,N_10784);
xor U13020 (N_13020,N_10985,N_10805);
or U13021 (N_13021,N_10722,N_10735);
nor U13022 (N_13022,N_10838,N_11046);
and U13023 (N_13023,N_10877,N_11351);
nand U13024 (N_13024,N_11133,N_11224);
nand U13025 (N_13025,N_11523,N_10564);
nand U13026 (N_13026,N_11211,N_11026);
xor U13027 (N_13027,N_11559,N_10853);
or U13028 (N_13028,N_11774,N_11236);
nand U13029 (N_13029,N_10811,N_11746);
nor U13030 (N_13030,N_11336,N_10875);
nand U13031 (N_13031,N_11204,N_11054);
nor U13032 (N_13032,N_11671,N_11436);
nor U13033 (N_13033,N_10862,N_11666);
nand U13034 (N_13034,N_10799,N_11742);
nand U13035 (N_13035,N_11504,N_10793);
or U13036 (N_13036,N_11605,N_11010);
or U13037 (N_13037,N_10928,N_10710);
nand U13038 (N_13038,N_11029,N_10658);
or U13039 (N_13039,N_10812,N_11932);
nor U13040 (N_13040,N_11154,N_11802);
nand U13041 (N_13041,N_11041,N_10676);
or U13042 (N_13042,N_10756,N_10917);
nand U13043 (N_13043,N_11974,N_11401);
nor U13044 (N_13044,N_10562,N_10549);
and U13045 (N_13045,N_11804,N_11226);
and U13046 (N_13046,N_11671,N_10569);
or U13047 (N_13047,N_11685,N_11333);
xnor U13048 (N_13048,N_11188,N_11311);
xor U13049 (N_13049,N_11872,N_11219);
xor U13050 (N_13050,N_11940,N_11754);
and U13051 (N_13051,N_11142,N_11526);
nand U13052 (N_13052,N_11634,N_11457);
and U13053 (N_13053,N_11234,N_10951);
nand U13054 (N_13054,N_11863,N_11145);
nor U13055 (N_13055,N_11050,N_11279);
and U13056 (N_13056,N_10694,N_11528);
and U13057 (N_13057,N_11793,N_11474);
or U13058 (N_13058,N_10582,N_10782);
nand U13059 (N_13059,N_11504,N_10953);
nor U13060 (N_13060,N_11456,N_11731);
nand U13061 (N_13061,N_11473,N_11359);
nand U13062 (N_13062,N_11427,N_11394);
and U13063 (N_13063,N_11610,N_11073);
or U13064 (N_13064,N_11581,N_11176);
nand U13065 (N_13065,N_11059,N_11228);
nor U13066 (N_13066,N_10610,N_11569);
nand U13067 (N_13067,N_10564,N_11042);
nand U13068 (N_13068,N_10950,N_11312);
nor U13069 (N_13069,N_11177,N_11943);
and U13070 (N_13070,N_11364,N_11750);
or U13071 (N_13071,N_10549,N_11203);
nor U13072 (N_13072,N_11374,N_11914);
xnor U13073 (N_13073,N_11851,N_11307);
xor U13074 (N_13074,N_11460,N_11684);
nand U13075 (N_13075,N_11682,N_11464);
and U13076 (N_13076,N_10796,N_10560);
and U13077 (N_13077,N_11100,N_11005);
nand U13078 (N_13078,N_11936,N_11947);
xnor U13079 (N_13079,N_11029,N_11774);
nor U13080 (N_13080,N_10809,N_10747);
xor U13081 (N_13081,N_11159,N_10868);
nor U13082 (N_13082,N_11704,N_10906);
nand U13083 (N_13083,N_10555,N_10842);
nand U13084 (N_13084,N_10844,N_11897);
or U13085 (N_13085,N_10985,N_10946);
nand U13086 (N_13086,N_11225,N_10808);
nand U13087 (N_13087,N_11591,N_11708);
or U13088 (N_13088,N_11312,N_10506);
xnor U13089 (N_13089,N_11893,N_11299);
nand U13090 (N_13090,N_11621,N_10658);
and U13091 (N_13091,N_11665,N_11460);
xnor U13092 (N_13092,N_11599,N_10912);
and U13093 (N_13093,N_11048,N_11892);
nor U13094 (N_13094,N_11003,N_10557);
nor U13095 (N_13095,N_10864,N_11587);
nand U13096 (N_13096,N_11513,N_10831);
and U13097 (N_13097,N_10842,N_11772);
or U13098 (N_13098,N_11977,N_11376);
and U13099 (N_13099,N_11033,N_11264);
nand U13100 (N_13100,N_11971,N_10776);
nor U13101 (N_13101,N_11041,N_10661);
or U13102 (N_13102,N_11967,N_11109);
xnor U13103 (N_13103,N_10731,N_11932);
xor U13104 (N_13104,N_10806,N_10530);
nor U13105 (N_13105,N_11970,N_11204);
xor U13106 (N_13106,N_11498,N_11855);
nand U13107 (N_13107,N_10517,N_11661);
or U13108 (N_13108,N_10615,N_10666);
or U13109 (N_13109,N_11868,N_11510);
or U13110 (N_13110,N_11508,N_11715);
xor U13111 (N_13111,N_10751,N_11929);
xnor U13112 (N_13112,N_11463,N_11877);
nand U13113 (N_13113,N_11248,N_10808);
nor U13114 (N_13114,N_10852,N_11088);
nor U13115 (N_13115,N_10856,N_11485);
nor U13116 (N_13116,N_11726,N_11459);
xor U13117 (N_13117,N_10879,N_10884);
or U13118 (N_13118,N_11569,N_11348);
or U13119 (N_13119,N_11614,N_10889);
nand U13120 (N_13120,N_11771,N_11728);
or U13121 (N_13121,N_10720,N_11107);
or U13122 (N_13122,N_10572,N_10604);
and U13123 (N_13123,N_10552,N_10701);
and U13124 (N_13124,N_10820,N_11782);
nor U13125 (N_13125,N_10785,N_11000);
and U13126 (N_13126,N_11364,N_11413);
xor U13127 (N_13127,N_11324,N_11087);
or U13128 (N_13128,N_11796,N_11712);
or U13129 (N_13129,N_10824,N_11757);
and U13130 (N_13130,N_10713,N_11229);
nand U13131 (N_13131,N_10988,N_10954);
or U13132 (N_13132,N_11471,N_10774);
xor U13133 (N_13133,N_11545,N_11389);
nor U13134 (N_13134,N_11680,N_10700);
or U13135 (N_13135,N_10764,N_11371);
xnor U13136 (N_13136,N_10695,N_11322);
or U13137 (N_13137,N_11714,N_10939);
nor U13138 (N_13138,N_11370,N_11037);
nand U13139 (N_13139,N_11299,N_10711);
nor U13140 (N_13140,N_10876,N_11365);
and U13141 (N_13141,N_10997,N_11986);
nor U13142 (N_13142,N_11009,N_11451);
xnor U13143 (N_13143,N_11715,N_11490);
and U13144 (N_13144,N_11282,N_11263);
and U13145 (N_13145,N_11329,N_10554);
and U13146 (N_13146,N_11012,N_10940);
xnor U13147 (N_13147,N_11627,N_11769);
and U13148 (N_13148,N_10908,N_10990);
and U13149 (N_13149,N_11006,N_10775);
nand U13150 (N_13150,N_11280,N_11577);
and U13151 (N_13151,N_11910,N_11337);
xor U13152 (N_13152,N_11010,N_10891);
and U13153 (N_13153,N_11474,N_10903);
or U13154 (N_13154,N_11198,N_11149);
xor U13155 (N_13155,N_11276,N_10809);
nand U13156 (N_13156,N_10573,N_11303);
and U13157 (N_13157,N_11588,N_11264);
xor U13158 (N_13158,N_11480,N_10563);
xnor U13159 (N_13159,N_11774,N_10676);
or U13160 (N_13160,N_11814,N_11301);
xnor U13161 (N_13161,N_10729,N_11911);
and U13162 (N_13162,N_11637,N_10981);
nor U13163 (N_13163,N_11092,N_11352);
nor U13164 (N_13164,N_11913,N_10975);
nor U13165 (N_13165,N_10794,N_10606);
and U13166 (N_13166,N_11087,N_11209);
xnor U13167 (N_13167,N_11530,N_10777);
xnor U13168 (N_13168,N_11763,N_10726);
nand U13169 (N_13169,N_10873,N_10945);
xnor U13170 (N_13170,N_11915,N_11850);
xnor U13171 (N_13171,N_11821,N_11805);
nor U13172 (N_13172,N_11755,N_11910);
and U13173 (N_13173,N_11105,N_10956);
nand U13174 (N_13174,N_11753,N_10732);
and U13175 (N_13175,N_10714,N_11407);
and U13176 (N_13176,N_11462,N_10500);
and U13177 (N_13177,N_11526,N_11560);
xor U13178 (N_13178,N_10885,N_11042);
or U13179 (N_13179,N_11362,N_10582);
and U13180 (N_13180,N_11100,N_11009);
xor U13181 (N_13181,N_11033,N_11503);
nor U13182 (N_13182,N_11343,N_11778);
nor U13183 (N_13183,N_10586,N_11294);
nand U13184 (N_13184,N_11003,N_11013);
nor U13185 (N_13185,N_10702,N_11063);
and U13186 (N_13186,N_11272,N_11179);
and U13187 (N_13187,N_11310,N_10597);
nand U13188 (N_13188,N_11640,N_11856);
nand U13189 (N_13189,N_11992,N_10690);
nand U13190 (N_13190,N_11031,N_11026);
nor U13191 (N_13191,N_11369,N_11192);
and U13192 (N_13192,N_11862,N_11234);
or U13193 (N_13193,N_10689,N_11879);
xnor U13194 (N_13194,N_11862,N_10817);
xor U13195 (N_13195,N_11210,N_11428);
nor U13196 (N_13196,N_11593,N_10515);
nor U13197 (N_13197,N_11616,N_11683);
or U13198 (N_13198,N_11177,N_11424);
and U13199 (N_13199,N_10685,N_10831);
nor U13200 (N_13200,N_10544,N_11336);
nor U13201 (N_13201,N_11849,N_11391);
or U13202 (N_13202,N_11062,N_10923);
xnor U13203 (N_13203,N_11691,N_11502);
or U13204 (N_13204,N_11735,N_11361);
and U13205 (N_13205,N_10755,N_10741);
and U13206 (N_13206,N_11874,N_11002);
xnor U13207 (N_13207,N_10648,N_10533);
xor U13208 (N_13208,N_10730,N_10807);
or U13209 (N_13209,N_11283,N_11240);
or U13210 (N_13210,N_11635,N_10725);
or U13211 (N_13211,N_11031,N_11965);
nand U13212 (N_13212,N_11780,N_11706);
or U13213 (N_13213,N_11696,N_11088);
nor U13214 (N_13214,N_11773,N_11390);
nand U13215 (N_13215,N_10833,N_11162);
nor U13216 (N_13216,N_10645,N_11883);
nand U13217 (N_13217,N_11288,N_10827);
and U13218 (N_13218,N_11451,N_11342);
and U13219 (N_13219,N_11388,N_10875);
nand U13220 (N_13220,N_11833,N_11294);
and U13221 (N_13221,N_11880,N_11597);
nor U13222 (N_13222,N_11302,N_10971);
nor U13223 (N_13223,N_11439,N_11374);
and U13224 (N_13224,N_11684,N_10918);
xor U13225 (N_13225,N_11921,N_10619);
xnor U13226 (N_13226,N_11159,N_11868);
and U13227 (N_13227,N_11415,N_11171);
nand U13228 (N_13228,N_11218,N_11259);
or U13229 (N_13229,N_10716,N_11453);
or U13230 (N_13230,N_11161,N_10615);
xor U13231 (N_13231,N_11096,N_10520);
nor U13232 (N_13232,N_10624,N_10956);
xor U13233 (N_13233,N_11577,N_10886);
xnor U13234 (N_13234,N_11416,N_11541);
and U13235 (N_13235,N_11597,N_10673);
and U13236 (N_13236,N_10835,N_11276);
nor U13237 (N_13237,N_10777,N_10762);
nand U13238 (N_13238,N_11640,N_11679);
nand U13239 (N_13239,N_11118,N_11615);
nor U13240 (N_13240,N_11954,N_10812);
nand U13241 (N_13241,N_11796,N_11624);
nor U13242 (N_13242,N_11938,N_11300);
xnor U13243 (N_13243,N_10807,N_11561);
nand U13244 (N_13244,N_11773,N_11780);
nand U13245 (N_13245,N_11486,N_11430);
and U13246 (N_13246,N_11957,N_10960);
nor U13247 (N_13247,N_10961,N_11473);
xnor U13248 (N_13248,N_10523,N_10939);
xnor U13249 (N_13249,N_10792,N_11505);
nand U13250 (N_13250,N_11633,N_11863);
nor U13251 (N_13251,N_10772,N_11125);
or U13252 (N_13252,N_11245,N_11892);
nand U13253 (N_13253,N_11572,N_10756);
nand U13254 (N_13254,N_11386,N_11249);
nand U13255 (N_13255,N_11889,N_11180);
or U13256 (N_13256,N_11173,N_10614);
or U13257 (N_13257,N_11941,N_11272);
xor U13258 (N_13258,N_11004,N_11756);
xnor U13259 (N_13259,N_10785,N_11769);
or U13260 (N_13260,N_11955,N_11345);
or U13261 (N_13261,N_11064,N_11622);
xor U13262 (N_13262,N_11113,N_11436);
and U13263 (N_13263,N_10968,N_11894);
or U13264 (N_13264,N_11241,N_11734);
or U13265 (N_13265,N_11474,N_10809);
nand U13266 (N_13266,N_11460,N_10711);
nand U13267 (N_13267,N_10651,N_11002);
or U13268 (N_13268,N_10650,N_11161);
nand U13269 (N_13269,N_10713,N_11332);
or U13270 (N_13270,N_11430,N_10533);
nor U13271 (N_13271,N_11263,N_11745);
nand U13272 (N_13272,N_11955,N_11273);
or U13273 (N_13273,N_11370,N_11638);
and U13274 (N_13274,N_10786,N_10996);
nor U13275 (N_13275,N_11681,N_11345);
xor U13276 (N_13276,N_10810,N_11320);
xor U13277 (N_13277,N_11559,N_10527);
nand U13278 (N_13278,N_11096,N_11591);
or U13279 (N_13279,N_11454,N_10975);
xnor U13280 (N_13280,N_11324,N_11932);
nor U13281 (N_13281,N_10553,N_11789);
xor U13282 (N_13282,N_11806,N_10559);
or U13283 (N_13283,N_10718,N_11615);
or U13284 (N_13284,N_11667,N_11479);
and U13285 (N_13285,N_10715,N_11126);
nor U13286 (N_13286,N_11798,N_11768);
nor U13287 (N_13287,N_11442,N_11874);
nor U13288 (N_13288,N_10792,N_11802);
nor U13289 (N_13289,N_11886,N_10632);
and U13290 (N_13290,N_11415,N_11721);
nor U13291 (N_13291,N_11491,N_11364);
and U13292 (N_13292,N_11407,N_11526);
nor U13293 (N_13293,N_10906,N_11558);
xor U13294 (N_13294,N_11406,N_10912);
xor U13295 (N_13295,N_11668,N_11871);
and U13296 (N_13296,N_10896,N_11746);
and U13297 (N_13297,N_11544,N_11765);
xnor U13298 (N_13298,N_11132,N_11669);
and U13299 (N_13299,N_11980,N_11099);
nor U13300 (N_13300,N_10706,N_10686);
nor U13301 (N_13301,N_10776,N_10985);
or U13302 (N_13302,N_11831,N_11684);
and U13303 (N_13303,N_11358,N_10647);
nor U13304 (N_13304,N_11400,N_11865);
nor U13305 (N_13305,N_11867,N_10937);
nand U13306 (N_13306,N_10890,N_10614);
nand U13307 (N_13307,N_11485,N_11643);
xor U13308 (N_13308,N_11027,N_10650);
and U13309 (N_13309,N_11409,N_11207);
nor U13310 (N_13310,N_11274,N_11484);
or U13311 (N_13311,N_10957,N_10898);
nor U13312 (N_13312,N_11845,N_11697);
and U13313 (N_13313,N_11293,N_11681);
nor U13314 (N_13314,N_10568,N_11963);
nand U13315 (N_13315,N_10752,N_11511);
xor U13316 (N_13316,N_11310,N_10652);
xor U13317 (N_13317,N_11111,N_11219);
xor U13318 (N_13318,N_10783,N_10931);
or U13319 (N_13319,N_11890,N_11966);
or U13320 (N_13320,N_11374,N_11514);
or U13321 (N_13321,N_11617,N_11078);
xor U13322 (N_13322,N_11738,N_11268);
and U13323 (N_13323,N_11690,N_11838);
nand U13324 (N_13324,N_10541,N_10875);
or U13325 (N_13325,N_11443,N_10981);
xor U13326 (N_13326,N_11057,N_11448);
nor U13327 (N_13327,N_10667,N_11169);
xor U13328 (N_13328,N_11326,N_10596);
xnor U13329 (N_13329,N_11202,N_11025);
nor U13330 (N_13330,N_11527,N_11007);
xnor U13331 (N_13331,N_11693,N_10755);
nor U13332 (N_13332,N_10802,N_10812);
xor U13333 (N_13333,N_10656,N_11772);
and U13334 (N_13334,N_11961,N_11828);
and U13335 (N_13335,N_10604,N_11613);
nand U13336 (N_13336,N_11163,N_11987);
xor U13337 (N_13337,N_11384,N_10706);
or U13338 (N_13338,N_10940,N_11625);
nor U13339 (N_13339,N_10567,N_10535);
and U13340 (N_13340,N_10505,N_11262);
nand U13341 (N_13341,N_10779,N_11515);
or U13342 (N_13342,N_11155,N_11019);
or U13343 (N_13343,N_11848,N_11463);
or U13344 (N_13344,N_11213,N_11011);
nand U13345 (N_13345,N_10841,N_11359);
nand U13346 (N_13346,N_11242,N_11535);
or U13347 (N_13347,N_11567,N_11277);
xor U13348 (N_13348,N_11146,N_11613);
nand U13349 (N_13349,N_10661,N_11096);
xor U13350 (N_13350,N_11837,N_11550);
xor U13351 (N_13351,N_11778,N_10746);
or U13352 (N_13352,N_10865,N_11825);
or U13353 (N_13353,N_11504,N_11763);
nand U13354 (N_13354,N_11881,N_11012);
or U13355 (N_13355,N_11407,N_10991);
or U13356 (N_13356,N_11973,N_10840);
or U13357 (N_13357,N_11926,N_11887);
xor U13358 (N_13358,N_10920,N_10776);
nor U13359 (N_13359,N_10979,N_11881);
nor U13360 (N_13360,N_11423,N_11436);
or U13361 (N_13361,N_10951,N_11333);
xnor U13362 (N_13362,N_10907,N_10913);
and U13363 (N_13363,N_11279,N_11392);
nor U13364 (N_13364,N_10834,N_11121);
nor U13365 (N_13365,N_10702,N_11443);
and U13366 (N_13366,N_10667,N_11028);
or U13367 (N_13367,N_10815,N_11586);
nand U13368 (N_13368,N_11245,N_11143);
nand U13369 (N_13369,N_10572,N_11833);
or U13370 (N_13370,N_11721,N_11965);
or U13371 (N_13371,N_11740,N_10606);
and U13372 (N_13372,N_11583,N_11862);
xnor U13373 (N_13373,N_11962,N_10924);
nor U13374 (N_13374,N_11342,N_11537);
and U13375 (N_13375,N_11210,N_11171);
nand U13376 (N_13376,N_10901,N_11617);
nor U13377 (N_13377,N_11678,N_10647);
nor U13378 (N_13378,N_11168,N_11409);
nor U13379 (N_13379,N_11858,N_11211);
or U13380 (N_13380,N_11902,N_11436);
and U13381 (N_13381,N_10862,N_10696);
nor U13382 (N_13382,N_11816,N_11792);
nor U13383 (N_13383,N_11788,N_11222);
xor U13384 (N_13384,N_10640,N_11442);
xnor U13385 (N_13385,N_10961,N_10530);
and U13386 (N_13386,N_11643,N_11289);
nand U13387 (N_13387,N_11882,N_10980);
and U13388 (N_13388,N_10753,N_10530);
nand U13389 (N_13389,N_11813,N_11042);
xor U13390 (N_13390,N_10583,N_11124);
or U13391 (N_13391,N_10574,N_11791);
nor U13392 (N_13392,N_11843,N_11803);
xor U13393 (N_13393,N_11134,N_10710);
or U13394 (N_13394,N_11288,N_11484);
xor U13395 (N_13395,N_10723,N_11574);
nand U13396 (N_13396,N_11004,N_11569);
or U13397 (N_13397,N_10842,N_11372);
and U13398 (N_13398,N_11411,N_10984);
nand U13399 (N_13399,N_11955,N_10688);
nand U13400 (N_13400,N_11640,N_11052);
nor U13401 (N_13401,N_11191,N_10581);
nand U13402 (N_13402,N_11024,N_11808);
or U13403 (N_13403,N_10873,N_10704);
nand U13404 (N_13404,N_11466,N_10825);
xnor U13405 (N_13405,N_11960,N_11433);
nor U13406 (N_13406,N_10594,N_11364);
nand U13407 (N_13407,N_10717,N_10828);
nand U13408 (N_13408,N_10959,N_11662);
and U13409 (N_13409,N_11062,N_11916);
and U13410 (N_13410,N_11359,N_11787);
nor U13411 (N_13411,N_10508,N_10509);
and U13412 (N_13412,N_11617,N_11025);
nand U13413 (N_13413,N_11849,N_10595);
xnor U13414 (N_13414,N_11696,N_11961);
nor U13415 (N_13415,N_11606,N_10558);
nand U13416 (N_13416,N_11673,N_11306);
nand U13417 (N_13417,N_11657,N_11538);
and U13418 (N_13418,N_11112,N_11921);
and U13419 (N_13419,N_11330,N_10898);
nand U13420 (N_13420,N_11290,N_10512);
nand U13421 (N_13421,N_10908,N_11699);
or U13422 (N_13422,N_11628,N_11062);
nor U13423 (N_13423,N_10633,N_10956);
or U13424 (N_13424,N_11990,N_10662);
nor U13425 (N_13425,N_10559,N_11164);
and U13426 (N_13426,N_10577,N_11626);
xnor U13427 (N_13427,N_11472,N_11111);
or U13428 (N_13428,N_10758,N_11061);
xor U13429 (N_13429,N_10969,N_10650);
nor U13430 (N_13430,N_10898,N_11059);
nand U13431 (N_13431,N_11094,N_11245);
xor U13432 (N_13432,N_11928,N_10718);
or U13433 (N_13433,N_10678,N_11064);
nor U13434 (N_13434,N_10772,N_11887);
and U13435 (N_13435,N_10510,N_10505);
or U13436 (N_13436,N_11797,N_11120);
xor U13437 (N_13437,N_10523,N_11705);
xor U13438 (N_13438,N_11154,N_10888);
nor U13439 (N_13439,N_11555,N_11195);
or U13440 (N_13440,N_10956,N_11140);
nor U13441 (N_13441,N_10752,N_11076);
nand U13442 (N_13442,N_10818,N_11529);
and U13443 (N_13443,N_11402,N_10540);
nor U13444 (N_13444,N_10506,N_11621);
and U13445 (N_13445,N_11384,N_11900);
nor U13446 (N_13446,N_10856,N_11427);
nor U13447 (N_13447,N_10580,N_11474);
nor U13448 (N_13448,N_10975,N_11101);
xor U13449 (N_13449,N_10597,N_10570);
nand U13450 (N_13450,N_10862,N_10812);
nand U13451 (N_13451,N_10531,N_10915);
nand U13452 (N_13452,N_11521,N_11952);
and U13453 (N_13453,N_11557,N_11270);
nor U13454 (N_13454,N_11566,N_10898);
nor U13455 (N_13455,N_10951,N_10677);
nor U13456 (N_13456,N_11750,N_10585);
xor U13457 (N_13457,N_11281,N_11242);
nand U13458 (N_13458,N_10555,N_11050);
and U13459 (N_13459,N_11323,N_11824);
or U13460 (N_13460,N_10627,N_11844);
and U13461 (N_13461,N_11881,N_11533);
nand U13462 (N_13462,N_11483,N_10501);
and U13463 (N_13463,N_10528,N_10853);
or U13464 (N_13464,N_11288,N_11040);
and U13465 (N_13465,N_10512,N_10841);
and U13466 (N_13466,N_10807,N_10907);
nor U13467 (N_13467,N_11294,N_10810);
nor U13468 (N_13468,N_11201,N_11725);
nor U13469 (N_13469,N_11799,N_11893);
or U13470 (N_13470,N_10613,N_11989);
xor U13471 (N_13471,N_11199,N_11995);
or U13472 (N_13472,N_11036,N_11169);
nand U13473 (N_13473,N_11062,N_10596);
nor U13474 (N_13474,N_10541,N_11195);
nor U13475 (N_13475,N_11367,N_11560);
and U13476 (N_13476,N_11131,N_10961);
nand U13477 (N_13477,N_11259,N_10508);
nor U13478 (N_13478,N_11534,N_11390);
and U13479 (N_13479,N_11986,N_10966);
nor U13480 (N_13480,N_10507,N_11545);
and U13481 (N_13481,N_11658,N_10959);
nand U13482 (N_13482,N_11826,N_11768);
and U13483 (N_13483,N_11621,N_11680);
nor U13484 (N_13484,N_11315,N_10935);
xnor U13485 (N_13485,N_10947,N_11735);
xor U13486 (N_13486,N_10537,N_10781);
xnor U13487 (N_13487,N_11888,N_10946);
or U13488 (N_13488,N_11704,N_11079);
nand U13489 (N_13489,N_11306,N_11777);
and U13490 (N_13490,N_11665,N_11835);
and U13491 (N_13491,N_11689,N_11686);
xnor U13492 (N_13492,N_10904,N_11499);
xor U13493 (N_13493,N_10992,N_11703);
nand U13494 (N_13494,N_11502,N_11734);
nand U13495 (N_13495,N_11248,N_10853);
or U13496 (N_13496,N_11654,N_11049);
xnor U13497 (N_13497,N_11177,N_10679);
xnor U13498 (N_13498,N_11451,N_11701);
nand U13499 (N_13499,N_11241,N_11313);
or U13500 (N_13500,N_13120,N_13008);
xor U13501 (N_13501,N_12237,N_12182);
nor U13502 (N_13502,N_12584,N_12671);
nor U13503 (N_13503,N_12355,N_13459);
nor U13504 (N_13504,N_12401,N_12185);
or U13505 (N_13505,N_13311,N_12985);
or U13506 (N_13506,N_13091,N_12716);
xnor U13507 (N_13507,N_12774,N_12411);
xnor U13508 (N_13508,N_12142,N_12277);
or U13509 (N_13509,N_13109,N_12440);
or U13510 (N_13510,N_12839,N_12112);
nand U13511 (N_13511,N_13148,N_13201);
or U13512 (N_13512,N_12626,N_13105);
and U13513 (N_13513,N_12271,N_13488);
nor U13514 (N_13514,N_13328,N_13001);
nor U13515 (N_13515,N_12836,N_13106);
nor U13516 (N_13516,N_12991,N_13002);
and U13517 (N_13517,N_12867,N_12254);
and U13518 (N_13518,N_13213,N_13416);
nor U13519 (N_13519,N_12431,N_12856);
and U13520 (N_13520,N_12187,N_13358);
nor U13521 (N_13521,N_13455,N_13077);
and U13522 (N_13522,N_12339,N_12345);
nand U13523 (N_13523,N_12283,N_12654);
and U13524 (N_13524,N_12305,N_12398);
nand U13525 (N_13525,N_12700,N_12371);
nand U13526 (N_13526,N_13344,N_13449);
xnor U13527 (N_13527,N_12472,N_13273);
nand U13528 (N_13528,N_12622,N_12065);
xor U13529 (N_13529,N_13014,N_12047);
and U13530 (N_13530,N_13301,N_13048);
nand U13531 (N_13531,N_12178,N_12586);
and U13532 (N_13532,N_13317,N_12155);
and U13533 (N_13533,N_12738,N_12282);
and U13534 (N_13534,N_12427,N_12695);
nand U13535 (N_13535,N_12138,N_13007);
nor U13536 (N_13536,N_13132,N_12893);
nand U13537 (N_13537,N_12368,N_12081);
xor U13538 (N_13538,N_13355,N_12354);
or U13539 (N_13539,N_12367,N_12147);
and U13540 (N_13540,N_13394,N_12559);
xor U13541 (N_13541,N_13202,N_12754);
xor U13542 (N_13542,N_12548,N_12640);
or U13543 (N_13543,N_13232,N_12811);
xnor U13544 (N_13544,N_13451,N_13147);
xor U13545 (N_13545,N_12188,N_12685);
and U13546 (N_13546,N_12647,N_12930);
and U13547 (N_13547,N_13432,N_12702);
and U13548 (N_13548,N_12909,N_12012);
xnor U13549 (N_13549,N_13239,N_13021);
xor U13550 (N_13550,N_12847,N_12332);
or U13551 (N_13551,N_12657,N_12574);
nand U13552 (N_13552,N_12883,N_12973);
nand U13553 (N_13553,N_13217,N_12236);
and U13554 (N_13554,N_12061,N_12826);
or U13555 (N_13555,N_13012,N_13032);
nand U13556 (N_13556,N_13495,N_12203);
and U13557 (N_13557,N_12479,N_13454);
and U13558 (N_13558,N_13203,N_13298);
nand U13559 (N_13559,N_12004,N_12334);
or U13560 (N_13560,N_13238,N_12885);
or U13561 (N_13561,N_12285,N_12200);
and U13562 (N_13562,N_12321,N_12891);
nor U13563 (N_13563,N_13304,N_13268);
xor U13564 (N_13564,N_12257,N_12797);
xnor U13565 (N_13565,N_12230,N_13179);
nand U13566 (N_13566,N_12504,N_12944);
or U13567 (N_13567,N_12445,N_12787);
xnor U13568 (N_13568,N_12425,N_13445);
and U13569 (N_13569,N_12999,N_12307);
nand U13570 (N_13570,N_13023,N_12825);
nor U13571 (N_13571,N_12190,N_12711);
nor U13572 (N_13572,N_12184,N_13128);
nand U13573 (N_13573,N_12405,N_12473);
xnor U13574 (N_13574,N_13189,N_13039);
nor U13575 (N_13575,N_12884,N_12925);
and U13576 (N_13576,N_12670,N_12476);
xor U13577 (N_13577,N_13093,N_13061);
xnor U13578 (N_13578,N_12980,N_12165);
or U13579 (N_13579,N_12274,N_12007);
nand U13580 (N_13580,N_12364,N_13255);
nand U13581 (N_13581,N_12673,N_12432);
nor U13582 (N_13582,N_12508,N_13422);
and U13583 (N_13583,N_12820,N_12128);
nor U13584 (N_13584,N_12728,N_12869);
xor U13585 (N_13585,N_13030,N_13045);
or U13586 (N_13586,N_13052,N_12886);
and U13587 (N_13587,N_13417,N_12535);
or U13588 (N_13588,N_12131,N_13053);
nor U13589 (N_13589,N_12449,N_12400);
and U13590 (N_13590,N_12189,N_13152);
nor U13591 (N_13591,N_12926,N_13080);
and U13592 (N_13592,N_12122,N_12620);
nor U13593 (N_13593,N_13293,N_12556);
nor U13594 (N_13594,N_12388,N_12998);
and U13595 (N_13595,N_12665,N_13302);
xnor U13596 (N_13596,N_12444,N_12846);
nor U13597 (N_13597,N_12934,N_12323);
or U13598 (N_13598,N_12870,N_12162);
xor U13599 (N_13599,N_12526,N_13240);
or U13600 (N_13600,N_12749,N_12814);
nand U13601 (N_13601,N_12319,N_13050);
and U13602 (N_13602,N_12880,N_12901);
nand U13603 (N_13603,N_12854,N_12874);
xnor U13604 (N_13604,N_12730,N_12404);
or U13605 (N_13605,N_12239,N_12519);
xor U13606 (N_13606,N_12067,N_13402);
nand U13607 (N_13607,N_13327,N_12450);
nor U13608 (N_13608,N_13252,N_13149);
or U13609 (N_13609,N_13462,N_13191);
or U13610 (N_13610,N_13139,N_13427);
nor U13611 (N_13611,N_12322,N_13108);
nand U13612 (N_13612,N_12558,N_12923);
and U13613 (N_13613,N_12579,N_13281);
or U13614 (N_13614,N_13164,N_13308);
nor U13615 (N_13615,N_13448,N_12443);
or U13616 (N_13616,N_12139,N_12624);
nor U13617 (N_13617,N_12872,N_12933);
or U13618 (N_13618,N_12484,N_13010);
and U13619 (N_13619,N_13218,N_13401);
nand U13620 (N_13620,N_12534,N_12659);
nor U13621 (N_13621,N_13078,N_13107);
nor U13622 (N_13622,N_12598,N_12919);
or U13623 (N_13623,N_13151,N_13435);
xor U13624 (N_13624,N_12114,N_12894);
nand U13625 (N_13625,N_12402,N_13387);
and U13626 (N_13626,N_12549,N_13250);
xnor U13627 (N_13627,N_12546,N_12003);
or U13628 (N_13628,N_12454,N_12758);
nand U13629 (N_13629,N_12756,N_12866);
nand U13630 (N_13630,N_12570,N_12107);
xor U13631 (N_13631,N_12699,N_12186);
or U13632 (N_13632,N_13270,N_12972);
nor U13633 (N_13633,N_12161,N_12168);
and U13634 (N_13634,N_12206,N_12042);
or U13635 (N_13635,N_12532,N_12198);
and U13636 (N_13636,N_12209,N_12785);
nor U13637 (N_13637,N_12648,N_12602);
nand U13638 (N_13638,N_12053,N_12135);
nand U13639 (N_13639,N_12093,N_12480);
xor U13640 (N_13640,N_13354,N_12735);
nor U13641 (N_13641,N_12151,N_12140);
or U13642 (N_13642,N_12050,N_12056);
nand U13643 (N_13643,N_12447,N_13366);
nor U13644 (N_13644,N_12009,N_12238);
and U13645 (N_13645,N_12038,N_12896);
nor U13646 (N_13646,N_12594,N_13058);
or U13647 (N_13647,N_12745,N_13400);
nor U13648 (N_13648,N_12538,N_13085);
nand U13649 (N_13649,N_12195,N_12290);
nand U13650 (N_13650,N_12907,N_13340);
and U13651 (N_13651,N_12459,N_12658);
or U13652 (N_13652,N_12023,N_12929);
nand U13653 (N_13653,N_13076,N_12679);
or U13654 (N_13654,N_12714,N_12202);
and U13655 (N_13655,N_12393,N_13277);
and U13656 (N_13656,N_12036,N_12396);
and U13657 (N_13657,N_12218,N_13011);
nand U13658 (N_13658,N_12408,N_12046);
nand U13659 (N_13659,N_13087,N_13180);
nor U13660 (N_13660,N_12750,N_12248);
nor U13661 (N_13661,N_13230,N_12493);
nor U13662 (N_13662,N_12337,N_12706);
or U13663 (N_13663,N_12413,N_12922);
and U13664 (N_13664,N_13113,N_13028);
or U13665 (N_13665,N_12041,N_12981);
nand U13666 (N_13666,N_12530,N_12642);
nor U13667 (N_13667,N_12076,N_12066);
nor U13668 (N_13668,N_13169,N_12013);
nor U13669 (N_13669,N_12935,N_12724);
and U13670 (N_13670,N_12808,N_12429);
or U13671 (N_13671,N_12439,N_13018);
and U13672 (N_13672,N_12361,N_13064);
or U13673 (N_13673,N_12563,N_12800);
xnor U13674 (N_13674,N_13090,N_12552);
or U13675 (N_13675,N_12469,N_12518);
or U13676 (N_13676,N_13300,N_13225);
nand U13677 (N_13677,N_12234,N_13258);
nand U13678 (N_13678,N_12099,N_12194);
and U13679 (N_13679,N_12106,N_13296);
and U13680 (N_13680,N_12996,N_12180);
or U13681 (N_13681,N_12141,N_12683);
and U13682 (N_13682,N_12680,N_12232);
and U13683 (N_13683,N_12297,N_12284);
and U13684 (N_13684,N_12214,N_13026);
nand U13685 (N_13685,N_12366,N_12158);
and U13686 (N_13686,N_13471,N_12689);
nor U13687 (N_13687,N_13036,N_12416);
xor U13688 (N_13688,N_13465,N_12941);
xor U13689 (N_13689,N_13484,N_12089);
and U13690 (N_13690,N_12357,N_13319);
or U13691 (N_13691,N_12636,N_13166);
nand U13692 (N_13692,N_13464,N_13329);
xnor U13693 (N_13693,N_12614,N_13360);
nor U13694 (N_13694,N_12294,N_13443);
or U13695 (N_13695,N_12129,N_12824);
or U13696 (N_13696,N_13346,N_12028);
nor U13697 (N_13697,N_13364,N_13199);
nand U13698 (N_13698,N_12729,N_12585);
and U13699 (N_13699,N_12537,N_12390);
and U13700 (N_13700,N_12174,N_12641);
nand U13701 (N_13701,N_12557,N_12664);
nand U13702 (N_13702,N_12747,N_12086);
xor U13703 (N_13703,N_12491,N_13075);
and U13704 (N_13704,N_12740,N_13129);
nor U13705 (N_13705,N_13242,N_13384);
or U13706 (N_13706,N_12529,N_13428);
and U13707 (N_13707,N_13216,N_13003);
and U13708 (N_13708,N_12804,N_13423);
and U13709 (N_13709,N_12525,N_12208);
nand U13710 (N_13710,N_12247,N_13368);
and U13711 (N_13711,N_13375,N_12022);
xnor U13712 (N_13712,N_13352,N_12121);
xor U13713 (N_13713,N_12270,N_12603);
xnor U13714 (N_13714,N_12905,N_12341);
and U13715 (N_13715,N_12815,N_12913);
or U13716 (N_13716,N_12109,N_13224);
nor U13717 (N_13717,N_13051,N_12181);
and U13718 (N_13718,N_12650,N_12881);
and U13719 (N_13719,N_13156,N_12490);
and U13720 (N_13720,N_12362,N_13100);
and U13721 (N_13721,N_12852,N_13309);
nand U13722 (N_13722,N_12115,N_13292);
nand U13723 (N_13723,N_12566,N_12433);
or U13724 (N_13724,N_12687,N_12349);
xnor U13725 (N_13725,N_12569,N_12327);
and U13726 (N_13726,N_13290,N_12233);
xor U13727 (N_13727,N_12144,N_13294);
nor U13728 (N_13728,N_13497,N_12353);
and U13729 (N_13729,N_12732,N_12019);
nand U13730 (N_13730,N_12596,N_13378);
or U13731 (N_13731,N_12211,N_12506);
and U13732 (N_13732,N_12564,N_12261);
or U13733 (N_13733,N_12851,N_13284);
and U13734 (N_13734,N_12250,N_13135);
nand U13735 (N_13735,N_12495,N_13372);
nand U13736 (N_13736,N_12701,N_13125);
nand U13737 (N_13737,N_12799,N_12103);
and U13738 (N_13738,N_12489,N_12173);
xor U13739 (N_13739,N_12948,N_12111);
xnor U13740 (N_13740,N_12821,N_12352);
and U13741 (N_13741,N_12742,N_12164);
xor U13742 (N_13742,N_12527,N_12474);
nor U13743 (N_13743,N_13483,N_12336);
nand U13744 (N_13744,N_13338,N_12049);
nor U13745 (N_13745,N_13193,N_12436);
or U13746 (N_13746,N_13493,N_12617);
and U13747 (N_13747,N_12054,N_12079);
or U13748 (N_13748,N_12682,N_12623);
and U13749 (N_13749,N_13110,N_12782);
and U13750 (N_13750,N_12374,N_12365);
and U13751 (N_13751,N_12906,N_12840);
nand U13752 (N_13752,N_13331,N_12545);
and U13753 (N_13753,N_12762,N_13207);
xnor U13754 (N_13754,N_12987,N_12844);
and U13755 (N_13755,N_13192,N_12798);
nor U13756 (N_13756,N_12150,N_12976);
nor U13757 (N_13757,N_12838,N_12561);
nand U13758 (N_13758,N_13006,N_12104);
nor U13759 (N_13759,N_12707,N_13289);
and U13760 (N_13760,N_13337,N_12006);
xnor U13761 (N_13761,N_12582,N_12997);
nand U13762 (N_13762,N_13343,N_13243);
nand U13763 (N_13763,N_12958,N_12389);
xor U13764 (N_13764,N_13138,N_12229);
nand U13765 (N_13765,N_12739,N_12580);
nand U13766 (N_13766,N_12303,N_12088);
nand U13767 (N_13767,N_13130,N_12394);
and U13768 (N_13768,N_12021,N_12817);
nand U13769 (N_13769,N_13220,N_13379);
and U13770 (N_13770,N_13414,N_13066);
and U13771 (N_13771,N_13163,N_12646);
nor U13772 (N_13772,N_12809,N_12843);
nor U13773 (N_13773,N_13084,N_12720);
xor U13774 (N_13774,N_12075,N_12967);
xnor U13775 (N_13775,N_13196,N_13334);
and U13776 (N_13776,N_12426,N_13278);
nor U13777 (N_13777,N_13453,N_12253);
nor U13778 (N_13778,N_13382,N_12986);
and U13779 (N_13779,N_12152,N_12159);
xor U13780 (N_13780,N_12882,N_12509);
nand U13781 (N_13781,N_12153,N_13131);
and U13782 (N_13782,N_12604,N_13208);
nand U13783 (N_13783,N_13436,N_12118);
or U13784 (N_13784,N_12904,N_12663);
xor U13785 (N_13785,N_12638,N_12568);
nor U13786 (N_13786,N_12678,N_12016);
and U13787 (N_13787,N_12764,N_12289);
and U13788 (N_13788,N_13370,N_12567);
or U13789 (N_13789,N_13441,N_12171);
xnor U13790 (N_13790,N_13380,N_13330);
nor U13791 (N_13791,N_12192,N_12094);
and U13792 (N_13792,N_13212,N_12618);
or U13793 (N_13793,N_12116,N_12793);
nand U13794 (N_13794,N_12029,N_12910);
nand U13795 (N_13795,N_13275,N_12377);
and U13796 (N_13796,N_13494,N_13349);
xnor U13797 (N_13797,N_13305,N_13412);
nand U13798 (N_13798,N_12358,N_13430);
or U13799 (N_13799,N_12412,N_12373);
nand U13800 (N_13800,N_13286,N_12727);
and U13801 (N_13801,N_12252,N_13282);
xnor U13802 (N_13802,N_12132,N_13403);
nor U13803 (N_13803,N_12768,N_12212);
nand U13804 (N_13804,N_13150,N_12746);
xor U13805 (N_13805,N_13117,N_12228);
and U13806 (N_13806,N_13063,N_13119);
nor U13807 (N_13807,N_12778,N_12421);
and U13808 (N_13808,N_13404,N_12571);
xnor U13809 (N_13809,N_12576,N_12256);
and U13810 (N_13810,N_12026,N_12483);
nand U13811 (N_13811,N_12481,N_12951);
xnor U13812 (N_13812,N_12759,N_12397);
or U13813 (N_13813,N_12235,N_12818);
and U13814 (N_13814,N_12514,N_12786);
or U13815 (N_13815,N_12040,N_12502);
nor U13816 (N_13816,N_12722,N_12417);
or U13817 (N_13817,N_12877,N_12988);
nand U13818 (N_13818,N_12064,N_12387);
or U13819 (N_13819,N_13348,N_12062);
xor U13820 (N_13820,N_12403,N_13136);
xnor U13821 (N_13821,N_13060,N_12243);
nor U13822 (N_13822,N_13478,N_13234);
nand U13823 (N_13823,N_13496,N_12515);
nor U13824 (N_13824,N_13457,N_12299);
nor U13825 (N_13825,N_12020,N_12110);
nand U13826 (N_13826,N_13272,N_12581);
xor U13827 (N_13827,N_12938,N_13127);
xor U13828 (N_13828,N_13211,N_12900);
nand U13829 (N_13829,N_12555,N_12953);
xor U13830 (N_13830,N_13178,N_13433);
xnor U13831 (N_13831,N_13069,N_13418);
nor U13832 (N_13832,N_12466,N_13126);
xor U13833 (N_13833,N_13173,N_13195);
xor U13834 (N_13834,N_12773,N_12547);
or U13835 (N_13835,N_12386,N_12292);
nor U13836 (N_13836,N_13235,N_13279);
nor U13837 (N_13837,N_13313,N_12697);
nand U13838 (N_13838,N_12704,N_13361);
or U13839 (N_13839,N_13363,N_12608);
or U13840 (N_13840,N_13046,N_13054);
or U13841 (N_13841,N_13137,N_12002);
nor U13842 (N_13842,N_12338,N_13068);
nor U13843 (N_13843,N_12280,N_12419);
nor U13844 (N_13844,N_13016,N_12677);
and U13845 (N_13845,N_12968,N_13262);
nand U13846 (N_13846,N_12462,N_13231);
xnor U13847 (N_13847,N_12272,N_12903);
xnor U13848 (N_13848,N_13165,N_13185);
and U13849 (N_13849,N_12875,N_13024);
or U13850 (N_13850,N_12709,N_12937);
and U13851 (N_13851,N_12315,N_13095);
or U13852 (N_13852,N_13221,N_12898);
nor U13853 (N_13853,N_12792,N_12035);
and U13854 (N_13854,N_13477,N_12308);
or U13855 (N_13855,N_13020,N_12849);
and U13856 (N_13856,N_13473,N_12989);
nand U13857 (N_13857,N_12583,N_13439);
nand U13858 (N_13858,N_13038,N_12959);
and U13859 (N_13859,N_12892,N_12616);
nand U13860 (N_13860,N_12126,N_13197);
nand U13861 (N_13861,N_13303,N_12897);
or U13862 (N_13862,N_13246,N_12442);
nor U13863 (N_13863,N_12298,N_12995);
and U13864 (N_13864,N_13381,N_12227);
nor U13865 (N_13865,N_12266,N_12333);
nand U13866 (N_13866,N_12231,N_12105);
nor U13867 (N_13867,N_12060,N_12376);
xor U13868 (N_13868,N_12521,N_12775);
nand U13869 (N_13869,N_12130,N_12761);
and U13870 (N_13870,N_12781,N_12179);
and U13871 (N_13871,N_13415,N_12096);
nand U13872 (N_13872,N_13490,N_13092);
nor U13873 (N_13873,N_13489,N_12176);
and U13874 (N_13874,N_12908,N_13411);
xnor U13875 (N_13875,N_12541,N_13316);
or U13876 (N_13876,N_12291,N_12656);
and U13877 (N_13877,N_13475,N_12859);
nor U13878 (N_13878,N_13098,N_12055);
nor U13879 (N_13879,N_12156,N_12562);
xor U13880 (N_13880,N_12273,N_13369);
xnor U13881 (N_13881,N_13264,N_13374);
xnor U13882 (N_13882,N_12855,N_12314);
xor U13883 (N_13883,N_12045,N_12631);
nand U13884 (N_13884,N_13336,N_13333);
xor U13885 (N_13885,N_12392,N_13086);
or U13886 (N_13886,N_13479,N_12628);
nor U13887 (N_13887,N_13388,N_12633);
nand U13888 (N_13888,N_12760,N_12845);
or U13889 (N_13889,N_13341,N_12795);
xor U13890 (N_13890,N_13037,N_13236);
nand U13891 (N_13891,N_13157,N_12471);
or U13892 (N_13892,N_12857,N_12240);
nand U13893 (N_13893,N_13446,N_13306);
or U13894 (N_13894,N_12606,N_12554);
nand U13895 (N_13895,N_12356,N_12034);
nand U13896 (N_13896,N_12921,N_12667);
xor U13897 (N_13897,N_12902,N_12383);
and U13898 (N_13898,N_12610,N_13249);
and U13899 (N_13899,N_12048,N_12499);
or U13900 (N_13900,N_13200,N_13397);
xor U13901 (N_13901,N_13392,N_13263);
or U13902 (N_13902,N_12101,N_12705);
xor U13903 (N_13903,N_12721,N_12438);
xor U13904 (N_13904,N_13116,N_13112);
nor U13905 (N_13905,N_12005,N_12098);
or U13906 (N_13906,N_13140,N_13160);
and U13907 (N_13907,N_12698,N_13421);
and U13908 (N_13908,N_12085,N_12952);
nand U13909 (N_13909,N_12643,N_12264);
nand U13910 (N_13910,N_12325,N_12649);
nor U13911 (N_13911,N_12599,N_12789);
or U13912 (N_13912,N_13383,N_13357);
xnor U13913 (N_13913,N_12889,N_13114);
nand U13914 (N_13914,N_13487,N_13251);
xnor U13915 (N_13915,N_12531,N_12223);
nor U13916 (N_13916,N_12441,N_13074);
and U13917 (N_13917,N_12133,N_13175);
or U13918 (N_13918,N_12860,N_12326);
nor U13919 (N_13919,N_12154,N_13040);
xor U13920 (N_13920,N_13314,N_12931);
or U13921 (N_13921,N_12391,N_13042);
or U13922 (N_13922,N_12207,N_13082);
nand U13923 (N_13923,N_12625,N_12832);
and U13924 (N_13924,N_13033,N_13350);
nand U13925 (N_13925,N_13143,N_12293);
and U13926 (N_13926,N_13009,N_13184);
xnor U13927 (N_13927,N_12964,N_12520);
nand U13928 (N_13928,N_12287,N_12148);
xor U13929 (N_13929,N_12213,N_13386);
nand U13930 (N_13930,N_12260,N_12309);
nor U13931 (N_13931,N_13083,N_12961);
and U13932 (N_13932,N_12220,N_13424);
or U13933 (N_13933,N_13025,N_12488);
and U13934 (N_13934,N_13013,N_12301);
nor U13935 (N_13935,N_13000,N_12578);
or U13936 (N_13936,N_12522,N_13295);
nand U13937 (N_13937,N_13183,N_12621);
nand U13938 (N_13938,N_12044,N_12876);
and U13939 (N_13939,N_12078,N_12791);
nand U13940 (N_13940,N_12828,N_12418);
xor U13941 (N_13941,N_13190,N_12225);
and U13942 (N_13942,N_13385,N_13261);
or U13943 (N_13943,N_13187,N_12043);
xnor U13944 (N_13944,N_12940,N_13288);
or U13945 (N_13945,N_12634,N_13492);
nor U13946 (N_13946,N_12304,N_12428);
or U13947 (N_13947,N_13413,N_13485);
xnor U13948 (N_13948,N_13267,N_13244);
nor U13949 (N_13949,N_12737,N_12406);
and U13950 (N_13950,N_12842,N_12505);
xnor U13951 (N_13951,N_13029,N_12873);
nor U13952 (N_13952,N_13017,N_12609);
nand U13953 (N_13953,N_12979,N_12651);
xor U13954 (N_13954,N_13463,N_12468);
xnor U13955 (N_13955,N_13390,N_12117);
nor U13956 (N_13956,N_12595,N_12464);
and U13957 (N_13957,N_12348,N_13121);
nor U13958 (N_13958,N_13276,N_13347);
or U13959 (N_13959,N_12494,N_12936);
xor U13960 (N_13960,N_12074,N_12517);
or U13961 (N_13961,N_12058,N_12039);
or U13962 (N_13962,N_12915,N_13219);
nor U13963 (N_13963,N_13227,N_12960);
and U13964 (N_13964,N_12607,N_12265);
and U13965 (N_13965,N_12059,N_12124);
nor U13966 (N_13966,N_12945,N_12070);
xnor U13967 (N_13967,N_12533,N_13438);
nand U13968 (N_13968,N_12091,N_13447);
or U13969 (N_13969,N_12848,N_12410);
and U13970 (N_13970,N_12027,N_12752);
nor U13971 (N_13971,N_12244,N_13229);
nor U13972 (N_13972,N_12071,N_12024);
nand U13973 (N_13973,N_12613,N_12977);
nor U13974 (N_13974,N_12957,N_13022);
nand U13975 (N_13975,N_13103,N_12458);
nor U13976 (N_13976,N_13332,N_12008);
nand U13977 (N_13977,N_12095,N_12946);
or U13978 (N_13978,N_12510,N_12661);
nor U13979 (N_13979,N_12037,N_12328);
xor U13980 (N_13980,N_13442,N_12703);
or U13981 (N_13981,N_12080,N_12263);
and U13982 (N_13982,N_12226,N_12970);
and U13983 (N_13983,N_12331,N_12267);
xnor U13984 (N_13984,N_12092,N_12696);
xnor U13985 (N_13985,N_12871,N_13222);
or U13986 (N_13986,N_12511,N_12381);
or U13987 (N_13987,N_13470,N_12715);
xnor U13988 (N_13988,N_12812,N_12424);
nor U13989 (N_13989,N_12259,N_13111);
or U13990 (N_13990,N_13254,N_12890);
nor U13991 (N_13991,N_12262,N_12949);
nor U13992 (N_13992,N_13248,N_13297);
and U13993 (N_13993,N_12822,N_13233);
nor U13994 (N_13994,N_13486,N_13425);
nand U13995 (N_13995,N_12805,N_13067);
or U13996 (N_13996,N_12993,N_12216);
nor U13997 (N_13997,N_12540,N_12430);
xnor U13998 (N_13998,N_13177,N_12279);
xnor U13999 (N_13999,N_13172,N_12312);
or U14000 (N_14000,N_13186,N_13118);
or U14001 (N_14001,N_13004,N_13367);
and U14002 (N_14002,N_13070,N_13458);
and U14003 (N_14003,N_13299,N_13480);
and U14004 (N_14004,N_13065,N_12077);
and U14005 (N_14005,N_12193,N_12317);
and U14006 (N_14006,N_12175,N_12145);
and U14007 (N_14007,N_13440,N_12681);
xor U14008 (N_14008,N_12478,N_13145);
nand U14009 (N_14009,N_12204,N_12984);
and U14010 (N_14010,N_12888,N_12587);
nor U14011 (N_14011,N_12772,N_12983);
and U14012 (N_14012,N_12435,N_12753);
xnor U14013 (N_14013,N_13041,N_12409);
nor U14014 (N_14014,N_12316,N_13049);
xor U14015 (N_14015,N_12784,N_12465);
nand U14016 (N_14016,N_12674,N_13481);
nor U14017 (N_14017,N_12407,N_12575);
and U14018 (N_14018,N_12482,N_12258);
nand U14019 (N_14019,N_12073,N_12249);
xnor U14020 (N_14020,N_13434,N_12379);
nor U14021 (N_14021,N_12748,N_12255);
nor U14022 (N_14022,N_13322,N_12166);
nor U14023 (N_14023,N_12169,N_13476);
or U14024 (N_14024,N_12911,N_13265);
nor U14025 (N_14025,N_13460,N_13312);
nand U14026 (N_14026,N_13431,N_12969);
nand U14027 (N_14027,N_12835,N_12780);
xor U14028 (N_14028,N_12551,N_12954);
and U14029 (N_14029,N_13182,N_12125);
nand U14030 (N_14030,N_12841,N_13287);
nor U14031 (N_14031,N_13044,N_13461);
and U14032 (N_14032,N_12572,N_12295);
xor U14033 (N_14033,N_12102,N_12955);
and U14034 (N_14034,N_12470,N_12767);
nor U14035 (N_14035,N_12736,N_12512);
or U14036 (N_14036,N_12597,N_12710);
nand U14037 (N_14037,N_13389,N_13469);
nor U14038 (N_14038,N_13362,N_13345);
xnor U14039 (N_14039,N_12217,N_12974);
xor U14040 (N_14040,N_12766,N_12467);
xor U14041 (N_14041,N_13356,N_12455);
xor U14042 (N_14042,N_12676,N_12895);
xor U14043 (N_14043,N_12688,N_13073);
xor U14044 (N_14044,N_13228,N_13204);
and U14045 (N_14045,N_12668,N_12830);
and U14046 (N_14046,N_12492,N_12879);
and U14047 (N_14047,N_12281,N_13426);
or U14048 (N_14048,N_13498,N_13393);
nor U14049 (N_14049,N_12928,N_13324);
nor U14050 (N_14050,N_12723,N_13123);
nand U14051 (N_14051,N_13198,N_12163);
nand U14052 (N_14052,N_12306,N_12448);
or U14053 (N_14053,N_12177,N_13059);
or U14054 (N_14054,N_13096,N_13474);
nor U14055 (N_14055,N_13491,N_13115);
or U14056 (N_14056,N_13055,N_13141);
or U14057 (N_14057,N_12612,N_13326);
or U14058 (N_14058,N_13408,N_12487);
and U14059 (N_14059,N_12813,N_12611);
nand U14060 (N_14060,N_12313,N_12982);
nor U14061 (N_14061,N_13122,N_12127);
nand U14062 (N_14062,N_13101,N_12210);
nor U14063 (N_14063,N_12485,N_12966);
nor U14064 (N_14064,N_13079,N_12629);
nor U14065 (N_14065,N_12965,N_12669);
nor U14066 (N_14066,N_12684,N_12963);
or U14067 (N_14067,N_13210,N_12655);
and U14068 (N_14068,N_13168,N_12242);
nand U14069 (N_14069,N_12384,N_13146);
nand U14070 (N_14070,N_13056,N_12539);
nor U14071 (N_14071,N_12637,N_13174);
nand U14072 (N_14072,N_13499,N_12523);
nor U14073 (N_14073,N_12311,N_12452);
xnor U14074 (N_14074,N_12743,N_12370);
nand U14075 (N_14075,N_12497,N_12167);
nor U14076 (N_14076,N_12300,N_12276);
xor U14077 (N_14077,N_13247,N_12807);
nor U14078 (N_14078,N_12224,N_12090);
xnor U14079 (N_14079,N_12829,N_12765);
nand U14080 (N_14080,N_13429,N_12378);
and U14081 (N_14081,N_13466,N_12201);
nor U14082 (N_14082,N_12052,N_12486);
nor U14083 (N_14083,N_13088,N_13171);
xor U14084 (N_14084,N_12082,N_12414);
xor U14085 (N_14085,N_12542,N_12268);
or U14086 (N_14086,N_12516,N_12858);
xnor U14087 (N_14087,N_12222,N_12573);
xor U14088 (N_14088,N_12010,N_12639);
or U14089 (N_14089,N_12296,N_12810);
or U14090 (N_14090,N_12865,N_12788);
nor U14091 (N_14091,N_12927,N_13019);
xor U14092 (N_14092,N_13241,N_13124);
or U14093 (N_14093,N_12717,N_12068);
nor U14094 (N_14094,N_12335,N_12120);
or U14095 (N_14095,N_12652,N_12000);
nand U14096 (N_14096,N_12108,N_12803);
nand U14097 (N_14097,N_12605,N_13161);
nand U14098 (N_14098,N_12119,N_12149);
nand U14099 (N_14099,N_12686,N_13396);
xor U14100 (N_14100,N_12544,N_13181);
nand U14101 (N_14101,N_12395,N_12302);
nor U14102 (N_14102,N_12343,N_12601);
or U14103 (N_14103,N_13409,N_13377);
nor U14104 (N_14104,N_12796,N_13398);
nor U14105 (N_14105,N_13335,N_12072);
or U14106 (N_14106,N_12025,N_13099);
nand U14107 (N_14107,N_12837,N_12589);
or U14108 (N_14108,N_12713,N_12536);
or U14109 (N_14109,N_12288,N_12032);
and U14110 (N_14110,N_12347,N_12917);
and U14111 (N_14111,N_12755,N_12769);
or U14112 (N_14112,N_12437,N_12565);
nand U14113 (N_14113,N_13405,N_12113);
nor U14114 (N_14114,N_13027,N_12318);
nand U14115 (N_14115,N_12507,N_13472);
and U14116 (N_14116,N_12183,N_12801);
and U14117 (N_14117,N_12051,N_13318);
nand U14118 (N_14118,N_13205,N_12017);
or U14119 (N_14119,N_13406,N_13209);
xor U14120 (N_14120,N_13047,N_12630);
and U14121 (N_14121,N_13194,N_13339);
xnor U14122 (N_14122,N_13062,N_12344);
nor U14123 (N_14123,N_12962,N_12916);
nand U14124 (N_14124,N_12215,N_13444);
nor U14125 (N_14125,N_12771,N_12446);
and U14126 (N_14126,N_13359,N_12600);
nand U14127 (N_14127,N_12456,N_13214);
or U14128 (N_14128,N_12457,N_12741);
nor U14129 (N_14129,N_12577,N_12653);
xnor U14130 (N_14130,N_13162,N_12863);
and U14131 (N_14131,N_13456,N_12477);
nand U14132 (N_14132,N_12172,N_12372);
or U14133 (N_14133,N_12553,N_13373);
xor U14134 (N_14134,N_12777,N_13188);
nor U14135 (N_14135,N_12744,N_13468);
nand U14136 (N_14136,N_12329,N_12712);
nor U14137 (N_14137,N_12588,N_13376);
or U14138 (N_14138,N_12199,N_12819);
and U14139 (N_14139,N_12590,N_12513);
nor U14140 (N_14140,N_13325,N_12463);
nand U14141 (N_14141,N_12205,N_12619);
xnor U14142 (N_14142,N_13154,N_12718);
nor U14143 (N_14143,N_13266,N_13419);
xnor U14144 (N_14144,N_12942,N_12790);
nand U14145 (N_14145,N_12143,N_13351);
nor U14146 (N_14146,N_12340,N_12733);
and U14147 (N_14147,N_12451,N_12324);
or U14148 (N_14148,N_12827,N_12350);
or U14149 (N_14149,N_13280,N_13089);
or U14150 (N_14150,N_12912,N_12868);
or U14151 (N_14151,N_12543,N_12100);
nand U14152 (N_14152,N_13081,N_12375);
nor U14153 (N_14153,N_13155,N_13307);
or U14154 (N_14154,N_12924,N_12146);
or U14155 (N_14155,N_12415,N_13206);
nand U14156 (N_14156,N_13104,N_12363);
nand U14157 (N_14157,N_13158,N_13260);
nor U14158 (N_14158,N_12528,N_12672);
and U14159 (N_14159,N_12939,N_12496);
or U14160 (N_14160,N_12802,N_12992);
and U14161 (N_14161,N_13153,N_12692);
nand U14162 (N_14162,N_12346,N_12351);
nand U14163 (N_14163,N_12726,N_12833);
xnor U14164 (N_14164,N_12030,N_12011);
xnor U14165 (N_14165,N_12751,N_12956);
nand U14166 (N_14166,N_12251,N_13253);
nand U14167 (N_14167,N_12420,N_13291);
and U14168 (N_14168,N_12069,N_13437);
xnor U14169 (N_14169,N_12015,N_12853);
or U14170 (N_14170,N_12001,N_12160);
nor U14171 (N_14171,N_12475,N_13310);
xnor U14172 (N_14172,N_12278,N_12170);
or U14173 (N_14173,N_12422,N_12693);
or U14174 (N_14174,N_12083,N_12219);
nor U14175 (N_14175,N_12360,N_13271);
xor U14176 (N_14176,N_12134,N_12694);
nand U14177 (N_14177,N_12990,N_12763);
xnor U14178 (N_14178,N_13071,N_12342);
or U14179 (N_14179,N_12097,N_13467);
xor U14180 (N_14180,N_13134,N_12918);
xor U14181 (N_14181,N_12503,N_13034);
nand U14182 (N_14182,N_13321,N_13133);
or U14183 (N_14183,N_12725,N_13353);
and U14184 (N_14184,N_12645,N_12783);
nand U14185 (N_14185,N_12823,N_12593);
or U14186 (N_14186,N_13159,N_12770);
nand U14187 (N_14187,N_12978,N_13450);
nand U14188 (N_14188,N_12500,N_12806);
and U14189 (N_14189,N_12932,N_12275);
xor U14190 (N_14190,N_13407,N_13223);
nor U14191 (N_14191,N_12943,N_13482);
or U14192 (N_14192,N_12320,N_13142);
xnor U14193 (N_14193,N_13031,N_12660);
xor U14194 (N_14194,N_12033,N_12221);
nand U14195 (N_14195,N_13410,N_12734);
nor U14196 (N_14196,N_13452,N_12887);
and U14197 (N_14197,N_12063,N_12550);
or U14198 (N_14198,N_12675,N_12310);
nor U14199 (N_14199,N_13094,N_13005);
nand U14200 (N_14200,N_13323,N_12560);
and U14201 (N_14201,N_12831,N_13170);
xnor U14202 (N_14202,N_12524,N_12779);
nand U14203 (N_14203,N_12794,N_12947);
or U14204 (N_14204,N_13057,N_12498);
and U14205 (N_14205,N_12014,N_12950);
nor U14206 (N_14206,N_12385,N_12269);
xor U14207 (N_14207,N_13365,N_12460);
and U14208 (N_14208,N_13215,N_13274);
nand U14209 (N_14209,N_12591,N_12018);
xor U14210 (N_14210,N_12434,N_13237);
and U14211 (N_14211,N_12196,N_12862);
xnor U14212 (N_14212,N_12137,N_13259);
or U14213 (N_14213,N_12087,N_12369);
and U14214 (N_14214,N_13256,N_12031);
xnor U14215 (N_14215,N_12834,N_12708);
and U14216 (N_14216,N_12635,N_13395);
nand U14217 (N_14217,N_13283,N_12399);
nand U14218 (N_14218,N_12920,N_12719);
and U14219 (N_14219,N_12627,N_13102);
nand U14220 (N_14220,N_12501,N_12878);
or U14221 (N_14221,N_13176,N_12666);
xnor U14222 (N_14222,N_12084,N_13144);
xnor U14223 (N_14223,N_12246,N_13167);
nand U14224 (N_14224,N_13245,N_13269);
nand U14225 (N_14225,N_12123,N_13226);
nor U14226 (N_14226,N_12644,N_12330);
xor U14227 (N_14227,N_12382,N_12136);
or U14228 (N_14228,N_12461,N_12899);
nor U14229 (N_14229,N_12592,N_13043);
and U14230 (N_14230,N_12615,N_12861);
nor U14231 (N_14231,N_12380,N_12731);
or U14232 (N_14232,N_13371,N_13342);
nor U14233 (N_14233,N_12971,N_12423);
nor U14234 (N_14234,N_13399,N_12691);
or U14235 (N_14235,N_13097,N_13320);
xnor U14236 (N_14236,N_13072,N_13285);
nor U14237 (N_14237,N_12197,N_12286);
or U14238 (N_14238,N_12453,N_12864);
nor U14239 (N_14239,N_12994,N_12757);
xor U14240 (N_14240,N_12157,N_13035);
or U14241 (N_14241,N_12816,N_12191);
or U14242 (N_14242,N_13015,N_13391);
xnor U14243 (N_14243,N_13315,N_13257);
or U14244 (N_14244,N_12975,N_12850);
and U14245 (N_14245,N_12690,N_12359);
nor U14246 (N_14246,N_12632,N_12914);
xor U14247 (N_14247,N_12057,N_12241);
nor U14248 (N_14248,N_12662,N_13420);
nand U14249 (N_14249,N_12245,N_12776);
nand U14250 (N_14250,N_12454,N_12244);
or U14251 (N_14251,N_13256,N_12001);
and U14252 (N_14252,N_12311,N_12014);
xnor U14253 (N_14253,N_12431,N_12907);
or U14254 (N_14254,N_12522,N_12426);
xnor U14255 (N_14255,N_13121,N_13313);
nor U14256 (N_14256,N_13438,N_12664);
xnor U14257 (N_14257,N_13147,N_12479);
or U14258 (N_14258,N_12781,N_13454);
nor U14259 (N_14259,N_13239,N_12937);
or U14260 (N_14260,N_13211,N_13281);
and U14261 (N_14261,N_12123,N_12609);
and U14262 (N_14262,N_12809,N_12706);
or U14263 (N_14263,N_13135,N_13351);
and U14264 (N_14264,N_13484,N_13301);
nor U14265 (N_14265,N_12345,N_13280);
xor U14266 (N_14266,N_12385,N_12156);
or U14267 (N_14267,N_12124,N_13240);
nor U14268 (N_14268,N_13250,N_12455);
xor U14269 (N_14269,N_13144,N_13422);
or U14270 (N_14270,N_12037,N_13112);
and U14271 (N_14271,N_13351,N_12638);
and U14272 (N_14272,N_12744,N_12559);
xor U14273 (N_14273,N_13212,N_13088);
and U14274 (N_14274,N_12707,N_12317);
and U14275 (N_14275,N_12686,N_13029);
nor U14276 (N_14276,N_12304,N_12858);
nor U14277 (N_14277,N_12441,N_12898);
nand U14278 (N_14278,N_13187,N_13307);
and U14279 (N_14279,N_12422,N_12466);
nand U14280 (N_14280,N_12106,N_12411);
nand U14281 (N_14281,N_12921,N_12817);
nand U14282 (N_14282,N_12180,N_12277);
or U14283 (N_14283,N_13262,N_13044);
or U14284 (N_14284,N_12710,N_13408);
nand U14285 (N_14285,N_12149,N_13437);
xor U14286 (N_14286,N_13039,N_12071);
and U14287 (N_14287,N_13154,N_13079);
and U14288 (N_14288,N_13050,N_13170);
and U14289 (N_14289,N_12040,N_13466);
nand U14290 (N_14290,N_12352,N_12005);
and U14291 (N_14291,N_13208,N_13236);
nand U14292 (N_14292,N_12117,N_12412);
nand U14293 (N_14293,N_12283,N_13330);
nor U14294 (N_14294,N_13307,N_12355);
and U14295 (N_14295,N_13263,N_12511);
or U14296 (N_14296,N_13190,N_12360);
nand U14297 (N_14297,N_13371,N_12779);
nand U14298 (N_14298,N_12064,N_13051);
xor U14299 (N_14299,N_12721,N_12846);
and U14300 (N_14300,N_12957,N_13131);
nor U14301 (N_14301,N_13436,N_12872);
and U14302 (N_14302,N_12995,N_12852);
and U14303 (N_14303,N_13337,N_13325);
or U14304 (N_14304,N_12919,N_12994);
nand U14305 (N_14305,N_13288,N_13009);
nor U14306 (N_14306,N_12135,N_13250);
nor U14307 (N_14307,N_13280,N_13105);
nand U14308 (N_14308,N_12279,N_12442);
nand U14309 (N_14309,N_12840,N_12336);
or U14310 (N_14310,N_12192,N_12967);
and U14311 (N_14311,N_12185,N_13082);
nor U14312 (N_14312,N_12769,N_13220);
nand U14313 (N_14313,N_13090,N_13117);
and U14314 (N_14314,N_12910,N_12815);
and U14315 (N_14315,N_12833,N_12779);
nor U14316 (N_14316,N_13076,N_12840);
xnor U14317 (N_14317,N_12834,N_12999);
nor U14318 (N_14318,N_12287,N_12953);
or U14319 (N_14319,N_12499,N_13179);
xnor U14320 (N_14320,N_13126,N_12031);
xor U14321 (N_14321,N_12007,N_12116);
nor U14322 (N_14322,N_12836,N_13056);
nor U14323 (N_14323,N_13127,N_13300);
or U14324 (N_14324,N_12782,N_12463);
nor U14325 (N_14325,N_13338,N_12674);
nor U14326 (N_14326,N_12673,N_12070);
or U14327 (N_14327,N_12296,N_12511);
or U14328 (N_14328,N_12390,N_12964);
nand U14329 (N_14329,N_13080,N_12220);
xor U14330 (N_14330,N_12175,N_12877);
or U14331 (N_14331,N_12594,N_13303);
nor U14332 (N_14332,N_12347,N_12859);
and U14333 (N_14333,N_12044,N_13361);
xor U14334 (N_14334,N_13281,N_12272);
or U14335 (N_14335,N_13402,N_12860);
and U14336 (N_14336,N_12890,N_12457);
and U14337 (N_14337,N_12454,N_13346);
nor U14338 (N_14338,N_12842,N_12015);
or U14339 (N_14339,N_13186,N_12582);
and U14340 (N_14340,N_13008,N_12381);
xor U14341 (N_14341,N_13405,N_13138);
or U14342 (N_14342,N_13021,N_13461);
and U14343 (N_14343,N_13339,N_12652);
or U14344 (N_14344,N_13302,N_13122);
nor U14345 (N_14345,N_12103,N_12288);
nand U14346 (N_14346,N_12924,N_12226);
nand U14347 (N_14347,N_12669,N_12981);
nor U14348 (N_14348,N_13402,N_12816);
nor U14349 (N_14349,N_12838,N_13082);
or U14350 (N_14350,N_13192,N_12076);
or U14351 (N_14351,N_12087,N_12709);
xor U14352 (N_14352,N_12460,N_13275);
nor U14353 (N_14353,N_12948,N_13154);
nor U14354 (N_14354,N_13081,N_12477);
and U14355 (N_14355,N_13047,N_12424);
nor U14356 (N_14356,N_12541,N_13324);
xor U14357 (N_14357,N_12763,N_12436);
nor U14358 (N_14358,N_13223,N_12214);
and U14359 (N_14359,N_12600,N_13192);
or U14360 (N_14360,N_12297,N_12597);
nor U14361 (N_14361,N_13160,N_12425);
nand U14362 (N_14362,N_12690,N_12074);
nand U14363 (N_14363,N_12905,N_12384);
and U14364 (N_14364,N_13445,N_13181);
and U14365 (N_14365,N_12227,N_12261);
and U14366 (N_14366,N_12929,N_12556);
nor U14367 (N_14367,N_13226,N_12494);
nor U14368 (N_14368,N_12784,N_12386);
or U14369 (N_14369,N_12814,N_13419);
nand U14370 (N_14370,N_12397,N_13494);
nor U14371 (N_14371,N_13175,N_12169);
xor U14372 (N_14372,N_13263,N_12099);
nor U14373 (N_14373,N_13445,N_12321);
and U14374 (N_14374,N_12729,N_12588);
or U14375 (N_14375,N_13087,N_13043);
or U14376 (N_14376,N_13125,N_13077);
nor U14377 (N_14377,N_13467,N_13157);
and U14378 (N_14378,N_13346,N_12542);
nand U14379 (N_14379,N_12389,N_12419);
nor U14380 (N_14380,N_13444,N_12521);
and U14381 (N_14381,N_13484,N_12649);
xor U14382 (N_14382,N_13282,N_12509);
and U14383 (N_14383,N_12605,N_12059);
xnor U14384 (N_14384,N_13205,N_12927);
nand U14385 (N_14385,N_12146,N_12994);
or U14386 (N_14386,N_12640,N_12367);
xor U14387 (N_14387,N_13316,N_12842);
nor U14388 (N_14388,N_13422,N_12092);
nand U14389 (N_14389,N_12965,N_13132);
nand U14390 (N_14390,N_13336,N_12520);
nand U14391 (N_14391,N_13462,N_12073);
or U14392 (N_14392,N_13217,N_12980);
nand U14393 (N_14393,N_12791,N_12394);
xnor U14394 (N_14394,N_12283,N_12942);
nor U14395 (N_14395,N_13102,N_13068);
or U14396 (N_14396,N_12428,N_12900);
and U14397 (N_14397,N_13432,N_12017);
nor U14398 (N_14398,N_12091,N_12459);
xor U14399 (N_14399,N_13195,N_12935);
nor U14400 (N_14400,N_13267,N_12927);
xnor U14401 (N_14401,N_12717,N_12332);
nand U14402 (N_14402,N_12874,N_12213);
nand U14403 (N_14403,N_12171,N_12505);
nand U14404 (N_14404,N_13085,N_12799);
or U14405 (N_14405,N_13170,N_12239);
nor U14406 (N_14406,N_13153,N_12547);
nand U14407 (N_14407,N_12315,N_12170);
nand U14408 (N_14408,N_12439,N_13108);
or U14409 (N_14409,N_12312,N_12789);
nor U14410 (N_14410,N_13054,N_12240);
xor U14411 (N_14411,N_13114,N_12807);
and U14412 (N_14412,N_12433,N_12542);
nand U14413 (N_14413,N_12211,N_12019);
and U14414 (N_14414,N_13426,N_12597);
or U14415 (N_14415,N_12623,N_12177);
or U14416 (N_14416,N_12604,N_12129);
nor U14417 (N_14417,N_12197,N_12443);
and U14418 (N_14418,N_12855,N_12884);
nor U14419 (N_14419,N_12104,N_12174);
xor U14420 (N_14420,N_13466,N_12432);
and U14421 (N_14421,N_12530,N_13026);
xor U14422 (N_14422,N_12583,N_13306);
nor U14423 (N_14423,N_12634,N_13119);
and U14424 (N_14424,N_13235,N_12318);
nand U14425 (N_14425,N_13471,N_13217);
or U14426 (N_14426,N_12861,N_13110);
or U14427 (N_14427,N_12140,N_12298);
nor U14428 (N_14428,N_13087,N_12628);
nor U14429 (N_14429,N_12020,N_12119);
and U14430 (N_14430,N_12392,N_12530);
or U14431 (N_14431,N_12627,N_12623);
nand U14432 (N_14432,N_12417,N_12105);
and U14433 (N_14433,N_12465,N_12540);
nor U14434 (N_14434,N_12403,N_12031);
xnor U14435 (N_14435,N_13219,N_12457);
nor U14436 (N_14436,N_13236,N_13437);
nor U14437 (N_14437,N_12861,N_12262);
nand U14438 (N_14438,N_12900,N_12097);
or U14439 (N_14439,N_12547,N_12907);
nand U14440 (N_14440,N_13368,N_13130);
nand U14441 (N_14441,N_12278,N_12123);
nand U14442 (N_14442,N_12226,N_12555);
nand U14443 (N_14443,N_12370,N_12626);
and U14444 (N_14444,N_12382,N_12145);
nor U14445 (N_14445,N_12053,N_12141);
xor U14446 (N_14446,N_12117,N_13366);
or U14447 (N_14447,N_12155,N_12773);
or U14448 (N_14448,N_12355,N_13461);
nor U14449 (N_14449,N_12493,N_12501);
and U14450 (N_14450,N_12525,N_13305);
and U14451 (N_14451,N_13181,N_12744);
and U14452 (N_14452,N_12825,N_12664);
xnor U14453 (N_14453,N_13045,N_12736);
and U14454 (N_14454,N_12460,N_13247);
nor U14455 (N_14455,N_12328,N_12056);
xor U14456 (N_14456,N_12427,N_12479);
xor U14457 (N_14457,N_12798,N_13114);
nand U14458 (N_14458,N_12214,N_12852);
and U14459 (N_14459,N_12002,N_13402);
or U14460 (N_14460,N_12929,N_12908);
nand U14461 (N_14461,N_12236,N_12147);
nor U14462 (N_14462,N_13260,N_13062);
or U14463 (N_14463,N_12709,N_12751);
xor U14464 (N_14464,N_12791,N_12084);
nand U14465 (N_14465,N_12781,N_13225);
or U14466 (N_14466,N_12554,N_13351);
and U14467 (N_14467,N_12285,N_13027);
nand U14468 (N_14468,N_13413,N_12048);
nor U14469 (N_14469,N_12724,N_12039);
nor U14470 (N_14470,N_12024,N_13136);
and U14471 (N_14471,N_12951,N_12118);
and U14472 (N_14472,N_12836,N_12100);
nor U14473 (N_14473,N_12531,N_12346);
nand U14474 (N_14474,N_13224,N_13480);
xnor U14475 (N_14475,N_12477,N_13045);
xor U14476 (N_14476,N_12438,N_13209);
xor U14477 (N_14477,N_13255,N_13484);
nor U14478 (N_14478,N_12673,N_12957);
or U14479 (N_14479,N_12619,N_13136);
xor U14480 (N_14480,N_13395,N_12650);
and U14481 (N_14481,N_12227,N_12032);
and U14482 (N_14482,N_12189,N_13374);
and U14483 (N_14483,N_12746,N_13264);
or U14484 (N_14484,N_13470,N_12745);
or U14485 (N_14485,N_13195,N_12088);
nand U14486 (N_14486,N_12119,N_13398);
nand U14487 (N_14487,N_12959,N_12127);
xnor U14488 (N_14488,N_12448,N_13482);
and U14489 (N_14489,N_12388,N_12872);
nand U14490 (N_14490,N_13342,N_13176);
nor U14491 (N_14491,N_12889,N_12911);
nand U14492 (N_14492,N_12645,N_12376);
nor U14493 (N_14493,N_12839,N_12024);
nor U14494 (N_14494,N_13074,N_12485);
xor U14495 (N_14495,N_13437,N_12322);
nand U14496 (N_14496,N_12019,N_13431);
xor U14497 (N_14497,N_13417,N_13349);
nand U14498 (N_14498,N_12819,N_12414);
xor U14499 (N_14499,N_13192,N_12041);
xor U14500 (N_14500,N_12379,N_13465);
and U14501 (N_14501,N_13122,N_12984);
or U14502 (N_14502,N_13225,N_13113);
or U14503 (N_14503,N_12165,N_12643);
nand U14504 (N_14504,N_12549,N_12722);
nor U14505 (N_14505,N_12136,N_12752);
xor U14506 (N_14506,N_12485,N_13273);
nor U14507 (N_14507,N_13110,N_12974);
xor U14508 (N_14508,N_12615,N_13376);
and U14509 (N_14509,N_13455,N_12760);
or U14510 (N_14510,N_12369,N_13278);
xnor U14511 (N_14511,N_12542,N_13102);
nand U14512 (N_14512,N_12928,N_12661);
nand U14513 (N_14513,N_13052,N_13005);
nand U14514 (N_14514,N_13309,N_12338);
nor U14515 (N_14515,N_12786,N_12901);
and U14516 (N_14516,N_12999,N_12600);
nor U14517 (N_14517,N_13465,N_12419);
and U14518 (N_14518,N_12519,N_13197);
xnor U14519 (N_14519,N_13292,N_12997);
and U14520 (N_14520,N_12698,N_12840);
xor U14521 (N_14521,N_13478,N_13180);
xnor U14522 (N_14522,N_12862,N_13202);
nor U14523 (N_14523,N_12867,N_12105);
nor U14524 (N_14524,N_12319,N_12203);
and U14525 (N_14525,N_13294,N_12983);
nand U14526 (N_14526,N_12246,N_12702);
xnor U14527 (N_14527,N_12335,N_12836);
nand U14528 (N_14528,N_13044,N_12113);
or U14529 (N_14529,N_12375,N_13423);
xor U14530 (N_14530,N_12371,N_12055);
xnor U14531 (N_14531,N_12032,N_13449);
nor U14532 (N_14532,N_12559,N_12927);
nor U14533 (N_14533,N_13472,N_12925);
nand U14534 (N_14534,N_12907,N_13132);
nor U14535 (N_14535,N_13093,N_13218);
and U14536 (N_14536,N_13140,N_12153);
and U14537 (N_14537,N_12716,N_12636);
nor U14538 (N_14538,N_12452,N_13428);
nor U14539 (N_14539,N_12413,N_13278);
or U14540 (N_14540,N_13327,N_13193);
nor U14541 (N_14541,N_12869,N_12550);
and U14542 (N_14542,N_12479,N_13270);
or U14543 (N_14543,N_13320,N_13173);
or U14544 (N_14544,N_13150,N_12400);
xor U14545 (N_14545,N_12677,N_12589);
nor U14546 (N_14546,N_12662,N_13493);
and U14547 (N_14547,N_12166,N_13020);
or U14548 (N_14548,N_13072,N_12833);
nor U14549 (N_14549,N_13449,N_12209);
xor U14550 (N_14550,N_12178,N_12927);
and U14551 (N_14551,N_12338,N_12289);
nand U14552 (N_14552,N_12118,N_12545);
xnor U14553 (N_14553,N_12093,N_12252);
or U14554 (N_14554,N_13232,N_13420);
xor U14555 (N_14555,N_13068,N_12640);
nand U14556 (N_14556,N_12270,N_12451);
nand U14557 (N_14557,N_13201,N_12900);
xor U14558 (N_14558,N_12294,N_13478);
xor U14559 (N_14559,N_13163,N_12091);
and U14560 (N_14560,N_12055,N_13196);
or U14561 (N_14561,N_12867,N_13073);
nand U14562 (N_14562,N_13160,N_12496);
and U14563 (N_14563,N_12536,N_12542);
nor U14564 (N_14564,N_12158,N_13144);
xnor U14565 (N_14565,N_12065,N_13184);
nor U14566 (N_14566,N_13091,N_12596);
or U14567 (N_14567,N_12064,N_12156);
and U14568 (N_14568,N_12208,N_13079);
nand U14569 (N_14569,N_13024,N_13116);
or U14570 (N_14570,N_12936,N_12298);
nand U14571 (N_14571,N_13396,N_12042);
nor U14572 (N_14572,N_13402,N_12967);
nand U14573 (N_14573,N_13122,N_13379);
nor U14574 (N_14574,N_13450,N_13294);
nand U14575 (N_14575,N_12542,N_12648);
or U14576 (N_14576,N_12369,N_12470);
or U14577 (N_14577,N_12908,N_12024);
nor U14578 (N_14578,N_13253,N_12233);
nor U14579 (N_14579,N_12405,N_12717);
and U14580 (N_14580,N_13330,N_12602);
or U14581 (N_14581,N_12618,N_12201);
nor U14582 (N_14582,N_12947,N_12172);
nand U14583 (N_14583,N_12158,N_12055);
or U14584 (N_14584,N_13429,N_13279);
or U14585 (N_14585,N_12000,N_13285);
xor U14586 (N_14586,N_12454,N_12236);
nor U14587 (N_14587,N_12199,N_12232);
nand U14588 (N_14588,N_12917,N_12406);
or U14589 (N_14589,N_13177,N_12282);
and U14590 (N_14590,N_12312,N_13325);
nor U14591 (N_14591,N_13401,N_12494);
nand U14592 (N_14592,N_12110,N_12527);
and U14593 (N_14593,N_13160,N_12819);
xor U14594 (N_14594,N_12938,N_13460);
nand U14595 (N_14595,N_13300,N_12221);
nor U14596 (N_14596,N_13110,N_12079);
nor U14597 (N_14597,N_12266,N_12808);
xnor U14598 (N_14598,N_13293,N_12091);
and U14599 (N_14599,N_13073,N_12236);
xor U14600 (N_14600,N_13119,N_12985);
and U14601 (N_14601,N_12627,N_12816);
nor U14602 (N_14602,N_12638,N_13261);
nor U14603 (N_14603,N_12022,N_12413);
or U14604 (N_14604,N_13401,N_12222);
nand U14605 (N_14605,N_13472,N_12115);
and U14606 (N_14606,N_13257,N_12290);
and U14607 (N_14607,N_12838,N_13441);
and U14608 (N_14608,N_12695,N_12141);
nor U14609 (N_14609,N_12904,N_12724);
nor U14610 (N_14610,N_13203,N_13365);
and U14611 (N_14611,N_13491,N_12513);
xor U14612 (N_14612,N_13296,N_12347);
xor U14613 (N_14613,N_12606,N_12803);
or U14614 (N_14614,N_12656,N_12815);
or U14615 (N_14615,N_12639,N_13267);
xor U14616 (N_14616,N_13284,N_12532);
xor U14617 (N_14617,N_13156,N_13142);
and U14618 (N_14618,N_12769,N_12275);
and U14619 (N_14619,N_12857,N_13246);
xnor U14620 (N_14620,N_12133,N_12342);
and U14621 (N_14621,N_12100,N_13137);
or U14622 (N_14622,N_13115,N_12637);
xnor U14623 (N_14623,N_13178,N_13163);
and U14624 (N_14624,N_12596,N_12531);
nand U14625 (N_14625,N_12152,N_12033);
xor U14626 (N_14626,N_13429,N_12769);
nand U14627 (N_14627,N_13425,N_12518);
or U14628 (N_14628,N_12436,N_12080);
nand U14629 (N_14629,N_12439,N_12985);
nor U14630 (N_14630,N_12178,N_13345);
nor U14631 (N_14631,N_12821,N_13145);
xnor U14632 (N_14632,N_13165,N_13340);
and U14633 (N_14633,N_12331,N_13306);
nand U14634 (N_14634,N_12229,N_13123);
nor U14635 (N_14635,N_12764,N_12077);
xor U14636 (N_14636,N_12077,N_13321);
nor U14637 (N_14637,N_12783,N_12658);
nor U14638 (N_14638,N_13002,N_12835);
xnor U14639 (N_14639,N_12854,N_12466);
xnor U14640 (N_14640,N_12875,N_13348);
xnor U14641 (N_14641,N_12955,N_13333);
nor U14642 (N_14642,N_13496,N_13089);
nor U14643 (N_14643,N_13363,N_13157);
nor U14644 (N_14644,N_13426,N_12908);
nor U14645 (N_14645,N_12650,N_12147);
nor U14646 (N_14646,N_12285,N_12892);
and U14647 (N_14647,N_12792,N_13309);
xnor U14648 (N_14648,N_13212,N_12608);
and U14649 (N_14649,N_12417,N_12894);
and U14650 (N_14650,N_12071,N_13149);
or U14651 (N_14651,N_12260,N_12474);
or U14652 (N_14652,N_12790,N_12823);
xor U14653 (N_14653,N_12697,N_13418);
or U14654 (N_14654,N_12344,N_12438);
and U14655 (N_14655,N_13260,N_12493);
and U14656 (N_14656,N_12867,N_12879);
nand U14657 (N_14657,N_12068,N_12490);
nand U14658 (N_14658,N_12510,N_12232);
and U14659 (N_14659,N_12340,N_13185);
nor U14660 (N_14660,N_12351,N_13080);
and U14661 (N_14661,N_12770,N_13241);
xnor U14662 (N_14662,N_12308,N_12205);
and U14663 (N_14663,N_12150,N_13351);
nor U14664 (N_14664,N_12040,N_12948);
and U14665 (N_14665,N_12210,N_12001);
nand U14666 (N_14666,N_12684,N_12331);
and U14667 (N_14667,N_12617,N_12050);
nor U14668 (N_14668,N_12224,N_12134);
and U14669 (N_14669,N_13270,N_12333);
nor U14670 (N_14670,N_12237,N_13069);
and U14671 (N_14671,N_13083,N_12746);
nor U14672 (N_14672,N_13373,N_13030);
or U14673 (N_14673,N_12860,N_12992);
or U14674 (N_14674,N_12876,N_12175);
or U14675 (N_14675,N_12137,N_12835);
xnor U14676 (N_14676,N_12209,N_12576);
xnor U14677 (N_14677,N_12520,N_13140);
nand U14678 (N_14678,N_12894,N_13097);
or U14679 (N_14679,N_12151,N_13452);
xor U14680 (N_14680,N_13208,N_12588);
or U14681 (N_14681,N_13170,N_12001);
and U14682 (N_14682,N_13353,N_12727);
nand U14683 (N_14683,N_12752,N_13093);
and U14684 (N_14684,N_13008,N_12675);
nand U14685 (N_14685,N_12217,N_12146);
or U14686 (N_14686,N_13050,N_13132);
xnor U14687 (N_14687,N_12328,N_12906);
xor U14688 (N_14688,N_12208,N_12919);
and U14689 (N_14689,N_13315,N_13163);
xor U14690 (N_14690,N_12737,N_13012);
and U14691 (N_14691,N_12168,N_13023);
or U14692 (N_14692,N_13201,N_13124);
nand U14693 (N_14693,N_12092,N_12733);
xnor U14694 (N_14694,N_12527,N_12832);
and U14695 (N_14695,N_12940,N_13058);
nor U14696 (N_14696,N_12079,N_13014);
or U14697 (N_14697,N_12154,N_12287);
or U14698 (N_14698,N_12803,N_12556);
xor U14699 (N_14699,N_13081,N_12165);
nand U14700 (N_14700,N_12131,N_12299);
nor U14701 (N_14701,N_13204,N_12401);
nor U14702 (N_14702,N_13414,N_12751);
and U14703 (N_14703,N_13118,N_12827);
and U14704 (N_14704,N_12140,N_13385);
and U14705 (N_14705,N_12792,N_12314);
nand U14706 (N_14706,N_12006,N_13307);
and U14707 (N_14707,N_12944,N_12948);
nand U14708 (N_14708,N_12071,N_12994);
xor U14709 (N_14709,N_13370,N_12739);
nor U14710 (N_14710,N_13146,N_12577);
or U14711 (N_14711,N_13195,N_12423);
or U14712 (N_14712,N_12113,N_13286);
or U14713 (N_14713,N_12810,N_12767);
nand U14714 (N_14714,N_12824,N_13439);
nand U14715 (N_14715,N_13170,N_13084);
nand U14716 (N_14716,N_12120,N_13057);
nand U14717 (N_14717,N_12367,N_12970);
and U14718 (N_14718,N_12351,N_12281);
nor U14719 (N_14719,N_13382,N_12547);
and U14720 (N_14720,N_12947,N_12017);
nor U14721 (N_14721,N_12609,N_12867);
and U14722 (N_14722,N_12576,N_12191);
or U14723 (N_14723,N_12368,N_13462);
nor U14724 (N_14724,N_12359,N_12283);
xor U14725 (N_14725,N_12422,N_12171);
nor U14726 (N_14726,N_12459,N_12632);
or U14727 (N_14727,N_13051,N_13251);
nor U14728 (N_14728,N_12828,N_12671);
and U14729 (N_14729,N_12517,N_12743);
xor U14730 (N_14730,N_12970,N_13076);
nor U14731 (N_14731,N_13143,N_13334);
and U14732 (N_14732,N_12956,N_13066);
nor U14733 (N_14733,N_13382,N_12255);
or U14734 (N_14734,N_12923,N_12509);
nor U14735 (N_14735,N_12275,N_13293);
nand U14736 (N_14736,N_12981,N_12434);
or U14737 (N_14737,N_12951,N_12342);
nor U14738 (N_14738,N_12207,N_12620);
or U14739 (N_14739,N_12837,N_13305);
nor U14740 (N_14740,N_12806,N_12761);
xnor U14741 (N_14741,N_12470,N_12885);
and U14742 (N_14742,N_12838,N_12362);
xnor U14743 (N_14743,N_12079,N_13138);
nor U14744 (N_14744,N_12710,N_13411);
xor U14745 (N_14745,N_13351,N_13227);
and U14746 (N_14746,N_12162,N_12339);
nor U14747 (N_14747,N_12204,N_13203);
xor U14748 (N_14748,N_12943,N_13270);
nor U14749 (N_14749,N_13091,N_12273);
or U14750 (N_14750,N_12318,N_13457);
nand U14751 (N_14751,N_12599,N_12214);
xor U14752 (N_14752,N_12816,N_12337);
nor U14753 (N_14753,N_12127,N_12331);
nand U14754 (N_14754,N_12888,N_13168);
and U14755 (N_14755,N_12793,N_13405);
nor U14756 (N_14756,N_12799,N_12229);
nor U14757 (N_14757,N_12934,N_12264);
nand U14758 (N_14758,N_13082,N_12829);
nand U14759 (N_14759,N_12055,N_13366);
or U14760 (N_14760,N_12378,N_13289);
nand U14761 (N_14761,N_12714,N_12164);
nor U14762 (N_14762,N_12320,N_12675);
nor U14763 (N_14763,N_12689,N_12732);
nor U14764 (N_14764,N_12906,N_13082);
nand U14765 (N_14765,N_13006,N_12460);
and U14766 (N_14766,N_12907,N_12504);
xnor U14767 (N_14767,N_12724,N_13194);
or U14768 (N_14768,N_12166,N_13202);
xnor U14769 (N_14769,N_12813,N_12658);
or U14770 (N_14770,N_13153,N_12841);
xor U14771 (N_14771,N_12896,N_12503);
or U14772 (N_14772,N_12156,N_13182);
and U14773 (N_14773,N_12608,N_13179);
xor U14774 (N_14774,N_12083,N_12574);
nand U14775 (N_14775,N_12897,N_13409);
nor U14776 (N_14776,N_12042,N_12736);
and U14777 (N_14777,N_13329,N_12282);
xnor U14778 (N_14778,N_12952,N_13150);
nand U14779 (N_14779,N_13426,N_12526);
xnor U14780 (N_14780,N_12324,N_12681);
or U14781 (N_14781,N_12965,N_13161);
or U14782 (N_14782,N_12787,N_12530);
or U14783 (N_14783,N_12939,N_12381);
xor U14784 (N_14784,N_12549,N_12602);
nand U14785 (N_14785,N_12413,N_13280);
or U14786 (N_14786,N_12761,N_12721);
and U14787 (N_14787,N_12605,N_12068);
xor U14788 (N_14788,N_12760,N_12952);
nand U14789 (N_14789,N_13313,N_12852);
and U14790 (N_14790,N_12618,N_12156);
nand U14791 (N_14791,N_12286,N_13163);
and U14792 (N_14792,N_12999,N_12489);
or U14793 (N_14793,N_12019,N_12941);
nand U14794 (N_14794,N_12919,N_12002);
xor U14795 (N_14795,N_13448,N_13205);
xor U14796 (N_14796,N_13257,N_13176);
or U14797 (N_14797,N_12381,N_12407);
and U14798 (N_14798,N_13020,N_12417);
and U14799 (N_14799,N_12704,N_12140);
or U14800 (N_14800,N_13272,N_12771);
nor U14801 (N_14801,N_12255,N_12651);
xor U14802 (N_14802,N_12253,N_13069);
nand U14803 (N_14803,N_12086,N_13289);
xor U14804 (N_14804,N_13380,N_12416);
xor U14805 (N_14805,N_12394,N_12995);
nand U14806 (N_14806,N_12380,N_13198);
or U14807 (N_14807,N_12359,N_12706);
nand U14808 (N_14808,N_12574,N_12924);
nand U14809 (N_14809,N_13278,N_12160);
and U14810 (N_14810,N_13162,N_13150);
and U14811 (N_14811,N_12957,N_12642);
or U14812 (N_14812,N_12992,N_13285);
and U14813 (N_14813,N_12720,N_12442);
and U14814 (N_14814,N_12928,N_13025);
nor U14815 (N_14815,N_13127,N_12242);
nor U14816 (N_14816,N_12737,N_12166);
or U14817 (N_14817,N_12585,N_12762);
or U14818 (N_14818,N_12145,N_12722);
or U14819 (N_14819,N_12183,N_12173);
nand U14820 (N_14820,N_12419,N_13310);
nand U14821 (N_14821,N_13383,N_12256);
xnor U14822 (N_14822,N_13197,N_12378);
and U14823 (N_14823,N_12028,N_12138);
xor U14824 (N_14824,N_13132,N_12784);
or U14825 (N_14825,N_12539,N_13434);
nand U14826 (N_14826,N_13226,N_12612);
xnor U14827 (N_14827,N_13216,N_12151);
nand U14828 (N_14828,N_12042,N_13246);
and U14829 (N_14829,N_12647,N_13318);
or U14830 (N_14830,N_12336,N_12080);
nor U14831 (N_14831,N_12953,N_12941);
xor U14832 (N_14832,N_12748,N_12449);
nor U14833 (N_14833,N_12322,N_13045);
and U14834 (N_14834,N_12674,N_12502);
and U14835 (N_14835,N_12809,N_12986);
nor U14836 (N_14836,N_12336,N_13096);
nor U14837 (N_14837,N_12036,N_12765);
xnor U14838 (N_14838,N_12749,N_12829);
nand U14839 (N_14839,N_12918,N_12034);
or U14840 (N_14840,N_12313,N_12262);
nor U14841 (N_14841,N_12319,N_12250);
or U14842 (N_14842,N_12963,N_13074);
nand U14843 (N_14843,N_13126,N_13342);
nand U14844 (N_14844,N_13207,N_13220);
nand U14845 (N_14845,N_12032,N_12546);
nand U14846 (N_14846,N_13080,N_12505);
xnor U14847 (N_14847,N_13291,N_12342);
nand U14848 (N_14848,N_12668,N_13125);
xnor U14849 (N_14849,N_12291,N_12177);
and U14850 (N_14850,N_12244,N_12369);
or U14851 (N_14851,N_13231,N_12998);
or U14852 (N_14852,N_12729,N_12792);
xor U14853 (N_14853,N_12602,N_12585);
and U14854 (N_14854,N_12210,N_12616);
nand U14855 (N_14855,N_13283,N_13317);
nand U14856 (N_14856,N_13052,N_12522);
nor U14857 (N_14857,N_13447,N_12667);
nor U14858 (N_14858,N_13199,N_12652);
and U14859 (N_14859,N_12251,N_13190);
and U14860 (N_14860,N_12006,N_12995);
xnor U14861 (N_14861,N_12962,N_13446);
or U14862 (N_14862,N_13151,N_12966);
and U14863 (N_14863,N_12007,N_12420);
and U14864 (N_14864,N_12266,N_12101);
nand U14865 (N_14865,N_12955,N_12033);
nand U14866 (N_14866,N_12844,N_12974);
xor U14867 (N_14867,N_12817,N_13102);
nand U14868 (N_14868,N_12367,N_12807);
nand U14869 (N_14869,N_12417,N_12151);
nor U14870 (N_14870,N_13023,N_12691);
and U14871 (N_14871,N_12542,N_13403);
nor U14872 (N_14872,N_12184,N_12582);
or U14873 (N_14873,N_13049,N_12643);
nand U14874 (N_14874,N_12553,N_13129);
nor U14875 (N_14875,N_12851,N_13047);
and U14876 (N_14876,N_12014,N_12484);
and U14877 (N_14877,N_12140,N_12084);
xnor U14878 (N_14878,N_12546,N_12473);
or U14879 (N_14879,N_12962,N_12842);
nand U14880 (N_14880,N_12092,N_12511);
xnor U14881 (N_14881,N_12372,N_13259);
or U14882 (N_14882,N_12536,N_12221);
nand U14883 (N_14883,N_12940,N_12299);
nor U14884 (N_14884,N_12605,N_12333);
and U14885 (N_14885,N_12349,N_12304);
nand U14886 (N_14886,N_12613,N_13094);
nor U14887 (N_14887,N_13414,N_12167);
and U14888 (N_14888,N_13023,N_12139);
nand U14889 (N_14889,N_13150,N_12104);
nand U14890 (N_14890,N_13181,N_12382);
and U14891 (N_14891,N_13047,N_12061);
xor U14892 (N_14892,N_13456,N_12168);
or U14893 (N_14893,N_12841,N_12731);
nor U14894 (N_14894,N_13091,N_12526);
and U14895 (N_14895,N_12404,N_12812);
nand U14896 (N_14896,N_12958,N_12659);
nand U14897 (N_14897,N_13246,N_12091);
xor U14898 (N_14898,N_12611,N_13268);
and U14899 (N_14899,N_12389,N_12002);
nor U14900 (N_14900,N_12223,N_13434);
xnor U14901 (N_14901,N_13323,N_12023);
xor U14902 (N_14902,N_12613,N_12609);
and U14903 (N_14903,N_13196,N_12897);
xor U14904 (N_14904,N_13242,N_12497);
xor U14905 (N_14905,N_12702,N_12262);
and U14906 (N_14906,N_12880,N_12196);
and U14907 (N_14907,N_12835,N_12206);
and U14908 (N_14908,N_12008,N_12254);
nor U14909 (N_14909,N_13416,N_12252);
and U14910 (N_14910,N_12702,N_13278);
xnor U14911 (N_14911,N_12907,N_12730);
xnor U14912 (N_14912,N_12273,N_13034);
xor U14913 (N_14913,N_13296,N_13392);
nor U14914 (N_14914,N_12168,N_12633);
nand U14915 (N_14915,N_13352,N_13001);
and U14916 (N_14916,N_12970,N_12022);
xor U14917 (N_14917,N_12365,N_12629);
and U14918 (N_14918,N_12799,N_13375);
nor U14919 (N_14919,N_13185,N_12997);
or U14920 (N_14920,N_13005,N_13400);
nand U14921 (N_14921,N_12229,N_12078);
nand U14922 (N_14922,N_12271,N_13202);
xor U14923 (N_14923,N_13117,N_12168);
xor U14924 (N_14924,N_12081,N_13286);
xnor U14925 (N_14925,N_12790,N_12143);
nor U14926 (N_14926,N_12185,N_12584);
xnor U14927 (N_14927,N_12947,N_12224);
nor U14928 (N_14928,N_12133,N_12385);
xor U14929 (N_14929,N_13397,N_13039);
or U14930 (N_14930,N_12167,N_13162);
or U14931 (N_14931,N_12422,N_12138);
or U14932 (N_14932,N_13417,N_12929);
xor U14933 (N_14933,N_13169,N_12705);
xnor U14934 (N_14934,N_12942,N_12688);
nand U14935 (N_14935,N_12869,N_12461);
or U14936 (N_14936,N_12338,N_12605);
nand U14937 (N_14937,N_13192,N_12218);
and U14938 (N_14938,N_12131,N_13341);
nand U14939 (N_14939,N_13460,N_13472);
or U14940 (N_14940,N_12693,N_12307);
and U14941 (N_14941,N_12663,N_12889);
xnor U14942 (N_14942,N_12196,N_12542);
and U14943 (N_14943,N_12386,N_12198);
nand U14944 (N_14944,N_12516,N_12998);
xnor U14945 (N_14945,N_12957,N_12634);
and U14946 (N_14946,N_12716,N_13090);
nand U14947 (N_14947,N_12915,N_12929);
nor U14948 (N_14948,N_13472,N_12378);
and U14949 (N_14949,N_12242,N_12623);
and U14950 (N_14950,N_12727,N_12950);
and U14951 (N_14951,N_13011,N_13053);
xor U14952 (N_14952,N_12920,N_12598);
and U14953 (N_14953,N_12663,N_12939);
xor U14954 (N_14954,N_12643,N_12423);
or U14955 (N_14955,N_13289,N_12560);
nor U14956 (N_14956,N_12378,N_12439);
nor U14957 (N_14957,N_13262,N_13220);
and U14958 (N_14958,N_12779,N_12013);
and U14959 (N_14959,N_13052,N_12400);
xor U14960 (N_14960,N_12809,N_12822);
or U14961 (N_14961,N_12919,N_13479);
nor U14962 (N_14962,N_13352,N_12639);
nand U14963 (N_14963,N_12743,N_13296);
nand U14964 (N_14964,N_12271,N_12484);
and U14965 (N_14965,N_12920,N_12000);
or U14966 (N_14966,N_13206,N_12456);
or U14967 (N_14967,N_12465,N_12885);
nand U14968 (N_14968,N_13093,N_12847);
nor U14969 (N_14969,N_12930,N_12812);
or U14970 (N_14970,N_12506,N_12064);
xnor U14971 (N_14971,N_13050,N_13005);
nand U14972 (N_14972,N_13228,N_12661);
xor U14973 (N_14973,N_13484,N_12630);
nor U14974 (N_14974,N_13417,N_12902);
xnor U14975 (N_14975,N_12627,N_12148);
nor U14976 (N_14976,N_12936,N_12046);
or U14977 (N_14977,N_13247,N_13272);
nand U14978 (N_14978,N_13087,N_12893);
or U14979 (N_14979,N_13081,N_13133);
nor U14980 (N_14980,N_12657,N_12728);
nor U14981 (N_14981,N_12010,N_12530);
nand U14982 (N_14982,N_13361,N_13079);
and U14983 (N_14983,N_13419,N_13420);
nand U14984 (N_14984,N_12740,N_12769);
xor U14985 (N_14985,N_12826,N_12940);
nand U14986 (N_14986,N_12319,N_12198);
xor U14987 (N_14987,N_12198,N_13388);
nand U14988 (N_14988,N_12335,N_12185);
and U14989 (N_14989,N_12788,N_12573);
or U14990 (N_14990,N_12126,N_12345);
xnor U14991 (N_14991,N_12759,N_13220);
and U14992 (N_14992,N_12936,N_13375);
xnor U14993 (N_14993,N_12515,N_12488);
and U14994 (N_14994,N_12143,N_12458);
and U14995 (N_14995,N_13310,N_13071);
xnor U14996 (N_14996,N_13160,N_12999);
or U14997 (N_14997,N_12741,N_12116);
and U14998 (N_14998,N_13372,N_12722);
nor U14999 (N_14999,N_12389,N_12921);
and UO_0 (O_0,N_13912,N_13755);
nand UO_1 (O_1,N_13794,N_14215);
or UO_2 (O_2,N_13838,N_14029);
or UO_3 (O_3,N_14532,N_14523);
and UO_4 (O_4,N_14928,N_14842);
nand UO_5 (O_5,N_14078,N_14915);
nor UO_6 (O_6,N_14982,N_14483);
and UO_7 (O_7,N_14767,N_14236);
and UO_8 (O_8,N_13573,N_13606);
nor UO_9 (O_9,N_13864,N_14542);
nand UO_10 (O_10,N_14299,N_14421);
and UO_11 (O_11,N_14693,N_14156);
nor UO_12 (O_12,N_13968,N_13586);
nor UO_13 (O_13,N_13682,N_13711);
or UO_14 (O_14,N_13665,N_14482);
and UO_15 (O_15,N_14081,N_13767);
and UO_16 (O_16,N_14487,N_14182);
xnor UO_17 (O_17,N_13523,N_14335);
xnor UO_18 (O_18,N_14748,N_13625);
nand UO_19 (O_19,N_13716,N_14402);
xor UO_20 (O_20,N_14471,N_14734);
xnor UO_21 (O_21,N_14418,N_14194);
or UO_22 (O_22,N_14746,N_14427);
nand UO_23 (O_23,N_14862,N_14010);
nor UO_24 (O_24,N_13563,N_14599);
nand UO_25 (O_25,N_14082,N_14525);
nand UO_26 (O_26,N_14229,N_14342);
nand UO_27 (O_27,N_14547,N_13661);
nor UO_28 (O_28,N_14661,N_13712);
nor UO_29 (O_29,N_13868,N_14319);
and UO_30 (O_30,N_14019,N_14390);
nor UO_31 (O_31,N_14637,N_14780);
or UO_32 (O_32,N_14347,N_14958);
or UO_33 (O_33,N_14283,N_14720);
nor UO_34 (O_34,N_14846,N_13527);
xnor UO_35 (O_35,N_14618,N_14646);
xnor UO_36 (O_36,N_14249,N_13690);
and UO_37 (O_37,N_13604,N_14442);
nand UO_38 (O_38,N_13674,N_14709);
nand UO_39 (O_39,N_14635,N_13706);
or UO_40 (O_40,N_13526,N_13939);
nor UO_41 (O_41,N_13766,N_14987);
and UO_42 (O_42,N_13559,N_13827);
xor UO_43 (O_43,N_13621,N_14821);
and UO_44 (O_44,N_14456,N_14682);
or UO_45 (O_45,N_14015,N_14929);
or UO_46 (O_46,N_14736,N_13929);
nand UO_47 (O_47,N_14341,N_14975);
or UO_48 (O_48,N_14159,N_13779);
nor UO_49 (O_49,N_14038,N_13544);
and UO_50 (O_50,N_13558,N_14680);
and UO_51 (O_51,N_14793,N_14073);
and UO_52 (O_52,N_13576,N_14104);
nor UO_53 (O_53,N_13956,N_14835);
nor UO_54 (O_54,N_14548,N_13948);
nand UO_55 (O_55,N_14932,N_14004);
and UO_56 (O_56,N_14927,N_14117);
and UO_57 (O_57,N_14819,N_14749);
xor UO_58 (O_58,N_14853,N_13572);
and UO_59 (O_59,N_13550,N_13699);
or UO_60 (O_60,N_13945,N_14624);
or UO_61 (O_61,N_14142,N_14559);
and UO_62 (O_62,N_14292,N_14764);
and UO_63 (O_63,N_13842,N_14383);
or UO_64 (O_64,N_14959,N_14552);
nand UO_65 (O_65,N_14450,N_14437);
or UO_66 (O_66,N_14477,N_14337);
xnor UO_67 (O_67,N_14707,N_14951);
nor UO_68 (O_68,N_14275,N_13640);
nand UO_69 (O_69,N_13598,N_14562);
nor UO_70 (O_70,N_14847,N_14742);
nor UO_71 (O_71,N_13782,N_14352);
and UO_72 (O_72,N_14502,N_14365);
xor UO_73 (O_73,N_14955,N_13618);
and UO_74 (O_74,N_13960,N_14815);
nor UO_75 (O_75,N_14705,N_13748);
nand UO_76 (O_76,N_13677,N_14211);
nand UO_77 (O_77,N_14409,N_13727);
nand UO_78 (O_78,N_14558,N_14568);
nor UO_79 (O_79,N_14290,N_14253);
or UO_80 (O_80,N_14565,N_13928);
nand UO_81 (O_81,N_13543,N_14270);
xnor UO_82 (O_82,N_13944,N_13796);
nor UO_83 (O_83,N_14630,N_14257);
nand UO_84 (O_84,N_14428,N_13565);
xnor UO_85 (O_85,N_14787,N_14580);
or UO_86 (O_86,N_14900,N_13505);
or UO_87 (O_87,N_13693,N_13547);
or UO_88 (O_88,N_14578,N_14322);
xnor UO_89 (O_89,N_13763,N_13892);
or UO_90 (O_90,N_14093,N_13684);
nor UO_91 (O_91,N_13740,N_14612);
nor UO_92 (O_92,N_14118,N_13687);
nand UO_93 (O_93,N_14687,N_14028);
and UO_94 (O_94,N_14632,N_13795);
and UO_95 (O_95,N_14834,N_14940);
xnor UO_96 (O_96,N_14917,N_13719);
or UO_97 (O_97,N_13847,N_14776);
and UO_98 (O_98,N_13504,N_14839);
xor UO_99 (O_99,N_14364,N_13869);
nor UO_100 (O_100,N_13774,N_13783);
and UO_101 (O_101,N_14030,N_14638);
and UO_102 (O_102,N_13828,N_13787);
xor UO_103 (O_103,N_14035,N_13646);
or UO_104 (O_104,N_13845,N_14094);
or UO_105 (O_105,N_13549,N_13958);
and UO_106 (O_106,N_13546,N_13679);
nand UO_107 (O_107,N_13932,N_13975);
or UO_108 (O_108,N_13871,N_14091);
nand UO_109 (O_109,N_14269,N_13867);
nor UO_110 (O_110,N_14317,N_14902);
nor UO_111 (O_111,N_14145,N_14563);
nor UO_112 (O_112,N_14763,N_14098);
and UO_113 (O_113,N_13894,N_13854);
or UO_114 (O_114,N_13822,N_14789);
or UO_115 (O_115,N_14704,N_13681);
nor UO_116 (O_116,N_13966,N_13715);
or UO_117 (O_117,N_13557,N_14325);
and UO_118 (O_118,N_14645,N_14235);
nand UO_119 (O_119,N_13610,N_14639);
and UO_120 (O_120,N_13694,N_13678);
or UO_121 (O_121,N_14058,N_14895);
or UO_122 (O_122,N_14907,N_14076);
nor UO_123 (O_123,N_14261,N_14198);
nor UO_124 (O_124,N_14306,N_14822);
or UO_125 (O_125,N_14621,N_13628);
nor UO_126 (O_126,N_14230,N_14738);
xor UO_127 (O_127,N_14491,N_14114);
and UO_128 (O_128,N_14173,N_14713);
nand UO_129 (O_129,N_14260,N_14263);
nand UO_130 (O_130,N_14202,N_14647);
nand UO_131 (O_131,N_14980,N_14121);
or UO_132 (O_132,N_14891,N_13617);
or UO_133 (O_133,N_14598,N_13751);
nor UO_134 (O_134,N_14254,N_14960);
nor UO_135 (O_135,N_14640,N_13756);
or UO_136 (O_136,N_13829,N_14659);
nor UO_137 (O_137,N_14488,N_14622);
xnor UO_138 (O_138,N_13629,N_14034);
nand UO_139 (O_139,N_14836,N_14675);
nand UO_140 (O_140,N_14494,N_14773);
and UO_141 (O_141,N_13962,N_14222);
xor UO_142 (O_142,N_14995,N_14313);
xnor UO_143 (O_143,N_14361,N_14054);
or UO_144 (O_144,N_14685,N_14324);
xor UO_145 (O_145,N_14810,N_14625);
or UO_146 (O_146,N_14459,N_14535);
and UO_147 (O_147,N_14554,N_14543);
xnor UO_148 (O_148,N_14381,N_14865);
nand UO_149 (O_149,N_13902,N_14095);
or UO_150 (O_150,N_13908,N_14237);
and UO_151 (O_151,N_14153,N_13930);
nor UO_152 (O_152,N_13667,N_14399);
or UO_153 (O_153,N_14965,N_14389);
or UO_154 (O_154,N_14392,N_13865);
nand UO_155 (O_155,N_14226,N_14188);
nor UO_156 (O_156,N_14144,N_14003);
or UO_157 (O_157,N_14654,N_14608);
and UO_158 (O_158,N_14728,N_13556);
xnor UO_159 (O_159,N_13512,N_13717);
nand UO_160 (O_160,N_13599,N_14688);
and UO_161 (O_161,N_14162,N_14820);
and UO_162 (O_162,N_14896,N_13809);
nand UO_163 (O_163,N_14681,N_13529);
xnor UO_164 (O_164,N_13605,N_13596);
or UO_165 (O_165,N_13722,N_13655);
and UO_166 (O_166,N_14122,N_13639);
nand UO_167 (O_167,N_13554,N_13891);
or UO_168 (O_168,N_13876,N_14777);
and UO_169 (O_169,N_14962,N_14400);
xnor UO_170 (O_170,N_14985,N_14885);
nand UO_171 (O_171,N_13843,N_14045);
nand UO_172 (O_172,N_14924,N_14379);
and UO_173 (O_173,N_14724,N_14234);
nand UO_174 (O_174,N_14462,N_14786);
xnor UO_175 (O_175,N_14683,N_14610);
nand UO_176 (O_176,N_13934,N_13768);
or UO_177 (O_177,N_14583,N_14997);
or UO_178 (O_178,N_14013,N_14336);
nand UO_179 (O_179,N_13824,N_14258);
xor UO_180 (O_180,N_14343,N_14219);
or UO_181 (O_181,N_14520,N_14022);
nor UO_182 (O_182,N_14047,N_14151);
nor UO_183 (O_183,N_14373,N_13832);
or UO_184 (O_184,N_13773,N_13710);
and UO_185 (O_185,N_13887,N_13642);
xnor UO_186 (O_186,N_14027,N_14199);
nand UO_187 (O_187,N_13582,N_14735);
nor UO_188 (O_188,N_14790,N_14143);
or UO_189 (O_189,N_14077,N_14575);
xor UO_190 (O_190,N_14075,N_14321);
nor UO_191 (O_191,N_14910,N_14760);
nor UO_192 (O_192,N_13612,N_14444);
or UO_193 (O_193,N_14613,N_14032);
and UO_194 (O_194,N_14248,N_14129);
xor UO_195 (O_195,N_14676,N_14544);
xor UO_196 (O_196,N_13519,N_14064);
nor UO_197 (O_197,N_13844,N_14939);
nor UO_198 (O_198,N_14089,N_14818);
nand UO_199 (O_199,N_13890,N_13652);
nor UO_200 (O_200,N_14983,N_14438);
and UO_201 (O_201,N_13630,N_13859);
or UO_202 (O_202,N_14863,N_13817);
nor UO_203 (O_203,N_14731,N_14148);
and UO_204 (O_204,N_14036,N_14696);
xnor UO_205 (O_205,N_13870,N_14545);
nand UO_206 (O_206,N_14870,N_13562);
or UO_207 (O_207,N_14062,N_13762);
nand UO_208 (O_208,N_14715,N_13744);
xor UO_209 (O_209,N_14137,N_13814);
and UO_210 (O_210,N_14376,N_14287);
and UO_211 (O_211,N_14800,N_14706);
and UO_212 (O_212,N_14577,N_14909);
nor UO_213 (O_213,N_14684,N_13726);
nor UO_214 (O_214,N_14455,N_13982);
xor UO_215 (O_215,N_13786,N_13996);
xor UO_216 (O_216,N_14918,N_14490);
nor UO_217 (O_217,N_14852,N_13953);
nor UO_218 (O_218,N_14353,N_13641);
nand UO_219 (O_219,N_14416,N_14296);
xnor UO_220 (O_220,N_13917,N_14553);
or UO_221 (O_221,N_14286,N_14701);
and UO_222 (O_222,N_13853,N_14623);
nor UO_223 (O_223,N_13728,N_14858);
nand UO_224 (O_224,N_13739,N_13607);
nand UO_225 (O_225,N_14061,N_13539);
nor UO_226 (O_226,N_14439,N_14627);
xnor UO_227 (O_227,N_14546,N_14006);
xnor UO_228 (O_228,N_14005,N_14468);
nor UO_229 (O_229,N_14138,N_13800);
nand UO_230 (O_230,N_14719,N_14328);
or UO_231 (O_231,N_14057,N_14653);
nor UO_232 (O_232,N_14050,N_13803);
nor UO_233 (O_233,N_13517,N_14743);
nand UO_234 (O_234,N_14887,N_14305);
xnor UO_235 (O_235,N_14864,N_13925);
xnor UO_236 (O_236,N_13935,N_14566);
and UO_237 (O_237,N_14241,N_13812);
nor UO_238 (O_238,N_14903,N_14316);
xor UO_239 (O_239,N_14043,N_13963);
nand UO_240 (O_240,N_14919,N_14830);
and UO_241 (O_241,N_13664,N_13899);
or UO_242 (O_242,N_14679,N_14528);
nor UO_243 (O_243,N_14425,N_14240);
xor UO_244 (O_244,N_14186,N_13993);
nor UO_245 (O_245,N_14424,N_13904);
xor UO_246 (O_246,N_13926,N_13988);
and UO_247 (O_247,N_14407,N_14880);
or UO_248 (O_248,N_13602,N_14904);
nand UO_249 (O_249,N_14849,N_14515);
xor UO_250 (O_250,N_13734,N_14377);
or UO_251 (O_251,N_14605,N_13542);
xnor UO_252 (O_252,N_13759,N_14218);
xnor UO_253 (O_253,N_13613,N_13709);
xor UO_254 (O_254,N_13695,N_14843);
xnor UO_255 (O_255,N_14185,N_14170);
xnor UO_256 (O_256,N_14898,N_14785);
xnor UO_257 (O_257,N_13737,N_13893);
xnor UO_258 (O_258,N_14517,N_14410);
and UO_259 (O_259,N_14309,N_14158);
and UO_260 (O_260,N_14912,N_14498);
or UO_261 (O_261,N_14658,N_14938);
and UO_262 (O_262,N_14856,N_14833);
or UO_263 (O_263,N_13634,N_14301);
or UO_264 (O_264,N_14448,N_13861);
nor UO_265 (O_265,N_13616,N_14059);
nand UO_266 (O_266,N_14534,N_14519);
or UO_267 (O_267,N_13910,N_14901);
xnor UO_268 (O_268,N_14990,N_14970);
or UO_269 (O_269,N_13878,N_13729);
or UO_270 (O_270,N_13658,N_14092);
nor UO_271 (O_271,N_13820,N_13707);
or UO_272 (O_272,N_14817,N_14845);
and UO_273 (O_273,N_13897,N_14044);
xor UO_274 (O_274,N_14323,N_14964);
nor UO_275 (O_275,N_14252,N_13839);
xor UO_276 (O_276,N_14116,N_14799);
xnor UO_277 (O_277,N_14616,N_14803);
xnor UO_278 (O_278,N_14443,N_14832);
nand UO_279 (O_279,N_13834,N_14641);
and UO_280 (O_280,N_13626,N_14436);
and UO_281 (O_281,N_14134,N_14741);
or UO_282 (O_282,N_13997,N_14503);
or UO_283 (O_283,N_13835,N_14505);
and UO_284 (O_284,N_13965,N_13638);
or UO_285 (O_285,N_14769,N_14284);
and UO_286 (O_286,N_14586,N_14048);
nand UO_287 (O_287,N_14518,N_14514);
nand UO_288 (O_288,N_14606,N_14812);
xnor UO_289 (O_289,N_13983,N_13672);
and UO_290 (O_290,N_14126,N_14572);
and UO_291 (O_291,N_14403,N_14355);
and UO_292 (O_292,N_14988,N_14067);
nor UO_293 (O_293,N_13849,N_14472);
xnor UO_294 (O_294,N_14239,N_14085);
nand UO_295 (O_295,N_14667,N_14191);
and UO_296 (O_296,N_14920,N_14366);
or UO_297 (O_297,N_14604,N_14140);
or UO_298 (O_298,N_13992,N_13662);
and UO_299 (O_299,N_13807,N_14972);
nand UO_300 (O_300,N_14851,N_13569);
nor UO_301 (O_301,N_13673,N_13752);
nor UO_302 (O_302,N_14860,N_14538);
nor UO_303 (O_303,N_14423,N_14181);
and UO_304 (O_304,N_13971,N_14691);
nor UO_305 (O_305,N_14349,N_14105);
or UO_306 (O_306,N_13951,N_13575);
or UO_307 (O_307,N_13730,N_14172);
and UO_308 (O_308,N_14937,N_14001);
nor UO_309 (O_309,N_14560,N_13866);
xnor UO_310 (O_310,N_14281,N_14146);
xnor UO_311 (O_311,N_14992,N_13981);
or UO_312 (O_312,N_13804,N_14530);
nand UO_313 (O_313,N_14051,N_14816);
or UO_314 (O_314,N_14584,N_14451);
nand UO_315 (O_315,N_14913,N_14265);
and UO_316 (O_316,N_14086,N_14778);
and UO_317 (O_317,N_14797,N_14978);
and UO_318 (O_318,N_13503,N_14406);
and UO_319 (O_319,N_14993,N_14948);
nor UO_320 (O_320,N_13647,N_14660);
xnor UO_321 (O_321,N_14168,N_14408);
xnor UO_322 (O_322,N_14065,N_14246);
xor UO_323 (O_323,N_13850,N_14233);
nor UO_324 (O_324,N_13903,N_14615);
nand UO_325 (O_325,N_14770,N_14729);
xor UO_326 (O_326,N_13561,N_14429);
nor UO_327 (O_327,N_13581,N_14332);
or UO_328 (O_328,N_13846,N_13521);
or UO_329 (O_329,N_13657,N_13656);
or UO_330 (O_330,N_13723,N_13594);
nand UO_331 (O_331,N_14155,N_14775);
or UO_332 (O_332,N_14204,N_13533);
and UO_333 (O_333,N_14824,N_14811);
or UO_334 (O_334,N_14351,N_13592);
nand UO_335 (O_335,N_14674,N_14650);
or UO_336 (O_336,N_13998,N_14695);
xnor UO_337 (O_337,N_14315,N_14657);
nand UO_338 (O_338,N_14522,N_14597);
nand UO_339 (O_339,N_14310,N_14282);
or UO_340 (O_340,N_13806,N_14678);
nor UO_341 (O_341,N_13636,N_13631);
and UO_342 (O_342,N_13949,N_14823);
nor UO_343 (O_343,N_14132,N_14765);
xor UO_344 (O_344,N_14698,N_13749);
or UO_345 (O_345,N_13659,N_14308);
or UO_346 (O_346,N_14884,N_13911);
nor UO_347 (O_347,N_14434,N_13508);
nor UO_348 (O_348,N_13964,N_14164);
nor UO_349 (O_349,N_13758,N_14348);
nand UO_350 (O_350,N_13689,N_14774);
nor UO_351 (O_351,N_13927,N_14387);
or UO_352 (O_352,N_14949,N_14943);
nor UO_353 (O_353,N_14807,N_14088);
xor UO_354 (O_354,N_14023,N_13648);
nor UO_355 (O_355,N_14298,N_14700);
or UO_356 (O_356,N_14711,N_14669);
xor UO_357 (O_357,N_14014,N_13921);
nand UO_358 (O_358,N_13972,N_13595);
nor UO_359 (O_359,N_14031,N_13879);
xor UO_360 (O_360,N_13551,N_14721);
or UO_361 (O_361,N_13761,N_14579);
xor UO_362 (O_362,N_14431,N_14644);
xor UO_363 (O_363,N_14320,N_14208);
and UO_364 (O_364,N_14374,N_14363);
nor UO_365 (O_365,N_14716,N_13528);
xnor UO_366 (O_366,N_13898,N_14723);
xor UO_367 (O_367,N_14485,N_14703);
nor UO_368 (O_368,N_13841,N_14386);
or UO_369 (O_369,N_14794,N_14504);
and UO_370 (O_370,N_14561,N_13645);
nor UO_371 (O_371,N_13885,N_13671);
nand UO_372 (O_372,N_14809,N_13946);
nand UO_373 (O_373,N_13651,N_13815);
nand UO_374 (O_374,N_13697,N_13770);
and UO_375 (O_375,N_13520,N_14521);
nand UO_376 (O_376,N_13905,N_14784);
nand UO_377 (O_377,N_13703,N_14634);
nor UO_378 (O_378,N_14344,N_14469);
xor UO_379 (O_379,N_13819,N_14694);
nor UO_380 (O_380,N_13784,N_14533);
nand UO_381 (O_381,N_14877,N_14021);
and UO_382 (O_382,N_14072,N_14489);
nand UO_383 (O_383,N_13637,N_13788);
nor UO_384 (O_384,N_13942,N_14607);
xor UO_385 (O_385,N_13781,N_14228);
nand UO_386 (O_386,N_14147,N_13793);
nor UO_387 (O_387,N_13955,N_14666);
nor UO_388 (O_388,N_14360,N_14190);
nor UO_389 (O_389,N_14274,N_13511);
nor UO_390 (O_390,N_14529,N_14025);
nor UO_391 (O_391,N_13852,N_14161);
or UO_392 (O_392,N_13797,N_14220);
nand UO_393 (O_393,N_14276,N_14259);
nor UO_394 (O_394,N_14739,N_14433);
xor UO_395 (O_395,N_14755,N_14113);
nand UO_396 (O_396,N_13745,N_13848);
or UO_397 (O_397,N_13531,N_14404);
nand UO_398 (O_398,N_13747,N_14189);
nand UO_399 (O_399,N_14484,N_14699);
and UO_400 (O_400,N_14730,N_14102);
nor UO_401 (O_401,N_13863,N_14060);
or UO_402 (O_402,N_14664,N_13877);
xnor UO_403 (O_403,N_14447,N_14278);
nor UO_404 (O_404,N_13514,N_14378);
and UO_405 (O_405,N_14672,N_14670);
xor UO_406 (O_406,N_13743,N_14180);
and UO_407 (O_407,N_14506,N_14592);
nand UO_408 (O_408,N_14339,N_14593);
nor UO_409 (O_409,N_14708,N_14453);
nand UO_410 (O_410,N_14976,N_14643);
xor UO_411 (O_411,N_13980,N_13660);
and UO_412 (O_412,N_13990,N_14123);
xnor UO_413 (O_413,N_14435,N_14908);
and UO_414 (O_414,N_14984,N_13913);
or UO_415 (O_415,N_14867,N_13959);
or UO_416 (O_416,N_13583,N_14131);
xnor UO_417 (O_417,N_14850,N_14686);
nor UO_418 (O_418,N_13686,N_13801);
nor UO_419 (O_419,N_14890,N_13650);
and UO_420 (O_420,N_13833,N_14074);
nand UO_421 (O_421,N_13915,N_14963);
and UO_422 (O_422,N_13669,N_13936);
or UO_423 (O_423,N_14130,N_14124);
nand UO_424 (O_424,N_13874,N_14590);
nor UO_425 (O_425,N_13775,N_14969);
xnor UO_426 (O_426,N_14411,N_14367);
and UO_427 (O_427,N_14798,N_14017);
nand UO_428 (O_428,N_14837,N_14537);
nand UO_429 (O_429,N_14508,N_14999);
or UO_430 (O_430,N_13813,N_14245);
and UO_431 (O_431,N_14855,N_14750);
xnor UO_432 (O_432,N_13978,N_13567);
or UO_433 (O_433,N_14087,N_13808);
or UO_434 (O_434,N_14271,N_14571);
xor UO_435 (O_435,N_14068,N_14649);
and UO_436 (O_436,N_13830,N_13916);
and UO_437 (O_437,N_13920,N_14805);
nor UO_438 (O_438,N_13805,N_14049);
or UO_439 (O_439,N_14854,N_14016);
nand UO_440 (O_440,N_14210,N_13516);
xnor UO_441 (O_441,N_14175,N_13931);
and UO_442 (O_442,N_14217,N_14930);
nor UO_443 (O_443,N_13705,N_14163);
and UO_444 (O_444,N_13714,N_14499);
xnor UO_445 (O_445,N_14971,N_14385);
xnor UO_446 (O_446,N_14398,N_14925);
xor UO_447 (O_447,N_14868,N_14633);
nand UO_448 (O_448,N_14779,N_14648);
nor UO_449 (O_449,N_14977,N_13746);
nor UO_450 (O_450,N_13940,N_14394);
nor UO_451 (O_451,N_14771,N_14289);
nand UO_452 (O_452,N_14268,N_13535);
or UO_453 (O_453,N_13889,N_14203);
nor UO_454 (O_454,N_13969,N_13560);
nand UO_455 (O_455,N_14629,N_14100);
nor UO_456 (O_456,N_13579,N_14187);
or UO_457 (O_457,N_13721,N_13973);
nor UO_458 (O_458,N_13574,N_14345);
and UO_459 (O_459,N_14710,N_13534);
or UO_460 (O_460,N_13633,N_14871);
and UO_461 (O_461,N_14338,N_13663);
nand UO_462 (O_462,N_14178,N_13875);
nor UO_463 (O_463,N_14556,N_14944);
nor UO_464 (O_464,N_14702,N_14464);
xor UO_465 (O_465,N_13541,N_13831);
nand UO_466 (O_466,N_14136,N_13591);
nor UO_467 (O_467,N_14619,N_14829);
or UO_468 (O_468,N_14751,N_13799);
nand UO_469 (O_469,N_14201,N_14492);
xor UO_470 (O_470,N_14112,N_13536);
nand UO_471 (O_471,N_14327,N_13622);
and UO_472 (O_472,N_14781,N_14465);
or UO_473 (O_473,N_14242,N_14594);
nand UO_474 (O_474,N_13950,N_13580);
and UO_475 (O_475,N_14934,N_14974);
xor UO_476 (O_476,N_14294,N_13666);
xor UO_477 (O_477,N_14446,N_13644);
and UO_478 (O_478,N_14454,N_13584);
nand UO_479 (O_479,N_13552,N_14596);
or UO_480 (O_480,N_14079,N_14279);
and UO_481 (O_481,N_14026,N_14002);
nand UO_482 (O_482,N_14573,N_14224);
xor UO_483 (O_483,N_14587,N_14848);
nor UO_484 (O_484,N_13957,N_14838);
nor UO_485 (O_485,N_14330,N_13670);
nor UO_486 (O_486,N_14954,N_14422);
nor UO_487 (O_487,N_13954,N_13914);
xor UO_488 (O_488,N_13810,N_14101);
and UO_489 (O_489,N_14569,N_14441);
xor UO_490 (O_490,N_14133,N_14782);
or UO_491 (O_491,N_13900,N_14602);
nand UO_492 (O_492,N_14382,N_13733);
nor UO_493 (O_493,N_13738,N_14359);
nand UO_494 (O_494,N_14052,N_13718);
nand UO_495 (O_495,N_14350,N_14166);
nand UO_496 (O_496,N_14397,N_14620);
xnor UO_497 (O_497,N_13943,N_13789);
nor UO_498 (O_498,N_14183,N_14549);
and UO_499 (O_499,N_14501,N_14717);
nand UO_500 (O_500,N_14762,N_14894);
xor UO_501 (O_501,N_14857,N_14412);
and UO_502 (O_502,N_14756,N_14631);
xnor UO_503 (O_503,N_13919,N_13961);
and UO_504 (O_504,N_14212,N_14952);
nor UO_505 (O_505,N_13589,N_14665);
nand UO_506 (O_506,N_13568,N_14950);
nand UO_507 (O_507,N_14574,N_14250);
nand UO_508 (O_508,N_13600,N_13704);
xnor UO_509 (O_509,N_13750,N_14426);
nor UO_510 (O_510,N_14346,N_13776);
or UO_511 (O_511,N_14888,N_14110);
xnor UO_512 (O_512,N_14063,N_14989);
xnor UO_513 (O_513,N_14831,N_14262);
nor UO_514 (O_514,N_14302,N_14041);
nor UO_515 (O_515,N_14961,N_14905);
nor UO_516 (O_516,N_14576,N_14801);
or UO_517 (O_517,N_14991,N_14527);
and UO_518 (O_518,N_13924,N_14589);
or UO_519 (O_519,N_14120,N_14152);
nor UO_520 (O_520,N_14221,N_14474);
xnor UO_521 (O_521,N_14956,N_13974);
and UO_522 (O_522,N_14526,N_14042);
nand UO_523 (O_523,N_14725,N_14024);
nand UO_524 (O_524,N_14998,N_14267);
xor UO_525 (O_525,N_13923,N_14923);
or UO_526 (O_526,N_14000,N_14994);
nor UO_527 (O_527,N_14968,N_14209);
nand UO_528 (O_528,N_14184,N_13873);
xnor UO_529 (O_529,N_14318,N_14628);
and UO_530 (O_530,N_14813,N_13995);
nand UO_531 (O_531,N_14295,N_14311);
or UO_532 (O_532,N_13609,N_13862);
nand UO_533 (O_533,N_13984,N_14996);
nor UO_534 (O_534,N_13922,N_13764);
nor UO_535 (O_535,N_13872,N_13700);
or UO_536 (O_536,N_14591,N_14967);
or UO_537 (O_537,N_13588,N_14914);
or UO_538 (O_538,N_14496,N_14280);
xnor UO_539 (O_539,N_13702,N_13624);
nor UO_540 (O_540,N_14802,N_14873);
nand UO_541 (O_541,N_13537,N_14882);
xnor UO_542 (O_542,N_14795,N_14935);
nand UO_543 (O_543,N_13724,N_14109);
xor UO_544 (O_544,N_14712,N_14759);
nand UO_545 (O_545,N_13851,N_14570);
xnor UO_546 (O_546,N_13593,N_14757);
xnor UO_547 (O_547,N_14177,N_14167);
nand UO_548 (O_548,N_13947,N_14277);
xor UO_549 (O_549,N_14354,N_13792);
nor UO_550 (O_550,N_14745,N_14405);
or UO_551 (O_551,N_14479,N_13888);
nand UO_552 (O_552,N_14766,N_14582);
or UO_553 (O_553,N_14369,N_14466);
and UO_554 (O_554,N_13510,N_13696);
nor UO_555 (O_555,N_14154,N_13668);
and UO_556 (O_556,N_14460,N_14886);
xor UO_557 (O_557,N_13675,N_14497);
nor UO_558 (O_558,N_14792,N_13577);
nor UO_559 (O_559,N_14103,N_14033);
nand UO_560 (O_560,N_14192,N_14476);
or UO_561 (O_561,N_14744,N_14911);
and UO_562 (O_562,N_13530,N_13698);
and UO_563 (O_563,N_14291,N_13985);
or UO_564 (O_564,N_13635,N_14733);
or UO_565 (O_565,N_13601,N_14371);
and UO_566 (O_566,N_14127,N_14106);
xnor UO_567 (O_567,N_13909,N_14358);
and UO_568 (O_568,N_13976,N_14722);
nor UO_569 (O_569,N_14018,N_14238);
nor UO_570 (O_570,N_13685,N_13735);
xor UO_571 (O_571,N_13725,N_14331);
and UO_572 (O_572,N_14196,N_13823);
nand UO_573 (O_573,N_14356,N_14334);
nor UO_574 (O_574,N_14273,N_14636);
nand UO_575 (O_575,N_14897,N_14141);
xor UO_576 (O_576,N_14340,N_14551);
nand UO_577 (O_577,N_14892,N_13676);
and UO_578 (O_578,N_13811,N_14677);
or UO_579 (O_579,N_14080,N_14171);
nor UO_580 (O_580,N_14304,N_14247);
or UO_581 (O_581,N_14899,N_14889);
or UO_582 (O_582,N_14285,N_13578);
nand UO_583 (O_583,N_14207,N_14804);
nor UO_584 (O_584,N_14826,N_14176);
and UO_585 (O_585,N_14288,N_14473);
nand UO_586 (O_586,N_13986,N_13882);
nand UO_587 (O_587,N_14157,N_14941);
xnor UO_588 (O_588,N_14714,N_14524);
nor UO_589 (O_589,N_13857,N_14009);
nor UO_590 (O_590,N_13713,N_14244);
nand UO_591 (O_591,N_14223,N_13515);
nor UO_592 (O_592,N_13691,N_14174);
xnor UO_593 (O_593,N_14243,N_14329);
nand UO_594 (O_594,N_13540,N_14642);
xor UO_595 (O_595,N_14981,N_14979);
xor UO_596 (O_596,N_13979,N_14791);
or UO_597 (O_597,N_14869,N_14541);
nand UO_598 (O_598,N_13856,N_13608);
nor UO_599 (O_599,N_13826,N_14946);
nor UO_600 (O_600,N_14933,N_13614);
xor UO_601 (O_601,N_13500,N_14752);
or UO_602 (O_602,N_14205,N_13785);
nand UO_603 (O_603,N_14690,N_14652);
xnor UO_604 (O_604,N_13896,N_14445);
xnor UO_605 (O_605,N_14264,N_14070);
and UO_606 (O_606,N_14747,N_14603);
or UO_607 (O_607,N_14084,N_14461);
or UO_608 (O_608,N_14370,N_14673);
xor UO_609 (O_609,N_13918,N_14216);
and UO_610 (O_610,N_14926,N_13731);
or UO_611 (O_611,N_14539,N_13692);
xnor UO_612 (O_612,N_14689,N_14357);
nand UO_613 (O_613,N_14071,N_14768);
xor UO_614 (O_614,N_14375,N_14772);
xnor UO_615 (O_615,N_13901,N_14139);
and UO_616 (O_616,N_14303,N_14881);
or UO_617 (O_617,N_14761,N_13502);
or UO_618 (O_618,N_14256,N_13825);
or UO_619 (O_619,N_13571,N_14942);
xor UO_620 (O_620,N_14957,N_14307);
nor UO_621 (O_621,N_13507,N_14825);
or UO_622 (O_622,N_14866,N_14040);
nand UO_623 (O_623,N_13952,N_14395);
xor UO_624 (O_624,N_13790,N_14195);
and UO_625 (O_625,N_14945,N_14160);
or UO_626 (O_626,N_14878,N_14449);
xnor UO_627 (O_627,N_13720,N_14135);
and UO_628 (O_628,N_14214,N_14844);
or UO_629 (O_629,N_14401,N_14536);
xor UO_630 (O_630,N_14372,N_14883);
xor UO_631 (O_631,N_13615,N_13532);
and UO_632 (O_632,N_14452,N_13818);
nor UO_633 (O_633,N_14922,N_14251);
nand UO_634 (O_634,N_13570,N_14614);
nor UO_635 (O_635,N_13736,N_14861);
nand UO_636 (O_636,N_14314,N_14663);
xnor UO_637 (O_637,N_14718,N_13778);
and UO_638 (O_638,N_14827,N_14165);
nor UO_639 (O_639,N_13836,N_14272);
xnor UO_640 (O_640,N_13632,N_14232);
and UO_641 (O_641,N_13880,N_13989);
xnor UO_642 (O_642,N_14225,N_14872);
nor UO_643 (O_643,N_13654,N_13741);
nand UO_644 (O_644,N_14213,N_14480);
xnor UO_645 (O_645,N_13884,N_14227);
or UO_646 (O_646,N_14169,N_14737);
nor UO_647 (O_647,N_13643,N_14107);
xnor UO_648 (O_648,N_14312,N_13907);
nor UO_649 (O_649,N_14333,N_14893);
and UO_650 (O_650,N_13597,N_14150);
or UO_651 (O_651,N_14326,N_14037);
or UO_652 (O_652,N_13837,N_14056);
and UO_653 (O_653,N_14115,N_14754);
nor UO_654 (O_654,N_14007,N_14732);
xor UO_655 (O_655,N_13701,N_14656);
nand UO_656 (O_656,N_14564,N_14806);
nand UO_657 (O_657,N_14697,N_13501);
or UO_658 (O_658,N_14783,N_14297);
nand UO_659 (O_659,N_13994,N_14513);
xor UO_660 (O_660,N_14111,N_14300);
or UO_661 (O_661,N_14193,N_14986);
xor UO_662 (O_662,N_14875,N_14531);
and UO_663 (O_663,N_14417,N_14097);
nand UO_664 (O_664,N_13545,N_13881);
nor UO_665 (O_665,N_13816,N_13585);
or UO_666 (O_666,N_14197,N_14510);
nand UO_667 (O_667,N_14415,N_14692);
and UO_668 (O_668,N_14493,N_14478);
nand UO_669 (O_669,N_13883,N_14090);
and UO_670 (O_670,N_14662,N_13590);
and UO_671 (O_671,N_13895,N_14758);
xor UO_672 (O_672,N_13970,N_14581);
and UO_673 (O_673,N_14511,N_14947);
nand UO_674 (O_674,N_14083,N_14481);
or UO_675 (O_675,N_14727,N_14393);
nor UO_676 (O_676,N_13933,N_14516);
nor UO_677 (O_677,N_14486,N_14206);
xor UO_678 (O_678,N_14600,N_14966);
xor UO_679 (O_679,N_13821,N_13937);
nand UO_680 (O_680,N_13753,N_14020);
xor UO_681 (O_681,N_14814,N_13509);
and UO_682 (O_682,N_14557,N_14828);
nor UO_683 (O_683,N_14396,N_14921);
or UO_684 (O_684,N_14796,N_13798);
nand UO_685 (O_685,N_13587,N_14108);
nand UO_686 (O_686,N_14179,N_14266);
nand UO_687 (O_687,N_13777,N_14430);
nor UO_688 (O_688,N_14149,N_14128);
nor UO_689 (O_689,N_13688,N_14053);
or UO_690 (O_690,N_14011,N_14231);
xor UO_691 (O_691,N_14540,N_13649);
xnor UO_692 (O_692,N_13858,N_14859);
nand UO_693 (O_693,N_14626,N_14008);
and UO_694 (O_694,N_14906,N_14841);
or UO_695 (O_695,N_14611,N_13772);
nand UO_696 (O_696,N_14507,N_14788);
nand UO_697 (O_697,N_13522,N_14726);
nor UO_698 (O_698,N_13708,N_14512);
xor UO_699 (O_699,N_13802,N_13991);
or UO_700 (O_700,N_14384,N_13603);
nor UO_701 (O_701,N_13683,N_14457);
or UO_702 (O_702,N_13765,N_13886);
nor UO_703 (O_703,N_14099,N_13999);
or UO_704 (O_704,N_14931,N_13620);
xnor UO_705 (O_705,N_14125,N_13555);
xor UO_706 (O_706,N_14874,N_14255);
nand UO_707 (O_707,N_14039,N_13754);
and UO_708 (O_708,N_13941,N_14420);
or UO_709 (O_709,N_14470,N_14419);
and UO_710 (O_710,N_13769,N_14585);
nor UO_711 (O_711,N_14808,N_14055);
nor UO_712 (O_712,N_14119,N_13987);
xor UO_713 (O_713,N_14671,N_14500);
xor UO_714 (O_714,N_13757,N_14293);
and UO_715 (O_715,N_13906,N_13977);
nor UO_716 (O_716,N_13732,N_13967);
nand UO_717 (O_717,N_14655,N_13619);
or UO_718 (O_718,N_13524,N_13548);
and UO_719 (O_719,N_13525,N_14550);
xnor UO_720 (O_720,N_14601,N_14588);
nor UO_721 (O_721,N_13791,N_13855);
nand UO_722 (O_722,N_13623,N_14368);
nand UO_723 (O_723,N_13771,N_13513);
nor UO_724 (O_724,N_14567,N_14668);
nand UO_725 (O_725,N_13742,N_14475);
nor UO_726 (O_726,N_14069,N_13653);
nor UO_727 (O_727,N_14753,N_14380);
xor UO_728 (O_728,N_14066,N_14953);
or UO_729 (O_729,N_13840,N_13506);
nand UO_730 (O_730,N_14432,N_14879);
and UO_731 (O_731,N_14046,N_14012);
nor UO_732 (O_732,N_14495,N_14876);
nand UO_733 (O_733,N_14936,N_13938);
nor UO_734 (O_734,N_14362,N_14200);
and UO_735 (O_735,N_14509,N_13553);
xnor UO_736 (O_736,N_13518,N_13680);
or UO_737 (O_737,N_13566,N_13760);
or UO_738 (O_738,N_14414,N_14467);
or UO_739 (O_739,N_13611,N_13538);
nor UO_740 (O_740,N_13780,N_14973);
nand UO_741 (O_741,N_14388,N_14458);
or UO_742 (O_742,N_13564,N_14463);
xor UO_743 (O_743,N_14096,N_14555);
nor UO_744 (O_744,N_14595,N_14617);
or UO_745 (O_745,N_14840,N_14651);
nor UO_746 (O_746,N_14391,N_13860);
and UO_747 (O_747,N_14916,N_14440);
and UO_748 (O_748,N_14609,N_13627);
or UO_749 (O_749,N_14740,N_14413);
or UO_750 (O_750,N_13512,N_14354);
or UO_751 (O_751,N_13647,N_13897);
and UO_752 (O_752,N_14164,N_14822);
or UO_753 (O_753,N_13842,N_14566);
or UO_754 (O_754,N_14196,N_14808);
or UO_755 (O_755,N_13664,N_14695);
and UO_756 (O_756,N_14382,N_14543);
nand UO_757 (O_757,N_14464,N_14071);
xor UO_758 (O_758,N_14988,N_14103);
and UO_759 (O_759,N_13594,N_14736);
xor UO_760 (O_760,N_14377,N_14087);
nand UO_761 (O_761,N_13618,N_14794);
or UO_762 (O_762,N_14678,N_13908);
nor UO_763 (O_763,N_14135,N_14209);
nor UO_764 (O_764,N_14877,N_14268);
nand UO_765 (O_765,N_13608,N_14803);
nor UO_766 (O_766,N_14600,N_13564);
and UO_767 (O_767,N_14108,N_14612);
xor UO_768 (O_768,N_13622,N_14597);
xnor UO_769 (O_769,N_14908,N_13520);
nand UO_770 (O_770,N_14757,N_14593);
and UO_771 (O_771,N_13890,N_14267);
or UO_772 (O_772,N_14776,N_14927);
and UO_773 (O_773,N_14603,N_14326);
xor UO_774 (O_774,N_13648,N_14161);
nand UO_775 (O_775,N_14680,N_14658);
nand UO_776 (O_776,N_13559,N_13870);
nor UO_777 (O_777,N_13562,N_14937);
and UO_778 (O_778,N_14149,N_14359);
nand UO_779 (O_779,N_14768,N_14430);
nor UO_780 (O_780,N_13693,N_14660);
nand UO_781 (O_781,N_13698,N_14206);
or UO_782 (O_782,N_13703,N_14003);
and UO_783 (O_783,N_13823,N_14578);
xnor UO_784 (O_784,N_13756,N_14245);
or UO_785 (O_785,N_14439,N_14576);
nor UO_786 (O_786,N_13926,N_13635);
nor UO_787 (O_787,N_13553,N_14047);
xnor UO_788 (O_788,N_14925,N_14215);
or UO_789 (O_789,N_14095,N_13729);
nor UO_790 (O_790,N_14762,N_13548);
xor UO_791 (O_791,N_13874,N_13702);
nand UO_792 (O_792,N_14226,N_13694);
or UO_793 (O_793,N_14962,N_13506);
nand UO_794 (O_794,N_13968,N_14289);
nor UO_795 (O_795,N_14758,N_14110);
nor UO_796 (O_796,N_14527,N_14252);
nand UO_797 (O_797,N_14805,N_14985);
xor UO_798 (O_798,N_13550,N_13796);
or UO_799 (O_799,N_14079,N_14982);
nand UO_800 (O_800,N_14362,N_13772);
nand UO_801 (O_801,N_14860,N_14592);
nor UO_802 (O_802,N_14005,N_13876);
nor UO_803 (O_803,N_14461,N_14874);
nand UO_804 (O_804,N_14175,N_13542);
nor UO_805 (O_805,N_14424,N_13968);
nor UO_806 (O_806,N_13889,N_14878);
nand UO_807 (O_807,N_13531,N_13786);
nor UO_808 (O_808,N_13521,N_13635);
or UO_809 (O_809,N_14297,N_14652);
nand UO_810 (O_810,N_13591,N_14107);
xnor UO_811 (O_811,N_14401,N_14552);
and UO_812 (O_812,N_14288,N_13993);
and UO_813 (O_813,N_14055,N_13580);
nand UO_814 (O_814,N_13776,N_14832);
nand UO_815 (O_815,N_14137,N_13687);
xor UO_816 (O_816,N_14080,N_14633);
or UO_817 (O_817,N_13887,N_14816);
nor UO_818 (O_818,N_13748,N_14448);
or UO_819 (O_819,N_14097,N_14322);
nor UO_820 (O_820,N_14630,N_14597);
nand UO_821 (O_821,N_14077,N_14932);
or UO_822 (O_822,N_14811,N_14010);
and UO_823 (O_823,N_14135,N_13595);
and UO_824 (O_824,N_13955,N_14720);
and UO_825 (O_825,N_14312,N_14482);
and UO_826 (O_826,N_14904,N_13930);
nand UO_827 (O_827,N_13682,N_13980);
nand UO_828 (O_828,N_14685,N_13787);
and UO_829 (O_829,N_14070,N_13970);
or UO_830 (O_830,N_14347,N_14417);
nor UO_831 (O_831,N_14629,N_14340);
xnor UO_832 (O_832,N_13736,N_14452);
nand UO_833 (O_833,N_14568,N_14815);
nor UO_834 (O_834,N_14922,N_14168);
nand UO_835 (O_835,N_14423,N_14523);
xor UO_836 (O_836,N_13886,N_13982);
nor UO_837 (O_837,N_13629,N_14530);
nor UO_838 (O_838,N_14720,N_14416);
nand UO_839 (O_839,N_13893,N_14601);
nand UO_840 (O_840,N_13590,N_13990);
nand UO_841 (O_841,N_14879,N_14999);
or UO_842 (O_842,N_13534,N_14347);
nand UO_843 (O_843,N_14355,N_14243);
and UO_844 (O_844,N_14696,N_14708);
xnor UO_845 (O_845,N_13574,N_13825);
nor UO_846 (O_846,N_14908,N_14211);
xnor UO_847 (O_847,N_13747,N_13803);
and UO_848 (O_848,N_14926,N_14761);
or UO_849 (O_849,N_14060,N_14731);
and UO_850 (O_850,N_14105,N_14426);
or UO_851 (O_851,N_14415,N_13981);
xnor UO_852 (O_852,N_14496,N_14254);
and UO_853 (O_853,N_14868,N_14768);
nor UO_854 (O_854,N_13997,N_14427);
nor UO_855 (O_855,N_14477,N_14182);
nor UO_856 (O_856,N_13937,N_14646);
nand UO_857 (O_857,N_13991,N_14897);
nor UO_858 (O_858,N_14579,N_13639);
and UO_859 (O_859,N_13881,N_13739);
nand UO_860 (O_860,N_13725,N_13555);
xor UO_861 (O_861,N_14073,N_14579);
and UO_862 (O_862,N_13565,N_13967);
and UO_863 (O_863,N_14840,N_14703);
nor UO_864 (O_864,N_14859,N_13819);
nor UO_865 (O_865,N_13870,N_13517);
nand UO_866 (O_866,N_13583,N_14614);
nand UO_867 (O_867,N_13513,N_14410);
or UO_868 (O_868,N_14101,N_13521);
xor UO_869 (O_869,N_14115,N_13996);
nor UO_870 (O_870,N_14918,N_13901);
nand UO_871 (O_871,N_14868,N_14199);
nor UO_872 (O_872,N_14161,N_13574);
and UO_873 (O_873,N_13610,N_13973);
nor UO_874 (O_874,N_14629,N_14888);
nand UO_875 (O_875,N_14642,N_13518);
nand UO_876 (O_876,N_13987,N_14366);
and UO_877 (O_877,N_14173,N_14296);
or UO_878 (O_878,N_13820,N_14731);
nor UO_879 (O_879,N_14286,N_14273);
or UO_880 (O_880,N_13630,N_14848);
nor UO_881 (O_881,N_13694,N_14784);
xnor UO_882 (O_882,N_13743,N_13868);
xor UO_883 (O_883,N_13691,N_14730);
nor UO_884 (O_884,N_14472,N_14786);
xor UO_885 (O_885,N_13676,N_13679);
nand UO_886 (O_886,N_14881,N_14555);
or UO_887 (O_887,N_14379,N_14186);
nand UO_888 (O_888,N_13971,N_13699);
or UO_889 (O_889,N_13855,N_14486);
nand UO_890 (O_890,N_14783,N_14851);
nor UO_891 (O_891,N_14038,N_14458);
or UO_892 (O_892,N_14582,N_13750);
xor UO_893 (O_893,N_14627,N_13704);
and UO_894 (O_894,N_13610,N_14147);
and UO_895 (O_895,N_14886,N_14341);
xor UO_896 (O_896,N_14384,N_14013);
or UO_897 (O_897,N_14196,N_13748);
xor UO_898 (O_898,N_14960,N_13554);
nand UO_899 (O_899,N_14480,N_14009);
and UO_900 (O_900,N_14678,N_14127);
nor UO_901 (O_901,N_14025,N_13894);
and UO_902 (O_902,N_13953,N_14240);
or UO_903 (O_903,N_14378,N_14523);
nor UO_904 (O_904,N_14980,N_13509);
or UO_905 (O_905,N_13962,N_13585);
and UO_906 (O_906,N_13521,N_14031);
nor UO_907 (O_907,N_13632,N_13782);
xnor UO_908 (O_908,N_14841,N_14832);
nand UO_909 (O_909,N_14971,N_14027);
or UO_910 (O_910,N_14006,N_14291);
nand UO_911 (O_911,N_14516,N_14335);
nand UO_912 (O_912,N_14985,N_14890);
nand UO_913 (O_913,N_14300,N_14289);
and UO_914 (O_914,N_14083,N_14828);
nor UO_915 (O_915,N_14866,N_14293);
or UO_916 (O_916,N_14302,N_13941);
xor UO_917 (O_917,N_14482,N_13547);
and UO_918 (O_918,N_14526,N_14757);
and UO_919 (O_919,N_14330,N_14880);
and UO_920 (O_920,N_13883,N_14187);
and UO_921 (O_921,N_14242,N_14532);
xor UO_922 (O_922,N_14243,N_13985);
and UO_923 (O_923,N_14456,N_13815);
nand UO_924 (O_924,N_13678,N_13890);
nor UO_925 (O_925,N_13938,N_13928);
or UO_926 (O_926,N_14388,N_14427);
nor UO_927 (O_927,N_13838,N_14635);
xor UO_928 (O_928,N_14671,N_14843);
and UO_929 (O_929,N_14363,N_14666);
or UO_930 (O_930,N_14683,N_14284);
nand UO_931 (O_931,N_14044,N_14809);
or UO_932 (O_932,N_14530,N_13964);
xor UO_933 (O_933,N_13614,N_13557);
xor UO_934 (O_934,N_14984,N_14554);
and UO_935 (O_935,N_13750,N_13773);
or UO_936 (O_936,N_14714,N_14756);
and UO_937 (O_937,N_13546,N_13867);
or UO_938 (O_938,N_13974,N_14881);
and UO_939 (O_939,N_14982,N_14921);
and UO_940 (O_940,N_13846,N_14055);
xnor UO_941 (O_941,N_13677,N_14086);
and UO_942 (O_942,N_14969,N_14290);
nor UO_943 (O_943,N_14212,N_14576);
nand UO_944 (O_944,N_14847,N_14884);
nor UO_945 (O_945,N_14322,N_14861);
nor UO_946 (O_946,N_13648,N_14076);
nor UO_947 (O_947,N_13766,N_14633);
xor UO_948 (O_948,N_13829,N_14119);
nand UO_949 (O_949,N_13783,N_13886);
and UO_950 (O_950,N_13963,N_14965);
or UO_951 (O_951,N_13951,N_14588);
nor UO_952 (O_952,N_14976,N_14083);
or UO_953 (O_953,N_13603,N_14342);
nor UO_954 (O_954,N_13711,N_14845);
nor UO_955 (O_955,N_13648,N_14493);
nor UO_956 (O_956,N_13755,N_14399);
nand UO_957 (O_957,N_14381,N_14222);
nand UO_958 (O_958,N_14835,N_14716);
and UO_959 (O_959,N_14238,N_14085);
nand UO_960 (O_960,N_14920,N_14415);
and UO_961 (O_961,N_14983,N_13821);
nor UO_962 (O_962,N_13718,N_13963);
and UO_963 (O_963,N_14825,N_13983);
and UO_964 (O_964,N_13563,N_14089);
xnor UO_965 (O_965,N_13989,N_14882);
or UO_966 (O_966,N_13999,N_13560);
and UO_967 (O_967,N_13777,N_13537);
nor UO_968 (O_968,N_14452,N_14599);
and UO_969 (O_969,N_14857,N_13821);
xor UO_970 (O_970,N_14759,N_13684);
nand UO_971 (O_971,N_14518,N_14060);
nor UO_972 (O_972,N_13610,N_14586);
and UO_973 (O_973,N_14773,N_14584);
and UO_974 (O_974,N_14299,N_14057);
nand UO_975 (O_975,N_14972,N_14120);
or UO_976 (O_976,N_14398,N_13722);
nor UO_977 (O_977,N_13783,N_14178);
xnor UO_978 (O_978,N_14922,N_14815);
nand UO_979 (O_979,N_13614,N_13822);
nor UO_980 (O_980,N_14463,N_14769);
nand UO_981 (O_981,N_14591,N_14182);
xor UO_982 (O_982,N_14688,N_14316);
nand UO_983 (O_983,N_14134,N_14617);
and UO_984 (O_984,N_14571,N_13742);
and UO_985 (O_985,N_14770,N_14492);
xor UO_986 (O_986,N_14073,N_13888);
nor UO_987 (O_987,N_13551,N_14010);
xnor UO_988 (O_988,N_14262,N_14348);
nor UO_989 (O_989,N_14653,N_13814);
or UO_990 (O_990,N_13774,N_14528);
xnor UO_991 (O_991,N_14382,N_14787);
xnor UO_992 (O_992,N_14002,N_14087);
nor UO_993 (O_993,N_14225,N_13936);
or UO_994 (O_994,N_13976,N_13913);
nor UO_995 (O_995,N_14840,N_14509);
or UO_996 (O_996,N_14331,N_14879);
nor UO_997 (O_997,N_13565,N_13660);
nand UO_998 (O_998,N_13948,N_14093);
nor UO_999 (O_999,N_13795,N_14339);
nand UO_1000 (O_1000,N_14385,N_14996);
xnor UO_1001 (O_1001,N_13550,N_14592);
and UO_1002 (O_1002,N_14789,N_14269);
xor UO_1003 (O_1003,N_13631,N_13934);
or UO_1004 (O_1004,N_14428,N_13696);
or UO_1005 (O_1005,N_14414,N_13678);
nand UO_1006 (O_1006,N_13701,N_13587);
nand UO_1007 (O_1007,N_14636,N_14028);
nand UO_1008 (O_1008,N_13547,N_13655);
nand UO_1009 (O_1009,N_14879,N_14035);
xor UO_1010 (O_1010,N_14255,N_13920);
xor UO_1011 (O_1011,N_13611,N_14533);
and UO_1012 (O_1012,N_13928,N_14887);
or UO_1013 (O_1013,N_14297,N_13752);
nor UO_1014 (O_1014,N_13792,N_14505);
nor UO_1015 (O_1015,N_13518,N_14853);
nor UO_1016 (O_1016,N_14735,N_13620);
xor UO_1017 (O_1017,N_13804,N_13962);
nand UO_1018 (O_1018,N_14830,N_14991);
nor UO_1019 (O_1019,N_14150,N_13761);
xnor UO_1020 (O_1020,N_14078,N_13664);
xor UO_1021 (O_1021,N_14416,N_14338);
xnor UO_1022 (O_1022,N_13766,N_13952);
or UO_1023 (O_1023,N_14558,N_13758);
nand UO_1024 (O_1024,N_14248,N_14493);
xor UO_1025 (O_1025,N_14030,N_13941);
or UO_1026 (O_1026,N_13628,N_13998);
nor UO_1027 (O_1027,N_14558,N_14145);
xor UO_1028 (O_1028,N_14329,N_14478);
xor UO_1029 (O_1029,N_14505,N_14669);
or UO_1030 (O_1030,N_14734,N_13515);
nor UO_1031 (O_1031,N_14932,N_13873);
nand UO_1032 (O_1032,N_14528,N_14570);
and UO_1033 (O_1033,N_14808,N_14217);
or UO_1034 (O_1034,N_14100,N_13614);
xnor UO_1035 (O_1035,N_14622,N_14768);
nand UO_1036 (O_1036,N_13883,N_14765);
nor UO_1037 (O_1037,N_13697,N_13881);
xor UO_1038 (O_1038,N_14582,N_14314);
nor UO_1039 (O_1039,N_14849,N_14811);
xnor UO_1040 (O_1040,N_13757,N_13642);
or UO_1041 (O_1041,N_13869,N_13867);
and UO_1042 (O_1042,N_14135,N_14773);
nand UO_1043 (O_1043,N_13998,N_13971);
nor UO_1044 (O_1044,N_13506,N_14344);
nor UO_1045 (O_1045,N_14418,N_14672);
xor UO_1046 (O_1046,N_14499,N_14590);
nor UO_1047 (O_1047,N_14125,N_13668);
or UO_1048 (O_1048,N_14461,N_13711);
and UO_1049 (O_1049,N_13895,N_14289);
and UO_1050 (O_1050,N_14009,N_13834);
or UO_1051 (O_1051,N_13723,N_13576);
nand UO_1052 (O_1052,N_14130,N_13508);
nor UO_1053 (O_1053,N_14751,N_14000);
and UO_1054 (O_1054,N_13704,N_14802);
or UO_1055 (O_1055,N_13621,N_14286);
nor UO_1056 (O_1056,N_14166,N_14187);
nor UO_1057 (O_1057,N_13546,N_14481);
xnor UO_1058 (O_1058,N_14269,N_14160);
nand UO_1059 (O_1059,N_14060,N_13530);
or UO_1060 (O_1060,N_14396,N_14398);
xor UO_1061 (O_1061,N_14148,N_13962);
and UO_1062 (O_1062,N_14342,N_14775);
nor UO_1063 (O_1063,N_13706,N_14296);
and UO_1064 (O_1064,N_14757,N_14244);
xnor UO_1065 (O_1065,N_14906,N_13892);
or UO_1066 (O_1066,N_13957,N_13596);
and UO_1067 (O_1067,N_13731,N_14109);
nor UO_1068 (O_1068,N_14321,N_14577);
nand UO_1069 (O_1069,N_14966,N_13616);
nand UO_1070 (O_1070,N_13791,N_14194);
nor UO_1071 (O_1071,N_14583,N_14683);
nand UO_1072 (O_1072,N_14589,N_14890);
nor UO_1073 (O_1073,N_14209,N_14292);
and UO_1074 (O_1074,N_14103,N_14981);
and UO_1075 (O_1075,N_14033,N_14360);
and UO_1076 (O_1076,N_13651,N_13721);
nand UO_1077 (O_1077,N_14054,N_14834);
nor UO_1078 (O_1078,N_14544,N_14766);
nor UO_1079 (O_1079,N_13621,N_14923);
nor UO_1080 (O_1080,N_13724,N_14386);
nand UO_1081 (O_1081,N_14658,N_13568);
nor UO_1082 (O_1082,N_13586,N_14481);
nor UO_1083 (O_1083,N_13793,N_14404);
nand UO_1084 (O_1084,N_13606,N_14615);
and UO_1085 (O_1085,N_14800,N_13702);
or UO_1086 (O_1086,N_13950,N_14176);
or UO_1087 (O_1087,N_14342,N_13992);
nor UO_1088 (O_1088,N_14610,N_14136);
nand UO_1089 (O_1089,N_14160,N_14246);
xnor UO_1090 (O_1090,N_13957,N_14814);
and UO_1091 (O_1091,N_13587,N_13559);
and UO_1092 (O_1092,N_14253,N_14415);
or UO_1093 (O_1093,N_14342,N_14704);
nand UO_1094 (O_1094,N_13708,N_14430);
nor UO_1095 (O_1095,N_14259,N_14437);
nor UO_1096 (O_1096,N_14412,N_14010);
nand UO_1097 (O_1097,N_14278,N_14597);
nand UO_1098 (O_1098,N_14952,N_14449);
or UO_1099 (O_1099,N_14550,N_13849);
xnor UO_1100 (O_1100,N_14065,N_13551);
or UO_1101 (O_1101,N_14291,N_13686);
and UO_1102 (O_1102,N_14577,N_13865);
xor UO_1103 (O_1103,N_14460,N_13753);
or UO_1104 (O_1104,N_14838,N_13967);
or UO_1105 (O_1105,N_13990,N_14681);
nand UO_1106 (O_1106,N_14609,N_13613);
nand UO_1107 (O_1107,N_14420,N_13802);
nand UO_1108 (O_1108,N_13507,N_14289);
nand UO_1109 (O_1109,N_13615,N_14399);
nand UO_1110 (O_1110,N_14470,N_14693);
and UO_1111 (O_1111,N_14267,N_13976);
nand UO_1112 (O_1112,N_14194,N_14790);
or UO_1113 (O_1113,N_13631,N_14140);
xor UO_1114 (O_1114,N_14655,N_14338);
nor UO_1115 (O_1115,N_13759,N_13611);
and UO_1116 (O_1116,N_13619,N_14174);
nor UO_1117 (O_1117,N_14578,N_14798);
or UO_1118 (O_1118,N_14094,N_13631);
and UO_1119 (O_1119,N_14030,N_14864);
nor UO_1120 (O_1120,N_14994,N_13627);
and UO_1121 (O_1121,N_14111,N_14335);
xor UO_1122 (O_1122,N_14296,N_13631);
and UO_1123 (O_1123,N_14390,N_14726);
nor UO_1124 (O_1124,N_13882,N_13804);
and UO_1125 (O_1125,N_13502,N_13986);
xnor UO_1126 (O_1126,N_13820,N_14477);
or UO_1127 (O_1127,N_13681,N_14589);
nor UO_1128 (O_1128,N_14208,N_14265);
nand UO_1129 (O_1129,N_13888,N_13972);
nand UO_1130 (O_1130,N_14958,N_14398);
or UO_1131 (O_1131,N_14766,N_14226);
and UO_1132 (O_1132,N_13596,N_13561);
or UO_1133 (O_1133,N_14327,N_14427);
nand UO_1134 (O_1134,N_14662,N_14369);
and UO_1135 (O_1135,N_14177,N_14789);
and UO_1136 (O_1136,N_14694,N_13931);
or UO_1137 (O_1137,N_14582,N_14380);
nor UO_1138 (O_1138,N_14785,N_14538);
xnor UO_1139 (O_1139,N_14690,N_14753);
nand UO_1140 (O_1140,N_14164,N_14954);
nand UO_1141 (O_1141,N_14399,N_14532);
or UO_1142 (O_1142,N_14696,N_13965);
and UO_1143 (O_1143,N_14134,N_14161);
or UO_1144 (O_1144,N_14820,N_13783);
or UO_1145 (O_1145,N_14090,N_14083);
nor UO_1146 (O_1146,N_14352,N_14112);
and UO_1147 (O_1147,N_14459,N_14195);
nor UO_1148 (O_1148,N_13677,N_13790);
and UO_1149 (O_1149,N_14273,N_13703);
and UO_1150 (O_1150,N_14592,N_13723);
xor UO_1151 (O_1151,N_14930,N_13887);
nand UO_1152 (O_1152,N_14899,N_13821);
xnor UO_1153 (O_1153,N_13933,N_13836);
nor UO_1154 (O_1154,N_14117,N_14267);
or UO_1155 (O_1155,N_14394,N_14302);
and UO_1156 (O_1156,N_14685,N_14768);
nand UO_1157 (O_1157,N_14918,N_13525);
nand UO_1158 (O_1158,N_14253,N_13500);
or UO_1159 (O_1159,N_14927,N_14173);
nand UO_1160 (O_1160,N_13640,N_14584);
xor UO_1161 (O_1161,N_14453,N_14693);
or UO_1162 (O_1162,N_13836,N_13502);
and UO_1163 (O_1163,N_14903,N_14387);
and UO_1164 (O_1164,N_13604,N_14267);
and UO_1165 (O_1165,N_13906,N_14904);
or UO_1166 (O_1166,N_14158,N_14532);
xor UO_1167 (O_1167,N_14458,N_14163);
and UO_1168 (O_1168,N_13515,N_14736);
or UO_1169 (O_1169,N_13619,N_14325);
xor UO_1170 (O_1170,N_14966,N_14853);
nor UO_1171 (O_1171,N_14492,N_13515);
and UO_1172 (O_1172,N_14785,N_14795);
nand UO_1173 (O_1173,N_14635,N_14770);
or UO_1174 (O_1174,N_14719,N_14802);
nor UO_1175 (O_1175,N_14658,N_14207);
xnor UO_1176 (O_1176,N_14158,N_14602);
nor UO_1177 (O_1177,N_13853,N_14387);
nand UO_1178 (O_1178,N_13562,N_14112);
nor UO_1179 (O_1179,N_13786,N_13767);
nand UO_1180 (O_1180,N_14923,N_14513);
xor UO_1181 (O_1181,N_14831,N_14469);
or UO_1182 (O_1182,N_14756,N_14816);
nor UO_1183 (O_1183,N_14184,N_14285);
xor UO_1184 (O_1184,N_14062,N_13741);
or UO_1185 (O_1185,N_14009,N_14749);
nand UO_1186 (O_1186,N_14091,N_14824);
nand UO_1187 (O_1187,N_14229,N_14685);
nor UO_1188 (O_1188,N_14414,N_14435);
and UO_1189 (O_1189,N_13962,N_14405);
nand UO_1190 (O_1190,N_14543,N_14561);
xor UO_1191 (O_1191,N_14871,N_13668);
xor UO_1192 (O_1192,N_14664,N_14504);
and UO_1193 (O_1193,N_14961,N_14758);
or UO_1194 (O_1194,N_13770,N_13809);
and UO_1195 (O_1195,N_14993,N_14918);
or UO_1196 (O_1196,N_13954,N_13969);
nand UO_1197 (O_1197,N_14146,N_14528);
and UO_1198 (O_1198,N_14971,N_13640);
xor UO_1199 (O_1199,N_14022,N_14413);
nor UO_1200 (O_1200,N_13930,N_14335);
nor UO_1201 (O_1201,N_13544,N_14395);
or UO_1202 (O_1202,N_13812,N_14129);
and UO_1203 (O_1203,N_14616,N_14763);
nand UO_1204 (O_1204,N_13775,N_14962);
nand UO_1205 (O_1205,N_14933,N_14644);
and UO_1206 (O_1206,N_14871,N_14141);
xnor UO_1207 (O_1207,N_13585,N_14401);
nand UO_1208 (O_1208,N_14927,N_13995);
xnor UO_1209 (O_1209,N_13862,N_14211);
or UO_1210 (O_1210,N_14898,N_14316);
nand UO_1211 (O_1211,N_14507,N_14158);
and UO_1212 (O_1212,N_14419,N_14908);
or UO_1213 (O_1213,N_13645,N_13725);
nand UO_1214 (O_1214,N_13732,N_14645);
nor UO_1215 (O_1215,N_14343,N_13766);
nor UO_1216 (O_1216,N_13909,N_13683);
nor UO_1217 (O_1217,N_14789,N_14864);
and UO_1218 (O_1218,N_14236,N_14912);
xor UO_1219 (O_1219,N_13594,N_13892);
nand UO_1220 (O_1220,N_14646,N_13811);
nand UO_1221 (O_1221,N_14252,N_14733);
nor UO_1222 (O_1222,N_13923,N_13638);
or UO_1223 (O_1223,N_13844,N_13654);
or UO_1224 (O_1224,N_14487,N_13613);
nand UO_1225 (O_1225,N_14962,N_14039);
nand UO_1226 (O_1226,N_13723,N_14672);
and UO_1227 (O_1227,N_14481,N_14456);
or UO_1228 (O_1228,N_13943,N_14194);
or UO_1229 (O_1229,N_14715,N_13631);
or UO_1230 (O_1230,N_14250,N_13614);
or UO_1231 (O_1231,N_14013,N_14984);
and UO_1232 (O_1232,N_14981,N_14896);
nor UO_1233 (O_1233,N_14010,N_13989);
and UO_1234 (O_1234,N_14799,N_14380);
or UO_1235 (O_1235,N_14167,N_14634);
or UO_1236 (O_1236,N_13940,N_13629);
nand UO_1237 (O_1237,N_13814,N_14386);
and UO_1238 (O_1238,N_13961,N_13504);
xor UO_1239 (O_1239,N_14415,N_14358);
nand UO_1240 (O_1240,N_14590,N_14009);
and UO_1241 (O_1241,N_13640,N_13631);
and UO_1242 (O_1242,N_14794,N_14192);
and UO_1243 (O_1243,N_14304,N_14826);
or UO_1244 (O_1244,N_14857,N_14993);
nor UO_1245 (O_1245,N_14283,N_13823);
xnor UO_1246 (O_1246,N_14910,N_14563);
nand UO_1247 (O_1247,N_14246,N_14951);
nor UO_1248 (O_1248,N_14800,N_14978);
and UO_1249 (O_1249,N_13523,N_14973);
nand UO_1250 (O_1250,N_13847,N_14993);
nor UO_1251 (O_1251,N_14683,N_14259);
xnor UO_1252 (O_1252,N_14710,N_14763);
or UO_1253 (O_1253,N_14457,N_13828);
nand UO_1254 (O_1254,N_14314,N_13697);
xor UO_1255 (O_1255,N_13876,N_13985);
and UO_1256 (O_1256,N_14257,N_14038);
and UO_1257 (O_1257,N_14474,N_13532);
and UO_1258 (O_1258,N_14034,N_14161);
or UO_1259 (O_1259,N_13949,N_14292);
nor UO_1260 (O_1260,N_13921,N_13749);
nor UO_1261 (O_1261,N_14716,N_14564);
nand UO_1262 (O_1262,N_14154,N_14443);
and UO_1263 (O_1263,N_13731,N_14754);
and UO_1264 (O_1264,N_13516,N_14685);
xor UO_1265 (O_1265,N_14799,N_14639);
nor UO_1266 (O_1266,N_14278,N_14873);
nor UO_1267 (O_1267,N_14481,N_14162);
nor UO_1268 (O_1268,N_14600,N_14812);
nor UO_1269 (O_1269,N_14798,N_13901);
xor UO_1270 (O_1270,N_13921,N_13931);
or UO_1271 (O_1271,N_14059,N_14337);
and UO_1272 (O_1272,N_14006,N_13552);
nand UO_1273 (O_1273,N_14295,N_13970);
and UO_1274 (O_1274,N_13997,N_14901);
or UO_1275 (O_1275,N_14351,N_13513);
nand UO_1276 (O_1276,N_14687,N_14389);
and UO_1277 (O_1277,N_14774,N_14467);
or UO_1278 (O_1278,N_13651,N_13751);
nand UO_1279 (O_1279,N_14784,N_14549);
xnor UO_1280 (O_1280,N_14046,N_14085);
xnor UO_1281 (O_1281,N_14016,N_14136);
nand UO_1282 (O_1282,N_14162,N_14134);
or UO_1283 (O_1283,N_13586,N_13985);
xnor UO_1284 (O_1284,N_14620,N_13997);
or UO_1285 (O_1285,N_14836,N_13903);
or UO_1286 (O_1286,N_14367,N_13858);
and UO_1287 (O_1287,N_13777,N_14910);
xor UO_1288 (O_1288,N_14420,N_14690);
xnor UO_1289 (O_1289,N_14472,N_14597);
nor UO_1290 (O_1290,N_14349,N_13791);
nand UO_1291 (O_1291,N_14392,N_13608);
or UO_1292 (O_1292,N_13774,N_14064);
or UO_1293 (O_1293,N_14169,N_14860);
and UO_1294 (O_1294,N_13888,N_13711);
nor UO_1295 (O_1295,N_14928,N_14940);
nor UO_1296 (O_1296,N_14735,N_13838);
nor UO_1297 (O_1297,N_14136,N_13777);
nand UO_1298 (O_1298,N_14176,N_13718);
nand UO_1299 (O_1299,N_14732,N_14775);
and UO_1300 (O_1300,N_14694,N_13979);
and UO_1301 (O_1301,N_13844,N_14504);
or UO_1302 (O_1302,N_14565,N_13987);
nor UO_1303 (O_1303,N_13932,N_13591);
nand UO_1304 (O_1304,N_14911,N_13820);
and UO_1305 (O_1305,N_13615,N_14843);
nand UO_1306 (O_1306,N_13534,N_14525);
and UO_1307 (O_1307,N_13851,N_14121);
nand UO_1308 (O_1308,N_14811,N_14393);
nor UO_1309 (O_1309,N_13516,N_13746);
nor UO_1310 (O_1310,N_14669,N_14065);
and UO_1311 (O_1311,N_14084,N_13956);
xnor UO_1312 (O_1312,N_14829,N_14124);
and UO_1313 (O_1313,N_14519,N_14720);
nor UO_1314 (O_1314,N_14079,N_14371);
xor UO_1315 (O_1315,N_13650,N_13576);
nand UO_1316 (O_1316,N_14163,N_13819);
and UO_1317 (O_1317,N_14477,N_14052);
xor UO_1318 (O_1318,N_14800,N_13771);
and UO_1319 (O_1319,N_14198,N_14763);
xor UO_1320 (O_1320,N_14138,N_14206);
nand UO_1321 (O_1321,N_13885,N_13746);
or UO_1322 (O_1322,N_14639,N_13574);
nand UO_1323 (O_1323,N_13928,N_14654);
nand UO_1324 (O_1324,N_14830,N_14645);
nor UO_1325 (O_1325,N_14969,N_14552);
and UO_1326 (O_1326,N_14597,N_13975);
or UO_1327 (O_1327,N_13812,N_14202);
or UO_1328 (O_1328,N_13950,N_14302);
and UO_1329 (O_1329,N_14830,N_14927);
nor UO_1330 (O_1330,N_14461,N_13956);
nand UO_1331 (O_1331,N_14385,N_13551);
nand UO_1332 (O_1332,N_13831,N_13869);
and UO_1333 (O_1333,N_14518,N_14735);
or UO_1334 (O_1334,N_13612,N_14750);
nand UO_1335 (O_1335,N_13908,N_14761);
xnor UO_1336 (O_1336,N_13853,N_14616);
or UO_1337 (O_1337,N_14981,N_14641);
xor UO_1338 (O_1338,N_13823,N_14721);
nand UO_1339 (O_1339,N_14671,N_13652);
nand UO_1340 (O_1340,N_14594,N_14556);
nor UO_1341 (O_1341,N_14536,N_14885);
nor UO_1342 (O_1342,N_14472,N_13716);
or UO_1343 (O_1343,N_14401,N_14147);
nand UO_1344 (O_1344,N_14190,N_14291);
xor UO_1345 (O_1345,N_14028,N_14368);
nand UO_1346 (O_1346,N_14482,N_14838);
or UO_1347 (O_1347,N_13569,N_14434);
nand UO_1348 (O_1348,N_14367,N_14187);
nand UO_1349 (O_1349,N_14981,N_14957);
and UO_1350 (O_1350,N_14800,N_13986);
nor UO_1351 (O_1351,N_14529,N_13654);
or UO_1352 (O_1352,N_14674,N_14564);
nor UO_1353 (O_1353,N_14640,N_14162);
nand UO_1354 (O_1354,N_13912,N_14188);
xnor UO_1355 (O_1355,N_13513,N_14999);
or UO_1356 (O_1356,N_13768,N_13773);
or UO_1357 (O_1357,N_13900,N_13642);
or UO_1358 (O_1358,N_14275,N_14463);
xor UO_1359 (O_1359,N_14093,N_13557);
or UO_1360 (O_1360,N_13540,N_14100);
nor UO_1361 (O_1361,N_13670,N_14583);
and UO_1362 (O_1362,N_14985,N_14370);
or UO_1363 (O_1363,N_14428,N_14251);
or UO_1364 (O_1364,N_14187,N_13744);
nand UO_1365 (O_1365,N_14046,N_13509);
xor UO_1366 (O_1366,N_13674,N_13728);
and UO_1367 (O_1367,N_14944,N_14316);
or UO_1368 (O_1368,N_14226,N_14335);
and UO_1369 (O_1369,N_14244,N_14956);
and UO_1370 (O_1370,N_14937,N_13854);
nand UO_1371 (O_1371,N_14850,N_14429);
nor UO_1372 (O_1372,N_14499,N_14817);
xnor UO_1373 (O_1373,N_14550,N_14202);
nor UO_1374 (O_1374,N_13722,N_13810);
and UO_1375 (O_1375,N_14640,N_14852);
xnor UO_1376 (O_1376,N_14302,N_14657);
nor UO_1377 (O_1377,N_14594,N_14779);
nor UO_1378 (O_1378,N_14384,N_14058);
nor UO_1379 (O_1379,N_13780,N_14061);
or UO_1380 (O_1380,N_13625,N_13692);
xor UO_1381 (O_1381,N_14491,N_14574);
nand UO_1382 (O_1382,N_13577,N_14690);
or UO_1383 (O_1383,N_14723,N_14389);
nor UO_1384 (O_1384,N_13792,N_14756);
or UO_1385 (O_1385,N_13752,N_14748);
nand UO_1386 (O_1386,N_14566,N_13976);
nor UO_1387 (O_1387,N_13801,N_14896);
xor UO_1388 (O_1388,N_13838,N_13966);
and UO_1389 (O_1389,N_14229,N_14672);
nand UO_1390 (O_1390,N_13925,N_13812);
and UO_1391 (O_1391,N_14679,N_14873);
nor UO_1392 (O_1392,N_14336,N_14282);
nand UO_1393 (O_1393,N_14397,N_14726);
nand UO_1394 (O_1394,N_14327,N_14784);
xnor UO_1395 (O_1395,N_14825,N_13947);
nor UO_1396 (O_1396,N_14669,N_14517);
and UO_1397 (O_1397,N_13509,N_14338);
nor UO_1398 (O_1398,N_14633,N_14758);
xnor UO_1399 (O_1399,N_13732,N_14469);
nor UO_1400 (O_1400,N_14165,N_13793);
nand UO_1401 (O_1401,N_13640,N_13735);
nand UO_1402 (O_1402,N_13520,N_14601);
nand UO_1403 (O_1403,N_14121,N_13893);
nand UO_1404 (O_1404,N_14644,N_14245);
nor UO_1405 (O_1405,N_13762,N_13987);
nor UO_1406 (O_1406,N_14562,N_13977);
or UO_1407 (O_1407,N_14849,N_14930);
or UO_1408 (O_1408,N_14711,N_14725);
xnor UO_1409 (O_1409,N_13958,N_14140);
and UO_1410 (O_1410,N_14945,N_14447);
or UO_1411 (O_1411,N_14883,N_13540);
or UO_1412 (O_1412,N_13552,N_14105);
or UO_1413 (O_1413,N_13625,N_13895);
nand UO_1414 (O_1414,N_13502,N_14858);
or UO_1415 (O_1415,N_13805,N_14188);
and UO_1416 (O_1416,N_13797,N_14856);
nor UO_1417 (O_1417,N_13505,N_14141);
nand UO_1418 (O_1418,N_14472,N_14198);
and UO_1419 (O_1419,N_14500,N_14774);
nor UO_1420 (O_1420,N_14958,N_14862);
nand UO_1421 (O_1421,N_13513,N_14520);
xnor UO_1422 (O_1422,N_14932,N_13671);
nor UO_1423 (O_1423,N_14142,N_13795);
nor UO_1424 (O_1424,N_14364,N_14825);
nor UO_1425 (O_1425,N_14012,N_13862);
xor UO_1426 (O_1426,N_13638,N_13937);
xnor UO_1427 (O_1427,N_13826,N_14877);
and UO_1428 (O_1428,N_13580,N_13588);
nor UO_1429 (O_1429,N_14356,N_13899);
nor UO_1430 (O_1430,N_14105,N_14594);
xor UO_1431 (O_1431,N_14945,N_14987);
and UO_1432 (O_1432,N_13620,N_14604);
and UO_1433 (O_1433,N_13792,N_13606);
or UO_1434 (O_1434,N_14887,N_14192);
or UO_1435 (O_1435,N_13831,N_14726);
and UO_1436 (O_1436,N_13598,N_14585);
nor UO_1437 (O_1437,N_14218,N_13992);
and UO_1438 (O_1438,N_13850,N_13664);
and UO_1439 (O_1439,N_14729,N_14679);
or UO_1440 (O_1440,N_14244,N_13938);
and UO_1441 (O_1441,N_13602,N_14875);
and UO_1442 (O_1442,N_14927,N_14599);
nand UO_1443 (O_1443,N_14952,N_14812);
and UO_1444 (O_1444,N_13758,N_14057);
and UO_1445 (O_1445,N_13871,N_13594);
nand UO_1446 (O_1446,N_14509,N_14337);
nor UO_1447 (O_1447,N_14623,N_14336);
xnor UO_1448 (O_1448,N_14267,N_13675);
nor UO_1449 (O_1449,N_14143,N_13986);
nor UO_1450 (O_1450,N_14712,N_13505);
xnor UO_1451 (O_1451,N_14219,N_14965);
or UO_1452 (O_1452,N_14199,N_14194);
nor UO_1453 (O_1453,N_13787,N_13600);
xor UO_1454 (O_1454,N_13886,N_14833);
xnor UO_1455 (O_1455,N_14254,N_14074);
or UO_1456 (O_1456,N_14891,N_14728);
nand UO_1457 (O_1457,N_13633,N_14142);
nor UO_1458 (O_1458,N_13797,N_13840);
and UO_1459 (O_1459,N_14519,N_13658);
and UO_1460 (O_1460,N_14299,N_14389);
xor UO_1461 (O_1461,N_14813,N_14250);
xnor UO_1462 (O_1462,N_13554,N_13676);
nor UO_1463 (O_1463,N_14261,N_13623);
or UO_1464 (O_1464,N_14442,N_14430);
and UO_1465 (O_1465,N_13502,N_14150);
xor UO_1466 (O_1466,N_14339,N_14865);
and UO_1467 (O_1467,N_13661,N_14468);
and UO_1468 (O_1468,N_14846,N_13890);
xnor UO_1469 (O_1469,N_13936,N_13697);
or UO_1470 (O_1470,N_14021,N_13683);
nand UO_1471 (O_1471,N_13690,N_14966);
and UO_1472 (O_1472,N_14976,N_14937);
xnor UO_1473 (O_1473,N_13820,N_13823);
and UO_1474 (O_1474,N_14865,N_14193);
nor UO_1475 (O_1475,N_14971,N_14940);
nor UO_1476 (O_1476,N_14425,N_14877);
xnor UO_1477 (O_1477,N_14233,N_14977);
or UO_1478 (O_1478,N_14775,N_13602);
nor UO_1479 (O_1479,N_14882,N_14600);
nand UO_1480 (O_1480,N_14510,N_14432);
xnor UO_1481 (O_1481,N_14855,N_14093);
xor UO_1482 (O_1482,N_14200,N_14044);
nand UO_1483 (O_1483,N_14672,N_14986);
and UO_1484 (O_1484,N_14922,N_14410);
nand UO_1485 (O_1485,N_14150,N_14811);
nand UO_1486 (O_1486,N_13575,N_14397);
xnor UO_1487 (O_1487,N_14758,N_13940);
and UO_1488 (O_1488,N_14781,N_13926);
or UO_1489 (O_1489,N_14279,N_14285);
and UO_1490 (O_1490,N_14638,N_14227);
xnor UO_1491 (O_1491,N_13710,N_14261);
nand UO_1492 (O_1492,N_13615,N_13957);
or UO_1493 (O_1493,N_14058,N_14031);
and UO_1494 (O_1494,N_13821,N_13526);
and UO_1495 (O_1495,N_14537,N_14417);
and UO_1496 (O_1496,N_14502,N_14943);
nor UO_1497 (O_1497,N_13551,N_13594);
and UO_1498 (O_1498,N_14153,N_13775);
and UO_1499 (O_1499,N_13517,N_14908);
and UO_1500 (O_1500,N_14196,N_14577);
nand UO_1501 (O_1501,N_13916,N_14097);
nor UO_1502 (O_1502,N_13809,N_13715);
nand UO_1503 (O_1503,N_14661,N_13963);
xnor UO_1504 (O_1504,N_14467,N_14306);
nor UO_1505 (O_1505,N_14444,N_14956);
nand UO_1506 (O_1506,N_13984,N_14834);
nand UO_1507 (O_1507,N_13747,N_14296);
nand UO_1508 (O_1508,N_14505,N_14066);
or UO_1509 (O_1509,N_14204,N_14239);
and UO_1510 (O_1510,N_14853,N_14017);
and UO_1511 (O_1511,N_14887,N_14112);
and UO_1512 (O_1512,N_14898,N_14862);
and UO_1513 (O_1513,N_13841,N_13623);
nor UO_1514 (O_1514,N_13978,N_13725);
nor UO_1515 (O_1515,N_14787,N_14104);
and UO_1516 (O_1516,N_14311,N_14762);
nor UO_1517 (O_1517,N_14025,N_14361);
xor UO_1518 (O_1518,N_13800,N_13668);
nand UO_1519 (O_1519,N_13791,N_13688);
xor UO_1520 (O_1520,N_14897,N_14338);
nor UO_1521 (O_1521,N_14229,N_14994);
or UO_1522 (O_1522,N_13752,N_13922);
or UO_1523 (O_1523,N_14808,N_14873);
nor UO_1524 (O_1524,N_13995,N_14898);
nand UO_1525 (O_1525,N_13552,N_14862);
xor UO_1526 (O_1526,N_13917,N_13517);
nand UO_1527 (O_1527,N_13962,N_14141);
nand UO_1528 (O_1528,N_13866,N_13657);
or UO_1529 (O_1529,N_14168,N_14603);
or UO_1530 (O_1530,N_14639,N_14985);
and UO_1531 (O_1531,N_14877,N_14538);
and UO_1532 (O_1532,N_13591,N_14268);
nor UO_1533 (O_1533,N_13629,N_13905);
or UO_1534 (O_1534,N_14613,N_13722);
and UO_1535 (O_1535,N_14106,N_14833);
xnor UO_1536 (O_1536,N_14639,N_13770);
nand UO_1537 (O_1537,N_13985,N_14347);
xnor UO_1538 (O_1538,N_13690,N_14097);
and UO_1539 (O_1539,N_14814,N_13721);
xnor UO_1540 (O_1540,N_13994,N_13657);
nand UO_1541 (O_1541,N_14302,N_14188);
nor UO_1542 (O_1542,N_13808,N_14297);
xnor UO_1543 (O_1543,N_14514,N_14730);
xor UO_1544 (O_1544,N_14654,N_14831);
nand UO_1545 (O_1545,N_14634,N_14917);
xnor UO_1546 (O_1546,N_14400,N_13588);
xor UO_1547 (O_1547,N_14954,N_14607);
nand UO_1548 (O_1548,N_14877,N_14907);
nand UO_1549 (O_1549,N_14631,N_14980);
nor UO_1550 (O_1550,N_14352,N_14223);
nand UO_1551 (O_1551,N_14960,N_13593);
or UO_1552 (O_1552,N_13919,N_13527);
nand UO_1553 (O_1553,N_14342,N_13527);
xnor UO_1554 (O_1554,N_14500,N_13903);
nor UO_1555 (O_1555,N_14682,N_13955);
and UO_1556 (O_1556,N_14471,N_13500);
nand UO_1557 (O_1557,N_14731,N_14958);
xnor UO_1558 (O_1558,N_14724,N_14893);
nor UO_1559 (O_1559,N_14496,N_13919);
xnor UO_1560 (O_1560,N_14680,N_14590);
nand UO_1561 (O_1561,N_14811,N_14034);
nand UO_1562 (O_1562,N_13686,N_14699);
nand UO_1563 (O_1563,N_13968,N_14048);
or UO_1564 (O_1564,N_14642,N_14055);
nor UO_1565 (O_1565,N_14078,N_13876);
or UO_1566 (O_1566,N_14761,N_14391);
xor UO_1567 (O_1567,N_13708,N_14130);
nand UO_1568 (O_1568,N_14385,N_13513);
or UO_1569 (O_1569,N_14093,N_14110);
xnor UO_1570 (O_1570,N_14216,N_14845);
and UO_1571 (O_1571,N_13584,N_14505);
and UO_1572 (O_1572,N_14914,N_13675);
or UO_1573 (O_1573,N_14859,N_13584);
or UO_1574 (O_1574,N_14302,N_13671);
and UO_1575 (O_1575,N_14823,N_14118);
and UO_1576 (O_1576,N_14119,N_13706);
or UO_1577 (O_1577,N_14215,N_14009);
or UO_1578 (O_1578,N_13871,N_14444);
nand UO_1579 (O_1579,N_14811,N_14323);
nor UO_1580 (O_1580,N_14039,N_13960);
xnor UO_1581 (O_1581,N_14891,N_14997);
and UO_1582 (O_1582,N_14830,N_13858);
xor UO_1583 (O_1583,N_14546,N_14242);
and UO_1584 (O_1584,N_13567,N_13696);
and UO_1585 (O_1585,N_13835,N_14817);
and UO_1586 (O_1586,N_13807,N_14256);
nor UO_1587 (O_1587,N_13567,N_14671);
or UO_1588 (O_1588,N_14508,N_13611);
and UO_1589 (O_1589,N_14155,N_14779);
and UO_1590 (O_1590,N_14475,N_14564);
nor UO_1591 (O_1591,N_14469,N_14771);
nor UO_1592 (O_1592,N_14824,N_14601);
and UO_1593 (O_1593,N_14456,N_14272);
and UO_1594 (O_1594,N_14887,N_14191);
xnor UO_1595 (O_1595,N_13701,N_14722);
xnor UO_1596 (O_1596,N_13970,N_13811);
xnor UO_1597 (O_1597,N_13797,N_14148);
and UO_1598 (O_1598,N_14119,N_14240);
or UO_1599 (O_1599,N_14497,N_14288);
nand UO_1600 (O_1600,N_14320,N_14936);
xnor UO_1601 (O_1601,N_14559,N_14579);
and UO_1602 (O_1602,N_13522,N_13702);
or UO_1603 (O_1603,N_14539,N_13880);
nand UO_1604 (O_1604,N_13617,N_14049);
nand UO_1605 (O_1605,N_13796,N_13808);
xnor UO_1606 (O_1606,N_13538,N_13809);
nand UO_1607 (O_1607,N_14123,N_14106);
xnor UO_1608 (O_1608,N_13857,N_13775);
nor UO_1609 (O_1609,N_14516,N_14193);
nand UO_1610 (O_1610,N_13903,N_13827);
or UO_1611 (O_1611,N_14557,N_14502);
and UO_1612 (O_1612,N_14012,N_14644);
nand UO_1613 (O_1613,N_14917,N_14717);
or UO_1614 (O_1614,N_14216,N_14950);
nand UO_1615 (O_1615,N_13608,N_14189);
and UO_1616 (O_1616,N_14675,N_14319);
and UO_1617 (O_1617,N_14165,N_14792);
or UO_1618 (O_1618,N_13815,N_14558);
or UO_1619 (O_1619,N_14921,N_14286);
xnor UO_1620 (O_1620,N_13695,N_14186);
nand UO_1621 (O_1621,N_14900,N_13907);
nor UO_1622 (O_1622,N_14295,N_14292);
xor UO_1623 (O_1623,N_14213,N_13834);
or UO_1624 (O_1624,N_13545,N_14389);
xor UO_1625 (O_1625,N_13818,N_14311);
nor UO_1626 (O_1626,N_14612,N_13989);
or UO_1627 (O_1627,N_13679,N_14982);
xnor UO_1628 (O_1628,N_14881,N_14008);
or UO_1629 (O_1629,N_14378,N_14244);
nor UO_1630 (O_1630,N_14534,N_14886);
and UO_1631 (O_1631,N_14381,N_14280);
nor UO_1632 (O_1632,N_14880,N_14893);
or UO_1633 (O_1633,N_14386,N_14795);
xnor UO_1634 (O_1634,N_14613,N_13862);
or UO_1635 (O_1635,N_13587,N_13817);
and UO_1636 (O_1636,N_13776,N_13718);
and UO_1637 (O_1637,N_13530,N_13608);
nand UO_1638 (O_1638,N_13912,N_14293);
xor UO_1639 (O_1639,N_14388,N_14882);
and UO_1640 (O_1640,N_14910,N_14386);
xor UO_1641 (O_1641,N_14904,N_13835);
or UO_1642 (O_1642,N_14793,N_13502);
and UO_1643 (O_1643,N_13516,N_13558);
xor UO_1644 (O_1644,N_14641,N_14953);
and UO_1645 (O_1645,N_14209,N_14572);
xnor UO_1646 (O_1646,N_14286,N_13738);
and UO_1647 (O_1647,N_13684,N_14571);
nand UO_1648 (O_1648,N_14822,N_13864);
or UO_1649 (O_1649,N_14760,N_13769);
nand UO_1650 (O_1650,N_14490,N_14888);
and UO_1651 (O_1651,N_14431,N_14928);
xnor UO_1652 (O_1652,N_13833,N_14558);
xor UO_1653 (O_1653,N_14367,N_13879);
xnor UO_1654 (O_1654,N_14188,N_14666);
and UO_1655 (O_1655,N_14258,N_14220);
and UO_1656 (O_1656,N_13618,N_14531);
and UO_1657 (O_1657,N_14463,N_14504);
nand UO_1658 (O_1658,N_14762,N_14540);
and UO_1659 (O_1659,N_14189,N_14344);
nand UO_1660 (O_1660,N_13863,N_14498);
and UO_1661 (O_1661,N_14271,N_13503);
and UO_1662 (O_1662,N_14837,N_14281);
xnor UO_1663 (O_1663,N_13763,N_13676);
xor UO_1664 (O_1664,N_14499,N_14289);
and UO_1665 (O_1665,N_13590,N_14605);
and UO_1666 (O_1666,N_14034,N_14211);
and UO_1667 (O_1667,N_14718,N_13887);
xor UO_1668 (O_1668,N_14390,N_13890);
nand UO_1669 (O_1669,N_14453,N_13991);
xor UO_1670 (O_1670,N_13513,N_14164);
nand UO_1671 (O_1671,N_14241,N_13932);
and UO_1672 (O_1672,N_14841,N_13666);
and UO_1673 (O_1673,N_14602,N_13922);
nor UO_1674 (O_1674,N_14897,N_13545);
nor UO_1675 (O_1675,N_14144,N_14612);
xnor UO_1676 (O_1676,N_13973,N_14194);
and UO_1677 (O_1677,N_14142,N_14054);
and UO_1678 (O_1678,N_14985,N_14608);
xor UO_1679 (O_1679,N_14085,N_14397);
and UO_1680 (O_1680,N_14318,N_13757);
or UO_1681 (O_1681,N_13705,N_13834);
or UO_1682 (O_1682,N_14815,N_14827);
nand UO_1683 (O_1683,N_14341,N_14438);
xnor UO_1684 (O_1684,N_14153,N_14564);
xor UO_1685 (O_1685,N_13698,N_14693);
and UO_1686 (O_1686,N_13703,N_14834);
or UO_1687 (O_1687,N_14155,N_14141);
or UO_1688 (O_1688,N_13760,N_13659);
and UO_1689 (O_1689,N_14454,N_13760);
or UO_1690 (O_1690,N_13833,N_13818);
and UO_1691 (O_1691,N_14280,N_14423);
nand UO_1692 (O_1692,N_14267,N_13658);
and UO_1693 (O_1693,N_14313,N_13733);
or UO_1694 (O_1694,N_14561,N_14184);
and UO_1695 (O_1695,N_14478,N_14925);
nor UO_1696 (O_1696,N_13581,N_14182);
nand UO_1697 (O_1697,N_13873,N_14947);
or UO_1698 (O_1698,N_14126,N_14774);
xor UO_1699 (O_1699,N_14242,N_14232);
nand UO_1700 (O_1700,N_14333,N_14323);
nand UO_1701 (O_1701,N_14433,N_14591);
and UO_1702 (O_1702,N_14247,N_13999);
nand UO_1703 (O_1703,N_13827,N_13549);
nand UO_1704 (O_1704,N_13828,N_14521);
nor UO_1705 (O_1705,N_14357,N_14585);
xor UO_1706 (O_1706,N_13837,N_14091);
and UO_1707 (O_1707,N_14924,N_13657);
and UO_1708 (O_1708,N_13542,N_13857);
or UO_1709 (O_1709,N_13882,N_14454);
nand UO_1710 (O_1710,N_14838,N_13865);
nor UO_1711 (O_1711,N_14036,N_14741);
nor UO_1712 (O_1712,N_14314,N_14867);
nor UO_1713 (O_1713,N_14120,N_13746);
or UO_1714 (O_1714,N_14018,N_14041);
xnor UO_1715 (O_1715,N_14450,N_14781);
and UO_1716 (O_1716,N_14957,N_14051);
or UO_1717 (O_1717,N_14876,N_14558);
or UO_1718 (O_1718,N_13798,N_13921);
nand UO_1719 (O_1719,N_14859,N_14353);
nand UO_1720 (O_1720,N_14442,N_14408);
xnor UO_1721 (O_1721,N_14760,N_13558);
nand UO_1722 (O_1722,N_14135,N_14701);
or UO_1723 (O_1723,N_14756,N_14296);
nor UO_1724 (O_1724,N_14317,N_14658);
and UO_1725 (O_1725,N_13504,N_14712);
or UO_1726 (O_1726,N_13658,N_14713);
xor UO_1727 (O_1727,N_14128,N_13558);
nor UO_1728 (O_1728,N_14421,N_13946);
nand UO_1729 (O_1729,N_14269,N_13822);
and UO_1730 (O_1730,N_13820,N_14424);
xor UO_1731 (O_1731,N_14226,N_14660);
nand UO_1732 (O_1732,N_13823,N_13642);
nand UO_1733 (O_1733,N_13702,N_13909);
nand UO_1734 (O_1734,N_13736,N_14633);
nor UO_1735 (O_1735,N_13835,N_13741);
nand UO_1736 (O_1736,N_14612,N_14615);
xor UO_1737 (O_1737,N_13579,N_14559);
or UO_1738 (O_1738,N_14564,N_14879);
xnor UO_1739 (O_1739,N_14462,N_14486);
and UO_1740 (O_1740,N_14565,N_14177);
nor UO_1741 (O_1741,N_14376,N_13550);
and UO_1742 (O_1742,N_14761,N_13719);
xor UO_1743 (O_1743,N_14842,N_13704);
xnor UO_1744 (O_1744,N_14590,N_14242);
xor UO_1745 (O_1745,N_13989,N_14518);
nor UO_1746 (O_1746,N_14041,N_14677);
or UO_1747 (O_1747,N_13548,N_14019);
nand UO_1748 (O_1748,N_14593,N_14591);
nand UO_1749 (O_1749,N_14556,N_13976);
or UO_1750 (O_1750,N_14458,N_13555);
or UO_1751 (O_1751,N_14932,N_13924);
nor UO_1752 (O_1752,N_13707,N_14690);
or UO_1753 (O_1753,N_14128,N_13571);
or UO_1754 (O_1754,N_13788,N_14641);
and UO_1755 (O_1755,N_13959,N_14665);
and UO_1756 (O_1756,N_13902,N_14735);
nor UO_1757 (O_1757,N_13850,N_14981);
nand UO_1758 (O_1758,N_14475,N_14610);
and UO_1759 (O_1759,N_13748,N_14164);
nor UO_1760 (O_1760,N_13825,N_13614);
and UO_1761 (O_1761,N_14874,N_13557);
nor UO_1762 (O_1762,N_14036,N_14825);
or UO_1763 (O_1763,N_13745,N_13510);
and UO_1764 (O_1764,N_14774,N_14492);
and UO_1765 (O_1765,N_13605,N_13932);
or UO_1766 (O_1766,N_14075,N_14389);
nand UO_1767 (O_1767,N_13518,N_14446);
nor UO_1768 (O_1768,N_14443,N_14289);
nor UO_1769 (O_1769,N_14940,N_13759);
nor UO_1770 (O_1770,N_13550,N_14268);
and UO_1771 (O_1771,N_13500,N_14703);
or UO_1772 (O_1772,N_13511,N_13851);
and UO_1773 (O_1773,N_14354,N_14998);
nor UO_1774 (O_1774,N_13940,N_13703);
nor UO_1775 (O_1775,N_14255,N_13593);
nor UO_1776 (O_1776,N_14443,N_14231);
xnor UO_1777 (O_1777,N_13814,N_13986);
nand UO_1778 (O_1778,N_14678,N_14884);
nand UO_1779 (O_1779,N_14194,N_13622);
and UO_1780 (O_1780,N_13917,N_14673);
nor UO_1781 (O_1781,N_14971,N_14932);
or UO_1782 (O_1782,N_14248,N_14878);
and UO_1783 (O_1783,N_13532,N_14421);
nor UO_1784 (O_1784,N_14635,N_14325);
and UO_1785 (O_1785,N_14073,N_14671);
xor UO_1786 (O_1786,N_14040,N_14191);
or UO_1787 (O_1787,N_14502,N_14727);
xor UO_1788 (O_1788,N_13930,N_14809);
nor UO_1789 (O_1789,N_13537,N_13877);
xnor UO_1790 (O_1790,N_14837,N_14345);
and UO_1791 (O_1791,N_14231,N_13687);
nor UO_1792 (O_1792,N_13725,N_14338);
nand UO_1793 (O_1793,N_13680,N_14170);
and UO_1794 (O_1794,N_14833,N_13871);
xor UO_1795 (O_1795,N_13969,N_13667);
or UO_1796 (O_1796,N_14841,N_14703);
nor UO_1797 (O_1797,N_14561,N_14009);
or UO_1798 (O_1798,N_14284,N_14594);
nor UO_1799 (O_1799,N_14188,N_13632);
nand UO_1800 (O_1800,N_14141,N_13691);
or UO_1801 (O_1801,N_14535,N_14925);
nor UO_1802 (O_1802,N_13990,N_14512);
and UO_1803 (O_1803,N_13772,N_13890);
nor UO_1804 (O_1804,N_14014,N_14006);
or UO_1805 (O_1805,N_13603,N_14308);
nor UO_1806 (O_1806,N_14393,N_13547);
nand UO_1807 (O_1807,N_13561,N_14282);
and UO_1808 (O_1808,N_13514,N_13792);
nand UO_1809 (O_1809,N_14471,N_13715);
xnor UO_1810 (O_1810,N_13787,N_14254);
nand UO_1811 (O_1811,N_13550,N_13775);
and UO_1812 (O_1812,N_14257,N_13726);
and UO_1813 (O_1813,N_14102,N_13708);
xor UO_1814 (O_1814,N_14496,N_14104);
nor UO_1815 (O_1815,N_13781,N_14209);
nor UO_1816 (O_1816,N_14809,N_14034);
or UO_1817 (O_1817,N_13616,N_14042);
and UO_1818 (O_1818,N_14664,N_13856);
or UO_1819 (O_1819,N_14561,N_14842);
and UO_1820 (O_1820,N_14881,N_14333);
nand UO_1821 (O_1821,N_13807,N_14722);
nand UO_1822 (O_1822,N_13742,N_13840);
or UO_1823 (O_1823,N_14903,N_14221);
nor UO_1824 (O_1824,N_13866,N_14665);
and UO_1825 (O_1825,N_13932,N_14340);
xnor UO_1826 (O_1826,N_13749,N_13677);
xor UO_1827 (O_1827,N_14807,N_13996);
xor UO_1828 (O_1828,N_14456,N_14222);
xor UO_1829 (O_1829,N_14389,N_14944);
and UO_1830 (O_1830,N_14617,N_14431);
xor UO_1831 (O_1831,N_13617,N_13949);
or UO_1832 (O_1832,N_13882,N_14348);
and UO_1833 (O_1833,N_13695,N_13748);
nand UO_1834 (O_1834,N_14473,N_13993);
and UO_1835 (O_1835,N_14819,N_14383);
and UO_1836 (O_1836,N_14439,N_13861);
xor UO_1837 (O_1837,N_13826,N_14413);
and UO_1838 (O_1838,N_13670,N_14821);
xnor UO_1839 (O_1839,N_14786,N_14332);
and UO_1840 (O_1840,N_14660,N_13939);
nand UO_1841 (O_1841,N_13594,N_13885);
nor UO_1842 (O_1842,N_14930,N_14346);
xnor UO_1843 (O_1843,N_14328,N_14737);
or UO_1844 (O_1844,N_14997,N_14974);
or UO_1845 (O_1845,N_13762,N_14968);
and UO_1846 (O_1846,N_14401,N_14886);
or UO_1847 (O_1847,N_14797,N_14347);
or UO_1848 (O_1848,N_14641,N_14571);
or UO_1849 (O_1849,N_13658,N_14685);
xnor UO_1850 (O_1850,N_13571,N_13620);
nand UO_1851 (O_1851,N_13967,N_13904);
nand UO_1852 (O_1852,N_14797,N_14424);
nor UO_1853 (O_1853,N_14049,N_14948);
nand UO_1854 (O_1854,N_14761,N_14044);
nor UO_1855 (O_1855,N_13728,N_14365);
xnor UO_1856 (O_1856,N_14691,N_14946);
nand UO_1857 (O_1857,N_13514,N_14065);
nor UO_1858 (O_1858,N_14898,N_14866);
or UO_1859 (O_1859,N_14666,N_14593);
nand UO_1860 (O_1860,N_13546,N_14181);
nand UO_1861 (O_1861,N_14067,N_13533);
and UO_1862 (O_1862,N_14996,N_14344);
and UO_1863 (O_1863,N_13941,N_14522);
or UO_1864 (O_1864,N_14300,N_14171);
xor UO_1865 (O_1865,N_13960,N_14521);
and UO_1866 (O_1866,N_14123,N_14384);
xor UO_1867 (O_1867,N_14904,N_13967);
nor UO_1868 (O_1868,N_14528,N_14398);
or UO_1869 (O_1869,N_13762,N_13986);
nor UO_1870 (O_1870,N_13972,N_14469);
xor UO_1871 (O_1871,N_13912,N_14395);
xor UO_1872 (O_1872,N_14007,N_13751);
nor UO_1873 (O_1873,N_14623,N_14595);
and UO_1874 (O_1874,N_14628,N_14215);
xnor UO_1875 (O_1875,N_14113,N_14546);
nor UO_1876 (O_1876,N_14514,N_14328);
and UO_1877 (O_1877,N_13747,N_14241);
or UO_1878 (O_1878,N_14409,N_14056);
or UO_1879 (O_1879,N_13913,N_14241);
and UO_1880 (O_1880,N_13678,N_14713);
nand UO_1881 (O_1881,N_14429,N_14297);
nand UO_1882 (O_1882,N_13761,N_13752);
and UO_1883 (O_1883,N_14700,N_13571);
or UO_1884 (O_1884,N_13913,N_14103);
or UO_1885 (O_1885,N_14736,N_14653);
and UO_1886 (O_1886,N_13514,N_14728);
and UO_1887 (O_1887,N_13781,N_14657);
or UO_1888 (O_1888,N_14755,N_14116);
or UO_1889 (O_1889,N_13561,N_14117);
nor UO_1890 (O_1890,N_14823,N_13607);
or UO_1891 (O_1891,N_14442,N_13758);
xnor UO_1892 (O_1892,N_14090,N_13870);
and UO_1893 (O_1893,N_13563,N_14305);
and UO_1894 (O_1894,N_14397,N_14037);
nand UO_1895 (O_1895,N_13742,N_13810);
and UO_1896 (O_1896,N_14105,N_14458);
nand UO_1897 (O_1897,N_13724,N_14017);
and UO_1898 (O_1898,N_13736,N_13572);
nor UO_1899 (O_1899,N_14235,N_14895);
nand UO_1900 (O_1900,N_13800,N_13536);
xnor UO_1901 (O_1901,N_14026,N_13813);
or UO_1902 (O_1902,N_14748,N_14083);
xor UO_1903 (O_1903,N_14556,N_13876);
or UO_1904 (O_1904,N_13813,N_13742);
xnor UO_1905 (O_1905,N_14414,N_14522);
nor UO_1906 (O_1906,N_14765,N_14479);
nand UO_1907 (O_1907,N_14206,N_14982);
or UO_1908 (O_1908,N_14466,N_14897);
nand UO_1909 (O_1909,N_13933,N_14634);
nor UO_1910 (O_1910,N_14391,N_14335);
and UO_1911 (O_1911,N_14333,N_14041);
nor UO_1912 (O_1912,N_14378,N_13829);
xor UO_1913 (O_1913,N_13931,N_14468);
nand UO_1914 (O_1914,N_13933,N_13884);
xnor UO_1915 (O_1915,N_13807,N_13604);
nor UO_1916 (O_1916,N_13858,N_13805);
nor UO_1917 (O_1917,N_13856,N_14958);
and UO_1918 (O_1918,N_14007,N_14672);
xnor UO_1919 (O_1919,N_14315,N_14020);
or UO_1920 (O_1920,N_14005,N_14144);
xnor UO_1921 (O_1921,N_13944,N_13745);
nor UO_1922 (O_1922,N_14689,N_14766);
or UO_1923 (O_1923,N_13511,N_14827);
and UO_1924 (O_1924,N_14009,N_14068);
nand UO_1925 (O_1925,N_14571,N_14506);
or UO_1926 (O_1926,N_13736,N_14173);
xnor UO_1927 (O_1927,N_14664,N_14349);
nand UO_1928 (O_1928,N_13825,N_14409);
nand UO_1929 (O_1929,N_14613,N_14538);
or UO_1930 (O_1930,N_13885,N_14281);
nor UO_1931 (O_1931,N_14283,N_14927);
nand UO_1932 (O_1932,N_13610,N_14833);
nand UO_1933 (O_1933,N_14102,N_14964);
and UO_1934 (O_1934,N_13648,N_14233);
nand UO_1935 (O_1935,N_14963,N_14063);
xnor UO_1936 (O_1936,N_14144,N_13788);
and UO_1937 (O_1937,N_14661,N_14814);
xor UO_1938 (O_1938,N_13655,N_13583);
nor UO_1939 (O_1939,N_14224,N_14092);
or UO_1940 (O_1940,N_13985,N_14651);
or UO_1941 (O_1941,N_13703,N_13773);
nor UO_1942 (O_1942,N_13852,N_13523);
or UO_1943 (O_1943,N_14006,N_13967);
xnor UO_1944 (O_1944,N_14422,N_14489);
and UO_1945 (O_1945,N_13585,N_14975);
nor UO_1946 (O_1946,N_13622,N_14074);
nand UO_1947 (O_1947,N_13880,N_14489);
or UO_1948 (O_1948,N_13515,N_13984);
nand UO_1949 (O_1949,N_14122,N_13801);
nand UO_1950 (O_1950,N_14976,N_13503);
or UO_1951 (O_1951,N_14968,N_13543);
nand UO_1952 (O_1952,N_13569,N_13602);
or UO_1953 (O_1953,N_13835,N_14623);
nand UO_1954 (O_1954,N_14517,N_14846);
nor UO_1955 (O_1955,N_14001,N_13638);
nand UO_1956 (O_1956,N_14127,N_14795);
and UO_1957 (O_1957,N_14539,N_13500);
nor UO_1958 (O_1958,N_13808,N_14472);
xnor UO_1959 (O_1959,N_14066,N_13971);
xnor UO_1960 (O_1960,N_13655,N_14924);
xor UO_1961 (O_1961,N_13857,N_14154);
or UO_1962 (O_1962,N_13937,N_14338);
or UO_1963 (O_1963,N_13616,N_13651);
xnor UO_1964 (O_1964,N_14699,N_14201);
nand UO_1965 (O_1965,N_14927,N_14250);
nor UO_1966 (O_1966,N_14514,N_13598);
or UO_1967 (O_1967,N_14952,N_14029);
nand UO_1968 (O_1968,N_14941,N_14398);
nand UO_1969 (O_1969,N_14876,N_13712);
or UO_1970 (O_1970,N_13622,N_14011);
and UO_1971 (O_1971,N_13560,N_14826);
and UO_1972 (O_1972,N_13552,N_13640);
xnor UO_1973 (O_1973,N_13614,N_13500);
nand UO_1974 (O_1974,N_14525,N_13793);
xor UO_1975 (O_1975,N_14815,N_14022);
xnor UO_1976 (O_1976,N_13665,N_14514);
or UO_1977 (O_1977,N_14138,N_14101);
nand UO_1978 (O_1978,N_14019,N_13863);
nand UO_1979 (O_1979,N_14801,N_14956);
or UO_1980 (O_1980,N_14639,N_13520);
xor UO_1981 (O_1981,N_13550,N_13626);
nor UO_1982 (O_1982,N_13603,N_13852);
or UO_1983 (O_1983,N_13905,N_14757);
xor UO_1984 (O_1984,N_13803,N_13753);
xor UO_1985 (O_1985,N_14575,N_14365);
xnor UO_1986 (O_1986,N_13744,N_14351);
xnor UO_1987 (O_1987,N_14269,N_14944);
and UO_1988 (O_1988,N_14342,N_14436);
nand UO_1989 (O_1989,N_14103,N_14963);
or UO_1990 (O_1990,N_13928,N_14008);
xnor UO_1991 (O_1991,N_14018,N_14100);
or UO_1992 (O_1992,N_14137,N_14417);
or UO_1993 (O_1993,N_14856,N_14240);
xor UO_1994 (O_1994,N_14042,N_13635);
nor UO_1995 (O_1995,N_13780,N_14109);
nor UO_1996 (O_1996,N_14639,N_14287);
or UO_1997 (O_1997,N_14854,N_13857);
nand UO_1998 (O_1998,N_14495,N_14801);
or UO_1999 (O_1999,N_14548,N_14770);
endmodule