module basic_2000_20000_2500_20_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_1606,In_1123);
nor U1 (N_1,In_1719,In_861);
nand U2 (N_2,In_1436,In_271);
and U3 (N_3,In_76,In_575);
xor U4 (N_4,In_1622,In_1638);
and U5 (N_5,In_338,In_1852);
nor U6 (N_6,In_9,In_1118);
and U7 (N_7,In_495,In_1280);
nor U8 (N_8,In_441,In_1432);
or U9 (N_9,In_1954,In_1505);
and U10 (N_10,In_1182,In_673);
xnor U11 (N_11,In_1600,In_1375);
or U12 (N_12,In_1336,In_1463);
nor U13 (N_13,In_925,In_966);
nand U14 (N_14,In_1973,In_114);
and U15 (N_15,In_1941,In_842);
xnor U16 (N_16,In_300,In_1823);
and U17 (N_17,In_778,In_1833);
xor U18 (N_18,In_866,In_1758);
xor U19 (N_19,In_1785,In_762);
and U20 (N_20,In_1437,In_480);
and U21 (N_21,In_474,In_1143);
or U22 (N_22,In_753,In_543);
and U23 (N_23,In_1316,In_1189);
xnor U24 (N_24,In_1510,In_72);
xor U25 (N_25,In_377,In_1443);
nor U26 (N_26,In_407,In_876);
nor U27 (N_27,In_1936,In_396);
nand U28 (N_28,In_1926,In_1836);
and U29 (N_29,In_1656,In_1482);
and U30 (N_30,In_505,In_157);
xor U31 (N_31,In_1916,In_428);
or U32 (N_32,In_1642,In_1745);
nor U33 (N_33,In_1035,In_36);
nor U34 (N_34,In_454,In_1038);
and U35 (N_35,In_874,In_134);
and U36 (N_36,In_1063,In_481);
xor U37 (N_37,In_164,In_101);
nand U38 (N_38,In_1131,In_1932);
and U39 (N_39,In_855,In_1746);
or U40 (N_40,In_754,In_1707);
or U41 (N_41,In_1085,In_1668);
or U42 (N_42,In_1697,In_295);
and U43 (N_43,In_282,In_639);
nand U44 (N_44,In_1019,In_1790);
xnor U45 (N_45,In_179,In_1200);
nand U46 (N_46,In_1552,In_989);
and U47 (N_47,In_1540,In_961);
or U48 (N_48,In_1160,In_1256);
xor U49 (N_49,In_1507,In_446);
and U50 (N_50,In_1636,In_1257);
and U51 (N_51,In_1012,In_468);
or U52 (N_52,In_1528,In_1365);
or U53 (N_53,In_805,In_1975);
or U54 (N_54,In_1420,In_435);
xnor U55 (N_55,In_689,In_1048);
and U56 (N_56,In_1494,In_491);
nand U57 (N_57,In_1457,In_1797);
nand U58 (N_58,In_378,In_276);
nor U59 (N_59,In_578,In_1736);
and U60 (N_60,In_1541,In_1831);
nor U61 (N_61,In_1146,In_401);
xor U62 (N_62,In_303,In_1405);
nand U63 (N_63,In_1914,In_1047);
xnor U64 (N_64,In_54,In_1379);
nand U65 (N_65,In_1276,In_644);
nand U66 (N_66,In_1088,In_14);
nand U67 (N_67,In_13,In_75);
xnor U68 (N_68,In_761,In_756);
and U69 (N_69,In_1391,In_1213);
nand U70 (N_70,In_1421,In_1979);
nor U71 (N_71,In_1079,In_133);
nand U72 (N_72,In_626,In_970);
nor U73 (N_73,In_12,In_1570);
or U74 (N_74,In_1206,In_414);
nand U75 (N_75,In_1748,In_417);
or U76 (N_76,In_78,In_1907);
nand U77 (N_77,In_1920,In_1524);
and U78 (N_78,In_26,In_1199);
and U79 (N_79,In_865,In_992);
and U80 (N_80,In_1655,In_801);
and U81 (N_81,In_1547,In_594);
and U82 (N_82,In_918,In_1468);
nand U83 (N_83,In_1119,In_1929);
and U84 (N_84,In_1589,In_1658);
xnor U85 (N_85,In_1779,In_1369);
xnor U86 (N_86,In_1575,In_261);
nand U87 (N_87,In_522,In_343);
nand U88 (N_88,In_252,In_1531);
xnor U89 (N_89,In_766,In_385);
xor U90 (N_90,In_1472,In_671);
and U91 (N_91,In_741,In_1627);
xor U92 (N_92,In_1176,In_541);
and U93 (N_93,In_1350,In_706);
and U94 (N_94,In_82,In_1065);
or U95 (N_95,In_342,In_1803);
nand U96 (N_96,In_1827,In_322);
or U97 (N_97,In_1765,In_1764);
xnor U98 (N_98,In_154,In_674);
or U99 (N_99,In_686,In_1599);
nor U100 (N_100,In_1159,In_77);
and U101 (N_101,In_166,In_582);
nor U102 (N_102,In_655,In_1837);
or U103 (N_103,In_1931,In_283);
xnor U104 (N_104,In_449,In_516);
or U105 (N_105,In_1234,In_56);
xnor U106 (N_106,In_1177,In_1426);
or U107 (N_107,In_816,In_1657);
nor U108 (N_108,In_846,In_1069);
xnor U109 (N_109,In_1989,In_1843);
nor U110 (N_110,In_1824,In_1112);
nand U111 (N_111,In_158,In_251);
nand U112 (N_112,In_422,In_199);
nand U113 (N_113,In_210,In_270);
xnor U114 (N_114,In_1043,In_145);
nor U115 (N_115,In_1191,In_1986);
nand U116 (N_116,In_203,In_826);
xor U117 (N_117,In_1485,In_1683);
xnor U118 (N_118,In_739,In_908);
xor U119 (N_119,In_990,In_952);
nor U120 (N_120,In_1586,In_650);
nor U121 (N_121,In_1462,In_1912);
nand U122 (N_122,In_744,In_654);
nand U123 (N_123,In_1927,In_539);
and U124 (N_124,In_28,In_1360);
xor U125 (N_125,In_897,In_745);
nand U126 (N_126,In_1110,In_714);
and U127 (N_127,In_1741,In_469);
nor U128 (N_128,In_953,In_1724);
nor U129 (N_129,In_1013,In_1471);
nand U130 (N_130,In_35,In_1641);
or U131 (N_131,In_891,In_1637);
and U132 (N_132,In_1195,In_1645);
nand U133 (N_133,In_1513,In_968);
and U134 (N_134,In_1704,In_1001);
or U135 (N_135,In_1714,In_152);
nor U136 (N_136,In_1574,In_1755);
nor U137 (N_137,In_796,In_1988);
nor U138 (N_138,In_1009,In_239);
and U139 (N_139,In_1382,In_433);
or U140 (N_140,In_1067,In_535);
and U141 (N_141,In_1080,In_171);
nand U142 (N_142,In_1474,In_1192);
nand U143 (N_143,In_1242,In_976);
nor U144 (N_144,In_1151,In_1971);
nor U145 (N_145,In_964,In_1684);
nand U146 (N_146,In_1811,In_1629);
or U147 (N_147,In_625,In_160);
xnor U148 (N_148,In_1533,In_364);
and U149 (N_149,In_841,In_734);
and U150 (N_150,In_220,In_1813);
and U151 (N_151,In_1572,In_643);
and U152 (N_152,In_1150,In_257);
and U153 (N_153,In_1686,In_1839);
or U154 (N_154,In_2,In_566);
and U155 (N_155,In_1096,In_603);
xor U156 (N_156,In_588,In_852);
and U157 (N_157,In_301,In_1265);
nand U158 (N_158,In_290,In_89);
nand U159 (N_159,In_888,In_1559);
or U160 (N_160,In_1408,In_965);
or U161 (N_161,In_1838,In_1963);
nor U162 (N_162,In_1041,In_1097);
nor U163 (N_163,In_1221,In_1105);
nand U164 (N_164,In_1720,In_799);
and U165 (N_165,In_906,In_1680);
xnor U166 (N_166,In_1300,In_723);
nand U167 (N_167,In_1732,In_279);
nand U168 (N_168,In_461,In_1671);
xor U169 (N_169,In_223,In_1654);
xnor U170 (N_170,In_629,In_911);
nand U171 (N_171,In_399,In_1923);
nor U172 (N_172,In_1278,In_1084);
nand U173 (N_173,In_1075,In_875);
nand U174 (N_174,In_949,In_1);
or U175 (N_175,In_904,In_1477);
nand U176 (N_176,In_467,In_138);
and U177 (N_177,In_559,In_1279);
and U178 (N_178,In_529,In_871);
or U179 (N_179,In_326,In_518);
nor U180 (N_180,In_752,In_306);
or U181 (N_181,In_46,In_605);
xnor U182 (N_182,In_498,In_662);
and U183 (N_183,In_1120,In_1835);
nand U184 (N_184,In_1938,In_1194);
or U185 (N_185,In_1733,In_1848);
xor U186 (N_186,In_116,In_1784);
or U187 (N_187,In_413,In_659);
xor U188 (N_188,In_1040,In_1698);
nor U189 (N_189,In_1174,In_331);
or U190 (N_190,In_738,In_19);
or U191 (N_191,In_1441,In_519);
and U192 (N_192,In_1446,In_1706);
and U193 (N_193,In_269,In_1701);
or U194 (N_194,In_144,In_509);
nor U195 (N_195,In_997,In_959);
nor U196 (N_196,In_452,In_254);
or U197 (N_197,In_1220,In_1996);
nand U198 (N_198,In_472,In_1325);
and U199 (N_199,In_1309,In_808);
or U200 (N_200,In_1202,In_242);
nand U201 (N_201,In_1321,In_471);
or U202 (N_202,In_1076,In_1111);
or U203 (N_203,In_515,In_488);
or U204 (N_204,In_48,In_1774);
or U205 (N_205,In_1530,In_363);
nand U206 (N_206,In_255,In_695);
and U207 (N_207,In_1165,In_767);
nand U208 (N_208,In_1252,In_137);
xor U209 (N_209,In_163,In_716);
or U210 (N_210,In_1277,In_309);
and U211 (N_211,In_190,In_649);
nand U212 (N_212,In_638,In_1427);
nand U213 (N_213,In_1224,In_1334);
and U214 (N_214,In_1503,In_1315);
and U215 (N_215,In_1526,In_1987);
or U216 (N_216,In_1361,In_704);
xor U217 (N_217,In_1699,In_1725);
nor U218 (N_218,In_464,In_1240);
nand U219 (N_219,In_416,In_1885);
xor U220 (N_220,In_1977,In_1121);
nor U221 (N_221,In_933,In_1125);
nor U222 (N_222,In_1549,In_1893);
nor U223 (N_223,In_889,In_1287);
xor U224 (N_224,In_533,In_1212);
nand U225 (N_225,In_49,In_1461);
or U226 (N_226,In_1208,In_1219);
xor U227 (N_227,In_1751,In_1281);
nand U228 (N_228,In_833,In_1509);
nand U229 (N_229,In_79,In_424);
nand U230 (N_230,In_1241,In_1819);
nand U231 (N_231,In_130,In_688);
xor U232 (N_232,In_1381,In_88);
or U233 (N_233,In_125,In_1367);
xor U234 (N_234,In_1849,In_18);
xnor U235 (N_235,In_1928,In_1267);
xor U236 (N_236,In_118,In_1608);
or U237 (N_237,In_677,In_1335);
or U238 (N_238,In_486,In_1856);
nand U239 (N_239,In_727,In_353);
or U240 (N_240,In_569,In_437);
xnor U241 (N_241,In_1868,In_1203);
and U242 (N_242,In_785,In_1138);
xor U243 (N_243,In_1229,In_366);
xor U244 (N_244,In_647,In_1245);
or U245 (N_245,In_1034,In_1995);
xor U246 (N_246,In_1635,In_1139);
or U247 (N_247,In_1007,In_1949);
and U248 (N_248,In_980,In_1883);
and U249 (N_249,In_549,In_737);
xnor U250 (N_250,In_1429,In_1005);
or U251 (N_251,In_1380,In_1945);
and U252 (N_252,In_1897,In_1127);
nor U253 (N_253,In_1372,In_560);
xnor U254 (N_254,In_574,In_1233);
nor U255 (N_255,In_1348,In_357);
xnor U256 (N_256,In_1491,In_1662);
nor U257 (N_257,In_1337,In_969);
or U258 (N_258,In_334,In_907);
nor U259 (N_259,In_1623,In_883);
xor U260 (N_260,In_419,In_1016);
xnor U261 (N_261,In_71,In_929);
or U262 (N_262,In_96,In_1866);
or U263 (N_263,In_1994,In_1809);
and U264 (N_264,In_863,In_1749);
and U265 (N_265,In_356,In_1435);
nand U266 (N_266,In_730,In_248);
or U267 (N_267,In_1157,In_487);
xnor U268 (N_268,In_1767,In_839);
nand U269 (N_269,In_576,In_293);
nand U270 (N_270,In_1665,In_1403);
and U271 (N_271,In_1042,In_100);
nor U272 (N_272,In_1935,In_1997);
nor U273 (N_273,In_87,In_1922);
and U274 (N_274,In_1341,In_760);
or U275 (N_275,In_665,In_405);
nand U276 (N_276,In_1685,In_460);
or U277 (N_277,In_409,In_1388);
xor U278 (N_278,In_1900,In_1306);
nor U279 (N_279,In_1478,In_408);
nand U280 (N_280,In_1404,In_1320);
or U281 (N_281,In_31,In_943);
nor U282 (N_282,In_479,In_1141);
nand U283 (N_283,In_1615,In_939);
nor U284 (N_284,In_86,In_824);
and U285 (N_285,In_172,In_1387);
nor U286 (N_286,In_1882,In_1310);
or U287 (N_287,In_854,In_1937);
and U288 (N_288,In_979,In_1296);
xor U289 (N_289,In_1061,In_1134);
xnor U290 (N_290,In_1129,In_1077);
nor U291 (N_291,In_1798,In_847);
or U292 (N_292,In_104,In_60);
nor U293 (N_293,In_517,In_264);
nor U294 (N_294,In_1142,In_857);
and U295 (N_295,In_1674,In_429);
or U296 (N_296,In_1425,In_432);
or U297 (N_297,In_1888,In_1498);
and U298 (N_298,In_1413,In_757);
nor U299 (N_299,In_1448,In_1616);
xor U300 (N_300,In_243,In_1564);
and U301 (N_301,In_1484,In_563);
xor U302 (N_302,In_1617,In_1032);
or U303 (N_303,In_1217,In_1205);
xor U304 (N_304,In_1844,In_1512);
and U305 (N_305,In_1740,In_1487);
nor U306 (N_306,In_607,In_1976);
nor U307 (N_307,In_958,In_860);
or U308 (N_308,In_602,In_1639);
or U309 (N_309,In_1169,In_1132);
xor U310 (N_310,In_1268,In_1308);
and U311 (N_311,In_1373,In_1517);
nor U312 (N_312,In_656,In_934);
or U313 (N_313,In_622,In_1990);
and U314 (N_314,In_807,In_1652);
and U315 (N_315,In_1021,In_570);
or U316 (N_316,In_1126,In_97);
xnor U317 (N_317,In_368,In_1679);
xor U318 (N_318,In_849,In_1626);
and U319 (N_319,In_456,In_721);
and U320 (N_320,In_63,In_38);
or U321 (N_321,In_371,In_691);
nand U322 (N_322,In_1480,In_151);
xor U323 (N_323,In_636,In_1948);
and U324 (N_324,In_1962,In_614);
nor U325 (N_325,In_214,In_1548);
xnor U326 (N_326,In_1793,In_848);
nor U327 (N_327,In_347,In_1416);
and U328 (N_328,In_1290,In_1322);
nor U329 (N_329,In_782,In_1311);
nand U330 (N_330,In_355,In_404);
and U331 (N_331,In_877,In_94);
xnor U332 (N_332,In_1460,In_170);
or U333 (N_333,In_1822,In_129);
xor U334 (N_334,In_1392,In_209);
nand U335 (N_335,In_617,In_1522);
or U336 (N_336,In_1190,In_1044);
xnor U337 (N_337,In_1397,In_201);
and U338 (N_338,In_735,In_1727);
nor U339 (N_339,In_827,In_1544);
xnor U340 (N_340,In_1921,In_1770);
or U341 (N_341,In_299,In_1317);
nand U342 (N_342,In_1282,In_387);
xor U343 (N_343,In_1913,In_176);
xnor U344 (N_344,In_1314,In_1394);
xor U345 (N_345,In_39,In_1781);
or U346 (N_346,In_561,In_1187);
and U347 (N_347,In_612,In_780);
nor U348 (N_348,In_121,In_1054);
and U349 (N_349,In_1560,In_287);
nor U350 (N_350,In_881,In_313);
nor U351 (N_351,In_1197,In_1612);
nor U352 (N_352,In_1087,In_29);
and U353 (N_353,In_593,In_259);
xnor U354 (N_354,In_775,In_333);
xor U355 (N_355,In_1892,In_1395);
and U356 (N_356,In_1231,In_20);
and U357 (N_357,In_384,In_1423);
xor U358 (N_358,In_1438,In_1663);
nor U359 (N_359,In_273,In_613);
or U360 (N_360,In_606,In_1525);
and U361 (N_361,In_710,In_971);
or U362 (N_362,In_1634,In_1539);
nor U363 (N_363,In_937,In_1292);
nand U364 (N_364,In_1017,In_1957);
nand U365 (N_365,In_661,In_542);
xnor U366 (N_366,In_1692,In_1853);
nand U367 (N_367,In_0,In_1004);
nor U368 (N_368,In_1008,In_1690);
nor U369 (N_369,In_1024,In_1542);
nor U370 (N_370,In_946,In_546);
nor U371 (N_371,In_65,In_351);
and U372 (N_372,In_1688,In_32);
or U373 (N_373,In_898,In_1237);
and U374 (N_374,In_1389,In_1855);
xnor U375 (N_375,In_892,In_1721);
nor U376 (N_376,In_608,In_224);
or U377 (N_377,In_1861,In_1687);
or U378 (N_378,In_1648,In_798);
nor U379 (N_379,In_7,In_69);
nor U380 (N_380,In_1368,In_1293);
nor U381 (N_381,In_879,In_1649);
and U382 (N_382,In_1737,In_1419);
or U383 (N_383,In_996,In_354);
or U384 (N_384,In_1434,In_553);
and U385 (N_385,In_110,In_470);
nor U386 (N_386,In_1068,In_554);
and U387 (N_387,In_676,In_149);
nand U388 (N_388,In_684,In_1998);
xnor U389 (N_389,In_1558,In_571);
nor U390 (N_390,In_978,In_1966);
nand U391 (N_391,In_1428,In_1625);
or U392 (N_392,In_1374,In_105);
xnor U393 (N_393,In_1073,In_503);
nor U394 (N_394,In_1284,In_1153);
and U395 (N_395,In_1595,In_818);
xnor U396 (N_396,In_1693,In_809);
xnor U397 (N_397,In_379,In_1919);
or U398 (N_398,In_1985,In_1624);
or U399 (N_399,In_308,In_1991);
nor U400 (N_400,In_592,In_944);
nand U401 (N_401,In_1376,In_858);
and U402 (N_402,In_1953,In_773);
xnor U403 (N_403,In_236,In_1891);
nor U404 (N_404,In_963,In_398);
nand U405 (N_405,In_1775,In_1248);
or U406 (N_406,In_1847,In_1884);
xor U407 (N_407,In_108,In_1418);
or U408 (N_408,In_713,In_1605);
xnor U409 (N_409,In_1584,In_1486);
and U410 (N_410,In_192,In_388);
and U411 (N_411,In_183,In_1653);
nor U412 (N_412,In_573,In_207);
nand U413 (N_413,In_1723,In_1804);
xnor U414 (N_414,In_330,In_823);
and U415 (N_415,In_1162,In_113);
and U416 (N_416,In_162,In_1841);
or U417 (N_417,In_289,In_169);
or U418 (N_418,In_1726,In_1225);
xnor U419 (N_419,In_1440,In_1058);
or U420 (N_420,In_1045,In_11);
or U421 (N_421,In_178,In_532);
nand U422 (N_422,In_1787,In_1274);
and U423 (N_423,In_143,In_1537);
nor U424 (N_424,In_1332,In_1845);
xnor U425 (N_425,In_736,In_1356);
nand U426 (N_426,In_931,In_1676);
and U427 (N_427,In_1064,In_499);
nor U428 (N_428,In_367,In_641);
or U429 (N_429,In_427,In_473);
or U430 (N_430,In_1091,In_870);
or U431 (N_431,In_418,In_1769);
xor U432 (N_432,In_1898,In_1585);
or U433 (N_433,In_1951,In_1890);
or U434 (N_434,In_475,In_1771);
and U435 (N_435,In_395,In_1786);
and U436 (N_436,In_1532,In_1304);
xnor U437 (N_437,In_1093,In_455);
and U438 (N_438,In_1496,In_423);
and U439 (N_439,In_394,In_1918);
nand U440 (N_440,In_564,In_1974);
or U441 (N_441,In_181,In_993);
nor U442 (N_442,In_1092,In_1609);
or U443 (N_443,In_204,In_1795);
nand U444 (N_444,In_30,In_272);
or U445 (N_445,In_572,In_731);
nor U446 (N_446,In_1878,In_402);
nand U447 (N_447,In_1902,In_1303);
xor U448 (N_448,In_896,In_135);
xnor U449 (N_449,In_635,In_450);
or U450 (N_450,In_266,In_1860);
and U451 (N_451,In_1062,In_987);
nor U452 (N_452,In_828,In_109);
nor U453 (N_453,In_537,In_1378);
xor U454 (N_454,In_159,In_813);
and U455 (N_455,In_604,In_728);
nand U456 (N_456,In_784,In_1894);
nor U457 (N_457,In_238,In_1579);
xnor U458 (N_458,In_955,In_1947);
nand U459 (N_459,In_619,In_1148);
or U460 (N_460,In_365,In_1659);
xor U461 (N_461,In_1896,In_168);
xor U462 (N_462,In_1535,In_1593);
nor U463 (N_463,In_658,In_1981);
xor U464 (N_464,In_350,In_1903);
or U465 (N_465,In_1980,In_1550);
nand U466 (N_466,In_972,In_591);
nor U467 (N_467,In_318,In_1270);
or U468 (N_468,In_16,In_781);
nand U469 (N_469,In_1571,In_1493);
nand U470 (N_470,In_1647,In_1555);
or U471 (N_471,In_768,In_584);
nor U472 (N_472,In_161,In_1810);
nor U473 (N_473,In_1604,In_1702);
nand U474 (N_474,In_814,In_1338);
nand U475 (N_475,In_648,In_234);
or U476 (N_476,In_631,In_1538);
or U477 (N_477,In_838,In_1851);
nor U478 (N_478,In_1551,In_1066);
and U479 (N_479,In_311,In_1459);
nand U480 (N_480,In_107,In_372);
or U481 (N_481,In_894,In_1501);
nand U482 (N_482,In_1266,In_500);
and U483 (N_483,In_493,In_1154);
or U484 (N_484,In_835,In_1239);
nand U485 (N_485,In_1840,In_1396);
nor U486 (N_486,In_587,In_1752);
or U487 (N_487,In_1098,In_250);
nor U488 (N_488,In_1523,In_262);
and U489 (N_489,In_1275,In_426);
and U490 (N_490,In_1911,In_797);
xnor U491 (N_491,In_589,In_1130);
xor U492 (N_492,In_899,In_1703);
nand U493 (N_493,In_451,In_991);
or U494 (N_494,In_1857,In_45);
and U495 (N_495,In_81,In_1215);
xnor U496 (N_496,In_941,In_1344);
nand U497 (N_497,In_146,In_103);
nand U498 (N_498,In_1670,In_93);
nor U499 (N_499,In_1832,In_1033);
nand U500 (N_500,In_1481,In_1346);
xnor U501 (N_501,In_1362,In_916);
and U502 (N_502,In_393,In_360);
nand U503 (N_503,In_256,In_502);
or U504 (N_504,In_683,In_1993);
nand U505 (N_505,In_200,In_193);
nor U506 (N_506,In_1667,In_1029);
and U507 (N_507,In_1789,In_74);
nor U508 (N_508,In_1956,In_600);
and U509 (N_509,In_1449,In_1877);
and U510 (N_510,In_1762,In_733);
nor U511 (N_511,In_1607,In_1881);
or U512 (N_512,In_1168,In_329);
or U513 (N_513,In_420,In_1036);
or U514 (N_514,In_1253,In_508);
xnor U515 (N_515,In_830,In_859);
xor U516 (N_516,In_1864,In_599);
xor U517 (N_517,In_40,In_1632);
nand U518 (N_518,In_869,In_1122);
nand U519 (N_519,In_173,In_1172);
nand U520 (N_520,In_1568,In_771);
or U521 (N_521,In_1052,In_1906);
nand U522 (N_522,In_278,In_1497);
and U523 (N_523,In_530,In_298);
nand U524 (N_524,In_924,In_187);
nor U525 (N_525,In_1327,In_1862);
and U526 (N_526,In_1454,In_1717);
nor U527 (N_527,In_1950,In_772);
nand U528 (N_528,In_1566,In_1519);
xnor U529 (N_529,In_5,In_1294);
nand U530 (N_530,In_1455,In_1490);
nor U531 (N_531,In_702,In_1155);
nor U532 (N_532,In_1716,In_206);
and U533 (N_533,In_1578,In_1651);
or U534 (N_534,In_1453,In_812);
and U535 (N_535,In_156,In_817);
and U536 (N_536,In_1089,In_672);
nor U537 (N_537,In_1136,In_1562);
nand U538 (N_538,In_267,In_265);
or U539 (N_539,In_235,In_175);
nand U540 (N_540,In_1992,In_177);
xnor U541 (N_541,In_1411,In_1761);
xnor U542 (N_542,In_339,In_1326);
or U543 (N_543,In_260,In_124);
and U544 (N_544,In_1511,In_319);
and U545 (N_545,In_751,In_1037);
xnor U546 (N_546,In_1263,In_923);
xnor U547 (N_547,In_1488,In_1982);
or U548 (N_548,In_1867,In_1152);
and U549 (N_549,In_1750,In_340);
nor U550 (N_550,In_729,In_912);
and U551 (N_551,In_485,In_186);
and U552 (N_552,In_803,In_776);
or U553 (N_553,In_637,In_174);
xnor U554 (N_554,In_227,In_1210);
and U555 (N_555,In_749,In_1871);
xor U556 (N_556,In_720,In_258);
nor U557 (N_557,In_1099,In_1520);
nor U558 (N_558,In_1661,In_1489);
nand U559 (N_559,In_1801,In_909);
or U560 (N_560,In_1082,In_1492);
xnor U561 (N_561,In_922,In_436);
or U562 (N_562,In_447,In_147);
nand U563 (N_563,In_380,In_577);
and U564 (N_564,In_1640,In_182);
or U565 (N_565,In_213,In_442);
nor U566 (N_566,In_1830,In_1958);
or U567 (N_567,In_61,In_1614);
xnor U568 (N_568,In_321,In_1700);
nand U569 (N_569,In_1621,In_868);
xnor U570 (N_570,In_701,In_595);
xnor U571 (N_571,In_1358,In_942);
nand U572 (N_572,In_1967,In_59);
or U573 (N_573,In_189,In_525);
and U574 (N_574,In_1788,In_1858);
nor U575 (N_575,In_1095,In_1385);
and U576 (N_576,In_1410,In_811);
or U577 (N_577,In_1430,In_1543);
xnor U578 (N_578,In_722,In_1518);
nand U579 (N_579,In_494,In_41);
and U580 (N_580,In_391,In_1620);
or U581 (N_581,In_1643,In_583);
xnor U582 (N_582,In_1880,In_1872);
nand U583 (N_583,In_932,In_1046);
or U584 (N_584,In_136,In_1483);
xnor U585 (N_585,In_55,In_1072);
or U586 (N_586,In_8,In_1401);
and U587 (N_587,In_1603,In_601);
and U588 (N_588,In_1826,In_1145);
xor U589 (N_589,In_1447,In_585);
and U590 (N_590,In_1582,In_85);
and U591 (N_591,In_618,In_1915);
nand U592 (N_592,In_957,In_307);
and U593 (N_593,In_905,In_1264);
nand U594 (N_594,In_579,In_1124);
and U595 (N_595,In_1960,In_443);
and U596 (N_596,In_586,In_1591);
or U597 (N_597,In_1709,In_1504);
nor U598 (N_598,In_1117,In_497);
xor U599 (N_599,In_316,In_590);
or U600 (N_600,In_1010,In_954);
nor U601 (N_601,In_822,In_247);
nor U602 (N_602,In_1534,In_774);
xor U603 (N_603,In_1283,In_862);
nor U604 (N_604,In_185,In_496);
nand U605 (N_605,In_275,In_787);
xnor U606 (N_606,In_1243,In_845);
nand U607 (N_607,In_682,In_1393);
nor U608 (N_608,In_1386,In_1407);
nand U609 (N_609,In_1128,In_1805);
nand U610 (N_610,In_1456,In_678);
xor U611 (N_611,In_1587,In_1020);
and U612 (N_612,In_1495,In_1102);
nand U613 (N_613,In_1227,In_1978);
and U614 (N_614,In_1964,In_57);
nand U615 (N_615,In_886,In_1027);
or U616 (N_616,In_712,In_540);
or U617 (N_617,In_598,In_538);
nor U618 (N_618,In_1944,In_715);
nand U619 (N_619,In_1870,In_374);
or U620 (N_620,In_1791,In_403);
and U621 (N_621,In_750,In_882);
or U622 (N_622,In_1100,In_218);
xor U623 (N_623,In_1000,In_726);
nand U624 (N_624,In_1228,In_1409);
nor U625 (N_625,In_349,In_960);
or U626 (N_626,In_1222,In_843);
and U627 (N_627,In_1815,In_127);
nor U628 (N_628,In_663,In_1756);
and U629 (N_629,In_1424,In_708);
or U630 (N_630,In_770,In_1450);
and U631 (N_631,In_1901,In_565);
and U632 (N_632,In_1984,In_1156);
or U633 (N_633,In_274,In_141);
and U634 (N_634,In_1238,In_1818);
and U635 (N_635,In_1713,In_80);
nand U636 (N_636,In_1768,In_1022);
and U637 (N_637,In_1464,In_1307);
nor U638 (N_638,In_216,In_920);
nand U639 (N_639,In_153,In_1766);
nor U640 (N_640,In_680,In_1646);
nor U641 (N_641,In_1955,In_382);
nor U642 (N_642,In_885,In_1295);
xor U643 (N_643,In_1193,In_1887);
nand U644 (N_644,In_1940,In_98);
nor U645 (N_645,In_112,In_1546);
xnor U646 (N_646,In_150,In_226);
nand U647 (N_647,In_253,In_596);
nand U648 (N_648,In_645,In_628);
nor U649 (N_649,In_476,In_901);
or U650 (N_650,In_1873,In_376);
nand U651 (N_651,In_707,In_1514);
or U652 (N_652,In_786,In_791);
or U653 (N_653,In_1414,In_392);
or U654 (N_654,In_47,In_1886);
nand U655 (N_655,In_975,In_1198);
or U656 (N_656,In_1086,In_1235);
xor U657 (N_657,In_370,In_1297);
nand U658 (N_658,In_793,In_1444);
nand U659 (N_659,In_783,In_1814);
xor U660 (N_660,In_1469,In_1342);
and U661 (N_661,In_51,In_523);
nor U662 (N_662,In_1247,In_1147);
and U663 (N_663,In_792,In_3);
nand U664 (N_664,In_653,In_245);
xor U665 (N_665,In_294,In_352);
and U666 (N_666,In_1272,In_795);
nand U667 (N_667,In_1014,In_1983);
nor U668 (N_668,In_1452,In_1794);
nor U669 (N_669,In_222,In_514);
or U670 (N_670,In_567,In_597);
nand U671 (N_671,In_790,In_1135);
nor U672 (N_672,In_1173,In_410);
nand U673 (N_673,In_821,In_375);
nand U674 (N_674,In_1596,In_1631);
nor U675 (N_675,In_928,In_1357);
xnor U676 (N_676,In_1672,In_652);
nor U677 (N_677,In_610,In_327);
xnor U678 (N_678,In_1925,In_1188);
nor U679 (N_679,In_1355,In_1343);
and U680 (N_680,In_73,In_998);
and U681 (N_681,In_1854,In_1285);
or U682 (N_682,In_690,In_195);
xnor U683 (N_683,In_430,In_1114);
nand U684 (N_684,In_632,In_1258);
nor U685 (N_685,In_844,In_1783);
or U686 (N_686,In_1133,In_940);
nor U687 (N_687,In_102,In_373);
and U688 (N_688,In_789,In_1113);
or U689 (N_689,In_291,In_1865);
or U690 (N_690,In_390,In_1644);
or U691 (N_691,In_1329,In_1628);
and U692 (N_692,In_24,In_1731);
nor U693 (N_693,In_646,In_1301);
or U694 (N_694,In_142,In_197);
or U695 (N_695,In_132,In_994);
or U696 (N_696,In_1108,In_501);
nor U697 (N_697,In_1415,In_44);
xor U698 (N_698,In_1006,In_956);
and U699 (N_699,In_281,In_510);
or U700 (N_700,In_155,In_288);
nor U701 (N_701,In_512,In_277);
nor U702 (N_702,In_1499,In_411);
nand U703 (N_703,In_1255,In_1875);
or U704 (N_704,In_856,In_1874);
nand U705 (N_705,In_1249,In_699);
nand U706 (N_706,In_37,In_884);
nor U707 (N_707,In_551,In_1972);
xor U708 (N_708,In_1056,In_4);
or U709 (N_709,In_1666,In_1942);
nor U710 (N_710,In_324,In_765);
and U711 (N_711,In_832,In_67);
xor U712 (N_712,In_1691,In_23);
xor U713 (N_713,In_120,In_581);
or U714 (N_714,In_1516,In_984);
or U715 (N_715,In_64,In_1179);
nand U716 (N_716,In_233,In_1305);
xor U717 (N_717,In_52,In_1952);
nor U718 (N_718,In_1782,In_90);
xor U719 (N_719,In_400,In_1298);
nand U720 (N_720,In_568,In_1026);
nand U721 (N_721,In_552,In_819);
xor U722 (N_722,In_709,In_1377);
xor U723 (N_723,In_229,In_747);
or U724 (N_724,In_634,In_1299);
nand U725 (N_725,In_128,In_1930);
and U726 (N_726,In_457,In_627);
nor U727 (N_727,In_1742,In_415);
or U728 (N_728,In_92,In_1103);
xor U729 (N_729,In_1500,In_1288);
nor U730 (N_730,In_221,In_1567);
nor U731 (N_731,In_232,In_1164);
and U732 (N_732,In_1476,In_337);
xor U733 (N_733,In_1601,In_1271);
nand U734 (N_734,In_1869,In_740);
nand U735 (N_735,In_640,In_1739);
xnor U736 (N_736,In_463,In_1816);
or U737 (N_737,In_490,In_1244);
xnor U738 (N_738,In_1715,In_412);
and U739 (N_739,In_544,In_165);
or U740 (N_740,In_1318,In_167);
or U741 (N_741,In_945,In_1465);
nand U742 (N_742,In_111,In_1214);
and U743 (N_743,In_1184,In_1023);
xor U744 (N_744,In_131,In_825);
xor U745 (N_745,In_1743,In_359);
nor U746 (N_746,In_630,In_1286);
nor U747 (N_747,In_1859,In_1689);
or U748 (N_748,In_815,In_902);
and U749 (N_749,In_1594,In_1695);
and U750 (N_750,In_53,In_346);
nor U751 (N_751,In_555,In_919);
nand U752 (N_752,In_1778,In_421);
xor U753 (N_753,In_1399,In_759);
xor U754 (N_754,In_1776,In_1158);
or U755 (N_755,In_1371,In_1879);
nor U756 (N_756,In_936,In_332);
nand U757 (N_757,In_225,In_717);
nand U758 (N_758,In_205,In_642);
nor U759 (N_759,In_1170,In_1850);
and U760 (N_760,In_1965,In_1780);
xnor U761 (N_761,In_1144,In_675);
and U762 (N_762,In_1754,In_1470);
nor U763 (N_763,In_1529,In_837);
nand U764 (N_764,In_1934,In_1613);
nand U765 (N_765,In_302,In_660);
or U766 (N_766,In_1402,In_527);
nand U767 (N_767,In_358,In_1431);
and U768 (N_768,In_1347,In_986);
nand U769 (N_769,In_50,In_938);
or U770 (N_770,In_434,In_1090);
or U771 (N_771,In_1999,In_679);
or U772 (N_772,In_1106,In_1031);
nand U773 (N_773,In_1515,In_1055);
or U774 (N_774,In_703,In_962);
xor U775 (N_775,In_558,In_431);
nand U776 (N_776,In_1181,In_1633);
xor U777 (N_777,In_1598,In_520);
nand U778 (N_778,In_1889,In_1028);
xor U779 (N_779,In_297,In_1412);
or U780 (N_780,In_1807,In_1137);
nand U781 (N_781,In_1057,In_1025);
and U782 (N_782,In_633,In_33);
nand U783 (N_783,In_725,In_536);
xnor U784 (N_784,In_1508,In_1506);
nand U785 (N_785,In_1664,In_1384);
nand U786 (N_786,In_1711,In_1149);
and U787 (N_787,In_1475,In_1094);
xor U788 (N_788,In_1289,In_386);
nor U789 (N_789,In_43,In_913);
nor U790 (N_790,In_1969,In_1536);
nor U791 (N_791,In_1821,In_1049);
nand U792 (N_792,In_1445,In_1223);
and U793 (N_793,In_700,In_1261);
and U794 (N_794,In_531,In_930);
nor U795 (N_795,In_915,In_804);
and U796 (N_796,In_1619,In_1422);
xor U797 (N_797,In_1050,In_1772);
and U798 (N_798,In_180,In_748);
and U799 (N_799,In_853,In_1796);
or U800 (N_800,In_215,In_657);
nor U801 (N_801,In_348,In_361);
and U802 (N_802,In_1003,In_1178);
nand U803 (N_803,In_1924,In_1760);
xnor U804 (N_804,In_1565,In_513);
xor U805 (N_805,In_927,In_1576);
nand U806 (N_806,In_240,In_526);
xnor U807 (N_807,In_280,In_1502);
nand U808 (N_808,In_196,In_829);
and U809 (N_809,In_1561,In_459);
and U810 (N_810,In_973,In_711);
and U811 (N_811,In_99,In_914);
xnor U812 (N_812,In_1051,In_381);
xor U813 (N_813,In_763,In_1345);
and U814 (N_814,In_1011,In_1580);
and U815 (N_815,In_1115,In_806);
or U816 (N_816,In_1390,In_478);
nor U817 (N_817,In_1825,In_208);
xor U818 (N_818,In_1939,In_550);
xnor U819 (N_819,In_140,In_462);
nand U820 (N_820,In_948,In_263);
nand U821 (N_821,In_1610,In_448);
or U822 (N_822,In_1353,In_191);
and U823 (N_823,In_1030,In_1186);
or U824 (N_824,In_268,In_947);
or U825 (N_825,In_1808,In_504);
xnor U826 (N_826,In_623,In_1398);
or U827 (N_827,In_524,In_1406);
and U828 (N_828,In_1351,In_465);
nand U829 (N_829,In_1829,In_1682);
and U830 (N_830,In_880,In_17);
nand U831 (N_831,In_1763,In_694);
nand U832 (N_832,In_1554,In_438);
xnor U833 (N_833,In_696,In_794);
or U834 (N_834,In_123,In_988);
or U835 (N_835,In_285,In_1340);
and U836 (N_836,In_1236,In_336);
nor U837 (N_837,In_506,In_687);
or U838 (N_838,In_548,In_230);
or U839 (N_839,In_1660,In_42);
nand U840 (N_840,In_698,In_1577);
nand U841 (N_841,In_202,In_1581);
and U842 (N_842,In_511,In_341);
nor U843 (N_843,In_1354,In_1207);
and U844 (N_844,In_820,In_1744);
and U845 (N_845,In_1442,In_1196);
nor U846 (N_846,In_482,In_325);
xnor U847 (N_847,In_895,In_21);
and U848 (N_848,In_1573,In_1705);
and U849 (N_849,In_1729,In_1753);
xor U850 (N_850,In_1201,In_1820);
nor U851 (N_851,In_1232,In_1211);
nor U852 (N_852,In_1269,In_1364);
and U853 (N_853,In_697,In_1728);
and U854 (N_854,In_237,In_1339);
or U855 (N_855,In_484,In_983);
and U856 (N_856,In_15,In_1324);
nor U857 (N_857,In_1933,In_425);
and U858 (N_858,In_1466,In_246);
xor U859 (N_859,In_83,In_362);
and U860 (N_860,In_1171,In_1273);
or U861 (N_861,In_685,In_864);
and U862 (N_862,In_1259,In_1718);
xnor U863 (N_863,In_534,In_620);
and U864 (N_864,In_58,In_1330);
xor U865 (N_865,In_310,In_184);
nand U866 (N_866,In_1333,In_1757);
and U867 (N_867,In_1553,In_249);
and U868 (N_868,In_758,In_624);
and U869 (N_869,In_802,In_439);
nor U870 (N_870,In_91,In_406);
nor U871 (N_871,In_1590,In_974);
xnor U872 (N_872,In_119,In_1712);
and U873 (N_873,In_231,In_557);
nor U874 (N_874,In_1291,In_1246);
nor U875 (N_875,In_1738,In_1773);
nor U876 (N_876,In_834,In_556);
xor U877 (N_877,In_62,In_788);
nand U878 (N_878,In_383,In_1078);
and U879 (N_879,In_1302,In_126);
and U880 (N_880,In_1060,In_1039);
nand U881 (N_881,In_389,In_1053);
nand U882 (N_882,In_1323,In_1071);
and U883 (N_883,In_1313,In_1943);
nor U884 (N_884,In_198,In_1569);
or U885 (N_885,In_669,In_1451);
or U886 (N_886,In_926,In_1183);
xor U887 (N_887,In_115,In_1905);
nor U888 (N_888,In_212,In_292);
nor U889 (N_889,In_800,In_1669);
xnor U890 (N_890,In_743,In_1015);
or U891 (N_891,In_724,In_1140);
and U892 (N_892,In_1545,In_1166);
nor U893 (N_893,In_1909,In_1910);
and U894 (N_894,In_917,In_445);
nor U895 (N_895,In_1262,In_507);
nand U896 (N_896,In_6,In_615);
nor U897 (N_897,In_1527,In_117);
or U898 (N_898,In_1230,In_1678);
xnor U899 (N_899,In_995,In_244);
and U900 (N_900,In_1204,In_296);
nand U901 (N_901,In_66,In_1250);
nor U902 (N_902,In_910,In_1968);
or U903 (N_903,In_1946,In_609);
nor U904 (N_904,In_68,In_1175);
nand U905 (N_905,In_779,In_440);
or U906 (N_906,In_1439,In_1349);
or U907 (N_907,In_777,In_139);
and U908 (N_908,In_492,In_25);
and U909 (N_909,In_982,In_95);
nor U910 (N_910,In_1583,In_489);
nand U911 (N_911,In_1319,In_521);
and U912 (N_912,In_528,In_1180);
nor U913 (N_913,In_873,In_1328);
nor U914 (N_914,In_1109,In_1167);
and U915 (N_915,In_1694,In_1863);
or U916 (N_916,In_1730,In_312);
and U917 (N_917,In_228,In_1473);
nand U918 (N_918,In_1722,In_122);
nor U919 (N_919,In_893,In_985);
xor U920 (N_920,In_84,In_1521);
nor U921 (N_921,In_1710,In_315);
or U922 (N_922,In_188,In_1366);
or U923 (N_923,In_836,In_323);
or U924 (N_924,In_219,In_305);
and U925 (N_925,In_562,In_746);
nor U926 (N_926,In_1018,In_900);
and U927 (N_927,In_1185,In_328);
xor U928 (N_928,In_304,In_1557);
nand U929 (N_929,In_1458,In_70);
and U930 (N_930,In_1735,In_1959);
xnor U931 (N_931,In_764,In_718);
nand U932 (N_932,In_1611,In_1216);
nand U933 (N_933,In_867,In_1734);
or U934 (N_934,In_1370,In_314);
nor U935 (N_935,In_1618,In_1602);
or U936 (N_936,In_1363,In_951);
nor U937 (N_937,In_1681,In_1400);
nand U938 (N_938,In_967,In_1163);
nor U939 (N_939,In_1226,In_1083);
xor U940 (N_940,In_681,In_217);
and U941 (N_941,In_1846,In_1895);
and U942 (N_942,In_651,In_458);
or U943 (N_943,In_1359,In_1254);
or U944 (N_944,In_1563,In_742);
and U945 (N_945,In_1904,In_1834);
xor U946 (N_946,In_840,In_1792);
nor U947 (N_947,In_887,In_664);
xnor U948 (N_948,In_1074,In_903);
nor U949 (N_949,In_670,In_1556);
and U950 (N_950,In_1417,In_1101);
and U951 (N_951,In_999,In_1777);
or U952 (N_952,In_1800,In_719);
or U953 (N_953,In_621,In_755);
or U954 (N_954,In_545,In_935);
xor U955 (N_955,In_1806,In_320);
nand U956 (N_956,In_1352,In_693);
and U957 (N_957,In_1961,In_950);
nand U958 (N_958,In_1209,In_1251);
xnor U959 (N_959,In_1467,In_890);
nor U960 (N_960,In_1588,In_1817);
or U961 (N_961,In_477,In_981);
nor U962 (N_962,In_1161,In_1799);
and U963 (N_963,In_831,In_453);
or U964 (N_964,In_10,In_344);
or U965 (N_965,In_1899,In_1677);
nor U966 (N_966,In_850,In_1104);
and U967 (N_967,In_1081,In_1812);
and U968 (N_968,In_921,In_547);
or U969 (N_969,In_466,In_810);
and U970 (N_970,In_1673,In_666);
xor U971 (N_971,In_878,In_284);
or U972 (N_972,In_148,In_1708);
and U973 (N_973,In_194,In_1479);
xor U974 (N_974,In_286,In_616);
or U975 (N_975,In_1116,In_1331);
nand U976 (N_976,In_580,In_211);
nand U977 (N_977,In_1002,In_1107);
xnor U978 (N_978,In_732,In_345);
nor U979 (N_979,In_692,In_1592);
xor U980 (N_980,In_34,In_444);
nor U981 (N_981,In_611,In_1759);
and U982 (N_982,In_667,In_1842);
nor U983 (N_983,In_1917,In_1597);
nand U984 (N_984,In_1630,In_1696);
and U985 (N_985,In_317,In_335);
nor U986 (N_986,In_977,In_483);
xor U987 (N_987,In_1802,In_1908);
and U988 (N_988,In_1260,In_872);
xor U989 (N_989,In_1828,In_851);
nor U990 (N_990,In_1970,In_22);
or U991 (N_991,In_241,In_668);
nor U992 (N_992,In_1650,In_369);
or U993 (N_993,In_1876,In_397);
and U994 (N_994,In_1675,In_1747);
nand U995 (N_995,In_106,In_27);
and U996 (N_996,In_1070,In_1433);
nand U997 (N_997,In_1312,In_1218);
and U998 (N_998,In_769,In_1383);
nor U999 (N_999,In_1059,In_705);
xor U1000 (N_1000,N_839,N_788);
or U1001 (N_1001,N_682,N_335);
or U1002 (N_1002,N_338,N_49);
and U1003 (N_1003,N_240,N_252);
xnor U1004 (N_1004,N_887,N_107);
xnor U1005 (N_1005,N_553,N_111);
and U1006 (N_1006,N_621,N_869);
and U1007 (N_1007,N_285,N_224);
nor U1008 (N_1008,N_376,N_593);
nor U1009 (N_1009,N_481,N_613);
and U1010 (N_1010,N_550,N_922);
nor U1011 (N_1011,N_628,N_436);
nand U1012 (N_1012,N_87,N_460);
or U1013 (N_1013,N_449,N_592);
and U1014 (N_1014,N_600,N_320);
xor U1015 (N_1015,N_42,N_323);
or U1016 (N_1016,N_982,N_685);
or U1017 (N_1017,N_80,N_871);
nand U1018 (N_1018,N_619,N_368);
nand U1019 (N_1019,N_640,N_693);
or U1020 (N_1020,N_511,N_399);
and U1021 (N_1021,N_2,N_974);
nand U1022 (N_1022,N_563,N_393);
nand U1023 (N_1023,N_343,N_23);
xor U1024 (N_1024,N_182,N_454);
nor U1025 (N_1025,N_318,N_45);
xnor U1026 (N_1026,N_911,N_832);
and U1027 (N_1027,N_505,N_325);
nor U1028 (N_1028,N_420,N_558);
and U1029 (N_1029,N_488,N_777);
or U1030 (N_1030,N_211,N_298);
or U1031 (N_1031,N_733,N_362);
or U1032 (N_1032,N_708,N_296);
or U1033 (N_1033,N_208,N_434);
and U1034 (N_1034,N_303,N_265);
nor U1035 (N_1035,N_177,N_422);
xor U1036 (N_1036,N_329,N_981);
xor U1037 (N_1037,N_122,N_227);
and U1038 (N_1038,N_664,N_366);
xor U1039 (N_1039,N_926,N_246);
and U1040 (N_1040,N_586,N_26);
and U1041 (N_1041,N_704,N_514);
nor U1042 (N_1042,N_221,N_548);
nand U1043 (N_1043,N_656,N_985);
nor U1044 (N_1044,N_372,N_521);
and U1045 (N_1045,N_123,N_602);
xor U1046 (N_1046,N_409,N_22);
or U1047 (N_1047,N_643,N_63);
or U1048 (N_1048,N_849,N_197);
or U1049 (N_1049,N_769,N_873);
or U1050 (N_1050,N_618,N_61);
nand U1051 (N_1051,N_465,N_357);
xnor U1052 (N_1052,N_520,N_353);
nand U1053 (N_1053,N_743,N_146);
nor U1054 (N_1054,N_858,N_248);
nand U1055 (N_1055,N_575,N_421);
xor U1056 (N_1056,N_863,N_400);
nand U1057 (N_1057,N_599,N_482);
or U1058 (N_1058,N_352,N_805);
nor U1059 (N_1059,N_220,N_569);
nand U1060 (N_1060,N_53,N_95);
or U1061 (N_1061,N_894,N_75);
nor U1062 (N_1062,N_844,N_311);
and U1063 (N_1063,N_48,N_897);
and U1064 (N_1064,N_786,N_31);
and U1065 (N_1065,N_412,N_949);
xnor U1066 (N_1066,N_756,N_155);
or U1067 (N_1067,N_314,N_179);
nand U1068 (N_1068,N_468,N_895);
nand U1069 (N_1069,N_652,N_712);
nand U1070 (N_1070,N_793,N_219);
nor U1071 (N_1071,N_251,N_681);
nor U1072 (N_1072,N_52,N_294);
or U1073 (N_1073,N_886,N_29);
or U1074 (N_1074,N_181,N_910);
xor U1075 (N_1075,N_459,N_138);
nand U1076 (N_1076,N_692,N_40);
xnor U1077 (N_1077,N_716,N_310);
nor U1078 (N_1078,N_626,N_730);
nand U1079 (N_1079,N_143,N_280);
or U1080 (N_1080,N_164,N_257);
xnor U1081 (N_1081,N_753,N_565);
nor U1082 (N_1082,N_171,N_776);
nor U1083 (N_1083,N_767,N_200);
xnor U1084 (N_1084,N_526,N_649);
nor U1085 (N_1085,N_903,N_97);
xor U1086 (N_1086,N_697,N_942);
xor U1087 (N_1087,N_115,N_491);
xor U1088 (N_1088,N_929,N_6);
xnor U1089 (N_1089,N_616,N_884);
and U1090 (N_1090,N_659,N_554);
and U1091 (N_1091,N_984,N_165);
nand U1092 (N_1092,N_113,N_501);
nor U1093 (N_1093,N_448,N_54);
nand U1094 (N_1094,N_108,N_378);
xor U1095 (N_1095,N_846,N_67);
nand U1096 (N_1096,N_0,N_126);
and U1097 (N_1097,N_636,N_142);
and U1098 (N_1098,N_27,N_383);
nor U1099 (N_1099,N_939,N_951);
nand U1100 (N_1100,N_110,N_291);
xor U1101 (N_1101,N_429,N_850);
nor U1102 (N_1102,N_167,N_689);
or U1103 (N_1103,N_721,N_212);
and U1104 (N_1104,N_633,N_477);
xnor U1105 (N_1105,N_9,N_504);
and U1106 (N_1106,N_315,N_83);
and U1107 (N_1107,N_557,N_135);
nand U1108 (N_1108,N_398,N_348);
xnor U1109 (N_1109,N_3,N_268);
nand U1110 (N_1110,N_415,N_589);
nand U1111 (N_1111,N_464,N_798);
and U1112 (N_1112,N_892,N_433);
xor U1113 (N_1113,N_527,N_379);
and U1114 (N_1114,N_46,N_568);
nor U1115 (N_1115,N_317,N_327);
nand U1116 (N_1116,N_322,N_474);
or U1117 (N_1117,N_316,N_408);
xnor U1118 (N_1118,N_486,N_672);
nand U1119 (N_1119,N_133,N_28);
and U1120 (N_1120,N_510,N_861);
and U1121 (N_1121,N_471,N_19);
or U1122 (N_1122,N_867,N_301);
nand U1123 (N_1123,N_363,N_288);
nand U1124 (N_1124,N_856,N_779);
or U1125 (N_1125,N_269,N_432);
nand U1126 (N_1126,N_117,N_161);
nand U1127 (N_1127,N_202,N_157);
xnor U1128 (N_1128,N_967,N_187);
nor U1129 (N_1129,N_341,N_866);
nand U1130 (N_1130,N_1,N_783);
nor U1131 (N_1131,N_85,N_609);
nor U1132 (N_1132,N_438,N_544);
xnor U1133 (N_1133,N_444,N_282);
nand U1134 (N_1134,N_971,N_403);
xnor U1135 (N_1135,N_330,N_347);
xnor U1136 (N_1136,N_765,N_306);
nor U1137 (N_1137,N_760,N_620);
nor U1138 (N_1138,N_817,N_210);
and U1139 (N_1139,N_965,N_611);
xor U1140 (N_1140,N_114,N_289);
nand U1141 (N_1141,N_79,N_795);
or U1142 (N_1142,N_843,N_847);
or U1143 (N_1143,N_908,N_43);
and U1144 (N_1144,N_577,N_349);
and U1145 (N_1145,N_734,N_705);
or U1146 (N_1146,N_830,N_792);
nand U1147 (N_1147,N_337,N_485);
nand U1148 (N_1148,N_770,N_152);
xor U1149 (N_1149,N_639,N_749);
nor U1150 (N_1150,N_836,N_519);
or U1151 (N_1151,N_979,N_174);
or U1152 (N_1152,N_747,N_324);
nor U1153 (N_1153,N_414,N_551);
nand U1154 (N_1154,N_617,N_160);
nand U1155 (N_1155,N_879,N_752);
nand U1156 (N_1156,N_972,N_71);
or U1157 (N_1157,N_148,N_562);
xnor U1158 (N_1158,N_105,N_748);
or U1159 (N_1159,N_522,N_102);
and U1160 (N_1160,N_21,N_145);
and U1161 (N_1161,N_232,N_881);
nand U1162 (N_1162,N_273,N_601);
nor U1163 (N_1163,N_304,N_371);
nor U1164 (N_1164,N_305,N_344);
xnor U1165 (N_1165,N_523,N_810);
xnor U1166 (N_1166,N_439,N_405);
xor U1167 (N_1167,N_823,N_901);
nand U1168 (N_1168,N_57,N_688);
xor U1169 (N_1169,N_955,N_226);
and U1170 (N_1170,N_651,N_647);
and U1171 (N_1171,N_456,N_713);
and U1172 (N_1172,N_62,N_552);
and U1173 (N_1173,N_194,N_274);
nand U1174 (N_1174,N_913,N_73);
xor U1175 (N_1175,N_116,N_888);
and U1176 (N_1176,N_17,N_430);
nor U1177 (N_1177,N_907,N_533);
xnor U1178 (N_1178,N_862,N_334);
or U1179 (N_1179,N_65,N_55);
nand U1180 (N_1180,N_136,N_898);
xnor U1181 (N_1181,N_851,N_916);
and U1182 (N_1182,N_82,N_931);
nor U1183 (N_1183,N_663,N_156);
nand U1184 (N_1184,N_935,N_178);
nor U1185 (N_1185,N_38,N_966);
xnor U1186 (N_1186,N_623,N_757);
and U1187 (N_1187,N_679,N_309);
or U1188 (N_1188,N_707,N_475);
nor U1189 (N_1189,N_691,N_826);
and U1190 (N_1190,N_258,N_646);
or U1191 (N_1191,N_782,N_119);
xnor U1192 (N_1192,N_350,N_124);
nor U1193 (N_1193,N_677,N_331);
and U1194 (N_1194,N_992,N_446);
nor U1195 (N_1195,N_295,N_802);
or U1196 (N_1196,N_263,N_94);
or U1197 (N_1197,N_775,N_650);
or U1198 (N_1198,N_231,N_824);
nand U1199 (N_1199,N_242,N_555);
nor U1200 (N_1200,N_896,N_883);
and U1201 (N_1201,N_134,N_808);
and U1202 (N_1202,N_937,N_809);
and U1203 (N_1203,N_128,N_358);
nand U1204 (N_1204,N_827,N_339);
xnor U1205 (N_1205,N_270,N_297);
or U1206 (N_1206,N_120,N_77);
nand U1207 (N_1207,N_696,N_489);
nand U1208 (N_1208,N_106,N_479);
nand U1209 (N_1209,N_396,N_799);
xor U1210 (N_1210,N_975,N_821);
and U1211 (N_1211,N_662,N_661);
xnor U1212 (N_1212,N_658,N_35);
xnor U1213 (N_1213,N_938,N_813);
xor U1214 (N_1214,N_946,N_912);
nor U1215 (N_1215,N_72,N_130);
and U1216 (N_1216,N_96,N_112);
or U1217 (N_1217,N_718,N_25);
nand U1218 (N_1218,N_854,N_591);
nor U1219 (N_1219,N_151,N_728);
xnor U1220 (N_1220,N_473,N_785);
nand U1221 (N_1221,N_498,N_675);
nand U1222 (N_1222,N_517,N_741);
and U1223 (N_1223,N_631,N_406);
nand U1224 (N_1224,N_153,N_528);
nand U1225 (N_1225,N_815,N_336);
nor U1226 (N_1226,N_542,N_507);
xor U1227 (N_1227,N_490,N_720);
nor U1228 (N_1228,N_667,N_78);
or U1229 (N_1229,N_431,N_225);
and U1230 (N_1230,N_855,N_882);
xnor U1231 (N_1231,N_192,N_207);
and U1232 (N_1232,N_125,N_902);
or U1233 (N_1233,N_402,N_803);
nand U1234 (N_1234,N_666,N_64);
nor U1235 (N_1235,N_277,N_947);
or U1236 (N_1236,N_228,N_587);
and U1237 (N_1237,N_745,N_169);
and U1238 (N_1238,N_204,N_13);
nor U1239 (N_1239,N_154,N_746);
nand U1240 (N_1240,N_950,N_333);
or U1241 (N_1241,N_763,N_90);
nor U1242 (N_1242,N_367,N_33);
or U1243 (N_1243,N_172,N_794);
nand U1244 (N_1244,N_196,N_321);
nor U1245 (N_1245,N_941,N_986);
nand U1246 (N_1246,N_714,N_300);
nand U1247 (N_1247,N_302,N_876);
xnor U1248 (N_1248,N_469,N_463);
or U1249 (N_1249,N_529,N_872);
xor U1250 (N_1250,N_515,N_253);
or U1251 (N_1251,N_996,N_583);
and U1252 (N_1252,N_870,N_924);
or U1253 (N_1253,N_754,N_772);
nor U1254 (N_1254,N_723,N_190);
nor U1255 (N_1255,N_822,N_701);
or U1256 (N_1256,N_973,N_797);
nand U1257 (N_1257,N_361,N_725);
or U1258 (N_1258,N_132,N_382);
xnor U1259 (N_1259,N_566,N_534);
and U1260 (N_1260,N_131,N_880);
xnor U1261 (N_1261,N_780,N_175);
or U1262 (N_1262,N_953,N_709);
nand U1263 (N_1263,N_499,N_14);
or U1264 (N_1264,N_217,N_370);
nor U1265 (N_1265,N_203,N_149);
xnor U1266 (N_1266,N_218,N_238);
nor U1267 (N_1267,N_91,N_990);
xor U1268 (N_1268,N_932,N_859);
or U1269 (N_1269,N_920,N_581);
xor U1270 (N_1270,N_622,N_954);
nand U1271 (N_1271,N_742,N_500);
nor U1272 (N_1272,N_607,N_416);
xor U1273 (N_1273,N_518,N_150);
or U1274 (N_1274,N_139,N_956);
nand U1275 (N_1275,N_670,N_271);
nor U1276 (N_1276,N_766,N_615);
nand U1277 (N_1277,N_272,N_657);
and U1278 (N_1278,N_874,N_539);
and U1279 (N_1279,N_989,N_428);
nand U1280 (N_1280,N_710,N_262);
or U1281 (N_1281,N_243,N_467);
xor U1282 (N_1282,N_627,N_308);
or U1283 (N_1283,N_5,N_214);
xor U1284 (N_1284,N_694,N_969);
or U1285 (N_1285,N_513,N_411);
or U1286 (N_1286,N_374,N_462);
nand U1287 (N_1287,N_461,N_635);
and U1288 (N_1288,N_761,N_995);
and U1289 (N_1289,N_159,N_629);
nand U1290 (N_1290,N_355,N_804);
or U1291 (N_1291,N_957,N_739);
nor U1292 (N_1292,N_380,N_493);
xnor U1293 (N_1293,N_759,N_286);
and U1294 (N_1294,N_144,N_385);
xor U1295 (N_1295,N_260,N_264);
and U1296 (N_1296,N_56,N_676);
xor U1297 (N_1297,N_744,N_837);
and U1298 (N_1298,N_373,N_877);
xor U1299 (N_1299,N_588,N_418);
and U1300 (N_1300,N_921,N_18);
or U1301 (N_1301,N_450,N_140);
or U1302 (N_1302,N_437,N_531);
xor U1303 (N_1303,N_549,N_841);
nor U1304 (N_1304,N_395,N_394);
and U1305 (N_1305,N_865,N_413);
or U1306 (N_1306,N_267,N_60);
nor U1307 (N_1307,N_768,N_81);
nand U1308 (N_1308,N_497,N_213);
and U1309 (N_1309,N_584,N_70);
and U1310 (N_1310,N_943,N_455);
xnor U1311 (N_1311,N_825,N_906);
nor U1312 (N_1312,N_440,N_998);
nand U1313 (N_1313,N_944,N_680);
nor U1314 (N_1314,N_624,N_12);
or U1315 (N_1315,N_419,N_483);
xor U1316 (N_1316,N_829,N_384);
or U1317 (N_1317,N_630,N_233);
and U1318 (N_1318,N_216,N_168);
or U1319 (N_1319,N_375,N_977);
nand U1320 (N_1320,N_386,N_209);
or U1321 (N_1321,N_442,N_988);
or U1322 (N_1322,N_724,N_560);
nand U1323 (N_1323,N_838,N_963);
xnor U1324 (N_1324,N_695,N_571);
xnor U1325 (N_1325,N_162,N_928);
xor U1326 (N_1326,N_698,N_237);
nand U1327 (N_1327,N_726,N_968);
and U1328 (N_1328,N_328,N_230);
nor U1329 (N_1329,N_451,N_678);
and U1330 (N_1330,N_994,N_641);
xor U1331 (N_1331,N_99,N_819);
nor U1332 (N_1332,N_645,N_934);
nand U1333 (N_1333,N_762,N_256);
nand U1334 (N_1334,N_925,N_100);
nor U1335 (N_1335,N_496,N_407);
or U1336 (N_1336,N_255,N_787);
nor U1337 (N_1337,N_983,N_885);
xnor U1338 (N_1338,N_790,N_509);
nor U1339 (N_1339,N_796,N_806);
and U1340 (N_1340,N_84,N_590);
or U1341 (N_1341,N_502,N_535);
nor U1342 (N_1342,N_241,N_351);
xor U1343 (N_1343,N_354,N_997);
or U1344 (N_1344,N_637,N_580);
nor U1345 (N_1345,N_598,N_512);
xor U1346 (N_1346,N_781,N_738);
nor U1347 (N_1347,N_466,N_261);
nor U1348 (N_1348,N_632,N_890);
and U1349 (N_1349,N_452,N_952);
xor U1350 (N_1350,N_275,N_722);
or U1351 (N_1351,N_634,N_684);
xnor U1352 (N_1352,N_900,N_845);
or U1353 (N_1353,N_76,N_812);
nand U1354 (N_1354,N_15,N_41);
xnor U1355 (N_1355,N_923,N_625);
and U1356 (N_1356,N_141,N_180);
or U1357 (N_1357,N_683,N_191);
and U1358 (N_1358,N_961,N_835);
nor U1359 (N_1359,N_915,N_905);
nor U1360 (N_1360,N_235,N_506);
xor U1361 (N_1361,N_914,N_188);
nand U1362 (N_1362,N_579,N_516);
nand U1363 (N_1363,N_546,N_648);
or U1364 (N_1364,N_183,N_572);
or U1365 (N_1365,N_47,N_109);
nor U1366 (N_1366,N_919,N_597);
or U1367 (N_1367,N_840,N_578);
xnor U1368 (N_1368,N_976,N_807);
nand U1369 (N_1369,N_736,N_457);
or U1370 (N_1370,N_381,N_254);
and U1371 (N_1371,N_917,N_312);
xnor U1372 (N_1372,N_24,N_435);
nand U1373 (N_1373,N_700,N_39);
nand U1374 (N_1374,N_687,N_816);
nand U1375 (N_1375,N_771,N_540);
nand U1376 (N_1376,N_732,N_669);
and U1377 (N_1377,N_74,N_959);
nor U1378 (N_1378,N_32,N_290);
and U1379 (N_1379,N_970,N_834);
nand U1380 (N_1380,N_778,N_68);
xnor U1381 (N_1381,N_147,N_706);
and U1382 (N_1382,N_284,N_129);
and U1383 (N_1383,N_731,N_764);
xor U1384 (N_1384,N_948,N_936);
nor U1385 (N_1385,N_472,N_564);
nor U1386 (N_1386,N_727,N_458);
or U1387 (N_1387,N_532,N_332);
and U1388 (N_1388,N_50,N_945);
xnor U1389 (N_1389,N_735,N_98);
and U1390 (N_1390,N_541,N_287);
nand U1391 (N_1391,N_37,N_538);
nand U1392 (N_1392,N_962,N_36);
and U1393 (N_1393,N_441,N_904);
nand U1394 (N_1394,N_980,N_958);
or U1395 (N_1395,N_346,N_30);
nand U1396 (N_1396,N_427,N_495);
xnor U1397 (N_1397,N_342,N_711);
nand U1398 (N_1398,N_58,N_993);
or U1399 (N_1399,N_89,N_703);
nor U1400 (N_1400,N_364,N_387);
or U1401 (N_1401,N_365,N_453);
xor U1402 (N_1402,N_279,N_614);
or U1403 (N_1403,N_66,N_377);
nor U1404 (N_1404,N_186,N_610);
xnor U1405 (N_1405,N_193,N_814);
or U1406 (N_1406,N_176,N_960);
nor U1407 (N_1407,N_715,N_909);
xnor U1408 (N_1408,N_401,N_101);
xnor U1409 (N_1409,N_573,N_878);
or U1410 (N_1410,N_424,N_199);
or U1411 (N_1411,N_831,N_478);
and U1412 (N_1412,N_576,N_717);
nor U1413 (N_1413,N_283,N_893);
nand U1414 (N_1414,N_487,N_567);
or U1415 (N_1415,N_299,N_93);
or U1416 (N_1416,N_868,N_556);
or U1417 (N_1417,N_999,N_820);
or U1418 (N_1418,N_987,N_127);
nand U1419 (N_1419,N_818,N_737);
and U1420 (N_1420,N_927,N_185);
and U1421 (N_1421,N_699,N_397);
nor U1422 (N_1422,N_654,N_86);
and U1423 (N_1423,N_118,N_536);
xnor U1424 (N_1424,N_653,N_447);
and U1425 (N_1425,N_852,N_392);
and U1426 (N_1426,N_356,N_121);
nand U1427 (N_1427,N_234,N_740);
nand U1428 (N_1428,N_606,N_789);
nor U1429 (N_1429,N_933,N_638);
nor U1430 (N_1430,N_751,N_222);
nand U1431 (N_1431,N_445,N_388);
or U1432 (N_1432,N_34,N_480);
or U1433 (N_1433,N_390,N_864);
or U1434 (N_1434,N_417,N_11);
nor U1435 (N_1435,N_773,N_828);
or U1436 (N_1436,N_574,N_899);
or U1437 (N_1437,N_281,N_404);
and U1438 (N_1438,N_791,N_690);
nor U1439 (N_1439,N_389,N_853);
xor U1440 (N_1440,N_758,N_750);
and U1441 (N_1441,N_7,N_668);
nor U1442 (N_1442,N_359,N_223);
or U1443 (N_1443,N_784,N_88);
and U1444 (N_1444,N_59,N_326);
and U1445 (N_1445,N_595,N_250);
nand U1446 (N_1446,N_476,N_660);
and U1447 (N_1447,N_215,N_889);
and U1448 (N_1448,N_547,N_369);
and U1449 (N_1449,N_292,N_801);
or U1450 (N_1450,N_307,N_605);
xor U1451 (N_1451,N_266,N_206);
nor U1452 (N_1452,N_158,N_978);
nand U1453 (N_1453,N_163,N_842);
nand U1454 (N_1454,N_426,N_166);
nand U1455 (N_1455,N_525,N_236);
and U1456 (N_1456,N_719,N_964);
nor U1457 (N_1457,N_603,N_671);
nand U1458 (N_1458,N_425,N_800);
nor U1459 (N_1459,N_655,N_604);
and U1460 (N_1460,N_561,N_774);
or U1461 (N_1461,N_857,N_391);
xnor U1462 (N_1462,N_494,N_249);
nor U1463 (N_1463,N_345,N_195);
xor U1464 (N_1464,N_860,N_8);
nand U1465 (N_1465,N_244,N_470);
nor U1466 (N_1466,N_340,N_702);
xor U1467 (N_1467,N_20,N_360);
or U1468 (N_1468,N_239,N_848);
xor U1469 (N_1469,N_319,N_508);
nand U1470 (N_1470,N_173,N_103);
or U1471 (N_1471,N_594,N_686);
xor U1472 (N_1472,N_16,N_570);
or U1473 (N_1473,N_596,N_259);
or U1474 (N_1474,N_991,N_423);
or U1475 (N_1475,N_559,N_198);
nor U1476 (N_1476,N_918,N_4);
or U1477 (N_1477,N_293,N_940);
or U1478 (N_1478,N_229,N_582);
or U1479 (N_1479,N_51,N_69);
nand U1480 (N_1480,N_543,N_443);
nand U1481 (N_1481,N_170,N_642);
nand U1482 (N_1482,N_665,N_612);
nor U1483 (N_1483,N_524,N_201);
or U1484 (N_1484,N_755,N_484);
nand U1485 (N_1485,N_10,N_545);
xnor U1486 (N_1486,N_585,N_104);
nor U1487 (N_1487,N_492,N_674);
nand U1488 (N_1488,N_410,N_313);
and U1489 (N_1489,N_245,N_811);
xnor U1490 (N_1490,N_644,N_92);
and U1491 (N_1491,N_537,N_729);
or U1492 (N_1492,N_278,N_673);
nand U1493 (N_1493,N_930,N_503);
and U1494 (N_1494,N_189,N_205);
nand U1495 (N_1495,N_44,N_184);
xnor U1496 (N_1496,N_137,N_875);
nor U1497 (N_1497,N_608,N_276);
nand U1498 (N_1498,N_530,N_891);
and U1499 (N_1499,N_247,N_833);
nand U1500 (N_1500,N_842,N_981);
or U1501 (N_1501,N_803,N_239);
and U1502 (N_1502,N_83,N_882);
xor U1503 (N_1503,N_551,N_536);
or U1504 (N_1504,N_855,N_962);
nand U1505 (N_1505,N_24,N_966);
xnor U1506 (N_1506,N_912,N_309);
nor U1507 (N_1507,N_818,N_276);
nor U1508 (N_1508,N_75,N_63);
and U1509 (N_1509,N_680,N_932);
nor U1510 (N_1510,N_842,N_627);
nor U1511 (N_1511,N_210,N_854);
xnor U1512 (N_1512,N_730,N_479);
nor U1513 (N_1513,N_909,N_524);
nor U1514 (N_1514,N_109,N_143);
or U1515 (N_1515,N_903,N_933);
xnor U1516 (N_1516,N_135,N_830);
and U1517 (N_1517,N_652,N_369);
xnor U1518 (N_1518,N_346,N_75);
nand U1519 (N_1519,N_757,N_204);
nand U1520 (N_1520,N_419,N_707);
and U1521 (N_1521,N_994,N_92);
nor U1522 (N_1522,N_273,N_883);
xnor U1523 (N_1523,N_705,N_382);
xnor U1524 (N_1524,N_363,N_825);
nand U1525 (N_1525,N_205,N_431);
nand U1526 (N_1526,N_580,N_308);
or U1527 (N_1527,N_66,N_326);
nand U1528 (N_1528,N_49,N_781);
nor U1529 (N_1529,N_109,N_706);
nand U1530 (N_1530,N_373,N_651);
and U1531 (N_1531,N_861,N_212);
or U1532 (N_1532,N_375,N_141);
xor U1533 (N_1533,N_885,N_463);
nand U1534 (N_1534,N_165,N_297);
nand U1535 (N_1535,N_840,N_773);
nor U1536 (N_1536,N_702,N_629);
xnor U1537 (N_1537,N_557,N_995);
and U1538 (N_1538,N_447,N_69);
or U1539 (N_1539,N_660,N_855);
xnor U1540 (N_1540,N_863,N_898);
and U1541 (N_1541,N_740,N_980);
nor U1542 (N_1542,N_100,N_271);
nand U1543 (N_1543,N_410,N_25);
nand U1544 (N_1544,N_660,N_260);
and U1545 (N_1545,N_382,N_206);
xor U1546 (N_1546,N_462,N_275);
or U1547 (N_1547,N_130,N_365);
nor U1548 (N_1548,N_600,N_324);
nand U1549 (N_1549,N_713,N_760);
nand U1550 (N_1550,N_185,N_26);
nand U1551 (N_1551,N_209,N_955);
xnor U1552 (N_1552,N_338,N_559);
nor U1553 (N_1553,N_726,N_674);
nor U1554 (N_1554,N_695,N_39);
nand U1555 (N_1555,N_516,N_345);
nand U1556 (N_1556,N_843,N_667);
and U1557 (N_1557,N_412,N_697);
nor U1558 (N_1558,N_380,N_79);
nor U1559 (N_1559,N_144,N_916);
nor U1560 (N_1560,N_741,N_732);
or U1561 (N_1561,N_447,N_251);
nand U1562 (N_1562,N_297,N_365);
nor U1563 (N_1563,N_418,N_623);
xnor U1564 (N_1564,N_255,N_244);
nand U1565 (N_1565,N_734,N_226);
xnor U1566 (N_1566,N_891,N_705);
and U1567 (N_1567,N_28,N_812);
nand U1568 (N_1568,N_293,N_649);
and U1569 (N_1569,N_543,N_758);
xnor U1570 (N_1570,N_157,N_241);
nand U1571 (N_1571,N_133,N_655);
xnor U1572 (N_1572,N_677,N_510);
and U1573 (N_1573,N_95,N_64);
and U1574 (N_1574,N_793,N_706);
and U1575 (N_1575,N_904,N_421);
or U1576 (N_1576,N_294,N_543);
nand U1577 (N_1577,N_803,N_585);
nand U1578 (N_1578,N_125,N_384);
nand U1579 (N_1579,N_984,N_396);
and U1580 (N_1580,N_221,N_438);
nand U1581 (N_1581,N_62,N_201);
xnor U1582 (N_1582,N_626,N_711);
or U1583 (N_1583,N_562,N_440);
or U1584 (N_1584,N_449,N_276);
nor U1585 (N_1585,N_300,N_643);
nor U1586 (N_1586,N_802,N_316);
xor U1587 (N_1587,N_10,N_58);
nand U1588 (N_1588,N_48,N_224);
nor U1589 (N_1589,N_31,N_673);
xnor U1590 (N_1590,N_598,N_544);
nor U1591 (N_1591,N_105,N_765);
or U1592 (N_1592,N_76,N_771);
nor U1593 (N_1593,N_136,N_135);
nand U1594 (N_1594,N_309,N_219);
and U1595 (N_1595,N_334,N_532);
nand U1596 (N_1596,N_79,N_417);
nor U1597 (N_1597,N_127,N_241);
or U1598 (N_1598,N_135,N_451);
or U1599 (N_1599,N_504,N_244);
xnor U1600 (N_1600,N_313,N_162);
nor U1601 (N_1601,N_656,N_26);
and U1602 (N_1602,N_170,N_656);
xor U1603 (N_1603,N_793,N_110);
xor U1604 (N_1604,N_457,N_721);
nand U1605 (N_1605,N_175,N_146);
nand U1606 (N_1606,N_119,N_44);
xor U1607 (N_1607,N_673,N_104);
nor U1608 (N_1608,N_671,N_82);
nand U1609 (N_1609,N_188,N_902);
or U1610 (N_1610,N_648,N_820);
xnor U1611 (N_1611,N_861,N_724);
nand U1612 (N_1612,N_841,N_71);
nand U1613 (N_1613,N_288,N_163);
xor U1614 (N_1614,N_283,N_168);
and U1615 (N_1615,N_809,N_555);
and U1616 (N_1616,N_122,N_304);
nor U1617 (N_1617,N_573,N_344);
xor U1618 (N_1618,N_981,N_102);
and U1619 (N_1619,N_596,N_151);
nor U1620 (N_1620,N_31,N_156);
xor U1621 (N_1621,N_406,N_309);
nand U1622 (N_1622,N_689,N_987);
nand U1623 (N_1623,N_401,N_253);
nand U1624 (N_1624,N_825,N_916);
nor U1625 (N_1625,N_699,N_799);
and U1626 (N_1626,N_615,N_199);
or U1627 (N_1627,N_885,N_52);
and U1628 (N_1628,N_479,N_286);
xnor U1629 (N_1629,N_781,N_564);
nor U1630 (N_1630,N_88,N_462);
nand U1631 (N_1631,N_882,N_600);
xor U1632 (N_1632,N_104,N_506);
and U1633 (N_1633,N_213,N_9);
xor U1634 (N_1634,N_603,N_5);
or U1635 (N_1635,N_18,N_584);
xor U1636 (N_1636,N_173,N_952);
xnor U1637 (N_1637,N_818,N_211);
and U1638 (N_1638,N_161,N_197);
nor U1639 (N_1639,N_395,N_581);
and U1640 (N_1640,N_353,N_620);
nand U1641 (N_1641,N_298,N_180);
nor U1642 (N_1642,N_164,N_692);
or U1643 (N_1643,N_527,N_182);
and U1644 (N_1644,N_833,N_765);
nor U1645 (N_1645,N_715,N_680);
or U1646 (N_1646,N_648,N_25);
and U1647 (N_1647,N_510,N_306);
and U1648 (N_1648,N_209,N_101);
and U1649 (N_1649,N_26,N_225);
nor U1650 (N_1650,N_350,N_775);
xnor U1651 (N_1651,N_808,N_425);
nand U1652 (N_1652,N_926,N_762);
or U1653 (N_1653,N_220,N_491);
nor U1654 (N_1654,N_264,N_189);
nand U1655 (N_1655,N_857,N_480);
and U1656 (N_1656,N_584,N_869);
xnor U1657 (N_1657,N_963,N_50);
nor U1658 (N_1658,N_272,N_961);
or U1659 (N_1659,N_35,N_287);
and U1660 (N_1660,N_771,N_900);
or U1661 (N_1661,N_942,N_115);
and U1662 (N_1662,N_872,N_468);
or U1663 (N_1663,N_294,N_902);
nor U1664 (N_1664,N_730,N_577);
nand U1665 (N_1665,N_537,N_429);
xor U1666 (N_1666,N_673,N_930);
nor U1667 (N_1667,N_314,N_373);
and U1668 (N_1668,N_575,N_568);
xor U1669 (N_1669,N_121,N_834);
nand U1670 (N_1670,N_619,N_630);
or U1671 (N_1671,N_235,N_807);
nor U1672 (N_1672,N_287,N_621);
nand U1673 (N_1673,N_175,N_918);
and U1674 (N_1674,N_510,N_197);
and U1675 (N_1675,N_784,N_67);
or U1676 (N_1676,N_55,N_229);
xnor U1677 (N_1677,N_589,N_479);
or U1678 (N_1678,N_198,N_412);
nand U1679 (N_1679,N_173,N_588);
and U1680 (N_1680,N_653,N_679);
and U1681 (N_1681,N_578,N_581);
or U1682 (N_1682,N_416,N_443);
or U1683 (N_1683,N_52,N_909);
or U1684 (N_1684,N_95,N_863);
xor U1685 (N_1685,N_388,N_394);
nor U1686 (N_1686,N_869,N_782);
nor U1687 (N_1687,N_528,N_926);
nor U1688 (N_1688,N_925,N_378);
nor U1689 (N_1689,N_162,N_576);
nor U1690 (N_1690,N_776,N_950);
or U1691 (N_1691,N_331,N_28);
and U1692 (N_1692,N_571,N_362);
or U1693 (N_1693,N_44,N_411);
nand U1694 (N_1694,N_912,N_848);
nor U1695 (N_1695,N_273,N_724);
nand U1696 (N_1696,N_728,N_398);
xnor U1697 (N_1697,N_574,N_959);
nand U1698 (N_1698,N_69,N_318);
or U1699 (N_1699,N_886,N_476);
nor U1700 (N_1700,N_396,N_568);
xnor U1701 (N_1701,N_956,N_539);
nand U1702 (N_1702,N_215,N_450);
nor U1703 (N_1703,N_79,N_158);
nor U1704 (N_1704,N_335,N_698);
xor U1705 (N_1705,N_297,N_839);
and U1706 (N_1706,N_107,N_717);
or U1707 (N_1707,N_146,N_996);
or U1708 (N_1708,N_738,N_903);
nand U1709 (N_1709,N_881,N_408);
nand U1710 (N_1710,N_626,N_407);
and U1711 (N_1711,N_232,N_242);
xor U1712 (N_1712,N_209,N_62);
xnor U1713 (N_1713,N_815,N_690);
or U1714 (N_1714,N_157,N_76);
nor U1715 (N_1715,N_494,N_655);
or U1716 (N_1716,N_803,N_789);
or U1717 (N_1717,N_570,N_551);
and U1718 (N_1718,N_882,N_488);
or U1719 (N_1719,N_352,N_856);
nor U1720 (N_1720,N_179,N_116);
xor U1721 (N_1721,N_310,N_385);
nand U1722 (N_1722,N_318,N_497);
nor U1723 (N_1723,N_151,N_243);
or U1724 (N_1724,N_565,N_827);
xnor U1725 (N_1725,N_595,N_499);
nand U1726 (N_1726,N_340,N_989);
xnor U1727 (N_1727,N_104,N_979);
and U1728 (N_1728,N_473,N_424);
nand U1729 (N_1729,N_402,N_486);
or U1730 (N_1730,N_949,N_886);
or U1731 (N_1731,N_817,N_974);
or U1732 (N_1732,N_307,N_264);
nand U1733 (N_1733,N_403,N_500);
xor U1734 (N_1734,N_189,N_98);
xnor U1735 (N_1735,N_606,N_101);
nand U1736 (N_1736,N_458,N_754);
nor U1737 (N_1737,N_208,N_201);
nand U1738 (N_1738,N_291,N_292);
and U1739 (N_1739,N_455,N_966);
xor U1740 (N_1740,N_271,N_423);
and U1741 (N_1741,N_926,N_763);
nand U1742 (N_1742,N_249,N_151);
or U1743 (N_1743,N_19,N_495);
nor U1744 (N_1744,N_821,N_948);
or U1745 (N_1745,N_996,N_798);
nor U1746 (N_1746,N_638,N_98);
nand U1747 (N_1747,N_366,N_826);
and U1748 (N_1748,N_331,N_586);
nor U1749 (N_1749,N_481,N_701);
or U1750 (N_1750,N_989,N_610);
xor U1751 (N_1751,N_161,N_293);
xnor U1752 (N_1752,N_103,N_442);
xor U1753 (N_1753,N_231,N_158);
and U1754 (N_1754,N_395,N_366);
nor U1755 (N_1755,N_587,N_546);
and U1756 (N_1756,N_243,N_494);
nand U1757 (N_1757,N_955,N_845);
nor U1758 (N_1758,N_567,N_780);
nand U1759 (N_1759,N_458,N_503);
or U1760 (N_1760,N_792,N_577);
xnor U1761 (N_1761,N_917,N_465);
and U1762 (N_1762,N_270,N_105);
nor U1763 (N_1763,N_645,N_586);
or U1764 (N_1764,N_516,N_436);
and U1765 (N_1765,N_261,N_165);
or U1766 (N_1766,N_952,N_14);
nor U1767 (N_1767,N_132,N_273);
nand U1768 (N_1768,N_795,N_674);
and U1769 (N_1769,N_427,N_487);
nor U1770 (N_1770,N_489,N_471);
nor U1771 (N_1771,N_693,N_411);
xor U1772 (N_1772,N_197,N_488);
and U1773 (N_1773,N_523,N_789);
xor U1774 (N_1774,N_910,N_813);
or U1775 (N_1775,N_151,N_443);
xor U1776 (N_1776,N_334,N_130);
or U1777 (N_1777,N_815,N_244);
nor U1778 (N_1778,N_772,N_155);
or U1779 (N_1779,N_105,N_46);
nor U1780 (N_1780,N_61,N_107);
and U1781 (N_1781,N_570,N_780);
and U1782 (N_1782,N_727,N_918);
nor U1783 (N_1783,N_816,N_241);
and U1784 (N_1784,N_879,N_367);
nand U1785 (N_1785,N_831,N_456);
nor U1786 (N_1786,N_622,N_558);
nand U1787 (N_1787,N_26,N_130);
and U1788 (N_1788,N_631,N_891);
and U1789 (N_1789,N_189,N_584);
or U1790 (N_1790,N_701,N_968);
nand U1791 (N_1791,N_779,N_798);
or U1792 (N_1792,N_780,N_863);
nand U1793 (N_1793,N_346,N_870);
nand U1794 (N_1794,N_142,N_885);
and U1795 (N_1795,N_752,N_500);
or U1796 (N_1796,N_864,N_433);
or U1797 (N_1797,N_89,N_294);
or U1798 (N_1798,N_4,N_392);
or U1799 (N_1799,N_792,N_307);
or U1800 (N_1800,N_109,N_324);
or U1801 (N_1801,N_980,N_599);
nand U1802 (N_1802,N_118,N_207);
xor U1803 (N_1803,N_436,N_620);
xor U1804 (N_1804,N_176,N_592);
and U1805 (N_1805,N_181,N_704);
and U1806 (N_1806,N_703,N_401);
and U1807 (N_1807,N_553,N_977);
or U1808 (N_1808,N_367,N_939);
xnor U1809 (N_1809,N_441,N_935);
nor U1810 (N_1810,N_484,N_223);
xnor U1811 (N_1811,N_879,N_888);
nor U1812 (N_1812,N_221,N_377);
xnor U1813 (N_1813,N_385,N_882);
or U1814 (N_1814,N_280,N_762);
nor U1815 (N_1815,N_632,N_777);
or U1816 (N_1816,N_988,N_523);
nor U1817 (N_1817,N_555,N_813);
nand U1818 (N_1818,N_797,N_389);
nor U1819 (N_1819,N_553,N_618);
nor U1820 (N_1820,N_267,N_75);
nand U1821 (N_1821,N_440,N_827);
and U1822 (N_1822,N_269,N_176);
and U1823 (N_1823,N_875,N_460);
xor U1824 (N_1824,N_238,N_836);
xnor U1825 (N_1825,N_619,N_622);
nand U1826 (N_1826,N_838,N_674);
xnor U1827 (N_1827,N_364,N_572);
xnor U1828 (N_1828,N_570,N_274);
or U1829 (N_1829,N_262,N_314);
nand U1830 (N_1830,N_665,N_821);
nand U1831 (N_1831,N_688,N_115);
or U1832 (N_1832,N_902,N_407);
nor U1833 (N_1833,N_158,N_46);
nor U1834 (N_1834,N_585,N_880);
and U1835 (N_1835,N_207,N_429);
nor U1836 (N_1836,N_305,N_607);
nor U1837 (N_1837,N_348,N_794);
nand U1838 (N_1838,N_21,N_91);
and U1839 (N_1839,N_40,N_78);
or U1840 (N_1840,N_515,N_107);
and U1841 (N_1841,N_224,N_742);
or U1842 (N_1842,N_548,N_60);
nand U1843 (N_1843,N_381,N_975);
and U1844 (N_1844,N_0,N_354);
xor U1845 (N_1845,N_370,N_315);
xor U1846 (N_1846,N_990,N_550);
and U1847 (N_1847,N_730,N_386);
nor U1848 (N_1848,N_416,N_274);
nand U1849 (N_1849,N_389,N_253);
and U1850 (N_1850,N_303,N_359);
or U1851 (N_1851,N_900,N_678);
xnor U1852 (N_1852,N_428,N_837);
xnor U1853 (N_1853,N_27,N_39);
xor U1854 (N_1854,N_133,N_351);
nor U1855 (N_1855,N_241,N_827);
or U1856 (N_1856,N_663,N_70);
or U1857 (N_1857,N_352,N_912);
and U1858 (N_1858,N_878,N_4);
nor U1859 (N_1859,N_255,N_901);
xnor U1860 (N_1860,N_730,N_65);
nor U1861 (N_1861,N_457,N_680);
nor U1862 (N_1862,N_980,N_881);
nor U1863 (N_1863,N_68,N_446);
nor U1864 (N_1864,N_42,N_436);
and U1865 (N_1865,N_936,N_870);
nor U1866 (N_1866,N_188,N_808);
and U1867 (N_1867,N_163,N_669);
nand U1868 (N_1868,N_690,N_981);
xnor U1869 (N_1869,N_590,N_536);
nand U1870 (N_1870,N_560,N_153);
and U1871 (N_1871,N_324,N_981);
and U1872 (N_1872,N_314,N_841);
nand U1873 (N_1873,N_395,N_479);
nor U1874 (N_1874,N_0,N_364);
nand U1875 (N_1875,N_553,N_13);
or U1876 (N_1876,N_216,N_612);
xnor U1877 (N_1877,N_179,N_395);
xnor U1878 (N_1878,N_440,N_452);
xor U1879 (N_1879,N_175,N_216);
and U1880 (N_1880,N_483,N_359);
or U1881 (N_1881,N_758,N_541);
nand U1882 (N_1882,N_443,N_379);
or U1883 (N_1883,N_883,N_441);
nand U1884 (N_1884,N_346,N_335);
nand U1885 (N_1885,N_340,N_402);
and U1886 (N_1886,N_44,N_376);
or U1887 (N_1887,N_452,N_495);
nand U1888 (N_1888,N_486,N_790);
or U1889 (N_1889,N_549,N_50);
xnor U1890 (N_1890,N_22,N_175);
xnor U1891 (N_1891,N_26,N_864);
nor U1892 (N_1892,N_637,N_689);
nand U1893 (N_1893,N_266,N_760);
xor U1894 (N_1894,N_620,N_502);
and U1895 (N_1895,N_424,N_998);
or U1896 (N_1896,N_165,N_877);
and U1897 (N_1897,N_296,N_287);
xor U1898 (N_1898,N_932,N_220);
xor U1899 (N_1899,N_919,N_231);
or U1900 (N_1900,N_156,N_815);
xnor U1901 (N_1901,N_205,N_20);
nor U1902 (N_1902,N_814,N_305);
and U1903 (N_1903,N_929,N_133);
nand U1904 (N_1904,N_262,N_291);
xor U1905 (N_1905,N_684,N_315);
nor U1906 (N_1906,N_827,N_937);
nand U1907 (N_1907,N_885,N_948);
and U1908 (N_1908,N_950,N_530);
or U1909 (N_1909,N_334,N_710);
or U1910 (N_1910,N_193,N_453);
nand U1911 (N_1911,N_137,N_920);
and U1912 (N_1912,N_373,N_337);
nor U1913 (N_1913,N_224,N_626);
xnor U1914 (N_1914,N_370,N_612);
and U1915 (N_1915,N_851,N_92);
or U1916 (N_1916,N_229,N_513);
nand U1917 (N_1917,N_801,N_201);
and U1918 (N_1918,N_878,N_525);
nand U1919 (N_1919,N_95,N_611);
nand U1920 (N_1920,N_364,N_151);
nand U1921 (N_1921,N_674,N_656);
nor U1922 (N_1922,N_889,N_797);
xor U1923 (N_1923,N_555,N_313);
nor U1924 (N_1924,N_332,N_713);
nand U1925 (N_1925,N_503,N_310);
or U1926 (N_1926,N_347,N_256);
xnor U1927 (N_1927,N_595,N_192);
or U1928 (N_1928,N_85,N_438);
nand U1929 (N_1929,N_550,N_94);
or U1930 (N_1930,N_576,N_301);
nand U1931 (N_1931,N_695,N_323);
or U1932 (N_1932,N_187,N_124);
xnor U1933 (N_1933,N_478,N_55);
xor U1934 (N_1934,N_88,N_905);
nand U1935 (N_1935,N_844,N_369);
xnor U1936 (N_1936,N_430,N_850);
xnor U1937 (N_1937,N_429,N_47);
nor U1938 (N_1938,N_290,N_127);
nand U1939 (N_1939,N_646,N_189);
or U1940 (N_1940,N_651,N_332);
and U1941 (N_1941,N_981,N_299);
and U1942 (N_1942,N_999,N_815);
xnor U1943 (N_1943,N_842,N_169);
xor U1944 (N_1944,N_702,N_936);
xnor U1945 (N_1945,N_121,N_420);
nand U1946 (N_1946,N_21,N_652);
or U1947 (N_1947,N_768,N_865);
or U1948 (N_1948,N_199,N_916);
or U1949 (N_1949,N_711,N_597);
or U1950 (N_1950,N_979,N_492);
or U1951 (N_1951,N_465,N_906);
nor U1952 (N_1952,N_677,N_372);
nor U1953 (N_1953,N_661,N_480);
nor U1954 (N_1954,N_936,N_444);
or U1955 (N_1955,N_469,N_322);
nor U1956 (N_1956,N_633,N_825);
xnor U1957 (N_1957,N_403,N_872);
nand U1958 (N_1958,N_547,N_201);
xor U1959 (N_1959,N_504,N_984);
nand U1960 (N_1960,N_177,N_733);
or U1961 (N_1961,N_789,N_379);
or U1962 (N_1962,N_381,N_910);
or U1963 (N_1963,N_591,N_419);
and U1964 (N_1964,N_607,N_54);
xnor U1965 (N_1965,N_817,N_930);
nor U1966 (N_1966,N_598,N_529);
and U1967 (N_1967,N_393,N_258);
xnor U1968 (N_1968,N_288,N_298);
nand U1969 (N_1969,N_476,N_781);
nand U1970 (N_1970,N_92,N_429);
or U1971 (N_1971,N_301,N_335);
xor U1972 (N_1972,N_124,N_426);
nor U1973 (N_1973,N_972,N_703);
and U1974 (N_1974,N_273,N_181);
xnor U1975 (N_1975,N_320,N_58);
nor U1976 (N_1976,N_754,N_830);
nand U1977 (N_1977,N_747,N_678);
nand U1978 (N_1978,N_778,N_285);
or U1979 (N_1979,N_670,N_70);
xor U1980 (N_1980,N_726,N_105);
nand U1981 (N_1981,N_759,N_957);
nor U1982 (N_1982,N_720,N_924);
or U1983 (N_1983,N_639,N_561);
or U1984 (N_1984,N_552,N_96);
nand U1985 (N_1985,N_148,N_131);
nor U1986 (N_1986,N_182,N_27);
nand U1987 (N_1987,N_325,N_277);
or U1988 (N_1988,N_27,N_824);
or U1989 (N_1989,N_182,N_400);
xnor U1990 (N_1990,N_3,N_321);
nand U1991 (N_1991,N_213,N_602);
or U1992 (N_1992,N_861,N_974);
xor U1993 (N_1993,N_76,N_985);
and U1994 (N_1994,N_40,N_794);
xor U1995 (N_1995,N_46,N_207);
xor U1996 (N_1996,N_170,N_583);
or U1997 (N_1997,N_988,N_658);
or U1998 (N_1998,N_680,N_64);
nand U1999 (N_1999,N_935,N_853);
and U2000 (N_2000,N_1963,N_1949);
xnor U2001 (N_2001,N_1910,N_1466);
nand U2002 (N_2002,N_1587,N_1840);
and U2003 (N_2003,N_1837,N_1340);
or U2004 (N_2004,N_1129,N_1810);
or U2005 (N_2005,N_1369,N_1254);
and U2006 (N_2006,N_1183,N_1990);
or U2007 (N_2007,N_1795,N_1181);
and U2008 (N_2008,N_1833,N_1812);
and U2009 (N_2009,N_1618,N_1332);
or U2010 (N_2010,N_1051,N_1668);
nor U2011 (N_2011,N_1237,N_1649);
and U2012 (N_2012,N_1221,N_1580);
and U2013 (N_2013,N_1718,N_1261);
nor U2014 (N_2014,N_1298,N_1291);
xnor U2015 (N_2015,N_1527,N_1199);
nor U2016 (N_2016,N_1585,N_1776);
nand U2017 (N_2017,N_1364,N_1187);
or U2018 (N_2018,N_1018,N_1617);
nor U2019 (N_2019,N_1371,N_1603);
nor U2020 (N_2020,N_1762,N_1307);
or U2021 (N_2021,N_1893,N_1520);
or U2022 (N_2022,N_1642,N_1176);
nor U2023 (N_2023,N_1194,N_1973);
nand U2024 (N_2024,N_1720,N_1211);
and U2025 (N_2025,N_1442,N_1621);
or U2026 (N_2026,N_1081,N_1447);
and U2027 (N_2027,N_1670,N_1247);
nor U2028 (N_2028,N_1420,N_1785);
nor U2029 (N_2029,N_1547,N_1351);
nor U2030 (N_2030,N_1532,N_1881);
xor U2031 (N_2031,N_1834,N_1700);
nand U2032 (N_2032,N_1461,N_1888);
nor U2033 (N_2033,N_1078,N_1429);
xor U2034 (N_2034,N_1962,N_1132);
nor U2035 (N_2035,N_1573,N_1170);
nand U2036 (N_2036,N_1731,N_1316);
nor U2037 (N_2037,N_1229,N_1948);
and U2038 (N_2038,N_1085,N_1534);
nand U2039 (N_2039,N_1519,N_1412);
nand U2040 (N_2040,N_1468,N_1748);
nor U2041 (N_2041,N_1713,N_1606);
and U2042 (N_2042,N_1958,N_1353);
nor U2043 (N_2043,N_1434,N_1164);
xnor U2044 (N_2044,N_1019,N_1804);
nand U2045 (N_2045,N_1414,N_1568);
or U2046 (N_2046,N_1093,N_1114);
xnor U2047 (N_2047,N_1627,N_1882);
nor U2048 (N_2048,N_1218,N_1441);
and U2049 (N_2049,N_1815,N_1197);
or U2050 (N_2050,N_1146,N_1417);
nand U2051 (N_2051,N_1565,N_1550);
or U2052 (N_2052,N_1913,N_1306);
or U2053 (N_2053,N_1022,N_1438);
xnor U2054 (N_2054,N_1168,N_1667);
nand U2055 (N_2055,N_1428,N_1435);
xnor U2056 (N_2056,N_1163,N_1540);
nand U2057 (N_2057,N_1681,N_1664);
nor U2058 (N_2058,N_1003,N_1781);
or U2059 (N_2059,N_1077,N_1308);
nor U2060 (N_2060,N_1203,N_1122);
xnor U2061 (N_2061,N_1657,N_1450);
nand U2062 (N_2062,N_1905,N_1265);
xor U2063 (N_2063,N_1212,N_1223);
nor U2064 (N_2064,N_1350,N_1270);
or U2065 (N_2065,N_1297,N_1898);
or U2066 (N_2066,N_1522,N_1370);
or U2067 (N_2067,N_1872,N_1766);
nand U2068 (N_2068,N_1752,N_1422);
and U2069 (N_2069,N_1242,N_1038);
and U2070 (N_2070,N_1286,N_1103);
nand U2071 (N_2071,N_1366,N_1994);
or U2072 (N_2072,N_1842,N_1145);
nor U2073 (N_2073,N_1562,N_1043);
xnor U2074 (N_2074,N_1656,N_1460);
and U2075 (N_2075,N_1249,N_1177);
nand U2076 (N_2076,N_1745,N_1880);
or U2077 (N_2077,N_1172,N_1281);
nand U2078 (N_2078,N_1788,N_1065);
xnor U2079 (N_2079,N_1269,N_1282);
nand U2080 (N_2080,N_1822,N_1205);
xor U2081 (N_2081,N_1566,N_1105);
or U2082 (N_2082,N_1467,N_1289);
xor U2083 (N_2083,N_1736,N_1989);
nand U2084 (N_2084,N_1684,N_1464);
xnor U2085 (N_2085,N_1919,N_1941);
and U2086 (N_2086,N_1315,N_1045);
and U2087 (N_2087,N_1650,N_1448);
nor U2088 (N_2088,N_1600,N_1518);
nor U2089 (N_2089,N_1739,N_1292);
nor U2090 (N_2090,N_1426,N_1719);
or U2091 (N_2091,N_1569,N_1789);
and U2092 (N_2092,N_1033,N_1180);
xor U2093 (N_2093,N_1988,N_1488);
nand U2094 (N_2094,N_1692,N_1946);
nor U2095 (N_2095,N_1641,N_1945);
xor U2096 (N_2096,N_1685,N_1452);
or U2097 (N_2097,N_1783,N_1272);
nand U2098 (N_2098,N_1219,N_1920);
or U2099 (N_2099,N_1127,N_1241);
or U2100 (N_2100,N_1537,N_1346);
or U2101 (N_2101,N_1931,N_1126);
and U2102 (N_2102,N_1956,N_1336);
or U2103 (N_2103,N_1407,N_1802);
nor U2104 (N_2104,N_1347,N_1960);
nor U2105 (N_2105,N_1119,N_1267);
or U2106 (N_2106,N_1157,N_1123);
nor U2107 (N_2107,N_1396,N_1144);
or U2108 (N_2108,N_1799,N_1635);
or U2109 (N_2109,N_1139,N_1699);
nor U2110 (N_2110,N_1220,N_1342);
nor U2111 (N_2111,N_1653,N_1208);
nand U2112 (N_2112,N_1302,N_1341);
and U2113 (N_2113,N_1944,N_1884);
nand U2114 (N_2114,N_1938,N_1803);
xor U2115 (N_2115,N_1453,N_1458);
nor U2116 (N_2116,N_1475,N_1849);
xor U2117 (N_2117,N_1026,N_1153);
nand U2118 (N_2118,N_1303,N_1102);
nor U2119 (N_2119,N_1996,N_1034);
and U2120 (N_2120,N_1222,N_1494);
nor U2121 (N_2121,N_1258,N_1143);
xnor U2122 (N_2122,N_1832,N_1375);
nand U2123 (N_2123,N_1597,N_1240);
xnor U2124 (N_2124,N_1362,N_1310);
and U2125 (N_2125,N_1848,N_1069);
xor U2126 (N_2126,N_1521,N_1955);
xnor U2127 (N_2127,N_1546,N_1725);
nor U2128 (N_2128,N_1445,N_1111);
xnor U2129 (N_2129,N_1391,N_1232);
or U2130 (N_2130,N_1735,N_1395);
and U2131 (N_2131,N_1909,N_1638);
or U2132 (N_2132,N_1987,N_1402);
or U2133 (N_2133,N_1980,N_1706);
nor U2134 (N_2134,N_1004,N_1868);
nand U2135 (N_2135,N_1405,N_1190);
xnor U2136 (N_2136,N_1885,N_1869);
or U2137 (N_2137,N_1485,N_1317);
or U2138 (N_2138,N_1064,N_1917);
xor U2139 (N_2139,N_1694,N_1588);
and U2140 (N_2140,N_1673,N_1586);
or U2141 (N_2141,N_1092,N_1490);
nor U2142 (N_2142,N_1818,N_1253);
and U2143 (N_2143,N_1264,N_1554);
nor U2144 (N_2144,N_1551,N_1397);
and U2145 (N_2145,N_1171,N_1155);
xor U2146 (N_2146,N_1054,N_1179);
nor U2147 (N_2147,N_1496,N_1174);
or U2148 (N_2148,N_1708,N_1124);
or U2149 (N_2149,N_1070,N_1000);
and U2150 (N_2150,N_1131,N_1844);
nor U2151 (N_2151,N_1671,N_1952);
or U2152 (N_2152,N_1549,N_1687);
and U2153 (N_2153,N_1437,N_1128);
nand U2154 (N_2154,N_1500,N_1764);
and U2155 (N_2155,N_1552,N_1440);
xnor U2156 (N_2156,N_1196,N_1192);
or U2157 (N_2157,N_1903,N_1021);
nand U2158 (N_2158,N_1243,N_1277);
or U2159 (N_2159,N_1563,N_1830);
and U2160 (N_2160,N_1031,N_1935);
and U2161 (N_2161,N_1011,N_1595);
and U2162 (N_2162,N_1951,N_1792);
xor U2163 (N_2163,N_1697,N_1015);
or U2164 (N_2164,N_1703,N_1978);
and U2165 (N_2165,N_1787,N_1985);
and U2166 (N_2166,N_1716,N_1968);
or U2167 (N_2167,N_1991,N_1487);
xnor U2168 (N_2168,N_1791,N_1099);
nor U2169 (N_2169,N_1060,N_1262);
nor U2170 (N_2170,N_1095,N_1101);
and U2171 (N_2171,N_1016,N_1614);
and U2172 (N_2172,N_1579,N_1071);
xnor U2173 (N_2173,N_1106,N_1999);
nand U2174 (N_2174,N_1189,N_1930);
nor U2175 (N_2175,N_1309,N_1966);
nand U2176 (N_2176,N_1936,N_1782);
nor U2177 (N_2177,N_1418,N_1294);
xor U2178 (N_2178,N_1098,N_1775);
nor U2179 (N_2179,N_1864,N_1046);
or U2180 (N_2180,N_1471,N_1423);
or U2181 (N_2181,N_1878,N_1747);
xor U2182 (N_2182,N_1184,N_1271);
xor U2183 (N_2183,N_1410,N_1030);
nand U2184 (N_2184,N_1559,N_1800);
xnor U2185 (N_2185,N_1628,N_1318);
nor U2186 (N_2186,N_1957,N_1977);
nand U2187 (N_2187,N_1854,N_1805);
nor U2188 (N_2188,N_1055,N_1964);
and U2189 (N_2189,N_1710,N_1959);
or U2190 (N_2190,N_1140,N_1645);
xnor U2191 (N_2191,N_1361,N_1701);
nor U2192 (N_2192,N_1202,N_1984);
and U2193 (N_2193,N_1686,N_1883);
nor U2194 (N_2194,N_1200,N_1724);
xnor U2195 (N_2195,N_1901,N_1463);
or U2196 (N_2196,N_1216,N_1760);
nand U2197 (N_2197,N_1075,N_1691);
and U2198 (N_2198,N_1149,N_1052);
xnor U2199 (N_2199,N_1511,N_1887);
nor U2200 (N_2200,N_1117,N_1602);
or U2201 (N_2201,N_1839,N_1943);
and U2202 (N_2202,N_1167,N_1032);
nand U2203 (N_2203,N_1427,N_1583);
or U2204 (N_2204,N_1714,N_1061);
or U2205 (N_2205,N_1301,N_1079);
nand U2206 (N_2206,N_1147,N_1571);
or U2207 (N_2207,N_1976,N_1436);
and U2208 (N_2208,N_1394,N_1063);
or U2209 (N_2209,N_1620,N_1625);
nor U2210 (N_2210,N_1877,N_1311);
nor U2211 (N_2211,N_1251,N_1678);
nand U2212 (N_2212,N_1195,N_1924);
nor U2213 (N_2213,N_1492,N_1239);
nand U2214 (N_2214,N_1377,N_1870);
nor U2215 (N_2215,N_1152,N_1087);
and U2216 (N_2216,N_1915,N_1321);
and U2217 (N_2217,N_1324,N_1539);
nor U2218 (N_2218,N_1501,N_1508);
and U2219 (N_2219,N_1275,N_1677);
nand U2220 (N_2220,N_1801,N_1769);
nor U2221 (N_2221,N_1290,N_1507);
or U2222 (N_2222,N_1698,N_1807);
or U2223 (N_2223,N_1393,N_1875);
nor U2224 (N_2224,N_1225,N_1244);
xnor U2225 (N_2225,N_1012,N_1413);
or U2226 (N_2226,N_1082,N_1767);
nor U2227 (N_2227,N_1740,N_1858);
and U2228 (N_2228,N_1874,N_1937);
xor U2229 (N_2229,N_1738,N_1182);
or U2230 (N_2230,N_1765,N_1835);
xor U2231 (N_2231,N_1743,N_1689);
xor U2232 (N_2232,N_1160,N_1940);
nand U2233 (N_2233,N_1204,N_1623);
xor U2234 (N_2234,N_1712,N_1419);
nand U2235 (N_2235,N_1227,N_1886);
nor U2236 (N_2236,N_1542,N_1669);
xnor U2237 (N_2237,N_1619,N_1853);
or U2238 (N_2238,N_1312,N_1567);
nand U2239 (N_2239,N_1974,N_1365);
and U2240 (N_2240,N_1048,N_1389);
xnor U2241 (N_2241,N_1481,N_1841);
and U2242 (N_2242,N_1325,N_1478);
nor U2243 (N_2243,N_1836,N_1538);
nor U2244 (N_2244,N_1536,N_1777);
nor U2245 (N_2245,N_1047,N_1383);
and U2246 (N_2246,N_1073,N_1904);
or U2247 (N_2247,N_1360,N_1557);
or U2248 (N_2248,N_1823,N_1912);
nand U2249 (N_2249,N_1751,N_1493);
nor U2250 (N_2250,N_1479,N_1217);
or U2251 (N_2251,N_1041,N_1173);
nor U2252 (N_2252,N_1257,N_1057);
and U2253 (N_2253,N_1454,N_1299);
xnor U2254 (N_2254,N_1416,N_1680);
nor U2255 (N_2255,N_1961,N_1564);
nand U2256 (N_2256,N_1861,N_1863);
and U2257 (N_2257,N_1088,N_1631);
nor U2258 (N_2258,N_1778,N_1295);
nor U2259 (N_2259,N_1774,N_1750);
nor U2260 (N_2260,N_1090,N_1986);
xor U2261 (N_2261,N_1280,N_1855);
nor U2262 (N_2262,N_1722,N_1582);
or U2263 (N_2263,N_1908,N_1509);
and U2264 (N_2264,N_1343,N_1333);
nand U2265 (N_2265,N_1923,N_1363);
nand U2266 (N_2266,N_1319,N_1729);
nand U2267 (N_2267,N_1663,N_1502);
or U2268 (N_2268,N_1338,N_1476);
and U2269 (N_2269,N_1866,N_1304);
nor U2270 (N_2270,N_1814,N_1288);
and U2271 (N_2271,N_1439,N_1577);
and U2272 (N_2272,N_1451,N_1352);
or U2273 (N_2273,N_1755,N_1797);
xor U2274 (N_2274,N_1516,N_1330);
nor U2275 (N_2275,N_1696,N_1089);
xnor U2276 (N_2276,N_1871,N_1918);
and U2277 (N_2277,N_1465,N_1828);
or U2278 (N_2278,N_1856,N_1495);
or U2279 (N_2279,N_1285,N_1942);
nor U2280 (N_2280,N_1598,N_1612);
or U2281 (N_2281,N_1646,N_1737);
and U2282 (N_2282,N_1409,N_1679);
nor U2283 (N_2283,N_1424,N_1378);
nor U2284 (N_2284,N_1850,N_1113);
nor U2285 (N_2285,N_1757,N_1889);
nand U2286 (N_2286,N_1624,N_1928);
nor U2287 (N_2287,N_1817,N_1857);
and U2288 (N_2288,N_1584,N_1198);
or U2289 (N_2289,N_1715,N_1560);
nor U2290 (N_2290,N_1761,N_1756);
or U2291 (N_2291,N_1161,N_1813);
or U2292 (N_2292,N_1406,N_1846);
xnor U2293 (N_2293,N_1867,N_1530);
nor U2294 (N_2294,N_1615,N_1334);
and U2295 (N_2295,N_1411,N_1138);
and U2296 (N_2296,N_1444,N_1006);
nand U2297 (N_2297,N_1820,N_1505);
nand U2298 (N_2298,N_1380,N_1385);
xnor U2299 (N_2299,N_1914,N_1036);
xor U2300 (N_2300,N_1023,N_1263);
or U2301 (N_2301,N_1008,N_1786);
nor U2302 (N_2302,N_1323,N_1296);
nand U2303 (N_2303,N_1510,N_1293);
nor U2304 (N_2304,N_1749,N_1432);
nand U2305 (N_2305,N_1503,N_1514);
xor U2306 (N_2306,N_1392,N_1517);
or U2307 (N_2307,N_1780,N_1592);
nand U2308 (N_2308,N_1742,N_1604);
nand U2309 (N_2309,N_1816,N_1166);
xor U2310 (N_2310,N_1035,N_1744);
nor U2311 (N_2311,N_1640,N_1860);
xnor U2312 (N_2312,N_1193,N_1734);
xor U2313 (N_2313,N_1808,N_1339);
nor U2314 (N_2314,N_1151,N_1354);
or U2315 (N_2315,N_1231,N_1278);
nand U2316 (N_2316,N_1136,N_1707);
and U2317 (N_2317,N_1274,N_1622);
and U2318 (N_2318,N_1121,N_1214);
xor U2319 (N_2319,N_1556,N_1793);
or U2320 (N_2320,N_1541,N_1590);
nor U2321 (N_2321,N_1044,N_1142);
nand U2322 (N_2322,N_1906,N_1683);
xnor U2323 (N_2323,N_1025,N_1056);
and U2324 (N_2324,N_1421,N_1233);
or U2325 (N_2325,N_1137,N_1215);
xor U2326 (N_2326,N_1643,N_1357);
and U2327 (N_2327,N_1859,N_1266);
and U2328 (N_2328,N_1753,N_1328);
nor U2329 (N_2329,N_1659,N_1236);
nor U2330 (N_2330,N_1482,N_1206);
nand U2331 (N_2331,N_1327,N_1376);
or U2332 (N_2332,N_1907,N_1368);
or U2333 (N_2333,N_1076,N_1548);
nor U2334 (N_2334,N_1578,N_1477);
and U2335 (N_2335,N_1238,N_1754);
xor U2336 (N_2336,N_1979,N_1462);
nor U2337 (N_2337,N_1576,N_1666);
nand U2338 (N_2338,N_1120,N_1609);
and U2339 (N_2339,N_1995,N_1007);
nor U2340 (N_2340,N_1954,N_1390);
xor U2341 (N_2341,N_1732,N_1072);
and U2342 (N_2342,N_1768,N_1226);
nor U2343 (N_2343,N_1356,N_1110);
nor U2344 (N_2344,N_1819,N_1305);
xnor U2345 (N_2345,N_1355,N_1480);
nand U2346 (N_2346,N_1373,N_1491);
xor U2347 (N_2347,N_1806,N_1345);
xnor U2348 (N_2348,N_1403,N_1284);
nor U2349 (N_2349,N_1965,N_1457);
xnor U2350 (N_2350,N_1273,N_1074);
or U2351 (N_2351,N_1388,N_1553);
or U2352 (N_2352,N_1268,N_1430);
nand U2353 (N_2353,N_1400,N_1335);
nand U2354 (N_2354,N_1693,N_1925);
and U2355 (N_2355,N_1705,N_1381);
nand U2356 (N_2356,N_1947,N_1349);
nor U2357 (N_2357,N_1675,N_1504);
and U2358 (N_2358,N_1498,N_1983);
and U2359 (N_2359,N_1545,N_1425);
and U2360 (N_2360,N_1058,N_1116);
nor U2361 (N_2361,N_1873,N_1825);
nor U2362 (N_2362,N_1067,N_1982);
xor U2363 (N_2363,N_1287,N_1790);
nand U2364 (N_2364,N_1824,N_1651);
nand U2365 (N_2365,N_1094,N_1459);
nor U2366 (N_2366,N_1314,N_1690);
or U2367 (N_2367,N_1637,N_1010);
xor U2368 (N_2368,N_1050,N_1300);
or U2369 (N_2369,N_1639,N_1770);
nor U2370 (N_2370,N_1037,N_1528);
or U2371 (N_2371,N_1446,N_1483);
xnor U2372 (N_2372,N_1727,N_1809);
nand U2373 (N_2373,N_1246,N_1831);
or U2374 (N_2374,N_1838,N_1644);
xor U2375 (N_2375,N_1695,N_1230);
and U2376 (N_2376,N_1443,N_1374);
and U2377 (N_2377,N_1484,N_1141);
xor U2378 (N_2378,N_1083,N_1993);
nand U2379 (N_2379,N_1178,N_1020);
or U2380 (N_2380,N_1162,N_1897);
and U2381 (N_2381,N_1027,N_1610);
nor U2382 (N_2382,N_1386,N_1506);
or U2383 (N_2383,N_1524,N_1248);
or U2384 (N_2384,N_1456,N_1845);
nand U2385 (N_2385,N_1759,N_1594);
xnor U2386 (N_2386,N_1097,N_1975);
or U2387 (N_2387,N_1523,N_1156);
and U2388 (N_2388,N_1711,N_1922);
nor U2389 (N_2389,N_1634,N_1159);
xnor U2390 (N_2390,N_1652,N_1283);
or U2391 (N_2391,N_1245,N_1647);
or U2392 (N_2392,N_1662,N_1613);
and U2393 (N_2393,N_1758,N_1148);
or U2394 (N_2394,N_1862,N_1902);
nor U2395 (N_2395,N_1062,N_1779);
nor U2396 (N_2396,N_1981,N_1186);
nand U2397 (N_2397,N_1191,N_1894);
xnor U2398 (N_2398,N_1763,N_1826);
nor U2399 (N_2399,N_1992,N_1771);
or U2400 (N_2400,N_1702,N_1939);
xor U2401 (N_2401,N_1660,N_1891);
and U2402 (N_2402,N_1473,N_1851);
nand U2403 (N_2403,N_1529,N_1276);
or U2404 (N_2404,N_1210,N_1387);
and U2405 (N_2405,N_1723,N_1513);
and U2406 (N_2406,N_1474,N_1154);
or U2407 (N_2407,N_1259,N_1028);
and U2408 (N_2408,N_1091,N_1672);
nand U2409 (N_2409,N_1039,N_1337);
nor U2410 (N_2410,N_1561,N_1108);
nand U2411 (N_2411,N_1911,N_1133);
or U2412 (N_2412,N_1581,N_1967);
or U2413 (N_2413,N_1100,N_1525);
nand U2414 (N_2414,N_1626,N_1213);
xnor U2415 (N_2415,N_1921,N_1175);
nand U2416 (N_2416,N_1704,N_1998);
or U2417 (N_2417,N_1228,N_1636);
and U2418 (N_2418,N_1326,N_1589);
or U2419 (N_2419,N_1224,N_1709);
and U2420 (N_2420,N_1107,N_1629);
or U2421 (N_2421,N_1401,N_1469);
nor U2422 (N_2422,N_1150,N_1852);
nor U2423 (N_2423,N_1398,N_1320);
or U2424 (N_2424,N_1125,N_1558);
or U2425 (N_2425,N_1741,N_1811);
xor U2426 (N_2426,N_1630,N_1379);
or U2427 (N_2427,N_1029,N_1433);
or U2428 (N_2428,N_1431,N_1572);
or U2429 (N_2429,N_1784,N_1367);
nor U2430 (N_2430,N_1449,N_1059);
nand U2431 (N_2431,N_1726,N_1531);
or U2432 (N_2432,N_1250,N_1158);
nand U2433 (N_2433,N_1486,N_1329);
and U2434 (N_2434,N_1895,N_1260);
and U2435 (N_2435,N_1489,N_1331);
nand U2436 (N_2436,N_1384,N_1399);
nor U2437 (N_2437,N_1601,N_1847);
nor U2438 (N_2438,N_1188,N_1515);
nand U2439 (N_2439,N_1934,N_1575);
xor U2440 (N_2440,N_1252,N_1201);
and U2441 (N_2441,N_1593,N_1608);
nand U2442 (N_2442,N_1115,N_1879);
nand U2443 (N_2443,N_1005,N_1865);
xnor U2444 (N_2444,N_1728,N_1717);
or U2445 (N_2445,N_1165,N_1929);
or U2446 (N_2446,N_1169,N_1794);
or U2447 (N_2447,N_1235,N_1084);
or U2448 (N_2448,N_1049,N_1599);
nand U2449 (N_2449,N_1927,N_1555);
and U2450 (N_2450,N_1255,N_1358);
nand U2451 (N_2451,N_1676,N_1499);
nor U2452 (N_2452,N_1130,N_1900);
or U2453 (N_2453,N_1933,N_1408);
or U2454 (N_2454,N_1688,N_1086);
or U2455 (N_2455,N_1533,N_1591);
nand U2456 (N_2456,N_1605,N_1279);
and U2457 (N_2457,N_1080,N_1543);
nor U2458 (N_2458,N_1526,N_1415);
xnor U2459 (N_2459,N_1470,N_1950);
nand U2460 (N_2460,N_1892,N_1721);
or U2461 (N_2461,N_1322,N_1040);
nand U2462 (N_2462,N_1876,N_1455);
xnor U2463 (N_2463,N_1574,N_1112);
nand U2464 (N_2464,N_1404,N_1997);
and U2465 (N_2465,N_1002,N_1843);
nand U2466 (N_2466,N_1916,N_1344);
xor U2467 (N_2467,N_1926,N_1118);
nand U2468 (N_2468,N_1969,N_1616);
nand U2469 (N_2469,N_1682,N_1472);
xor U2470 (N_2470,N_1053,N_1256);
or U2471 (N_2471,N_1207,N_1674);
xor U2472 (N_2472,N_1512,N_1665);
nor U2473 (N_2473,N_1570,N_1648);
xor U2474 (N_2474,N_1209,N_1658);
xnor U2475 (N_2475,N_1234,N_1773);
and U2476 (N_2476,N_1359,N_1596);
and U2477 (N_2477,N_1066,N_1009);
and U2478 (N_2478,N_1970,N_1013);
xor U2479 (N_2479,N_1953,N_1932);
nand U2480 (N_2480,N_1654,N_1890);
and U2481 (N_2481,N_1971,N_1896);
nand U2482 (N_2482,N_1633,N_1042);
nand U2483 (N_2483,N_1104,N_1611);
nand U2484 (N_2484,N_1185,N_1798);
or U2485 (N_2485,N_1772,N_1661);
or U2486 (N_2486,N_1096,N_1827);
or U2487 (N_2487,N_1733,N_1655);
or U2488 (N_2488,N_1014,N_1796);
xnor U2489 (N_2489,N_1972,N_1109);
xor U2490 (N_2490,N_1544,N_1017);
and U2491 (N_2491,N_1730,N_1746);
and U2492 (N_2492,N_1348,N_1382);
nand U2493 (N_2493,N_1001,N_1497);
and U2494 (N_2494,N_1829,N_1135);
nand U2495 (N_2495,N_1372,N_1068);
and U2496 (N_2496,N_1313,N_1134);
xnor U2497 (N_2497,N_1821,N_1632);
xnor U2498 (N_2498,N_1607,N_1899);
nor U2499 (N_2499,N_1024,N_1535);
xnor U2500 (N_2500,N_1380,N_1707);
and U2501 (N_2501,N_1357,N_1958);
or U2502 (N_2502,N_1783,N_1649);
nor U2503 (N_2503,N_1804,N_1459);
nand U2504 (N_2504,N_1581,N_1567);
nand U2505 (N_2505,N_1338,N_1856);
and U2506 (N_2506,N_1617,N_1008);
or U2507 (N_2507,N_1967,N_1996);
and U2508 (N_2508,N_1138,N_1315);
xnor U2509 (N_2509,N_1231,N_1309);
nand U2510 (N_2510,N_1912,N_1522);
or U2511 (N_2511,N_1259,N_1442);
and U2512 (N_2512,N_1596,N_1654);
and U2513 (N_2513,N_1742,N_1753);
nand U2514 (N_2514,N_1503,N_1934);
or U2515 (N_2515,N_1612,N_1735);
or U2516 (N_2516,N_1999,N_1642);
nor U2517 (N_2517,N_1450,N_1709);
nand U2518 (N_2518,N_1696,N_1608);
or U2519 (N_2519,N_1248,N_1392);
nor U2520 (N_2520,N_1734,N_1148);
nand U2521 (N_2521,N_1309,N_1108);
xor U2522 (N_2522,N_1448,N_1002);
and U2523 (N_2523,N_1129,N_1967);
nor U2524 (N_2524,N_1802,N_1632);
xor U2525 (N_2525,N_1432,N_1100);
nor U2526 (N_2526,N_1953,N_1464);
and U2527 (N_2527,N_1676,N_1937);
nand U2528 (N_2528,N_1719,N_1893);
and U2529 (N_2529,N_1301,N_1613);
nor U2530 (N_2530,N_1961,N_1181);
nor U2531 (N_2531,N_1107,N_1814);
or U2532 (N_2532,N_1362,N_1736);
nand U2533 (N_2533,N_1553,N_1288);
nand U2534 (N_2534,N_1954,N_1090);
or U2535 (N_2535,N_1800,N_1147);
nand U2536 (N_2536,N_1656,N_1812);
xor U2537 (N_2537,N_1763,N_1581);
nand U2538 (N_2538,N_1947,N_1980);
and U2539 (N_2539,N_1132,N_1332);
and U2540 (N_2540,N_1511,N_1669);
nand U2541 (N_2541,N_1399,N_1120);
nor U2542 (N_2542,N_1913,N_1062);
or U2543 (N_2543,N_1256,N_1319);
nand U2544 (N_2544,N_1725,N_1006);
xor U2545 (N_2545,N_1637,N_1840);
and U2546 (N_2546,N_1900,N_1896);
xnor U2547 (N_2547,N_1103,N_1379);
xnor U2548 (N_2548,N_1983,N_1811);
nand U2549 (N_2549,N_1894,N_1337);
xor U2550 (N_2550,N_1170,N_1770);
or U2551 (N_2551,N_1134,N_1083);
or U2552 (N_2552,N_1812,N_1979);
nor U2553 (N_2553,N_1726,N_1232);
or U2554 (N_2554,N_1620,N_1092);
and U2555 (N_2555,N_1055,N_1177);
nand U2556 (N_2556,N_1851,N_1707);
or U2557 (N_2557,N_1286,N_1351);
and U2558 (N_2558,N_1111,N_1337);
or U2559 (N_2559,N_1661,N_1747);
or U2560 (N_2560,N_1052,N_1990);
xor U2561 (N_2561,N_1116,N_1573);
nand U2562 (N_2562,N_1214,N_1145);
xnor U2563 (N_2563,N_1614,N_1958);
and U2564 (N_2564,N_1872,N_1507);
nor U2565 (N_2565,N_1483,N_1992);
nand U2566 (N_2566,N_1432,N_1811);
nor U2567 (N_2567,N_1928,N_1470);
and U2568 (N_2568,N_1100,N_1910);
or U2569 (N_2569,N_1267,N_1553);
nor U2570 (N_2570,N_1024,N_1674);
xnor U2571 (N_2571,N_1557,N_1443);
nor U2572 (N_2572,N_1778,N_1191);
nor U2573 (N_2573,N_1628,N_1352);
and U2574 (N_2574,N_1806,N_1649);
or U2575 (N_2575,N_1606,N_1341);
nand U2576 (N_2576,N_1756,N_1479);
or U2577 (N_2577,N_1929,N_1046);
nor U2578 (N_2578,N_1074,N_1674);
and U2579 (N_2579,N_1468,N_1864);
and U2580 (N_2580,N_1192,N_1323);
nor U2581 (N_2581,N_1028,N_1554);
nand U2582 (N_2582,N_1824,N_1372);
nor U2583 (N_2583,N_1557,N_1300);
and U2584 (N_2584,N_1914,N_1332);
xnor U2585 (N_2585,N_1451,N_1947);
or U2586 (N_2586,N_1209,N_1835);
or U2587 (N_2587,N_1842,N_1966);
nand U2588 (N_2588,N_1564,N_1934);
xnor U2589 (N_2589,N_1379,N_1987);
nor U2590 (N_2590,N_1257,N_1143);
or U2591 (N_2591,N_1978,N_1709);
xnor U2592 (N_2592,N_1220,N_1815);
xor U2593 (N_2593,N_1605,N_1072);
xor U2594 (N_2594,N_1703,N_1079);
nor U2595 (N_2595,N_1387,N_1147);
nand U2596 (N_2596,N_1188,N_1479);
and U2597 (N_2597,N_1146,N_1421);
nor U2598 (N_2598,N_1112,N_1741);
or U2599 (N_2599,N_1866,N_1640);
and U2600 (N_2600,N_1165,N_1525);
nand U2601 (N_2601,N_1848,N_1528);
and U2602 (N_2602,N_1346,N_1445);
nand U2603 (N_2603,N_1340,N_1091);
nor U2604 (N_2604,N_1312,N_1830);
nor U2605 (N_2605,N_1649,N_1277);
nor U2606 (N_2606,N_1128,N_1248);
xnor U2607 (N_2607,N_1548,N_1516);
xnor U2608 (N_2608,N_1775,N_1563);
or U2609 (N_2609,N_1651,N_1017);
and U2610 (N_2610,N_1883,N_1320);
or U2611 (N_2611,N_1697,N_1770);
nor U2612 (N_2612,N_1154,N_1479);
nor U2613 (N_2613,N_1330,N_1752);
nand U2614 (N_2614,N_1477,N_1597);
or U2615 (N_2615,N_1652,N_1227);
xnor U2616 (N_2616,N_1794,N_1790);
xor U2617 (N_2617,N_1233,N_1718);
nand U2618 (N_2618,N_1860,N_1495);
xnor U2619 (N_2619,N_1561,N_1010);
nor U2620 (N_2620,N_1395,N_1964);
nand U2621 (N_2621,N_1138,N_1983);
xor U2622 (N_2622,N_1173,N_1597);
xnor U2623 (N_2623,N_1972,N_1852);
nor U2624 (N_2624,N_1729,N_1110);
xor U2625 (N_2625,N_1369,N_1142);
and U2626 (N_2626,N_1342,N_1396);
xor U2627 (N_2627,N_1732,N_1022);
nor U2628 (N_2628,N_1813,N_1758);
nor U2629 (N_2629,N_1132,N_1323);
and U2630 (N_2630,N_1321,N_1139);
or U2631 (N_2631,N_1812,N_1167);
or U2632 (N_2632,N_1996,N_1400);
and U2633 (N_2633,N_1329,N_1306);
nand U2634 (N_2634,N_1876,N_1309);
and U2635 (N_2635,N_1795,N_1991);
or U2636 (N_2636,N_1439,N_1398);
xnor U2637 (N_2637,N_1241,N_1412);
xor U2638 (N_2638,N_1808,N_1798);
and U2639 (N_2639,N_1809,N_1906);
xor U2640 (N_2640,N_1130,N_1021);
and U2641 (N_2641,N_1594,N_1244);
or U2642 (N_2642,N_1678,N_1900);
nor U2643 (N_2643,N_1832,N_1851);
nand U2644 (N_2644,N_1021,N_1705);
xor U2645 (N_2645,N_1564,N_1359);
or U2646 (N_2646,N_1985,N_1087);
and U2647 (N_2647,N_1589,N_1849);
or U2648 (N_2648,N_1758,N_1792);
xnor U2649 (N_2649,N_1054,N_1377);
or U2650 (N_2650,N_1959,N_1061);
xnor U2651 (N_2651,N_1568,N_1098);
and U2652 (N_2652,N_1660,N_1987);
and U2653 (N_2653,N_1266,N_1692);
and U2654 (N_2654,N_1402,N_1144);
and U2655 (N_2655,N_1540,N_1437);
nand U2656 (N_2656,N_1585,N_1595);
or U2657 (N_2657,N_1273,N_1772);
or U2658 (N_2658,N_1629,N_1008);
and U2659 (N_2659,N_1072,N_1602);
or U2660 (N_2660,N_1085,N_1857);
or U2661 (N_2661,N_1188,N_1787);
nor U2662 (N_2662,N_1710,N_1392);
nor U2663 (N_2663,N_1348,N_1540);
nor U2664 (N_2664,N_1973,N_1955);
xnor U2665 (N_2665,N_1164,N_1058);
nand U2666 (N_2666,N_1526,N_1161);
nand U2667 (N_2667,N_1119,N_1793);
xor U2668 (N_2668,N_1887,N_1241);
and U2669 (N_2669,N_1735,N_1313);
xnor U2670 (N_2670,N_1102,N_1237);
or U2671 (N_2671,N_1750,N_1099);
nor U2672 (N_2672,N_1756,N_1365);
nor U2673 (N_2673,N_1144,N_1369);
and U2674 (N_2674,N_1591,N_1574);
or U2675 (N_2675,N_1993,N_1005);
or U2676 (N_2676,N_1513,N_1375);
xor U2677 (N_2677,N_1378,N_1272);
xnor U2678 (N_2678,N_1362,N_1996);
or U2679 (N_2679,N_1514,N_1427);
and U2680 (N_2680,N_1007,N_1591);
or U2681 (N_2681,N_1894,N_1787);
or U2682 (N_2682,N_1999,N_1740);
nand U2683 (N_2683,N_1539,N_1807);
or U2684 (N_2684,N_1692,N_1501);
nor U2685 (N_2685,N_1431,N_1340);
nand U2686 (N_2686,N_1016,N_1876);
nor U2687 (N_2687,N_1587,N_1820);
nor U2688 (N_2688,N_1959,N_1747);
nor U2689 (N_2689,N_1303,N_1281);
nor U2690 (N_2690,N_1755,N_1053);
nand U2691 (N_2691,N_1504,N_1893);
nor U2692 (N_2692,N_1423,N_1823);
and U2693 (N_2693,N_1661,N_1783);
and U2694 (N_2694,N_1645,N_1969);
xor U2695 (N_2695,N_1432,N_1520);
xnor U2696 (N_2696,N_1065,N_1774);
or U2697 (N_2697,N_1707,N_1179);
nor U2698 (N_2698,N_1916,N_1037);
xor U2699 (N_2699,N_1277,N_1883);
nor U2700 (N_2700,N_1104,N_1452);
nor U2701 (N_2701,N_1377,N_1680);
and U2702 (N_2702,N_1188,N_1347);
nand U2703 (N_2703,N_1747,N_1123);
and U2704 (N_2704,N_1853,N_1640);
or U2705 (N_2705,N_1501,N_1275);
or U2706 (N_2706,N_1214,N_1031);
or U2707 (N_2707,N_1106,N_1551);
nor U2708 (N_2708,N_1748,N_1065);
nand U2709 (N_2709,N_1811,N_1231);
or U2710 (N_2710,N_1688,N_1756);
or U2711 (N_2711,N_1696,N_1163);
or U2712 (N_2712,N_1522,N_1930);
xor U2713 (N_2713,N_1401,N_1241);
nand U2714 (N_2714,N_1532,N_1208);
nor U2715 (N_2715,N_1479,N_1528);
nor U2716 (N_2716,N_1245,N_1325);
and U2717 (N_2717,N_1610,N_1402);
or U2718 (N_2718,N_1784,N_1115);
nand U2719 (N_2719,N_1242,N_1761);
xnor U2720 (N_2720,N_1318,N_1180);
or U2721 (N_2721,N_1789,N_1363);
or U2722 (N_2722,N_1085,N_1961);
nor U2723 (N_2723,N_1375,N_1623);
xnor U2724 (N_2724,N_1879,N_1747);
nand U2725 (N_2725,N_1143,N_1667);
xnor U2726 (N_2726,N_1977,N_1816);
and U2727 (N_2727,N_1689,N_1926);
and U2728 (N_2728,N_1249,N_1032);
and U2729 (N_2729,N_1813,N_1532);
nor U2730 (N_2730,N_1644,N_1045);
and U2731 (N_2731,N_1628,N_1885);
nand U2732 (N_2732,N_1701,N_1064);
or U2733 (N_2733,N_1489,N_1691);
or U2734 (N_2734,N_1805,N_1036);
nand U2735 (N_2735,N_1755,N_1061);
nor U2736 (N_2736,N_1388,N_1951);
xnor U2737 (N_2737,N_1868,N_1992);
and U2738 (N_2738,N_1684,N_1355);
nand U2739 (N_2739,N_1935,N_1671);
xnor U2740 (N_2740,N_1035,N_1737);
nand U2741 (N_2741,N_1662,N_1717);
or U2742 (N_2742,N_1560,N_1576);
xnor U2743 (N_2743,N_1717,N_1157);
xnor U2744 (N_2744,N_1444,N_1848);
and U2745 (N_2745,N_1511,N_1740);
or U2746 (N_2746,N_1651,N_1643);
nand U2747 (N_2747,N_1611,N_1994);
nor U2748 (N_2748,N_1766,N_1590);
or U2749 (N_2749,N_1003,N_1997);
or U2750 (N_2750,N_1926,N_1138);
nor U2751 (N_2751,N_1983,N_1065);
nand U2752 (N_2752,N_1474,N_1198);
nand U2753 (N_2753,N_1360,N_1294);
xnor U2754 (N_2754,N_1356,N_1807);
nand U2755 (N_2755,N_1474,N_1312);
nand U2756 (N_2756,N_1288,N_1393);
xor U2757 (N_2757,N_1278,N_1362);
xnor U2758 (N_2758,N_1378,N_1081);
and U2759 (N_2759,N_1867,N_1780);
xnor U2760 (N_2760,N_1692,N_1493);
nor U2761 (N_2761,N_1608,N_1485);
nand U2762 (N_2762,N_1148,N_1667);
or U2763 (N_2763,N_1419,N_1145);
nand U2764 (N_2764,N_1750,N_1063);
xor U2765 (N_2765,N_1544,N_1788);
and U2766 (N_2766,N_1778,N_1228);
nor U2767 (N_2767,N_1458,N_1845);
or U2768 (N_2768,N_1878,N_1400);
xor U2769 (N_2769,N_1135,N_1767);
xor U2770 (N_2770,N_1751,N_1146);
and U2771 (N_2771,N_1188,N_1897);
nor U2772 (N_2772,N_1596,N_1072);
xor U2773 (N_2773,N_1175,N_1081);
nor U2774 (N_2774,N_1235,N_1140);
nand U2775 (N_2775,N_1682,N_1791);
and U2776 (N_2776,N_1898,N_1378);
nand U2777 (N_2777,N_1894,N_1238);
nor U2778 (N_2778,N_1806,N_1563);
nor U2779 (N_2779,N_1870,N_1615);
xnor U2780 (N_2780,N_1791,N_1513);
nand U2781 (N_2781,N_1266,N_1747);
nand U2782 (N_2782,N_1452,N_1667);
xor U2783 (N_2783,N_1760,N_1712);
nor U2784 (N_2784,N_1316,N_1543);
or U2785 (N_2785,N_1210,N_1649);
and U2786 (N_2786,N_1807,N_1781);
xor U2787 (N_2787,N_1718,N_1174);
nand U2788 (N_2788,N_1741,N_1787);
or U2789 (N_2789,N_1240,N_1941);
nand U2790 (N_2790,N_1010,N_1133);
and U2791 (N_2791,N_1888,N_1774);
and U2792 (N_2792,N_1136,N_1249);
nand U2793 (N_2793,N_1103,N_1229);
xor U2794 (N_2794,N_1977,N_1085);
xnor U2795 (N_2795,N_1790,N_1892);
nand U2796 (N_2796,N_1566,N_1631);
and U2797 (N_2797,N_1766,N_1554);
nor U2798 (N_2798,N_1162,N_1489);
nand U2799 (N_2799,N_1599,N_1553);
xnor U2800 (N_2800,N_1470,N_1533);
nand U2801 (N_2801,N_1637,N_1588);
nand U2802 (N_2802,N_1951,N_1808);
nor U2803 (N_2803,N_1080,N_1590);
nor U2804 (N_2804,N_1093,N_1327);
and U2805 (N_2805,N_1217,N_1379);
nand U2806 (N_2806,N_1308,N_1965);
and U2807 (N_2807,N_1681,N_1676);
nand U2808 (N_2808,N_1672,N_1719);
nand U2809 (N_2809,N_1507,N_1258);
or U2810 (N_2810,N_1090,N_1994);
xnor U2811 (N_2811,N_1277,N_1301);
xor U2812 (N_2812,N_1312,N_1313);
xnor U2813 (N_2813,N_1758,N_1345);
and U2814 (N_2814,N_1043,N_1495);
and U2815 (N_2815,N_1549,N_1970);
or U2816 (N_2816,N_1874,N_1351);
xor U2817 (N_2817,N_1236,N_1190);
and U2818 (N_2818,N_1501,N_1605);
or U2819 (N_2819,N_1274,N_1937);
nand U2820 (N_2820,N_1930,N_1110);
or U2821 (N_2821,N_1459,N_1562);
nor U2822 (N_2822,N_1094,N_1345);
or U2823 (N_2823,N_1280,N_1528);
or U2824 (N_2824,N_1123,N_1585);
or U2825 (N_2825,N_1735,N_1821);
xor U2826 (N_2826,N_1069,N_1395);
nor U2827 (N_2827,N_1780,N_1318);
and U2828 (N_2828,N_1325,N_1313);
nor U2829 (N_2829,N_1756,N_1869);
and U2830 (N_2830,N_1265,N_1028);
and U2831 (N_2831,N_1732,N_1258);
or U2832 (N_2832,N_1867,N_1986);
nand U2833 (N_2833,N_1048,N_1127);
and U2834 (N_2834,N_1537,N_1462);
or U2835 (N_2835,N_1945,N_1478);
xnor U2836 (N_2836,N_1661,N_1118);
and U2837 (N_2837,N_1191,N_1677);
nand U2838 (N_2838,N_1400,N_1311);
nor U2839 (N_2839,N_1297,N_1831);
nand U2840 (N_2840,N_1532,N_1210);
nor U2841 (N_2841,N_1975,N_1170);
nand U2842 (N_2842,N_1286,N_1907);
nor U2843 (N_2843,N_1255,N_1326);
xor U2844 (N_2844,N_1377,N_1942);
nor U2845 (N_2845,N_1705,N_1235);
or U2846 (N_2846,N_1758,N_1186);
xnor U2847 (N_2847,N_1094,N_1075);
or U2848 (N_2848,N_1780,N_1752);
xor U2849 (N_2849,N_1111,N_1310);
and U2850 (N_2850,N_1571,N_1981);
nand U2851 (N_2851,N_1344,N_1498);
nand U2852 (N_2852,N_1056,N_1627);
xnor U2853 (N_2853,N_1917,N_1611);
xnor U2854 (N_2854,N_1333,N_1660);
nor U2855 (N_2855,N_1414,N_1860);
and U2856 (N_2856,N_1372,N_1506);
nand U2857 (N_2857,N_1403,N_1915);
nand U2858 (N_2858,N_1348,N_1313);
xor U2859 (N_2859,N_1188,N_1858);
or U2860 (N_2860,N_1987,N_1836);
xor U2861 (N_2861,N_1441,N_1267);
or U2862 (N_2862,N_1924,N_1680);
nand U2863 (N_2863,N_1310,N_1164);
xor U2864 (N_2864,N_1028,N_1677);
nor U2865 (N_2865,N_1754,N_1730);
or U2866 (N_2866,N_1288,N_1305);
xnor U2867 (N_2867,N_1607,N_1844);
and U2868 (N_2868,N_1476,N_1168);
nor U2869 (N_2869,N_1019,N_1420);
or U2870 (N_2870,N_1799,N_1900);
or U2871 (N_2871,N_1431,N_1072);
and U2872 (N_2872,N_1252,N_1168);
and U2873 (N_2873,N_1757,N_1001);
xor U2874 (N_2874,N_1257,N_1780);
and U2875 (N_2875,N_1812,N_1820);
or U2876 (N_2876,N_1476,N_1876);
nor U2877 (N_2877,N_1544,N_1376);
xor U2878 (N_2878,N_1727,N_1660);
xor U2879 (N_2879,N_1093,N_1719);
nand U2880 (N_2880,N_1685,N_1616);
and U2881 (N_2881,N_1440,N_1748);
and U2882 (N_2882,N_1151,N_1646);
and U2883 (N_2883,N_1728,N_1802);
or U2884 (N_2884,N_1789,N_1001);
xnor U2885 (N_2885,N_1415,N_1613);
and U2886 (N_2886,N_1430,N_1686);
or U2887 (N_2887,N_1405,N_1479);
xnor U2888 (N_2888,N_1748,N_1087);
nor U2889 (N_2889,N_1418,N_1004);
nand U2890 (N_2890,N_1882,N_1901);
nand U2891 (N_2891,N_1205,N_1773);
and U2892 (N_2892,N_1535,N_1814);
and U2893 (N_2893,N_1441,N_1485);
xnor U2894 (N_2894,N_1516,N_1986);
and U2895 (N_2895,N_1717,N_1533);
nand U2896 (N_2896,N_1082,N_1357);
or U2897 (N_2897,N_1627,N_1103);
nor U2898 (N_2898,N_1384,N_1491);
and U2899 (N_2899,N_1007,N_1940);
nor U2900 (N_2900,N_1259,N_1187);
or U2901 (N_2901,N_1318,N_1650);
and U2902 (N_2902,N_1401,N_1860);
nor U2903 (N_2903,N_1564,N_1887);
and U2904 (N_2904,N_1645,N_1876);
or U2905 (N_2905,N_1457,N_1730);
or U2906 (N_2906,N_1250,N_1427);
and U2907 (N_2907,N_1208,N_1567);
nand U2908 (N_2908,N_1442,N_1105);
and U2909 (N_2909,N_1123,N_1511);
or U2910 (N_2910,N_1818,N_1974);
xor U2911 (N_2911,N_1504,N_1505);
and U2912 (N_2912,N_1779,N_1399);
xor U2913 (N_2913,N_1464,N_1019);
nor U2914 (N_2914,N_1588,N_1823);
or U2915 (N_2915,N_1752,N_1814);
nor U2916 (N_2916,N_1649,N_1721);
xnor U2917 (N_2917,N_1183,N_1765);
or U2918 (N_2918,N_1769,N_1266);
and U2919 (N_2919,N_1903,N_1682);
or U2920 (N_2920,N_1212,N_1026);
and U2921 (N_2921,N_1969,N_1838);
nor U2922 (N_2922,N_1222,N_1794);
nand U2923 (N_2923,N_1559,N_1348);
xnor U2924 (N_2924,N_1446,N_1502);
and U2925 (N_2925,N_1819,N_1518);
nand U2926 (N_2926,N_1668,N_1609);
xor U2927 (N_2927,N_1525,N_1115);
or U2928 (N_2928,N_1376,N_1589);
and U2929 (N_2929,N_1483,N_1387);
or U2930 (N_2930,N_1321,N_1824);
and U2931 (N_2931,N_1399,N_1393);
nor U2932 (N_2932,N_1676,N_1066);
xnor U2933 (N_2933,N_1305,N_1586);
or U2934 (N_2934,N_1420,N_1258);
xnor U2935 (N_2935,N_1930,N_1552);
and U2936 (N_2936,N_1168,N_1147);
xor U2937 (N_2937,N_1523,N_1852);
nand U2938 (N_2938,N_1150,N_1162);
and U2939 (N_2939,N_1862,N_1955);
or U2940 (N_2940,N_1053,N_1016);
nor U2941 (N_2941,N_1393,N_1207);
and U2942 (N_2942,N_1634,N_1709);
nor U2943 (N_2943,N_1246,N_1274);
nor U2944 (N_2944,N_1637,N_1969);
and U2945 (N_2945,N_1832,N_1059);
xor U2946 (N_2946,N_1174,N_1765);
or U2947 (N_2947,N_1317,N_1861);
xor U2948 (N_2948,N_1685,N_1314);
and U2949 (N_2949,N_1055,N_1556);
or U2950 (N_2950,N_1541,N_1340);
and U2951 (N_2951,N_1561,N_1219);
nand U2952 (N_2952,N_1277,N_1491);
and U2953 (N_2953,N_1535,N_1761);
nor U2954 (N_2954,N_1997,N_1036);
xor U2955 (N_2955,N_1489,N_1501);
or U2956 (N_2956,N_1182,N_1492);
nor U2957 (N_2957,N_1173,N_1500);
xnor U2958 (N_2958,N_1882,N_1218);
xnor U2959 (N_2959,N_1843,N_1595);
xnor U2960 (N_2960,N_1945,N_1414);
nor U2961 (N_2961,N_1874,N_1268);
and U2962 (N_2962,N_1792,N_1073);
or U2963 (N_2963,N_1570,N_1411);
xnor U2964 (N_2964,N_1536,N_1500);
or U2965 (N_2965,N_1569,N_1165);
and U2966 (N_2966,N_1859,N_1286);
xnor U2967 (N_2967,N_1772,N_1096);
nand U2968 (N_2968,N_1423,N_1447);
or U2969 (N_2969,N_1118,N_1230);
nor U2970 (N_2970,N_1352,N_1350);
or U2971 (N_2971,N_1794,N_1707);
and U2972 (N_2972,N_1328,N_1205);
and U2973 (N_2973,N_1685,N_1756);
and U2974 (N_2974,N_1713,N_1499);
and U2975 (N_2975,N_1273,N_1968);
nor U2976 (N_2976,N_1679,N_1238);
or U2977 (N_2977,N_1353,N_1073);
xor U2978 (N_2978,N_1555,N_1073);
or U2979 (N_2979,N_1848,N_1389);
and U2980 (N_2980,N_1297,N_1491);
and U2981 (N_2981,N_1725,N_1012);
nand U2982 (N_2982,N_1628,N_1835);
and U2983 (N_2983,N_1823,N_1871);
and U2984 (N_2984,N_1119,N_1570);
nor U2985 (N_2985,N_1232,N_1484);
nand U2986 (N_2986,N_1810,N_1852);
xor U2987 (N_2987,N_1138,N_1230);
nor U2988 (N_2988,N_1235,N_1281);
or U2989 (N_2989,N_1115,N_1677);
nand U2990 (N_2990,N_1092,N_1666);
or U2991 (N_2991,N_1461,N_1946);
and U2992 (N_2992,N_1339,N_1366);
nor U2993 (N_2993,N_1415,N_1495);
nor U2994 (N_2994,N_1778,N_1534);
nand U2995 (N_2995,N_1598,N_1223);
and U2996 (N_2996,N_1061,N_1398);
nor U2997 (N_2997,N_1211,N_1597);
or U2998 (N_2998,N_1522,N_1125);
nor U2999 (N_2999,N_1812,N_1583);
xnor U3000 (N_3000,N_2533,N_2504);
and U3001 (N_3001,N_2791,N_2688);
or U3002 (N_3002,N_2200,N_2498);
or U3003 (N_3003,N_2662,N_2199);
nor U3004 (N_3004,N_2234,N_2870);
and U3005 (N_3005,N_2613,N_2677);
nand U3006 (N_3006,N_2718,N_2044);
nand U3007 (N_3007,N_2787,N_2620);
and U3008 (N_3008,N_2207,N_2535);
and U3009 (N_3009,N_2736,N_2125);
xor U3010 (N_3010,N_2365,N_2699);
xor U3011 (N_3011,N_2850,N_2352);
xor U3012 (N_3012,N_2858,N_2776);
and U3013 (N_3013,N_2424,N_2090);
or U3014 (N_3014,N_2060,N_2720);
nor U3015 (N_3015,N_2817,N_2384);
nor U3016 (N_3016,N_2781,N_2947);
nand U3017 (N_3017,N_2807,N_2182);
xnor U3018 (N_3018,N_2785,N_2484);
xnor U3019 (N_3019,N_2208,N_2697);
or U3020 (N_3020,N_2531,N_2844);
and U3021 (N_3021,N_2944,N_2464);
xnor U3022 (N_3022,N_2370,N_2545);
nand U3023 (N_3023,N_2655,N_2307);
and U3024 (N_3024,N_2784,N_2762);
or U3025 (N_3025,N_2281,N_2193);
nand U3026 (N_3026,N_2511,N_2777);
nand U3027 (N_3027,N_2242,N_2339);
or U3028 (N_3028,N_2948,N_2894);
or U3029 (N_3029,N_2843,N_2745);
or U3030 (N_3030,N_2441,N_2458);
nand U3031 (N_3031,N_2626,N_2457);
and U3032 (N_3032,N_2790,N_2104);
nor U3033 (N_3033,N_2961,N_2757);
nand U3034 (N_3034,N_2335,N_2711);
nand U3035 (N_3035,N_2707,N_2342);
or U3036 (N_3036,N_2916,N_2225);
nor U3037 (N_3037,N_2279,N_2656);
or U3038 (N_3038,N_2316,N_2582);
xor U3039 (N_3039,N_2192,N_2322);
and U3040 (N_3040,N_2270,N_2338);
nand U3041 (N_3041,N_2179,N_2379);
and U3042 (N_3042,N_2717,N_2703);
nor U3043 (N_3043,N_2428,N_2911);
or U3044 (N_3044,N_2884,N_2495);
and U3045 (N_3045,N_2183,N_2506);
and U3046 (N_3046,N_2128,N_2546);
xnor U3047 (N_3047,N_2489,N_2853);
nor U3048 (N_3048,N_2398,N_2111);
nand U3049 (N_3049,N_2882,N_2601);
and U3050 (N_3050,N_2002,N_2468);
or U3051 (N_3051,N_2501,N_2153);
or U3052 (N_3052,N_2009,N_2743);
and U3053 (N_3053,N_2015,N_2425);
xnor U3054 (N_3054,N_2624,N_2516);
and U3055 (N_3055,N_2888,N_2140);
and U3056 (N_3056,N_2979,N_2692);
nand U3057 (N_3057,N_2347,N_2746);
xor U3058 (N_3058,N_2170,N_2678);
and U3059 (N_3059,N_2098,N_2008);
nand U3060 (N_3060,N_2891,N_2760);
nand U3061 (N_3061,N_2303,N_2324);
nand U3062 (N_3062,N_2175,N_2215);
nor U3063 (N_3063,N_2328,N_2726);
nand U3064 (N_3064,N_2851,N_2589);
or U3065 (N_3065,N_2124,N_2114);
and U3066 (N_3066,N_2750,N_2217);
xnor U3067 (N_3067,N_2754,N_2863);
and U3068 (N_3068,N_2459,N_2701);
and U3069 (N_3069,N_2089,N_2551);
and U3070 (N_3070,N_2237,N_2910);
and U3071 (N_3071,N_2845,N_2454);
xnor U3072 (N_3072,N_2930,N_2239);
and U3073 (N_3073,N_2728,N_2210);
nand U3074 (N_3074,N_2245,N_2075);
xor U3075 (N_3075,N_2197,N_2665);
and U3076 (N_3076,N_2395,N_2928);
nand U3077 (N_3077,N_2221,N_2621);
nor U3078 (N_3078,N_2940,N_2019);
or U3079 (N_3079,N_2740,N_2190);
nand U3080 (N_3080,N_2936,N_2020);
and U3081 (N_3081,N_2082,N_2137);
nand U3082 (N_3082,N_2487,N_2660);
xor U3083 (N_3083,N_2917,N_2646);
and U3084 (N_3084,N_2393,N_2704);
nand U3085 (N_3085,N_2377,N_2938);
or U3086 (N_3086,N_2311,N_2181);
nor U3087 (N_3087,N_2046,N_2808);
nand U3088 (N_3088,N_2528,N_2856);
xor U3089 (N_3089,N_2522,N_2344);
nand U3090 (N_3090,N_2450,N_2864);
nand U3091 (N_3091,N_2722,N_2602);
or U3092 (N_3092,N_2941,N_2157);
and U3093 (N_3093,N_2134,N_2449);
and U3094 (N_3094,N_2951,N_2500);
or U3095 (N_3095,N_2686,N_2974);
and U3096 (N_3096,N_2912,N_2879);
or U3097 (N_3097,N_2466,N_2779);
nand U3098 (N_3098,N_2759,N_2399);
xnor U3099 (N_3099,N_2854,N_2364);
and U3100 (N_3100,N_2166,N_2645);
nand U3101 (N_3101,N_2542,N_2893);
xor U3102 (N_3102,N_2136,N_2422);
nand U3103 (N_3103,N_2356,N_2148);
nor U3104 (N_3104,N_2194,N_2016);
or U3105 (N_3105,N_2418,N_2191);
or U3106 (N_3106,N_2741,N_2982);
or U3107 (N_3107,N_2387,N_2249);
nand U3108 (N_3108,N_2868,N_2625);
xnor U3109 (N_3109,N_2345,N_2117);
and U3110 (N_3110,N_2878,N_2603);
nand U3111 (N_3111,N_2106,N_2548);
xnor U3112 (N_3112,N_2109,N_2608);
xor U3113 (N_3113,N_2820,N_2374);
nand U3114 (N_3114,N_2641,N_2954);
or U3115 (N_3115,N_2460,N_2556);
and U3116 (N_3116,N_2559,N_2873);
nor U3117 (N_3117,N_2381,N_2348);
or U3118 (N_3118,N_2415,N_2482);
or U3119 (N_3119,N_2828,N_2473);
or U3120 (N_3120,N_2354,N_2369);
nor U3121 (N_3121,N_2472,N_2569);
or U3122 (N_3122,N_2097,N_2923);
or U3123 (N_3123,N_2475,N_2451);
nor U3124 (N_3124,N_2276,N_2080);
or U3125 (N_3125,N_2924,N_2195);
nand U3126 (N_3126,N_2043,N_2107);
or U3127 (N_3127,N_2965,N_2386);
and U3128 (N_3128,N_2032,N_2667);
and U3129 (N_3129,N_2229,N_2251);
and U3130 (N_3130,N_2086,N_2886);
xor U3131 (N_3131,N_2039,N_2184);
nor U3132 (N_3132,N_2058,N_2513);
or U3133 (N_3133,N_2919,N_2793);
nor U3134 (N_3134,N_2629,N_2518);
and U3135 (N_3135,N_2816,N_2609);
nor U3136 (N_3136,N_2969,N_2634);
and U3137 (N_3137,N_2123,N_2768);
xor U3138 (N_3138,N_2702,N_2842);
and U3139 (N_3139,N_2801,N_2616);
or U3140 (N_3140,N_2588,N_2986);
and U3141 (N_3141,N_2054,N_2427);
and U3142 (N_3142,N_2481,N_2146);
nor U3143 (N_3143,N_2756,N_2710);
and U3144 (N_3144,N_2031,N_2292);
or U3145 (N_3145,N_2812,N_2375);
nor U3146 (N_3146,N_2942,N_2248);
and U3147 (N_3147,N_2837,N_2337);
or U3148 (N_3148,N_2929,N_2874);
or U3149 (N_3149,N_2789,N_2897);
and U3150 (N_3150,N_2599,N_2186);
or U3151 (N_3151,N_2265,N_2100);
and U3152 (N_3152,N_2168,N_2105);
nor U3153 (N_3153,N_2406,N_2231);
nand U3154 (N_3154,N_2981,N_2445);
and U3155 (N_3155,N_2714,N_2685);
or U3156 (N_3156,N_2617,N_2433);
xor U3157 (N_3157,N_2505,N_2230);
nor U3158 (N_3158,N_2669,N_2607);
or U3159 (N_3159,N_2524,N_2770);
nand U3160 (N_3160,N_2675,N_2120);
and U3161 (N_3161,N_2453,N_2680);
nor U3162 (N_3162,N_2351,N_2510);
nor U3163 (N_3163,N_2895,N_2730);
nand U3164 (N_3164,N_2663,N_2957);
or U3165 (N_3165,N_2050,N_2549);
xor U3166 (N_3166,N_2112,N_2295);
and U3167 (N_3167,N_2380,N_2313);
xnor U3168 (N_3168,N_2962,N_2698);
or U3169 (N_3169,N_2341,N_2538);
nor U3170 (N_3170,N_2640,N_2113);
xnor U3171 (N_3171,N_2417,N_2803);
or U3172 (N_3172,N_2547,N_2437);
and U3173 (N_3173,N_2595,N_2973);
and U3174 (N_3174,N_2088,N_2782);
or U3175 (N_3175,N_2918,N_2361);
or U3176 (N_3176,N_2521,N_2333);
or U3177 (N_3177,N_2411,N_2610);
nand U3178 (N_3178,N_2706,N_2169);
nor U3179 (N_3179,N_2966,N_2304);
and U3180 (N_3180,N_2805,N_2096);
or U3181 (N_3181,N_2110,N_2889);
xor U3182 (N_3182,N_2491,N_2389);
nand U3183 (N_3183,N_2036,N_2243);
and U3184 (N_3184,N_2885,N_2277);
nand U3185 (N_3185,N_2151,N_2065);
and U3186 (N_3186,N_2187,N_2848);
xnor U3187 (N_3187,N_2223,N_2026);
and U3188 (N_3188,N_2636,N_2078);
nor U3189 (N_3189,N_2494,N_2534);
or U3190 (N_3190,N_2907,N_2896);
nand U3191 (N_3191,N_2390,N_2519);
nand U3192 (N_3192,N_2975,N_2285);
and U3193 (N_3193,N_2822,N_2980);
and U3194 (N_3194,N_2672,N_2288);
and U3195 (N_3195,N_2264,N_2159);
and U3196 (N_3196,N_2984,N_2695);
and U3197 (N_3197,N_2226,N_2751);
or U3198 (N_3198,N_2727,N_2438);
or U3199 (N_3199,N_2130,N_2405);
and U3200 (N_3200,N_2371,N_2585);
and U3201 (N_3201,N_2362,N_2832);
and U3202 (N_3202,N_2849,N_2946);
and U3203 (N_3203,N_2092,N_2052);
or U3204 (N_3204,N_2250,N_2799);
nor U3205 (N_3205,N_2116,N_2034);
nor U3206 (N_3206,N_2129,N_2119);
nor U3207 (N_3207,N_2977,N_2282);
or U3208 (N_3208,N_2763,N_2527);
nor U3209 (N_3209,N_2280,N_2363);
nand U3210 (N_3210,N_2469,N_2953);
or U3211 (N_3211,N_2875,N_2788);
or U3212 (N_3212,N_2598,N_2994);
xor U3213 (N_3213,N_2829,N_2048);
xor U3214 (N_3214,N_2985,N_2715);
or U3215 (N_3215,N_2014,N_2865);
nor U3216 (N_3216,N_2053,N_2914);
nand U3217 (N_3217,N_2644,N_2566);
and U3218 (N_3218,N_2834,N_2431);
xor U3219 (N_3219,N_2859,N_2880);
nor U3220 (N_3220,N_2543,N_2594);
nand U3221 (N_3221,N_2963,N_2293);
or U3222 (N_3222,N_2876,N_2643);
nand U3223 (N_3223,N_2541,N_2811);
or U3224 (N_3224,N_2814,N_2045);
nor U3225 (N_3225,N_2298,N_2263);
or U3226 (N_3226,N_2758,N_2087);
and U3227 (N_3227,N_2121,N_2557);
xor U3228 (N_3228,N_2841,N_2318);
xor U3229 (N_3229,N_2135,N_2448);
nor U3230 (N_3230,N_2971,N_2723);
nand U3231 (N_3231,N_2302,N_2887);
and U3232 (N_3232,N_2290,N_2622);
xnor U3233 (N_3233,N_2143,N_2471);
and U3234 (N_3234,N_2964,N_2666);
nand U3235 (N_3235,N_2041,N_2206);
xor U3236 (N_3236,N_2978,N_2131);
or U3237 (N_3237,N_2299,N_2198);
xor U3238 (N_3238,N_2103,N_2508);
and U3239 (N_3239,N_2765,N_2490);
nor U3240 (N_3240,N_2262,N_2689);
or U3241 (N_3241,N_2650,N_2514);
and U3242 (N_3242,N_2806,N_2319);
xnor U3243 (N_3243,N_2553,N_2839);
or U3244 (N_3244,N_2001,N_2496);
nand U3245 (N_3245,N_2783,N_2988);
or U3246 (N_3246,N_2796,N_2838);
nand U3247 (N_3247,N_2890,N_2881);
or U3248 (N_3248,N_2353,N_2639);
nand U3249 (N_3249,N_2385,N_2647);
xnor U3250 (N_3250,N_2430,N_2523);
nand U3251 (N_3251,N_2410,N_2631);
or U3252 (N_3252,N_2778,N_2580);
xor U3253 (N_3253,N_2483,N_2612);
and U3254 (N_3254,N_2819,N_2004);
xnor U3255 (N_3255,N_2188,N_2567);
xnor U3256 (N_3256,N_2220,N_2359);
nand U3257 (N_3257,N_2479,N_2266);
nand U3258 (N_3258,N_2637,N_2224);
nor U3259 (N_3259,N_2679,N_2797);
and U3260 (N_3260,N_2826,N_2115);
or U3261 (N_3261,N_2142,N_2145);
nor U3262 (N_3262,N_2259,N_2877);
nand U3263 (N_3263,N_2925,N_2550);
or U3264 (N_3264,N_2139,N_2712);
xor U3265 (N_3265,N_2657,N_2872);
nor U3266 (N_3266,N_2767,N_2561);
and U3267 (N_3267,N_2150,N_2544);
nor U3268 (N_3268,N_2898,N_2840);
or U3269 (N_3269,N_2989,N_2520);
and U3270 (N_3270,N_2126,N_2492);
xor U3271 (N_3271,N_2772,N_2164);
nand U3272 (N_3272,N_2042,N_2604);
nand U3273 (N_3273,N_2138,N_2416);
and U3274 (N_3274,N_2211,N_2570);
nand U3275 (N_3275,N_2586,N_2252);
and U3276 (N_3276,N_2771,N_2012);
xor U3277 (N_3277,N_2540,N_2809);
nand U3278 (N_3278,N_2798,N_2273);
nor U3279 (N_3279,N_2382,N_2857);
xnor U3280 (N_3280,N_2499,N_2670);
nand U3281 (N_3281,N_2400,N_2795);
or U3282 (N_3282,N_2794,N_2530);
nor U3283 (N_3283,N_2572,N_2584);
xor U3284 (N_3284,N_2301,N_2325);
and U3285 (N_3285,N_2003,N_2600);
or U3286 (N_3286,N_2436,N_2284);
and U3287 (N_3287,N_2420,N_2247);
nor U3288 (N_3288,N_2018,N_2581);
xor U3289 (N_3289,N_2291,N_2755);
or U3290 (N_3290,N_2824,N_2493);
and U3291 (N_3291,N_2439,N_2007);
or U3292 (N_3292,N_2388,N_2274);
nand U3293 (N_3293,N_2228,N_2900);
and U3294 (N_3294,N_2470,N_2509);
and U3295 (N_3295,N_2651,N_2959);
nor U3296 (N_3296,N_2654,N_2958);
nand U3297 (N_3297,N_2397,N_2476);
xor U3298 (N_3298,N_2764,N_2869);
and U3299 (N_3299,N_2346,N_2413);
xor U3300 (N_3300,N_2235,N_2827);
nor U3301 (N_3301,N_2158,N_2774);
and U3302 (N_3302,N_2611,N_2972);
nand U3303 (N_3303,N_2721,N_2414);
or U3304 (N_3304,N_2005,N_2246);
xnor U3305 (N_3305,N_2664,N_2577);
or U3306 (N_3306,N_2683,N_2308);
nand U3307 (N_3307,N_2724,N_2057);
xor U3308 (N_3308,N_2079,N_2592);
nand U3309 (N_3309,N_2267,N_2578);
nor U3310 (N_3310,N_2681,N_2905);
or U3311 (N_3311,N_2310,N_2635);
or U3312 (N_3312,N_2283,N_2573);
nand U3313 (N_3313,N_2214,N_2071);
nor U3314 (N_3314,N_2605,N_2349);
nand U3315 (N_3315,N_2006,N_2571);
and U3316 (N_3316,N_2227,N_2434);
nor U3317 (N_3317,N_2147,N_2687);
xor U3318 (N_3318,N_2378,N_2172);
and U3319 (N_3319,N_2769,N_2674);
or U3320 (N_3320,N_2825,N_2871);
xor U3321 (N_3321,N_2892,N_2899);
and U3322 (N_3322,N_2073,N_2321);
nor U3323 (N_3323,N_2070,N_2013);
xor U3324 (N_3324,N_2628,N_2336);
and U3325 (N_3325,N_2102,N_2465);
and U3326 (N_3326,N_2932,N_2537);
nor U3327 (N_3327,N_2272,N_2461);
or U3328 (N_3328,N_2419,N_2462);
nor U3329 (N_3329,N_2709,N_2440);
or U3330 (N_3330,N_2922,N_2945);
and U3331 (N_3331,N_2861,N_2144);
or U3332 (N_3332,N_2030,N_2554);
or U3333 (N_3333,N_2976,N_2761);
nand U3334 (N_3334,N_2821,N_2312);
xnor U3335 (N_3335,N_2485,N_2529);
xor U3336 (N_3336,N_2368,N_2309);
nor U3337 (N_3337,N_2040,N_2253);
xor U3338 (N_3338,N_2023,N_2627);
nand U3339 (N_3339,N_2810,N_2038);
nor U3340 (N_3340,N_2452,N_2331);
nand U3341 (N_3341,N_2056,N_2512);
or U3342 (N_3342,N_2326,N_2401);
and U3343 (N_3343,N_2132,N_2160);
or U3344 (N_3344,N_2261,N_2503);
nand U3345 (N_3345,N_2708,N_2334);
xor U3346 (N_3346,N_2463,N_2067);
or U3347 (N_3347,N_2022,N_2196);
or U3348 (N_3348,N_2737,N_2992);
nand U3349 (N_3349,N_2939,N_2920);
xnor U3350 (N_3350,N_2081,N_2507);
nor U3351 (N_3351,N_2101,N_2412);
nand U3352 (N_3352,N_2268,N_2069);
nand U3353 (N_3353,N_2367,N_2987);
or U3354 (N_3354,N_2011,N_2024);
nor U3355 (N_3355,N_2659,N_2202);
nand U3356 (N_3356,N_2804,N_2502);
and U3357 (N_3357,N_2576,N_2456);
nand U3358 (N_3358,N_2565,N_2536);
or U3359 (N_3359,N_2350,N_2652);
xor U3360 (N_3360,N_2355,N_2590);
nand U3361 (N_3361,N_2661,N_2835);
or U3362 (N_3362,N_2360,N_2269);
xor U3363 (N_3363,N_2133,N_2515);
nor U3364 (N_3364,N_2673,N_2775);
xor U3365 (N_3365,N_2244,N_2236);
or U3366 (N_3366,N_2676,N_2357);
and U3367 (N_3367,N_2391,N_2731);
nor U3368 (N_3368,N_2085,N_2099);
xnor U3369 (N_3369,N_2062,N_2167);
nand U3370 (N_3370,N_2327,N_2421);
xnor U3371 (N_3371,N_2860,N_2447);
and U3372 (N_3372,N_2862,N_2408);
xnor U3373 (N_3373,N_2035,N_2474);
nand U3374 (N_3374,N_2562,N_2021);
and U3375 (N_3375,N_2122,N_2830);
xnor U3376 (N_3376,N_2693,N_2432);
or U3377 (N_3377,N_2480,N_2563);
nor U3378 (N_3378,N_2028,N_2943);
nand U3379 (N_3379,N_2077,N_2162);
nand U3380 (N_3380,N_2323,N_2780);
or U3381 (N_3381,N_2921,N_2615);
and U3382 (N_3382,N_2995,N_2671);
nor U3383 (N_3383,N_2802,N_2061);
nor U3384 (N_3384,N_2638,N_2189);
nor U3385 (N_3385,N_2329,N_2185);
or U3386 (N_3386,N_2950,N_2847);
xor U3387 (N_3387,N_2068,N_2084);
nand U3388 (N_3388,N_2642,N_2998);
nor U3389 (N_3389,N_2340,N_2619);
nor U3390 (N_3390,N_2725,N_2317);
xor U3391 (N_3391,N_2552,N_2937);
nor U3392 (N_3392,N_2933,N_2118);
and U3393 (N_3393,N_2154,N_2000);
nor U3394 (N_3394,N_2256,N_2343);
xnor U3395 (N_3395,N_2064,N_2171);
nor U3396 (N_3396,N_2684,N_2591);
or U3397 (N_3397,N_2213,N_2402);
nor U3398 (N_3398,N_2033,N_2752);
xnor U3399 (N_3399,N_2955,N_2867);
xor U3400 (N_3400,N_2564,N_2127);
xnor U3401 (N_3401,N_2314,N_2967);
nand U3402 (N_3402,N_2606,N_2883);
xnor U3403 (N_3403,N_2255,N_2108);
nand U3404 (N_3404,N_2063,N_2271);
xnor U3405 (N_3405,N_2903,N_2792);
xnor U3406 (N_3406,N_2539,N_2532);
xnor U3407 (N_3407,N_2156,N_2165);
nor U3408 (N_3408,N_2748,N_2583);
and U3409 (N_3409,N_2394,N_2999);
nor U3410 (N_3410,N_2525,N_2155);
nand U3411 (N_3411,N_2330,N_2823);
and U3412 (N_3412,N_2178,N_2558);
xnor U3413 (N_3413,N_2435,N_2332);
nand U3414 (N_3414,N_2855,N_2747);
nand U3415 (N_3415,N_2051,N_2729);
or U3416 (N_3416,N_2913,N_2993);
nand U3417 (N_3417,N_2927,N_2204);
nor U3418 (N_3418,N_2209,N_2218);
nand U3419 (N_3419,N_2222,N_2467);
nand U3420 (N_3420,N_2478,N_2488);
nor U3421 (N_3421,N_2593,N_2296);
nand U3422 (N_3422,N_2091,N_2297);
and U3423 (N_3423,N_2444,N_2396);
or U3424 (N_3424,N_2025,N_2815);
nor U3425 (N_3425,N_2066,N_2149);
or U3426 (N_3426,N_2596,N_2749);
nand U3427 (N_3427,N_2205,N_2059);
nor U3428 (N_3428,N_2152,N_2904);
and U3429 (N_3429,N_2161,N_2426);
or U3430 (N_3430,N_2176,N_2700);
nand U3431 (N_3431,N_2094,N_2734);
xnor U3432 (N_3432,N_2083,N_2833);
nor U3433 (N_3433,N_2668,N_2970);
nand U3434 (N_3434,N_2423,N_2648);
xor U3435 (N_3435,N_2901,N_2409);
and U3436 (N_3436,N_2597,N_2201);
nor U3437 (N_3437,N_2983,N_2173);
nor U3438 (N_3438,N_2935,N_2934);
and U3439 (N_3439,N_2739,N_2497);
and U3440 (N_3440,N_2649,N_2831);
and U3441 (N_3441,N_2254,N_2278);
nor U3442 (N_3442,N_2902,N_2180);
xnor U3443 (N_3443,N_2238,N_2836);
nand U3444 (N_3444,N_2455,N_2076);
and U3445 (N_3445,N_2047,N_2163);
nand U3446 (N_3446,N_2568,N_2753);
nor U3447 (N_3447,N_2072,N_2909);
xnor U3448 (N_3448,N_2653,N_2141);
nand U3449 (N_3449,N_2372,N_2719);
nor U3450 (N_3450,N_2575,N_2358);
or U3451 (N_3451,N_2813,N_2996);
nor U3452 (N_3452,N_2174,N_2404);
and U3453 (N_3453,N_2579,N_2691);
and U3454 (N_3454,N_2010,N_2713);
nor U3455 (N_3455,N_2733,N_2287);
and U3456 (N_3456,N_2260,N_2305);
nand U3457 (N_3457,N_2429,N_2614);
nor U3458 (N_3458,N_2786,N_2027);
nor U3459 (N_3459,N_2956,N_2017);
nand U3460 (N_3460,N_2232,N_2818);
nor U3461 (N_3461,N_2526,N_2219);
xor U3462 (N_3462,N_2732,N_2952);
xnor U3463 (N_3463,N_2300,N_2392);
and U3464 (N_3464,N_2906,N_2968);
and U3465 (N_3465,N_2443,N_2555);
and U3466 (N_3466,N_2306,N_2630);
and U3467 (N_3467,N_2240,N_2633);
nor U3468 (N_3468,N_2658,N_2212);
nand U3469 (N_3469,N_2037,N_2990);
nor U3470 (N_3470,N_2407,N_2632);
xor U3471 (N_3471,N_2682,N_2477);
nand U3472 (N_3472,N_2320,N_2258);
nor U3473 (N_3473,N_2093,N_2742);
nor U3474 (N_3474,N_2800,N_2366);
nor U3475 (N_3475,N_2690,N_2315);
nor U3476 (N_3476,N_2623,N_2373);
nand U3477 (N_3477,N_2997,N_2049);
xor U3478 (N_3478,N_2766,N_2074);
nand U3479 (N_3479,N_2289,N_2383);
xnor U3480 (N_3480,N_2442,N_2286);
and U3481 (N_3481,N_2203,N_2587);
and U3482 (N_3482,N_2517,N_2029);
xor U3483 (N_3483,N_2931,N_2055);
nor U3484 (N_3484,N_2095,N_2846);
or U3485 (N_3485,N_2960,N_2908);
or U3486 (N_3486,N_2560,N_2744);
xor U3487 (N_3487,N_2738,N_2446);
or U3488 (N_3488,N_2216,N_2852);
and U3489 (N_3489,N_2403,N_2949);
nand U3490 (N_3490,N_2705,N_2177);
nor U3491 (N_3491,N_2486,N_2257);
xnor U3492 (N_3492,N_2716,N_2696);
xnor U3493 (N_3493,N_2866,N_2694);
xnor U3494 (N_3494,N_2735,N_2241);
nand U3495 (N_3495,N_2294,N_2618);
nand U3496 (N_3496,N_2233,N_2926);
xnor U3497 (N_3497,N_2376,N_2574);
nand U3498 (N_3498,N_2915,N_2773);
xnor U3499 (N_3499,N_2275,N_2991);
and U3500 (N_3500,N_2096,N_2040);
nand U3501 (N_3501,N_2052,N_2837);
and U3502 (N_3502,N_2137,N_2418);
and U3503 (N_3503,N_2225,N_2172);
xnor U3504 (N_3504,N_2671,N_2907);
nand U3505 (N_3505,N_2806,N_2527);
and U3506 (N_3506,N_2052,N_2276);
or U3507 (N_3507,N_2778,N_2002);
nor U3508 (N_3508,N_2667,N_2609);
nand U3509 (N_3509,N_2099,N_2540);
nor U3510 (N_3510,N_2216,N_2589);
nor U3511 (N_3511,N_2711,N_2776);
nor U3512 (N_3512,N_2258,N_2483);
nand U3513 (N_3513,N_2124,N_2033);
nor U3514 (N_3514,N_2498,N_2614);
and U3515 (N_3515,N_2944,N_2175);
nor U3516 (N_3516,N_2004,N_2273);
nor U3517 (N_3517,N_2184,N_2356);
and U3518 (N_3518,N_2523,N_2718);
xnor U3519 (N_3519,N_2011,N_2428);
or U3520 (N_3520,N_2621,N_2703);
nor U3521 (N_3521,N_2515,N_2006);
or U3522 (N_3522,N_2165,N_2544);
or U3523 (N_3523,N_2716,N_2326);
nand U3524 (N_3524,N_2395,N_2768);
nand U3525 (N_3525,N_2436,N_2344);
and U3526 (N_3526,N_2450,N_2303);
nor U3527 (N_3527,N_2220,N_2540);
or U3528 (N_3528,N_2047,N_2475);
and U3529 (N_3529,N_2277,N_2025);
nor U3530 (N_3530,N_2512,N_2878);
xor U3531 (N_3531,N_2830,N_2136);
and U3532 (N_3532,N_2019,N_2632);
nand U3533 (N_3533,N_2096,N_2767);
and U3534 (N_3534,N_2369,N_2899);
nand U3535 (N_3535,N_2716,N_2386);
xor U3536 (N_3536,N_2324,N_2709);
xnor U3537 (N_3537,N_2115,N_2818);
or U3538 (N_3538,N_2428,N_2553);
and U3539 (N_3539,N_2509,N_2214);
nand U3540 (N_3540,N_2009,N_2379);
nor U3541 (N_3541,N_2110,N_2094);
and U3542 (N_3542,N_2280,N_2966);
xnor U3543 (N_3543,N_2146,N_2316);
or U3544 (N_3544,N_2496,N_2565);
nor U3545 (N_3545,N_2783,N_2293);
or U3546 (N_3546,N_2308,N_2222);
xnor U3547 (N_3547,N_2793,N_2337);
xor U3548 (N_3548,N_2326,N_2832);
or U3549 (N_3549,N_2701,N_2942);
or U3550 (N_3550,N_2190,N_2973);
xor U3551 (N_3551,N_2555,N_2428);
nand U3552 (N_3552,N_2010,N_2403);
xor U3553 (N_3553,N_2019,N_2602);
nor U3554 (N_3554,N_2244,N_2560);
or U3555 (N_3555,N_2162,N_2825);
or U3556 (N_3556,N_2068,N_2445);
and U3557 (N_3557,N_2316,N_2029);
xor U3558 (N_3558,N_2986,N_2197);
or U3559 (N_3559,N_2782,N_2349);
and U3560 (N_3560,N_2273,N_2477);
nor U3561 (N_3561,N_2966,N_2814);
or U3562 (N_3562,N_2588,N_2609);
xor U3563 (N_3563,N_2904,N_2287);
xnor U3564 (N_3564,N_2297,N_2095);
nor U3565 (N_3565,N_2621,N_2930);
or U3566 (N_3566,N_2561,N_2514);
xor U3567 (N_3567,N_2375,N_2432);
and U3568 (N_3568,N_2280,N_2741);
nor U3569 (N_3569,N_2340,N_2538);
xor U3570 (N_3570,N_2735,N_2599);
or U3571 (N_3571,N_2771,N_2209);
or U3572 (N_3572,N_2286,N_2699);
nor U3573 (N_3573,N_2115,N_2902);
nand U3574 (N_3574,N_2441,N_2249);
nor U3575 (N_3575,N_2622,N_2153);
nand U3576 (N_3576,N_2940,N_2817);
nor U3577 (N_3577,N_2203,N_2223);
nand U3578 (N_3578,N_2413,N_2586);
and U3579 (N_3579,N_2652,N_2461);
and U3580 (N_3580,N_2248,N_2614);
xor U3581 (N_3581,N_2108,N_2410);
nor U3582 (N_3582,N_2089,N_2066);
nor U3583 (N_3583,N_2318,N_2257);
nand U3584 (N_3584,N_2155,N_2146);
nor U3585 (N_3585,N_2025,N_2634);
or U3586 (N_3586,N_2606,N_2748);
nor U3587 (N_3587,N_2596,N_2387);
nor U3588 (N_3588,N_2330,N_2179);
and U3589 (N_3589,N_2256,N_2082);
nand U3590 (N_3590,N_2559,N_2909);
xnor U3591 (N_3591,N_2007,N_2374);
nand U3592 (N_3592,N_2075,N_2330);
xor U3593 (N_3593,N_2905,N_2029);
nand U3594 (N_3594,N_2165,N_2224);
nor U3595 (N_3595,N_2945,N_2784);
or U3596 (N_3596,N_2363,N_2986);
nand U3597 (N_3597,N_2204,N_2809);
and U3598 (N_3598,N_2006,N_2071);
nand U3599 (N_3599,N_2318,N_2190);
xor U3600 (N_3600,N_2099,N_2621);
nor U3601 (N_3601,N_2751,N_2352);
and U3602 (N_3602,N_2055,N_2957);
nor U3603 (N_3603,N_2367,N_2402);
nor U3604 (N_3604,N_2685,N_2256);
nor U3605 (N_3605,N_2618,N_2092);
nor U3606 (N_3606,N_2204,N_2984);
nor U3607 (N_3607,N_2823,N_2636);
nor U3608 (N_3608,N_2768,N_2834);
xor U3609 (N_3609,N_2163,N_2442);
nor U3610 (N_3610,N_2194,N_2979);
nand U3611 (N_3611,N_2050,N_2513);
nor U3612 (N_3612,N_2738,N_2788);
and U3613 (N_3613,N_2948,N_2213);
nand U3614 (N_3614,N_2934,N_2764);
and U3615 (N_3615,N_2315,N_2671);
nand U3616 (N_3616,N_2614,N_2062);
and U3617 (N_3617,N_2985,N_2718);
nand U3618 (N_3618,N_2302,N_2954);
nand U3619 (N_3619,N_2733,N_2704);
or U3620 (N_3620,N_2995,N_2834);
xnor U3621 (N_3621,N_2044,N_2986);
or U3622 (N_3622,N_2683,N_2285);
xnor U3623 (N_3623,N_2661,N_2626);
nor U3624 (N_3624,N_2720,N_2722);
nor U3625 (N_3625,N_2901,N_2721);
and U3626 (N_3626,N_2494,N_2523);
and U3627 (N_3627,N_2221,N_2790);
xnor U3628 (N_3628,N_2075,N_2015);
nand U3629 (N_3629,N_2688,N_2984);
and U3630 (N_3630,N_2411,N_2509);
and U3631 (N_3631,N_2493,N_2719);
nand U3632 (N_3632,N_2632,N_2264);
nand U3633 (N_3633,N_2702,N_2774);
and U3634 (N_3634,N_2842,N_2426);
and U3635 (N_3635,N_2858,N_2987);
nor U3636 (N_3636,N_2447,N_2492);
nor U3637 (N_3637,N_2599,N_2323);
and U3638 (N_3638,N_2237,N_2166);
nand U3639 (N_3639,N_2586,N_2636);
nand U3640 (N_3640,N_2233,N_2741);
and U3641 (N_3641,N_2453,N_2194);
and U3642 (N_3642,N_2923,N_2628);
nor U3643 (N_3643,N_2703,N_2953);
xnor U3644 (N_3644,N_2203,N_2093);
and U3645 (N_3645,N_2554,N_2770);
xor U3646 (N_3646,N_2072,N_2493);
and U3647 (N_3647,N_2577,N_2331);
xor U3648 (N_3648,N_2710,N_2350);
xnor U3649 (N_3649,N_2903,N_2390);
nand U3650 (N_3650,N_2859,N_2659);
or U3651 (N_3651,N_2647,N_2048);
nand U3652 (N_3652,N_2413,N_2153);
or U3653 (N_3653,N_2194,N_2917);
xor U3654 (N_3654,N_2272,N_2528);
nor U3655 (N_3655,N_2936,N_2072);
nor U3656 (N_3656,N_2555,N_2664);
nor U3657 (N_3657,N_2071,N_2249);
nand U3658 (N_3658,N_2857,N_2946);
nor U3659 (N_3659,N_2194,N_2334);
nand U3660 (N_3660,N_2317,N_2458);
or U3661 (N_3661,N_2195,N_2531);
nand U3662 (N_3662,N_2055,N_2282);
and U3663 (N_3663,N_2551,N_2101);
nand U3664 (N_3664,N_2996,N_2478);
and U3665 (N_3665,N_2326,N_2871);
nand U3666 (N_3666,N_2720,N_2577);
nor U3667 (N_3667,N_2926,N_2608);
or U3668 (N_3668,N_2534,N_2587);
xnor U3669 (N_3669,N_2761,N_2929);
nand U3670 (N_3670,N_2873,N_2980);
or U3671 (N_3671,N_2365,N_2240);
or U3672 (N_3672,N_2173,N_2662);
and U3673 (N_3673,N_2131,N_2363);
xor U3674 (N_3674,N_2591,N_2235);
xor U3675 (N_3675,N_2192,N_2371);
xnor U3676 (N_3676,N_2029,N_2200);
nand U3677 (N_3677,N_2855,N_2981);
nor U3678 (N_3678,N_2839,N_2968);
nor U3679 (N_3679,N_2674,N_2307);
nor U3680 (N_3680,N_2772,N_2480);
and U3681 (N_3681,N_2288,N_2823);
or U3682 (N_3682,N_2412,N_2402);
nor U3683 (N_3683,N_2424,N_2236);
nor U3684 (N_3684,N_2608,N_2687);
xor U3685 (N_3685,N_2998,N_2013);
and U3686 (N_3686,N_2797,N_2042);
nor U3687 (N_3687,N_2891,N_2081);
nand U3688 (N_3688,N_2342,N_2131);
nor U3689 (N_3689,N_2400,N_2670);
nor U3690 (N_3690,N_2790,N_2608);
and U3691 (N_3691,N_2042,N_2972);
nor U3692 (N_3692,N_2291,N_2585);
or U3693 (N_3693,N_2585,N_2961);
and U3694 (N_3694,N_2922,N_2202);
and U3695 (N_3695,N_2580,N_2840);
xor U3696 (N_3696,N_2873,N_2892);
or U3697 (N_3697,N_2452,N_2146);
nor U3698 (N_3698,N_2536,N_2430);
or U3699 (N_3699,N_2460,N_2665);
and U3700 (N_3700,N_2053,N_2309);
and U3701 (N_3701,N_2422,N_2896);
nor U3702 (N_3702,N_2416,N_2534);
and U3703 (N_3703,N_2586,N_2752);
nand U3704 (N_3704,N_2081,N_2268);
nand U3705 (N_3705,N_2966,N_2294);
nand U3706 (N_3706,N_2344,N_2554);
or U3707 (N_3707,N_2011,N_2140);
and U3708 (N_3708,N_2932,N_2023);
nor U3709 (N_3709,N_2870,N_2989);
xnor U3710 (N_3710,N_2281,N_2936);
xor U3711 (N_3711,N_2252,N_2359);
nand U3712 (N_3712,N_2764,N_2942);
nor U3713 (N_3713,N_2562,N_2300);
xor U3714 (N_3714,N_2132,N_2153);
xor U3715 (N_3715,N_2746,N_2011);
or U3716 (N_3716,N_2410,N_2346);
xnor U3717 (N_3717,N_2033,N_2586);
or U3718 (N_3718,N_2997,N_2300);
xor U3719 (N_3719,N_2357,N_2293);
or U3720 (N_3720,N_2024,N_2545);
nand U3721 (N_3721,N_2784,N_2017);
xnor U3722 (N_3722,N_2519,N_2938);
xor U3723 (N_3723,N_2481,N_2856);
nand U3724 (N_3724,N_2374,N_2030);
and U3725 (N_3725,N_2862,N_2205);
nor U3726 (N_3726,N_2809,N_2045);
xor U3727 (N_3727,N_2236,N_2262);
or U3728 (N_3728,N_2990,N_2548);
nor U3729 (N_3729,N_2352,N_2542);
nand U3730 (N_3730,N_2892,N_2208);
and U3731 (N_3731,N_2076,N_2837);
nand U3732 (N_3732,N_2840,N_2869);
or U3733 (N_3733,N_2026,N_2845);
nor U3734 (N_3734,N_2932,N_2639);
nand U3735 (N_3735,N_2647,N_2118);
nor U3736 (N_3736,N_2337,N_2366);
or U3737 (N_3737,N_2665,N_2036);
or U3738 (N_3738,N_2846,N_2723);
nor U3739 (N_3739,N_2725,N_2228);
and U3740 (N_3740,N_2053,N_2285);
nand U3741 (N_3741,N_2036,N_2125);
and U3742 (N_3742,N_2508,N_2811);
or U3743 (N_3743,N_2272,N_2642);
nor U3744 (N_3744,N_2501,N_2630);
or U3745 (N_3745,N_2616,N_2296);
nand U3746 (N_3746,N_2755,N_2440);
nor U3747 (N_3747,N_2721,N_2434);
nor U3748 (N_3748,N_2063,N_2225);
or U3749 (N_3749,N_2267,N_2751);
xor U3750 (N_3750,N_2565,N_2903);
or U3751 (N_3751,N_2258,N_2260);
nand U3752 (N_3752,N_2198,N_2922);
or U3753 (N_3753,N_2628,N_2294);
or U3754 (N_3754,N_2421,N_2958);
nand U3755 (N_3755,N_2678,N_2406);
or U3756 (N_3756,N_2305,N_2759);
nor U3757 (N_3757,N_2430,N_2626);
xnor U3758 (N_3758,N_2441,N_2690);
nand U3759 (N_3759,N_2623,N_2528);
or U3760 (N_3760,N_2187,N_2127);
nand U3761 (N_3761,N_2472,N_2844);
or U3762 (N_3762,N_2485,N_2899);
nand U3763 (N_3763,N_2702,N_2657);
and U3764 (N_3764,N_2014,N_2238);
or U3765 (N_3765,N_2967,N_2960);
nand U3766 (N_3766,N_2859,N_2924);
nor U3767 (N_3767,N_2957,N_2867);
and U3768 (N_3768,N_2819,N_2278);
and U3769 (N_3769,N_2016,N_2057);
nand U3770 (N_3770,N_2643,N_2989);
and U3771 (N_3771,N_2096,N_2651);
xor U3772 (N_3772,N_2596,N_2914);
or U3773 (N_3773,N_2922,N_2676);
nand U3774 (N_3774,N_2971,N_2677);
or U3775 (N_3775,N_2630,N_2312);
nand U3776 (N_3776,N_2313,N_2977);
and U3777 (N_3777,N_2006,N_2772);
and U3778 (N_3778,N_2664,N_2814);
nor U3779 (N_3779,N_2524,N_2880);
or U3780 (N_3780,N_2806,N_2875);
and U3781 (N_3781,N_2788,N_2661);
xor U3782 (N_3782,N_2605,N_2618);
xnor U3783 (N_3783,N_2157,N_2643);
xor U3784 (N_3784,N_2349,N_2206);
or U3785 (N_3785,N_2429,N_2688);
nand U3786 (N_3786,N_2564,N_2341);
or U3787 (N_3787,N_2941,N_2546);
xor U3788 (N_3788,N_2504,N_2195);
and U3789 (N_3789,N_2461,N_2951);
nand U3790 (N_3790,N_2057,N_2346);
nand U3791 (N_3791,N_2752,N_2198);
or U3792 (N_3792,N_2282,N_2371);
or U3793 (N_3793,N_2474,N_2918);
nand U3794 (N_3794,N_2549,N_2852);
or U3795 (N_3795,N_2645,N_2715);
nor U3796 (N_3796,N_2140,N_2724);
or U3797 (N_3797,N_2731,N_2928);
or U3798 (N_3798,N_2671,N_2665);
nor U3799 (N_3799,N_2011,N_2057);
and U3800 (N_3800,N_2262,N_2846);
or U3801 (N_3801,N_2686,N_2039);
and U3802 (N_3802,N_2324,N_2169);
xnor U3803 (N_3803,N_2846,N_2297);
or U3804 (N_3804,N_2486,N_2954);
and U3805 (N_3805,N_2286,N_2353);
or U3806 (N_3806,N_2704,N_2996);
nor U3807 (N_3807,N_2097,N_2306);
or U3808 (N_3808,N_2778,N_2248);
xnor U3809 (N_3809,N_2474,N_2466);
and U3810 (N_3810,N_2074,N_2711);
xnor U3811 (N_3811,N_2397,N_2693);
nor U3812 (N_3812,N_2085,N_2732);
nand U3813 (N_3813,N_2983,N_2741);
or U3814 (N_3814,N_2907,N_2824);
or U3815 (N_3815,N_2756,N_2515);
and U3816 (N_3816,N_2667,N_2347);
xnor U3817 (N_3817,N_2604,N_2400);
xnor U3818 (N_3818,N_2960,N_2364);
and U3819 (N_3819,N_2552,N_2140);
and U3820 (N_3820,N_2919,N_2698);
and U3821 (N_3821,N_2887,N_2175);
nand U3822 (N_3822,N_2757,N_2913);
nand U3823 (N_3823,N_2097,N_2570);
or U3824 (N_3824,N_2912,N_2689);
xor U3825 (N_3825,N_2590,N_2274);
nand U3826 (N_3826,N_2061,N_2636);
nand U3827 (N_3827,N_2319,N_2808);
or U3828 (N_3828,N_2661,N_2737);
xor U3829 (N_3829,N_2667,N_2258);
nor U3830 (N_3830,N_2015,N_2424);
nor U3831 (N_3831,N_2316,N_2261);
xor U3832 (N_3832,N_2609,N_2056);
xor U3833 (N_3833,N_2338,N_2480);
nor U3834 (N_3834,N_2606,N_2200);
and U3835 (N_3835,N_2405,N_2926);
xnor U3836 (N_3836,N_2936,N_2786);
nor U3837 (N_3837,N_2782,N_2327);
nand U3838 (N_3838,N_2084,N_2587);
nand U3839 (N_3839,N_2562,N_2574);
or U3840 (N_3840,N_2144,N_2990);
or U3841 (N_3841,N_2100,N_2415);
nor U3842 (N_3842,N_2724,N_2943);
or U3843 (N_3843,N_2668,N_2007);
and U3844 (N_3844,N_2975,N_2417);
nand U3845 (N_3845,N_2771,N_2248);
and U3846 (N_3846,N_2295,N_2954);
nand U3847 (N_3847,N_2356,N_2719);
nor U3848 (N_3848,N_2862,N_2245);
nand U3849 (N_3849,N_2619,N_2609);
nor U3850 (N_3850,N_2154,N_2028);
xor U3851 (N_3851,N_2594,N_2690);
or U3852 (N_3852,N_2762,N_2454);
nor U3853 (N_3853,N_2334,N_2536);
and U3854 (N_3854,N_2933,N_2218);
and U3855 (N_3855,N_2578,N_2247);
and U3856 (N_3856,N_2864,N_2428);
or U3857 (N_3857,N_2573,N_2590);
nor U3858 (N_3858,N_2316,N_2697);
nor U3859 (N_3859,N_2437,N_2532);
or U3860 (N_3860,N_2667,N_2205);
xnor U3861 (N_3861,N_2785,N_2827);
nand U3862 (N_3862,N_2608,N_2698);
nor U3863 (N_3863,N_2072,N_2670);
nand U3864 (N_3864,N_2645,N_2491);
or U3865 (N_3865,N_2362,N_2695);
nand U3866 (N_3866,N_2639,N_2757);
or U3867 (N_3867,N_2540,N_2866);
or U3868 (N_3868,N_2458,N_2960);
or U3869 (N_3869,N_2839,N_2540);
nor U3870 (N_3870,N_2353,N_2100);
and U3871 (N_3871,N_2252,N_2072);
xor U3872 (N_3872,N_2977,N_2070);
or U3873 (N_3873,N_2041,N_2511);
nand U3874 (N_3874,N_2192,N_2918);
nand U3875 (N_3875,N_2658,N_2528);
nor U3876 (N_3876,N_2796,N_2744);
and U3877 (N_3877,N_2985,N_2319);
or U3878 (N_3878,N_2205,N_2749);
or U3879 (N_3879,N_2282,N_2452);
nand U3880 (N_3880,N_2496,N_2882);
xor U3881 (N_3881,N_2814,N_2230);
and U3882 (N_3882,N_2219,N_2159);
nor U3883 (N_3883,N_2168,N_2320);
or U3884 (N_3884,N_2754,N_2477);
nand U3885 (N_3885,N_2683,N_2982);
or U3886 (N_3886,N_2440,N_2716);
or U3887 (N_3887,N_2895,N_2189);
nand U3888 (N_3888,N_2127,N_2100);
xor U3889 (N_3889,N_2324,N_2140);
or U3890 (N_3890,N_2929,N_2922);
nand U3891 (N_3891,N_2627,N_2503);
nor U3892 (N_3892,N_2462,N_2729);
xnor U3893 (N_3893,N_2914,N_2625);
nand U3894 (N_3894,N_2039,N_2155);
xnor U3895 (N_3895,N_2833,N_2382);
nand U3896 (N_3896,N_2174,N_2223);
or U3897 (N_3897,N_2598,N_2765);
nor U3898 (N_3898,N_2326,N_2452);
xnor U3899 (N_3899,N_2166,N_2528);
nand U3900 (N_3900,N_2055,N_2704);
nor U3901 (N_3901,N_2287,N_2828);
nor U3902 (N_3902,N_2444,N_2090);
nor U3903 (N_3903,N_2540,N_2362);
xnor U3904 (N_3904,N_2938,N_2511);
xnor U3905 (N_3905,N_2734,N_2365);
and U3906 (N_3906,N_2555,N_2885);
nand U3907 (N_3907,N_2822,N_2168);
nand U3908 (N_3908,N_2484,N_2198);
xor U3909 (N_3909,N_2478,N_2986);
or U3910 (N_3910,N_2616,N_2650);
and U3911 (N_3911,N_2041,N_2325);
nor U3912 (N_3912,N_2546,N_2572);
and U3913 (N_3913,N_2291,N_2827);
nand U3914 (N_3914,N_2112,N_2512);
and U3915 (N_3915,N_2910,N_2735);
xor U3916 (N_3916,N_2012,N_2097);
xor U3917 (N_3917,N_2043,N_2080);
xor U3918 (N_3918,N_2489,N_2996);
nand U3919 (N_3919,N_2125,N_2601);
xor U3920 (N_3920,N_2203,N_2926);
nand U3921 (N_3921,N_2413,N_2194);
nor U3922 (N_3922,N_2409,N_2742);
nand U3923 (N_3923,N_2871,N_2427);
or U3924 (N_3924,N_2571,N_2250);
nand U3925 (N_3925,N_2120,N_2818);
xor U3926 (N_3926,N_2112,N_2550);
xor U3927 (N_3927,N_2399,N_2655);
nor U3928 (N_3928,N_2407,N_2558);
or U3929 (N_3929,N_2254,N_2782);
and U3930 (N_3930,N_2309,N_2973);
or U3931 (N_3931,N_2076,N_2801);
nor U3932 (N_3932,N_2211,N_2931);
and U3933 (N_3933,N_2437,N_2317);
nor U3934 (N_3934,N_2557,N_2726);
nor U3935 (N_3935,N_2917,N_2881);
and U3936 (N_3936,N_2138,N_2552);
nand U3937 (N_3937,N_2593,N_2416);
or U3938 (N_3938,N_2065,N_2144);
xor U3939 (N_3939,N_2774,N_2952);
nand U3940 (N_3940,N_2302,N_2829);
or U3941 (N_3941,N_2211,N_2733);
nand U3942 (N_3942,N_2348,N_2974);
nand U3943 (N_3943,N_2444,N_2833);
or U3944 (N_3944,N_2627,N_2192);
or U3945 (N_3945,N_2851,N_2426);
xor U3946 (N_3946,N_2336,N_2377);
nand U3947 (N_3947,N_2220,N_2630);
and U3948 (N_3948,N_2642,N_2352);
nor U3949 (N_3949,N_2117,N_2339);
nor U3950 (N_3950,N_2095,N_2910);
nand U3951 (N_3951,N_2475,N_2721);
nand U3952 (N_3952,N_2908,N_2670);
and U3953 (N_3953,N_2424,N_2342);
xor U3954 (N_3954,N_2460,N_2700);
nand U3955 (N_3955,N_2047,N_2760);
and U3956 (N_3956,N_2297,N_2309);
and U3957 (N_3957,N_2268,N_2065);
nor U3958 (N_3958,N_2105,N_2991);
and U3959 (N_3959,N_2588,N_2933);
and U3960 (N_3960,N_2766,N_2500);
nor U3961 (N_3961,N_2979,N_2691);
xnor U3962 (N_3962,N_2488,N_2088);
xor U3963 (N_3963,N_2399,N_2419);
nand U3964 (N_3964,N_2186,N_2719);
nor U3965 (N_3965,N_2698,N_2494);
nor U3966 (N_3966,N_2243,N_2628);
and U3967 (N_3967,N_2618,N_2986);
nand U3968 (N_3968,N_2957,N_2348);
nand U3969 (N_3969,N_2041,N_2166);
nand U3970 (N_3970,N_2930,N_2332);
nor U3971 (N_3971,N_2089,N_2496);
and U3972 (N_3972,N_2800,N_2927);
nand U3973 (N_3973,N_2700,N_2468);
xnor U3974 (N_3974,N_2488,N_2880);
and U3975 (N_3975,N_2794,N_2019);
or U3976 (N_3976,N_2847,N_2022);
or U3977 (N_3977,N_2603,N_2984);
nor U3978 (N_3978,N_2406,N_2096);
and U3979 (N_3979,N_2287,N_2013);
nor U3980 (N_3980,N_2415,N_2275);
nand U3981 (N_3981,N_2245,N_2836);
xor U3982 (N_3982,N_2978,N_2994);
nor U3983 (N_3983,N_2540,N_2143);
and U3984 (N_3984,N_2936,N_2269);
or U3985 (N_3985,N_2540,N_2080);
xnor U3986 (N_3986,N_2276,N_2422);
and U3987 (N_3987,N_2375,N_2524);
nor U3988 (N_3988,N_2929,N_2932);
xnor U3989 (N_3989,N_2789,N_2832);
nand U3990 (N_3990,N_2051,N_2879);
nor U3991 (N_3991,N_2117,N_2033);
nor U3992 (N_3992,N_2444,N_2376);
nor U3993 (N_3993,N_2081,N_2826);
nand U3994 (N_3994,N_2526,N_2135);
nor U3995 (N_3995,N_2604,N_2029);
xor U3996 (N_3996,N_2426,N_2176);
xnor U3997 (N_3997,N_2713,N_2256);
or U3998 (N_3998,N_2964,N_2909);
or U3999 (N_3999,N_2885,N_2288);
nor U4000 (N_4000,N_3012,N_3945);
nor U4001 (N_4001,N_3070,N_3785);
nor U4002 (N_4002,N_3352,N_3601);
xor U4003 (N_4003,N_3103,N_3984);
xnor U4004 (N_4004,N_3048,N_3738);
nand U4005 (N_4005,N_3681,N_3983);
or U4006 (N_4006,N_3504,N_3730);
nand U4007 (N_4007,N_3162,N_3752);
nand U4008 (N_4008,N_3028,N_3694);
xnor U4009 (N_4009,N_3045,N_3650);
nand U4010 (N_4010,N_3896,N_3203);
nand U4011 (N_4011,N_3724,N_3978);
nor U4012 (N_4012,N_3033,N_3473);
nand U4013 (N_4013,N_3538,N_3566);
or U4014 (N_4014,N_3409,N_3178);
and U4015 (N_4015,N_3112,N_3800);
nand U4016 (N_4016,N_3116,N_3884);
or U4017 (N_4017,N_3224,N_3902);
nor U4018 (N_4018,N_3961,N_3227);
and U4019 (N_4019,N_3964,N_3057);
or U4020 (N_4020,N_3361,N_3561);
nand U4021 (N_4021,N_3830,N_3758);
xnor U4022 (N_4022,N_3906,N_3963);
nand U4023 (N_4023,N_3153,N_3711);
nor U4024 (N_4024,N_3856,N_3069);
and U4025 (N_4025,N_3787,N_3250);
or U4026 (N_4026,N_3607,N_3438);
xnor U4027 (N_4027,N_3167,N_3705);
and U4028 (N_4028,N_3560,N_3622);
nor U4029 (N_4029,N_3736,N_3096);
and U4030 (N_4030,N_3129,N_3570);
xor U4031 (N_4031,N_3229,N_3633);
nand U4032 (N_4032,N_3986,N_3833);
nand U4033 (N_4033,N_3423,N_3547);
xor U4034 (N_4034,N_3443,N_3992);
or U4035 (N_4035,N_3185,N_3389);
and U4036 (N_4036,N_3578,N_3075);
xor U4037 (N_4037,N_3631,N_3590);
or U4038 (N_4038,N_3756,N_3411);
xnor U4039 (N_4039,N_3287,N_3598);
and U4040 (N_4040,N_3994,N_3357);
nand U4041 (N_4041,N_3059,N_3067);
nand U4042 (N_4042,N_3559,N_3356);
xor U4043 (N_4043,N_3524,N_3933);
nor U4044 (N_4044,N_3776,N_3662);
and U4045 (N_4045,N_3737,N_3646);
nand U4046 (N_4046,N_3380,N_3119);
or U4047 (N_4047,N_3377,N_3821);
or U4048 (N_4048,N_3217,N_3324);
nor U4049 (N_4049,N_3759,N_3915);
nand U4050 (N_4050,N_3818,N_3859);
xor U4051 (N_4051,N_3734,N_3778);
or U4052 (N_4052,N_3422,N_3703);
or U4053 (N_4053,N_3874,N_3797);
and U4054 (N_4054,N_3184,N_3247);
nand U4055 (N_4055,N_3231,N_3729);
xnor U4056 (N_4056,N_3472,N_3238);
and U4057 (N_4057,N_3009,N_3495);
nand U4058 (N_4058,N_3670,N_3755);
nor U4059 (N_4059,N_3304,N_3201);
and U4060 (N_4060,N_3366,N_3228);
nand U4061 (N_4061,N_3824,N_3853);
nor U4062 (N_4062,N_3714,N_3880);
nand U4063 (N_4063,N_3801,N_3505);
or U4064 (N_4064,N_3054,N_3867);
nand U4065 (N_4065,N_3010,N_3501);
nand U4066 (N_4066,N_3465,N_3279);
xor U4067 (N_4067,N_3487,N_3606);
and U4068 (N_4068,N_3000,N_3368);
xor U4069 (N_4069,N_3689,N_3490);
nand U4070 (N_4070,N_3225,N_3174);
or U4071 (N_4071,N_3353,N_3351);
and U4072 (N_4072,N_3691,N_3795);
nand U4073 (N_4073,N_3100,N_3466);
nor U4074 (N_4074,N_3843,N_3222);
or U4075 (N_4075,N_3249,N_3521);
nand U4076 (N_4076,N_3006,N_3783);
and U4077 (N_4077,N_3491,N_3136);
nand U4078 (N_4078,N_3403,N_3323);
and U4079 (N_4079,N_3642,N_3927);
or U4080 (N_4080,N_3733,N_3643);
nor U4081 (N_4081,N_3047,N_3897);
xor U4082 (N_4082,N_3557,N_3692);
or U4083 (N_4083,N_3367,N_3617);
nand U4084 (N_4084,N_3823,N_3725);
nor U4085 (N_4085,N_3866,N_3111);
and U4086 (N_4086,N_3651,N_3040);
xnor U4087 (N_4087,N_3518,N_3425);
nor U4088 (N_4088,N_3256,N_3087);
xor U4089 (N_4089,N_3898,N_3804);
and U4090 (N_4090,N_3799,N_3344);
xnor U4091 (N_4091,N_3298,N_3637);
nor U4092 (N_4092,N_3158,N_3142);
or U4093 (N_4093,N_3499,N_3159);
nor U4094 (N_4094,N_3267,N_3126);
nand U4095 (N_4095,N_3663,N_3290);
nand U4096 (N_4096,N_3816,N_3084);
xor U4097 (N_4097,N_3550,N_3342);
nor U4098 (N_4098,N_3675,N_3770);
and U4099 (N_4099,N_3468,N_3132);
xor U4100 (N_4100,N_3782,N_3024);
nand U4101 (N_4101,N_3751,N_3749);
or U4102 (N_4102,N_3372,N_3831);
xnor U4103 (N_4103,N_3620,N_3464);
nor U4104 (N_4104,N_3427,N_3001);
nor U4105 (N_4105,N_3396,N_3318);
nand U4106 (N_4106,N_3168,N_3194);
and U4107 (N_4107,N_3043,N_3810);
nand U4108 (N_4108,N_3282,N_3241);
or U4109 (N_4109,N_3808,N_3876);
nand U4110 (N_4110,N_3710,N_3712);
xor U4111 (N_4111,N_3364,N_3039);
and U4112 (N_4112,N_3430,N_3450);
xor U4113 (N_4113,N_3102,N_3190);
and U4114 (N_4114,N_3922,N_3615);
and U4115 (N_4115,N_3664,N_3672);
nand U4116 (N_4116,N_3264,N_3721);
and U4117 (N_4117,N_3176,N_3164);
or U4118 (N_4118,N_3996,N_3894);
nand U4119 (N_4119,N_3972,N_3037);
xnor U4120 (N_4120,N_3639,N_3141);
xnor U4121 (N_4121,N_3358,N_3846);
xnor U4122 (N_4122,N_3858,N_3294);
xnor U4123 (N_4123,N_3932,N_3875);
and U4124 (N_4124,N_3883,N_3826);
nor U4125 (N_4125,N_3786,N_3827);
nand U4126 (N_4126,N_3143,N_3791);
nand U4127 (N_4127,N_3273,N_3426);
or U4128 (N_4128,N_3117,N_3979);
or U4129 (N_4129,N_3726,N_3140);
and U4130 (N_4130,N_3708,N_3431);
nor U4131 (N_4131,N_3486,N_3837);
xnor U4132 (N_4132,N_3391,N_3613);
xor U4133 (N_4133,N_3289,N_3952);
nand U4134 (N_4134,N_3108,N_3763);
xnor U4135 (N_4135,N_3101,N_3929);
nor U4136 (N_4136,N_3137,N_3072);
and U4137 (N_4137,N_3240,N_3453);
and U4138 (N_4138,N_3610,N_3947);
and U4139 (N_4139,N_3232,N_3154);
xor U4140 (N_4140,N_3761,N_3854);
xnor U4141 (N_4141,N_3905,N_3397);
or U4142 (N_4142,N_3700,N_3481);
and U4143 (N_4143,N_3839,N_3540);
or U4144 (N_4144,N_3326,N_3196);
xor U4145 (N_4145,N_3461,N_3005);
or U4146 (N_4146,N_3098,N_3571);
or U4147 (N_4147,N_3625,N_3888);
xnor U4148 (N_4148,N_3525,N_3363);
nand U4149 (N_4149,N_3206,N_3113);
nor U4150 (N_4150,N_3115,N_3599);
xor U4151 (N_4151,N_3032,N_3446);
nand U4152 (N_4152,N_3221,N_3912);
nor U4153 (N_4153,N_3569,N_3017);
or U4154 (N_4154,N_3161,N_3666);
nand U4155 (N_4155,N_3056,N_3781);
or U4156 (N_4156,N_3616,N_3698);
xnor U4157 (N_4157,N_3375,N_3951);
nor U4158 (N_4158,N_3647,N_3895);
and U4159 (N_4159,N_3489,N_3448);
and U4160 (N_4160,N_3765,N_3857);
and U4161 (N_4161,N_3415,N_3845);
xnor U4162 (N_4162,N_3748,N_3311);
and U4163 (N_4163,N_3935,N_3667);
nand U4164 (N_4164,N_3439,N_3175);
and U4165 (N_4165,N_3893,N_3385);
nor U4166 (N_4166,N_3274,N_3627);
nor U4167 (N_4167,N_3302,N_3528);
nand U4168 (N_4168,N_3124,N_3676);
nand U4169 (N_4169,N_3388,N_3003);
and U4170 (N_4170,N_3587,N_3440);
or U4171 (N_4171,N_3496,N_3412);
nor U4172 (N_4172,N_3974,N_3508);
or U4173 (N_4173,N_3657,N_3924);
nand U4174 (N_4174,N_3624,N_3475);
and U4175 (N_4175,N_3923,N_3469);
nand U4176 (N_4176,N_3970,N_3339);
xor U4177 (N_4177,N_3930,N_3463);
nor U4178 (N_4178,N_3235,N_3063);
nor U4179 (N_4179,N_3429,N_3960);
nand U4180 (N_4180,N_3456,N_3152);
nor U4181 (N_4181,N_3413,N_3621);
and U4182 (N_4182,N_3903,N_3855);
and U4183 (N_4183,N_3322,N_3731);
and U4184 (N_4184,N_3519,N_3399);
and U4185 (N_4185,N_3648,N_3901);
xor U4186 (N_4186,N_3913,N_3707);
or U4187 (N_4187,N_3041,N_3139);
nand U4188 (N_4188,N_3940,N_3805);
and U4189 (N_4189,N_3515,N_3661);
xor U4190 (N_4190,N_3343,N_3219);
xor U4191 (N_4191,N_3026,N_3534);
xor U4192 (N_4192,N_3205,N_3565);
nor U4193 (N_4193,N_3654,N_3788);
and U4194 (N_4194,N_3767,N_3938);
nor U4195 (N_4195,N_3742,N_3746);
xor U4196 (N_4196,N_3673,N_3555);
or U4197 (N_4197,N_3146,N_3634);
nor U4198 (N_4198,N_3744,N_3248);
and U4199 (N_4199,N_3183,N_3309);
nor U4200 (N_4200,N_3644,N_3236);
nand U4201 (N_4201,N_3189,N_3636);
nand U4202 (N_4202,N_3815,N_3580);
or U4203 (N_4203,N_3813,N_3659);
nor U4204 (N_4204,N_3275,N_3739);
nand U4205 (N_4205,N_3046,N_3207);
nand U4206 (N_4206,N_3197,N_3085);
and U4207 (N_4207,N_3680,N_3990);
and U4208 (N_4208,N_3702,N_3995);
and U4209 (N_4209,N_3460,N_3128);
nand U4210 (N_4210,N_3471,N_3878);
and U4211 (N_4211,N_3891,N_3114);
nand U4212 (N_4212,N_3576,N_3334);
nand U4213 (N_4213,N_3595,N_3941);
and U4214 (N_4214,N_3445,N_3498);
or U4215 (N_4215,N_3918,N_3243);
nor U4216 (N_4216,N_3629,N_3757);
and U4217 (N_4217,N_3864,N_3474);
nand U4218 (N_4218,N_3280,N_3150);
xnor U4219 (N_4219,N_3536,N_3562);
nand U4220 (N_4220,N_3244,N_3436);
and U4221 (N_4221,N_3572,N_3946);
and U4222 (N_4222,N_3485,N_3532);
and U4223 (N_4223,N_3747,N_3683);
or U4224 (N_4224,N_3283,N_3220);
xnor U4225 (N_4225,N_3467,N_3626);
nor U4226 (N_4226,N_3568,N_3779);
nand U4227 (N_4227,N_3789,N_3957);
xnor U4228 (N_4228,N_3278,N_3899);
and U4229 (N_4229,N_3817,N_3764);
nand U4230 (N_4230,N_3277,N_3081);
nor U4231 (N_4231,N_3286,N_3589);
or U4232 (N_4232,N_3198,N_3774);
nor U4233 (N_4233,N_3709,N_3181);
and U4234 (N_4234,N_3186,N_3768);
and U4235 (N_4235,N_3271,N_3812);
xnor U4236 (N_4236,N_3674,N_3687);
or U4237 (N_4237,N_3792,N_3382);
or U4238 (N_4238,N_3192,N_3863);
nand U4239 (N_4239,N_3936,N_3985);
xor U4240 (N_4240,N_3969,N_3074);
nor U4241 (N_4241,N_3829,N_3596);
nor U4242 (N_4242,N_3999,N_3819);
and U4243 (N_4243,N_3263,N_3612);
nand U4244 (N_4244,N_3981,N_3349);
and U4245 (N_4245,N_3753,N_3144);
xnor U4246 (N_4246,N_3355,N_3226);
or U4247 (N_4247,N_3060,N_3347);
and U4248 (N_4248,N_3061,N_3807);
nor U4249 (N_4249,N_3488,N_3890);
nor U4250 (N_4250,N_3077,N_3345);
xor U4251 (N_4251,N_3021,N_3825);
and U4252 (N_4252,N_3771,N_3877);
xor U4253 (N_4253,N_3563,N_3530);
nor U4254 (N_4254,N_3165,N_3310);
nor U4255 (N_4255,N_3257,N_3766);
and U4256 (N_4256,N_3105,N_3531);
and U4257 (N_4257,N_3020,N_3400);
or U4258 (N_4258,N_3954,N_3038);
nand U4259 (N_4259,N_3847,N_3370);
and U4260 (N_4260,N_3512,N_3640);
nand U4261 (N_4261,N_3394,N_3328);
nand U4262 (N_4262,N_3953,N_3959);
nand U4263 (N_4263,N_3420,N_3234);
nand U4264 (N_4264,N_3171,N_3262);
nor U4265 (N_4265,N_3457,N_3193);
xor U4266 (N_4266,N_3732,N_3567);
xor U4267 (N_4267,N_3015,N_3007);
nand U4268 (N_4268,N_3494,N_3870);
nand U4269 (N_4269,N_3684,N_3034);
and U4270 (N_4270,N_3329,N_3838);
and U4271 (N_4271,N_3321,N_3796);
nor U4272 (N_4272,N_3369,N_3239);
xnor U4273 (N_4273,N_3073,N_3018);
nand U4274 (N_4274,N_3522,N_3359);
nor U4275 (N_4275,N_3579,N_3251);
nor U4276 (N_4276,N_3374,N_3254);
or U4277 (N_4277,N_3583,N_3089);
or U4278 (N_4278,N_3402,N_3123);
xnor U4279 (N_4279,N_3641,N_3188);
xnor U4280 (N_4280,N_3078,N_3166);
xnor U4281 (N_4281,N_3862,N_3083);
nand U4282 (N_4282,N_3973,N_3305);
nor U4283 (N_4283,N_3545,N_3451);
and U4284 (N_4284,N_3079,N_3348);
xnor U4285 (N_4285,N_3346,N_3836);
and U4286 (N_4286,N_3437,N_3179);
nor U4287 (N_4287,N_3029,N_3265);
or U4288 (N_4288,N_3118,N_3916);
nor U4289 (N_4289,N_3956,N_3245);
nand U4290 (N_4290,N_3506,N_3065);
or U4291 (N_4291,N_3741,N_3517);
xor U4292 (N_4292,N_3597,N_3772);
nand U4293 (N_4293,N_3281,N_3331);
or U4294 (N_4294,N_3852,N_3784);
xnor U4295 (N_4295,N_3909,N_3134);
nor U4296 (N_4296,N_3419,N_3529);
or U4297 (N_4297,N_3030,N_3145);
nand U4298 (N_4298,N_3503,N_3255);
xor U4299 (N_4299,N_3887,N_3130);
or U4300 (N_4300,N_3308,N_3713);
and U4301 (N_4301,N_3301,N_3080);
xnor U4302 (N_4302,N_3449,N_3454);
nor U4303 (N_4303,N_3276,N_3542);
xnor U4304 (N_4304,N_3881,N_3628);
xor U4305 (N_4305,N_3340,N_3803);
and U4306 (N_4306,N_3320,N_3968);
or U4307 (N_4307,N_3050,N_3076);
or U4308 (N_4308,N_3051,N_3966);
or U4309 (N_4309,N_3293,N_3148);
nor U4310 (N_4310,N_3693,N_3980);
nand U4311 (N_4311,N_3019,N_3258);
xnor U4312 (N_4312,N_3811,N_3333);
nand U4313 (N_4313,N_3588,N_3407);
and U4314 (N_4314,N_3987,N_3976);
nor U4315 (N_4315,N_3291,N_3790);
and U4316 (N_4316,N_3434,N_3169);
nor U4317 (N_4317,N_3209,N_3520);
nand U4318 (N_4318,N_3548,N_3025);
nand U4319 (N_4319,N_3760,N_3036);
and U4320 (N_4320,N_3350,N_3093);
and U4321 (N_4321,N_3338,N_3327);
nor U4322 (N_4322,N_3246,N_3086);
nor U4323 (N_4323,N_3828,N_3109);
nor U4324 (N_4324,N_3092,N_3398);
and U4325 (N_4325,N_3510,N_3948);
and U4326 (N_4326,N_3163,N_3848);
xnor U4327 (N_4327,N_3851,N_3989);
and U4328 (N_4328,N_3421,N_3762);
nor U4329 (N_4329,N_3135,N_3653);
nor U4330 (N_4330,N_3266,N_3920);
nand U4331 (N_4331,N_3717,N_3172);
xnor U4332 (N_4332,N_3410,N_3546);
nor U4333 (N_4333,N_3997,N_3885);
nand U4334 (N_4334,N_3720,N_3406);
or U4335 (N_4335,N_3850,N_3458);
or U4336 (N_4336,N_3660,N_3216);
or U4337 (N_4337,N_3949,N_3042);
or U4338 (N_4338,N_3022,N_3478);
or U4339 (N_4339,N_3950,N_3230);
nand U4340 (N_4340,N_3998,N_3261);
and U4341 (N_4341,N_3424,N_3392);
or U4342 (N_4342,N_3535,N_3253);
or U4343 (N_4343,N_3943,N_3719);
or U4344 (N_4344,N_3182,N_3270);
xnor U4345 (N_4345,N_3873,N_3330);
nand U4346 (N_4346,N_3002,N_3064);
or U4347 (N_4347,N_3872,N_3649);
or U4348 (N_4348,N_3669,N_3455);
or U4349 (N_4349,N_3476,N_3295);
nor U4350 (N_4350,N_3284,N_3242);
or U4351 (N_4351,N_3543,N_3509);
nand U4352 (N_4352,N_3632,N_3053);
nand U4353 (N_4353,N_3016,N_3865);
or U4354 (N_4354,N_3671,N_3630);
nand U4355 (N_4355,N_3993,N_3104);
xor U4356 (N_4356,N_3917,N_3582);
and U4357 (N_4357,N_3581,N_3655);
nand U4358 (N_4358,N_3470,N_3099);
or U4359 (N_4359,N_3317,N_3527);
nor U4360 (N_4360,N_3868,N_3593);
xor U4361 (N_4361,N_3871,N_3337);
nor U4362 (N_4362,N_3919,N_3091);
nor U4363 (N_4363,N_3841,N_3665);
xnor U4364 (N_4364,N_3611,N_3939);
and U4365 (N_4365,N_3614,N_3210);
or U4366 (N_4366,N_3414,N_3011);
and U4367 (N_4367,N_3603,N_3395);
nand U4368 (N_4368,N_3780,N_3507);
and U4369 (N_4369,N_3214,N_3658);
xor U4370 (N_4370,N_3052,N_3180);
and U4371 (N_4371,N_3944,N_3699);
or U4372 (N_4372,N_3727,N_3055);
and U4373 (N_4373,N_3432,N_3695);
nor U4374 (N_4374,N_3312,N_3444);
and U4375 (N_4375,N_3701,N_3911);
nor U4376 (N_4376,N_3259,N_3500);
xor U4377 (N_4377,N_3237,N_3967);
or U4378 (N_4378,N_3325,N_3442);
or U4379 (N_4379,N_3023,N_3299);
xnor U4380 (N_4380,N_3552,N_3482);
nor U4381 (N_4381,N_3840,N_3594);
or U4382 (N_4382,N_3218,N_3716);
nand U4383 (N_4383,N_3832,N_3386);
and U4384 (N_4384,N_3558,N_3549);
nor U4385 (N_4385,N_3435,N_3638);
nor U4386 (N_4386,N_3769,N_3131);
nand U4387 (N_4387,N_3914,N_3750);
nand U4388 (N_4388,N_3269,N_3497);
or U4389 (N_4389,N_3288,N_3513);
and U4390 (N_4390,N_3441,N_3044);
nand U4391 (N_4391,N_3354,N_3988);
or U4392 (N_4392,N_3537,N_3834);
nor U4393 (N_4393,N_3121,N_3127);
or U4394 (N_4394,N_3608,N_3635);
nor U4395 (N_4395,N_3202,N_3907);
xor U4396 (N_4396,N_3155,N_3991);
and U4397 (N_4397,N_3199,N_3307);
nand U4398 (N_4398,N_3223,N_3160);
nor U4399 (N_4399,N_3493,N_3211);
and U4400 (N_4400,N_3685,N_3332);
nor U4401 (N_4401,N_3379,N_3384);
and U4402 (N_4402,N_3533,N_3605);
and U4403 (N_4403,N_3900,N_3904);
xor U4404 (N_4404,N_3822,N_3315);
nor U4405 (N_4405,N_3447,N_3802);
xnor U4406 (N_4406,N_3314,N_3013);
nor U4407 (N_4407,N_3842,N_3459);
or U4408 (N_4408,N_3008,N_3584);
xnor U4409 (N_4409,N_3926,N_3452);
nand U4410 (N_4410,N_3718,N_3609);
and U4411 (N_4411,N_3151,N_3319);
nand U4412 (N_4412,N_3715,N_3690);
and U4413 (N_4413,N_3004,N_3793);
nor U4414 (N_4414,N_3296,N_3173);
or U4415 (N_4415,N_3260,N_3931);
and U4416 (N_4416,N_3157,N_3068);
xnor U4417 (N_4417,N_3861,N_3416);
nor U4418 (N_4418,N_3585,N_3297);
and U4419 (N_4419,N_3097,N_3523);
nand U4420 (N_4420,N_3618,N_3303);
nor U4421 (N_4421,N_3806,N_3982);
or U4422 (N_4422,N_3300,N_3908);
and U4423 (N_4423,N_3604,N_3809);
or U4424 (N_4424,N_3735,N_3697);
xor U4425 (N_4425,N_3962,N_3365);
or U4426 (N_4426,N_3574,N_3600);
xnor U4427 (N_4427,N_3591,N_3728);
and U4428 (N_4428,N_3360,N_3492);
nor U4429 (N_4429,N_3682,N_3378);
xor U4430 (N_4430,N_3886,N_3285);
and U4431 (N_4431,N_3433,N_3937);
xnor U4432 (N_4432,N_3090,N_3928);
or U4433 (N_4433,N_3428,N_3213);
xnor U4434 (N_4434,N_3208,N_3526);
nor U4435 (N_4435,N_3942,N_3775);
and U4436 (N_4436,N_3313,N_3754);
xnor U4437 (N_4437,N_3740,N_3335);
nand U4438 (N_4438,N_3035,N_3479);
and U4439 (N_4439,N_3688,N_3484);
nand U4440 (N_4440,N_3882,N_3556);
or U4441 (N_4441,N_3773,N_3138);
and U4442 (N_4442,N_3170,N_3195);
xnor U4443 (N_4443,N_3514,N_3149);
nor U4444 (N_4444,N_3212,N_3272);
and U4445 (N_4445,N_3577,N_3652);
or U4446 (N_4446,N_3575,N_3417);
or U4447 (N_4447,N_3551,N_3110);
nor U4448 (N_4448,N_3677,N_3058);
nand U4449 (N_4449,N_3156,N_3133);
nand U4450 (N_4450,N_3373,N_3921);
nor U4451 (N_4451,N_3879,N_3200);
nand U4452 (N_4452,N_3745,N_3623);
and U4453 (N_4453,N_3204,N_3462);
nor U4454 (N_4454,N_3722,N_3958);
nand U4455 (N_4455,N_3706,N_3592);
nand U4456 (N_4456,N_3849,N_3602);
and U4457 (N_4457,N_3820,N_3686);
and U4458 (N_4458,N_3066,N_3934);
or U4459 (N_4459,N_3723,N_3656);
and U4460 (N_4460,N_3404,N_3645);
nor U4461 (N_4461,N_3122,N_3798);
xor U4462 (N_4462,N_3147,N_3107);
xor U4463 (N_4463,N_3477,N_3120);
and U4464 (N_4464,N_3955,N_3027);
or U4465 (N_4465,N_3376,N_3977);
or U4466 (N_4466,N_3553,N_3668);
nor U4467 (N_4467,N_3362,N_3777);
or U4468 (N_4468,N_3844,N_3619);
nor U4469 (N_4469,N_3088,N_3252);
or U4470 (N_4470,N_3586,N_3975);
or U4471 (N_4471,N_3405,N_3704);
xor U4472 (N_4472,N_3125,N_3062);
xor U4473 (N_4473,N_3292,N_3965);
xnor U4474 (N_4474,N_3187,N_3215);
or U4475 (N_4475,N_3268,N_3480);
or U4476 (N_4476,N_3860,N_3925);
xnor U4477 (N_4477,N_3106,N_3316);
nor U4478 (N_4478,N_3554,N_3341);
and U4479 (N_4479,N_3336,N_3511);
nor U4480 (N_4480,N_3393,N_3971);
nor U4481 (N_4481,N_3049,N_3835);
and U4482 (N_4482,N_3573,N_3516);
or U4483 (N_4483,N_3306,N_3483);
nor U4484 (N_4484,N_3696,N_3889);
and U4485 (N_4485,N_3892,N_3390);
and U4486 (N_4486,N_3743,N_3094);
or U4487 (N_4487,N_3071,N_3177);
and U4488 (N_4488,N_3381,N_3418);
and U4489 (N_4489,N_3539,N_3678);
or U4490 (N_4490,N_3082,N_3910);
and U4491 (N_4491,N_3541,N_3502);
xor U4492 (N_4492,N_3408,N_3869);
and U4493 (N_4493,N_3014,N_3233);
nor U4494 (N_4494,N_3371,N_3794);
nor U4495 (N_4495,N_3387,N_3401);
and U4496 (N_4496,N_3191,N_3814);
or U4497 (N_4497,N_3383,N_3544);
nor U4498 (N_4498,N_3564,N_3679);
xor U4499 (N_4499,N_3095,N_3031);
nand U4500 (N_4500,N_3074,N_3055);
and U4501 (N_4501,N_3399,N_3097);
or U4502 (N_4502,N_3983,N_3426);
nand U4503 (N_4503,N_3599,N_3399);
xor U4504 (N_4504,N_3962,N_3336);
nand U4505 (N_4505,N_3722,N_3019);
nor U4506 (N_4506,N_3339,N_3803);
and U4507 (N_4507,N_3073,N_3767);
or U4508 (N_4508,N_3258,N_3010);
and U4509 (N_4509,N_3716,N_3826);
and U4510 (N_4510,N_3050,N_3638);
nand U4511 (N_4511,N_3113,N_3004);
xnor U4512 (N_4512,N_3751,N_3329);
nor U4513 (N_4513,N_3878,N_3752);
nand U4514 (N_4514,N_3794,N_3119);
or U4515 (N_4515,N_3655,N_3190);
nor U4516 (N_4516,N_3338,N_3599);
nand U4517 (N_4517,N_3559,N_3613);
nor U4518 (N_4518,N_3297,N_3780);
or U4519 (N_4519,N_3535,N_3437);
and U4520 (N_4520,N_3483,N_3543);
or U4521 (N_4521,N_3677,N_3236);
and U4522 (N_4522,N_3587,N_3232);
xnor U4523 (N_4523,N_3799,N_3770);
nor U4524 (N_4524,N_3262,N_3589);
xor U4525 (N_4525,N_3311,N_3146);
xnor U4526 (N_4526,N_3785,N_3972);
nor U4527 (N_4527,N_3782,N_3281);
and U4528 (N_4528,N_3855,N_3326);
and U4529 (N_4529,N_3822,N_3425);
nor U4530 (N_4530,N_3858,N_3388);
or U4531 (N_4531,N_3133,N_3842);
nand U4532 (N_4532,N_3511,N_3060);
or U4533 (N_4533,N_3158,N_3904);
or U4534 (N_4534,N_3516,N_3734);
and U4535 (N_4535,N_3921,N_3007);
nor U4536 (N_4536,N_3084,N_3966);
and U4537 (N_4537,N_3015,N_3269);
or U4538 (N_4538,N_3539,N_3409);
nor U4539 (N_4539,N_3692,N_3972);
nor U4540 (N_4540,N_3416,N_3988);
nand U4541 (N_4541,N_3210,N_3986);
nor U4542 (N_4542,N_3052,N_3165);
or U4543 (N_4543,N_3570,N_3285);
nor U4544 (N_4544,N_3455,N_3207);
or U4545 (N_4545,N_3525,N_3583);
xor U4546 (N_4546,N_3083,N_3427);
nand U4547 (N_4547,N_3470,N_3799);
or U4548 (N_4548,N_3171,N_3495);
nand U4549 (N_4549,N_3755,N_3284);
nor U4550 (N_4550,N_3423,N_3537);
nor U4551 (N_4551,N_3247,N_3485);
and U4552 (N_4552,N_3553,N_3090);
nor U4553 (N_4553,N_3069,N_3066);
and U4554 (N_4554,N_3875,N_3470);
xor U4555 (N_4555,N_3336,N_3063);
nand U4556 (N_4556,N_3501,N_3528);
xnor U4557 (N_4557,N_3382,N_3033);
xnor U4558 (N_4558,N_3516,N_3413);
nand U4559 (N_4559,N_3453,N_3062);
or U4560 (N_4560,N_3698,N_3464);
or U4561 (N_4561,N_3269,N_3678);
nor U4562 (N_4562,N_3105,N_3483);
xor U4563 (N_4563,N_3006,N_3423);
or U4564 (N_4564,N_3684,N_3231);
xnor U4565 (N_4565,N_3675,N_3328);
nor U4566 (N_4566,N_3782,N_3094);
xor U4567 (N_4567,N_3441,N_3594);
xnor U4568 (N_4568,N_3634,N_3993);
xnor U4569 (N_4569,N_3428,N_3239);
or U4570 (N_4570,N_3892,N_3490);
and U4571 (N_4571,N_3725,N_3822);
or U4572 (N_4572,N_3848,N_3192);
and U4573 (N_4573,N_3089,N_3873);
or U4574 (N_4574,N_3333,N_3030);
or U4575 (N_4575,N_3708,N_3933);
xnor U4576 (N_4576,N_3562,N_3059);
or U4577 (N_4577,N_3106,N_3598);
or U4578 (N_4578,N_3899,N_3910);
nand U4579 (N_4579,N_3411,N_3479);
and U4580 (N_4580,N_3373,N_3304);
or U4581 (N_4581,N_3484,N_3850);
and U4582 (N_4582,N_3908,N_3241);
or U4583 (N_4583,N_3179,N_3704);
and U4584 (N_4584,N_3508,N_3315);
nor U4585 (N_4585,N_3049,N_3536);
xnor U4586 (N_4586,N_3569,N_3044);
nand U4587 (N_4587,N_3486,N_3164);
and U4588 (N_4588,N_3596,N_3884);
nand U4589 (N_4589,N_3559,N_3616);
and U4590 (N_4590,N_3092,N_3815);
and U4591 (N_4591,N_3829,N_3184);
nand U4592 (N_4592,N_3159,N_3387);
nor U4593 (N_4593,N_3085,N_3322);
or U4594 (N_4594,N_3637,N_3131);
nor U4595 (N_4595,N_3171,N_3028);
nor U4596 (N_4596,N_3593,N_3909);
and U4597 (N_4597,N_3674,N_3464);
xnor U4598 (N_4598,N_3824,N_3997);
xor U4599 (N_4599,N_3783,N_3339);
or U4600 (N_4600,N_3827,N_3425);
or U4601 (N_4601,N_3908,N_3071);
nand U4602 (N_4602,N_3123,N_3645);
and U4603 (N_4603,N_3216,N_3361);
xnor U4604 (N_4604,N_3684,N_3142);
xnor U4605 (N_4605,N_3093,N_3986);
nor U4606 (N_4606,N_3302,N_3692);
nand U4607 (N_4607,N_3615,N_3541);
or U4608 (N_4608,N_3711,N_3114);
and U4609 (N_4609,N_3911,N_3102);
and U4610 (N_4610,N_3563,N_3588);
nand U4611 (N_4611,N_3492,N_3171);
and U4612 (N_4612,N_3074,N_3011);
and U4613 (N_4613,N_3555,N_3516);
xnor U4614 (N_4614,N_3606,N_3989);
nor U4615 (N_4615,N_3029,N_3146);
or U4616 (N_4616,N_3077,N_3812);
or U4617 (N_4617,N_3052,N_3990);
xnor U4618 (N_4618,N_3679,N_3996);
and U4619 (N_4619,N_3528,N_3333);
or U4620 (N_4620,N_3606,N_3153);
nor U4621 (N_4621,N_3148,N_3266);
and U4622 (N_4622,N_3730,N_3374);
nor U4623 (N_4623,N_3965,N_3695);
or U4624 (N_4624,N_3150,N_3326);
or U4625 (N_4625,N_3173,N_3153);
nand U4626 (N_4626,N_3084,N_3104);
and U4627 (N_4627,N_3342,N_3701);
or U4628 (N_4628,N_3492,N_3306);
xor U4629 (N_4629,N_3745,N_3129);
or U4630 (N_4630,N_3897,N_3436);
and U4631 (N_4631,N_3765,N_3888);
nand U4632 (N_4632,N_3521,N_3297);
nand U4633 (N_4633,N_3582,N_3122);
xnor U4634 (N_4634,N_3254,N_3990);
or U4635 (N_4635,N_3186,N_3866);
and U4636 (N_4636,N_3549,N_3371);
nor U4637 (N_4637,N_3788,N_3686);
or U4638 (N_4638,N_3745,N_3711);
nor U4639 (N_4639,N_3301,N_3746);
nand U4640 (N_4640,N_3890,N_3081);
and U4641 (N_4641,N_3558,N_3566);
xnor U4642 (N_4642,N_3176,N_3102);
nor U4643 (N_4643,N_3096,N_3429);
nand U4644 (N_4644,N_3927,N_3114);
nor U4645 (N_4645,N_3490,N_3150);
nor U4646 (N_4646,N_3010,N_3053);
xnor U4647 (N_4647,N_3651,N_3834);
nor U4648 (N_4648,N_3053,N_3771);
nand U4649 (N_4649,N_3981,N_3043);
and U4650 (N_4650,N_3544,N_3108);
and U4651 (N_4651,N_3452,N_3467);
and U4652 (N_4652,N_3637,N_3437);
nor U4653 (N_4653,N_3470,N_3926);
nor U4654 (N_4654,N_3481,N_3041);
nor U4655 (N_4655,N_3911,N_3487);
and U4656 (N_4656,N_3967,N_3287);
nor U4657 (N_4657,N_3041,N_3761);
and U4658 (N_4658,N_3611,N_3350);
nor U4659 (N_4659,N_3344,N_3946);
nor U4660 (N_4660,N_3665,N_3655);
or U4661 (N_4661,N_3527,N_3856);
or U4662 (N_4662,N_3960,N_3990);
and U4663 (N_4663,N_3481,N_3477);
nor U4664 (N_4664,N_3289,N_3584);
xnor U4665 (N_4665,N_3768,N_3359);
nand U4666 (N_4666,N_3393,N_3789);
nand U4667 (N_4667,N_3701,N_3470);
nor U4668 (N_4668,N_3271,N_3327);
nor U4669 (N_4669,N_3889,N_3856);
and U4670 (N_4670,N_3829,N_3562);
and U4671 (N_4671,N_3209,N_3833);
nor U4672 (N_4672,N_3261,N_3135);
xnor U4673 (N_4673,N_3477,N_3845);
and U4674 (N_4674,N_3139,N_3163);
or U4675 (N_4675,N_3657,N_3033);
or U4676 (N_4676,N_3941,N_3132);
and U4677 (N_4677,N_3755,N_3438);
nor U4678 (N_4678,N_3639,N_3081);
and U4679 (N_4679,N_3517,N_3659);
or U4680 (N_4680,N_3558,N_3533);
and U4681 (N_4681,N_3078,N_3752);
or U4682 (N_4682,N_3326,N_3950);
xor U4683 (N_4683,N_3752,N_3756);
nor U4684 (N_4684,N_3944,N_3219);
and U4685 (N_4685,N_3891,N_3307);
nor U4686 (N_4686,N_3257,N_3730);
or U4687 (N_4687,N_3439,N_3914);
and U4688 (N_4688,N_3734,N_3272);
or U4689 (N_4689,N_3739,N_3377);
nor U4690 (N_4690,N_3666,N_3657);
xor U4691 (N_4691,N_3606,N_3447);
nor U4692 (N_4692,N_3386,N_3248);
xnor U4693 (N_4693,N_3845,N_3032);
xor U4694 (N_4694,N_3570,N_3593);
or U4695 (N_4695,N_3292,N_3745);
and U4696 (N_4696,N_3572,N_3598);
xnor U4697 (N_4697,N_3453,N_3718);
and U4698 (N_4698,N_3510,N_3354);
nand U4699 (N_4699,N_3172,N_3642);
and U4700 (N_4700,N_3883,N_3703);
and U4701 (N_4701,N_3378,N_3128);
and U4702 (N_4702,N_3759,N_3318);
and U4703 (N_4703,N_3213,N_3431);
nor U4704 (N_4704,N_3886,N_3072);
or U4705 (N_4705,N_3570,N_3480);
nor U4706 (N_4706,N_3878,N_3161);
and U4707 (N_4707,N_3258,N_3163);
or U4708 (N_4708,N_3627,N_3430);
nor U4709 (N_4709,N_3738,N_3831);
and U4710 (N_4710,N_3347,N_3586);
nor U4711 (N_4711,N_3596,N_3564);
or U4712 (N_4712,N_3827,N_3296);
xor U4713 (N_4713,N_3245,N_3898);
nor U4714 (N_4714,N_3726,N_3016);
or U4715 (N_4715,N_3537,N_3742);
nor U4716 (N_4716,N_3929,N_3267);
xor U4717 (N_4717,N_3414,N_3309);
xor U4718 (N_4718,N_3400,N_3472);
nor U4719 (N_4719,N_3794,N_3568);
nand U4720 (N_4720,N_3094,N_3009);
and U4721 (N_4721,N_3513,N_3549);
nor U4722 (N_4722,N_3490,N_3789);
nor U4723 (N_4723,N_3616,N_3113);
or U4724 (N_4724,N_3499,N_3674);
or U4725 (N_4725,N_3195,N_3823);
and U4726 (N_4726,N_3602,N_3732);
nor U4727 (N_4727,N_3810,N_3352);
nand U4728 (N_4728,N_3768,N_3567);
xor U4729 (N_4729,N_3242,N_3717);
xnor U4730 (N_4730,N_3100,N_3612);
and U4731 (N_4731,N_3789,N_3683);
xor U4732 (N_4732,N_3645,N_3003);
or U4733 (N_4733,N_3613,N_3436);
xor U4734 (N_4734,N_3717,N_3845);
nor U4735 (N_4735,N_3723,N_3598);
xor U4736 (N_4736,N_3948,N_3665);
and U4737 (N_4737,N_3552,N_3884);
and U4738 (N_4738,N_3503,N_3008);
nand U4739 (N_4739,N_3089,N_3751);
or U4740 (N_4740,N_3177,N_3545);
or U4741 (N_4741,N_3609,N_3073);
xor U4742 (N_4742,N_3908,N_3748);
nor U4743 (N_4743,N_3154,N_3307);
and U4744 (N_4744,N_3896,N_3097);
or U4745 (N_4745,N_3522,N_3724);
or U4746 (N_4746,N_3998,N_3225);
xor U4747 (N_4747,N_3835,N_3019);
xnor U4748 (N_4748,N_3350,N_3961);
nor U4749 (N_4749,N_3379,N_3775);
xor U4750 (N_4750,N_3507,N_3535);
nor U4751 (N_4751,N_3302,N_3189);
nor U4752 (N_4752,N_3941,N_3487);
or U4753 (N_4753,N_3480,N_3463);
xor U4754 (N_4754,N_3865,N_3767);
xor U4755 (N_4755,N_3750,N_3467);
nand U4756 (N_4756,N_3736,N_3215);
xor U4757 (N_4757,N_3461,N_3324);
nor U4758 (N_4758,N_3340,N_3879);
or U4759 (N_4759,N_3365,N_3024);
nand U4760 (N_4760,N_3559,N_3574);
and U4761 (N_4761,N_3711,N_3788);
nor U4762 (N_4762,N_3621,N_3092);
xor U4763 (N_4763,N_3910,N_3984);
nor U4764 (N_4764,N_3439,N_3249);
xor U4765 (N_4765,N_3487,N_3338);
nor U4766 (N_4766,N_3451,N_3333);
nor U4767 (N_4767,N_3854,N_3061);
or U4768 (N_4768,N_3876,N_3160);
nand U4769 (N_4769,N_3174,N_3248);
xnor U4770 (N_4770,N_3438,N_3339);
and U4771 (N_4771,N_3679,N_3323);
nor U4772 (N_4772,N_3630,N_3803);
nand U4773 (N_4773,N_3509,N_3580);
and U4774 (N_4774,N_3971,N_3048);
and U4775 (N_4775,N_3729,N_3610);
nor U4776 (N_4776,N_3708,N_3089);
xor U4777 (N_4777,N_3170,N_3374);
nand U4778 (N_4778,N_3829,N_3992);
nor U4779 (N_4779,N_3235,N_3068);
nand U4780 (N_4780,N_3476,N_3749);
and U4781 (N_4781,N_3339,N_3804);
nor U4782 (N_4782,N_3150,N_3256);
or U4783 (N_4783,N_3186,N_3066);
nor U4784 (N_4784,N_3157,N_3917);
nor U4785 (N_4785,N_3160,N_3444);
and U4786 (N_4786,N_3963,N_3164);
nand U4787 (N_4787,N_3740,N_3379);
and U4788 (N_4788,N_3316,N_3847);
and U4789 (N_4789,N_3435,N_3020);
nor U4790 (N_4790,N_3320,N_3920);
and U4791 (N_4791,N_3183,N_3121);
and U4792 (N_4792,N_3808,N_3052);
and U4793 (N_4793,N_3141,N_3026);
or U4794 (N_4794,N_3140,N_3116);
nor U4795 (N_4795,N_3305,N_3240);
nor U4796 (N_4796,N_3829,N_3959);
and U4797 (N_4797,N_3430,N_3356);
or U4798 (N_4798,N_3999,N_3021);
and U4799 (N_4799,N_3469,N_3251);
and U4800 (N_4800,N_3045,N_3151);
xor U4801 (N_4801,N_3360,N_3264);
and U4802 (N_4802,N_3570,N_3803);
or U4803 (N_4803,N_3809,N_3382);
nand U4804 (N_4804,N_3967,N_3106);
xnor U4805 (N_4805,N_3390,N_3884);
or U4806 (N_4806,N_3475,N_3157);
nor U4807 (N_4807,N_3503,N_3748);
nor U4808 (N_4808,N_3021,N_3071);
nand U4809 (N_4809,N_3201,N_3197);
nor U4810 (N_4810,N_3928,N_3897);
nor U4811 (N_4811,N_3178,N_3791);
xor U4812 (N_4812,N_3834,N_3339);
nand U4813 (N_4813,N_3961,N_3792);
nor U4814 (N_4814,N_3440,N_3384);
and U4815 (N_4815,N_3141,N_3580);
or U4816 (N_4816,N_3622,N_3355);
nor U4817 (N_4817,N_3842,N_3468);
xor U4818 (N_4818,N_3279,N_3977);
nor U4819 (N_4819,N_3198,N_3948);
or U4820 (N_4820,N_3175,N_3965);
or U4821 (N_4821,N_3774,N_3816);
nor U4822 (N_4822,N_3808,N_3815);
xor U4823 (N_4823,N_3120,N_3712);
or U4824 (N_4824,N_3661,N_3411);
and U4825 (N_4825,N_3280,N_3376);
xnor U4826 (N_4826,N_3269,N_3922);
nor U4827 (N_4827,N_3124,N_3518);
nor U4828 (N_4828,N_3548,N_3982);
and U4829 (N_4829,N_3165,N_3579);
or U4830 (N_4830,N_3966,N_3632);
xnor U4831 (N_4831,N_3279,N_3781);
nand U4832 (N_4832,N_3587,N_3729);
nor U4833 (N_4833,N_3983,N_3503);
nor U4834 (N_4834,N_3162,N_3319);
nand U4835 (N_4835,N_3674,N_3062);
nand U4836 (N_4836,N_3995,N_3733);
or U4837 (N_4837,N_3004,N_3643);
nor U4838 (N_4838,N_3824,N_3987);
xnor U4839 (N_4839,N_3822,N_3501);
xor U4840 (N_4840,N_3213,N_3659);
nand U4841 (N_4841,N_3397,N_3899);
nand U4842 (N_4842,N_3309,N_3609);
xnor U4843 (N_4843,N_3364,N_3770);
nand U4844 (N_4844,N_3833,N_3627);
and U4845 (N_4845,N_3135,N_3269);
nor U4846 (N_4846,N_3564,N_3403);
or U4847 (N_4847,N_3878,N_3662);
and U4848 (N_4848,N_3664,N_3112);
nand U4849 (N_4849,N_3083,N_3999);
or U4850 (N_4850,N_3950,N_3252);
or U4851 (N_4851,N_3562,N_3237);
xor U4852 (N_4852,N_3461,N_3541);
nand U4853 (N_4853,N_3913,N_3718);
nand U4854 (N_4854,N_3954,N_3642);
xor U4855 (N_4855,N_3412,N_3892);
xnor U4856 (N_4856,N_3646,N_3746);
nand U4857 (N_4857,N_3216,N_3451);
nor U4858 (N_4858,N_3065,N_3720);
xor U4859 (N_4859,N_3555,N_3125);
xnor U4860 (N_4860,N_3887,N_3515);
nor U4861 (N_4861,N_3033,N_3348);
and U4862 (N_4862,N_3044,N_3668);
or U4863 (N_4863,N_3216,N_3423);
or U4864 (N_4864,N_3172,N_3330);
and U4865 (N_4865,N_3437,N_3983);
or U4866 (N_4866,N_3720,N_3377);
nand U4867 (N_4867,N_3843,N_3571);
xor U4868 (N_4868,N_3414,N_3391);
or U4869 (N_4869,N_3031,N_3878);
nor U4870 (N_4870,N_3637,N_3619);
nand U4871 (N_4871,N_3567,N_3572);
or U4872 (N_4872,N_3859,N_3260);
or U4873 (N_4873,N_3004,N_3530);
xnor U4874 (N_4874,N_3005,N_3399);
nand U4875 (N_4875,N_3196,N_3635);
xnor U4876 (N_4876,N_3175,N_3576);
and U4877 (N_4877,N_3951,N_3554);
nor U4878 (N_4878,N_3701,N_3201);
and U4879 (N_4879,N_3661,N_3454);
xor U4880 (N_4880,N_3002,N_3416);
or U4881 (N_4881,N_3874,N_3764);
nand U4882 (N_4882,N_3367,N_3406);
or U4883 (N_4883,N_3030,N_3667);
and U4884 (N_4884,N_3663,N_3660);
and U4885 (N_4885,N_3869,N_3172);
xnor U4886 (N_4886,N_3748,N_3273);
or U4887 (N_4887,N_3036,N_3427);
xnor U4888 (N_4888,N_3392,N_3126);
nor U4889 (N_4889,N_3966,N_3752);
and U4890 (N_4890,N_3253,N_3951);
or U4891 (N_4891,N_3720,N_3474);
or U4892 (N_4892,N_3057,N_3259);
and U4893 (N_4893,N_3629,N_3579);
nor U4894 (N_4894,N_3978,N_3305);
and U4895 (N_4895,N_3004,N_3473);
and U4896 (N_4896,N_3451,N_3067);
xnor U4897 (N_4897,N_3938,N_3034);
or U4898 (N_4898,N_3330,N_3882);
xnor U4899 (N_4899,N_3205,N_3365);
and U4900 (N_4900,N_3046,N_3911);
nor U4901 (N_4901,N_3704,N_3107);
and U4902 (N_4902,N_3441,N_3429);
and U4903 (N_4903,N_3326,N_3085);
xor U4904 (N_4904,N_3346,N_3361);
nand U4905 (N_4905,N_3815,N_3932);
nor U4906 (N_4906,N_3120,N_3972);
nor U4907 (N_4907,N_3462,N_3345);
or U4908 (N_4908,N_3571,N_3402);
xor U4909 (N_4909,N_3191,N_3980);
or U4910 (N_4910,N_3146,N_3353);
xor U4911 (N_4911,N_3249,N_3950);
xnor U4912 (N_4912,N_3643,N_3591);
or U4913 (N_4913,N_3812,N_3100);
xnor U4914 (N_4914,N_3361,N_3646);
nor U4915 (N_4915,N_3208,N_3824);
or U4916 (N_4916,N_3165,N_3652);
nor U4917 (N_4917,N_3789,N_3086);
nor U4918 (N_4918,N_3481,N_3340);
nand U4919 (N_4919,N_3953,N_3912);
nand U4920 (N_4920,N_3014,N_3819);
or U4921 (N_4921,N_3996,N_3828);
nand U4922 (N_4922,N_3240,N_3129);
or U4923 (N_4923,N_3061,N_3431);
and U4924 (N_4924,N_3356,N_3535);
xor U4925 (N_4925,N_3322,N_3379);
or U4926 (N_4926,N_3106,N_3269);
nand U4927 (N_4927,N_3791,N_3142);
nor U4928 (N_4928,N_3418,N_3492);
or U4929 (N_4929,N_3140,N_3720);
nand U4930 (N_4930,N_3912,N_3737);
and U4931 (N_4931,N_3741,N_3141);
or U4932 (N_4932,N_3159,N_3857);
xnor U4933 (N_4933,N_3858,N_3682);
nand U4934 (N_4934,N_3071,N_3147);
or U4935 (N_4935,N_3221,N_3379);
xnor U4936 (N_4936,N_3966,N_3571);
nor U4937 (N_4937,N_3624,N_3677);
or U4938 (N_4938,N_3870,N_3894);
xor U4939 (N_4939,N_3321,N_3894);
xnor U4940 (N_4940,N_3825,N_3482);
xor U4941 (N_4941,N_3577,N_3282);
nand U4942 (N_4942,N_3144,N_3229);
nor U4943 (N_4943,N_3491,N_3122);
or U4944 (N_4944,N_3560,N_3598);
xnor U4945 (N_4945,N_3694,N_3752);
and U4946 (N_4946,N_3303,N_3033);
nor U4947 (N_4947,N_3029,N_3390);
xnor U4948 (N_4948,N_3017,N_3120);
or U4949 (N_4949,N_3348,N_3879);
nand U4950 (N_4950,N_3890,N_3578);
or U4951 (N_4951,N_3691,N_3582);
or U4952 (N_4952,N_3668,N_3382);
xnor U4953 (N_4953,N_3245,N_3957);
nand U4954 (N_4954,N_3334,N_3287);
or U4955 (N_4955,N_3330,N_3995);
and U4956 (N_4956,N_3699,N_3488);
nand U4957 (N_4957,N_3586,N_3041);
or U4958 (N_4958,N_3380,N_3778);
nand U4959 (N_4959,N_3939,N_3009);
nor U4960 (N_4960,N_3981,N_3601);
nand U4961 (N_4961,N_3062,N_3099);
xnor U4962 (N_4962,N_3456,N_3785);
nor U4963 (N_4963,N_3758,N_3539);
and U4964 (N_4964,N_3485,N_3273);
nor U4965 (N_4965,N_3533,N_3399);
nor U4966 (N_4966,N_3366,N_3298);
and U4967 (N_4967,N_3993,N_3156);
xnor U4968 (N_4968,N_3564,N_3687);
nor U4969 (N_4969,N_3680,N_3973);
nor U4970 (N_4970,N_3338,N_3150);
nor U4971 (N_4971,N_3922,N_3812);
or U4972 (N_4972,N_3618,N_3446);
or U4973 (N_4973,N_3675,N_3902);
nor U4974 (N_4974,N_3726,N_3304);
nand U4975 (N_4975,N_3522,N_3447);
nor U4976 (N_4976,N_3539,N_3978);
xnor U4977 (N_4977,N_3679,N_3417);
or U4978 (N_4978,N_3466,N_3684);
xor U4979 (N_4979,N_3696,N_3059);
or U4980 (N_4980,N_3076,N_3683);
xor U4981 (N_4981,N_3243,N_3098);
xor U4982 (N_4982,N_3421,N_3770);
xor U4983 (N_4983,N_3425,N_3488);
xor U4984 (N_4984,N_3737,N_3153);
nand U4985 (N_4985,N_3992,N_3148);
xor U4986 (N_4986,N_3488,N_3652);
nand U4987 (N_4987,N_3218,N_3273);
nor U4988 (N_4988,N_3360,N_3939);
or U4989 (N_4989,N_3427,N_3059);
nand U4990 (N_4990,N_3534,N_3898);
xor U4991 (N_4991,N_3354,N_3850);
nor U4992 (N_4992,N_3833,N_3045);
nand U4993 (N_4993,N_3807,N_3160);
or U4994 (N_4994,N_3124,N_3367);
nand U4995 (N_4995,N_3307,N_3538);
xor U4996 (N_4996,N_3505,N_3097);
or U4997 (N_4997,N_3996,N_3057);
nand U4998 (N_4998,N_3883,N_3017);
or U4999 (N_4999,N_3249,N_3365);
and U5000 (N_5000,N_4541,N_4346);
or U5001 (N_5001,N_4332,N_4792);
nor U5002 (N_5002,N_4480,N_4246);
xnor U5003 (N_5003,N_4007,N_4723);
nor U5004 (N_5004,N_4789,N_4185);
nor U5005 (N_5005,N_4021,N_4492);
or U5006 (N_5006,N_4065,N_4570);
nand U5007 (N_5007,N_4746,N_4728);
or U5008 (N_5008,N_4549,N_4520);
and U5009 (N_5009,N_4749,N_4691);
nor U5010 (N_5010,N_4055,N_4219);
xor U5011 (N_5011,N_4840,N_4880);
xnor U5012 (N_5012,N_4551,N_4743);
or U5013 (N_5013,N_4407,N_4504);
nor U5014 (N_5014,N_4121,N_4854);
nand U5015 (N_5015,N_4587,N_4049);
or U5016 (N_5016,N_4560,N_4113);
nor U5017 (N_5017,N_4629,N_4242);
or U5018 (N_5018,N_4986,N_4639);
and U5019 (N_5019,N_4171,N_4195);
or U5020 (N_5020,N_4714,N_4952);
xnor U5021 (N_5021,N_4321,N_4444);
nor U5022 (N_5022,N_4883,N_4062);
and U5023 (N_5023,N_4561,N_4735);
nand U5024 (N_5024,N_4773,N_4200);
xor U5025 (N_5025,N_4668,N_4134);
xnor U5026 (N_5026,N_4665,N_4331);
or U5027 (N_5027,N_4759,N_4433);
nor U5028 (N_5028,N_4542,N_4944);
or U5029 (N_5029,N_4973,N_4058);
nor U5030 (N_5030,N_4093,N_4945);
and U5031 (N_5031,N_4566,N_4879);
nor U5032 (N_5032,N_4718,N_4920);
xnor U5033 (N_5033,N_4388,N_4969);
nand U5034 (N_5034,N_4553,N_4226);
nor U5035 (N_5035,N_4696,N_4163);
and U5036 (N_5036,N_4605,N_4913);
or U5037 (N_5037,N_4027,N_4387);
xnor U5038 (N_5038,N_4032,N_4656);
xor U5039 (N_5039,N_4820,N_4647);
and U5040 (N_5040,N_4715,N_4698);
or U5041 (N_5041,N_4413,N_4596);
nor U5042 (N_5042,N_4369,N_4104);
xor U5043 (N_5043,N_4653,N_4812);
nand U5044 (N_5044,N_4244,N_4807);
xor U5045 (N_5045,N_4706,N_4237);
and U5046 (N_5046,N_4804,N_4288);
nor U5047 (N_5047,N_4175,N_4394);
xor U5048 (N_5048,N_4004,N_4261);
nor U5049 (N_5049,N_4344,N_4724);
and U5050 (N_5050,N_4236,N_4708);
or U5051 (N_5051,N_4164,N_4046);
xnor U5052 (N_5052,N_4671,N_4029);
or U5053 (N_5053,N_4834,N_4657);
nand U5054 (N_5054,N_4469,N_4811);
or U5055 (N_5055,N_4584,N_4833);
nand U5056 (N_5056,N_4962,N_4005);
or U5057 (N_5057,N_4417,N_4866);
or U5058 (N_5058,N_4679,N_4930);
or U5059 (N_5059,N_4926,N_4109);
nand U5060 (N_5060,N_4410,N_4270);
xor U5061 (N_5061,N_4375,N_4563);
xnor U5062 (N_5062,N_4318,N_4893);
xnor U5063 (N_5063,N_4736,N_4465);
xor U5064 (N_5064,N_4090,N_4450);
or U5065 (N_5065,N_4608,N_4153);
nor U5066 (N_5066,N_4509,N_4474);
or U5067 (N_5067,N_4212,N_4742);
and U5068 (N_5068,N_4946,N_4786);
nand U5069 (N_5069,N_4774,N_4564);
nand U5070 (N_5070,N_4468,N_4501);
and U5071 (N_5071,N_4592,N_4285);
and U5072 (N_5072,N_4430,N_4690);
nor U5073 (N_5073,N_4333,N_4071);
or U5074 (N_5074,N_4953,N_4950);
and U5075 (N_5075,N_4799,N_4516);
xnor U5076 (N_5076,N_4737,N_4421);
or U5077 (N_5077,N_4456,N_4087);
and U5078 (N_5078,N_4284,N_4081);
nand U5079 (N_5079,N_4280,N_4967);
and U5080 (N_5080,N_4012,N_4511);
nor U5081 (N_5081,N_4684,N_4047);
xnor U5082 (N_5082,N_4882,N_4255);
nand U5083 (N_5083,N_4623,N_4573);
or U5084 (N_5084,N_4576,N_4241);
xor U5085 (N_5085,N_4901,N_4364);
or U5086 (N_5086,N_4199,N_4341);
nor U5087 (N_5087,N_4156,N_4905);
nand U5088 (N_5088,N_4102,N_4061);
and U5089 (N_5089,N_4727,N_4157);
nor U5090 (N_5090,N_4627,N_4338);
or U5091 (N_5091,N_4726,N_4381);
or U5092 (N_5092,N_4748,N_4326);
nor U5093 (N_5093,N_4253,N_4921);
and U5094 (N_5094,N_4386,N_4779);
xnor U5095 (N_5095,N_4734,N_4303);
xor U5096 (N_5096,N_4568,N_4855);
nand U5097 (N_5097,N_4074,N_4125);
nand U5098 (N_5098,N_4458,N_4149);
and U5099 (N_5099,N_4194,N_4756);
or U5100 (N_5100,N_4556,N_4207);
or U5101 (N_5101,N_4397,N_4764);
nor U5102 (N_5102,N_4814,N_4939);
and U5103 (N_5103,N_4546,N_4116);
or U5104 (N_5104,N_4853,N_4794);
nand U5105 (N_5105,N_4009,N_4354);
nor U5106 (N_5106,N_4739,N_4152);
or U5107 (N_5107,N_4427,N_4536);
or U5108 (N_5108,N_4716,N_4825);
nor U5109 (N_5109,N_4750,N_4871);
nand U5110 (N_5110,N_4110,N_4223);
and U5111 (N_5111,N_4637,N_4440);
and U5112 (N_5112,N_4725,N_4403);
xnor U5113 (N_5113,N_4972,N_4186);
nor U5114 (N_5114,N_4365,N_4589);
xor U5115 (N_5115,N_4126,N_4131);
or U5116 (N_5116,N_4574,N_4521);
xor U5117 (N_5117,N_4028,N_4069);
nand U5118 (N_5118,N_4819,N_4582);
or U5119 (N_5119,N_4254,N_4655);
or U5120 (N_5120,N_4291,N_4707);
and U5121 (N_5121,N_4642,N_4632);
nand U5122 (N_5122,N_4203,N_4654);
xnor U5123 (N_5123,N_4890,N_4167);
xor U5124 (N_5124,N_4687,N_4868);
nand U5125 (N_5125,N_4362,N_4772);
nor U5126 (N_5126,N_4620,N_4686);
nor U5127 (N_5127,N_4290,N_4377);
nand U5128 (N_5128,N_4558,N_4624);
or U5129 (N_5129,N_4385,N_4765);
xnor U5130 (N_5130,N_4697,N_4399);
xnor U5131 (N_5131,N_4429,N_4795);
and U5132 (N_5132,N_4809,N_4777);
nand U5133 (N_5133,N_4320,N_4705);
nor U5134 (N_5134,N_4722,N_4958);
nor U5135 (N_5135,N_4192,N_4517);
and U5136 (N_5136,N_4328,N_4769);
nand U5137 (N_5137,N_4154,N_4785);
nor U5138 (N_5138,N_4720,N_4494);
and U5139 (N_5139,N_4190,N_4122);
nor U5140 (N_5140,N_4416,N_4128);
xnor U5141 (N_5141,N_4678,N_4273);
and U5142 (N_5142,N_4788,N_4783);
nor U5143 (N_5143,N_4670,N_4857);
nor U5144 (N_5144,N_4887,N_4111);
or U5145 (N_5145,N_4514,N_4776);
nand U5146 (N_5146,N_4052,N_4595);
nand U5147 (N_5147,N_4196,N_4076);
or U5148 (N_5148,N_4601,N_4079);
nor U5149 (N_5149,N_4626,N_4873);
or U5150 (N_5150,N_4144,N_4051);
xor U5151 (N_5151,N_4949,N_4233);
xnor U5152 (N_5152,N_4538,N_4393);
xor U5153 (N_5153,N_4250,N_4170);
and U5154 (N_5154,N_4851,N_4348);
nand U5155 (N_5155,N_4446,N_4982);
or U5156 (N_5156,N_4150,N_4597);
or U5157 (N_5157,N_4912,N_4650);
and U5158 (N_5158,N_4680,N_4903);
nor U5159 (N_5159,N_4137,N_4455);
nand U5160 (N_5160,N_4611,N_4409);
nand U5161 (N_5161,N_4941,N_4984);
and U5162 (N_5162,N_4208,N_4402);
and U5163 (N_5163,N_4347,N_4666);
xnor U5164 (N_5164,N_4197,N_4523);
or U5165 (N_5165,N_4907,N_4165);
or U5166 (N_5166,N_4518,N_4638);
and U5167 (N_5167,N_4428,N_4527);
and U5168 (N_5168,N_4847,N_4389);
and U5169 (N_5169,N_4002,N_4470);
xnor U5170 (N_5170,N_4900,N_4540);
xnor U5171 (N_5171,N_4987,N_4881);
nand U5172 (N_5172,N_4761,N_4897);
and U5173 (N_5173,N_4496,N_4436);
and U5174 (N_5174,N_4443,N_4633);
nand U5175 (N_5175,N_4800,N_4619);
nor U5176 (N_5176,N_4020,N_4826);
nor U5177 (N_5177,N_4554,N_4581);
nand U5178 (N_5178,N_4374,N_4781);
nor U5179 (N_5179,N_4198,N_4618);
or U5180 (N_5180,N_4204,N_4395);
and U5181 (N_5181,N_4844,N_4983);
or U5182 (N_5182,N_4439,N_4505);
nor U5183 (N_5183,N_4583,N_4302);
and U5184 (N_5184,N_4422,N_4050);
nor U5185 (N_5185,N_4221,N_4401);
and U5186 (N_5186,N_4092,N_4934);
and U5187 (N_5187,N_4106,N_4559);
nor U5188 (N_5188,N_4989,N_4497);
or U5189 (N_5189,N_4992,N_4041);
and U5190 (N_5190,N_4675,N_4392);
nor U5191 (N_5191,N_4733,N_4938);
nand U5192 (N_5192,N_4179,N_4418);
and U5193 (N_5193,N_4565,N_4771);
and U5194 (N_5194,N_4995,N_4117);
nand U5195 (N_5195,N_4214,N_4297);
and U5196 (N_5196,N_4658,N_4831);
nand U5197 (N_5197,N_4869,N_4937);
xor U5198 (N_5198,N_4043,N_4317);
xor U5199 (N_5199,N_4606,N_4307);
nand U5200 (N_5200,N_4711,N_4817);
or U5201 (N_5201,N_4053,N_4437);
xnor U5202 (N_5202,N_4598,N_4645);
nor U5203 (N_5203,N_4649,N_4139);
xnor U5204 (N_5204,N_4299,N_4420);
nor U5205 (N_5205,N_4202,N_4822);
and U5206 (N_5206,N_4024,N_4008);
xor U5207 (N_5207,N_4217,N_4447);
nor U5208 (N_5208,N_4095,N_4425);
nor U5209 (N_5209,N_4547,N_4238);
or U5210 (N_5210,N_4755,N_4482);
and U5211 (N_5211,N_4042,N_4211);
xnor U5212 (N_5212,N_4940,N_4909);
or U5213 (N_5213,N_4463,N_4486);
and U5214 (N_5214,N_4507,N_4575);
nand U5215 (N_5215,N_4925,N_4350);
nand U5216 (N_5216,N_4183,N_4979);
nand U5217 (N_5217,N_4088,N_4974);
or U5218 (N_5218,N_4823,N_4719);
nand U5219 (N_5219,N_4569,N_4448);
nor U5220 (N_5220,N_4222,N_4703);
nand U5221 (N_5221,N_4562,N_4506);
and U5222 (N_5222,N_4683,N_4232);
xor U5223 (N_5223,N_4841,N_4457);
xnor U5224 (N_5224,N_4904,N_4075);
or U5225 (N_5225,N_4567,N_4461);
or U5226 (N_5226,N_4166,N_4271);
nand U5227 (N_5227,N_4345,N_4685);
or U5228 (N_5228,N_4481,N_4681);
xor U5229 (N_5229,N_4266,N_4304);
and U5230 (N_5230,N_4181,N_4013);
xnor U5231 (N_5231,N_4096,N_4682);
or U5232 (N_5232,N_4867,N_4923);
xor U5233 (N_5233,N_4651,N_4862);
xnor U5234 (N_5234,N_4070,N_4089);
xor U5235 (N_5235,N_4329,N_4612);
nor U5236 (N_5236,N_4966,N_4355);
and U5237 (N_5237,N_4366,N_4129);
nor U5238 (N_5238,N_4182,N_4955);
nor U5239 (N_5239,N_4502,N_4778);
nand U5240 (N_5240,N_4745,N_4688);
xor U5241 (N_5241,N_4265,N_4015);
and U5242 (N_5242,N_4339,N_4766);
nor U5243 (N_5243,N_4085,N_4352);
nand U5244 (N_5244,N_4602,N_4180);
nand U5245 (N_5245,N_4054,N_4373);
and U5246 (N_5246,N_4997,N_4340);
xor U5247 (N_5247,N_4752,N_4634);
nand U5248 (N_5248,N_4702,N_4114);
nor U5249 (N_5249,N_4815,N_4856);
nand U5250 (N_5250,N_4802,N_4895);
or U5251 (N_5251,N_4249,N_4943);
nor U5252 (N_5252,N_4648,N_4312);
or U5253 (N_5253,N_4325,N_4248);
nor U5254 (N_5254,N_4545,N_4442);
and U5255 (N_5255,N_4022,N_4292);
nand U5256 (N_5256,N_4915,N_4206);
or U5257 (N_5257,N_4740,N_4193);
xnor U5258 (N_5258,N_4676,N_4239);
and U5259 (N_5259,N_4874,N_4935);
and U5260 (N_5260,N_4790,N_4390);
nor U5261 (N_5261,N_4594,N_4404);
and U5262 (N_5262,N_4172,N_4641);
nand U5263 (N_5263,N_4296,N_4431);
or U5264 (N_5264,N_4229,N_4808);
and U5265 (N_5265,N_4479,N_4908);
or U5266 (N_5266,N_4363,N_4342);
nand U5267 (N_5267,N_4978,N_4080);
nor U5268 (N_5268,N_4701,N_4892);
xor U5269 (N_5269,N_4435,N_4911);
and U5270 (N_5270,N_4030,N_4294);
xor U5271 (N_5271,N_4976,N_4591);
nand U5272 (N_5272,N_4098,N_4490);
and U5273 (N_5273,N_4311,N_4228);
or U5274 (N_5274,N_4484,N_4309);
nand U5275 (N_5275,N_4033,N_4493);
nand U5276 (N_5276,N_4510,N_4784);
and U5277 (N_5277,N_4003,N_4801);
xor U5278 (N_5278,N_4625,N_4636);
nor U5279 (N_5279,N_4942,N_4278);
and U5280 (N_5280,N_4732,N_4586);
and U5281 (N_5281,N_4452,N_4010);
or U5282 (N_5282,N_4617,N_4132);
nand U5283 (N_5283,N_4933,N_4295);
nand U5284 (N_5284,N_4975,N_4860);
nand U5285 (N_5285,N_4947,N_4391);
nand U5286 (N_5286,N_4017,N_4048);
nand U5287 (N_5287,N_4337,N_4824);
and U5288 (N_5288,N_4123,N_4260);
nor U5289 (N_5289,N_4286,N_4130);
xor U5290 (N_5290,N_4793,N_4533);
xor U5291 (N_5291,N_4018,N_4693);
nor U5292 (N_5292,N_4405,N_4251);
nand U5293 (N_5293,N_4888,N_4960);
and U5294 (N_5294,N_4672,N_4257);
or U5295 (N_5295,N_4082,N_4169);
nor U5296 (N_5296,N_4334,N_4539);
and U5297 (N_5297,N_4865,N_4552);
and U5298 (N_5298,N_4159,N_4689);
and U5299 (N_5299,N_4530,N_4717);
nor U5300 (N_5300,N_4961,N_4991);
and U5301 (N_5301,N_4613,N_4610);
and U5302 (N_5302,N_4981,N_4245);
and U5303 (N_5303,N_4848,N_4664);
xor U5304 (N_5304,N_4891,N_4314);
nor U5305 (N_5305,N_4875,N_4850);
or U5306 (N_5306,N_4603,N_4100);
and U5307 (N_5307,N_4931,N_4039);
xor U5308 (N_5308,N_4408,N_4068);
and U5309 (N_5309,N_4262,N_4529);
xor U5310 (N_5310,N_4803,N_4160);
xor U5311 (N_5311,N_4158,N_4000);
or U5312 (N_5312,N_4301,N_4579);
or U5313 (N_5313,N_4877,N_4741);
or U5314 (N_5314,N_4839,N_4599);
xor U5315 (N_5315,N_4016,N_4957);
nand U5316 (N_5316,N_4336,N_4322);
or U5317 (N_5317,N_4057,N_4234);
nand U5318 (N_5318,N_4896,N_4449);
xor U5319 (N_5319,N_4188,N_4578);
and U5320 (N_5320,N_4604,N_4327);
nand U5321 (N_5321,N_4209,N_4063);
and U5322 (N_5322,N_4064,N_4673);
or U5323 (N_5323,N_4730,N_4240);
nor U5324 (N_5324,N_4956,N_4376);
xor U5325 (N_5325,N_4555,N_4298);
and U5326 (N_5326,N_4744,N_4335);
nand U5327 (N_5327,N_4146,N_4951);
or U5328 (N_5328,N_4256,N_4147);
or U5329 (N_5329,N_4990,N_4994);
and U5330 (N_5330,N_4964,N_4380);
xnor U5331 (N_5331,N_4475,N_4872);
nand U5332 (N_5332,N_4532,N_4631);
xor U5333 (N_5333,N_4281,N_4434);
nor U5334 (N_5334,N_4215,N_4924);
xor U5335 (N_5335,N_4646,N_4709);
or U5336 (N_5336,N_4036,N_4138);
or U5337 (N_5337,N_4396,N_4534);
xor U5338 (N_5338,N_4806,N_4699);
xnor U5339 (N_5339,N_4531,N_4550);
or U5340 (N_5340,N_4644,N_4615);
and U5341 (N_5341,N_4487,N_4999);
or U5342 (N_5342,N_4537,N_4899);
or U5343 (N_5343,N_4916,N_4073);
xor U5344 (N_5344,N_4423,N_4889);
nand U5345 (N_5345,N_4289,N_4600);
and U5346 (N_5346,N_4025,N_4863);
nand U5347 (N_5347,N_4067,N_4379);
nand U5348 (N_5348,N_4034,N_4971);
nand U5349 (N_5349,N_4384,N_4970);
xnor U5350 (N_5350,N_4635,N_4220);
or U5351 (N_5351,N_4370,N_4174);
or U5352 (N_5352,N_4023,N_4513);
nand U5353 (N_5353,N_4323,N_4258);
nand U5354 (N_5354,N_4628,N_4072);
xor U5355 (N_5355,N_4998,N_4928);
xnor U5356 (N_5356,N_4412,N_4464);
nor U5357 (N_5357,N_4133,N_4500);
nor U5358 (N_5358,N_4512,N_4524);
and U5359 (N_5359,N_4544,N_4607);
xnor U5360 (N_5360,N_4279,N_4127);
nand U5361 (N_5361,N_4115,N_4993);
xor U5362 (N_5362,N_4276,N_4996);
xor U5363 (N_5363,N_4099,N_4343);
and U5364 (N_5364,N_4667,N_4832);
and U5365 (N_5365,N_4227,N_4168);
and U5366 (N_5366,N_4622,N_4731);
xor U5367 (N_5367,N_4078,N_4108);
and U5368 (N_5368,N_4191,N_4571);
and U5369 (N_5369,N_4210,N_4593);
and U5370 (N_5370,N_4488,N_4515);
nand U5371 (N_5371,N_4796,N_4218);
or U5372 (N_5372,N_4243,N_4148);
and U5373 (N_5373,N_4526,N_4415);
nor U5374 (N_5374,N_4398,N_4356);
xnor U5375 (N_5375,N_4224,N_4780);
nor U5376 (N_5376,N_4489,N_4189);
nand U5377 (N_5377,N_4438,N_4040);
nand U5378 (N_5378,N_4838,N_4810);
nand U5379 (N_5379,N_4936,N_4274);
nor U5380 (N_5380,N_4758,N_4713);
nand U5381 (N_5381,N_4313,N_4472);
and U5382 (N_5382,N_4151,N_4315);
and U5383 (N_5383,N_4830,N_4060);
nand U5384 (N_5384,N_4609,N_4821);
or U5385 (N_5385,N_4621,N_4798);
and U5386 (N_5386,N_4886,N_4852);
nand U5387 (N_5387,N_4259,N_4454);
and U5388 (N_5388,N_4585,N_4173);
and U5389 (N_5389,N_4885,N_4827);
and U5390 (N_5390,N_4287,N_4580);
nor U5391 (N_5391,N_4837,N_4922);
or U5392 (N_5392,N_4519,N_4704);
xor U5393 (N_5393,N_4495,N_4176);
or U5394 (N_5394,N_4006,N_4498);
xnor U5395 (N_5395,N_4894,N_4859);
or U5396 (N_5396,N_4721,N_4101);
or U5397 (N_5397,N_4383,N_4358);
nand U5398 (N_5398,N_4216,N_4828);
nand U5399 (N_5399,N_4753,N_4674);
nor U5400 (N_5400,N_4272,N_4948);
nor U5401 (N_5401,N_4652,N_4963);
or U5402 (N_5402,N_4441,N_4588);
and U5403 (N_5403,N_4614,N_4044);
and U5404 (N_5404,N_4959,N_4184);
nor U5405 (N_5405,N_4965,N_4548);
xor U5406 (N_5406,N_4406,N_4927);
xor U5407 (N_5407,N_4453,N_4980);
or U5408 (N_5408,N_4084,N_4932);
xor U5409 (N_5409,N_4919,N_4143);
and U5410 (N_5410,N_4359,N_4662);
and U5411 (N_5411,N_4118,N_4277);
or U5412 (N_5412,N_4577,N_4902);
and U5413 (N_5413,N_4797,N_4103);
nor U5414 (N_5414,N_4135,N_4112);
or U5415 (N_5415,N_4091,N_4787);
nand U5416 (N_5416,N_4107,N_4451);
nand U5417 (N_5417,N_4066,N_4861);
nor U5418 (N_5418,N_4884,N_4059);
and U5419 (N_5419,N_4768,N_4424);
nor U5420 (N_5420,N_4119,N_4471);
and U5421 (N_5421,N_4710,N_4762);
nand U5422 (N_5422,N_4459,N_4400);
or U5423 (N_5423,N_4268,N_4590);
xnor U5424 (N_5424,N_4700,N_4011);
nor U5425 (N_5425,N_4001,N_4269);
nor U5426 (N_5426,N_4086,N_4105);
xor U5427 (N_5427,N_4306,N_4864);
or U5428 (N_5428,N_4525,N_4813);
nand U5429 (N_5429,N_4283,N_4426);
and U5430 (N_5430,N_4231,N_4445);
nand U5431 (N_5431,N_4842,N_4432);
or U5432 (N_5432,N_4077,N_4661);
or U5433 (N_5433,N_4843,N_4988);
and U5434 (N_5434,N_4818,N_4142);
nand U5435 (N_5435,N_4572,N_4985);
nand U5436 (N_5436,N_4914,N_4316);
xnor U5437 (N_5437,N_4910,N_4378);
or U5438 (N_5438,N_4754,N_4460);
nor U5439 (N_5439,N_4829,N_4045);
xnor U5440 (N_5440,N_4037,N_4213);
nor U5441 (N_5441,N_4097,N_4712);
and U5442 (N_5442,N_4161,N_4177);
xnor U5443 (N_5443,N_4264,N_4929);
xor U5444 (N_5444,N_4324,N_4977);
and U5445 (N_5445,N_4491,N_4031);
or U5446 (N_5446,N_4019,N_4476);
or U5447 (N_5447,N_4477,N_4124);
nand U5448 (N_5448,N_4918,N_4499);
nand U5449 (N_5449,N_4630,N_4791);
nand U5450 (N_5450,N_4738,N_4187);
nand U5451 (N_5451,N_4467,N_4305);
or U5452 (N_5452,N_4205,N_4247);
and U5453 (N_5453,N_4816,N_4162);
or U5454 (N_5454,N_4663,N_4845);
or U5455 (N_5455,N_4310,N_4751);
nor U5456 (N_5456,N_4267,N_4263);
nor U5457 (N_5457,N_4178,N_4643);
nor U5458 (N_5458,N_4528,N_4419);
nand U5459 (N_5459,N_4835,N_4659);
and U5460 (N_5460,N_4917,N_4140);
nand U5461 (N_5461,N_4669,N_4145);
or U5462 (N_5462,N_4535,N_4483);
or U5463 (N_5463,N_4371,N_4775);
or U5464 (N_5464,N_4382,N_4293);
nor U5465 (N_5465,N_4485,N_4543);
or U5466 (N_5466,N_4201,N_4729);
nor U5467 (N_5467,N_4141,N_4660);
xnor U5468 (N_5468,N_4906,N_4330);
or U5469 (N_5469,N_4308,N_4035);
and U5470 (N_5470,N_4275,N_4026);
and U5471 (N_5471,N_4677,N_4694);
or U5472 (N_5472,N_4747,N_4640);
nor U5473 (N_5473,N_4763,N_4155);
nand U5474 (N_5474,N_4014,N_4770);
nand U5475 (N_5475,N_4805,N_4235);
nor U5476 (N_5476,N_4695,N_4083);
xor U5477 (N_5477,N_4557,N_4056);
xor U5478 (N_5478,N_4954,N_4367);
and U5479 (N_5479,N_4968,N_4760);
xor U5480 (N_5480,N_4411,N_4870);
nand U5481 (N_5481,N_4616,N_4319);
nor U5482 (N_5482,N_4349,N_4522);
nand U5483 (N_5483,N_4478,N_4282);
nor U5484 (N_5484,N_4757,N_4878);
xnor U5485 (N_5485,N_4136,N_4692);
nand U5486 (N_5486,N_4368,N_4252);
xnor U5487 (N_5487,N_4782,N_4225);
xor U5488 (N_5488,N_4503,N_4473);
nand U5489 (N_5489,N_4353,N_4230);
xnor U5490 (N_5490,N_4120,N_4361);
or U5491 (N_5491,N_4898,N_4300);
or U5492 (N_5492,N_4767,N_4462);
and U5493 (N_5493,N_4360,N_4858);
nor U5494 (N_5494,N_4836,N_4846);
or U5495 (N_5495,N_4466,N_4508);
and U5496 (N_5496,N_4094,N_4351);
nand U5497 (N_5497,N_4038,N_4414);
xnor U5498 (N_5498,N_4849,N_4357);
and U5499 (N_5499,N_4372,N_4876);
xor U5500 (N_5500,N_4540,N_4447);
nor U5501 (N_5501,N_4689,N_4422);
and U5502 (N_5502,N_4844,N_4177);
and U5503 (N_5503,N_4132,N_4711);
nand U5504 (N_5504,N_4512,N_4730);
and U5505 (N_5505,N_4881,N_4976);
nand U5506 (N_5506,N_4352,N_4312);
nor U5507 (N_5507,N_4134,N_4674);
xnor U5508 (N_5508,N_4984,N_4995);
nor U5509 (N_5509,N_4939,N_4557);
and U5510 (N_5510,N_4256,N_4874);
xnor U5511 (N_5511,N_4870,N_4161);
xor U5512 (N_5512,N_4607,N_4236);
xnor U5513 (N_5513,N_4858,N_4920);
xor U5514 (N_5514,N_4272,N_4882);
or U5515 (N_5515,N_4667,N_4981);
nand U5516 (N_5516,N_4042,N_4056);
and U5517 (N_5517,N_4007,N_4150);
xor U5518 (N_5518,N_4269,N_4763);
xor U5519 (N_5519,N_4413,N_4661);
or U5520 (N_5520,N_4325,N_4145);
xor U5521 (N_5521,N_4189,N_4785);
or U5522 (N_5522,N_4370,N_4583);
nand U5523 (N_5523,N_4284,N_4059);
nand U5524 (N_5524,N_4304,N_4888);
nor U5525 (N_5525,N_4941,N_4665);
nor U5526 (N_5526,N_4553,N_4264);
or U5527 (N_5527,N_4281,N_4323);
xnor U5528 (N_5528,N_4928,N_4372);
xor U5529 (N_5529,N_4699,N_4013);
xnor U5530 (N_5530,N_4114,N_4467);
nand U5531 (N_5531,N_4873,N_4354);
nor U5532 (N_5532,N_4057,N_4253);
and U5533 (N_5533,N_4215,N_4954);
nor U5534 (N_5534,N_4752,N_4222);
and U5535 (N_5535,N_4167,N_4432);
and U5536 (N_5536,N_4790,N_4505);
or U5537 (N_5537,N_4278,N_4692);
nor U5538 (N_5538,N_4495,N_4480);
nor U5539 (N_5539,N_4271,N_4451);
nor U5540 (N_5540,N_4375,N_4223);
or U5541 (N_5541,N_4787,N_4384);
and U5542 (N_5542,N_4709,N_4868);
and U5543 (N_5543,N_4889,N_4546);
nor U5544 (N_5544,N_4794,N_4724);
nor U5545 (N_5545,N_4148,N_4806);
and U5546 (N_5546,N_4070,N_4551);
nand U5547 (N_5547,N_4346,N_4263);
nand U5548 (N_5548,N_4353,N_4300);
nand U5549 (N_5549,N_4970,N_4701);
xnor U5550 (N_5550,N_4713,N_4050);
nand U5551 (N_5551,N_4575,N_4726);
xor U5552 (N_5552,N_4409,N_4313);
or U5553 (N_5553,N_4677,N_4409);
xor U5554 (N_5554,N_4074,N_4204);
or U5555 (N_5555,N_4768,N_4966);
and U5556 (N_5556,N_4258,N_4961);
or U5557 (N_5557,N_4155,N_4393);
nand U5558 (N_5558,N_4803,N_4830);
nor U5559 (N_5559,N_4645,N_4980);
xor U5560 (N_5560,N_4338,N_4622);
nand U5561 (N_5561,N_4756,N_4471);
xor U5562 (N_5562,N_4846,N_4300);
nor U5563 (N_5563,N_4394,N_4347);
nand U5564 (N_5564,N_4618,N_4659);
nor U5565 (N_5565,N_4214,N_4334);
or U5566 (N_5566,N_4859,N_4054);
and U5567 (N_5567,N_4837,N_4868);
nand U5568 (N_5568,N_4973,N_4006);
nand U5569 (N_5569,N_4031,N_4954);
xnor U5570 (N_5570,N_4034,N_4074);
nand U5571 (N_5571,N_4941,N_4091);
nand U5572 (N_5572,N_4690,N_4050);
xor U5573 (N_5573,N_4859,N_4541);
or U5574 (N_5574,N_4197,N_4266);
xor U5575 (N_5575,N_4899,N_4119);
nand U5576 (N_5576,N_4448,N_4637);
and U5577 (N_5577,N_4933,N_4262);
xnor U5578 (N_5578,N_4541,N_4493);
nand U5579 (N_5579,N_4779,N_4027);
xnor U5580 (N_5580,N_4824,N_4200);
nand U5581 (N_5581,N_4847,N_4123);
nand U5582 (N_5582,N_4175,N_4837);
xnor U5583 (N_5583,N_4500,N_4269);
or U5584 (N_5584,N_4614,N_4906);
or U5585 (N_5585,N_4931,N_4426);
xor U5586 (N_5586,N_4390,N_4580);
or U5587 (N_5587,N_4944,N_4864);
xnor U5588 (N_5588,N_4439,N_4522);
nor U5589 (N_5589,N_4383,N_4043);
xor U5590 (N_5590,N_4907,N_4412);
and U5591 (N_5591,N_4617,N_4526);
nand U5592 (N_5592,N_4174,N_4696);
nand U5593 (N_5593,N_4710,N_4186);
nand U5594 (N_5594,N_4572,N_4839);
and U5595 (N_5595,N_4219,N_4210);
nand U5596 (N_5596,N_4574,N_4212);
nand U5597 (N_5597,N_4427,N_4050);
or U5598 (N_5598,N_4694,N_4936);
xnor U5599 (N_5599,N_4533,N_4107);
and U5600 (N_5600,N_4849,N_4158);
xnor U5601 (N_5601,N_4622,N_4118);
and U5602 (N_5602,N_4269,N_4143);
xor U5603 (N_5603,N_4748,N_4096);
xnor U5604 (N_5604,N_4784,N_4828);
and U5605 (N_5605,N_4065,N_4524);
nor U5606 (N_5606,N_4968,N_4560);
and U5607 (N_5607,N_4426,N_4621);
nand U5608 (N_5608,N_4353,N_4960);
and U5609 (N_5609,N_4772,N_4064);
and U5610 (N_5610,N_4322,N_4107);
xor U5611 (N_5611,N_4411,N_4568);
nand U5612 (N_5612,N_4792,N_4489);
or U5613 (N_5613,N_4046,N_4763);
or U5614 (N_5614,N_4725,N_4374);
nand U5615 (N_5615,N_4092,N_4752);
nand U5616 (N_5616,N_4347,N_4075);
xnor U5617 (N_5617,N_4496,N_4256);
xor U5618 (N_5618,N_4702,N_4953);
and U5619 (N_5619,N_4961,N_4333);
and U5620 (N_5620,N_4004,N_4793);
or U5621 (N_5621,N_4625,N_4686);
nor U5622 (N_5622,N_4596,N_4313);
nor U5623 (N_5623,N_4025,N_4028);
nor U5624 (N_5624,N_4351,N_4461);
or U5625 (N_5625,N_4137,N_4086);
nand U5626 (N_5626,N_4285,N_4902);
xnor U5627 (N_5627,N_4279,N_4635);
nor U5628 (N_5628,N_4266,N_4722);
nand U5629 (N_5629,N_4653,N_4430);
nor U5630 (N_5630,N_4348,N_4068);
and U5631 (N_5631,N_4038,N_4941);
and U5632 (N_5632,N_4906,N_4470);
nor U5633 (N_5633,N_4285,N_4539);
nand U5634 (N_5634,N_4064,N_4227);
and U5635 (N_5635,N_4142,N_4112);
and U5636 (N_5636,N_4898,N_4670);
nor U5637 (N_5637,N_4285,N_4074);
xor U5638 (N_5638,N_4406,N_4167);
nand U5639 (N_5639,N_4141,N_4559);
nand U5640 (N_5640,N_4431,N_4085);
nor U5641 (N_5641,N_4991,N_4739);
nor U5642 (N_5642,N_4265,N_4825);
or U5643 (N_5643,N_4244,N_4567);
nand U5644 (N_5644,N_4854,N_4867);
or U5645 (N_5645,N_4213,N_4822);
and U5646 (N_5646,N_4755,N_4309);
or U5647 (N_5647,N_4138,N_4703);
and U5648 (N_5648,N_4312,N_4150);
xnor U5649 (N_5649,N_4284,N_4373);
xnor U5650 (N_5650,N_4356,N_4592);
or U5651 (N_5651,N_4956,N_4580);
or U5652 (N_5652,N_4626,N_4441);
and U5653 (N_5653,N_4228,N_4060);
nand U5654 (N_5654,N_4220,N_4412);
or U5655 (N_5655,N_4595,N_4434);
xnor U5656 (N_5656,N_4666,N_4240);
nor U5657 (N_5657,N_4332,N_4925);
nand U5658 (N_5658,N_4831,N_4929);
and U5659 (N_5659,N_4843,N_4048);
nand U5660 (N_5660,N_4489,N_4533);
nand U5661 (N_5661,N_4648,N_4148);
nor U5662 (N_5662,N_4827,N_4025);
nand U5663 (N_5663,N_4031,N_4178);
nor U5664 (N_5664,N_4636,N_4495);
nor U5665 (N_5665,N_4177,N_4799);
xor U5666 (N_5666,N_4633,N_4501);
or U5667 (N_5667,N_4424,N_4337);
or U5668 (N_5668,N_4233,N_4083);
and U5669 (N_5669,N_4962,N_4683);
and U5670 (N_5670,N_4046,N_4159);
and U5671 (N_5671,N_4095,N_4490);
or U5672 (N_5672,N_4553,N_4268);
and U5673 (N_5673,N_4170,N_4619);
nand U5674 (N_5674,N_4719,N_4417);
nor U5675 (N_5675,N_4369,N_4850);
nand U5676 (N_5676,N_4357,N_4455);
nand U5677 (N_5677,N_4655,N_4991);
nor U5678 (N_5678,N_4089,N_4602);
nor U5679 (N_5679,N_4332,N_4718);
or U5680 (N_5680,N_4087,N_4789);
xor U5681 (N_5681,N_4117,N_4036);
nand U5682 (N_5682,N_4846,N_4181);
or U5683 (N_5683,N_4027,N_4262);
nor U5684 (N_5684,N_4274,N_4875);
nor U5685 (N_5685,N_4421,N_4007);
and U5686 (N_5686,N_4255,N_4251);
nor U5687 (N_5687,N_4553,N_4677);
and U5688 (N_5688,N_4123,N_4587);
or U5689 (N_5689,N_4269,N_4429);
nor U5690 (N_5690,N_4550,N_4591);
xor U5691 (N_5691,N_4243,N_4956);
xor U5692 (N_5692,N_4407,N_4322);
or U5693 (N_5693,N_4211,N_4560);
nand U5694 (N_5694,N_4616,N_4205);
nand U5695 (N_5695,N_4034,N_4022);
nor U5696 (N_5696,N_4764,N_4235);
nor U5697 (N_5697,N_4779,N_4418);
or U5698 (N_5698,N_4496,N_4943);
and U5699 (N_5699,N_4360,N_4665);
nor U5700 (N_5700,N_4867,N_4978);
and U5701 (N_5701,N_4136,N_4126);
or U5702 (N_5702,N_4156,N_4825);
nor U5703 (N_5703,N_4387,N_4592);
nand U5704 (N_5704,N_4185,N_4277);
and U5705 (N_5705,N_4164,N_4475);
or U5706 (N_5706,N_4442,N_4418);
nand U5707 (N_5707,N_4660,N_4504);
or U5708 (N_5708,N_4692,N_4924);
nor U5709 (N_5709,N_4447,N_4665);
xnor U5710 (N_5710,N_4765,N_4191);
nand U5711 (N_5711,N_4022,N_4674);
or U5712 (N_5712,N_4590,N_4975);
xor U5713 (N_5713,N_4913,N_4203);
or U5714 (N_5714,N_4920,N_4768);
nor U5715 (N_5715,N_4438,N_4675);
nand U5716 (N_5716,N_4769,N_4119);
xnor U5717 (N_5717,N_4220,N_4126);
and U5718 (N_5718,N_4024,N_4594);
nand U5719 (N_5719,N_4204,N_4335);
and U5720 (N_5720,N_4212,N_4628);
or U5721 (N_5721,N_4713,N_4911);
xnor U5722 (N_5722,N_4105,N_4853);
and U5723 (N_5723,N_4225,N_4686);
nor U5724 (N_5724,N_4460,N_4698);
and U5725 (N_5725,N_4110,N_4220);
nand U5726 (N_5726,N_4624,N_4606);
and U5727 (N_5727,N_4318,N_4300);
or U5728 (N_5728,N_4753,N_4523);
and U5729 (N_5729,N_4675,N_4412);
xnor U5730 (N_5730,N_4644,N_4608);
nor U5731 (N_5731,N_4565,N_4011);
and U5732 (N_5732,N_4577,N_4539);
or U5733 (N_5733,N_4339,N_4616);
nand U5734 (N_5734,N_4774,N_4636);
or U5735 (N_5735,N_4133,N_4193);
xnor U5736 (N_5736,N_4820,N_4300);
xor U5737 (N_5737,N_4418,N_4280);
nor U5738 (N_5738,N_4853,N_4161);
nand U5739 (N_5739,N_4197,N_4981);
xor U5740 (N_5740,N_4981,N_4965);
nor U5741 (N_5741,N_4509,N_4951);
nand U5742 (N_5742,N_4533,N_4536);
nand U5743 (N_5743,N_4195,N_4890);
or U5744 (N_5744,N_4732,N_4028);
and U5745 (N_5745,N_4037,N_4196);
and U5746 (N_5746,N_4206,N_4385);
or U5747 (N_5747,N_4306,N_4588);
xor U5748 (N_5748,N_4631,N_4350);
and U5749 (N_5749,N_4996,N_4781);
nand U5750 (N_5750,N_4905,N_4235);
or U5751 (N_5751,N_4258,N_4238);
nand U5752 (N_5752,N_4769,N_4451);
nand U5753 (N_5753,N_4785,N_4452);
and U5754 (N_5754,N_4389,N_4585);
or U5755 (N_5755,N_4636,N_4043);
nor U5756 (N_5756,N_4196,N_4703);
nor U5757 (N_5757,N_4514,N_4320);
and U5758 (N_5758,N_4384,N_4442);
nand U5759 (N_5759,N_4924,N_4720);
and U5760 (N_5760,N_4960,N_4160);
and U5761 (N_5761,N_4433,N_4236);
nor U5762 (N_5762,N_4795,N_4328);
nand U5763 (N_5763,N_4307,N_4617);
xnor U5764 (N_5764,N_4857,N_4493);
and U5765 (N_5765,N_4741,N_4315);
xnor U5766 (N_5766,N_4829,N_4570);
xnor U5767 (N_5767,N_4943,N_4313);
and U5768 (N_5768,N_4408,N_4392);
or U5769 (N_5769,N_4364,N_4797);
and U5770 (N_5770,N_4699,N_4641);
and U5771 (N_5771,N_4042,N_4478);
xnor U5772 (N_5772,N_4356,N_4812);
xor U5773 (N_5773,N_4199,N_4990);
xnor U5774 (N_5774,N_4887,N_4582);
or U5775 (N_5775,N_4527,N_4917);
and U5776 (N_5776,N_4747,N_4145);
xor U5777 (N_5777,N_4791,N_4442);
nor U5778 (N_5778,N_4943,N_4426);
nor U5779 (N_5779,N_4264,N_4584);
nor U5780 (N_5780,N_4873,N_4697);
nand U5781 (N_5781,N_4282,N_4732);
nor U5782 (N_5782,N_4584,N_4404);
and U5783 (N_5783,N_4869,N_4730);
or U5784 (N_5784,N_4934,N_4508);
nand U5785 (N_5785,N_4437,N_4446);
nor U5786 (N_5786,N_4613,N_4099);
nand U5787 (N_5787,N_4980,N_4134);
or U5788 (N_5788,N_4975,N_4210);
and U5789 (N_5789,N_4113,N_4692);
nand U5790 (N_5790,N_4086,N_4496);
nor U5791 (N_5791,N_4152,N_4011);
and U5792 (N_5792,N_4660,N_4686);
or U5793 (N_5793,N_4507,N_4822);
xnor U5794 (N_5794,N_4086,N_4414);
and U5795 (N_5795,N_4443,N_4191);
or U5796 (N_5796,N_4863,N_4889);
nand U5797 (N_5797,N_4219,N_4347);
xnor U5798 (N_5798,N_4705,N_4520);
xnor U5799 (N_5799,N_4798,N_4837);
nor U5800 (N_5800,N_4390,N_4087);
and U5801 (N_5801,N_4950,N_4334);
nor U5802 (N_5802,N_4127,N_4234);
or U5803 (N_5803,N_4765,N_4482);
xor U5804 (N_5804,N_4861,N_4793);
nor U5805 (N_5805,N_4974,N_4815);
xor U5806 (N_5806,N_4835,N_4815);
and U5807 (N_5807,N_4597,N_4750);
nand U5808 (N_5808,N_4659,N_4806);
xor U5809 (N_5809,N_4157,N_4387);
and U5810 (N_5810,N_4248,N_4518);
xnor U5811 (N_5811,N_4370,N_4578);
xor U5812 (N_5812,N_4758,N_4561);
or U5813 (N_5813,N_4417,N_4725);
nor U5814 (N_5814,N_4286,N_4225);
or U5815 (N_5815,N_4047,N_4200);
or U5816 (N_5816,N_4100,N_4739);
xor U5817 (N_5817,N_4829,N_4634);
nor U5818 (N_5818,N_4133,N_4261);
nand U5819 (N_5819,N_4941,N_4579);
nor U5820 (N_5820,N_4439,N_4370);
and U5821 (N_5821,N_4911,N_4372);
or U5822 (N_5822,N_4659,N_4611);
and U5823 (N_5823,N_4452,N_4434);
and U5824 (N_5824,N_4368,N_4677);
or U5825 (N_5825,N_4135,N_4394);
nand U5826 (N_5826,N_4773,N_4043);
and U5827 (N_5827,N_4170,N_4117);
or U5828 (N_5828,N_4495,N_4803);
xor U5829 (N_5829,N_4973,N_4550);
and U5830 (N_5830,N_4889,N_4115);
xor U5831 (N_5831,N_4722,N_4014);
nor U5832 (N_5832,N_4113,N_4973);
nor U5833 (N_5833,N_4592,N_4032);
or U5834 (N_5834,N_4017,N_4621);
nand U5835 (N_5835,N_4628,N_4301);
and U5836 (N_5836,N_4956,N_4245);
or U5837 (N_5837,N_4973,N_4686);
nor U5838 (N_5838,N_4091,N_4136);
nand U5839 (N_5839,N_4062,N_4207);
and U5840 (N_5840,N_4657,N_4226);
nor U5841 (N_5841,N_4568,N_4976);
xor U5842 (N_5842,N_4980,N_4013);
or U5843 (N_5843,N_4234,N_4530);
nor U5844 (N_5844,N_4763,N_4230);
xor U5845 (N_5845,N_4571,N_4465);
nand U5846 (N_5846,N_4354,N_4505);
and U5847 (N_5847,N_4295,N_4616);
or U5848 (N_5848,N_4328,N_4045);
and U5849 (N_5849,N_4621,N_4481);
and U5850 (N_5850,N_4393,N_4632);
or U5851 (N_5851,N_4526,N_4343);
nor U5852 (N_5852,N_4129,N_4494);
nor U5853 (N_5853,N_4955,N_4987);
nor U5854 (N_5854,N_4742,N_4609);
and U5855 (N_5855,N_4725,N_4256);
nor U5856 (N_5856,N_4618,N_4063);
xor U5857 (N_5857,N_4201,N_4055);
nand U5858 (N_5858,N_4892,N_4106);
xor U5859 (N_5859,N_4626,N_4432);
nand U5860 (N_5860,N_4373,N_4163);
nand U5861 (N_5861,N_4137,N_4899);
nor U5862 (N_5862,N_4981,N_4918);
nor U5863 (N_5863,N_4028,N_4565);
or U5864 (N_5864,N_4973,N_4549);
nor U5865 (N_5865,N_4712,N_4539);
or U5866 (N_5866,N_4986,N_4624);
nor U5867 (N_5867,N_4098,N_4167);
nor U5868 (N_5868,N_4388,N_4216);
xnor U5869 (N_5869,N_4485,N_4129);
and U5870 (N_5870,N_4573,N_4033);
nand U5871 (N_5871,N_4676,N_4534);
xnor U5872 (N_5872,N_4124,N_4435);
xor U5873 (N_5873,N_4521,N_4724);
and U5874 (N_5874,N_4252,N_4225);
nor U5875 (N_5875,N_4871,N_4984);
nand U5876 (N_5876,N_4784,N_4994);
nand U5877 (N_5877,N_4648,N_4470);
and U5878 (N_5878,N_4779,N_4359);
nor U5879 (N_5879,N_4473,N_4373);
xnor U5880 (N_5880,N_4261,N_4307);
or U5881 (N_5881,N_4525,N_4786);
nand U5882 (N_5882,N_4401,N_4844);
xnor U5883 (N_5883,N_4421,N_4996);
nor U5884 (N_5884,N_4946,N_4820);
or U5885 (N_5885,N_4698,N_4612);
xor U5886 (N_5886,N_4340,N_4366);
nor U5887 (N_5887,N_4074,N_4088);
or U5888 (N_5888,N_4235,N_4232);
or U5889 (N_5889,N_4918,N_4985);
or U5890 (N_5890,N_4386,N_4717);
or U5891 (N_5891,N_4386,N_4039);
nand U5892 (N_5892,N_4756,N_4334);
and U5893 (N_5893,N_4196,N_4850);
or U5894 (N_5894,N_4180,N_4884);
or U5895 (N_5895,N_4526,N_4246);
or U5896 (N_5896,N_4123,N_4043);
xnor U5897 (N_5897,N_4595,N_4103);
nand U5898 (N_5898,N_4144,N_4950);
nor U5899 (N_5899,N_4806,N_4422);
nor U5900 (N_5900,N_4073,N_4058);
nor U5901 (N_5901,N_4806,N_4160);
and U5902 (N_5902,N_4046,N_4873);
or U5903 (N_5903,N_4621,N_4496);
nand U5904 (N_5904,N_4208,N_4702);
and U5905 (N_5905,N_4649,N_4063);
xnor U5906 (N_5906,N_4604,N_4839);
nand U5907 (N_5907,N_4418,N_4520);
nand U5908 (N_5908,N_4229,N_4745);
nand U5909 (N_5909,N_4803,N_4421);
nand U5910 (N_5910,N_4989,N_4153);
nand U5911 (N_5911,N_4313,N_4049);
and U5912 (N_5912,N_4202,N_4137);
nor U5913 (N_5913,N_4300,N_4021);
nand U5914 (N_5914,N_4150,N_4019);
and U5915 (N_5915,N_4939,N_4565);
nand U5916 (N_5916,N_4809,N_4917);
xnor U5917 (N_5917,N_4719,N_4564);
or U5918 (N_5918,N_4479,N_4523);
xor U5919 (N_5919,N_4045,N_4053);
nor U5920 (N_5920,N_4719,N_4374);
or U5921 (N_5921,N_4794,N_4648);
or U5922 (N_5922,N_4299,N_4789);
or U5923 (N_5923,N_4096,N_4492);
xnor U5924 (N_5924,N_4958,N_4065);
nor U5925 (N_5925,N_4067,N_4511);
nor U5926 (N_5926,N_4613,N_4934);
xnor U5927 (N_5927,N_4208,N_4366);
and U5928 (N_5928,N_4722,N_4999);
nor U5929 (N_5929,N_4267,N_4623);
nor U5930 (N_5930,N_4566,N_4711);
xor U5931 (N_5931,N_4123,N_4706);
nor U5932 (N_5932,N_4569,N_4496);
xor U5933 (N_5933,N_4775,N_4705);
and U5934 (N_5934,N_4458,N_4183);
and U5935 (N_5935,N_4982,N_4907);
nand U5936 (N_5936,N_4764,N_4936);
nor U5937 (N_5937,N_4535,N_4964);
nand U5938 (N_5938,N_4518,N_4967);
nand U5939 (N_5939,N_4018,N_4727);
nand U5940 (N_5940,N_4277,N_4748);
and U5941 (N_5941,N_4281,N_4926);
xnor U5942 (N_5942,N_4244,N_4026);
nand U5943 (N_5943,N_4717,N_4060);
nand U5944 (N_5944,N_4132,N_4291);
nor U5945 (N_5945,N_4179,N_4530);
nand U5946 (N_5946,N_4913,N_4276);
nand U5947 (N_5947,N_4995,N_4873);
or U5948 (N_5948,N_4635,N_4126);
nand U5949 (N_5949,N_4054,N_4378);
or U5950 (N_5950,N_4351,N_4087);
nor U5951 (N_5951,N_4652,N_4183);
xnor U5952 (N_5952,N_4565,N_4500);
nor U5953 (N_5953,N_4051,N_4809);
or U5954 (N_5954,N_4910,N_4418);
nor U5955 (N_5955,N_4283,N_4573);
xnor U5956 (N_5956,N_4841,N_4440);
nand U5957 (N_5957,N_4924,N_4519);
nor U5958 (N_5958,N_4148,N_4832);
xnor U5959 (N_5959,N_4788,N_4648);
or U5960 (N_5960,N_4757,N_4675);
or U5961 (N_5961,N_4991,N_4394);
and U5962 (N_5962,N_4095,N_4850);
nor U5963 (N_5963,N_4147,N_4574);
or U5964 (N_5964,N_4770,N_4639);
nand U5965 (N_5965,N_4782,N_4281);
and U5966 (N_5966,N_4432,N_4942);
and U5967 (N_5967,N_4597,N_4788);
or U5968 (N_5968,N_4003,N_4680);
or U5969 (N_5969,N_4752,N_4769);
xnor U5970 (N_5970,N_4538,N_4333);
xnor U5971 (N_5971,N_4708,N_4489);
nand U5972 (N_5972,N_4576,N_4808);
nor U5973 (N_5973,N_4902,N_4221);
nand U5974 (N_5974,N_4209,N_4747);
xor U5975 (N_5975,N_4737,N_4639);
xnor U5976 (N_5976,N_4943,N_4487);
xor U5977 (N_5977,N_4110,N_4278);
or U5978 (N_5978,N_4736,N_4554);
xnor U5979 (N_5979,N_4626,N_4976);
or U5980 (N_5980,N_4247,N_4468);
nor U5981 (N_5981,N_4752,N_4732);
nor U5982 (N_5982,N_4111,N_4493);
and U5983 (N_5983,N_4900,N_4048);
and U5984 (N_5984,N_4780,N_4918);
nand U5985 (N_5985,N_4496,N_4159);
nor U5986 (N_5986,N_4540,N_4778);
nand U5987 (N_5987,N_4970,N_4481);
nand U5988 (N_5988,N_4045,N_4215);
xor U5989 (N_5989,N_4484,N_4532);
and U5990 (N_5990,N_4482,N_4528);
xor U5991 (N_5991,N_4190,N_4080);
nand U5992 (N_5992,N_4225,N_4406);
nor U5993 (N_5993,N_4366,N_4251);
or U5994 (N_5994,N_4284,N_4906);
nand U5995 (N_5995,N_4298,N_4733);
and U5996 (N_5996,N_4203,N_4407);
nand U5997 (N_5997,N_4836,N_4988);
or U5998 (N_5998,N_4005,N_4182);
nand U5999 (N_5999,N_4308,N_4349);
nor U6000 (N_6000,N_5015,N_5571);
nor U6001 (N_6001,N_5565,N_5859);
xor U6002 (N_6002,N_5937,N_5832);
nor U6003 (N_6003,N_5659,N_5610);
or U6004 (N_6004,N_5947,N_5851);
and U6005 (N_6005,N_5356,N_5514);
or U6006 (N_6006,N_5127,N_5734);
nor U6007 (N_6007,N_5095,N_5504);
nor U6008 (N_6008,N_5846,N_5310);
nor U6009 (N_6009,N_5838,N_5191);
and U6010 (N_6010,N_5938,N_5032);
xor U6011 (N_6011,N_5968,N_5377);
and U6012 (N_6012,N_5136,N_5464);
or U6013 (N_6013,N_5804,N_5645);
or U6014 (N_6014,N_5570,N_5281);
or U6015 (N_6015,N_5409,N_5339);
xnor U6016 (N_6016,N_5400,N_5745);
xnor U6017 (N_6017,N_5080,N_5455);
and U6018 (N_6018,N_5288,N_5608);
xor U6019 (N_6019,N_5213,N_5410);
nor U6020 (N_6020,N_5665,N_5830);
nor U6021 (N_6021,N_5017,N_5332);
and U6022 (N_6022,N_5869,N_5777);
nor U6023 (N_6023,N_5207,N_5901);
nand U6024 (N_6024,N_5704,N_5681);
nor U6025 (N_6025,N_5496,N_5367);
or U6026 (N_6026,N_5249,N_5722);
nand U6027 (N_6027,N_5396,N_5972);
and U6028 (N_6028,N_5931,N_5460);
nor U6029 (N_6029,N_5557,N_5754);
xor U6030 (N_6030,N_5865,N_5466);
nand U6031 (N_6031,N_5391,N_5178);
nor U6032 (N_6032,N_5533,N_5150);
and U6033 (N_6033,N_5701,N_5203);
and U6034 (N_6034,N_5781,N_5442);
nor U6035 (N_6035,N_5172,N_5697);
nor U6036 (N_6036,N_5433,N_5501);
nand U6037 (N_6037,N_5662,N_5634);
nand U6038 (N_6038,N_5138,N_5027);
xor U6039 (N_6039,N_5583,N_5439);
nand U6040 (N_6040,N_5489,N_5685);
nor U6041 (N_6041,N_5591,N_5967);
nor U6042 (N_6042,N_5341,N_5147);
or U6043 (N_6043,N_5301,N_5067);
and U6044 (N_6044,N_5115,N_5040);
nand U6045 (N_6045,N_5860,N_5693);
and U6046 (N_6046,N_5295,N_5957);
and U6047 (N_6047,N_5453,N_5037);
nand U6048 (N_6048,N_5355,N_5787);
nor U6049 (N_6049,N_5520,N_5075);
nand U6050 (N_6050,N_5818,N_5952);
nand U6051 (N_6051,N_5181,N_5467);
xnor U6052 (N_6052,N_5373,N_5440);
or U6053 (N_6053,N_5180,N_5058);
xor U6054 (N_6054,N_5156,N_5048);
or U6055 (N_6055,N_5904,N_5737);
nand U6056 (N_6056,N_5993,N_5354);
nor U6057 (N_6057,N_5992,N_5555);
xor U6058 (N_6058,N_5061,N_5709);
and U6059 (N_6059,N_5255,N_5268);
xnor U6060 (N_6060,N_5060,N_5184);
or U6061 (N_6061,N_5674,N_5280);
nor U6062 (N_6062,N_5019,N_5471);
nand U6063 (N_6063,N_5870,N_5873);
nand U6064 (N_6064,N_5366,N_5344);
nand U6065 (N_6065,N_5198,N_5554);
or U6066 (N_6066,N_5678,N_5331);
or U6067 (N_6067,N_5448,N_5238);
or U6068 (N_6068,N_5390,N_5862);
xnor U6069 (N_6069,N_5943,N_5969);
and U6070 (N_6070,N_5402,N_5076);
or U6071 (N_6071,N_5602,N_5918);
and U6072 (N_6072,N_5707,N_5145);
nand U6073 (N_6073,N_5793,N_5105);
xnor U6074 (N_6074,N_5671,N_5603);
or U6075 (N_6075,N_5677,N_5960);
or U6076 (N_6076,N_5796,N_5511);
nor U6077 (N_6077,N_5168,N_5985);
xor U6078 (N_6078,N_5413,N_5124);
nor U6079 (N_6079,N_5126,N_5179);
or U6080 (N_6080,N_5979,N_5007);
xor U6081 (N_6081,N_5392,N_5300);
nand U6082 (N_6082,N_5617,N_5654);
nand U6083 (N_6083,N_5166,N_5908);
and U6084 (N_6084,N_5534,N_5286);
nor U6085 (N_6085,N_5899,N_5429);
xor U6086 (N_6086,N_5578,N_5732);
or U6087 (N_6087,N_5944,N_5463);
nand U6088 (N_6088,N_5443,N_5399);
nand U6089 (N_6089,N_5503,N_5766);
nand U6090 (N_6090,N_5562,N_5327);
xnor U6091 (N_6091,N_5680,N_5871);
or U6092 (N_6092,N_5199,N_5539);
or U6093 (N_6093,N_5164,N_5119);
and U6094 (N_6094,N_5498,N_5990);
xnor U6095 (N_6095,N_5461,N_5560);
or U6096 (N_6096,N_5529,N_5921);
and U6097 (N_6097,N_5389,N_5093);
and U6098 (N_6098,N_5275,N_5326);
xor U6099 (N_6099,N_5381,N_5933);
or U6100 (N_6100,N_5369,N_5744);
nand U6101 (N_6101,N_5306,N_5502);
xnor U6102 (N_6102,N_5710,N_5879);
or U6103 (N_6103,N_5430,N_5222);
nand U6104 (N_6104,N_5053,N_5891);
and U6105 (N_6105,N_5973,N_5609);
nor U6106 (N_6106,N_5927,N_5508);
and U6107 (N_6107,N_5417,N_5196);
or U6108 (N_6108,N_5371,N_5308);
xnor U6109 (N_6109,N_5597,N_5867);
nand U6110 (N_6110,N_5346,N_5641);
or U6111 (N_6111,N_5739,N_5197);
xnor U6112 (N_6112,N_5393,N_5692);
nor U6113 (N_6113,N_5094,N_5506);
nor U6114 (N_6114,N_5995,N_5585);
xor U6115 (N_6115,N_5436,N_5828);
or U6116 (N_6116,N_5526,N_5507);
nor U6117 (N_6117,N_5230,N_5619);
xnor U6118 (N_6118,N_5073,N_5458);
nand U6119 (N_6119,N_5167,N_5427);
nand U6120 (N_6120,N_5253,N_5765);
nand U6121 (N_6121,N_5111,N_5205);
xnor U6122 (N_6122,N_5621,N_5157);
and U6123 (N_6123,N_5270,N_5449);
nand U6124 (N_6124,N_5258,N_5378);
xor U6125 (N_6125,N_5160,N_5232);
or U6126 (N_6126,N_5140,N_5065);
nor U6127 (N_6127,N_5472,N_5782);
xor U6128 (N_6128,N_5117,N_5630);
or U6129 (N_6129,N_5083,N_5850);
nor U6130 (N_6130,N_5013,N_5182);
xor U6131 (N_6131,N_5260,N_5866);
or U6132 (N_6132,N_5236,N_5579);
or U6133 (N_6133,N_5043,N_5062);
or U6134 (N_6134,N_5081,N_5741);
or U6135 (N_6135,N_5349,N_5755);
xor U6136 (N_6136,N_5546,N_5883);
nand U6137 (N_6137,N_5102,N_5868);
and U6138 (N_6138,N_5171,N_5971);
xnor U6139 (N_6139,N_5499,N_5452);
nand U6140 (N_6140,N_5801,N_5760);
xor U6141 (N_6141,N_5437,N_5002);
nand U6142 (N_6142,N_5233,N_5623);
or U6143 (N_6143,N_5468,N_5844);
and U6144 (N_6144,N_5494,N_5008);
nand U6145 (N_6145,N_5715,N_5450);
or U6146 (N_6146,N_5813,N_5807);
or U6147 (N_6147,N_5465,N_5663);
nand U6148 (N_6148,N_5816,N_5613);
or U6149 (N_6149,N_5438,N_5042);
nand U6150 (N_6150,N_5107,N_5989);
nor U6151 (N_6151,N_5540,N_5314);
and U6152 (N_6152,N_5978,N_5601);
xor U6153 (N_6153,N_5895,N_5379);
and U6154 (N_6154,N_5840,N_5731);
or U6155 (N_6155,N_5342,N_5764);
nand U6156 (N_6156,N_5997,N_5955);
nor U6157 (N_6157,N_5375,N_5607);
nor U6158 (N_6158,N_5423,N_5114);
nand U6159 (N_6159,N_5185,N_5950);
or U6160 (N_6160,N_5551,N_5626);
nor U6161 (N_6161,N_5852,N_5872);
and U6162 (N_6162,N_5970,N_5987);
or U6163 (N_6163,N_5477,N_5118);
nand U6164 (N_6164,N_5194,N_5202);
or U6165 (N_6165,N_5545,N_5330);
nand U6166 (N_6166,N_5885,N_5385);
xnor U6167 (N_6167,N_5337,N_5475);
xnor U6168 (N_6168,N_5652,N_5237);
and U6169 (N_6169,N_5387,N_5509);
xor U6170 (N_6170,N_5264,N_5047);
and U6171 (N_6171,N_5163,N_5836);
xor U6172 (N_6172,N_5404,N_5549);
xor U6173 (N_6173,N_5696,N_5414);
nor U6174 (N_6174,N_5915,N_5292);
xor U6175 (N_6175,N_5352,N_5650);
or U6176 (N_6176,N_5541,N_5077);
and U6177 (N_6177,N_5577,N_5309);
or U6178 (N_6178,N_5024,N_5316);
nor U6179 (N_6179,N_5815,N_5220);
xnor U6180 (N_6180,N_5240,N_5112);
nor U6181 (N_6181,N_5071,N_5620);
and U6182 (N_6182,N_5018,N_5359);
or U6183 (N_6183,N_5996,N_5384);
nor U6184 (N_6184,N_5717,N_5149);
and U6185 (N_6185,N_5099,N_5357);
nand U6186 (N_6186,N_5824,N_5833);
nand U6187 (N_6187,N_5778,N_5667);
and U6188 (N_6188,N_5587,N_5687);
or U6189 (N_6189,N_5211,N_5057);
nor U6190 (N_6190,N_5962,N_5311);
xnor U6191 (N_6191,N_5842,N_5016);
or U6192 (N_6192,N_5059,N_5487);
nor U6193 (N_6193,N_5284,N_5383);
nor U6194 (N_6194,N_5447,N_5478);
and U6195 (N_6195,N_5805,N_5473);
or U6196 (N_6196,N_5274,N_5939);
nand U6197 (N_6197,N_5817,N_5774);
xnor U6198 (N_6198,N_5605,N_5748);
nand U6199 (N_6199,N_5435,N_5064);
nor U6200 (N_6200,N_5561,N_5757);
nor U6201 (N_6201,N_5513,N_5044);
nor U6202 (N_6202,N_5001,N_5457);
and U6203 (N_6203,N_5700,N_5797);
xnor U6204 (N_6204,N_5906,N_5874);
nand U6205 (N_6205,N_5627,N_5820);
or U6206 (N_6206,N_5313,N_5209);
and U6207 (N_6207,N_5082,N_5364);
nand U6208 (N_6208,N_5679,N_5034);
or U6209 (N_6209,N_5718,N_5532);
or U6210 (N_6210,N_5515,N_5011);
nor U6211 (N_6211,N_5988,N_5576);
nand U6212 (N_6212,N_5454,N_5505);
nand U6213 (N_6213,N_5252,N_5103);
nor U6214 (N_6214,N_5776,N_5386);
and U6215 (N_6215,N_5733,N_5293);
nand U6216 (N_6216,N_5090,N_5257);
and U6217 (N_6217,N_5312,N_5175);
or U6218 (N_6218,N_5703,N_5829);
xnor U6219 (N_6219,N_5497,N_5854);
or U6220 (N_6220,N_5265,N_5035);
nand U6221 (N_6221,N_5686,N_5033);
or U6222 (N_6222,N_5474,N_5097);
or U6223 (N_6223,N_5319,N_5800);
and U6224 (N_6224,N_5289,N_5631);
and U6225 (N_6225,N_5122,N_5495);
and U6226 (N_6226,N_5451,N_5537);
nand U6227 (N_6227,N_5742,N_5078);
xor U6228 (N_6228,N_5266,N_5759);
or U6229 (N_6229,N_5790,N_5961);
xor U6230 (N_6230,N_5282,N_5050);
nor U6231 (N_6231,N_5304,N_5045);
xor U6232 (N_6232,N_5155,N_5618);
or U6233 (N_6233,N_5231,N_5900);
and U6234 (N_6234,N_5923,N_5821);
nand U6235 (N_6235,N_5169,N_5596);
xor U6236 (N_6236,N_5638,N_5177);
nor U6237 (N_6237,N_5022,N_5669);
and U6238 (N_6238,N_5750,N_5806);
or U6239 (N_6239,N_5930,N_5758);
nand U6240 (N_6240,N_5553,N_5984);
nand U6241 (N_6241,N_5317,N_5581);
nor U6242 (N_6242,N_5695,N_5738);
nand U6243 (N_6243,N_5370,N_5843);
nor U6244 (N_6244,N_5910,N_5153);
nand U6245 (N_6245,N_5643,N_5835);
xnor U6246 (N_6246,N_5142,N_5857);
nor U6247 (N_6247,N_5676,N_5418);
xor U6248 (N_6248,N_5000,N_5794);
or U6249 (N_6249,N_5350,N_5644);
nand U6250 (N_6250,N_5227,N_5148);
nor U6251 (N_6251,N_5706,N_5134);
and U6252 (N_6252,N_5010,N_5974);
or U6253 (N_6253,N_5586,N_5049);
or U6254 (N_6254,N_5861,N_5212);
and U6255 (N_6255,N_5791,N_5360);
and U6256 (N_6256,N_5642,N_5522);
and U6257 (N_6257,N_5006,N_5711);
xor U6258 (N_6258,N_5298,N_5510);
nand U6259 (N_6259,N_5420,N_5285);
or U6260 (N_6260,N_5792,N_5544);
and U6261 (N_6261,N_5085,N_5951);
nand U6262 (N_6262,N_5550,N_5982);
xnor U6263 (N_6263,N_5320,N_5247);
nand U6264 (N_6264,N_5855,N_5566);
nor U6265 (N_6265,N_5176,N_5219);
and U6266 (N_6266,N_5538,N_5720);
and U6267 (N_6267,N_5143,N_5195);
or U6268 (N_6268,N_5116,N_5485);
xnor U6269 (N_6269,N_5547,N_5023);
or U6270 (N_6270,N_5848,N_5096);
nor U6271 (N_6271,N_5432,N_5315);
and U6272 (N_6272,N_5876,N_5535);
nand U6273 (N_6273,N_5651,N_5214);
xnor U6274 (N_6274,N_5481,N_5347);
xor U6275 (N_6275,N_5031,N_5936);
nor U6276 (N_6276,N_5500,N_5159);
and U6277 (N_6277,N_5810,N_5382);
nand U6278 (N_6278,N_5524,N_5411);
or U6279 (N_6279,N_5629,N_5291);
nand U6280 (N_6280,N_5029,N_5958);
nand U6281 (N_6281,N_5849,N_5753);
nand U6282 (N_6282,N_5580,N_5063);
or U6283 (N_6283,N_5421,N_5215);
and U6284 (N_6284,N_5137,N_5132);
xor U6285 (N_6285,N_5523,N_5056);
or U6286 (N_6286,N_5917,N_5615);
xnor U6287 (N_6287,N_5784,N_5959);
nand U6288 (N_6288,N_5991,N_5834);
and U6289 (N_6289,N_5726,N_5636);
nand U6290 (N_6290,N_5548,N_5558);
and U6291 (N_6291,N_5600,N_5980);
nor U6292 (N_6292,N_5660,N_5491);
xnor U6293 (N_6293,N_5953,N_5809);
nor U6294 (N_6294,N_5922,N_5469);
nand U6295 (N_6295,N_5273,N_5694);
or U6296 (N_6296,N_5814,N_5217);
or U6297 (N_6297,N_5092,N_5763);
nand U6298 (N_6298,N_5756,N_5186);
nand U6299 (N_6299,N_5747,N_5584);
nor U6300 (N_6300,N_5261,N_5878);
nor U6301 (N_6301,N_5788,N_5445);
xnor U6302 (N_6302,N_5530,N_5599);
nor U6303 (N_6303,N_5446,N_5303);
xnor U6304 (N_6304,N_5569,N_5305);
nand U6305 (N_6305,N_5574,N_5831);
and U6306 (N_6306,N_5907,N_5892);
xnor U6307 (N_6307,N_5789,N_5552);
xnor U6308 (N_6308,N_5779,N_5089);
nand U6309 (N_6309,N_5072,N_5785);
xor U6310 (N_6310,N_5087,N_5276);
or U6311 (N_6311,N_5682,N_5318);
or U6312 (N_6312,N_5259,N_5129);
nor U6313 (N_6313,N_5716,N_5604);
nor U6314 (N_6314,N_5307,N_5690);
and U6315 (N_6315,N_5773,N_5684);
nor U6316 (N_6316,N_5322,N_5190);
xnor U6317 (N_6317,N_5724,N_5877);
or U6318 (N_6318,N_5456,N_5909);
xor U6319 (N_6319,N_5655,N_5484);
xnor U6320 (N_6320,N_5647,N_5141);
xnor U6321 (N_6321,N_5903,N_5424);
and U6322 (N_6322,N_5568,N_5896);
xnor U6323 (N_6323,N_5070,N_5088);
or U6324 (N_6324,N_5795,N_5054);
or U6325 (N_6325,N_5911,N_5752);
nor U6326 (N_6326,N_5898,N_5395);
xnor U6327 (N_6327,N_5106,N_5702);
or U6328 (N_6328,N_5165,N_5727);
xor U6329 (N_6329,N_5372,N_5986);
and U6330 (N_6330,N_5287,N_5130);
nand U6331 (N_6331,N_5086,N_5296);
and U6332 (N_6332,N_5735,N_5334);
and U6333 (N_6333,N_5902,N_5527);
xnor U6334 (N_6334,N_5775,N_5225);
xor U6335 (N_6335,N_5368,N_5812);
or U6336 (N_6336,N_5021,N_5929);
and U6337 (N_6337,N_5786,N_5653);
xor U6338 (N_6338,N_5633,N_5808);
or U6339 (N_6339,N_5761,N_5799);
and U6340 (N_6340,N_5003,N_5193);
or U6341 (N_6341,N_5245,N_5210);
and U6342 (N_6342,N_5740,N_5912);
xnor U6343 (N_6343,N_5241,N_5632);
nand U6344 (N_6344,N_5407,N_5769);
nand U6345 (N_6345,N_5039,N_5161);
nor U6346 (N_6346,N_5234,N_5590);
xnor U6347 (N_6347,N_5595,N_5736);
nor U6348 (N_6348,N_5277,N_5323);
nor U6349 (N_6349,N_5128,N_5052);
nand U6350 (N_6350,N_5925,N_5123);
nor U6351 (N_6351,N_5428,N_5598);
nand U6352 (N_6352,N_5699,N_5847);
or U6353 (N_6353,N_5672,N_5675);
nor U6354 (N_6354,N_5256,N_5622);
nor U6355 (N_6355,N_5068,N_5783);
and U6356 (N_6356,N_5459,N_5888);
or U6357 (N_6357,N_5336,N_5624);
or U6358 (N_6358,N_5593,N_5994);
and U6359 (N_6359,N_5920,N_5218);
and U6360 (N_6360,N_5353,N_5826);
nor U6361 (N_6361,N_5963,N_5490);
or U6362 (N_6362,N_5188,N_5966);
xnor U6363 (N_6363,N_5723,N_5954);
xnor U6364 (N_6364,N_5762,N_5041);
xnor U6365 (N_6365,N_5154,N_5625);
and U6366 (N_6366,N_5248,N_5964);
nand U6367 (N_6367,N_5030,N_5144);
or U6368 (N_6368,N_5856,N_5894);
xor U6369 (N_6369,N_5983,N_5721);
and U6370 (N_6370,N_5708,N_5683);
or U6371 (N_6371,N_5380,N_5542);
or U6372 (N_6372,N_5434,N_5657);
nor U6373 (N_6373,N_5251,N_5528);
or U6374 (N_6374,N_5361,N_5751);
nor U6375 (N_6375,N_5668,N_5516);
or U6376 (N_6376,N_5426,N_5839);
xor U6377 (N_6377,N_5493,N_5229);
or U6378 (N_6378,N_5567,N_5882);
or U6379 (N_6379,N_5208,N_5333);
and U6380 (N_6380,N_5940,N_5729);
nand U6381 (N_6381,N_5228,N_5131);
nand U6382 (N_6382,N_5269,N_5412);
nand U6383 (N_6383,N_5109,N_5345);
nor U6384 (N_6384,N_5321,N_5004);
or U6385 (N_6385,N_5946,N_5572);
or U6386 (N_6386,N_5363,N_5698);
and U6387 (N_6387,N_5730,N_5556);
xor U6388 (N_6388,N_5594,N_5290);
and U6389 (N_6389,N_5863,N_5376);
nand U6390 (N_6390,N_5913,N_5243);
and U6391 (N_6391,N_5246,N_5005);
or U6392 (N_6392,N_5559,N_5640);
nand U6393 (N_6393,N_5374,N_5173);
or U6394 (N_6394,N_5803,N_5462);
and U6395 (N_6395,N_5479,N_5771);
xnor U6396 (N_6396,N_5250,N_5670);
and U6397 (N_6397,N_5074,N_5827);
xnor U6398 (N_6398,N_5351,N_5798);
nand U6399 (N_6399,N_5201,N_5325);
and U6400 (N_6400,N_5661,N_5531);
nor U6401 (N_6401,N_5837,N_5588);
nor U6402 (N_6402,N_5924,N_5388);
and U6403 (N_6403,N_5853,N_5408);
xor U6404 (N_6404,N_5612,N_5880);
xor U6405 (N_6405,N_5934,N_5294);
nor U6406 (N_6406,N_5046,N_5328);
xnor U6407 (N_6407,N_5406,N_5575);
and U6408 (N_6408,N_5822,N_5066);
nor U6409 (N_6409,N_5932,N_5401);
and U6410 (N_6410,N_5151,N_5705);
or U6411 (N_6411,N_5614,N_5444);
nand U6412 (N_6412,N_5398,N_5025);
nand U6413 (N_6413,N_5884,N_5101);
nor U6414 (N_6414,N_5152,N_5014);
or U6415 (N_6415,N_5483,N_5965);
and U6416 (N_6416,N_5656,N_5324);
or U6417 (N_6417,N_5864,N_5422);
nand U6418 (N_6418,N_5226,N_5297);
and U6419 (N_6419,N_5646,N_5135);
xnor U6420 (N_6420,N_5975,N_5518);
nor U6421 (N_6421,N_5441,N_5713);
nand U6422 (N_6422,N_5365,N_5881);
or U6423 (N_6423,N_5926,N_5712);
and U6424 (N_6424,N_5886,N_5767);
or U6425 (N_6425,N_5512,N_5139);
xor U6426 (N_6426,N_5028,N_5725);
or U6427 (N_6427,N_5121,N_5564);
nor U6428 (N_6428,N_5343,N_5875);
or U6429 (N_6429,N_5492,N_5020);
or U6430 (N_6430,N_5714,N_5329);
and U6431 (N_6431,N_5893,N_5768);
nor U6432 (N_6432,N_5948,N_5905);
or U6433 (N_6433,N_5525,N_5486);
xnor U6434 (N_6434,N_5976,N_5942);
nand U6435 (N_6435,N_5611,N_5649);
nor U6436 (N_6436,N_5916,N_5267);
xnor U6437 (N_6437,N_5397,N_5666);
and U6438 (N_6438,N_5235,N_5819);
nand U6439 (N_6439,N_5224,N_5802);
and U6440 (N_6440,N_5935,N_5914);
or U6441 (N_6441,N_5519,N_5302);
xor U6442 (N_6442,N_5482,N_5606);
nor U6443 (N_6443,N_5858,N_5338);
and U6444 (N_6444,N_5887,N_5981);
and U6445 (N_6445,N_5949,N_5691);
and U6446 (N_6446,N_5146,N_5394);
nor U6447 (N_6447,N_5823,N_5012);
and U6448 (N_6448,N_5480,N_5100);
nand U6449 (N_6449,N_5582,N_5162);
or U6450 (N_6450,N_5091,N_5084);
and U6451 (N_6451,N_5897,N_5746);
or U6452 (N_6452,N_5416,N_5271);
xor U6453 (N_6453,N_5928,N_5592);
or U6454 (N_6454,N_5223,N_5299);
nand U6455 (N_6455,N_5216,N_5113);
nand U6456 (N_6456,N_5919,N_5728);
or U6457 (N_6457,N_5108,N_5637);
and U6458 (N_6458,N_5780,N_5104);
or U6459 (N_6459,N_5689,N_5956);
nand U6460 (N_6460,N_5476,N_5069);
nor U6461 (N_6461,N_5348,N_5200);
or U6462 (N_6462,N_5340,N_5616);
or U6463 (N_6463,N_5573,N_5415);
or U6464 (N_6464,N_5536,N_5628);
and U6465 (N_6465,N_5998,N_5405);
and U6466 (N_6466,N_5335,N_5770);
nor U6467 (N_6467,N_5825,N_5719);
nand U6468 (N_6468,N_5009,N_5183);
nand U6469 (N_6469,N_5563,N_5125);
nand U6470 (N_6470,N_5192,N_5036);
xnor U6471 (N_6471,N_5244,N_5811);
xor U6472 (N_6472,N_5889,N_5890);
nand U6473 (N_6473,N_5589,N_5488);
nor U6474 (N_6474,N_5977,N_5051);
xor U6475 (N_6475,N_5425,N_5279);
xor U6476 (N_6476,N_5945,N_5079);
or U6477 (N_6477,N_5204,N_5026);
nor U6478 (N_6478,N_5263,N_5470);
and U6479 (N_6479,N_5110,N_5120);
and U6480 (N_6480,N_5187,N_5221);
nand U6481 (N_6481,N_5431,N_5262);
nor U6482 (N_6482,N_5206,N_5688);
nor U6483 (N_6483,N_5648,N_5664);
and U6484 (N_6484,N_5658,N_5133);
nand U6485 (N_6485,N_5743,N_5098);
xor U6486 (N_6486,N_5358,N_5845);
xor U6487 (N_6487,N_5055,N_5403);
or U6488 (N_6488,N_5841,N_5170);
nand U6489 (N_6489,N_5239,N_5174);
and U6490 (N_6490,N_5941,N_5189);
or U6491 (N_6491,N_5272,N_5517);
xor U6492 (N_6492,N_5254,N_5158);
xor U6493 (N_6493,N_5543,N_5639);
xor U6494 (N_6494,N_5278,N_5521);
and U6495 (N_6495,N_5283,N_5242);
nand U6496 (N_6496,N_5772,N_5999);
and U6497 (N_6497,N_5419,N_5635);
nor U6498 (N_6498,N_5362,N_5749);
and U6499 (N_6499,N_5673,N_5038);
and U6500 (N_6500,N_5353,N_5761);
or U6501 (N_6501,N_5838,N_5386);
nor U6502 (N_6502,N_5096,N_5870);
or U6503 (N_6503,N_5301,N_5177);
or U6504 (N_6504,N_5254,N_5443);
nor U6505 (N_6505,N_5076,N_5791);
xnor U6506 (N_6506,N_5311,N_5350);
nand U6507 (N_6507,N_5627,N_5915);
or U6508 (N_6508,N_5406,N_5931);
nand U6509 (N_6509,N_5294,N_5337);
nor U6510 (N_6510,N_5136,N_5736);
or U6511 (N_6511,N_5574,N_5434);
nand U6512 (N_6512,N_5889,N_5604);
xnor U6513 (N_6513,N_5468,N_5504);
or U6514 (N_6514,N_5203,N_5109);
or U6515 (N_6515,N_5291,N_5141);
xor U6516 (N_6516,N_5240,N_5592);
nor U6517 (N_6517,N_5566,N_5658);
and U6518 (N_6518,N_5906,N_5123);
or U6519 (N_6519,N_5975,N_5341);
xor U6520 (N_6520,N_5114,N_5553);
nor U6521 (N_6521,N_5598,N_5906);
xor U6522 (N_6522,N_5703,N_5317);
nand U6523 (N_6523,N_5731,N_5577);
or U6524 (N_6524,N_5726,N_5643);
or U6525 (N_6525,N_5678,N_5227);
or U6526 (N_6526,N_5577,N_5068);
xor U6527 (N_6527,N_5774,N_5978);
or U6528 (N_6528,N_5215,N_5623);
nand U6529 (N_6529,N_5147,N_5428);
nor U6530 (N_6530,N_5812,N_5168);
nor U6531 (N_6531,N_5686,N_5298);
nand U6532 (N_6532,N_5887,N_5693);
and U6533 (N_6533,N_5094,N_5021);
xnor U6534 (N_6534,N_5947,N_5659);
nand U6535 (N_6535,N_5799,N_5220);
xnor U6536 (N_6536,N_5409,N_5731);
nor U6537 (N_6537,N_5583,N_5365);
xnor U6538 (N_6538,N_5694,N_5221);
and U6539 (N_6539,N_5953,N_5623);
xnor U6540 (N_6540,N_5416,N_5293);
nand U6541 (N_6541,N_5907,N_5002);
nor U6542 (N_6542,N_5116,N_5456);
nand U6543 (N_6543,N_5828,N_5533);
or U6544 (N_6544,N_5200,N_5933);
or U6545 (N_6545,N_5785,N_5963);
nand U6546 (N_6546,N_5429,N_5123);
nor U6547 (N_6547,N_5733,N_5161);
and U6548 (N_6548,N_5098,N_5518);
and U6549 (N_6549,N_5557,N_5618);
nand U6550 (N_6550,N_5173,N_5212);
xor U6551 (N_6551,N_5995,N_5965);
and U6552 (N_6552,N_5357,N_5432);
and U6553 (N_6553,N_5505,N_5217);
nand U6554 (N_6554,N_5814,N_5249);
xnor U6555 (N_6555,N_5625,N_5178);
and U6556 (N_6556,N_5217,N_5833);
and U6557 (N_6557,N_5220,N_5983);
xor U6558 (N_6558,N_5397,N_5969);
or U6559 (N_6559,N_5903,N_5153);
nor U6560 (N_6560,N_5088,N_5381);
nor U6561 (N_6561,N_5081,N_5651);
and U6562 (N_6562,N_5013,N_5323);
nand U6563 (N_6563,N_5014,N_5409);
nand U6564 (N_6564,N_5965,N_5773);
xnor U6565 (N_6565,N_5160,N_5588);
nor U6566 (N_6566,N_5110,N_5075);
xnor U6567 (N_6567,N_5347,N_5643);
and U6568 (N_6568,N_5060,N_5967);
or U6569 (N_6569,N_5785,N_5731);
and U6570 (N_6570,N_5171,N_5197);
and U6571 (N_6571,N_5268,N_5148);
and U6572 (N_6572,N_5522,N_5282);
nor U6573 (N_6573,N_5628,N_5303);
xor U6574 (N_6574,N_5131,N_5480);
and U6575 (N_6575,N_5008,N_5410);
and U6576 (N_6576,N_5268,N_5430);
and U6577 (N_6577,N_5906,N_5107);
and U6578 (N_6578,N_5035,N_5455);
xnor U6579 (N_6579,N_5550,N_5062);
and U6580 (N_6580,N_5937,N_5865);
xor U6581 (N_6581,N_5234,N_5657);
xnor U6582 (N_6582,N_5904,N_5456);
nor U6583 (N_6583,N_5763,N_5094);
xnor U6584 (N_6584,N_5234,N_5542);
and U6585 (N_6585,N_5058,N_5720);
nor U6586 (N_6586,N_5805,N_5096);
and U6587 (N_6587,N_5252,N_5645);
nor U6588 (N_6588,N_5992,N_5050);
or U6589 (N_6589,N_5651,N_5121);
xnor U6590 (N_6590,N_5045,N_5873);
nand U6591 (N_6591,N_5631,N_5673);
nor U6592 (N_6592,N_5140,N_5288);
nor U6593 (N_6593,N_5557,N_5707);
nor U6594 (N_6594,N_5142,N_5701);
nor U6595 (N_6595,N_5952,N_5991);
or U6596 (N_6596,N_5799,N_5892);
nand U6597 (N_6597,N_5384,N_5688);
and U6598 (N_6598,N_5139,N_5597);
xor U6599 (N_6599,N_5368,N_5733);
or U6600 (N_6600,N_5064,N_5247);
nor U6601 (N_6601,N_5193,N_5408);
xor U6602 (N_6602,N_5586,N_5387);
and U6603 (N_6603,N_5666,N_5750);
nand U6604 (N_6604,N_5507,N_5308);
and U6605 (N_6605,N_5776,N_5023);
nand U6606 (N_6606,N_5623,N_5181);
and U6607 (N_6607,N_5760,N_5236);
or U6608 (N_6608,N_5988,N_5930);
nand U6609 (N_6609,N_5776,N_5468);
or U6610 (N_6610,N_5682,N_5679);
and U6611 (N_6611,N_5892,N_5838);
nand U6612 (N_6612,N_5048,N_5829);
nor U6613 (N_6613,N_5113,N_5569);
nand U6614 (N_6614,N_5374,N_5714);
or U6615 (N_6615,N_5862,N_5606);
nor U6616 (N_6616,N_5856,N_5812);
nor U6617 (N_6617,N_5077,N_5712);
nand U6618 (N_6618,N_5000,N_5775);
nand U6619 (N_6619,N_5269,N_5242);
or U6620 (N_6620,N_5175,N_5237);
or U6621 (N_6621,N_5763,N_5224);
nand U6622 (N_6622,N_5425,N_5380);
or U6623 (N_6623,N_5174,N_5175);
xnor U6624 (N_6624,N_5214,N_5737);
and U6625 (N_6625,N_5335,N_5671);
nand U6626 (N_6626,N_5003,N_5349);
and U6627 (N_6627,N_5869,N_5720);
and U6628 (N_6628,N_5376,N_5385);
nor U6629 (N_6629,N_5541,N_5732);
and U6630 (N_6630,N_5603,N_5567);
nand U6631 (N_6631,N_5574,N_5541);
or U6632 (N_6632,N_5684,N_5399);
or U6633 (N_6633,N_5146,N_5180);
xor U6634 (N_6634,N_5131,N_5939);
or U6635 (N_6635,N_5002,N_5191);
xor U6636 (N_6636,N_5572,N_5677);
or U6637 (N_6637,N_5408,N_5866);
and U6638 (N_6638,N_5436,N_5383);
or U6639 (N_6639,N_5402,N_5594);
nand U6640 (N_6640,N_5354,N_5416);
nor U6641 (N_6641,N_5331,N_5594);
nor U6642 (N_6642,N_5022,N_5133);
nor U6643 (N_6643,N_5825,N_5795);
nand U6644 (N_6644,N_5615,N_5214);
or U6645 (N_6645,N_5264,N_5719);
and U6646 (N_6646,N_5195,N_5973);
xnor U6647 (N_6647,N_5005,N_5510);
nor U6648 (N_6648,N_5454,N_5144);
or U6649 (N_6649,N_5945,N_5693);
and U6650 (N_6650,N_5299,N_5043);
nor U6651 (N_6651,N_5448,N_5393);
or U6652 (N_6652,N_5198,N_5353);
or U6653 (N_6653,N_5002,N_5464);
or U6654 (N_6654,N_5254,N_5948);
and U6655 (N_6655,N_5440,N_5863);
and U6656 (N_6656,N_5892,N_5915);
nand U6657 (N_6657,N_5803,N_5059);
or U6658 (N_6658,N_5812,N_5354);
nand U6659 (N_6659,N_5196,N_5080);
nor U6660 (N_6660,N_5935,N_5085);
nor U6661 (N_6661,N_5293,N_5663);
nor U6662 (N_6662,N_5908,N_5676);
nor U6663 (N_6663,N_5036,N_5682);
and U6664 (N_6664,N_5789,N_5534);
nand U6665 (N_6665,N_5101,N_5129);
nand U6666 (N_6666,N_5679,N_5874);
nor U6667 (N_6667,N_5059,N_5185);
and U6668 (N_6668,N_5970,N_5917);
nor U6669 (N_6669,N_5000,N_5027);
or U6670 (N_6670,N_5133,N_5229);
nand U6671 (N_6671,N_5286,N_5930);
xor U6672 (N_6672,N_5741,N_5931);
nor U6673 (N_6673,N_5332,N_5909);
xnor U6674 (N_6674,N_5200,N_5454);
nor U6675 (N_6675,N_5956,N_5279);
nor U6676 (N_6676,N_5536,N_5082);
xnor U6677 (N_6677,N_5518,N_5523);
or U6678 (N_6678,N_5602,N_5164);
xor U6679 (N_6679,N_5120,N_5012);
xnor U6680 (N_6680,N_5978,N_5624);
nor U6681 (N_6681,N_5580,N_5856);
nor U6682 (N_6682,N_5673,N_5690);
xor U6683 (N_6683,N_5277,N_5717);
nand U6684 (N_6684,N_5887,N_5013);
nand U6685 (N_6685,N_5660,N_5976);
and U6686 (N_6686,N_5867,N_5561);
or U6687 (N_6687,N_5542,N_5434);
or U6688 (N_6688,N_5986,N_5065);
nor U6689 (N_6689,N_5840,N_5816);
nand U6690 (N_6690,N_5787,N_5477);
xnor U6691 (N_6691,N_5153,N_5907);
xnor U6692 (N_6692,N_5441,N_5717);
or U6693 (N_6693,N_5829,N_5082);
and U6694 (N_6694,N_5656,N_5691);
xnor U6695 (N_6695,N_5280,N_5865);
nor U6696 (N_6696,N_5529,N_5643);
nand U6697 (N_6697,N_5013,N_5017);
and U6698 (N_6698,N_5295,N_5403);
and U6699 (N_6699,N_5303,N_5475);
and U6700 (N_6700,N_5609,N_5926);
nand U6701 (N_6701,N_5689,N_5329);
and U6702 (N_6702,N_5771,N_5589);
xor U6703 (N_6703,N_5270,N_5489);
and U6704 (N_6704,N_5111,N_5088);
nand U6705 (N_6705,N_5419,N_5630);
or U6706 (N_6706,N_5033,N_5538);
and U6707 (N_6707,N_5606,N_5810);
and U6708 (N_6708,N_5071,N_5297);
and U6709 (N_6709,N_5770,N_5665);
or U6710 (N_6710,N_5016,N_5326);
or U6711 (N_6711,N_5827,N_5793);
and U6712 (N_6712,N_5341,N_5861);
xor U6713 (N_6713,N_5547,N_5636);
nor U6714 (N_6714,N_5556,N_5962);
or U6715 (N_6715,N_5792,N_5657);
and U6716 (N_6716,N_5690,N_5922);
nand U6717 (N_6717,N_5471,N_5920);
xnor U6718 (N_6718,N_5897,N_5588);
and U6719 (N_6719,N_5805,N_5011);
xnor U6720 (N_6720,N_5340,N_5908);
nor U6721 (N_6721,N_5577,N_5256);
and U6722 (N_6722,N_5480,N_5137);
nor U6723 (N_6723,N_5144,N_5957);
and U6724 (N_6724,N_5113,N_5406);
xnor U6725 (N_6725,N_5391,N_5838);
or U6726 (N_6726,N_5325,N_5697);
or U6727 (N_6727,N_5278,N_5026);
or U6728 (N_6728,N_5272,N_5688);
or U6729 (N_6729,N_5242,N_5362);
nand U6730 (N_6730,N_5787,N_5144);
or U6731 (N_6731,N_5915,N_5883);
or U6732 (N_6732,N_5176,N_5139);
or U6733 (N_6733,N_5654,N_5609);
nand U6734 (N_6734,N_5883,N_5834);
nor U6735 (N_6735,N_5573,N_5164);
nand U6736 (N_6736,N_5596,N_5570);
nor U6737 (N_6737,N_5661,N_5950);
xnor U6738 (N_6738,N_5353,N_5354);
or U6739 (N_6739,N_5173,N_5178);
xnor U6740 (N_6740,N_5056,N_5377);
nand U6741 (N_6741,N_5036,N_5284);
or U6742 (N_6742,N_5723,N_5990);
and U6743 (N_6743,N_5413,N_5389);
nor U6744 (N_6744,N_5762,N_5808);
or U6745 (N_6745,N_5379,N_5292);
xnor U6746 (N_6746,N_5786,N_5000);
or U6747 (N_6747,N_5572,N_5492);
and U6748 (N_6748,N_5001,N_5532);
or U6749 (N_6749,N_5960,N_5841);
nand U6750 (N_6750,N_5464,N_5728);
or U6751 (N_6751,N_5700,N_5268);
nor U6752 (N_6752,N_5270,N_5319);
xor U6753 (N_6753,N_5627,N_5290);
or U6754 (N_6754,N_5127,N_5517);
xor U6755 (N_6755,N_5149,N_5479);
or U6756 (N_6756,N_5285,N_5641);
nand U6757 (N_6757,N_5662,N_5809);
nand U6758 (N_6758,N_5845,N_5688);
and U6759 (N_6759,N_5870,N_5700);
nand U6760 (N_6760,N_5946,N_5466);
or U6761 (N_6761,N_5877,N_5968);
and U6762 (N_6762,N_5100,N_5350);
xor U6763 (N_6763,N_5844,N_5062);
and U6764 (N_6764,N_5916,N_5544);
and U6765 (N_6765,N_5425,N_5426);
nand U6766 (N_6766,N_5246,N_5912);
nand U6767 (N_6767,N_5008,N_5069);
and U6768 (N_6768,N_5222,N_5386);
and U6769 (N_6769,N_5051,N_5464);
nor U6770 (N_6770,N_5355,N_5351);
xor U6771 (N_6771,N_5924,N_5221);
or U6772 (N_6772,N_5841,N_5658);
nand U6773 (N_6773,N_5569,N_5183);
and U6774 (N_6774,N_5197,N_5547);
nand U6775 (N_6775,N_5515,N_5648);
or U6776 (N_6776,N_5052,N_5730);
or U6777 (N_6777,N_5562,N_5421);
and U6778 (N_6778,N_5594,N_5829);
xor U6779 (N_6779,N_5309,N_5709);
xnor U6780 (N_6780,N_5973,N_5109);
xnor U6781 (N_6781,N_5632,N_5223);
or U6782 (N_6782,N_5993,N_5853);
and U6783 (N_6783,N_5351,N_5838);
or U6784 (N_6784,N_5080,N_5493);
nor U6785 (N_6785,N_5508,N_5292);
or U6786 (N_6786,N_5758,N_5129);
and U6787 (N_6787,N_5683,N_5621);
nand U6788 (N_6788,N_5618,N_5428);
nand U6789 (N_6789,N_5073,N_5124);
and U6790 (N_6790,N_5382,N_5877);
or U6791 (N_6791,N_5188,N_5457);
nand U6792 (N_6792,N_5104,N_5129);
nor U6793 (N_6793,N_5535,N_5558);
nor U6794 (N_6794,N_5215,N_5635);
and U6795 (N_6795,N_5959,N_5520);
or U6796 (N_6796,N_5619,N_5375);
or U6797 (N_6797,N_5552,N_5489);
nor U6798 (N_6798,N_5669,N_5754);
or U6799 (N_6799,N_5840,N_5102);
nand U6800 (N_6800,N_5203,N_5524);
or U6801 (N_6801,N_5055,N_5089);
and U6802 (N_6802,N_5304,N_5058);
and U6803 (N_6803,N_5083,N_5160);
xnor U6804 (N_6804,N_5945,N_5624);
xnor U6805 (N_6805,N_5928,N_5640);
xnor U6806 (N_6806,N_5823,N_5129);
xnor U6807 (N_6807,N_5919,N_5199);
nand U6808 (N_6808,N_5636,N_5135);
or U6809 (N_6809,N_5663,N_5093);
xnor U6810 (N_6810,N_5198,N_5089);
and U6811 (N_6811,N_5872,N_5097);
or U6812 (N_6812,N_5580,N_5270);
nand U6813 (N_6813,N_5141,N_5036);
and U6814 (N_6814,N_5801,N_5303);
nor U6815 (N_6815,N_5304,N_5300);
or U6816 (N_6816,N_5917,N_5726);
or U6817 (N_6817,N_5102,N_5948);
or U6818 (N_6818,N_5240,N_5858);
xnor U6819 (N_6819,N_5469,N_5830);
nand U6820 (N_6820,N_5059,N_5691);
and U6821 (N_6821,N_5478,N_5070);
xor U6822 (N_6822,N_5094,N_5433);
xnor U6823 (N_6823,N_5515,N_5725);
and U6824 (N_6824,N_5632,N_5536);
and U6825 (N_6825,N_5560,N_5815);
nand U6826 (N_6826,N_5513,N_5316);
nand U6827 (N_6827,N_5875,N_5998);
nor U6828 (N_6828,N_5104,N_5597);
and U6829 (N_6829,N_5290,N_5680);
nor U6830 (N_6830,N_5044,N_5046);
nor U6831 (N_6831,N_5393,N_5565);
and U6832 (N_6832,N_5489,N_5014);
and U6833 (N_6833,N_5976,N_5670);
nor U6834 (N_6834,N_5199,N_5742);
and U6835 (N_6835,N_5631,N_5105);
and U6836 (N_6836,N_5609,N_5498);
or U6837 (N_6837,N_5955,N_5995);
and U6838 (N_6838,N_5680,N_5389);
nand U6839 (N_6839,N_5466,N_5857);
nand U6840 (N_6840,N_5692,N_5400);
or U6841 (N_6841,N_5064,N_5832);
and U6842 (N_6842,N_5364,N_5263);
and U6843 (N_6843,N_5735,N_5328);
nor U6844 (N_6844,N_5886,N_5050);
xnor U6845 (N_6845,N_5733,N_5304);
nand U6846 (N_6846,N_5208,N_5004);
and U6847 (N_6847,N_5000,N_5883);
xnor U6848 (N_6848,N_5639,N_5951);
and U6849 (N_6849,N_5622,N_5104);
or U6850 (N_6850,N_5756,N_5057);
and U6851 (N_6851,N_5045,N_5671);
xor U6852 (N_6852,N_5042,N_5300);
nor U6853 (N_6853,N_5543,N_5360);
and U6854 (N_6854,N_5611,N_5950);
and U6855 (N_6855,N_5782,N_5175);
xor U6856 (N_6856,N_5513,N_5661);
xor U6857 (N_6857,N_5154,N_5691);
and U6858 (N_6858,N_5373,N_5863);
nor U6859 (N_6859,N_5038,N_5744);
nand U6860 (N_6860,N_5047,N_5679);
nand U6861 (N_6861,N_5418,N_5494);
nand U6862 (N_6862,N_5728,N_5941);
or U6863 (N_6863,N_5898,N_5493);
nor U6864 (N_6864,N_5052,N_5193);
or U6865 (N_6865,N_5406,N_5256);
xnor U6866 (N_6866,N_5684,N_5581);
or U6867 (N_6867,N_5484,N_5027);
nor U6868 (N_6868,N_5417,N_5206);
or U6869 (N_6869,N_5225,N_5503);
nor U6870 (N_6870,N_5645,N_5523);
nand U6871 (N_6871,N_5748,N_5889);
or U6872 (N_6872,N_5060,N_5509);
and U6873 (N_6873,N_5541,N_5122);
xor U6874 (N_6874,N_5553,N_5291);
and U6875 (N_6875,N_5229,N_5128);
xor U6876 (N_6876,N_5635,N_5437);
or U6877 (N_6877,N_5064,N_5186);
nor U6878 (N_6878,N_5537,N_5403);
nor U6879 (N_6879,N_5303,N_5474);
and U6880 (N_6880,N_5441,N_5744);
nor U6881 (N_6881,N_5918,N_5654);
nor U6882 (N_6882,N_5427,N_5271);
nor U6883 (N_6883,N_5513,N_5028);
nor U6884 (N_6884,N_5390,N_5039);
or U6885 (N_6885,N_5805,N_5302);
nor U6886 (N_6886,N_5318,N_5344);
and U6887 (N_6887,N_5402,N_5637);
and U6888 (N_6888,N_5764,N_5060);
xnor U6889 (N_6889,N_5192,N_5313);
nor U6890 (N_6890,N_5410,N_5175);
and U6891 (N_6891,N_5792,N_5036);
nor U6892 (N_6892,N_5333,N_5362);
or U6893 (N_6893,N_5729,N_5834);
and U6894 (N_6894,N_5489,N_5288);
and U6895 (N_6895,N_5670,N_5416);
and U6896 (N_6896,N_5153,N_5726);
or U6897 (N_6897,N_5109,N_5625);
nor U6898 (N_6898,N_5980,N_5484);
xnor U6899 (N_6899,N_5828,N_5627);
nor U6900 (N_6900,N_5764,N_5080);
nand U6901 (N_6901,N_5927,N_5928);
nand U6902 (N_6902,N_5310,N_5896);
nand U6903 (N_6903,N_5991,N_5120);
nor U6904 (N_6904,N_5926,N_5035);
and U6905 (N_6905,N_5859,N_5447);
or U6906 (N_6906,N_5117,N_5969);
and U6907 (N_6907,N_5258,N_5243);
nand U6908 (N_6908,N_5315,N_5049);
nand U6909 (N_6909,N_5921,N_5160);
nand U6910 (N_6910,N_5587,N_5109);
or U6911 (N_6911,N_5296,N_5286);
and U6912 (N_6912,N_5530,N_5952);
and U6913 (N_6913,N_5660,N_5208);
nor U6914 (N_6914,N_5505,N_5917);
xor U6915 (N_6915,N_5769,N_5050);
xor U6916 (N_6916,N_5343,N_5003);
or U6917 (N_6917,N_5533,N_5907);
or U6918 (N_6918,N_5860,N_5337);
xor U6919 (N_6919,N_5167,N_5417);
and U6920 (N_6920,N_5865,N_5207);
or U6921 (N_6921,N_5478,N_5746);
nor U6922 (N_6922,N_5274,N_5948);
or U6923 (N_6923,N_5093,N_5320);
or U6924 (N_6924,N_5087,N_5154);
nand U6925 (N_6925,N_5157,N_5781);
nor U6926 (N_6926,N_5817,N_5559);
nand U6927 (N_6927,N_5684,N_5750);
or U6928 (N_6928,N_5261,N_5091);
nor U6929 (N_6929,N_5627,N_5651);
or U6930 (N_6930,N_5143,N_5090);
xnor U6931 (N_6931,N_5976,N_5838);
nor U6932 (N_6932,N_5602,N_5257);
nand U6933 (N_6933,N_5311,N_5836);
and U6934 (N_6934,N_5790,N_5616);
nor U6935 (N_6935,N_5564,N_5617);
or U6936 (N_6936,N_5801,N_5044);
or U6937 (N_6937,N_5944,N_5937);
nand U6938 (N_6938,N_5158,N_5150);
or U6939 (N_6939,N_5843,N_5299);
xnor U6940 (N_6940,N_5094,N_5054);
nor U6941 (N_6941,N_5175,N_5205);
and U6942 (N_6942,N_5301,N_5790);
xor U6943 (N_6943,N_5235,N_5396);
xor U6944 (N_6944,N_5521,N_5164);
nor U6945 (N_6945,N_5544,N_5510);
nor U6946 (N_6946,N_5743,N_5459);
nor U6947 (N_6947,N_5859,N_5956);
or U6948 (N_6948,N_5624,N_5507);
and U6949 (N_6949,N_5267,N_5134);
and U6950 (N_6950,N_5107,N_5164);
xnor U6951 (N_6951,N_5706,N_5287);
and U6952 (N_6952,N_5972,N_5184);
and U6953 (N_6953,N_5416,N_5346);
and U6954 (N_6954,N_5778,N_5765);
xor U6955 (N_6955,N_5684,N_5628);
nand U6956 (N_6956,N_5757,N_5702);
or U6957 (N_6957,N_5216,N_5793);
and U6958 (N_6958,N_5524,N_5491);
and U6959 (N_6959,N_5418,N_5261);
or U6960 (N_6960,N_5151,N_5192);
or U6961 (N_6961,N_5303,N_5554);
nor U6962 (N_6962,N_5299,N_5704);
nor U6963 (N_6963,N_5964,N_5446);
and U6964 (N_6964,N_5617,N_5681);
or U6965 (N_6965,N_5297,N_5920);
or U6966 (N_6966,N_5388,N_5537);
nand U6967 (N_6967,N_5904,N_5005);
or U6968 (N_6968,N_5179,N_5158);
and U6969 (N_6969,N_5171,N_5108);
or U6970 (N_6970,N_5174,N_5997);
xor U6971 (N_6971,N_5337,N_5018);
and U6972 (N_6972,N_5893,N_5804);
and U6973 (N_6973,N_5089,N_5929);
nor U6974 (N_6974,N_5490,N_5286);
nor U6975 (N_6975,N_5864,N_5235);
xnor U6976 (N_6976,N_5792,N_5356);
or U6977 (N_6977,N_5281,N_5392);
and U6978 (N_6978,N_5868,N_5353);
nor U6979 (N_6979,N_5394,N_5962);
or U6980 (N_6980,N_5701,N_5540);
nor U6981 (N_6981,N_5768,N_5118);
and U6982 (N_6982,N_5707,N_5920);
and U6983 (N_6983,N_5674,N_5703);
and U6984 (N_6984,N_5072,N_5218);
or U6985 (N_6985,N_5145,N_5369);
nand U6986 (N_6986,N_5738,N_5496);
and U6987 (N_6987,N_5301,N_5902);
nand U6988 (N_6988,N_5708,N_5478);
nor U6989 (N_6989,N_5970,N_5402);
nand U6990 (N_6990,N_5203,N_5377);
and U6991 (N_6991,N_5933,N_5911);
and U6992 (N_6992,N_5735,N_5272);
xor U6993 (N_6993,N_5766,N_5210);
or U6994 (N_6994,N_5532,N_5048);
nor U6995 (N_6995,N_5663,N_5139);
nand U6996 (N_6996,N_5185,N_5246);
nand U6997 (N_6997,N_5741,N_5705);
or U6998 (N_6998,N_5220,N_5514);
or U6999 (N_6999,N_5966,N_5923);
nand U7000 (N_7000,N_6557,N_6824);
or U7001 (N_7001,N_6599,N_6860);
nor U7002 (N_7002,N_6590,N_6332);
nor U7003 (N_7003,N_6565,N_6719);
nand U7004 (N_7004,N_6456,N_6201);
nand U7005 (N_7005,N_6002,N_6229);
and U7006 (N_7006,N_6180,N_6173);
xor U7007 (N_7007,N_6676,N_6512);
nand U7008 (N_7008,N_6667,N_6145);
nor U7009 (N_7009,N_6837,N_6602);
nor U7010 (N_7010,N_6699,N_6897);
nor U7011 (N_7011,N_6049,N_6207);
xor U7012 (N_7012,N_6464,N_6490);
xnor U7013 (N_7013,N_6252,N_6521);
xnor U7014 (N_7014,N_6193,N_6756);
and U7015 (N_7015,N_6064,N_6636);
or U7016 (N_7016,N_6781,N_6955);
or U7017 (N_7017,N_6610,N_6624);
and U7018 (N_7018,N_6966,N_6698);
xor U7019 (N_7019,N_6838,N_6903);
xor U7020 (N_7020,N_6678,N_6627);
or U7021 (N_7021,N_6928,N_6352);
xnor U7022 (N_7022,N_6005,N_6017);
nand U7023 (N_7023,N_6471,N_6329);
xnor U7024 (N_7024,N_6254,N_6309);
nand U7025 (N_7025,N_6162,N_6104);
nand U7026 (N_7026,N_6295,N_6703);
or U7027 (N_7027,N_6028,N_6444);
nand U7028 (N_7028,N_6062,N_6405);
or U7029 (N_7029,N_6333,N_6109);
nor U7030 (N_7030,N_6630,N_6688);
xor U7031 (N_7031,N_6281,N_6510);
or U7032 (N_7032,N_6076,N_6712);
and U7033 (N_7033,N_6604,N_6169);
xnor U7034 (N_7034,N_6043,N_6215);
nand U7035 (N_7035,N_6312,N_6155);
or U7036 (N_7036,N_6905,N_6972);
and U7037 (N_7037,N_6096,N_6434);
nand U7038 (N_7038,N_6470,N_6337);
xor U7039 (N_7039,N_6407,N_6122);
nor U7040 (N_7040,N_6716,N_6568);
or U7041 (N_7041,N_6596,N_6642);
nor U7042 (N_7042,N_6025,N_6419);
xnor U7043 (N_7043,N_6694,N_6945);
nor U7044 (N_7044,N_6219,N_6858);
and U7045 (N_7045,N_6098,N_6878);
or U7046 (N_7046,N_6266,N_6527);
nand U7047 (N_7047,N_6030,N_6450);
nand U7048 (N_7048,N_6168,N_6090);
and U7049 (N_7049,N_6531,N_6754);
xor U7050 (N_7050,N_6526,N_6035);
and U7051 (N_7051,N_6992,N_6567);
nand U7052 (N_7052,N_6745,N_6555);
nand U7053 (N_7053,N_6755,N_6380);
or U7054 (N_7054,N_6544,N_6425);
nor U7055 (N_7055,N_6112,N_6317);
or U7056 (N_7056,N_6374,N_6366);
nand U7057 (N_7057,N_6165,N_6186);
xnor U7058 (N_7058,N_6908,N_6232);
and U7059 (N_7059,N_6718,N_6282);
nand U7060 (N_7060,N_6664,N_6074);
xnor U7061 (N_7061,N_6340,N_6351);
nor U7062 (N_7062,N_6999,N_6902);
nor U7063 (N_7063,N_6396,N_6223);
or U7064 (N_7064,N_6154,N_6733);
and U7065 (N_7065,N_6543,N_6750);
xnor U7066 (N_7066,N_6373,N_6068);
nand U7067 (N_7067,N_6491,N_6650);
nand U7068 (N_7068,N_6272,N_6323);
and U7069 (N_7069,N_6259,N_6801);
or U7070 (N_7070,N_6575,N_6150);
xor U7071 (N_7071,N_6131,N_6939);
and U7072 (N_7072,N_6845,N_6654);
or U7073 (N_7073,N_6263,N_6420);
and U7074 (N_7074,N_6560,N_6920);
nand U7075 (N_7075,N_6623,N_6414);
or U7076 (N_7076,N_6012,N_6832);
nand U7077 (N_7077,N_6658,N_6742);
and U7078 (N_7078,N_6107,N_6707);
and U7079 (N_7079,N_6585,N_6302);
or U7080 (N_7080,N_6917,N_6923);
and U7081 (N_7081,N_6632,N_6629);
nor U7082 (N_7082,N_6181,N_6504);
or U7083 (N_7083,N_6408,N_6690);
nand U7084 (N_7084,N_6486,N_6620);
xnor U7085 (N_7085,N_6887,N_6569);
nand U7086 (N_7086,N_6645,N_6951);
nor U7087 (N_7087,N_6370,N_6976);
or U7088 (N_7088,N_6392,N_6727);
or U7089 (N_7089,N_6182,N_6192);
nand U7090 (N_7090,N_6124,N_6741);
or U7091 (N_7091,N_6533,N_6494);
xnor U7092 (N_7092,N_6705,N_6037);
or U7093 (N_7093,N_6589,N_6009);
xnor U7094 (N_7094,N_6156,N_6102);
nor U7095 (N_7095,N_6812,N_6199);
or U7096 (N_7096,N_6835,N_6278);
nor U7097 (N_7097,N_6236,N_6379);
nand U7098 (N_7098,N_6572,N_6672);
and U7099 (N_7099,N_6586,N_6296);
nand U7100 (N_7100,N_6482,N_6360);
xor U7101 (N_7101,N_6428,N_6031);
nand U7102 (N_7102,N_6840,N_6611);
nor U7103 (N_7103,N_6844,N_6211);
nor U7104 (N_7104,N_6775,N_6046);
or U7105 (N_7105,N_6178,N_6409);
or U7106 (N_7106,N_6591,N_6984);
xnor U7107 (N_7107,N_6398,N_6113);
xor U7108 (N_7108,N_6865,N_6873);
nand U7109 (N_7109,N_6200,N_6634);
and U7110 (N_7110,N_6481,N_6447);
nand U7111 (N_7111,N_6530,N_6465);
xnor U7112 (N_7112,N_6209,N_6509);
nand U7113 (N_7113,N_6904,N_6000);
xor U7114 (N_7114,N_6751,N_6054);
or U7115 (N_7115,N_6077,N_6190);
and U7116 (N_7116,N_6338,N_6391);
nand U7117 (N_7117,N_6545,N_6042);
nand U7118 (N_7118,N_6790,N_6235);
xor U7119 (N_7119,N_6950,N_6144);
nand U7120 (N_7120,N_6082,N_6948);
or U7121 (N_7121,N_6711,N_6151);
nor U7122 (N_7122,N_6542,N_6683);
nor U7123 (N_7123,N_6652,N_6831);
and U7124 (N_7124,N_6899,N_6176);
xor U7125 (N_7125,N_6541,N_6141);
or U7126 (N_7126,N_6301,N_6417);
and U7127 (N_7127,N_6324,N_6969);
nand U7128 (N_7128,N_6679,N_6639);
xor U7129 (N_7129,N_6217,N_6292);
xor U7130 (N_7130,N_6286,N_6411);
or U7131 (N_7131,N_6003,N_6594);
xor U7132 (N_7132,N_6856,N_6306);
nand U7133 (N_7133,N_6094,N_6888);
or U7134 (N_7134,N_6095,N_6539);
xor U7135 (N_7135,N_6498,N_6101);
and U7136 (N_7136,N_6558,N_6519);
nand U7137 (N_7137,N_6427,N_6033);
nand U7138 (N_7138,N_6331,N_6534);
or U7139 (N_7139,N_6435,N_6262);
or U7140 (N_7140,N_6965,N_6140);
nand U7141 (N_7141,N_6912,N_6280);
nor U7142 (N_7142,N_6105,N_6906);
and U7143 (N_7143,N_6473,N_6884);
nor U7144 (N_7144,N_6053,N_6422);
xnor U7145 (N_7145,N_6163,N_6597);
nand U7146 (N_7146,N_6161,N_6593);
and U7147 (N_7147,N_6746,N_6648);
or U7148 (N_7148,N_6430,N_6172);
or U7149 (N_7149,N_6401,N_6174);
or U7150 (N_7150,N_6327,N_6857);
nand U7151 (N_7151,N_6460,N_6925);
xor U7152 (N_7152,N_6210,N_6919);
nor U7153 (N_7153,N_6039,N_6100);
nand U7154 (N_7154,N_6245,N_6655);
xnor U7155 (N_7155,N_6106,N_6686);
and U7156 (N_7156,N_6298,N_6792);
and U7157 (N_7157,N_6023,N_6047);
xor U7158 (N_7158,N_6212,N_6365);
xor U7159 (N_7159,N_6221,N_6868);
nand U7160 (N_7160,N_6111,N_6191);
xor U7161 (N_7161,N_6063,N_6115);
nor U7162 (N_7162,N_6890,N_6977);
xor U7163 (N_7163,N_6294,N_6179);
or U7164 (N_7164,N_6454,N_6684);
nand U7165 (N_7165,N_6717,N_6852);
and U7166 (N_7166,N_6901,N_6830);
and U7167 (N_7167,N_6795,N_6345);
nor U7168 (N_7168,N_6413,N_6319);
nor U7169 (N_7169,N_6749,N_6126);
or U7170 (N_7170,N_6866,N_6721);
or U7171 (N_7171,N_6116,N_6458);
and U7172 (N_7172,N_6603,N_6404);
or U7173 (N_7173,N_6135,N_6320);
and U7174 (N_7174,N_6022,N_6618);
or U7175 (N_7175,N_6070,N_6438);
and U7176 (N_7176,N_6861,N_6522);
xor U7177 (N_7177,N_6097,N_6314);
and U7178 (N_7178,N_6477,N_6429);
and U7179 (N_7179,N_6635,N_6363);
xnor U7180 (N_7180,N_6723,N_6441);
nor U7181 (N_7181,N_6501,N_6796);
and U7182 (N_7182,N_6574,N_6990);
and U7183 (N_7183,N_6625,N_6706);
nor U7184 (N_7184,N_6249,N_6788);
xor U7185 (N_7185,N_6388,N_6783);
nor U7186 (N_7186,N_6768,N_6308);
nand U7187 (N_7187,N_6961,N_6239);
nor U7188 (N_7188,N_6930,N_6549);
and U7189 (N_7189,N_6440,N_6159);
xor U7190 (N_7190,N_6685,N_6728);
nand U7191 (N_7191,N_6382,N_6934);
xnor U7192 (N_7192,N_6536,N_6563);
nor U7193 (N_7193,N_6052,N_6216);
nand U7194 (N_7194,N_6540,N_6318);
and U7195 (N_7195,N_6394,N_6621);
nand U7196 (N_7196,N_6980,N_6493);
xnor U7197 (N_7197,N_6137,N_6968);
xnor U7198 (N_7198,N_6595,N_6782);
nand U7199 (N_7199,N_6244,N_6007);
or U7200 (N_7200,N_6784,N_6433);
nand U7201 (N_7201,N_6128,N_6778);
and U7202 (N_7202,N_6187,N_6631);
nand U7203 (N_7203,N_6061,N_6571);
or U7204 (N_7204,N_6810,N_6626);
xnor U7205 (N_7205,N_6547,N_6358);
or U7206 (N_7206,N_6475,N_6213);
xor U7207 (N_7207,N_6316,N_6663);
nor U7208 (N_7208,N_6643,N_6987);
nand U7209 (N_7209,N_6204,N_6171);
nand U7210 (N_7210,N_6896,N_6462);
or U7211 (N_7211,N_6825,N_6771);
and U7212 (N_7212,N_6507,N_6395);
xor U7213 (N_7213,N_6850,N_6436);
xnor U7214 (N_7214,N_6400,N_6764);
or U7215 (N_7215,N_6633,N_6581);
nand U7216 (N_7216,N_6160,N_6696);
and U7217 (N_7217,N_6989,N_6828);
and U7218 (N_7218,N_6864,N_6709);
nand U7219 (N_7219,N_6303,N_6225);
or U7220 (N_7220,N_6587,N_6132);
and U7221 (N_7221,N_6015,N_6451);
or U7222 (N_7222,N_6787,N_6253);
xor U7223 (N_7223,N_6666,N_6378);
or U7224 (N_7224,N_6867,N_6524);
or U7225 (N_7225,N_6001,N_6562);
or U7226 (N_7226,N_6148,N_6243);
and U7227 (N_7227,N_6900,N_6234);
xnor U7228 (N_7228,N_6087,N_6321);
or U7229 (N_7229,N_6582,N_6670);
xnor U7230 (N_7230,N_6995,N_6882);
xnor U7231 (N_7231,N_6779,N_6157);
nor U7232 (N_7232,N_6819,N_6886);
and U7233 (N_7233,N_6883,N_6843);
xnor U7234 (N_7234,N_6431,N_6993);
nand U7235 (N_7235,N_6459,N_6578);
and U7236 (N_7236,N_6681,N_6637);
and U7237 (N_7237,N_6326,N_6393);
or U7238 (N_7238,N_6982,N_6300);
xor U7239 (N_7239,N_6067,N_6305);
nor U7240 (N_7240,N_6285,N_6220);
nor U7241 (N_7241,N_6827,N_6083);
and U7242 (N_7242,N_6389,N_6255);
nor U7243 (N_7243,N_6601,N_6752);
nand U7244 (N_7244,N_6123,N_6013);
and U7245 (N_7245,N_6099,N_6335);
nand U7246 (N_7246,N_6876,N_6416);
nand U7247 (N_7247,N_6836,N_6091);
nor U7248 (N_7248,N_6598,N_6986);
nor U7249 (N_7249,N_6088,N_6988);
or U7250 (N_7250,N_6791,N_6556);
nor U7251 (N_7251,N_6189,N_6461);
and U7252 (N_7252,N_6240,N_6975);
nor U7253 (N_7253,N_6250,N_6277);
and U7254 (N_7254,N_6793,N_6849);
or U7255 (N_7255,N_6763,N_6103);
and U7256 (N_7256,N_6138,N_6364);
and U7257 (N_7257,N_6677,N_6963);
nor U7258 (N_7258,N_6289,N_6268);
and U7259 (N_7259,N_6566,N_6889);
or U7260 (N_7260,N_6962,N_6503);
xor U7261 (N_7261,N_6820,N_6251);
or U7262 (N_7262,N_6767,N_6120);
nand U7263 (N_7263,N_6343,N_6817);
or U7264 (N_7264,N_6072,N_6660);
or U7265 (N_7265,N_6084,N_6348);
xor U7266 (N_7266,N_6092,N_6937);
nand U7267 (N_7267,N_6121,N_6553);
and U7268 (N_7268,N_6080,N_6938);
xor U7269 (N_7269,N_6693,N_6862);
and U7270 (N_7270,N_6474,N_6484);
nand U7271 (N_7271,N_6695,N_6387);
and U7272 (N_7272,N_6377,N_6915);
or U7273 (N_7273,N_6818,N_6073);
nor U7274 (N_7274,N_6761,N_6117);
or U7275 (N_7275,N_6500,N_6985);
xnor U7276 (N_7276,N_6615,N_6368);
or U7277 (N_7277,N_6922,N_6349);
and U7278 (N_7278,N_6048,N_6375);
or U7279 (N_7279,N_6342,N_6227);
nor U7280 (N_7280,N_6502,N_6508);
xor U7281 (N_7281,N_6584,N_6933);
xnor U7282 (N_7282,N_6619,N_6385);
and U7283 (N_7283,N_6926,N_6846);
and U7284 (N_7284,N_6580,N_6233);
or U7285 (N_7285,N_6735,N_6789);
xor U7286 (N_7286,N_6537,N_6564);
xor U7287 (N_7287,N_6469,N_6954);
xor U7288 (N_7288,N_6075,N_6515);
nor U7289 (N_7289,N_6164,N_6525);
xor U7290 (N_7290,N_6757,N_6806);
nor U7291 (N_7291,N_6758,N_6994);
and U7292 (N_7292,N_6523,N_6224);
xor U7293 (N_7293,N_6269,N_6260);
and U7294 (N_7294,N_6410,N_6026);
nand U7295 (N_7295,N_6725,N_6576);
and U7296 (N_7296,N_6439,N_6871);
or U7297 (N_7297,N_6893,N_6202);
nor U7298 (N_7298,N_6513,N_6967);
or U7299 (N_7299,N_6205,N_6143);
or U7300 (N_7300,N_6559,N_6492);
and U7301 (N_7301,N_6606,N_6038);
xor U7302 (N_7302,N_6907,N_6946);
nand U7303 (N_7303,N_6467,N_6600);
xnor U7304 (N_7304,N_6086,N_6264);
and U7305 (N_7305,N_6609,N_6814);
nor U7306 (N_7306,N_6853,N_6715);
and U7307 (N_7307,N_6010,N_6518);
and U7308 (N_7308,N_6724,N_6894);
and U7309 (N_7309,N_6455,N_6668);
nand U7310 (N_7310,N_6403,N_6241);
and U7311 (N_7311,N_6798,N_6270);
xnor U7312 (N_7312,N_6479,N_6271);
nor U7313 (N_7313,N_6029,N_6821);
xnor U7314 (N_7314,N_6386,N_6532);
or U7315 (N_7315,N_6996,N_6855);
xnor U7316 (N_7316,N_6307,N_6371);
nand U7317 (N_7317,N_6057,N_6628);
xnor U7318 (N_7318,N_6472,N_6583);
nand U7319 (N_7319,N_6823,N_6800);
and U7320 (N_7320,N_6605,N_6021);
or U7321 (N_7321,N_6018,N_6811);
nand U7322 (N_7322,N_6517,N_6446);
and U7323 (N_7323,N_6649,N_6208);
nor U7324 (N_7324,N_6376,N_6813);
or U7325 (N_7325,N_6287,N_6981);
xnor U7326 (N_7326,N_6734,N_6974);
and U7327 (N_7327,N_6284,N_6740);
and U7328 (N_7328,N_6739,N_6027);
xor U7329 (N_7329,N_6288,N_6432);
or U7330 (N_7330,N_6125,N_6108);
xnor U7331 (N_7331,N_6701,N_6669);
xnor U7332 (N_7332,N_6998,N_6311);
nor U7333 (N_7333,N_6448,N_6949);
and U7334 (N_7334,N_6879,N_6874);
or U7335 (N_7335,N_6913,N_6310);
nand U7336 (N_7336,N_6765,N_6265);
nor U7337 (N_7337,N_6040,N_6956);
nand U7338 (N_7338,N_6384,N_6177);
nor U7339 (N_7339,N_6274,N_6708);
nand U7340 (N_7340,N_6118,N_6799);
nor U7341 (N_7341,N_6110,N_6055);
nand U7342 (N_7342,N_6426,N_6423);
nand U7343 (N_7343,N_6916,N_6032);
nand U7344 (N_7344,N_6129,N_6056);
xnor U7345 (N_7345,N_6704,N_6644);
nor U7346 (N_7346,N_6198,N_6194);
xnor U7347 (N_7347,N_6673,N_6834);
nor U7348 (N_7348,N_6918,N_6592);
nand U7349 (N_7349,N_6561,N_6226);
and U7350 (N_7350,N_6891,N_6315);
nor U7351 (N_7351,N_6952,N_6929);
or U7352 (N_7352,N_6065,N_6114);
and U7353 (N_7353,N_6346,N_6877);
nand U7354 (N_7354,N_6641,N_6020);
or U7355 (N_7355,N_6892,N_6804);
or U7356 (N_7356,N_6506,N_6702);
nor U7357 (N_7357,N_6059,N_6869);
or U7358 (N_7358,N_6196,N_6230);
or U7359 (N_7359,N_6737,N_6738);
nand U7360 (N_7360,N_6661,N_6924);
and U7361 (N_7361,N_6158,N_6927);
xor U7362 (N_7362,N_6730,N_6214);
and U7363 (N_7363,N_6722,N_6466);
nor U7364 (N_7364,N_6570,N_6895);
xnor U7365 (N_7365,N_6726,N_6483);
nand U7366 (N_7366,N_6554,N_6659);
xor U7367 (N_7367,N_6079,N_6489);
nand U7368 (N_7368,N_6700,N_6197);
and U7369 (N_7369,N_6942,N_6089);
nor U7370 (N_7370,N_6044,N_6297);
nand U7371 (N_7371,N_6833,N_6069);
nor U7372 (N_7372,N_6538,N_6514);
xor U7373 (N_7373,N_6816,N_6499);
nand U7374 (N_7374,N_6347,N_6185);
xor U7375 (N_7375,N_6780,N_6119);
nand U7376 (N_7376,N_6146,N_6206);
nand U7377 (N_7377,N_6516,N_6675);
xor U7378 (N_7378,N_6944,N_6361);
or U7379 (N_7379,N_6914,N_6293);
nor U7380 (N_7380,N_6747,N_6004);
or U7381 (N_7381,N_6851,N_6607);
xnor U7382 (N_7382,N_6957,N_6136);
or U7383 (N_7383,N_6328,N_6267);
nand U7384 (N_7384,N_6369,N_6355);
and U7385 (N_7385,N_6935,N_6203);
xnor U7386 (N_7386,N_6662,N_6881);
nor U7387 (N_7387,N_6979,N_6273);
nor U7388 (N_7388,N_6983,N_6766);
and U7389 (N_7389,N_6991,N_6714);
xnor U7390 (N_7390,N_6931,N_6797);
nor U7391 (N_7391,N_6520,N_6680);
xor U7392 (N_7392,N_6078,N_6008);
or U7393 (N_7393,N_6006,N_6732);
xnor U7394 (N_7394,N_6424,N_6697);
nor U7395 (N_7395,N_6943,N_6362);
nor U7396 (N_7396,N_6959,N_6256);
and U7397 (N_7397,N_6153,N_6166);
xnor U7398 (N_7398,N_6147,N_6222);
and U7399 (N_7399,N_6152,N_6184);
nor U7400 (N_7400,N_6195,N_6653);
and U7401 (N_7401,N_6910,N_6248);
xnor U7402 (N_7402,N_6535,N_6936);
nor U7403 (N_7403,N_6638,N_6066);
nor U7404 (N_7404,N_6353,N_6276);
or U7405 (N_7405,N_6612,N_6505);
nor U7406 (N_7406,N_6133,N_6183);
or U7407 (N_7407,N_6743,N_6336);
or U7408 (N_7408,N_6218,N_6445);
nor U7409 (N_7409,N_6339,N_6231);
xor U7410 (N_7410,N_6016,N_6579);
xor U7411 (N_7411,N_6546,N_6748);
xor U7412 (N_7412,N_6729,N_6050);
or U7413 (N_7413,N_6847,N_6552);
nand U7414 (N_7414,N_6720,N_6011);
nor U7415 (N_7415,N_6651,N_6051);
nor U7416 (N_7416,N_6870,N_6188);
or U7417 (N_7417,N_6608,N_6372);
or U7418 (N_7418,N_6776,N_6665);
nand U7419 (N_7419,N_6921,N_6247);
xnor U7420 (N_7420,N_6909,N_6495);
and U7421 (N_7421,N_6859,N_6970);
and U7422 (N_7422,N_6334,N_6682);
nand U7423 (N_7423,N_6863,N_6794);
or U7424 (N_7424,N_6497,N_6397);
or U7425 (N_7425,N_6304,N_6770);
nand U7426 (N_7426,N_6657,N_6744);
nor U7427 (N_7427,N_6325,N_6826);
and U7428 (N_7428,N_6953,N_6085);
xnor U7429 (N_7429,N_6528,N_6656);
xnor U7430 (N_7430,N_6885,N_6774);
xnor U7431 (N_7431,N_6753,N_6736);
and U7432 (N_7432,N_6291,N_6551);
nor U7433 (N_7433,N_6468,N_6449);
nand U7434 (N_7434,N_6691,N_6452);
nor U7435 (N_7435,N_6261,N_6399);
xor U7436 (N_7436,N_6367,N_6875);
xnor U7437 (N_7437,N_6854,N_6588);
nor U7438 (N_7438,N_6805,N_6093);
and U7439 (N_7439,N_6689,N_6773);
xnor U7440 (N_7440,N_6390,N_6496);
or U7441 (N_7441,N_6674,N_6488);
nor U7442 (N_7442,N_6616,N_6759);
or U7443 (N_7443,N_6170,N_6617);
nand U7444 (N_7444,N_6383,N_6457);
and U7445 (N_7445,N_6071,N_6228);
xnor U7446 (N_7446,N_6573,N_6283);
and U7447 (N_7447,N_6443,N_6036);
or U7448 (N_7448,N_6418,N_6622);
nor U7449 (N_7449,N_6341,N_6613);
and U7450 (N_7450,N_6808,N_6299);
or U7451 (N_7451,N_6415,N_6713);
or U7452 (N_7452,N_6354,N_6257);
nor U7453 (N_7453,N_6971,N_6421);
xnor U7454 (N_7454,N_6550,N_6898);
nand U7455 (N_7455,N_6731,N_6548);
xnor U7456 (N_7456,N_6973,N_6019);
and U7457 (N_7457,N_6344,N_6330);
xnor U7458 (N_7458,N_6777,N_6142);
nand U7459 (N_7459,N_6692,N_6127);
or U7460 (N_7460,N_6175,N_6577);
nor U7461 (N_7461,N_6978,N_6829);
xnor U7462 (N_7462,N_6356,N_6246);
nor U7463 (N_7463,N_6478,N_6412);
nor U7464 (N_7464,N_6841,N_6480);
nand U7465 (N_7465,N_6640,N_6710);
nor U7466 (N_7466,N_6060,N_6815);
xnor U7467 (N_7467,N_6167,N_6041);
nor U7468 (N_7468,N_6941,N_6081);
nor U7469 (N_7469,N_6149,N_6014);
and U7470 (N_7470,N_6453,N_6960);
nor U7471 (N_7471,N_6687,N_6760);
or U7472 (N_7472,N_6529,N_6785);
nand U7473 (N_7473,N_6511,N_6058);
nand U7474 (N_7474,N_6964,N_6487);
nor U7475 (N_7475,N_6242,N_6275);
and U7476 (N_7476,N_6932,N_6807);
and U7477 (N_7477,N_6034,N_6359);
nor U7478 (N_7478,N_6406,N_6997);
or U7479 (N_7479,N_6238,N_6322);
and U7480 (N_7480,N_6258,N_6839);
nor U7481 (N_7481,N_6802,N_6350);
xor U7482 (N_7482,N_6772,N_6822);
and U7483 (N_7483,N_6786,N_6463);
and U7484 (N_7484,N_6947,N_6485);
xnor U7485 (N_7485,N_6646,N_6437);
xnor U7486 (N_7486,N_6848,N_6442);
and U7487 (N_7487,N_6614,N_6313);
or U7488 (N_7488,N_6357,N_6940);
nor U7489 (N_7489,N_6803,N_6809);
xnor U7490 (N_7490,N_6237,N_6842);
or U7491 (N_7491,N_6476,N_6402);
xnor U7492 (N_7492,N_6139,N_6381);
xnor U7493 (N_7493,N_6647,N_6872);
and U7494 (N_7494,N_6671,N_6134);
or U7495 (N_7495,N_6130,N_6880);
and U7496 (N_7496,N_6024,N_6762);
nor U7497 (N_7497,N_6279,N_6911);
xnor U7498 (N_7498,N_6290,N_6958);
or U7499 (N_7499,N_6769,N_6045);
nor U7500 (N_7500,N_6858,N_6443);
and U7501 (N_7501,N_6929,N_6445);
or U7502 (N_7502,N_6987,N_6950);
nor U7503 (N_7503,N_6902,N_6690);
xor U7504 (N_7504,N_6207,N_6095);
or U7505 (N_7505,N_6068,N_6763);
xor U7506 (N_7506,N_6135,N_6313);
xor U7507 (N_7507,N_6391,N_6528);
nand U7508 (N_7508,N_6104,N_6022);
nand U7509 (N_7509,N_6020,N_6104);
nor U7510 (N_7510,N_6518,N_6117);
or U7511 (N_7511,N_6230,N_6238);
xnor U7512 (N_7512,N_6166,N_6468);
nor U7513 (N_7513,N_6062,N_6396);
and U7514 (N_7514,N_6528,N_6764);
or U7515 (N_7515,N_6448,N_6761);
or U7516 (N_7516,N_6492,N_6580);
or U7517 (N_7517,N_6944,N_6692);
and U7518 (N_7518,N_6711,N_6969);
and U7519 (N_7519,N_6711,N_6765);
xnor U7520 (N_7520,N_6763,N_6290);
or U7521 (N_7521,N_6391,N_6889);
and U7522 (N_7522,N_6168,N_6281);
xnor U7523 (N_7523,N_6145,N_6493);
nand U7524 (N_7524,N_6433,N_6757);
nand U7525 (N_7525,N_6066,N_6412);
or U7526 (N_7526,N_6137,N_6280);
xnor U7527 (N_7527,N_6100,N_6368);
and U7528 (N_7528,N_6920,N_6184);
xor U7529 (N_7529,N_6782,N_6901);
and U7530 (N_7530,N_6214,N_6131);
or U7531 (N_7531,N_6044,N_6455);
or U7532 (N_7532,N_6658,N_6971);
nand U7533 (N_7533,N_6969,N_6252);
and U7534 (N_7534,N_6332,N_6792);
nand U7535 (N_7535,N_6821,N_6823);
nand U7536 (N_7536,N_6643,N_6603);
xnor U7537 (N_7537,N_6601,N_6015);
xnor U7538 (N_7538,N_6648,N_6798);
xnor U7539 (N_7539,N_6072,N_6264);
and U7540 (N_7540,N_6231,N_6730);
nor U7541 (N_7541,N_6290,N_6951);
nand U7542 (N_7542,N_6548,N_6113);
and U7543 (N_7543,N_6505,N_6253);
nor U7544 (N_7544,N_6510,N_6942);
xnor U7545 (N_7545,N_6125,N_6640);
xnor U7546 (N_7546,N_6844,N_6932);
or U7547 (N_7547,N_6636,N_6577);
and U7548 (N_7548,N_6452,N_6706);
nor U7549 (N_7549,N_6038,N_6759);
nand U7550 (N_7550,N_6313,N_6749);
or U7551 (N_7551,N_6962,N_6230);
and U7552 (N_7552,N_6373,N_6618);
nor U7553 (N_7553,N_6163,N_6357);
nand U7554 (N_7554,N_6139,N_6048);
and U7555 (N_7555,N_6443,N_6837);
and U7556 (N_7556,N_6491,N_6304);
and U7557 (N_7557,N_6784,N_6953);
and U7558 (N_7558,N_6873,N_6098);
nor U7559 (N_7559,N_6351,N_6064);
xnor U7560 (N_7560,N_6375,N_6039);
nor U7561 (N_7561,N_6408,N_6311);
and U7562 (N_7562,N_6007,N_6359);
nor U7563 (N_7563,N_6778,N_6473);
xnor U7564 (N_7564,N_6667,N_6797);
nor U7565 (N_7565,N_6086,N_6005);
and U7566 (N_7566,N_6041,N_6567);
nor U7567 (N_7567,N_6334,N_6299);
or U7568 (N_7568,N_6902,N_6128);
and U7569 (N_7569,N_6009,N_6418);
or U7570 (N_7570,N_6072,N_6529);
xnor U7571 (N_7571,N_6085,N_6489);
or U7572 (N_7572,N_6796,N_6876);
or U7573 (N_7573,N_6383,N_6362);
or U7574 (N_7574,N_6395,N_6706);
xor U7575 (N_7575,N_6799,N_6832);
nand U7576 (N_7576,N_6405,N_6222);
nor U7577 (N_7577,N_6099,N_6393);
and U7578 (N_7578,N_6740,N_6817);
xnor U7579 (N_7579,N_6900,N_6203);
or U7580 (N_7580,N_6206,N_6215);
xnor U7581 (N_7581,N_6667,N_6411);
or U7582 (N_7582,N_6646,N_6269);
nand U7583 (N_7583,N_6606,N_6435);
or U7584 (N_7584,N_6869,N_6135);
xor U7585 (N_7585,N_6301,N_6742);
xor U7586 (N_7586,N_6854,N_6907);
and U7587 (N_7587,N_6584,N_6798);
or U7588 (N_7588,N_6850,N_6176);
nor U7589 (N_7589,N_6188,N_6736);
and U7590 (N_7590,N_6161,N_6723);
nand U7591 (N_7591,N_6501,N_6899);
or U7592 (N_7592,N_6122,N_6488);
or U7593 (N_7593,N_6630,N_6385);
or U7594 (N_7594,N_6284,N_6909);
xor U7595 (N_7595,N_6374,N_6404);
nand U7596 (N_7596,N_6838,N_6672);
and U7597 (N_7597,N_6759,N_6635);
nor U7598 (N_7598,N_6259,N_6072);
nor U7599 (N_7599,N_6935,N_6421);
nand U7600 (N_7600,N_6401,N_6203);
nand U7601 (N_7601,N_6852,N_6739);
nand U7602 (N_7602,N_6267,N_6101);
or U7603 (N_7603,N_6037,N_6774);
nor U7604 (N_7604,N_6270,N_6330);
xor U7605 (N_7605,N_6236,N_6799);
xnor U7606 (N_7606,N_6347,N_6073);
and U7607 (N_7607,N_6260,N_6371);
nand U7608 (N_7608,N_6203,N_6904);
and U7609 (N_7609,N_6082,N_6231);
or U7610 (N_7610,N_6833,N_6263);
nor U7611 (N_7611,N_6775,N_6162);
and U7612 (N_7612,N_6085,N_6020);
nor U7613 (N_7613,N_6032,N_6141);
and U7614 (N_7614,N_6431,N_6297);
and U7615 (N_7615,N_6531,N_6153);
nor U7616 (N_7616,N_6931,N_6088);
xnor U7617 (N_7617,N_6871,N_6953);
or U7618 (N_7618,N_6796,N_6995);
and U7619 (N_7619,N_6706,N_6741);
or U7620 (N_7620,N_6552,N_6470);
nand U7621 (N_7621,N_6091,N_6277);
and U7622 (N_7622,N_6033,N_6594);
nor U7623 (N_7623,N_6871,N_6522);
nand U7624 (N_7624,N_6854,N_6815);
xor U7625 (N_7625,N_6359,N_6058);
and U7626 (N_7626,N_6455,N_6185);
nor U7627 (N_7627,N_6807,N_6090);
nand U7628 (N_7628,N_6415,N_6728);
or U7629 (N_7629,N_6835,N_6126);
nor U7630 (N_7630,N_6254,N_6927);
nor U7631 (N_7631,N_6593,N_6846);
xnor U7632 (N_7632,N_6786,N_6278);
xnor U7633 (N_7633,N_6607,N_6888);
nand U7634 (N_7634,N_6548,N_6013);
nand U7635 (N_7635,N_6822,N_6138);
or U7636 (N_7636,N_6058,N_6747);
nand U7637 (N_7637,N_6357,N_6848);
nor U7638 (N_7638,N_6103,N_6779);
nand U7639 (N_7639,N_6726,N_6688);
nand U7640 (N_7640,N_6774,N_6584);
nand U7641 (N_7641,N_6191,N_6538);
or U7642 (N_7642,N_6510,N_6990);
and U7643 (N_7643,N_6846,N_6240);
xor U7644 (N_7644,N_6205,N_6886);
nand U7645 (N_7645,N_6999,N_6862);
nor U7646 (N_7646,N_6498,N_6361);
nor U7647 (N_7647,N_6738,N_6457);
nor U7648 (N_7648,N_6401,N_6338);
and U7649 (N_7649,N_6623,N_6841);
xnor U7650 (N_7650,N_6671,N_6527);
and U7651 (N_7651,N_6718,N_6008);
or U7652 (N_7652,N_6751,N_6163);
xor U7653 (N_7653,N_6920,N_6063);
or U7654 (N_7654,N_6931,N_6454);
nand U7655 (N_7655,N_6288,N_6297);
nand U7656 (N_7656,N_6048,N_6811);
nor U7657 (N_7657,N_6500,N_6186);
or U7658 (N_7658,N_6112,N_6326);
or U7659 (N_7659,N_6515,N_6674);
or U7660 (N_7660,N_6860,N_6709);
nand U7661 (N_7661,N_6103,N_6181);
xnor U7662 (N_7662,N_6866,N_6220);
xnor U7663 (N_7663,N_6288,N_6233);
nor U7664 (N_7664,N_6515,N_6028);
nor U7665 (N_7665,N_6255,N_6083);
xor U7666 (N_7666,N_6704,N_6535);
or U7667 (N_7667,N_6631,N_6517);
nor U7668 (N_7668,N_6572,N_6834);
and U7669 (N_7669,N_6636,N_6073);
nor U7670 (N_7670,N_6579,N_6114);
nor U7671 (N_7671,N_6988,N_6309);
and U7672 (N_7672,N_6495,N_6053);
nor U7673 (N_7673,N_6032,N_6819);
nand U7674 (N_7674,N_6424,N_6922);
and U7675 (N_7675,N_6491,N_6480);
nand U7676 (N_7676,N_6731,N_6965);
nand U7677 (N_7677,N_6841,N_6674);
and U7678 (N_7678,N_6066,N_6598);
nand U7679 (N_7679,N_6576,N_6442);
or U7680 (N_7680,N_6753,N_6668);
nand U7681 (N_7681,N_6873,N_6675);
nor U7682 (N_7682,N_6865,N_6270);
xnor U7683 (N_7683,N_6791,N_6188);
nor U7684 (N_7684,N_6922,N_6225);
or U7685 (N_7685,N_6845,N_6545);
or U7686 (N_7686,N_6489,N_6946);
nand U7687 (N_7687,N_6771,N_6760);
nand U7688 (N_7688,N_6166,N_6140);
xor U7689 (N_7689,N_6215,N_6809);
nor U7690 (N_7690,N_6035,N_6138);
or U7691 (N_7691,N_6866,N_6358);
nand U7692 (N_7692,N_6600,N_6450);
nand U7693 (N_7693,N_6134,N_6867);
or U7694 (N_7694,N_6869,N_6728);
nand U7695 (N_7695,N_6243,N_6721);
xor U7696 (N_7696,N_6959,N_6542);
and U7697 (N_7697,N_6465,N_6387);
xor U7698 (N_7698,N_6175,N_6668);
nor U7699 (N_7699,N_6865,N_6956);
and U7700 (N_7700,N_6592,N_6689);
and U7701 (N_7701,N_6202,N_6952);
nor U7702 (N_7702,N_6379,N_6464);
nor U7703 (N_7703,N_6471,N_6554);
and U7704 (N_7704,N_6545,N_6090);
and U7705 (N_7705,N_6088,N_6316);
nor U7706 (N_7706,N_6148,N_6809);
nand U7707 (N_7707,N_6817,N_6664);
xnor U7708 (N_7708,N_6480,N_6380);
and U7709 (N_7709,N_6619,N_6065);
xnor U7710 (N_7710,N_6212,N_6566);
xnor U7711 (N_7711,N_6190,N_6754);
or U7712 (N_7712,N_6174,N_6127);
and U7713 (N_7713,N_6749,N_6395);
or U7714 (N_7714,N_6076,N_6529);
and U7715 (N_7715,N_6729,N_6100);
nand U7716 (N_7716,N_6945,N_6016);
nor U7717 (N_7717,N_6022,N_6450);
and U7718 (N_7718,N_6001,N_6837);
nand U7719 (N_7719,N_6048,N_6438);
xor U7720 (N_7720,N_6388,N_6584);
xor U7721 (N_7721,N_6021,N_6119);
and U7722 (N_7722,N_6779,N_6055);
and U7723 (N_7723,N_6352,N_6323);
and U7724 (N_7724,N_6557,N_6490);
and U7725 (N_7725,N_6267,N_6727);
and U7726 (N_7726,N_6057,N_6761);
nand U7727 (N_7727,N_6215,N_6141);
xor U7728 (N_7728,N_6936,N_6552);
xor U7729 (N_7729,N_6746,N_6234);
and U7730 (N_7730,N_6473,N_6752);
nor U7731 (N_7731,N_6903,N_6121);
or U7732 (N_7732,N_6003,N_6988);
xnor U7733 (N_7733,N_6195,N_6231);
nand U7734 (N_7734,N_6256,N_6048);
xnor U7735 (N_7735,N_6708,N_6701);
nor U7736 (N_7736,N_6159,N_6416);
nand U7737 (N_7737,N_6299,N_6828);
xnor U7738 (N_7738,N_6440,N_6133);
and U7739 (N_7739,N_6677,N_6651);
and U7740 (N_7740,N_6324,N_6953);
nand U7741 (N_7741,N_6527,N_6741);
nor U7742 (N_7742,N_6271,N_6230);
or U7743 (N_7743,N_6163,N_6192);
and U7744 (N_7744,N_6465,N_6817);
or U7745 (N_7745,N_6981,N_6795);
or U7746 (N_7746,N_6710,N_6918);
xor U7747 (N_7747,N_6311,N_6892);
and U7748 (N_7748,N_6006,N_6233);
or U7749 (N_7749,N_6762,N_6050);
and U7750 (N_7750,N_6222,N_6507);
or U7751 (N_7751,N_6022,N_6482);
nand U7752 (N_7752,N_6487,N_6654);
xnor U7753 (N_7753,N_6903,N_6639);
nand U7754 (N_7754,N_6239,N_6070);
or U7755 (N_7755,N_6994,N_6573);
nor U7756 (N_7756,N_6910,N_6405);
xor U7757 (N_7757,N_6856,N_6767);
or U7758 (N_7758,N_6497,N_6354);
nand U7759 (N_7759,N_6545,N_6873);
nor U7760 (N_7760,N_6833,N_6912);
xnor U7761 (N_7761,N_6985,N_6073);
xor U7762 (N_7762,N_6888,N_6854);
and U7763 (N_7763,N_6518,N_6358);
nor U7764 (N_7764,N_6893,N_6790);
xnor U7765 (N_7765,N_6084,N_6709);
xnor U7766 (N_7766,N_6790,N_6189);
xor U7767 (N_7767,N_6519,N_6049);
and U7768 (N_7768,N_6387,N_6193);
or U7769 (N_7769,N_6865,N_6217);
and U7770 (N_7770,N_6630,N_6032);
nor U7771 (N_7771,N_6140,N_6569);
nor U7772 (N_7772,N_6835,N_6228);
nand U7773 (N_7773,N_6351,N_6111);
nor U7774 (N_7774,N_6128,N_6696);
nor U7775 (N_7775,N_6821,N_6446);
or U7776 (N_7776,N_6101,N_6282);
and U7777 (N_7777,N_6680,N_6954);
and U7778 (N_7778,N_6757,N_6966);
or U7779 (N_7779,N_6247,N_6661);
nand U7780 (N_7780,N_6088,N_6770);
nand U7781 (N_7781,N_6204,N_6806);
or U7782 (N_7782,N_6278,N_6660);
nand U7783 (N_7783,N_6157,N_6466);
and U7784 (N_7784,N_6644,N_6423);
nor U7785 (N_7785,N_6170,N_6549);
xnor U7786 (N_7786,N_6251,N_6696);
nand U7787 (N_7787,N_6042,N_6029);
xnor U7788 (N_7788,N_6535,N_6260);
or U7789 (N_7789,N_6370,N_6030);
xor U7790 (N_7790,N_6207,N_6123);
and U7791 (N_7791,N_6755,N_6090);
xnor U7792 (N_7792,N_6498,N_6647);
nor U7793 (N_7793,N_6729,N_6964);
xor U7794 (N_7794,N_6466,N_6909);
or U7795 (N_7795,N_6085,N_6775);
nor U7796 (N_7796,N_6857,N_6306);
nor U7797 (N_7797,N_6214,N_6612);
nor U7798 (N_7798,N_6510,N_6973);
nand U7799 (N_7799,N_6987,N_6336);
and U7800 (N_7800,N_6444,N_6412);
nand U7801 (N_7801,N_6831,N_6193);
and U7802 (N_7802,N_6216,N_6399);
or U7803 (N_7803,N_6180,N_6375);
or U7804 (N_7804,N_6402,N_6834);
xor U7805 (N_7805,N_6093,N_6062);
nor U7806 (N_7806,N_6563,N_6651);
nand U7807 (N_7807,N_6890,N_6759);
or U7808 (N_7808,N_6878,N_6128);
nor U7809 (N_7809,N_6463,N_6807);
nor U7810 (N_7810,N_6332,N_6337);
xnor U7811 (N_7811,N_6293,N_6137);
nand U7812 (N_7812,N_6028,N_6069);
nand U7813 (N_7813,N_6183,N_6070);
nor U7814 (N_7814,N_6408,N_6175);
or U7815 (N_7815,N_6779,N_6597);
and U7816 (N_7816,N_6055,N_6271);
and U7817 (N_7817,N_6014,N_6771);
nor U7818 (N_7818,N_6575,N_6882);
and U7819 (N_7819,N_6030,N_6657);
and U7820 (N_7820,N_6218,N_6084);
xor U7821 (N_7821,N_6268,N_6961);
xor U7822 (N_7822,N_6082,N_6969);
xnor U7823 (N_7823,N_6439,N_6194);
nor U7824 (N_7824,N_6247,N_6317);
or U7825 (N_7825,N_6493,N_6192);
or U7826 (N_7826,N_6680,N_6975);
nand U7827 (N_7827,N_6132,N_6336);
and U7828 (N_7828,N_6769,N_6682);
xor U7829 (N_7829,N_6362,N_6923);
nand U7830 (N_7830,N_6720,N_6928);
nor U7831 (N_7831,N_6310,N_6093);
nand U7832 (N_7832,N_6055,N_6530);
and U7833 (N_7833,N_6349,N_6785);
or U7834 (N_7834,N_6794,N_6799);
and U7835 (N_7835,N_6664,N_6516);
and U7836 (N_7836,N_6922,N_6755);
nand U7837 (N_7837,N_6987,N_6337);
nor U7838 (N_7838,N_6711,N_6147);
nor U7839 (N_7839,N_6376,N_6742);
nand U7840 (N_7840,N_6715,N_6596);
xor U7841 (N_7841,N_6641,N_6313);
nand U7842 (N_7842,N_6135,N_6618);
nor U7843 (N_7843,N_6004,N_6178);
and U7844 (N_7844,N_6222,N_6943);
and U7845 (N_7845,N_6125,N_6646);
nor U7846 (N_7846,N_6172,N_6459);
xor U7847 (N_7847,N_6199,N_6183);
or U7848 (N_7848,N_6875,N_6954);
xor U7849 (N_7849,N_6847,N_6693);
or U7850 (N_7850,N_6089,N_6051);
xnor U7851 (N_7851,N_6599,N_6259);
xnor U7852 (N_7852,N_6974,N_6503);
and U7853 (N_7853,N_6538,N_6807);
xor U7854 (N_7854,N_6240,N_6437);
or U7855 (N_7855,N_6525,N_6268);
nand U7856 (N_7856,N_6803,N_6030);
or U7857 (N_7857,N_6807,N_6159);
nor U7858 (N_7858,N_6933,N_6861);
and U7859 (N_7859,N_6166,N_6620);
or U7860 (N_7860,N_6883,N_6590);
or U7861 (N_7861,N_6593,N_6198);
and U7862 (N_7862,N_6963,N_6471);
xor U7863 (N_7863,N_6298,N_6554);
nand U7864 (N_7864,N_6510,N_6120);
nor U7865 (N_7865,N_6034,N_6299);
nand U7866 (N_7866,N_6039,N_6714);
or U7867 (N_7867,N_6038,N_6154);
xor U7868 (N_7868,N_6628,N_6344);
nor U7869 (N_7869,N_6274,N_6882);
xor U7870 (N_7870,N_6636,N_6516);
or U7871 (N_7871,N_6778,N_6697);
nand U7872 (N_7872,N_6604,N_6011);
and U7873 (N_7873,N_6208,N_6182);
or U7874 (N_7874,N_6369,N_6963);
nor U7875 (N_7875,N_6141,N_6174);
or U7876 (N_7876,N_6239,N_6258);
nand U7877 (N_7877,N_6166,N_6055);
xor U7878 (N_7878,N_6187,N_6692);
nand U7879 (N_7879,N_6940,N_6115);
nand U7880 (N_7880,N_6194,N_6303);
or U7881 (N_7881,N_6071,N_6416);
or U7882 (N_7882,N_6004,N_6453);
and U7883 (N_7883,N_6123,N_6884);
xor U7884 (N_7884,N_6734,N_6465);
or U7885 (N_7885,N_6826,N_6803);
nor U7886 (N_7886,N_6576,N_6574);
and U7887 (N_7887,N_6578,N_6402);
xor U7888 (N_7888,N_6009,N_6901);
and U7889 (N_7889,N_6946,N_6947);
or U7890 (N_7890,N_6211,N_6858);
or U7891 (N_7891,N_6393,N_6768);
nand U7892 (N_7892,N_6247,N_6301);
nand U7893 (N_7893,N_6164,N_6223);
or U7894 (N_7894,N_6733,N_6543);
or U7895 (N_7895,N_6139,N_6093);
and U7896 (N_7896,N_6205,N_6430);
nor U7897 (N_7897,N_6851,N_6566);
and U7898 (N_7898,N_6142,N_6474);
nor U7899 (N_7899,N_6886,N_6405);
nand U7900 (N_7900,N_6235,N_6440);
or U7901 (N_7901,N_6666,N_6513);
xnor U7902 (N_7902,N_6954,N_6067);
nor U7903 (N_7903,N_6637,N_6048);
nor U7904 (N_7904,N_6345,N_6911);
nand U7905 (N_7905,N_6202,N_6314);
nand U7906 (N_7906,N_6540,N_6234);
or U7907 (N_7907,N_6048,N_6224);
nand U7908 (N_7908,N_6040,N_6683);
nor U7909 (N_7909,N_6032,N_6285);
nor U7910 (N_7910,N_6262,N_6573);
and U7911 (N_7911,N_6236,N_6270);
nor U7912 (N_7912,N_6205,N_6069);
xnor U7913 (N_7913,N_6282,N_6459);
and U7914 (N_7914,N_6983,N_6626);
or U7915 (N_7915,N_6790,N_6631);
nor U7916 (N_7916,N_6399,N_6125);
nor U7917 (N_7917,N_6361,N_6009);
xnor U7918 (N_7918,N_6483,N_6120);
nor U7919 (N_7919,N_6668,N_6456);
nor U7920 (N_7920,N_6578,N_6680);
and U7921 (N_7921,N_6375,N_6774);
or U7922 (N_7922,N_6217,N_6412);
xnor U7923 (N_7923,N_6565,N_6445);
nand U7924 (N_7924,N_6612,N_6603);
nor U7925 (N_7925,N_6033,N_6739);
xor U7926 (N_7926,N_6532,N_6654);
and U7927 (N_7927,N_6499,N_6496);
or U7928 (N_7928,N_6375,N_6892);
or U7929 (N_7929,N_6482,N_6009);
nor U7930 (N_7930,N_6259,N_6730);
nor U7931 (N_7931,N_6905,N_6077);
nand U7932 (N_7932,N_6076,N_6975);
or U7933 (N_7933,N_6861,N_6316);
xnor U7934 (N_7934,N_6009,N_6780);
or U7935 (N_7935,N_6002,N_6368);
nand U7936 (N_7936,N_6208,N_6010);
and U7937 (N_7937,N_6897,N_6139);
nand U7938 (N_7938,N_6487,N_6580);
nand U7939 (N_7939,N_6447,N_6157);
xnor U7940 (N_7940,N_6151,N_6877);
xnor U7941 (N_7941,N_6748,N_6507);
and U7942 (N_7942,N_6842,N_6051);
nor U7943 (N_7943,N_6465,N_6874);
nor U7944 (N_7944,N_6681,N_6848);
nand U7945 (N_7945,N_6275,N_6197);
nor U7946 (N_7946,N_6844,N_6834);
nand U7947 (N_7947,N_6347,N_6718);
and U7948 (N_7948,N_6825,N_6476);
xor U7949 (N_7949,N_6647,N_6178);
nand U7950 (N_7950,N_6137,N_6481);
nand U7951 (N_7951,N_6161,N_6034);
nor U7952 (N_7952,N_6589,N_6297);
nand U7953 (N_7953,N_6808,N_6452);
and U7954 (N_7954,N_6804,N_6295);
or U7955 (N_7955,N_6486,N_6999);
nor U7956 (N_7956,N_6462,N_6650);
xnor U7957 (N_7957,N_6616,N_6802);
xor U7958 (N_7958,N_6217,N_6408);
or U7959 (N_7959,N_6565,N_6454);
nor U7960 (N_7960,N_6649,N_6873);
xnor U7961 (N_7961,N_6170,N_6298);
and U7962 (N_7962,N_6638,N_6057);
and U7963 (N_7963,N_6881,N_6996);
or U7964 (N_7964,N_6479,N_6610);
xor U7965 (N_7965,N_6083,N_6134);
nor U7966 (N_7966,N_6431,N_6093);
nand U7967 (N_7967,N_6768,N_6287);
and U7968 (N_7968,N_6952,N_6205);
nand U7969 (N_7969,N_6301,N_6908);
xnor U7970 (N_7970,N_6420,N_6816);
and U7971 (N_7971,N_6163,N_6149);
nor U7972 (N_7972,N_6483,N_6178);
xnor U7973 (N_7973,N_6292,N_6855);
and U7974 (N_7974,N_6328,N_6273);
or U7975 (N_7975,N_6918,N_6486);
and U7976 (N_7976,N_6676,N_6606);
nand U7977 (N_7977,N_6423,N_6344);
nor U7978 (N_7978,N_6700,N_6277);
nor U7979 (N_7979,N_6192,N_6663);
nand U7980 (N_7980,N_6604,N_6970);
or U7981 (N_7981,N_6578,N_6827);
nor U7982 (N_7982,N_6825,N_6300);
and U7983 (N_7983,N_6736,N_6233);
nand U7984 (N_7984,N_6168,N_6397);
and U7985 (N_7985,N_6579,N_6561);
nor U7986 (N_7986,N_6168,N_6999);
and U7987 (N_7987,N_6190,N_6842);
and U7988 (N_7988,N_6266,N_6907);
nand U7989 (N_7989,N_6751,N_6992);
nand U7990 (N_7990,N_6428,N_6418);
nor U7991 (N_7991,N_6004,N_6512);
and U7992 (N_7992,N_6685,N_6008);
nor U7993 (N_7993,N_6689,N_6197);
and U7994 (N_7994,N_6708,N_6726);
and U7995 (N_7995,N_6341,N_6227);
nor U7996 (N_7996,N_6281,N_6257);
xnor U7997 (N_7997,N_6568,N_6992);
nor U7998 (N_7998,N_6559,N_6353);
nor U7999 (N_7999,N_6337,N_6422);
and U8000 (N_8000,N_7750,N_7892);
or U8001 (N_8001,N_7417,N_7996);
and U8002 (N_8002,N_7576,N_7574);
nor U8003 (N_8003,N_7936,N_7336);
and U8004 (N_8004,N_7265,N_7715);
nor U8005 (N_8005,N_7186,N_7605);
xor U8006 (N_8006,N_7058,N_7876);
nor U8007 (N_8007,N_7707,N_7304);
nand U8008 (N_8008,N_7433,N_7077);
nand U8009 (N_8009,N_7423,N_7473);
nor U8010 (N_8010,N_7994,N_7967);
xnor U8011 (N_8011,N_7158,N_7611);
nand U8012 (N_8012,N_7462,N_7407);
or U8013 (N_8013,N_7248,N_7298);
xnor U8014 (N_8014,N_7213,N_7926);
or U8015 (N_8015,N_7237,N_7736);
nand U8016 (N_8016,N_7831,N_7500);
or U8017 (N_8017,N_7722,N_7579);
and U8018 (N_8018,N_7993,N_7343);
and U8019 (N_8019,N_7073,N_7119);
or U8020 (N_8020,N_7698,N_7641);
or U8021 (N_8021,N_7367,N_7839);
nor U8022 (N_8022,N_7911,N_7045);
nor U8023 (N_8023,N_7710,N_7215);
or U8024 (N_8024,N_7814,N_7016);
or U8025 (N_8025,N_7866,N_7513);
xnor U8026 (N_8026,N_7446,N_7759);
xnor U8027 (N_8027,N_7506,N_7673);
xnor U8028 (N_8028,N_7036,N_7120);
nand U8029 (N_8029,N_7572,N_7081);
or U8030 (N_8030,N_7100,N_7915);
nand U8031 (N_8031,N_7218,N_7365);
nand U8032 (N_8032,N_7087,N_7477);
nand U8033 (N_8033,N_7226,N_7459);
nand U8034 (N_8034,N_7929,N_7803);
or U8035 (N_8035,N_7686,N_7674);
xor U8036 (N_8036,N_7053,N_7559);
xnor U8037 (N_8037,N_7313,N_7984);
xnor U8038 (N_8038,N_7653,N_7429);
and U8039 (N_8039,N_7162,N_7648);
xor U8040 (N_8040,N_7819,N_7028);
or U8041 (N_8041,N_7895,N_7905);
xnor U8042 (N_8042,N_7622,N_7052);
and U8043 (N_8043,N_7359,N_7899);
nand U8044 (N_8044,N_7230,N_7428);
nor U8045 (N_8045,N_7614,N_7564);
nor U8046 (N_8046,N_7840,N_7533);
or U8047 (N_8047,N_7591,N_7980);
xnor U8048 (N_8048,N_7509,N_7140);
nor U8049 (N_8049,N_7727,N_7725);
xnor U8050 (N_8050,N_7330,N_7118);
or U8051 (N_8051,N_7370,N_7160);
nor U8052 (N_8052,N_7373,N_7882);
xnor U8053 (N_8053,N_7885,N_7387);
and U8054 (N_8054,N_7691,N_7247);
nor U8055 (N_8055,N_7130,N_7512);
xnor U8056 (N_8056,N_7449,N_7078);
and U8057 (N_8057,N_7689,N_7794);
nor U8058 (N_8058,N_7971,N_7595);
and U8059 (N_8059,N_7632,N_7626);
and U8060 (N_8060,N_7867,N_7761);
xor U8061 (N_8061,N_7744,N_7390);
or U8062 (N_8062,N_7999,N_7953);
or U8063 (N_8063,N_7930,N_7811);
xor U8064 (N_8064,N_7068,N_7117);
nand U8065 (N_8065,N_7034,N_7849);
nand U8066 (N_8066,N_7221,N_7402);
and U8067 (N_8067,N_7029,N_7862);
nand U8068 (N_8068,N_7392,N_7280);
xor U8069 (N_8069,N_7085,N_7709);
nand U8070 (N_8070,N_7272,N_7664);
nor U8071 (N_8071,N_7630,N_7601);
nand U8072 (N_8072,N_7244,N_7870);
xor U8073 (N_8073,N_7793,N_7854);
or U8074 (N_8074,N_7471,N_7510);
and U8075 (N_8075,N_7483,N_7812);
nor U8076 (N_8076,N_7655,N_7652);
nor U8077 (N_8077,N_7333,N_7779);
nand U8078 (N_8078,N_7475,N_7421);
xnor U8079 (N_8079,N_7657,N_7598);
xnor U8080 (N_8080,N_7954,N_7735);
and U8081 (N_8081,N_7056,N_7565);
nor U8082 (N_8082,N_7419,N_7238);
or U8083 (N_8083,N_7554,N_7193);
nand U8084 (N_8084,N_7478,N_7562);
or U8085 (N_8085,N_7381,N_7532);
nor U8086 (N_8086,N_7852,N_7426);
and U8087 (N_8087,N_7216,N_7089);
and U8088 (N_8088,N_7939,N_7873);
xor U8089 (N_8089,N_7252,N_7302);
nand U8090 (N_8090,N_7150,N_7138);
xnor U8091 (N_8091,N_7638,N_7733);
or U8092 (N_8092,N_7306,N_7753);
nand U8093 (N_8093,N_7716,N_7080);
nand U8094 (N_8094,N_7714,N_7325);
nor U8095 (N_8095,N_7484,N_7185);
xor U8096 (N_8096,N_7338,N_7377);
or U8097 (N_8097,N_7051,N_7164);
xnor U8098 (N_8098,N_7422,N_7724);
or U8099 (N_8099,N_7127,N_7297);
nor U8100 (N_8100,N_7692,N_7846);
or U8101 (N_8101,N_7728,N_7476);
or U8102 (N_8102,N_7181,N_7444);
or U8103 (N_8103,N_7502,N_7227);
nor U8104 (N_8104,N_7030,N_7091);
or U8105 (N_8105,N_7524,N_7871);
nor U8106 (N_8106,N_7437,N_7439);
and U8107 (N_8107,N_7159,N_7411);
nor U8108 (N_8108,N_7115,N_7869);
or U8109 (N_8109,N_7389,N_7983);
nor U8110 (N_8110,N_7264,N_7789);
or U8111 (N_8111,N_7038,N_7308);
or U8112 (N_8112,N_7182,N_7580);
or U8113 (N_8113,N_7799,N_7401);
and U8114 (N_8114,N_7253,N_7575);
xnor U8115 (N_8115,N_7263,N_7763);
nand U8116 (N_8116,N_7166,N_7545);
and U8117 (N_8117,N_7589,N_7331);
and U8118 (N_8118,N_7132,N_7382);
nand U8119 (N_8119,N_7944,N_7555);
and U8120 (N_8120,N_7225,N_7084);
xnor U8121 (N_8121,N_7332,N_7925);
and U8122 (N_8122,N_7588,N_7109);
nand U8123 (N_8123,N_7898,N_7070);
nand U8124 (N_8124,N_7146,N_7742);
and U8125 (N_8125,N_7619,N_7531);
xor U8126 (N_8126,N_7291,N_7661);
nand U8127 (N_8127,N_7153,N_7918);
xor U8128 (N_8128,N_7875,N_7455);
and U8129 (N_8129,N_7299,N_7734);
nand U8130 (N_8130,N_7538,N_7995);
xor U8131 (N_8131,N_7678,N_7520);
nand U8132 (N_8132,N_7813,N_7222);
or U8133 (N_8133,N_7443,N_7639);
nand U8134 (N_8134,N_7284,N_7550);
or U8135 (N_8135,N_7800,N_7825);
nor U8136 (N_8136,N_7457,N_7792);
nor U8137 (N_8137,N_7771,N_7540);
and U8138 (N_8138,N_7324,N_7516);
nand U8139 (N_8139,N_7514,N_7631);
nor U8140 (N_8140,N_7064,N_7864);
and U8141 (N_8141,N_7416,N_7860);
xor U8142 (N_8142,N_7818,N_7234);
or U8143 (N_8143,N_7277,N_7289);
xnor U8144 (N_8144,N_7775,N_7910);
nand U8145 (N_8145,N_7287,N_7394);
nand U8146 (N_8146,N_7749,N_7354);
nor U8147 (N_8147,N_7326,N_7179);
and U8148 (N_8148,N_7436,N_7530);
and U8149 (N_8149,N_7693,N_7095);
and U8150 (N_8150,N_7738,N_7337);
xor U8151 (N_8151,N_7801,N_7434);
or U8152 (N_8152,N_7442,N_7711);
nor U8153 (N_8153,N_7178,N_7209);
and U8154 (N_8154,N_7041,N_7743);
xnor U8155 (N_8155,N_7582,N_7278);
xor U8156 (N_8156,N_7927,N_7395);
nor U8157 (N_8157,N_7857,N_7345);
nor U8158 (N_8158,N_7680,N_7460);
and U8159 (N_8159,N_7152,N_7438);
or U8160 (N_8160,N_7566,N_7900);
nand U8161 (N_8161,N_7820,N_7561);
nor U8162 (N_8162,N_7257,N_7031);
or U8163 (N_8163,N_7398,N_7685);
or U8164 (N_8164,N_7951,N_7184);
and U8165 (N_8165,N_7061,N_7069);
nor U8166 (N_8166,N_7328,N_7773);
or U8167 (N_8167,N_7785,N_7766);
nand U8168 (N_8168,N_7379,N_7223);
and U8169 (N_8169,N_7526,N_7380);
or U8170 (N_8170,N_7656,N_7042);
or U8171 (N_8171,N_7039,N_7805);
and U8172 (N_8172,N_7616,N_7891);
or U8173 (N_8173,N_7323,N_7646);
nand U8174 (N_8174,N_7780,N_7625);
xnor U8175 (N_8175,N_7977,N_7249);
xnor U8176 (N_8176,N_7102,N_7283);
xnor U8177 (N_8177,N_7916,N_7292);
nor U8178 (N_8178,N_7001,N_7096);
xor U8179 (N_8179,N_7956,N_7063);
nand U8180 (N_8180,N_7143,N_7023);
or U8181 (N_8181,N_7720,N_7634);
or U8182 (N_8182,N_7467,N_7665);
or U8183 (N_8183,N_7836,N_7107);
or U8184 (N_8184,N_7482,N_7155);
nand U8185 (N_8185,N_7239,N_7784);
and U8186 (N_8186,N_7912,N_7981);
xor U8187 (N_8187,N_7020,N_7347);
or U8188 (N_8188,N_7650,N_7364);
and U8189 (N_8189,N_7676,N_7568);
or U8190 (N_8190,N_7335,N_7368);
and U8191 (N_8191,N_7106,N_7004);
nand U8192 (N_8192,N_7266,N_7511);
and U8193 (N_8193,N_7696,N_7060);
or U8194 (N_8194,N_7172,N_7961);
and U8195 (N_8195,N_7383,N_7469);
xor U8196 (N_8196,N_7047,N_7404);
xor U8197 (N_8197,N_7319,N_7214);
xor U8198 (N_8198,N_7282,N_7755);
nand U8199 (N_8199,N_7139,N_7960);
or U8200 (N_8200,N_7486,N_7732);
xnor U8201 (N_8201,N_7991,N_7826);
and U8202 (N_8202,N_7731,N_7168);
or U8203 (N_8203,N_7942,N_7537);
xor U8204 (N_8204,N_7441,N_7125);
nor U8205 (N_8205,N_7659,N_7192);
nor U8206 (N_8206,N_7397,N_7649);
nand U8207 (N_8207,N_7592,N_7878);
or U8208 (N_8208,N_7342,N_7212);
and U8209 (N_8209,N_7975,N_7872);
and U8210 (N_8210,N_7134,N_7447);
or U8211 (N_8211,N_7704,N_7346);
or U8212 (N_8212,N_7590,N_7494);
or U8213 (N_8213,N_7741,N_7048);
xor U8214 (N_8214,N_7809,N_7262);
nand U8215 (N_8215,N_7640,N_7933);
nand U8216 (N_8216,N_7002,N_7830);
nor U8217 (N_8217,N_7019,N_7504);
xor U8218 (N_8218,N_7986,N_7288);
or U8219 (N_8219,N_7585,N_7211);
xor U8220 (N_8220,N_7348,N_7705);
nor U8221 (N_8221,N_7388,N_7105);
or U8222 (N_8222,N_7260,N_7154);
xor U8223 (N_8223,N_7316,N_7480);
and U8224 (N_8224,N_7362,N_7396);
xor U8225 (N_8225,N_7987,N_7391);
and U8226 (N_8226,N_7834,N_7551);
nor U8227 (N_8227,N_7190,N_7874);
nand U8228 (N_8228,N_7197,N_7843);
nand U8229 (N_8229,N_7848,N_7353);
nand U8230 (N_8230,N_7205,N_7199);
or U8231 (N_8231,N_7121,N_7970);
xor U8232 (N_8232,N_7046,N_7523);
and U8233 (N_8233,N_7093,N_7706);
or U8234 (N_8234,N_7414,N_7075);
and U8235 (N_8235,N_7082,N_7274);
or U8236 (N_8236,N_7189,N_7712);
nand U8237 (N_8237,N_7907,N_7018);
nand U8238 (N_8238,N_7112,N_7094);
and U8239 (N_8239,N_7007,N_7982);
xor U8240 (N_8240,N_7492,N_7145);
or U8241 (N_8241,N_7740,N_7235);
xor U8242 (N_8242,N_7098,N_7050);
nand U8243 (N_8243,N_7463,N_7989);
or U8244 (N_8244,N_7695,N_7005);
xnor U8245 (N_8245,N_7880,N_7853);
xnor U8246 (N_8246,N_7195,N_7418);
nand U8247 (N_8247,N_7726,N_7969);
or U8248 (N_8248,N_7300,N_7156);
xnor U8249 (N_8249,N_7952,N_7642);
nand U8250 (N_8250,N_7790,N_7810);
and U8251 (N_8251,N_7948,N_7546);
and U8252 (N_8252,N_7578,N_7116);
nor U8253 (N_8253,N_7497,N_7838);
nor U8254 (N_8254,N_7481,N_7188);
and U8255 (N_8255,N_7147,N_7913);
xor U8256 (N_8256,N_7668,N_7856);
nand U8257 (N_8257,N_7934,N_7947);
xnor U8258 (N_8258,N_7043,N_7774);
nand U8259 (N_8259,N_7548,N_7795);
or U8260 (N_8260,N_7610,N_7307);
and U8261 (N_8261,N_7806,N_7972);
or U8262 (N_8262,N_7133,N_7747);
nand U8263 (N_8263,N_7142,N_7006);
or U8264 (N_8264,N_7889,N_7489);
nor U8265 (N_8265,N_7553,N_7279);
or U8266 (N_8266,N_7405,N_7203);
xnor U8267 (N_8267,N_7472,N_7083);
or U8268 (N_8268,N_7352,N_7276);
or U8269 (N_8269,N_7009,N_7600);
nor U8270 (N_8270,N_7758,N_7713);
xnor U8271 (N_8271,N_7943,N_7752);
or U8272 (N_8272,N_7543,N_7552);
and U8273 (N_8273,N_7493,N_7914);
xnor U8274 (N_8274,N_7978,N_7011);
or U8275 (N_8275,N_7470,N_7563);
nand U8276 (N_8276,N_7966,N_7861);
nor U8277 (N_8277,N_7584,N_7123);
or U8278 (N_8278,N_7988,N_7474);
and U8279 (N_8279,N_7832,N_7255);
nor U8280 (N_8280,N_7267,N_7355);
or U8281 (N_8281,N_7356,N_7660);
and U8282 (N_8282,N_7224,N_7985);
and U8283 (N_8283,N_7157,N_7863);
or U8284 (N_8284,N_7902,N_7904);
xnor U8285 (N_8285,N_7310,N_7458);
and U8286 (N_8286,N_7108,N_7903);
nand U8287 (N_8287,N_7859,N_7850);
xor U8288 (N_8288,N_7651,N_7453);
and U8289 (N_8289,N_7173,N_7496);
and U8290 (N_8290,N_7240,N_7541);
or U8291 (N_8291,N_7938,N_7901);
or U8292 (N_8292,N_7964,N_7535);
nand U8293 (N_8293,N_7022,N_7827);
nand U8294 (N_8294,N_7448,N_7637);
and U8295 (N_8295,N_7066,N_7430);
and U8296 (N_8296,N_7770,N_7415);
or U8297 (N_8297,N_7618,N_7717);
xor U8298 (N_8298,N_7886,N_7896);
nand U8299 (N_8299,N_7887,N_7440);
or U8300 (N_8300,N_7594,N_7945);
nand U8301 (N_8301,N_7339,N_7329);
nand U8302 (N_8302,N_7816,N_7645);
or U8303 (N_8303,N_7177,N_7037);
nand U8304 (N_8304,N_7167,N_7386);
or U8305 (N_8305,N_7644,N_7583);
and U8306 (N_8306,N_7466,N_7014);
xor U8307 (N_8307,N_7044,N_7236);
and U8308 (N_8308,N_7054,N_7521);
nor U8309 (N_8309,N_7376,N_7748);
xnor U8310 (N_8310,N_7729,N_7294);
nor U8311 (N_8311,N_7684,N_7270);
xnor U8312 (N_8312,N_7090,N_7627);
nor U8313 (N_8313,N_7932,N_7435);
xnor U8314 (N_8314,N_7135,N_7424);
nor U8315 (N_8315,N_7450,N_7208);
nor U8316 (N_8316,N_7220,N_7783);
nor U8317 (N_8317,N_7890,N_7671);
nor U8318 (N_8318,N_7824,N_7596);
xor U8319 (N_8319,N_7241,N_7427);
and U8320 (N_8320,N_7454,N_7242);
and U8321 (N_8321,N_7250,N_7515);
nor U8322 (N_8322,N_7719,N_7363);
or U8323 (N_8323,N_7519,N_7357);
and U8324 (N_8324,N_7025,N_7754);
and U8325 (N_8325,N_7350,N_7126);
and U8326 (N_8326,N_7615,N_7767);
and U8327 (N_8327,N_7577,N_7488);
or U8328 (N_8328,N_7269,N_7917);
nor U8329 (N_8329,N_7635,N_7593);
nand U8330 (N_8330,N_7040,N_7321);
or U8331 (N_8331,N_7919,N_7174);
or U8332 (N_8332,N_7499,N_7908);
and U8333 (N_8333,N_7950,N_7024);
xor U8334 (N_8334,N_7219,N_7703);
nor U8335 (N_8335,N_7990,N_7161);
and U8336 (N_8336,N_7431,N_7293);
or U8337 (N_8337,N_7522,N_7957);
nand U8338 (N_8338,N_7032,N_7008);
or U8339 (N_8339,N_7361,N_7788);
nor U8340 (N_8340,N_7739,N_7525);
xnor U8341 (N_8341,N_7968,N_7688);
and U8342 (N_8342,N_7670,N_7768);
and U8343 (N_8343,N_7372,N_7104);
nand U8344 (N_8344,N_7847,N_7194);
nor U8345 (N_8345,N_7808,N_7074);
xor U8346 (N_8346,N_7452,N_7737);
or U8347 (N_8347,N_7647,N_7567);
xor U8348 (N_8348,N_7305,N_7406);
and U8349 (N_8349,N_7662,N_7807);
nand U8350 (N_8350,N_7959,N_7017);
nor U8351 (N_8351,N_7400,N_7701);
nand U8352 (N_8352,N_7245,N_7974);
and U8353 (N_8353,N_7271,N_7015);
or U8354 (N_8354,N_7349,N_7268);
xnor U8355 (N_8355,N_7062,N_7101);
and U8356 (N_8356,N_7682,N_7201);
or U8357 (N_8357,N_7920,N_7769);
and U8358 (N_8358,N_7320,N_7922);
or U8359 (N_8359,N_7010,N_7965);
xnor U8360 (N_8360,N_7229,N_7581);
xnor U8361 (N_8361,N_7384,N_7318);
nor U8362 (N_8362,N_7196,N_7787);
and U8363 (N_8363,N_7835,N_7612);
or U8364 (N_8364,N_7765,N_7071);
xor U8365 (N_8365,N_7171,N_7327);
nor U8366 (N_8366,N_7000,N_7207);
or U8367 (N_8367,N_7169,N_7344);
nand U8368 (N_8368,N_7613,N_7149);
nor U8369 (N_8369,N_7776,N_7621);
and U8370 (N_8370,N_7629,N_7340);
or U8371 (N_8371,N_7412,N_7675);
and U8372 (N_8372,N_7931,N_7527);
and U8373 (N_8373,N_7508,N_7962);
or U8374 (N_8374,N_7569,N_7351);
and U8375 (N_8375,N_7111,N_7425);
nand U8376 (N_8376,N_7558,N_7003);
nor U8377 (N_8377,N_7573,N_7777);
nor U8378 (N_8378,N_7841,N_7833);
or U8379 (N_8379,N_7296,N_7358);
xnor U8380 (N_8380,N_7700,N_7233);
or U8381 (N_8381,N_7165,N_7817);
or U8382 (N_8382,N_7491,N_7501);
or U8383 (N_8383,N_7941,N_7254);
nand U8384 (N_8384,N_7557,N_7183);
or U8385 (N_8385,N_7366,N_7888);
or U8386 (N_8386,N_7609,N_7597);
or U8387 (N_8387,N_7822,N_7796);
nand U8388 (N_8388,N_7322,N_7851);
nor U8389 (N_8389,N_7163,N_7539);
or U8390 (N_8390,N_7694,N_7536);
or U8391 (N_8391,N_7529,N_7033);
or U8392 (N_8392,N_7528,N_7175);
nor U8393 (N_8393,N_7517,N_7868);
nand U8394 (N_8394,N_7667,N_7072);
nor U8395 (N_8395,N_7503,N_7092);
or U8396 (N_8396,N_7923,N_7113);
nor U8397 (N_8397,N_7256,N_7403);
xor U8398 (N_8398,N_7883,N_7456);
or U8399 (N_8399,N_7067,N_7385);
and U8400 (N_8400,N_7607,N_7187);
or U8401 (N_8401,N_7587,N_7314);
or U8402 (N_8402,N_7955,N_7928);
or U8403 (N_8403,N_7290,N_7815);
nand U8404 (N_8404,N_7858,N_7495);
xor U8405 (N_8405,N_7285,N_7751);
xnor U8406 (N_8406,N_7821,N_7408);
or U8407 (N_8407,N_7451,N_7603);
nand U8408 (N_8408,N_7781,N_7312);
or U8409 (N_8409,N_7180,N_7251);
xnor U8410 (N_8410,N_7097,N_7823);
xnor U8411 (N_8411,N_7798,N_7301);
nor U8412 (N_8412,N_7746,N_7399);
xor U8413 (N_8413,N_7136,N_7893);
and U8414 (N_8414,N_7586,N_7026);
or U8415 (N_8415,N_7697,N_7206);
nand U8416 (N_8416,N_7413,N_7341);
xor U8417 (N_8417,N_7231,N_7804);
or U8418 (N_8418,N_7261,N_7702);
nand U8419 (N_8419,N_7170,N_7842);
or U8420 (N_8420,N_7721,N_7756);
nor U8421 (N_8421,N_7672,N_7683);
nor U8422 (N_8422,N_7487,N_7103);
nand U8423 (N_8423,N_7949,N_7628);
xor U8424 (N_8424,N_7369,N_7542);
xor U8425 (N_8425,N_7829,N_7654);
or U8426 (N_8426,N_7534,N_7623);
nor U8427 (N_8427,N_7124,N_7723);
nor U8428 (N_8428,N_7643,N_7420);
xor U8429 (N_8429,N_7958,N_7217);
or U8430 (N_8430,N_7498,N_7079);
xor U8431 (N_8431,N_7375,N_7275);
or U8432 (N_8432,N_7604,N_7129);
nor U8433 (N_8433,N_7273,N_7490);
or U8434 (N_8434,N_7802,N_7485);
xor U8435 (N_8435,N_7303,N_7937);
xnor U8436 (N_8436,N_7881,N_7243);
nand U8437 (N_8437,N_7393,N_7059);
nand U8438 (N_8438,N_7110,N_7764);
nand U8439 (N_8439,N_7099,N_7571);
or U8440 (N_8440,N_7049,N_7035);
nand U8441 (N_8441,N_7176,N_7730);
nor U8442 (N_8442,N_7371,N_7148);
or U8443 (N_8443,N_7828,N_7295);
or U8444 (N_8444,N_7973,N_7012);
and U8445 (N_8445,N_7465,N_7258);
and U8446 (N_8446,N_7602,N_7556);
xor U8447 (N_8447,N_7549,N_7131);
xnor U8448 (N_8448,N_7879,N_7570);
or U8449 (N_8449,N_7606,N_7246);
and U8450 (N_8450,N_7445,N_7762);
and U8451 (N_8451,N_7461,N_7151);
or U8452 (N_8452,N_7315,N_7141);
xnor U8453 (N_8453,N_7877,N_7432);
xnor U8454 (N_8454,N_7547,N_7374);
and U8455 (N_8455,N_7198,N_7979);
or U8456 (N_8456,N_7021,N_7894);
nor U8457 (N_8457,N_7200,N_7128);
nand U8458 (N_8458,N_7317,N_7617);
or U8459 (N_8459,N_7505,N_7760);
nand U8460 (N_8460,N_7281,N_7624);
xor U8461 (N_8461,N_7608,N_7507);
or U8462 (N_8462,N_7309,N_7409);
and U8463 (N_8463,N_7786,N_7921);
or U8464 (N_8464,N_7013,N_7679);
or U8465 (N_8465,N_7410,N_7086);
nor U8466 (N_8466,N_7782,N_7334);
nand U8467 (N_8467,N_7076,N_7636);
nand U8468 (N_8468,N_7906,N_7837);
xor U8469 (N_8469,N_7976,N_7464);
nand U8470 (N_8470,N_7518,N_7055);
nand U8471 (N_8471,N_7057,N_7468);
or U8472 (N_8472,N_7963,N_7757);
or U8473 (N_8473,N_7620,N_7228);
or U8474 (N_8474,N_7663,N_7088);
xor U8475 (N_8475,N_7772,N_7778);
xnor U8476 (N_8476,N_7378,N_7992);
nand U8477 (N_8477,N_7360,N_7259);
xnor U8478 (N_8478,N_7666,N_7909);
nand U8479 (N_8479,N_7122,N_7897);
xor U8480 (N_8480,N_7998,N_7677);
nor U8481 (N_8481,N_7924,N_7946);
or U8482 (N_8482,N_7599,N_7544);
xnor U8483 (N_8483,N_7286,N_7311);
nand U8484 (N_8484,N_7202,N_7114);
nor U8485 (N_8485,N_7658,N_7855);
nand U8486 (N_8486,N_7690,N_7797);
xnor U8487 (N_8487,N_7940,N_7844);
xor U8488 (N_8488,N_7791,N_7137);
xnor U8489 (N_8489,N_7669,N_7845);
and U8490 (N_8490,N_7997,N_7699);
nand U8491 (N_8491,N_7633,N_7027);
nor U8492 (N_8492,N_7232,N_7191);
nand U8493 (N_8493,N_7745,N_7718);
nand U8494 (N_8494,N_7204,N_7687);
or U8495 (N_8495,N_7210,N_7681);
nor U8496 (N_8496,N_7560,N_7865);
or U8497 (N_8497,N_7479,N_7884);
nand U8498 (N_8498,N_7144,N_7935);
nor U8499 (N_8499,N_7065,N_7708);
or U8500 (N_8500,N_7161,N_7199);
nand U8501 (N_8501,N_7572,N_7045);
nor U8502 (N_8502,N_7966,N_7844);
nand U8503 (N_8503,N_7901,N_7660);
or U8504 (N_8504,N_7752,N_7745);
nor U8505 (N_8505,N_7400,N_7929);
xnor U8506 (N_8506,N_7750,N_7232);
nor U8507 (N_8507,N_7767,N_7572);
nand U8508 (N_8508,N_7405,N_7530);
nor U8509 (N_8509,N_7998,N_7495);
and U8510 (N_8510,N_7203,N_7272);
and U8511 (N_8511,N_7440,N_7389);
nor U8512 (N_8512,N_7491,N_7374);
and U8513 (N_8513,N_7248,N_7338);
or U8514 (N_8514,N_7404,N_7849);
and U8515 (N_8515,N_7421,N_7419);
and U8516 (N_8516,N_7796,N_7921);
nand U8517 (N_8517,N_7761,N_7255);
nor U8518 (N_8518,N_7017,N_7565);
xor U8519 (N_8519,N_7758,N_7316);
and U8520 (N_8520,N_7175,N_7721);
and U8521 (N_8521,N_7939,N_7988);
nor U8522 (N_8522,N_7861,N_7217);
xor U8523 (N_8523,N_7493,N_7478);
nand U8524 (N_8524,N_7013,N_7140);
nand U8525 (N_8525,N_7442,N_7456);
and U8526 (N_8526,N_7856,N_7991);
xnor U8527 (N_8527,N_7090,N_7523);
and U8528 (N_8528,N_7110,N_7122);
nor U8529 (N_8529,N_7763,N_7715);
nand U8530 (N_8530,N_7654,N_7221);
nand U8531 (N_8531,N_7040,N_7171);
nor U8532 (N_8532,N_7615,N_7953);
and U8533 (N_8533,N_7450,N_7668);
or U8534 (N_8534,N_7778,N_7954);
nand U8535 (N_8535,N_7617,N_7541);
or U8536 (N_8536,N_7862,N_7632);
nand U8537 (N_8537,N_7056,N_7362);
or U8538 (N_8538,N_7899,N_7076);
nor U8539 (N_8539,N_7657,N_7061);
and U8540 (N_8540,N_7941,N_7750);
nand U8541 (N_8541,N_7575,N_7172);
nand U8542 (N_8542,N_7887,N_7482);
xor U8543 (N_8543,N_7516,N_7120);
nand U8544 (N_8544,N_7630,N_7174);
and U8545 (N_8545,N_7174,N_7767);
nor U8546 (N_8546,N_7039,N_7273);
or U8547 (N_8547,N_7236,N_7391);
nor U8548 (N_8548,N_7825,N_7167);
nor U8549 (N_8549,N_7344,N_7821);
and U8550 (N_8550,N_7867,N_7515);
or U8551 (N_8551,N_7165,N_7259);
xnor U8552 (N_8552,N_7246,N_7095);
nand U8553 (N_8553,N_7649,N_7027);
xnor U8554 (N_8554,N_7406,N_7520);
and U8555 (N_8555,N_7521,N_7383);
xnor U8556 (N_8556,N_7765,N_7064);
and U8557 (N_8557,N_7252,N_7494);
or U8558 (N_8558,N_7469,N_7824);
and U8559 (N_8559,N_7419,N_7153);
or U8560 (N_8560,N_7247,N_7110);
and U8561 (N_8561,N_7016,N_7064);
xor U8562 (N_8562,N_7339,N_7113);
and U8563 (N_8563,N_7970,N_7943);
or U8564 (N_8564,N_7631,N_7188);
nand U8565 (N_8565,N_7109,N_7317);
and U8566 (N_8566,N_7761,N_7239);
nand U8567 (N_8567,N_7668,N_7558);
and U8568 (N_8568,N_7367,N_7964);
nor U8569 (N_8569,N_7519,N_7951);
nor U8570 (N_8570,N_7835,N_7650);
nor U8571 (N_8571,N_7571,N_7595);
and U8572 (N_8572,N_7437,N_7685);
nand U8573 (N_8573,N_7467,N_7697);
nand U8574 (N_8574,N_7968,N_7845);
or U8575 (N_8575,N_7765,N_7560);
or U8576 (N_8576,N_7908,N_7749);
nand U8577 (N_8577,N_7914,N_7482);
xnor U8578 (N_8578,N_7561,N_7893);
nor U8579 (N_8579,N_7881,N_7836);
nor U8580 (N_8580,N_7352,N_7896);
nand U8581 (N_8581,N_7517,N_7365);
or U8582 (N_8582,N_7105,N_7784);
and U8583 (N_8583,N_7555,N_7629);
and U8584 (N_8584,N_7928,N_7778);
or U8585 (N_8585,N_7654,N_7435);
nand U8586 (N_8586,N_7735,N_7597);
xor U8587 (N_8587,N_7974,N_7933);
nand U8588 (N_8588,N_7933,N_7894);
nand U8589 (N_8589,N_7341,N_7309);
nor U8590 (N_8590,N_7243,N_7860);
xor U8591 (N_8591,N_7712,N_7099);
nor U8592 (N_8592,N_7526,N_7923);
xor U8593 (N_8593,N_7202,N_7826);
or U8594 (N_8594,N_7153,N_7190);
nand U8595 (N_8595,N_7585,N_7044);
nor U8596 (N_8596,N_7591,N_7888);
and U8597 (N_8597,N_7898,N_7014);
or U8598 (N_8598,N_7641,N_7662);
or U8599 (N_8599,N_7026,N_7769);
or U8600 (N_8600,N_7889,N_7261);
xnor U8601 (N_8601,N_7514,N_7207);
nand U8602 (N_8602,N_7829,N_7539);
nand U8603 (N_8603,N_7275,N_7028);
nand U8604 (N_8604,N_7745,N_7220);
or U8605 (N_8605,N_7909,N_7763);
xnor U8606 (N_8606,N_7067,N_7696);
nor U8607 (N_8607,N_7725,N_7554);
and U8608 (N_8608,N_7887,N_7464);
nor U8609 (N_8609,N_7935,N_7859);
or U8610 (N_8610,N_7084,N_7530);
nand U8611 (N_8611,N_7264,N_7074);
and U8612 (N_8612,N_7293,N_7231);
or U8613 (N_8613,N_7174,N_7904);
and U8614 (N_8614,N_7379,N_7411);
nand U8615 (N_8615,N_7626,N_7876);
or U8616 (N_8616,N_7588,N_7302);
or U8617 (N_8617,N_7424,N_7205);
xor U8618 (N_8618,N_7694,N_7533);
nand U8619 (N_8619,N_7979,N_7819);
nand U8620 (N_8620,N_7132,N_7428);
or U8621 (N_8621,N_7976,N_7056);
nand U8622 (N_8622,N_7642,N_7516);
and U8623 (N_8623,N_7356,N_7051);
nor U8624 (N_8624,N_7498,N_7268);
xnor U8625 (N_8625,N_7357,N_7585);
nand U8626 (N_8626,N_7044,N_7053);
nor U8627 (N_8627,N_7732,N_7583);
nand U8628 (N_8628,N_7565,N_7331);
xor U8629 (N_8629,N_7461,N_7816);
nor U8630 (N_8630,N_7942,N_7293);
nor U8631 (N_8631,N_7698,N_7545);
nand U8632 (N_8632,N_7235,N_7728);
nor U8633 (N_8633,N_7636,N_7109);
or U8634 (N_8634,N_7638,N_7554);
nor U8635 (N_8635,N_7101,N_7427);
nor U8636 (N_8636,N_7620,N_7517);
nor U8637 (N_8637,N_7788,N_7288);
or U8638 (N_8638,N_7256,N_7194);
nor U8639 (N_8639,N_7089,N_7068);
or U8640 (N_8640,N_7323,N_7957);
xor U8641 (N_8641,N_7441,N_7900);
xor U8642 (N_8642,N_7113,N_7603);
and U8643 (N_8643,N_7123,N_7062);
nand U8644 (N_8644,N_7084,N_7642);
xor U8645 (N_8645,N_7174,N_7185);
or U8646 (N_8646,N_7005,N_7665);
and U8647 (N_8647,N_7069,N_7088);
nor U8648 (N_8648,N_7471,N_7876);
nand U8649 (N_8649,N_7498,N_7449);
and U8650 (N_8650,N_7958,N_7698);
or U8651 (N_8651,N_7781,N_7733);
and U8652 (N_8652,N_7490,N_7286);
or U8653 (N_8653,N_7855,N_7885);
and U8654 (N_8654,N_7874,N_7595);
or U8655 (N_8655,N_7797,N_7852);
nand U8656 (N_8656,N_7329,N_7094);
nand U8657 (N_8657,N_7618,N_7789);
nand U8658 (N_8658,N_7018,N_7132);
or U8659 (N_8659,N_7754,N_7911);
or U8660 (N_8660,N_7319,N_7366);
xnor U8661 (N_8661,N_7770,N_7171);
and U8662 (N_8662,N_7861,N_7617);
nor U8663 (N_8663,N_7200,N_7253);
and U8664 (N_8664,N_7477,N_7381);
nand U8665 (N_8665,N_7210,N_7926);
and U8666 (N_8666,N_7176,N_7789);
nor U8667 (N_8667,N_7730,N_7761);
nor U8668 (N_8668,N_7052,N_7821);
xnor U8669 (N_8669,N_7420,N_7182);
nand U8670 (N_8670,N_7908,N_7794);
nand U8671 (N_8671,N_7216,N_7330);
and U8672 (N_8672,N_7108,N_7074);
and U8673 (N_8673,N_7466,N_7792);
nand U8674 (N_8674,N_7237,N_7366);
and U8675 (N_8675,N_7544,N_7718);
nor U8676 (N_8676,N_7692,N_7279);
or U8677 (N_8677,N_7821,N_7616);
or U8678 (N_8678,N_7928,N_7465);
nor U8679 (N_8679,N_7397,N_7478);
xnor U8680 (N_8680,N_7377,N_7296);
and U8681 (N_8681,N_7435,N_7962);
nand U8682 (N_8682,N_7033,N_7346);
xnor U8683 (N_8683,N_7129,N_7925);
or U8684 (N_8684,N_7057,N_7842);
and U8685 (N_8685,N_7572,N_7396);
nand U8686 (N_8686,N_7047,N_7336);
xnor U8687 (N_8687,N_7028,N_7712);
nor U8688 (N_8688,N_7423,N_7668);
xor U8689 (N_8689,N_7147,N_7326);
nand U8690 (N_8690,N_7879,N_7885);
xor U8691 (N_8691,N_7803,N_7459);
nand U8692 (N_8692,N_7327,N_7973);
nor U8693 (N_8693,N_7134,N_7469);
and U8694 (N_8694,N_7199,N_7023);
or U8695 (N_8695,N_7317,N_7619);
and U8696 (N_8696,N_7142,N_7201);
nand U8697 (N_8697,N_7504,N_7156);
xor U8698 (N_8698,N_7049,N_7996);
or U8699 (N_8699,N_7027,N_7063);
nor U8700 (N_8700,N_7690,N_7427);
xnor U8701 (N_8701,N_7446,N_7488);
or U8702 (N_8702,N_7064,N_7725);
or U8703 (N_8703,N_7754,N_7896);
and U8704 (N_8704,N_7589,N_7421);
and U8705 (N_8705,N_7523,N_7887);
and U8706 (N_8706,N_7098,N_7729);
or U8707 (N_8707,N_7396,N_7421);
nand U8708 (N_8708,N_7920,N_7782);
nor U8709 (N_8709,N_7955,N_7649);
nor U8710 (N_8710,N_7063,N_7775);
and U8711 (N_8711,N_7919,N_7683);
xnor U8712 (N_8712,N_7129,N_7146);
or U8713 (N_8713,N_7610,N_7618);
and U8714 (N_8714,N_7099,N_7942);
nand U8715 (N_8715,N_7566,N_7016);
nor U8716 (N_8716,N_7933,N_7452);
or U8717 (N_8717,N_7911,N_7351);
nor U8718 (N_8718,N_7009,N_7988);
or U8719 (N_8719,N_7823,N_7767);
nand U8720 (N_8720,N_7000,N_7764);
nor U8721 (N_8721,N_7533,N_7067);
and U8722 (N_8722,N_7246,N_7964);
and U8723 (N_8723,N_7980,N_7713);
nand U8724 (N_8724,N_7704,N_7967);
and U8725 (N_8725,N_7875,N_7938);
xor U8726 (N_8726,N_7420,N_7974);
nand U8727 (N_8727,N_7813,N_7068);
nor U8728 (N_8728,N_7412,N_7747);
nand U8729 (N_8729,N_7999,N_7131);
nor U8730 (N_8730,N_7047,N_7658);
xnor U8731 (N_8731,N_7287,N_7828);
xor U8732 (N_8732,N_7780,N_7165);
and U8733 (N_8733,N_7258,N_7127);
xnor U8734 (N_8734,N_7302,N_7398);
nand U8735 (N_8735,N_7214,N_7561);
nand U8736 (N_8736,N_7979,N_7501);
nor U8737 (N_8737,N_7206,N_7798);
nand U8738 (N_8738,N_7061,N_7079);
nor U8739 (N_8739,N_7014,N_7975);
or U8740 (N_8740,N_7511,N_7951);
nand U8741 (N_8741,N_7507,N_7233);
and U8742 (N_8742,N_7837,N_7572);
and U8743 (N_8743,N_7528,N_7144);
nor U8744 (N_8744,N_7771,N_7031);
xnor U8745 (N_8745,N_7321,N_7202);
nor U8746 (N_8746,N_7522,N_7845);
nor U8747 (N_8747,N_7458,N_7153);
xnor U8748 (N_8748,N_7617,N_7868);
or U8749 (N_8749,N_7641,N_7142);
and U8750 (N_8750,N_7136,N_7430);
nand U8751 (N_8751,N_7437,N_7572);
or U8752 (N_8752,N_7772,N_7909);
or U8753 (N_8753,N_7961,N_7400);
or U8754 (N_8754,N_7776,N_7705);
nand U8755 (N_8755,N_7303,N_7123);
xnor U8756 (N_8756,N_7097,N_7771);
or U8757 (N_8757,N_7607,N_7851);
xor U8758 (N_8758,N_7580,N_7801);
nor U8759 (N_8759,N_7933,N_7418);
or U8760 (N_8760,N_7360,N_7689);
nand U8761 (N_8761,N_7280,N_7852);
and U8762 (N_8762,N_7632,N_7854);
xnor U8763 (N_8763,N_7333,N_7398);
xnor U8764 (N_8764,N_7157,N_7500);
xor U8765 (N_8765,N_7157,N_7339);
or U8766 (N_8766,N_7999,N_7657);
nand U8767 (N_8767,N_7653,N_7970);
or U8768 (N_8768,N_7861,N_7828);
xor U8769 (N_8769,N_7707,N_7897);
nor U8770 (N_8770,N_7640,N_7312);
xnor U8771 (N_8771,N_7825,N_7796);
nor U8772 (N_8772,N_7613,N_7741);
and U8773 (N_8773,N_7881,N_7608);
nand U8774 (N_8774,N_7860,N_7452);
nand U8775 (N_8775,N_7660,N_7723);
or U8776 (N_8776,N_7010,N_7087);
or U8777 (N_8777,N_7885,N_7309);
and U8778 (N_8778,N_7036,N_7440);
nand U8779 (N_8779,N_7212,N_7086);
nand U8780 (N_8780,N_7286,N_7757);
xnor U8781 (N_8781,N_7645,N_7334);
or U8782 (N_8782,N_7457,N_7886);
or U8783 (N_8783,N_7059,N_7732);
nand U8784 (N_8784,N_7344,N_7505);
and U8785 (N_8785,N_7251,N_7405);
or U8786 (N_8786,N_7827,N_7600);
nand U8787 (N_8787,N_7820,N_7939);
xnor U8788 (N_8788,N_7669,N_7984);
and U8789 (N_8789,N_7094,N_7686);
nand U8790 (N_8790,N_7667,N_7016);
nand U8791 (N_8791,N_7018,N_7462);
nor U8792 (N_8792,N_7237,N_7612);
or U8793 (N_8793,N_7350,N_7651);
or U8794 (N_8794,N_7926,N_7150);
nand U8795 (N_8795,N_7772,N_7055);
nand U8796 (N_8796,N_7533,N_7352);
xnor U8797 (N_8797,N_7269,N_7422);
xor U8798 (N_8798,N_7535,N_7398);
xnor U8799 (N_8799,N_7806,N_7772);
xor U8800 (N_8800,N_7988,N_7640);
nand U8801 (N_8801,N_7263,N_7445);
and U8802 (N_8802,N_7976,N_7083);
xnor U8803 (N_8803,N_7044,N_7030);
or U8804 (N_8804,N_7176,N_7923);
xor U8805 (N_8805,N_7335,N_7494);
xnor U8806 (N_8806,N_7629,N_7481);
nand U8807 (N_8807,N_7271,N_7362);
xor U8808 (N_8808,N_7504,N_7835);
and U8809 (N_8809,N_7078,N_7546);
or U8810 (N_8810,N_7544,N_7749);
nor U8811 (N_8811,N_7642,N_7557);
nor U8812 (N_8812,N_7546,N_7749);
nor U8813 (N_8813,N_7431,N_7878);
nand U8814 (N_8814,N_7824,N_7564);
nor U8815 (N_8815,N_7219,N_7480);
xnor U8816 (N_8816,N_7528,N_7996);
nor U8817 (N_8817,N_7305,N_7625);
xnor U8818 (N_8818,N_7075,N_7043);
nor U8819 (N_8819,N_7384,N_7984);
nand U8820 (N_8820,N_7403,N_7973);
or U8821 (N_8821,N_7760,N_7313);
nor U8822 (N_8822,N_7048,N_7355);
xor U8823 (N_8823,N_7068,N_7081);
or U8824 (N_8824,N_7615,N_7063);
and U8825 (N_8825,N_7522,N_7360);
or U8826 (N_8826,N_7592,N_7278);
or U8827 (N_8827,N_7271,N_7126);
nor U8828 (N_8828,N_7096,N_7044);
or U8829 (N_8829,N_7477,N_7287);
and U8830 (N_8830,N_7073,N_7197);
or U8831 (N_8831,N_7509,N_7994);
or U8832 (N_8832,N_7855,N_7107);
xnor U8833 (N_8833,N_7073,N_7203);
nand U8834 (N_8834,N_7721,N_7879);
or U8835 (N_8835,N_7307,N_7282);
nor U8836 (N_8836,N_7593,N_7293);
xnor U8837 (N_8837,N_7668,N_7469);
nor U8838 (N_8838,N_7491,N_7191);
or U8839 (N_8839,N_7446,N_7572);
or U8840 (N_8840,N_7382,N_7276);
nand U8841 (N_8841,N_7096,N_7772);
and U8842 (N_8842,N_7753,N_7727);
or U8843 (N_8843,N_7414,N_7983);
xnor U8844 (N_8844,N_7093,N_7229);
xor U8845 (N_8845,N_7949,N_7083);
or U8846 (N_8846,N_7868,N_7896);
and U8847 (N_8847,N_7929,N_7155);
nand U8848 (N_8848,N_7558,N_7134);
nor U8849 (N_8849,N_7328,N_7445);
xnor U8850 (N_8850,N_7543,N_7890);
xor U8851 (N_8851,N_7078,N_7324);
nor U8852 (N_8852,N_7636,N_7591);
and U8853 (N_8853,N_7518,N_7300);
nand U8854 (N_8854,N_7131,N_7085);
nand U8855 (N_8855,N_7340,N_7928);
nand U8856 (N_8856,N_7701,N_7690);
xor U8857 (N_8857,N_7642,N_7449);
and U8858 (N_8858,N_7198,N_7649);
nand U8859 (N_8859,N_7260,N_7520);
or U8860 (N_8860,N_7894,N_7576);
nand U8861 (N_8861,N_7762,N_7331);
xnor U8862 (N_8862,N_7504,N_7513);
or U8863 (N_8863,N_7162,N_7649);
and U8864 (N_8864,N_7363,N_7945);
nor U8865 (N_8865,N_7889,N_7600);
and U8866 (N_8866,N_7529,N_7858);
xnor U8867 (N_8867,N_7682,N_7737);
or U8868 (N_8868,N_7885,N_7089);
or U8869 (N_8869,N_7692,N_7592);
xor U8870 (N_8870,N_7689,N_7438);
and U8871 (N_8871,N_7510,N_7145);
xor U8872 (N_8872,N_7449,N_7311);
and U8873 (N_8873,N_7853,N_7651);
and U8874 (N_8874,N_7011,N_7529);
or U8875 (N_8875,N_7036,N_7685);
nand U8876 (N_8876,N_7386,N_7659);
nand U8877 (N_8877,N_7051,N_7923);
and U8878 (N_8878,N_7412,N_7902);
nand U8879 (N_8879,N_7315,N_7974);
or U8880 (N_8880,N_7799,N_7661);
nor U8881 (N_8881,N_7948,N_7070);
nand U8882 (N_8882,N_7430,N_7831);
nand U8883 (N_8883,N_7979,N_7292);
nand U8884 (N_8884,N_7395,N_7050);
nor U8885 (N_8885,N_7692,N_7852);
and U8886 (N_8886,N_7294,N_7810);
or U8887 (N_8887,N_7095,N_7242);
or U8888 (N_8888,N_7345,N_7753);
or U8889 (N_8889,N_7789,N_7352);
nor U8890 (N_8890,N_7090,N_7671);
and U8891 (N_8891,N_7419,N_7152);
and U8892 (N_8892,N_7142,N_7491);
nor U8893 (N_8893,N_7209,N_7021);
or U8894 (N_8894,N_7246,N_7127);
or U8895 (N_8895,N_7889,N_7498);
nor U8896 (N_8896,N_7024,N_7507);
nand U8897 (N_8897,N_7700,N_7807);
nand U8898 (N_8898,N_7848,N_7472);
or U8899 (N_8899,N_7580,N_7472);
xor U8900 (N_8900,N_7892,N_7347);
nand U8901 (N_8901,N_7275,N_7368);
nor U8902 (N_8902,N_7794,N_7150);
and U8903 (N_8903,N_7979,N_7997);
xnor U8904 (N_8904,N_7806,N_7977);
nand U8905 (N_8905,N_7882,N_7922);
or U8906 (N_8906,N_7951,N_7645);
or U8907 (N_8907,N_7481,N_7852);
nor U8908 (N_8908,N_7585,N_7139);
and U8909 (N_8909,N_7660,N_7535);
nand U8910 (N_8910,N_7406,N_7733);
nand U8911 (N_8911,N_7677,N_7826);
xor U8912 (N_8912,N_7734,N_7330);
nor U8913 (N_8913,N_7725,N_7676);
nor U8914 (N_8914,N_7557,N_7269);
and U8915 (N_8915,N_7915,N_7571);
or U8916 (N_8916,N_7806,N_7732);
or U8917 (N_8917,N_7382,N_7682);
nor U8918 (N_8918,N_7890,N_7835);
xnor U8919 (N_8919,N_7646,N_7893);
or U8920 (N_8920,N_7197,N_7020);
or U8921 (N_8921,N_7390,N_7644);
xor U8922 (N_8922,N_7234,N_7170);
or U8923 (N_8923,N_7260,N_7412);
or U8924 (N_8924,N_7988,N_7425);
and U8925 (N_8925,N_7461,N_7367);
nand U8926 (N_8926,N_7526,N_7204);
xnor U8927 (N_8927,N_7314,N_7575);
or U8928 (N_8928,N_7147,N_7725);
nor U8929 (N_8929,N_7883,N_7528);
and U8930 (N_8930,N_7724,N_7199);
nand U8931 (N_8931,N_7629,N_7619);
nor U8932 (N_8932,N_7504,N_7717);
nor U8933 (N_8933,N_7812,N_7088);
nor U8934 (N_8934,N_7404,N_7980);
xor U8935 (N_8935,N_7148,N_7631);
xor U8936 (N_8936,N_7766,N_7236);
nand U8937 (N_8937,N_7063,N_7695);
and U8938 (N_8938,N_7995,N_7690);
and U8939 (N_8939,N_7660,N_7481);
or U8940 (N_8940,N_7017,N_7312);
nor U8941 (N_8941,N_7638,N_7062);
nor U8942 (N_8942,N_7866,N_7358);
or U8943 (N_8943,N_7867,N_7315);
nor U8944 (N_8944,N_7253,N_7027);
and U8945 (N_8945,N_7170,N_7883);
or U8946 (N_8946,N_7725,N_7372);
xor U8947 (N_8947,N_7650,N_7219);
xor U8948 (N_8948,N_7899,N_7132);
and U8949 (N_8949,N_7140,N_7598);
xor U8950 (N_8950,N_7189,N_7369);
nor U8951 (N_8951,N_7775,N_7214);
nor U8952 (N_8952,N_7455,N_7731);
nor U8953 (N_8953,N_7587,N_7181);
or U8954 (N_8954,N_7080,N_7499);
nand U8955 (N_8955,N_7452,N_7438);
xor U8956 (N_8956,N_7242,N_7034);
xnor U8957 (N_8957,N_7345,N_7376);
nand U8958 (N_8958,N_7392,N_7401);
and U8959 (N_8959,N_7111,N_7216);
or U8960 (N_8960,N_7345,N_7832);
xnor U8961 (N_8961,N_7280,N_7843);
xor U8962 (N_8962,N_7567,N_7806);
or U8963 (N_8963,N_7928,N_7499);
xor U8964 (N_8964,N_7776,N_7201);
xnor U8965 (N_8965,N_7878,N_7009);
and U8966 (N_8966,N_7872,N_7481);
nor U8967 (N_8967,N_7225,N_7625);
xnor U8968 (N_8968,N_7718,N_7823);
or U8969 (N_8969,N_7547,N_7561);
or U8970 (N_8970,N_7583,N_7806);
or U8971 (N_8971,N_7768,N_7630);
nand U8972 (N_8972,N_7605,N_7596);
nor U8973 (N_8973,N_7002,N_7265);
nor U8974 (N_8974,N_7538,N_7582);
nand U8975 (N_8975,N_7522,N_7268);
xnor U8976 (N_8976,N_7423,N_7853);
or U8977 (N_8977,N_7207,N_7851);
xnor U8978 (N_8978,N_7402,N_7519);
and U8979 (N_8979,N_7413,N_7171);
or U8980 (N_8980,N_7131,N_7863);
nand U8981 (N_8981,N_7067,N_7930);
nor U8982 (N_8982,N_7044,N_7566);
nor U8983 (N_8983,N_7498,N_7683);
nand U8984 (N_8984,N_7257,N_7634);
or U8985 (N_8985,N_7642,N_7364);
nor U8986 (N_8986,N_7307,N_7047);
and U8987 (N_8987,N_7356,N_7117);
xor U8988 (N_8988,N_7571,N_7634);
nor U8989 (N_8989,N_7931,N_7113);
or U8990 (N_8990,N_7394,N_7923);
xor U8991 (N_8991,N_7027,N_7861);
or U8992 (N_8992,N_7695,N_7965);
nand U8993 (N_8993,N_7844,N_7107);
and U8994 (N_8994,N_7304,N_7553);
and U8995 (N_8995,N_7403,N_7757);
nand U8996 (N_8996,N_7161,N_7317);
nand U8997 (N_8997,N_7724,N_7553);
or U8998 (N_8998,N_7828,N_7176);
xnor U8999 (N_8999,N_7072,N_7099);
and U9000 (N_9000,N_8431,N_8678);
and U9001 (N_9001,N_8663,N_8981);
or U9002 (N_9002,N_8381,N_8156);
or U9003 (N_9003,N_8579,N_8417);
nor U9004 (N_9004,N_8573,N_8113);
and U9005 (N_9005,N_8641,N_8829);
or U9006 (N_9006,N_8031,N_8264);
xnor U9007 (N_9007,N_8250,N_8058);
nor U9008 (N_9008,N_8336,N_8041);
nand U9009 (N_9009,N_8762,N_8931);
xnor U9010 (N_9010,N_8209,N_8363);
and U9011 (N_9011,N_8481,N_8295);
or U9012 (N_9012,N_8406,N_8290);
nor U9013 (N_9013,N_8890,N_8834);
nand U9014 (N_9014,N_8909,N_8107);
and U9015 (N_9015,N_8294,N_8769);
and U9016 (N_9016,N_8649,N_8096);
nor U9017 (N_9017,N_8744,N_8202);
and U9018 (N_9018,N_8053,N_8100);
nor U9019 (N_9019,N_8459,N_8742);
nor U9020 (N_9020,N_8609,N_8748);
or U9021 (N_9021,N_8439,N_8135);
nor U9022 (N_9022,N_8035,N_8559);
or U9023 (N_9023,N_8389,N_8997);
or U9024 (N_9024,N_8804,N_8089);
nand U9025 (N_9025,N_8975,N_8359);
and U9026 (N_9026,N_8668,N_8013);
xor U9027 (N_9027,N_8042,N_8913);
nor U9028 (N_9028,N_8916,N_8048);
or U9029 (N_9029,N_8241,N_8868);
xor U9030 (N_9030,N_8011,N_8985);
and U9031 (N_9031,N_8647,N_8409);
or U9032 (N_9032,N_8937,N_8966);
xor U9033 (N_9033,N_8211,N_8343);
xnor U9034 (N_9034,N_8765,N_8725);
xnor U9035 (N_9035,N_8059,N_8116);
xnor U9036 (N_9036,N_8236,N_8587);
xor U9037 (N_9037,N_8703,N_8301);
nand U9038 (N_9038,N_8963,N_8738);
and U9039 (N_9039,N_8557,N_8495);
xor U9040 (N_9040,N_8606,N_8847);
xnor U9041 (N_9041,N_8940,N_8252);
nand U9042 (N_9042,N_8821,N_8124);
xor U9043 (N_9043,N_8243,N_8379);
nand U9044 (N_9044,N_8915,N_8869);
xnor U9045 (N_9045,N_8518,N_8531);
nand U9046 (N_9046,N_8297,N_8191);
and U9047 (N_9047,N_8127,N_8111);
or U9048 (N_9048,N_8945,N_8427);
and U9049 (N_9049,N_8911,N_8581);
nand U9050 (N_9050,N_8094,N_8622);
or U9051 (N_9051,N_8272,N_8240);
xnor U9052 (N_9052,N_8192,N_8049);
xor U9053 (N_9053,N_8207,N_8313);
and U9054 (N_9054,N_8793,N_8285);
or U9055 (N_9055,N_8176,N_8060);
and U9056 (N_9056,N_8522,N_8684);
nand U9057 (N_9057,N_8882,N_8688);
or U9058 (N_9058,N_8469,N_8012);
nand U9059 (N_9059,N_8160,N_8619);
and U9060 (N_9060,N_8922,N_8104);
xnor U9061 (N_9061,N_8468,N_8449);
and U9062 (N_9062,N_8970,N_8547);
and U9063 (N_9063,N_8450,N_8351);
and U9064 (N_9064,N_8624,N_8292);
nand U9065 (N_9065,N_8014,N_8134);
or U9066 (N_9066,N_8648,N_8463);
or U9067 (N_9067,N_8232,N_8877);
nor U9068 (N_9068,N_8885,N_8528);
nor U9069 (N_9069,N_8561,N_8539);
nor U9070 (N_9070,N_8411,N_8355);
or U9071 (N_9071,N_8628,N_8457);
or U9072 (N_9072,N_8125,N_8630);
and U9073 (N_9073,N_8052,N_8639);
xor U9074 (N_9074,N_8075,N_8269);
and U9075 (N_9075,N_8387,N_8825);
nor U9076 (N_9076,N_8588,N_8967);
xnor U9077 (N_9077,N_8289,N_8291);
or U9078 (N_9078,N_8896,N_8398);
and U9079 (N_9079,N_8442,N_8118);
or U9080 (N_9080,N_8245,N_8867);
or U9081 (N_9081,N_8563,N_8800);
and U9082 (N_9082,N_8412,N_8194);
xnor U9083 (N_9083,N_8597,N_8173);
nor U9084 (N_9084,N_8978,N_8991);
and U9085 (N_9085,N_8430,N_8872);
and U9086 (N_9086,N_8679,N_8914);
xor U9087 (N_9087,N_8831,N_8101);
nor U9088 (N_9088,N_8905,N_8006);
xor U9089 (N_9089,N_8939,N_8919);
and U9090 (N_9090,N_8165,N_8370);
or U9091 (N_9091,N_8485,N_8345);
or U9092 (N_9092,N_8889,N_8705);
xnor U9093 (N_9093,N_8000,N_8397);
nand U9094 (N_9094,N_8566,N_8342);
nand U9095 (N_9095,N_8399,N_8188);
xor U9096 (N_9096,N_8895,N_8611);
xor U9097 (N_9097,N_8731,N_8815);
or U9098 (N_9098,N_8613,N_8246);
nor U9099 (N_9099,N_8779,N_8848);
xnor U9100 (N_9100,N_8030,N_8064);
nand U9101 (N_9101,N_8591,N_8808);
or U9102 (N_9102,N_8316,N_8095);
and U9103 (N_9103,N_8008,N_8820);
and U9104 (N_9104,N_8857,N_8824);
and U9105 (N_9105,N_8015,N_8632);
or U9106 (N_9106,N_8129,N_8323);
nand U9107 (N_9107,N_8025,N_8498);
or U9108 (N_9108,N_8019,N_8876);
and U9109 (N_9109,N_8403,N_8056);
nand U9110 (N_9110,N_8852,N_8595);
and U9111 (N_9111,N_8608,N_8474);
and U9112 (N_9112,N_8426,N_8137);
or U9113 (N_9113,N_8667,N_8259);
nor U9114 (N_9114,N_8612,N_8879);
and U9115 (N_9115,N_8371,N_8061);
nor U9116 (N_9116,N_8594,N_8423);
or U9117 (N_9117,N_8733,N_8500);
and U9118 (N_9118,N_8103,N_8768);
nor U9119 (N_9119,N_8128,N_8216);
and U9120 (N_9120,N_8860,N_8925);
nand U9121 (N_9121,N_8620,N_8954);
xor U9122 (N_9122,N_8923,N_8842);
nor U9123 (N_9123,N_8535,N_8339);
nor U9124 (N_9124,N_8082,N_8664);
nor U9125 (N_9125,N_8887,N_8709);
or U9126 (N_9126,N_8550,N_8642);
and U9127 (N_9127,N_8473,N_8471);
xnor U9128 (N_9128,N_8974,N_8968);
xor U9129 (N_9129,N_8132,N_8607);
nand U9130 (N_9130,N_8517,N_8377);
or U9131 (N_9131,N_8537,N_8215);
and U9132 (N_9132,N_8745,N_8117);
nor U9133 (N_9133,N_8273,N_8136);
or U9134 (N_9134,N_8982,N_8179);
nor U9135 (N_9135,N_8907,N_8276);
xnor U9136 (N_9136,N_8254,N_8233);
nand U9137 (N_9137,N_8766,N_8479);
and U9138 (N_9138,N_8715,N_8263);
or U9139 (N_9139,N_8458,N_8033);
nor U9140 (N_9140,N_8166,N_8078);
nor U9141 (N_9141,N_8706,N_8454);
nor U9142 (N_9142,N_8516,N_8027);
or U9143 (N_9143,N_8849,N_8206);
and U9144 (N_9144,N_8984,N_8728);
xor U9145 (N_9145,N_8328,N_8392);
xor U9146 (N_9146,N_8112,N_8177);
and U9147 (N_9147,N_8146,N_8433);
or U9148 (N_9148,N_8776,N_8455);
and U9149 (N_9149,N_8636,N_8335);
or U9150 (N_9150,N_8900,N_8186);
xnor U9151 (N_9151,N_8674,N_8873);
and U9152 (N_9152,N_8115,N_8088);
nor U9153 (N_9153,N_8366,N_8741);
nor U9154 (N_9154,N_8770,N_8610);
and U9155 (N_9155,N_8452,N_8456);
nor U9156 (N_9156,N_8901,N_8929);
and U9157 (N_9157,N_8330,N_8773);
xor U9158 (N_9158,N_8099,N_8390);
nor U9159 (N_9159,N_8141,N_8029);
and U9160 (N_9160,N_8864,N_8955);
and U9161 (N_9161,N_8749,N_8348);
nand U9162 (N_9162,N_8614,N_8950);
nor U9163 (N_9163,N_8859,N_8902);
and U9164 (N_9164,N_8927,N_8076);
xnor U9165 (N_9165,N_8712,N_8546);
and U9166 (N_9166,N_8760,N_8629);
nand U9167 (N_9167,N_8230,N_8168);
nand U9168 (N_9168,N_8999,N_8756);
nand U9169 (N_9169,N_8279,N_8908);
xor U9170 (N_9170,N_8846,N_8508);
xnor U9171 (N_9171,N_8713,N_8038);
xor U9172 (N_9172,N_8781,N_8585);
and U9173 (N_9173,N_8511,N_8843);
or U9174 (N_9174,N_8865,N_8384);
nor U9175 (N_9175,N_8444,N_8214);
or U9176 (N_9176,N_8306,N_8005);
and U9177 (N_9177,N_8790,N_8792);
and U9178 (N_9178,N_8899,N_8957);
and U9179 (N_9179,N_8282,N_8802);
nand U9180 (N_9180,N_8691,N_8106);
or U9181 (N_9181,N_8462,N_8298);
and U9182 (N_9182,N_8257,N_8332);
or U9183 (N_9183,N_8540,N_8942);
nor U9184 (N_9184,N_8791,N_8998);
nand U9185 (N_9185,N_8601,N_8312);
xnor U9186 (N_9186,N_8480,N_8231);
nor U9187 (N_9187,N_8080,N_8840);
xor U9188 (N_9188,N_8977,N_8881);
or U9189 (N_9189,N_8219,N_8797);
or U9190 (N_9190,N_8670,N_8521);
and U9191 (N_9191,N_8258,N_8841);
nand U9192 (N_9192,N_8185,N_8799);
nand U9193 (N_9193,N_8190,N_8627);
or U9194 (N_9194,N_8801,N_8973);
xor U9195 (N_9195,N_8036,N_8711);
or U9196 (N_9196,N_8972,N_8930);
nand U9197 (N_9197,N_8296,N_8986);
or U9198 (N_9198,N_8415,N_8525);
nor U9199 (N_9199,N_8349,N_8600);
xnor U9200 (N_9200,N_8421,N_8928);
xor U9201 (N_9201,N_8416,N_8658);
and U9202 (N_9202,N_8388,N_8178);
xnor U9203 (N_9203,N_8813,N_8380);
and U9204 (N_9204,N_8063,N_8193);
nand U9205 (N_9205,N_8783,N_8677);
and U9206 (N_9206,N_8396,N_8098);
xnor U9207 (N_9207,N_8716,N_8739);
nor U9208 (N_9208,N_8839,N_8855);
nand U9209 (N_9209,N_8570,N_8623);
xnor U9210 (N_9210,N_8989,N_8302);
nor U9211 (N_9211,N_8861,N_8673);
or U9212 (N_9212,N_8943,N_8314);
xnor U9213 (N_9213,N_8949,N_8680);
or U9214 (N_9214,N_8325,N_8180);
and U9215 (N_9215,N_8007,N_8119);
or U9216 (N_9216,N_8835,N_8441);
xor U9217 (N_9217,N_8992,N_8714);
xor U9218 (N_9218,N_8753,N_8666);
or U9219 (N_9219,N_8621,N_8143);
nand U9220 (N_9220,N_8362,N_8309);
nand U9221 (N_9221,N_8552,N_8482);
nand U9222 (N_9222,N_8130,N_8515);
nor U9223 (N_9223,N_8281,N_8858);
and U9224 (N_9224,N_8681,N_8247);
nor U9225 (N_9225,N_8555,N_8572);
and U9226 (N_9226,N_8347,N_8447);
xnor U9227 (N_9227,N_8488,N_8701);
or U9228 (N_9228,N_8478,N_8150);
nor U9229 (N_9229,N_8196,N_8886);
xor U9230 (N_9230,N_8871,N_8475);
nand U9231 (N_9231,N_8034,N_8169);
nand U9232 (N_9232,N_8401,N_8017);
nand U9233 (N_9233,N_8726,N_8428);
xnor U9234 (N_9234,N_8344,N_8054);
xor U9235 (N_9235,N_8331,N_8081);
or U9236 (N_9236,N_8505,N_8544);
nand U9237 (N_9237,N_8153,N_8159);
nor U9238 (N_9238,N_8814,N_8534);
nor U9239 (N_9239,N_8962,N_8811);
or U9240 (N_9240,N_8883,N_8467);
nor U9241 (N_9241,N_8434,N_8200);
or U9242 (N_9242,N_8365,N_8655);
or U9243 (N_9243,N_8964,N_8271);
and U9244 (N_9244,N_8757,N_8483);
and U9245 (N_9245,N_8039,N_8960);
and U9246 (N_9246,N_8201,N_8529);
nand U9247 (N_9247,N_8599,N_8832);
or U9248 (N_9248,N_8683,N_8503);
nand U9249 (N_9249,N_8110,N_8322);
xor U9250 (N_9250,N_8492,N_8223);
xnor U9251 (N_9251,N_8287,N_8333);
and U9252 (N_9252,N_8736,N_8070);
nor U9253 (N_9253,N_8237,N_8994);
nor U9254 (N_9254,N_8720,N_8329);
xnor U9255 (N_9255,N_8777,N_8513);
and U9256 (N_9256,N_8723,N_8951);
nor U9257 (N_9257,N_8575,N_8952);
nor U9258 (N_9258,N_8538,N_8374);
nor U9259 (N_9259,N_8734,N_8284);
xnor U9260 (N_9260,N_8874,N_8265);
or U9261 (N_9261,N_8533,N_8617);
nand U9262 (N_9262,N_8527,N_8565);
xor U9263 (N_9263,N_8353,N_8499);
nor U9264 (N_9264,N_8050,N_8317);
and U9265 (N_9265,N_8198,N_8502);
nand U9266 (N_9266,N_8569,N_8308);
xor U9267 (N_9267,N_8926,N_8248);
or U9268 (N_9268,N_8553,N_8838);
or U9269 (N_9269,N_8429,N_8217);
or U9270 (N_9270,N_8163,N_8512);
nor U9271 (N_9271,N_8625,N_8717);
nand U9272 (N_9272,N_8091,N_8148);
and U9273 (N_9273,N_8073,N_8018);
nand U9274 (N_9274,N_8807,N_8220);
xor U9275 (N_9275,N_8844,N_8536);
xor U9276 (N_9276,N_8995,N_8438);
nor U9277 (N_9277,N_8778,N_8586);
and U9278 (N_9278,N_8700,N_8944);
nand U9279 (N_9279,N_8126,N_8420);
nor U9280 (N_9280,N_8404,N_8826);
and U9281 (N_9281,N_8138,N_8817);
and U9282 (N_9282,N_8558,N_8242);
nor U9283 (N_9283,N_8210,N_8976);
xnor U9284 (N_9284,N_8771,N_8491);
nand U9285 (N_9285,N_8708,N_8805);
xnor U9286 (N_9286,N_8554,N_8631);
nand U9287 (N_9287,N_8947,N_8320);
and U9288 (N_9288,N_8659,N_8626);
nand U9289 (N_9289,N_8315,N_8675);
nand U9290 (N_9290,N_8671,N_8361);
nand U9291 (N_9291,N_8501,N_8568);
xnor U9292 (N_9292,N_8519,N_8171);
nor U9293 (N_9293,N_8418,N_8722);
nand U9294 (N_9294,N_8310,N_8470);
or U9295 (N_9295,N_8996,N_8743);
nand U9296 (N_9296,N_8045,N_8637);
and U9297 (N_9297,N_8551,N_8604);
xnor U9298 (N_9298,N_8239,N_8436);
xor U9299 (N_9299,N_8616,N_8354);
xnor U9300 (N_9300,N_8238,N_8542);
and U9301 (N_9301,N_8319,N_8752);
or U9302 (N_9302,N_8833,N_8147);
xor U9303 (N_9303,N_8109,N_8465);
xor U9304 (N_9304,N_8918,N_8634);
and U9305 (N_9305,N_8530,N_8003);
and U9306 (N_9306,N_8507,N_8938);
and U9307 (N_9307,N_8695,N_8891);
or U9308 (N_9308,N_8123,N_8174);
nor U9309 (N_9309,N_8584,N_8692);
xor U9310 (N_9310,N_8615,N_8448);
xnor U9311 (N_9311,N_8274,N_8786);
nor U9312 (N_9312,N_8376,N_8645);
nor U9313 (N_9313,N_8803,N_8293);
nor U9314 (N_9314,N_8924,N_8221);
nand U9315 (N_9315,N_8917,N_8338);
or U9316 (N_9316,N_8772,N_8391);
or U9317 (N_9317,N_8763,N_8828);
xor U9318 (N_9318,N_8506,N_8046);
nor U9319 (N_9319,N_8114,N_8445);
nand U9320 (N_9320,N_8727,N_8443);
or U9321 (N_9321,N_8057,N_8055);
or U9322 (N_9322,N_8224,N_8262);
nor U9323 (N_9323,N_8571,N_8307);
xnor U9324 (N_9324,N_8761,N_8936);
nor U9325 (N_9325,N_8526,N_8935);
xnor U9326 (N_9326,N_8341,N_8906);
xor U9327 (N_9327,N_8424,N_8767);
and U9328 (N_9328,N_8044,N_8382);
and U9329 (N_9329,N_8020,N_8532);
nand U9330 (N_9330,N_8228,N_8853);
xnor U9331 (N_9331,N_8504,N_8486);
or U9332 (N_9332,N_8267,N_8866);
or U9333 (N_9333,N_8490,N_8676);
nor U9334 (N_9334,N_8661,N_8729);
nor U9335 (N_9335,N_8698,N_8288);
xnor U9336 (N_9336,N_8090,N_8592);
xor U9337 (N_9337,N_8602,N_8646);
and U9338 (N_9338,N_8199,N_8654);
nor U9339 (N_9339,N_8085,N_8707);
xor U9340 (N_9340,N_8493,N_8582);
nor U9341 (N_9341,N_8142,N_8368);
nor U9342 (N_9342,N_8787,N_8665);
nor U9343 (N_9343,N_8253,N_8732);
xor U9344 (N_9344,N_8633,N_8286);
and U9345 (N_9345,N_8062,N_8836);
or U9346 (N_9346,N_8244,N_8266);
xor U9347 (N_9347,N_8432,N_8066);
or U9348 (N_9348,N_8785,N_8580);
nand U9349 (N_9349,N_8959,N_8352);
and U9350 (N_9350,N_8300,N_8461);
nand U9351 (N_9351,N_8775,N_8162);
xor U9352 (N_9352,N_8910,N_8097);
xnor U9353 (N_9353,N_8660,N_8605);
xor U9354 (N_9354,N_8494,N_8464);
nor U9355 (N_9355,N_8229,N_8897);
xor U9356 (N_9356,N_8249,N_8395);
nor U9357 (N_9357,N_8932,N_8346);
nand U9358 (N_9358,N_8001,N_8809);
nor U9359 (N_9359,N_8022,N_8140);
xnor U9360 (N_9360,N_8203,N_8796);
xor U9361 (N_9361,N_8225,N_8750);
nor U9362 (N_9362,N_8375,N_8685);
nor U9363 (N_9363,N_8167,N_8472);
nand U9364 (N_9364,N_8862,N_8618);
and U9365 (N_9365,N_8643,N_8933);
xnor U9366 (N_9366,N_8305,N_8795);
nor U9367 (N_9367,N_8875,N_8578);
xor U9368 (N_9368,N_8987,N_8567);
nor U9369 (N_9369,N_8183,N_8983);
and U9370 (N_9370,N_8696,N_8638);
nor U9371 (N_9371,N_8912,N_8686);
or U9372 (N_9372,N_8863,N_8884);
xor U9373 (N_9373,N_8870,N_8878);
xnor U9374 (N_9374,N_8422,N_8851);
nand U9375 (N_9375,N_8514,N_8644);
xor U9376 (N_9376,N_8710,N_8822);
or U9377 (N_9377,N_8043,N_8598);
nand U9378 (N_9378,N_8364,N_8131);
nand U9379 (N_9379,N_8187,N_8311);
nor U9380 (N_9380,N_8155,N_8067);
and U9381 (N_9381,N_8358,N_8260);
nor U9382 (N_9382,N_8961,N_8151);
xnor U9383 (N_9383,N_8425,N_8373);
nor U9384 (N_9384,N_8072,N_8327);
xor U9385 (N_9385,N_8222,N_8888);
or U9386 (N_9386,N_8721,N_8032);
nor U9387 (N_9387,N_8121,N_8234);
nor U9388 (N_9388,N_8894,N_8133);
nand U9389 (N_9389,N_8212,N_8740);
nor U9390 (N_9390,N_8593,N_8197);
nor U9391 (N_9391,N_8277,N_8953);
and U9392 (N_9392,N_8324,N_8774);
nor U9393 (N_9393,N_8524,N_8496);
xor U9394 (N_9394,N_8789,N_8576);
and U9395 (N_9395,N_8487,N_8026);
nor U9396 (N_9396,N_8798,N_8383);
nand U9397 (N_9397,N_8405,N_8357);
or U9398 (N_9398,N_8990,N_8235);
or U9399 (N_9399,N_8816,N_8971);
nand U9400 (N_9400,N_8662,N_8549);
or U9401 (N_9401,N_8830,N_8653);
and U9402 (N_9402,N_8690,N_8719);
nor U9403 (N_9403,N_8360,N_8704);
nand U9404 (N_9404,N_8182,N_8735);
nand U9405 (N_9405,N_8509,N_8693);
nor U9406 (N_9406,N_8920,N_8651);
nand U9407 (N_9407,N_8724,N_8079);
or U9408 (N_9408,N_8845,N_8189);
nand U9409 (N_9409,N_8476,N_8784);
or U9410 (N_9410,N_8002,N_8369);
and U9411 (N_9411,N_8213,N_8904);
nor U9412 (N_9412,N_8161,N_8780);
and U9413 (N_9413,N_8181,N_8946);
or U9414 (N_9414,N_8993,N_8051);
nor U9415 (N_9415,N_8340,N_8023);
xnor U9416 (N_9416,N_8969,N_8755);
xnor U9417 (N_9417,N_8299,N_8394);
nand U9418 (N_9418,N_8965,N_8737);
xor U9419 (N_9419,N_8226,N_8083);
nor U9420 (N_9420,N_8794,N_8069);
xor U9421 (N_9421,N_8669,N_8367);
nand U9422 (N_9422,N_8218,N_8650);
or U9423 (N_9423,N_8818,N_8084);
xor U9424 (N_9424,N_8880,N_8195);
xor U9425 (N_9425,N_8980,N_8021);
or U9426 (N_9426,N_8988,N_8921);
nand U9427 (N_9427,N_8682,N_8275);
xor U9428 (N_9428,N_8419,N_8184);
nand U9429 (N_9429,N_8556,N_8837);
and U9430 (N_9430,N_8270,N_8460);
nand U9431 (N_9431,N_8510,N_8564);
or U9432 (N_9432,N_8577,N_8958);
nand U9433 (N_9433,N_8172,N_8764);
nand U9434 (N_9434,N_8074,N_8256);
xor U9435 (N_9435,N_8788,N_8408);
nand U9436 (N_9436,N_8687,N_8497);
nor U9437 (N_9437,N_8850,N_8278);
xnor U9438 (N_9438,N_8854,N_8672);
or U9439 (N_9439,N_8157,N_8453);
nor U9440 (N_9440,N_8004,N_8758);
nor U9441 (N_9441,N_8941,N_8385);
xnor U9442 (N_9442,N_8893,N_8334);
xnor U9443 (N_9443,N_8466,N_8640);
nand U9444 (N_9444,N_8145,N_8105);
xor U9445 (N_9445,N_8144,N_8979);
nor U9446 (N_9446,N_8158,N_8268);
xnor U9447 (N_9447,N_8303,N_8321);
xnor U9448 (N_9448,N_8437,N_8175);
nand U9449 (N_9449,N_8170,N_8718);
or U9450 (N_9450,N_8730,N_8204);
xnor U9451 (N_9451,N_8446,N_8635);
nor U9452 (N_9452,N_8451,N_8697);
nand U9453 (N_9453,N_8574,N_8541);
and U9454 (N_9454,N_8400,N_8092);
nand U9455 (N_9455,N_8548,N_8283);
or U9456 (N_9456,N_8948,N_8037);
nor U9457 (N_9457,N_8656,N_8543);
or U9458 (N_9458,N_8261,N_8139);
nor U9459 (N_9459,N_8956,N_8393);
nand U9460 (N_9460,N_8372,N_8093);
and U9461 (N_9461,N_8652,N_8208);
nor U9462 (N_9462,N_8164,N_8823);
nand U9463 (N_9463,N_8122,N_8477);
nand U9464 (N_9464,N_8077,N_8280);
xor U9465 (N_9465,N_8154,N_8523);
xnor U9466 (N_9466,N_8657,N_8746);
and U9467 (N_9467,N_8589,N_8856);
nor U9468 (N_9468,N_8040,N_8028);
xnor U9469 (N_9469,N_8819,N_8152);
and U9470 (N_9470,N_8251,N_8892);
and U9471 (N_9471,N_8010,N_8751);
nor U9472 (N_9472,N_8694,N_8545);
xnor U9473 (N_9473,N_8806,N_8350);
and U9474 (N_9474,N_8410,N_8603);
or U9475 (N_9475,N_8356,N_8440);
or U9476 (N_9476,N_8898,N_8120);
and U9477 (N_9477,N_8326,N_8596);
or U9478 (N_9478,N_8903,N_8149);
and U9479 (N_9479,N_8205,N_8747);
or U9480 (N_9480,N_8489,N_8378);
xnor U9481 (N_9481,N_8827,N_8108);
nand U9482 (N_9482,N_8754,N_8689);
nor U9483 (N_9483,N_8484,N_8227);
or U9484 (N_9484,N_8562,N_8810);
xnor U9485 (N_9485,N_8065,N_8699);
and U9486 (N_9486,N_8016,N_8414);
or U9487 (N_9487,N_8583,N_8520);
nor U9488 (N_9488,N_8304,N_8068);
nor U9489 (N_9489,N_8812,N_8759);
nor U9490 (N_9490,N_8087,N_8386);
or U9491 (N_9491,N_8102,N_8318);
xnor U9492 (N_9492,N_8402,N_8934);
and U9493 (N_9493,N_8009,N_8782);
or U9494 (N_9494,N_8413,N_8407);
and U9495 (N_9495,N_8590,N_8560);
and U9496 (N_9496,N_8047,N_8337);
nor U9497 (N_9497,N_8435,N_8086);
nor U9498 (N_9498,N_8071,N_8024);
or U9499 (N_9499,N_8702,N_8255);
and U9500 (N_9500,N_8448,N_8466);
xnor U9501 (N_9501,N_8691,N_8070);
or U9502 (N_9502,N_8038,N_8009);
xnor U9503 (N_9503,N_8496,N_8049);
and U9504 (N_9504,N_8037,N_8177);
and U9505 (N_9505,N_8458,N_8802);
or U9506 (N_9506,N_8340,N_8617);
or U9507 (N_9507,N_8863,N_8748);
nand U9508 (N_9508,N_8524,N_8953);
nor U9509 (N_9509,N_8643,N_8416);
and U9510 (N_9510,N_8140,N_8357);
xor U9511 (N_9511,N_8873,N_8300);
nor U9512 (N_9512,N_8967,N_8487);
or U9513 (N_9513,N_8567,N_8794);
or U9514 (N_9514,N_8035,N_8960);
and U9515 (N_9515,N_8592,N_8290);
nand U9516 (N_9516,N_8459,N_8112);
xor U9517 (N_9517,N_8965,N_8557);
and U9518 (N_9518,N_8885,N_8494);
nand U9519 (N_9519,N_8837,N_8640);
nor U9520 (N_9520,N_8126,N_8682);
nand U9521 (N_9521,N_8597,N_8668);
nand U9522 (N_9522,N_8748,N_8813);
and U9523 (N_9523,N_8265,N_8162);
nor U9524 (N_9524,N_8463,N_8706);
nand U9525 (N_9525,N_8077,N_8317);
nand U9526 (N_9526,N_8865,N_8535);
and U9527 (N_9527,N_8996,N_8371);
nor U9528 (N_9528,N_8305,N_8575);
nand U9529 (N_9529,N_8394,N_8756);
and U9530 (N_9530,N_8898,N_8794);
and U9531 (N_9531,N_8703,N_8600);
xnor U9532 (N_9532,N_8511,N_8660);
or U9533 (N_9533,N_8788,N_8572);
xnor U9534 (N_9534,N_8446,N_8372);
nand U9535 (N_9535,N_8273,N_8217);
xor U9536 (N_9536,N_8049,N_8099);
nand U9537 (N_9537,N_8141,N_8807);
nor U9538 (N_9538,N_8021,N_8440);
and U9539 (N_9539,N_8326,N_8499);
and U9540 (N_9540,N_8041,N_8732);
nand U9541 (N_9541,N_8317,N_8196);
or U9542 (N_9542,N_8148,N_8371);
or U9543 (N_9543,N_8587,N_8246);
or U9544 (N_9544,N_8913,N_8457);
or U9545 (N_9545,N_8264,N_8630);
or U9546 (N_9546,N_8552,N_8362);
or U9547 (N_9547,N_8447,N_8804);
xnor U9548 (N_9548,N_8155,N_8760);
or U9549 (N_9549,N_8474,N_8018);
or U9550 (N_9550,N_8500,N_8325);
or U9551 (N_9551,N_8443,N_8075);
nand U9552 (N_9552,N_8017,N_8740);
and U9553 (N_9553,N_8936,N_8270);
nor U9554 (N_9554,N_8107,N_8935);
and U9555 (N_9555,N_8362,N_8739);
nand U9556 (N_9556,N_8197,N_8861);
nor U9557 (N_9557,N_8481,N_8285);
nor U9558 (N_9558,N_8776,N_8663);
nand U9559 (N_9559,N_8078,N_8475);
xor U9560 (N_9560,N_8010,N_8945);
xor U9561 (N_9561,N_8420,N_8757);
xor U9562 (N_9562,N_8512,N_8149);
and U9563 (N_9563,N_8220,N_8686);
and U9564 (N_9564,N_8072,N_8816);
and U9565 (N_9565,N_8630,N_8918);
and U9566 (N_9566,N_8050,N_8222);
and U9567 (N_9567,N_8254,N_8831);
nand U9568 (N_9568,N_8714,N_8674);
nor U9569 (N_9569,N_8661,N_8573);
or U9570 (N_9570,N_8128,N_8718);
xnor U9571 (N_9571,N_8721,N_8861);
xor U9572 (N_9572,N_8788,N_8472);
xor U9573 (N_9573,N_8436,N_8232);
and U9574 (N_9574,N_8199,N_8600);
nand U9575 (N_9575,N_8402,N_8675);
nor U9576 (N_9576,N_8076,N_8817);
nor U9577 (N_9577,N_8028,N_8157);
nand U9578 (N_9578,N_8285,N_8115);
xnor U9579 (N_9579,N_8353,N_8009);
or U9580 (N_9580,N_8012,N_8690);
nor U9581 (N_9581,N_8431,N_8417);
or U9582 (N_9582,N_8495,N_8442);
nand U9583 (N_9583,N_8743,N_8311);
nand U9584 (N_9584,N_8287,N_8665);
xnor U9585 (N_9585,N_8812,N_8220);
and U9586 (N_9586,N_8016,N_8067);
xnor U9587 (N_9587,N_8015,N_8335);
and U9588 (N_9588,N_8288,N_8608);
nand U9589 (N_9589,N_8931,N_8924);
or U9590 (N_9590,N_8991,N_8809);
nand U9591 (N_9591,N_8091,N_8366);
xnor U9592 (N_9592,N_8249,N_8664);
nand U9593 (N_9593,N_8618,N_8732);
nand U9594 (N_9594,N_8967,N_8407);
nor U9595 (N_9595,N_8062,N_8245);
nor U9596 (N_9596,N_8421,N_8039);
nand U9597 (N_9597,N_8429,N_8644);
and U9598 (N_9598,N_8651,N_8770);
nand U9599 (N_9599,N_8647,N_8821);
or U9600 (N_9600,N_8592,N_8195);
nor U9601 (N_9601,N_8585,N_8691);
nand U9602 (N_9602,N_8467,N_8562);
or U9603 (N_9603,N_8944,N_8396);
and U9604 (N_9604,N_8309,N_8186);
and U9605 (N_9605,N_8255,N_8096);
xor U9606 (N_9606,N_8766,N_8499);
xor U9607 (N_9607,N_8291,N_8725);
xor U9608 (N_9608,N_8454,N_8503);
xnor U9609 (N_9609,N_8274,N_8122);
nand U9610 (N_9610,N_8345,N_8833);
xor U9611 (N_9611,N_8555,N_8827);
nor U9612 (N_9612,N_8820,N_8687);
xor U9613 (N_9613,N_8004,N_8479);
nor U9614 (N_9614,N_8140,N_8480);
nand U9615 (N_9615,N_8143,N_8050);
nor U9616 (N_9616,N_8949,N_8718);
nand U9617 (N_9617,N_8801,N_8734);
and U9618 (N_9618,N_8393,N_8976);
nand U9619 (N_9619,N_8651,N_8870);
xnor U9620 (N_9620,N_8673,N_8816);
and U9621 (N_9621,N_8297,N_8160);
nand U9622 (N_9622,N_8636,N_8455);
xor U9623 (N_9623,N_8178,N_8503);
nor U9624 (N_9624,N_8400,N_8435);
nor U9625 (N_9625,N_8870,N_8486);
xor U9626 (N_9626,N_8405,N_8421);
and U9627 (N_9627,N_8949,N_8115);
or U9628 (N_9628,N_8104,N_8722);
xnor U9629 (N_9629,N_8780,N_8597);
nand U9630 (N_9630,N_8664,N_8867);
and U9631 (N_9631,N_8875,N_8720);
and U9632 (N_9632,N_8587,N_8697);
nor U9633 (N_9633,N_8950,N_8970);
and U9634 (N_9634,N_8432,N_8627);
or U9635 (N_9635,N_8770,N_8366);
or U9636 (N_9636,N_8745,N_8317);
nor U9637 (N_9637,N_8502,N_8210);
xnor U9638 (N_9638,N_8469,N_8292);
nand U9639 (N_9639,N_8763,N_8143);
or U9640 (N_9640,N_8603,N_8787);
or U9641 (N_9641,N_8154,N_8054);
nor U9642 (N_9642,N_8517,N_8561);
and U9643 (N_9643,N_8945,N_8773);
nand U9644 (N_9644,N_8620,N_8441);
nand U9645 (N_9645,N_8789,N_8612);
or U9646 (N_9646,N_8781,N_8307);
and U9647 (N_9647,N_8224,N_8568);
or U9648 (N_9648,N_8485,N_8190);
or U9649 (N_9649,N_8826,N_8824);
xor U9650 (N_9650,N_8737,N_8625);
or U9651 (N_9651,N_8734,N_8051);
nor U9652 (N_9652,N_8386,N_8055);
nor U9653 (N_9653,N_8105,N_8442);
and U9654 (N_9654,N_8814,N_8564);
nor U9655 (N_9655,N_8145,N_8192);
xnor U9656 (N_9656,N_8551,N_8117);
xnor U9657 (N_9657,N_8873,N_8328);
or U9658 (N_9658,N_8071,N_8215);
and U9659 (N_9659,N_8214,N_8398);
xnor U9660 (N_9660,N_8379,N_8224);
and U9661 (N_9661,N_8839,N_8879);
nor U9662 (N_9662,N_8780,N_8103);
xnor U9663 (N_9663,N_8746,N_8563);
and U9664 (N_9664,N_8441,N_8243);
nor U9665 (N_9665,N_8399,N_8590);
or U9666 (N_9666,N_8037,N_8689);
xnor U9667 (N_9667,N_8137,N_8792);
nand U9668 (N_9668,N_8561,N_8411);
nor U9669 (N_9669,N_8661,N_8603);
and U9670 (N_9670,N_8415,N_8953);
nand U9671 (N_9671,N_8807,N_8354);
nor U9672 (N_9672,N_8994,N_8805);
nor U9673 (N_9673,N_8634,N_8833);
xnor U9674 (N_9674,N_8979,N_8449);
nor U9675 (N_9675,N_8704,N_8330);
nand U9676 (N_9676,N_8703,N_8524);
and U9677 (N_9677,N_8572,N_8917);
or U9678 (N_9678,N_8656,N_8824);
xnor U9679 (N_9679,N_8455,N_8265);
nor U9680 (N_9680,N_8437,N_8177);
or U9681 (N_9681,N_8611,N_8107);
or U9682 (N_9682,N_8156,N_8682);
and U9683 (N_9683,N_8650,N_8829);
and U9684 (N_9684,N_8825,N_8083);
and U9685 (N_9685,N_8324,N_8222);
nand U9686 (N_9686,N_8558,N_8388);
or U9687 (N_9687,N_8243,N_8772);
or U9688 (N_9688,N_8942,N_8400);
nand U9689 (N_9689,N_8372,N_8674);
nand U9690 (N_9690,N_8471,N_8272);
and U9691 (N_9691,N_8882,N_8546);
xor U9692 (N_9692,N_8014,N_8082);
xor U9693 (N_9693,N_8810,N_8428);
and U9694 (N_9694,N_8066,N_8456);
xnor U9695 (N_9695,N_8413,N_8129);
nor U9696 (N_9696,N_8114,N_8329);
nor U9697 (N_9697,N_8070,N_8636);
xnor U9698 (N_9698,N_8796,N_8464);
nand U9699 (N_9699,N_8684,N_8035);
and U9700 (N_9700,N_8100,N_8745);
nand U9701 (N_9701,N_8541,N_8716);
xor U9702 (N_9702,N_8201,N_8774);
nand U9703 (N_9703,N_8664,N_8848);
xnor U9704 (N_9704,N_8462,N_8156);
or U9705 (N_9705,N_8907,N_8588);
xnor U9706 (N_9706,N_8398,N_8506);
and U9707 (N_9707,N_8765,N_8649);
and U9708 (N_9708,N_8459,N_8077);
xnor U9709 (N_9709,N_8799,N_8706);
nand U9710 (N_9710,N_8881,N_8420);
and U9711 (N_9711,N_8585,N_8436);
and U9712 (N_9712,N_8289,N_8097);
nor U9713 (N_9713,N_8218,N_8502);
and U9714 (N_9714,N_8268,N_8041);
nor U9715 (N_9715,N_8354,N_8364);
xor U9716 (N_9716,N_8891,N_8056);
nor U9717 (N_9717,N_8334,N_8993);
and U9718 (N_9718,N_8044,N_8808);
or U9719 (N_9719,N_8476,N_8666);
nor U9720 (N_9720,N_8302,N_8482);
xor U9721 (N_9721,N_8984,N_8003);
nor U9722 (N_9722,N_8777,N_8945);
or U9723 (N_9723,N_8570,N_8000);
nor U9724 (N_9724,N_8320,N_8120);
and U9725 (N_9725,N_8507,N_8033);
nand U9726 (N_9726,N_8445,N_8975);
or U9727 (N_9727,N_8856,N_8280);
nor U9728 (N_9728,N_8827,N_8700);
nand U9729 (N_9729,N_8263,N_8456);
xnor U9730 (N_9730,N_8374,N_8748);
xor U9731 (N_9731,N_8850,N_8162);
xnor U9732 (N_9732,N_8842,N_8044);
nor U9733 (N_9733,N_8635,N_8943);
nor U9734 (N_9734,N_8815,N_8990);
xnor U9735 (N_9735,N_8779,N_8908);
xnor U9736 (N_9736,N_8909,N_8917);
nand U9737 (N_9737,N_8814,N_8533);
nand U9738 (N_9738,N_8733,N_8752);
nor U9739 (N_9739,N_8277,N_8543);
nand U9740 (N_9740,N_8001,N_8804);
xnor U9741 (N_9741,N_8532,N_8247);
nand U9742 (N_9742,N_8292,N_8706);
xnor U9743 (N_9743,N_8910,N_8804);
nand U9744 (N_9744,N_8297,N_8961);
nand U9745 (N_9745,N_8939,N_8850);
nor U9746 (N_9746,N_8233,N_8926);
and U9747 (N_9747,N_8084,N_8000);
and U9748 (N_9748,N_8652,N_8073);
xnor U9749 (N_9749,N_8590,N_8964);
xor U9750 (N_9750,N_8772,N_8382);
and U9751 (N_9751,N_8979,N_8390);
and U9752 (N_9752,N_8011,N_8532);
xor U9753 (N_9753,N_8386,N_8222);
nand U9754 (N_9754,N_8545,N_8935);
nor U9755 (N_9755,N_8985,N_8907);
xor U9756 (N_9756,N_8037,N_8798);
or U9757 (N_9757,N_8210,N_8646);
nor U9758 (N_9758,N_8634,N_8832);
xor U9759 (N_9759,N_8371,N_8180);
xnor U9760 (N_9760,N_8339,N_8891);
or U9761 (N_9761,N_8838,N_8013);
nand U9762 (N_9762,N_8172,N_8463);
and U9763 (N_9763,N_8076,N_8951);
xor U9764 (N_9764,N_8342,N_8306);
nand U9765 (N_9765,N_8601,N_8385);
xnor U9766 (N_9766,N_8363,N_8429);
and U9767 (N_9767,N_8726,N_8153);
nor U9768 (N_9768,N_8365,N_8530);
nand U9769 (N_9769,N_8032,N_8014);
or U9770 (N_9770,N_8209,N_8737);
or U9771 (N_9771,N_8291,N_8794);
nand U9772 (N_9772,N_8857,N_8388);
nor U9773 (N_9773,N_8330,N_8216);
and U9774 (N_9774,N_8190,N_8777);
nand U9775 (N_9775,N_8155,N_8200);
xor U9776 (N_9776,N_8397,N_8935);
nand U9777 (N_9777,N_8039,N_8625);
or U9778 (N_9778,N_8698,N_8891);
nand U9779 (N_9779,N_8500,N_8718);
nand U9780 (N_9780,N_8098,N_8554);
nor U9781 (N_9781,N_8137,N_8172);
nand U9782 (N_9782,N_8508,N_8443);
nand U9783 (N_9783,N_8281,N_8189);
nor U9784 (N_9784,N_8839,N_8847);
nor U9785 (N_9785,N_8172,N_8856);
xor U9786 (N_9786,N_8632,N_8941);
nand U9787 (N_9787,N_8883,N_8177);
or U9788 (N_9788,N_8528,N_8041);
nand U9789 (N_9789,N_8971,N_8889);
xnor U9790 (N_9790,N_8113,N_8562);
nor U9791 (N_9791,N_8999,N_8267);
or U9792 (N_9792,N_8658,N_8618);
and U9793 (N_9793,N_8966,N_8131);
nor U9794 (N_9794,N_8391,N_8958);
nand U9795 (N_9795,N_8291,N_8066);
xor U9796 (N_9796,N_8822,N_8169);
nor U9797 (N_9797,N_8444,N_8250);
nor U9798 (N_9798,N_8823,N_8639);
or U9799 (N_9799,N_8966,N_8107);
xor U9800 (N_9800,N_8115,N_8292);
or U9801 (N_9801,N_8484,N_8375);
or U9802 (N_9802,N_8748,N_8841);
nor U9803 (N_9803,N_8320,N_8707);
xor U9804 (N_9804,N_8258,N_8095);
nor U9805 (N_9805,N_8189,N_8294);
xor U9806 (N_9806,N_8532,N_8762);
and U9807 (N_9807,N_8020,N_8763);
nand U9808 (N_9808,N_8850,N_8878);
xor U9809 (N_9809,N_8577,N_8225);
or U9810 (N_9810,N_8986,N_8969);
and U9811 (N_9811,N_8007,N_8864);
nor U9812 (N_9812,N_8844,N_8819);
and U9813 (N_9813,N_8860,N_8884);
or U9814 (N_9814,N_8217,N_8839);
nor U9815 (N_9815,N_8486,N_8152);
nand U9816 (N_9816,N_8087,N_8416);
nand U9817 (N_9817,N_8027,N_8894);
and U9818 (N_9818,N_8692,N_8102);
and U9819 (N_9819,N_8872,N_8066);
and U9820 (N_9820,N_8115,N_8948);
or U9821 (N_9821,N_8551,N_8171);
and U9822 (N_9822,N_8237,N_8474);
and U9823 (N_9823,N_8714,N_8237);
or U9824 (N_9824,N_8270,N_8421);
nand U9825 (N_9825,N_8919,N_8847);
and U9826 (N_9826,N_8315,N_8402);
xor U9827 (N_9827,N_8831,N_8274);
or U9828 (N_9828,N_8022,N_8277);
or U9829 (N_9829,N_8494,N_8378);
and U9830 (N_9830,N_8854,N_8138);
and U9831 (N_9831,N_8892,N_8291);
or U9832 (N_9832,N_8952,N_8980);
or U9833 (N_9833,N_8638,N_8392);
nor U9834 (N_9834,N_8571,N_8505);
nor U9835 (N_9835,N_8918,N_8554);
nor U9836 (N_9836,N_8338,N_8138);
nor U9837 (N_9837,N_8141,N_8279);
nand U9838 (N_9838,N_8825,N_8778);
and U9839 (N_9839,N_8188,N_8751);
nor U9840 (N_9840,N_8542,N_8791);
xnor U9841 (N_9841,N_8840,N_8348);
or U9842 (N_9842,N_8095,N_8544);
or U9843 (N_9843,N_8576,N_8902);
and U9844 (N_9844,N_8713,N_8826);
nor U9845 (N_9845,N_8297,N_8335);
or U9846 (N_9846,N_8959,N_8455);
nor U9847 (N_9847,N_8452,N_8410);
and U9848 (N_9848,N_8916,N_8909);
nor U9849 (N_9849,N_8796,N_8024);
or U9850 (N_9850,N_8418,N_8463);
nor U9851 (N_9851,N_8995,N_8609);
nand U9852 (N_9852,N_8319,N_8435);
and U9853 (N_9853,N_8280,N_8417);
xnor U9854 (N_9854,N_8609,N_8603);
or U9855 (N_9855,N_8971,N_8473);
nand U9856 (N_9856,N_8379,N_8981);
or U9857 (N_9857,N_8872,N_8125);
nor U9858 (N_9858,N_8559,N_8794);
nand U9859 (N_9859,N_8331,N_8874);
and U9860 (N_9860,N_8639,N_8348);
xnor U9861 (N_9861,N_8293,N_8315);
xor U9862 (N_9862,N_8812,N_8967);
nand U9863 (N_9863,N_8902,N_8968);
nor U9864 (N_9864,N_8609,N_8393);
and U9865 (N_9865,N_8620,N_8016);
nor U9866 (N_9866,N_8264,N_8891);
xnor U9867 (N_9867,N_8300,N_8997);
or U9868 (N_9868,N_8631,N_8044);
and U9869 (N_9869,N_8271,N_8723);
nor U9870 (N_9870,N_8547,N_8546);
or U9871 (N_9871,N_8187,N_8839);
or U9872 (N_9872,N_8537,N_8071);
and U9873 (N_9873,N_8421,N_8021);
xnor U9874 (N_9874,N_8661,N_8293);
xor U9875 (N_9875,N_8133,N_8109);
or U9876 (N_9876,N_8639,N_8265);
and U9877 (N_9877,N_8749,N_8414);
nand U9878 (N_9878,N_8135,N_8678);
xnor U9879 (N_9879,N_8767,N_8911);
nor U9880 (N_9880,N_8608,N_8306);
nor U9881 (N_9881,N_8942,N_8127);
nor U9882 (N_9882,N_8823,N_8873);
xor U9883 (N_9883,N_8029,N_8622);
nand U9884 (N_9884,N_8534,N_8964);
or U9885 (N_9885,N_8123,N_8716);
nand U9886 (N_9886,N_8458,N_8951);
xnor U9887 (N_9887,N_8351,N_8252);
and U9888 (N_9888,N_8377,N_8065);
or U9889 (N_9889,N_8891,N_8964);
or U9890 (N_9890,N_8857,N_8939);
and U9891 (N_9891,N_8402,N_8854);
or U9892 (N_9892,N_8678,N_8731);
xor U9893 (N_9893,N_8883,N_8602);
or U9894 (N_9894,N_8417,N_8483);
and U9895 (N_9895,N_8498,N_8678);
and U9896 (N_9896,N_8889,N_8043);
nand U9897 (N_9897,N_8711,N_8559);
or U9898 (N_9898,N_8601,N_8231);
nor U9899 (N_9899,N_8708,N_8866);
or U9900 (N_9900,N_8677,N_8225);
nor U9901 (N_9901,N_8188,N_8190);
or U9902 (N_9902,N_8837,N_8168);
or U9903 (N_9903,N_8435,N_8909);
and U9904 (N_9904,N_8096,N_8344);
nor U9905 (N_9905,N_8382,N_8226);
or U9906 (N_9906,N_8048,N_8166);
nand U9907 (N_9907,N_8295,N_8159);
nor U9908 (N_9908,N_8736,N_8981);
nor U9909 (N_9909,N_8667,N_8462);
nor U9910 (N_9910,N_8839,N_8351);
nor U9911 (N_9911,N_8863,N_8197);
xor U9912 (N_9912,N_8350,N_8436);
nor U9913 (N_9913,N_8112,N_8912);
nand U9914 (N_9914,N_8848,N_8288);
nor U9915 (N_9915,N_8637,N_8280);
nand U9916 (N_9916,N_8776,N_8726);
or U9917 (N_9917,N_8975,N_8149);
nor U9918 (N_9918,N_8242,N_8534);
nand U9919 (N_9919,N_8186,N_8120);
and U9920 (N_9920,N_8279,N_8669);
nor U9921 (N_9921,N_8922,N_8053);
or U9922 (N_9922,N_8972,N_8950);
and U9923 (N_9923,N_8950,N_8848);
nor U9924 (N_9924,N_8048,N_8382);
and U9925 (N_9925,N_8903,N_8942);
and U9926 (N_9926,N_8633,N_8544);
and U9927 (N_9927,N_8358,N_8574);
nor U9928 (N_9928,N_8583,N_8207);
nor U9929 (N_9929,N_8824,N_8112);
and U9930 (N_9930,N_8295,N_8968);
xor U9931 (N_9931,N_8748,N_8567);
nand U9932 (N_9932,N_8243,N_8193);
or U9933 (N_9933,N_8538,N_8585);
nor U9934 (N_9934,N_8878,N_8481);
or U9935 (N_9935,N_8343,N_8615);
or U9936 (N_9936,N_8302,N_8631);
and U9937 (N_9937,N_8092,N_8746);
nor U9938 (N_9938,N_8631,N_8984);
and U9939 (N_9939,N_8892,N_8678);
nand U9940 (N_9940,N_8169,N_8013);
or U9941 (N_9941,N_8631,N_8893);
nor U9942 (N_9942,N_8186,N_8957);
nand U9943 (N_9943,N_8994,N_8139);
xnor U9944 (N_9944,N_8587,N_8814);
nand U9945 (N_9945,N_8823,N_8991);
nand U9946 (N_9946,N_8453,N_8974);
and U9947 (N_9947,N_8587,N_8797);
nand U9948 (N_9948,N_8581,N_8985);
and U9949 (N_9949,N_8486,N_8957);
and U9950 (N_9950,N_8281,N_8272);
or U9951 (N_9951,N_8959,N_8166);
nor U9952 (N_9952,N_8163,N_8613);
xnor U9953 (N_9953,N_8191,N_8920);
nor U9954 (N_9954,N_8779,N_8438);
xor U9955 (N_9955,N_8937,N_8239);
or U9956 (N_9956,N_8757,N_8101);
and U9957 (N_9957,N_8123,N_8508);
or U9958 (N_9958,N_8120,N_8178);
nor U9959 (N_9959,N_8696,N_8684);
nand U9960 (N_9960,N_8491,N_8908);
or U9961 (N_9961,N_8359,N_8583);
nand U9962 (N_9962,N_8285,N_8042);
nor U9963 (N_9963,N_8889,N_8798);
and U9964 (N_9964,N_8135,N_8576);
nor U9965 (N_9965,N_8691,N_8767);
xnor U9966 (N_9966,N_8816,N_8502);
or U9967 (N_9967,N_8268,N_8542);
xor U9968 (N_9968,N_8627,N_8936);
and U9969 (N_9969,N_8663,N_8082);
or U9970 (N_9970,N_8795,N_8660);
or U9971 (N_9971,N_8042,N_8184);
and U9972 (N_9972,N_8454,N_8487);
xnor U9973 (N_9973,N_8497,N_8816);
nor U9974 (N_9974,N_8602,N_8176);
or U9975 (N_9975,N_8272,N_8176);
nand U9976 (N_9976,N_8088,N_8245);
and U9977 (N_9977,N_8704,N_8865);
and U9978 (N_9978,N_8226,N_8314);
nand U9979 (N_9979,N_8028,N_8413);
nand U9980 (N_9980,N_8309,N_8092);
nor U9981 (N_9981,N_8431,N_8966);
xnor U9982 (N_9982,N_8740,N_8346);
and U9983 (N_9983,N_8683,N_8132);
nand U9984 (N_9984,N_8640,N_8915);
nor U9985 (N_9985,N_8932,N_8634);
or U9986 (N_9986,N_8422,N_8955);
xnor U9987 (N_9987,N_8115,N_8746);
xnor U9988 (N_9988,N_8951,N_8364);
nor U9989 (N_9989,N_8718,N_8674);
or U9990 (N_9990,N_8602,N_8205);
xor U9991 (N_9991,N_8357,N_8708);
nand U9992 (N_9992,N_8766,N_8429);
nor U9993 (N_9993,N_8350,N_8170);
and U9994 (N_9994,N_8438,N_8906);
and U9995 (N_9995,N_8836,N_8701);
nand U9996 (N_9996,N_8990,N_8610);
nand U9997 (N_9997,N_8556,N_8772);
and U9998 (N_9998,N_8939,N_8345);
or U9999 (N_9999,N_8841,N_8120);
xnor U10000 (N_10000,N_9277,N_9226);
nand U10001 (N_10001,N_9938,N_9025);
nor U10002 (N_10002,N_9154,N_9906);
xor U10003 (N_10003,N_9323,N_9376);
or U10004 (N_10004,N_9197,N_9644);
nor U10005 (N_10005,N_9517,N_9211);
nor U10006 (N_10006,N_9045,N_9335);
and U10007 (N_10007,N_9032,N_9426);
and U10008 (N_10008,N_9996,N_9676);
nor U10009 (N_10009,N_9221,N_9178);
nor U10010 (N_10010,N_9368,N_9217);
or U10011 (N_10011,N_9546,N_9822);
and U10012 (N_10012,N_9340,N_9412);
nand U10013 (N_10013,N_9894,N_9188);
xnor U10014 (N_10014,N_9717,N_9963);
nor U10015 (N_10015,N_9504,N_9862);
and U10016 (N_10016,N_9556,N_9236);
xnor U10017 (N_10017,N_9258,N_9400);
and U10018 (N_10018,N_9776,N_9849);
nor U10019 (N_10019,N_9878,N_9633);
or U10020 (N_10020,N_9010,N_9165);
xnor U10021 (N_10021,N_9840,N_9251);
or U10022 (N_10022,N_9626,N_9692);
xnor U10023 (N_10023,N_9103,N_9986);
xor U10024 (N_10024,N_9471,N_9017);
or U10025 (N_10025,N_9509,N_9716);
nor U10026 (N_10026,N_9729,N_9027);
or U10027 (N_10027,N_9179,N_9681);
xor U10028 (N_10028,N_9508,N_9072);
nor U10029 (N_10029,N_9555,N_9111);
xnor U10030 (N_10030,N_9638,N_9263);
nor U10031 (N_10031,N_9587,N_9004);
xor U10032 (N_10032,N_9430,N_9930);
or U10033 (N_10033,N_9389,N_9558);
or U10034 (N_10034,N_9553,N_9466);
xor U10035 (N_10035,N_9199,N_9428);
xor U10036 (N_10036,N_9708,N_9808);
nor U10037 (N_10037,N_9629,N_9053);
and U10038 (N_10038,N_9722,N_9015);
nand U10039 (N_10039,N_9564,N_9177);
and U10040 (N_10040,N_9078,N_9614);
and U10041 (N_10041,N_9102,N_9084);
or U10042 (N_10042,N_9715,N_9521);
and U10043 (N_10043,N_9486,N_9700);
and U10044 (N_10044,N_9668,N_9268);
xnor U10045 (N_10045,N_9750,N_9924);
nand U10046 (N_10046,N_9185,N_9462);
nor U10047 (N_10047,N_9275,N_9020);
nand U10048 (N_10048,N_9397,N_9040);
and U10049 (N_10049,N_9813,N_9636);
nor U10050 (N_10050,N_9173,N_9175);
or U10051 (N_10051,N_9460,N_9190);
xor U10052 (N_10052,N_9921,N_9818);
xor U10053 (N_10053,N_9519,N_9588);
and U10054 (N_10054,N_9195,N_9186);
xor U10055 (N_10055,N_9227,N_9828);
nor U10056 (N_10056,N_9007,N_9745);
and U10057 (N_10057,N_9654,N_9893);
nand U10058 (N_10058,N_9671,N_9884);
xnor U10059 (N_10059,N_9002,N_9161);
or U10060 (N_10060,N_9413,N_9094);
or U10061 (N_10061,N_9077,N_9838);
and U10062 (N_10062,N_9615,N_9892);
nand U10063 (N_10063,N_9435,N_9312);
nor U10064 (N_10064,N_9507,N_9203);
or U10065 (N_10065,N_9730,N_9087);
nand U10066 (N_10066,N_9839,N_9837);
nand U10067 (N_10067,N_9667,N_9575);
nand U10068 (N_10068,N_9806,N_9794);
and U10069 (N_10069,N_9993,N_9887);
nand U10070 (N_10070,N_9324,N_9765);
nor U10071 (N_10071,N_9542,N_9797);
xor U10072 (N_10072,N_9239,N_9176);
nor U10073 (N_10073,N_9992,N_9696);
nand U10074 (N_10074,N_9751,N_9309);
and U10075 (N_10075,N_9600,N_9968);
nand U10076 (N_10076,N_9721,N_9461);
or U10077 (N_10077,N_9130,N_9689);
and U10078 (N_10078,N_9207,N_9115);
and U10079 (N_10079,N_9364,N_9448);
nand U10080 (N_10080,N_9018,N_9550);
xor U10081 (N_10081,N_9138,N_9945);
or U10082 (N_10082,N_9349,N_9695);
nand U10083 (N_10083,N_9650,N_9476);
xor U10084 (N_10084,N_9999,N_9387);
or U10085 (N_10085,N_9854,N_9089);
or U10086 (N_10086,N_9363,N_9757);
or U10087 (N_10087,N_9423,N_9889);
or U10088 (N_10088,N_9358,N_9116);
nand U10089 (N_10089,N_9863,N_9422);
nor U10090 (N_10090,N_9622,N_9901);
nand U10091 (N_10091,N_9562,N_9779);
and U10092 (N_10092,N_9909,N_9286);
or U10093 (N_10093,N_9752,N_9080);
nor U10094 (N_10094,N_9578,N_9143);
nor U10095 (N_10095,N_9260,N_9058);
nor U10096 (N_10096,N_9810,N_9005);
and U10097 (N_10097,N_9569,N_9557);
or U10098 (N_10098,N_9725,N_9408);
xnor U10099 (N_10099,N_9665,N_9494);
and U10100 (N_10100,N_9705,N_9441);
nand U10101 (N_10101,N_9361,N_9811);
xnor U10102 (N_10102,N_9383,N_9118);
nor U10103 (N_10103,N_9060,N_9153);
and U10104 (N_10104,N_9381,N_9497);
nand U10105 (N_10105,N_9657,N_9308);
xor U10106 (N_10106,N_9613,N_9157);
nor U10107 (N_10107,N_9595,N_9880);
xor U10108 (N_10108,N_9205,N_9835);
and U10109 (N_10109,N_9534,N_9604);
nor U10110 (N_10110,N_9997,N_9000);
or U10111 (N_10111,N_9307,N_9821);
xnor U10112 (N_10112,N_9784,N_9451);
nor U10113 (N_10113,N_9233,N_9908);
nor U10114 (N_10114,N_9474,N_9473);
xnor U10115 (N_10115,N_9971,N_9617);
nor U10116 (N_10116,N_9951,N_9257);
and U10117 (N_10117,N_9946,N_9455);
and U10118 (N_10118,N_9867,N_9888);
or U10119 (N_10119,N_9127,N_9287);
nand U10120 (N_10120,N_9651,N_9823);
and U10121 (N_10121,N_9647,N_9314);
nor U10122 (N_10122,N_9998,N_9360);
or U10123 (N_10123,N_9772,N_9687);
or U10124 (N_10124,N_9061,N_9649);
nand U10125 (N_10125,N_9911,N_9510);
and U10126 (N_10126,N_9490,N_9431);
or U10127 (N_10127,N_9146,N_9660);
nor U10128 (N_10128,N_9276,N_9182);
or U10129 (N_10129,N_9516,N_9628);
xor U10130 (N_10130,N_9741,N_9799);
nor U10131 (N_10131,N_9869,N_9142);
xor U10132 (N_10132,N_9573,N_9560);
nor U10133 (N_10133,N_9978,N_9068);
or U10134 (N_10134,N_9278,N_9805);
or U10135 (N_10135,N_9602,N_9082);
or U10136 (N_10136,N_9902,N_9382);
and U10137 (N_10137,N_9230,N_9552);
xor U10138 (N_10138,N_9913,N_9975);
and U10139 (N_10139,N_9044,N_9261);
and U10140 (N_10140,N_9538,N_9104);
nand U10141 (N_10141,N_9265,N_9062);
nand U10142 (N_10142,N_9073,N_9145);
nor U10143 (N_10143,N_9694,N_9229);
nand U10144 (N_10144,N_9088,N_9762);
and U10145 (N_10145,N_9707,N_9531);
or U10146 (N_10146,N_9955,N_9591);
nand U10147 (N_10147,N_9270,N_9895);
or U10148 (N_10148,N_9498,N_9661);
and U10149 (N_10149,N_9882,N_9488);
nand U10150 (N_10150,N_9789,N_9155);
nor U10151 (N_10151,N_9576,N_9281);
xor U10152 (N_10152,N_9350,N_9656);
nor U10153 (N_10153,N_9738,N_9592);
xnor U10154 (N_10154,N_9320,N_9989);
nand U10155 (N_10155,N_9329,N_9874);
or U10156 (N_10156,N_9965,N_9401);
and U10157 (N_10157,N_9450,N_9150);
xor U10158 (N_10158,N_9006,N_9876);
nand U10159 (N_10159,N_9559,N_9362);
nand U10160 (N_10160,N_9995,N_9758);
and U10161 (N_10161,N_9056,N_9480);
and U10162 (N_10162,N_9711,N_9332);
nand U10163 (N_10163,N_9063,N_9561);
or U10164 (N_10164,N_9926,N_9873);
xnor U10165 (N_10165,N_9599,N_9310);
or U10166 (N_10166,N_9643,N_9174);
nor U10167 (N_10167,N_9790,N_9123);
xor U10168 (N_10168,N_9013,N_9343);
and U10169 (N_10169,N_9030,N_9583);
or U10170 (N_10170,N_9054,N_9528);
nor U10171 (N_10171,N_9446,N_9706);
nand U10172 (N_10172,N_9424,N_9345);
or U10173 (N_10173,N_9632,N_9033);
xor U10174 (N_10174,N_9537,N_9303);
and U10175 (N_10175,N_9411,N_9704);
and U10176 (N_10176,N_9927,N_9843);
and U10177 (N_10177,N_9481,N_9608);
or U10178 (N_10178,N_9781,N_9680);
xnor U10179 (N_10179,N_9934,N_9658);
or U10180 (N_10180,N_9929,N_9917);
nor U10181 (N_10181,N_9204,N_9634);
nand U10182 (N_10182,N_9742,N_9305);
or U10183 (N_10183,N_9645,N_9213);
nor U10184 (N_10184,N_9904,N_9825);
and U10185 (N_10185,N_9067,N_9817);
xor U10186 (N_10186,N_9394,N_9131);
and U10187 (N_10187,N_9845,N_9269);
or U10188 (N_10188,N_9607,N_9732);
xor U10189 (N_10189,N_9041,N_9983);
nor U10190 (N_10190,N_9941,N_9520);
xnor U10191 (N_10191,N_9379,N_9686);
nand U10192 (N_10192,N_9120,N_9390);
xor U10193 (N_10193,N_9731,N_9183);
nand U10194 (N_10194,N_9452,N_9306);
and U10195 (N_10195,N_9141,N_9442);
nand U10196 (N_10196,N_9726,N_9565);
nor U10197 (N_10197,N_9864,N_9812);
xnor U10198 (N_10198,N_9271,N_9858);
or U10199 (N_10199,N_9091,N_9284);
and U10200 (N_10200,N_9099,N_9948);
and U10201 (N_10201,N_9853,N_9279);
xor U10202 (N_10202,N_9727,N_9831);
nor U10203 (N_10203,N_9372,N_9655);
and U10204 (N_10204,N_9219,N_9495);
nand U10205 (N_10205,N_9833,N_9639);
xor U10206 (N_10206,N_9851,N_9697);
and U10207 (N_10207,N_9386,N_9107);
nand U10208 (N_10208,N_9266,N_9684);
or U10209 (N_10209,N_9807,N_9189);
or U10210 (N_10210,N_9896,N_9566);
and U10211 (N_10211,N_9682,N_9767);
xor U10212 (N_10212,N_9855,N_9815);
nor U10213 (N_10213,N_9148,N_9981);
nor U10214 (N_10214,N_9974,N_9919);
xnor U10215 (N_10215,N_9167,N_9406);
nand U10216 (N_10216,N_9014,N_9404);
nand U10217 (N_10217,N_9168,N_9949);
nand U10218 (N_10218,N_9250,N_9871);
or U10219 (N_10219,N_9011,N_9693);
nor U10220 (N_10220,N_9128,N_9283);
or U10221 (N_10221,N_9513,N_9976);
nand U10222 (N_10222,N_9191,N_9137);
nand U10223 (N_10223,N_9834,N_9786);
or U10224 (N_10224,N_9097,N_9366);
and U10225 (N_10225,N_9016,N_9957);
nand U10226 (N_10226,N_9961,N_9605);
nor U10227 (N_10227,N_9770,N_9803);
nor U10228 (N_10228,N_9581,N_9222);
or U10229 (N_10229,N_9187,N_9610);
nor U10230 (N_10230,N_9021,N_9761);
xor U10231 (N_10231,N_9549,N_9527);
or U10232 (N_10232,N_9532,N_9551);
xnor U10233 (N_10233,N_9457,N_9967);
nor U10234 (N_10234,N_9046,N_9105);
or U10235 (N_10235,N_9209,N_9859);
and U10236 (N_10236,N_9856,N_9925);
nand U10237 (N_10237,N_9392,N_9749);
nand U10238 (N_10238,N_9313,N_9857);
or U10239 (N_10239,N_9365,N_9539);
nand U10240 (N_10240,N_9210,N_9031);
and U10241 (N_10241,N_9733,N_9900);
or U10242 (N_10242,N_9380,N_9456);
and U10243 (N_10243,N_9641,N_9234);
and U10244 (N_10244,N_9954,N_9415);
nand U10245 (N_10245,N_9136,N_9915);
nand U10246 (N_10246,N_9347,N_9586);
nand U10247 (N_10247,N_9870,N_9069);
xnor U10248 (N_10248,N_9920,N_9228);
nor U10249 (N_10249,N_9619,N_9095);
nor U10250 (N_10250,N_9254,N_9543);
or U10251 (N_10251,N_9029,N_9800);
and U10252 (N_10252,N_9296,N_9417);
xnor U10253 (N_10253,N_9410,N_9375);
nor U10254 (N_10254,N_9724,N_9117);
xnor U10255 (N_10255,N_9096,N_9756);
xor U10256 (N_10256,N_9215,N_9964);
nor U10257 (N_10257,N_9454,N_9568);
nor U10258 (N_10258,N_9544,N_9846);
xnor U10259 (N_10259,N_9769,N_9966);
nor U10260 (N_10260,N_9438,N_9289);
or U10261 (N_10261,N_9598,N_9293);
and U10262 (N_10262,N_9122,N_9235);
nand U10263 (N_10263,N_9709,N_9262);
xor U10264 (N_10264,N_9231,N_9333);
nand U10265 (N_10265,N_9463,N_9133);
nor U10266 (N_10266,N_9304,N_9152);
nor U10267 (N_10267,N_9026,N_9736);
and U10268 (N_10268,N_9574,N_9960);
xnor U10269 (N_10269,N_9760,N_9860);
nand U10270 (N_10270,N_9047,N_9712);
and U10271 (N_10271,N_9766,N_9816);
and U10272 (N_10272,N_9330,N_9311);
nor U10273 (N_10273,N_9472,N_9514);
nor U10274 (N_10274,N_9255,N_9425);
nand U10275 (N_10275,N_9485,N_9285);
or U10276 (N_10276,N_9242,N_9370);
nand U10277 (N_10277,N_9249,N_9049);
nor U10278 (N_10278,N_9334,N_9541);
nor U10279 (N_10279,N_9618,N_9479);
nand U10280 (N_10280,N_9500,N_9664);
and U10281 (N_10281,N_9164,N_9414);
and U10282 (N_10282,N_9678,N_9196);
xnor U10283 (N_10283,N_9830,N_9172);
xor U10284 (N_10284,N_9601,N_9391);
or U10285 (N_10285,N_9836,N_9935);
or U10286 (N_10286,N_9151,N_9264);
nor U10287 (N_10287,N_9348,N_9198);
nand U10288 (N_10288,N_9972,N_9958);
and U10289 (N_10289,N_9288,N_9418);
nand U10290 (N_10290,N_9147,N_9540);
nor U10291 (N_10291,N_9988,N_9496);
and U10292 (N_10292,N_9405,N_9432);
xnor U10293 (N_10293,N_9819,N_9523);
or U10294 (N_10294,N_9193,N_9563);
and U10295 (N_10295,N_9652,N_9085);
nor U10296 (N_10296,N_9318,N_9028);
or U10297 (N_10297,N_9458,N_9582);
or U10298 (N_10298,N_9627,N_9522);
or U10299 (N_10299,N_9554,N_9524);
nor U10300 (N_10300,N_9070,N_9872);
xor U10301 (N_10301,N_9052,N_9009);
and U10302 (N_10302,N_9043,N_9337);
nor U10303 (N_10303,N_9589,N_9804);
and U10304 (N_10304,N_9325,N_9388);
xor U10305 (N_10305,N_9208,N_9090);
and U10306 (N_10306,N_9735,N_9910);
xor U10307 (N_10307,N_9877,N_9850);
xnor U10308 (N_10308,N_9942,N_9922);
nand U10309 (N_10309,N_9898,N_9606);
nand U10310 (N_10310,N_9399,N_9701);
xor U10311 (N_10311,N_9714,N_9319);
xnor U10312 (N_10312,N_9844,N_9739);
nor U10313 (N_10313,N_9445,N_9653);
nand U10314 (N_10314,N_9272,N_9526);
or U10315 (N_10315,N_9247,N_9897);
or U10316 (N_10316,N_9489,N_9108);
or U10317 (N_10317,N_9979,N_9001);
and U10318 (N_10318,N_9980,N_9977);
xnor U10319 (N_10319,N_9890,N_9673);
nand U10320 (N_10320,N_9923,N_9371);
nor U10321 (N_10321,N_9224,N_9212);
nor U10322 (N_10322,N_9385,N_9875);
nor U10323 (N_10323,N_9703,N_9253);
nor U10324 (N_10324,N_9530,N_9570);
and U10325 (N_10325,N_9774,N_9436);
nand U10326 (N_10326,N_9135,N_9809);
and U10327 (N_10327,N_9132,N_9747);
and U10328 (N_10328,N_9847,N_9491);
and U10329 (N_10329,N_9244,N_9352);
nor U10330 (N_10330,N_9237,N_9710);
or U10331 (N_10331,N_9535,N_9912);
and U10332 (N_10332,N_9918,N_9753);
or U10333 (N_10333,N_9801,N_9274);
nand U10334 (N_10334,N_9126,N_9331);
and U10335 (N_10335,N_9612,N_9321);
and U10336 (N_10336,N_9171,N_9775);
or U10337 (N_10337,N_9216,N_9113);
nor U10338 (N_10338,N_9192,N_9338);
nand U10339 (N_10339,N_9950,N_9434);
nand U10340 (N_10340,N_9577,N_9648);
nor U10341 (N_10341,N_9071,N_9719);
nand U10342 (N_10342,N_9914,N_9351);
nand U10343 (N_10343,N_9503,N_9003);
nor U10344 (N_10344,N_9140,N_9868);
and U10345 (N_10345,N_9625,N_9962);
and U10346 (N_10346,N_9223,N_9593);
nand U10347 (N_10347,N_9746,N_9827);
or U10348 (N_10348,N_9672,N_9158);
nor U10349 (N_10349,N_9698,N_9075);
or U10350 (N_10350,N_9200,N_9984);
or U10351 (N_10351,N_9384,N_9502);
and U10352 (N_10352,N_9723,N_9139);
nor U10353 (N_10353,N_9952,N_9616);
nor U10354 (N_10354,N_9034,N_9737);
or U10355 (N_10355,N_9437,N_9038);
or U10356 (N_10356,N_9768,N_9064);
nor U10357 (N_10357,N_9484,N_9449);
or U10358 (N_10358,N_9246,N_9891);
nand U10359 (N_10359,N_9734,N_9114);
and U10360 (N_10360,N_9580,N_9771);
xnor U10361 (N_10361,N_9478,N_9119);
nand U10362 (N_10362,N_9690,N_9459);
and U10363 (N_10363,N_9548,N_9373);
xor U10364 (N_10364,N_9374,N_9245);
nor U10365 (N_10365,N_9206,N_9842);
and U10366 (N_10366,N_9378,N_9100);
or U10367 (N_10367,N_9039,N_9336);
xor U10368 (N_10368,N_9506,N_9969);
xor U10369 (N_10369,N_9416,N_9778);
nand U10370 (N_10370,N_9050,N_9074);
or U10371 (N_10371,N_9252,N_9674);
and U10372 (N_10372,N_9160,N_9916);
nand U10373 (N_10373,N_9933,N_9782);
or U10374 (N_10374,N_9640,N_9427);
nor U10375 (N_10375,N_9093,N_9947);
or U10376 (N_10376,N_9763,N_9443);
or U10377 (N_10377,N_9169,N_9603);
and U10378 (N_10378,N_9985,N_9248);
xnor U10379 (N_10379,N_9092,N_9881);
nor U10380 (N_10380,N_9110,N_9317);
nor U10381 (N_10381,N_9396,N_9675);
or U10382 (N_10382,N_9970,N_9584);
or U10383 (N_10383,N_9865,N_9295);
or U10384 (N_10384,N_9783,N_9101);
and U10385 (N_10385,N_9944,N_9826);
nand U10386 (N_10386,N_9785,N_9795);
xor U10387 (N_10387,N_9243,N_9112);
nand U10388 (N_10388,N_9515,N_9787);
and U10389 (N_10389,N_9755,N_9545);
nand U10390 (N_10390,N_9467,N_9023);
nand U10391 (N_10391,N_9066,N_9369);
xnor U10392 (N_10392,N_9525,N_9290);
nor U10393 (N_10393,N_9691,N_9780);
nand U10394 (N_10394,N_9791,N_9240);
nand U10395 (N_10395,N_9125,N_9511);
or U10396 (N_10396,N_9302,N_9499);
and U10397 (N_10397,N_9081,N_9596);
or U10398 (N_10398,N_9956,N_9773);
xnor U10399 (N_10399,N_9720,N_9163);
nor U10400 (N_10400,N_9642,N_9659);
xor U10401 (N_10401,N_9403,N_9798);
nor U10402 (N_10402,N_9907,N_9482);
nor U10403 (N_10403,N_9994,N_9409);
xor U10404 (N_10404,N_9829,N_9547);
nor U10405 (N_10405,N_9841,N_9611);
nand U10406 (N_10406,N_9764,N_9621);
and U10407 (N_10407,N_9579,N_9065);
nor U10408 (N_10408,N_9273,N_9624);
or U10409 (N_10409,N_9008,N_9848);
or U10410 (N_10410,N_9328,N_9076);
nand U10411 (N_10411,N_9936,N_9940);
and U10412 (N_10412,N_9035,N_9398);
nor U10413 (N_10413,N_9086,N_9037);
and U10414 (N_10414,N_9444,N_9267);
xor U10415 (N_10415,N_9590,N_9662);
and U10416 (N_10416,N_9493,N_9012);
xor U10417 (N_10417,N_9820,N_9792);
nor U10418 (N_10418,N_9754,N_9341);
or U10419 (N_10419,N_9156,N_9623);
and U10420 (N_10420,N_9679,N_9483);
nand U10421 (N_10421,N_9106,N_9433);
nor U10422 (N_10422,N_9280,N_9470);
xnor U10423 (N_10423,N_9518,N_9937);
nor U10424 (N_10424,N_9170,N_9959);
nor U10425 (N_10425,N_9646,N_9928);
nor U10426 (N_10426,N_9718,N_9487);
nand U10427 (N_10427,N_9594,N_9464);
nand U10428 (N_10428,N_9740,N_9759);
xor U10429 (N_10429,N_9905,N_9297);
xor U10430 (N_10430,N_9059,N_9567);
nor U10431 (N_10431,N_9241,N_9301);
xor U10432 (N_10432,N_9042,N_9180);
nor U10433 (N_10433,N_9788,N_9620);
nand U10434 (N_10434,N_9098,N_9630);
xnor U10435 (N_10435,N_9688,N_9201);
nand U10436 (N_10436,N_9796,N_9149);
or U10437 (N_10437,N_9953,N_9505);
nor U10438 (N_10438,N_9669,N_9468);
xnor U10439 (N_10439,N_9299,N_9124);
xor U10440 (N_10440,N_9162,N_9079);
nor U10441 (N_10441,N_9990,N_9453);
and U10442 (N_10442,N_9429,N_9666);
nand U10443 (N_10443,N_9024,N_9744);
and U10444 (N_10444,N_9282,N_9571);
or U10445 (N_10445,N_9475,N_9943);
xnor U10446 (N_10446,N_9814,N_9932);
or U10447 (N_10447,N_9802,N_9291);
xor U10448 (N_10448,N_9346,N_9036);
nor U10449 (N_10449,N_9683,N_9218);
nor U10450 (N_10450,N_9677,N_9699);
or U10451 (N_10451,N_9109,N_9356);
nor U10452 (N_10452,N_9477,N_9327);
nand U10453 (N_10453,N_9057,N_9326);
nand U10454 (N_10454,N_9220,N_9259);
nand U10455 (N_10455,N_9440,N_9144);
and U10456 (N_10456,N_9469,N_9879);
nand U10457 (N_10457,N_9292,N_9357);
and U10458 (N_10458,N_9609,N_9055);
or U10459 (N_10459,N_9393,N_9939);
or U10460 (N_10460,N_9903,N_9344);
or U10461 (N_10461,N_9533,N_9512);
nand U10462 (N_10462,N_9420,N_9402);
nor U10463 (N_10463,N_9899,N_9225);
xor U10464 (N_10464,N_9377,N_9166);
nand U10465 (N_10465,N_9353,N_9316);
xor U10466 (N_10466,N_9685,N_9713);
nand U10467 (N_10467,N_9728,N_9631);
and U10468 (N_10468,N_9083,N_9051);
nor U10469 (N_10469,N_9355,N_9447);
nor U10470 (N_10470,N_9824,N_9194);
nor U10471 (N_10471,N_9407,N_9019);
nand U10472 (N_10472,N_9294,N_9885);
nand U10473 (N_10473,N_9987,N_9048);
or U10474 (N_10474,N_9300,N_9202);
nand U10475 (N_10475,N_9501,N_9743);
nand U10476 (N_10476,N_9232,N_9982);
nand U10477 (N_10477,N_9536,N_9931);
xnor U10478 (N_10478,N_9861,N_9238);
nand U10479 (N_10479,N_9121,N_9663);
or U10480 (N_10480,N_9214,N_9637);
xor U10481 (N_10481,N_9866,N_9367);
and U10482 (N_10482,N_9883,N_9991);
nand U10483 (N_10483,N_9184,N_9777);
and U10484 (N_10484,N_9159,N_9597);
and U10485 (N_10485,N_9529,N_9395);
nand U10486 (N_10486,N_9585,N_9572);
nand U10487 (N_10487,N_9670,N_9315);
nand U10488 (N_10488,N_9359,N_9322);
xor U10489 (N_10489,N_9748,N_9421);
and U10490 (N_10490,N_9419,N_9793);
nor U10491 (N_10491,N_9886,N_9702);
xnor U10492 (N_10492,N_9852,N_9635);
xor U10493 (N_10493,N_9339,N_9354);
nor U10494 (N_10494,N_9129,N_9134);
xnor U10495 (N_10495,N_9256,N_9022);
xnor U10496 (N_10496,N_9465,N_9181);
and U10497 (N_10497,N_9439,N_9973);
or U10498 (N_10498,N_9832,N_9492);
or U10499 (N_10499,N_9298,N_9342);
nor U10500 (N_10500,N_9038,N_9410);
and U10501 (N_10501,N_9217,N_9448);
nor U10502 (N_10502,N_9654,N_9530);
xor U10503 (N_10503,N_9360,N_9610);
nand U10504 (N_10504,N_9731,N_9662);
xor U10505 (N_10505,N_9521,N_9092);
nor U10506 (N_10506,N_9321,N_9708);
nand U10507 (N_10507,N_9973,N_9721);
nand U10508 (N_10508,N_9921,N_9213);
nor U10509 (N_10509,N_9531,N_9683);
and U10510 (N_10510,N_9223,N_9016);
xnor U10511 (N_10511,N_9819,N_9233);
and U10512 (N_10512,N_9176,N_9985);
nand U10513 (N_10513,N_9597,N_9363);
xor U10514 (N_10514,N_9051,N_9082);
or U10515 (N_10515,N_9479,N_9351);
xnor U10516 (N_10516,N_9810,N_9660);
nand U10517 (N_10517,N_9918,N_9402);
xor U10518 (N_10518,N_9410,N_9402);
nor U10519 (N_10519,N_9695,N_9857);
or U10520 (N_10520,N_9782,N_9108);
xor U10521 (N_10521,N_9344,N_9747);
or U10522 (N_10522,N_9816,N_9417);
nor U10523 (N_10523,N_9627,N_9281);
xor U10524 (N_10524,N_9808,N_9619);
and U10525 (N_10525,N_9680,N_9352);
xor U10526 (N_10526,N_9873,N_9515);
or U10527 (N_10527,N_9266,N_9132);
and U10528 (N_10528,N_9766,N_9502);
or U10529 (N_10529,N_9754,N_9967);
and U10530 (N_10530,N_9737,N_9394);
and U10531 (N_10531,N_9402,N_9107);
nand U10532 (N_10532,N_9968,N_9636);
or U10533 (N_10533,N_9281,N_9900);
or U10534 (N_10534,N_9644,N_9738);
nor U10535 (N_10535,N_9500,N_9413);
nand U10536 (N_10536,N_9177,N_9446);
nor U10537 (N_10537,N_9471,N_9988);
nand U10538 (N_10538,N_9101,N_9800);
nand U10539 (N_10539,N_9068,N_9975);
nor U10540 (N_10540,N_9508,N_9393);
or U10541 (N_10541,N_9654,N_9413);
or U10542 (N_10542,N_9649,N_9942);
or U10543 (N_10543,N_9791,N_9645);
nor U10544 (N_10544,N_9773,N_9740);
nor U10545 (N_10545,N_9996,N_9546);
nand U10546 (N_10546,N_9400,N_9038);
and U10547 (N_10547,N_9716,N_9022);
nand U10548 (N_10548,N_9531,N_9848);
and U10549 (N_10549,N_9594,N_9162);
nor U10550 (N_10550,N_9964,N_9082);
nand U10551 (N_10551,N_9414,N_9511);
xnor U10552 (N_10552,N_9815,N_9062);
nor U10553 (N_10553,N_9363,N_9843);
nor U10554 (N_10554,N_9369,N_9497);
nor U10555 (N_10555,N_9740,N_9962);
or U10556 (N_10556,N_9089,N_9508);
or U10557 (N_10557,N_9612,N_9592);
nand U10558 (N_10558,N_9416,N_9022);
xor U10559 (N_10559,N_9128,N_9993);
nor U10560 (N_10560,N_9616,N_9314);
nor U10561 (N_10561,N_9019,N_9758);
or U10562 (N_10562,N_9636,N_9184);
nand U10563 (N_10563,N_9240,N_9008);
nor U10564 (N_10564,N_9047,N_9677);
nor U10565 (N_10565,N_9962,N_9426);
nand U10566 (N_10566,N_9560,N_9873);
xor U10567 (N_10567,N_9896,N_9413);
nor U10568 (N_10568,N_9005,N_9689);
xnor U10569 (N_10569,N_9047,N_9744);
nand U10570 (N_10570,N_9324,N_9234);
or U10571 (N_10571,N_9957,N_9840);
xnor U10572 (N_10572,N_9343,N_9817);
or U10573 (N_10573,N_9649,N_9037);
xor U10574 (N_10574,N_9335,N_9205);
or U10575 (N_10575,N_9335,N_9312);
xnor U10576 (N_10576,N_9131,N_9989);
and U10577 (N_10577,N_9588,N_9615);
or U10578 (N_10578,N_9322,N_9381);
xor U10579 (N_10579,N_9852,N_9050);
xor U10580 (N_10580,N_9784,N_9667);
nand U10581 (N_10581,N_9228,N_9620);
nor U10582 (N_10582,N_9442,N_9905);
nand U10583 (N_10583,N_9234,N_9655);
xor U10584 (N_10584,N_9248,N_9656);
or U10585 (N_10585,N_9388,N_9767);
nand U10586 (N_10586,N_9345,N_9238);
nor U10587 (N_10587,N_9331,N_9795);
xor U10588 (N_10588,N_9824,N_9727);
nand U10589 (N_10589,N_9508,N_9168);
xor U10590 (N_10590,N_9572,N_9846);
nor U10591 (N_10591,N_9939,N_9711);
and U10592 (N_10592,N_9933,N_9993);
and U10593 (N_10593,N_9996,N_9449);
and U10594 (N_10594,N_9893,N_9418);
xor U10595 (N_10595,N_9160,N_9217);
or U10596 (N_10596,N_9726,N_9052);
and U10597 (N_10597,N_9584,N_9088);
nor U10598 (N_10598,N_9207,N_9014);
nand U10599 (N_10599,N_9516,N_9202);
nor U10600 (N_10600,N_9434,N_9121);
and U10601 (N_10601,N_9827,N_9694);
nand U10602 (N_10602,N_9634,N_9073);
and U10603 (N_10603,N_9394,N_9976);
and U10604 (N_10604,N_9295,N_9477);
nand U10605 (N_10605,N_9143,N_9218);
nor U10606 (N_10606,N_9399,N_9629);
and U10607 (N_10607,N_9986,N_9055);
or U10608 (N_10608,N_9509,N_9789);
or U10609 (N_10609,N_9107,N_9201);
and U10610 (N_10610,N_9408,N_9206);
and U10611 (N_10611,N_9649,N_9744);
xor U10612 (N_10612,N_9365,N_9603);
nor U10613 (N_10613,N_9159,N_9844);
or U10614 (N_10614,N_9934,N_9830);
and U10615 (N_10615,N_9947,N_9832);
xor U10616 (N_10616,N_9248,N_9129);
nor U10617 (N_10617,N_9381,N_9566);
xnor U10618 (N_10618,N_9875,N_9263);
or U10619 (N_10619,N_9867,N_9080);
nor U10620 (N_10620,N_9222,N_9274);
and U10621 (N_10621,N_9831,N_9406);
or U10622 (N_10622,N_9776,N_9556);
nand U10623 (N_10623,N_9055,N_9021);
nand U10624 (N_10624,N_9177,N_9031);
nor U10625 (N_10625,N_9408,N_9884);
nor U10626 (N_10626,N_9897,N_9833);
nand U10627 (N_10627,N_9730,N_9375);
nand U10628 (N_10628,N_9432,N_9641);
and U10629 (N_10629,N_9064,N_9953);
or U10630 (N_10630,N_9559,N_9020);
nand U10631 (N_10631,N_9093,N_9767);
or U10632 (N_10632,N_9752,N_9167);
or U10633 (N_10633,N_9055,N_9735);
xor U10634 (N_10634,N_9558,N_9352);
nor U10635 (N_10635,N_9745,N_9423);
xnor U10636 (N_10636,N_9831,N_9547);
nor U10637 (N_10637,N_9517,N_9656);
nand U10638 (N_10638,N_9275,N_9283);
and U10639 (N_10639,N_9456,N_9181);
nand U10640 (N_10640,N_9811,N_9097);
nand U10641 (N_10641,N_9811,N_9957);
xnor U10642 (N_10642,N_9793,N_9393);
nand U10643 (N_10643,N_9189,N_9071);
and U10644 (N_10644,N_9865,N_9453);
xnor U10645 (N_10645,N_9041,N_9682);
and U10646 (N_10646,N_9544,N_9918);
nand U10647 (N_10647,N_9934,N_9590);
nor U10648 (N_10648,N_9539,N_9596);
and U10649 (N_10649,N_9357,N_9449);
xnor U10650 (N_10650,N_9566,N_9515);
or U10651 (N_10651,N_9116,N_9867);
nor U10652 (N_10652,N_9993,N_9832);
nor U10653 (N_10653,N_9898,N_9429);
nor U10654 (N_10654,N_9057,N_9831);
and U10655 (N_10655,N_9302,N_9043);
or U10656 (N_10656,N_9631,N_9778);
xor U10657 (N_10657,N_9024,N_9848);
xor U10658 (N_10658,N_9583,N_9702);
or U10659 (N_10659,N_9174,N_9804);
xor U10660 (N_10660,N_9847,N_9944);
nor U10661 (N_10661,N_9068,N_9516);
xor U10662 (N_10662,N_9599,N_9421);
or U10663 (N_10663,N_9288,N_9759);
and U10664 (N_10664,N_9414,N_9433);
and U10665 (N_10665,N_9888,N_9476);
or U10666 (N_10666,N_9938,N_9522);
and U10667 (N_10667,N_9033,N_9480);
xnor U10668 (N_10668,N_9667,N_9137);
and U10669 (N_10669,N_9668,N_9286);
nor U10670 (N_10670,N_9329,N_9079);
and U10671 (N_10671,N_9806,N_9084);
and U10672 (N_10672,N_9372,N_9339);
xor U10673 (N_10673,N_9251,N_9012);
or U10674 (N_10674,N_9256,N_9667);
or U10675 (N_10675,N_9970,N_9972);
or U10676 (N_10676,N_9073,N_9643);
xnor U10677 (N_10677,N_9798,N_9688);
nand U10678 (N_10678,N_9371,N_9377);
nor U10679 (N_10679,N_9825,N_9508);
nand U10680 (N_10680,N_9960,N_9969);
nand U10681 (N_10681,N_9854,N_9544);
nor U10682 (N_10682,N_9695,N_9917);
or U10683 (N_10683,N_9661,N_9698);
xor U10684 (N_10684,N_9760,N_9863);
nand U10685 (N_10685,N_9437,N_9101);
nand U10686 (N_10686,N_9274,N_9890);
and U10687 (N_10687,N_9404,N_9615);
or U10688 (N_10688,N_9965,N_9487);
or U10689 (N_10689,N_9746,N_9586);
xnor U10690 (N_10690,N_9556,N_9816);
or U10691 (N_10691,N_9104,N_9007);
and U10692 (N_10692,N_9496,N_9784);
nor U10693 (N_10693,N_9619,N_9119);
xnor U10694 (N_10694,N_9811,N_9214);
and U10695 (N_10695,N_9948,N_9835);
nand U10696 (N_10696,N_9667,N_9875);
nand U10697 (N_10697,N_9210,N_9590);
nand U10698 (N_10698,N_9220,N_9569);
nand U10699 (N_10699,N_9396,N_9827);
or U10700 (N_10700,N_9844,N_9983);
nand U10701 (N_10701,N_9564,N_9374);
xor U10702 (N_10702,N_9545,N_9692);
xor U10703 (N_10703,N_9120,N_9203);
nand U10704 (N_10704,N_9968,N_9897);
nor U10705 (N_10705,N_9154,N_9239);
nand U10706 (N_10706,N_9070,N_9913);
nand U10707 (N_10707,N_9542,N_9068);
xnor U10708 (N_10708,N_9761,N_9639);
nor U10709 (N_10709,N_9249,N_9891);
xnor U10710 (N_10710,N_9843,N_9813);
or U10711 (N_10711,N_9379,N_9911);
xor U10712 (N_10712,N_9244,N_9726);
xnor U10713 (N_10713,N_9994,N_9794);
xnor U10714 (N_10714,N_9936,N_9859);
nand U10715 (N_10715,N_9647,N_9560);
or U10716 (N_10716,N_9469,N_9096);
or U10717 (N_10717,N_9746,N_9418);
nor U10718 (N_10718,N_9384,N_9172);
nor U10719 (N_10719,N_9543,N_9335);
or U10720 (N_10720,N_9386,N_9793);
xor U10721 (N_10721,N_9537,N_9606);
nand U10722 (N_10722,N_9119,N_9191);
xor U10723 (N_10723,N_9809,N_9478);
or U10724 (N_10724,N_9757,N_9787);
or U10725 (N_10725,N_9943,N_9224);
and U10726 (N_10726,N_9870,N_9407);
or U10727 (N_10727,N_9733,N_9801);
nor U10728 (N_10728,N_9301,N_9260);
and U10729 (N_10729,N_9868,N_9257);
or U10730 (N_10730,N_9415,N_9483);
nor U10731 (N_10731,N_9146,N_9039);
and U10732 (N_10732,N_9489,N_9925);
xnor U10733 (N_10733,N_9543,N_9570);
or U10734 (N_10734,N_9897,N_9182);
nor U10735 (N_10735,N_9938,N_9411);
and U10736 (N_10736,N_9477,N_9795);
nor U10737 (N_10737,N_9307,N_9518);
or U10738 (N_10738,N_9895,N_9833);
nand U10739 (N_10739,N_9748,N_9192);
and U10740 (N_10740,N_9670,N_9693);
and U10741 (N_10741,N_9904,N_9024);
or U10742 (N_10742,N_9825,N_9496);
nand U10743 (N_10743,N_9943,N_9237);
or U10744 (N_10744,N_9198,N_9327);
or U10745 (N_10745,N_9717,N_9228);
nor U10746 (N_10746,N_9629,N_9049);
nor U10747 (N_10747,N_9375,N_9845);
xnor U10748 (N_10748,N_9665,N_9503);
or U10749 (N_10749,N_9184,N_9140);
nand U10750 (N_10750,N_9297,N_9038);
xor U10751 (N_10751,N_9600,N_9079);
or U10752 (N_10752,N_9630,N_9058);
xnor U10753 (N_10753,N_9942,N_9768);
xnor U10754 (N_10754,N_9099,N_9801);
xor U10755 (N_10755,N_9048,N_9999);
or U10756 (N_10756,N_9573,N_9840);
or U10757 (N_10757,N_9854,N_9721);
nand U10758 (N_10758,N_9732,N_9276);
or U10759 (N_10759,N_9843,N_9571);
nand U10760 (N_10760,N_9851,N_9047);
xor U10761 (N_10761,N_9892,N_9749);
nand U10762 (N_10762,N_9024,N_9605);
xor U10763 (N_10763,N_9263,N_9253);
nand U10764 (N_10764,N_9093,N_9192);
and U10765 (N_10765,N_9846,N_9543);
nor U10766 (N_10766,N_9293,N_9360);
and U10767 (N_10767,N_9066,N_9601);
and U10768 (N_10768,N_9088,N_9308);
nand U10769 (N_10769,N_9521,N_9267);
and U10770 (N_10770,N_9998,N_9570);
nor U10771 (N_10771,N_9062,N_9383);
nand U10772 (N_10772,N_9101,N_9290);
or U10773 (N_10773,N_9918,N_9777);
nand U10774 (N_10774,N_9999,N_9421);
nand U10775 (N_10775,N_9305,N_9911);
nor U10776 (N_10776,N_9640,N_9864);
xor U10777 (N_10777,N_9002,N_9140);
nand U10778 (N_10778,N_9152,N_9005);
nand U10779 (N_10779,N_9946,N_9650);
nor U10780 (N_10780,N_9016,N_9586);
nor U10781 (N_10781,N_9278,N_9019);
or U10782 (N_10782,N_9885,N_9298);
or U10783 (N_10783,N_9202,N_9648);
nor U10784 (N_10784,N_9873,N_9666);
nor U10785 (N_10785,N_9112,N_9208);
xor U10786 (N_10786,N_9220,N_9780);
and U10787 (N_10787,N_9014,N_9639);
xnor U10788 (N_10788,N_9553,N_9029);
nand U10789 (N_10789,N_9755,N_9479);
or U10790 (N_10790,N_9515,N_9343);
nor U10791 (N_10791,N_9770,N_9225);
or U10792 (N_10792,N_9986,N_9339);
xor U10793 (N_10793,N_9978,N_9641);
nand U10794 (N_10794,N_9421,N_9857);
and U10795 (N_10795,N_9914,N_9218);
nor U10796 (N_10796,N_9957,N_9323);
or U10797 (N_10797,N_9881,N_9784);
nand U10798 (N_10798,N_9826,N_9260);
or U10799 (N_10799,N_9430,N_9612);
and U10800 (N_10800,N_9547,N_9426);
and U10801 (N_10801,N_9163,N_9436);
nor U10802 (N_10802,N_9137,N_9538);
nand U10803 (N_10803,N_9335,N_9375);
nor U10804 (N_10804,N_9150,N_9612);
nor U10805 (N_10805,N_9101,N_9451);
xnor U10806 (N_10806,N_9520,N_9903);
or U10807 (N_10807,N_9921,N_9002);
and U10808 (N_10808,N_9433,N_9812);
nand U10809 (N_10809,N_9750,N_9175);
nor U10810 (N_10810,N_9163,N_9203);
xnor U10811 (N_10811,N_9274,N_9778);
nor U10812 (N_10812,N_9078,N_9233);
or U10813 (N_10813,N_9184,N_9992);
xnor U10814 (N_10814,N_9226,N_9243);
or U10815 (N_10815,N_9160,N_9853);
or U10816 (N_10816,N_9574,N_9524);
nor U10817 (N_10817,N_9809,N_9374);
nand U10818 (N_10818,N_9818,N_9378);
nor U10819 (N_10819,N_9411,N_9962);
or U10820 (N_10820,N_9148,N_9583);
nand U10821 (N_10821,N_9546,N_9076);
xor U10822 (N_10822,N_9668,N_9908);
xor U10823 (N_10823,N_9765,N_9581);
xor U10824 (N_10824,N_9864,N_9970);
xor U10825 (N_10825,N_9099,N_9569);
or U10826 (N_10826,N_9593,N_9060);
or U10827 (N_10827,N_9169,N_9577);
xnor U10828 (N_10828,N_9453,N_9451);
and U10829 (N_10829,N_9335,N_9988);
xor U10830 (N_10830,N_9255,N_9373);
or U10831 (N_10831,N_9385,N_9275);
nand U10832 (N_10832,N_9128,N_9514);
nand U10833 (N_10833,N_9889,N_9414);
nor U10834 (N_10834,N_9730,N_9086);
and U10835 (N_10835,N_9734,N_9066);
xnor U10836 (N_10836,N_9324,N_9908);
xnor U10837 (N_10837,N_9950,N_9432);
or U10838 (N_10838,N_9946,N_9547);
and U10839 (N_10839,N_9688,N_9253);
and U10840 (N_10840,N_9512,N_9303);
nand U10841 (N_10841,N_9463,N_9720);
nor U10842 (N_10842,N_9570,N_9586);
nand U10843 (N_10843,N_9880,N_9745);
nor U10844 (N_10844,N_9994,N_9540);
nand U10845 (N_10845,N_9487,N_9217);
or U10846 (N_10846,N_9292,N_9829);
nor U10847 (N_10847,N_9379,N_9014);
nor U10848 (N_10848,N_9206,N_9349);
nor U10849 (N_10849,N_9425,N_9723);
nor U10850 (N_10850,N_9135,N_9072);
xnor U10851 (N_10851,N_9920,N_9454);
and U10852 (N_10852,N_9382,N_9363);
xor U10853 (N_10853,N_9439,N_9825);
xnor U10854 (N_10854,N_9765,N_9545);
nand U10855 (N_10855,N_9211,N_9969);
or U10856 (N_10856,N_9512,N_9445);
and U10857 (N_10857,N_9796,N_9637);
xnor U10858 (N_10858,N_9922,N_9066);
nand U10859 (N_10859,N_9566,N_9706);
nor U10860 (N_10860,N_9840,N_9749);
nor U10861 (N_10861,N_9237,N_9647);
nand U10862 (N_10862,N_9315,N_9932);
nor U10863 (N_10863,N_9314,N_9587);
nor U10864 (N_10864,N_9054,N_9808);
or U10865 (N_10865,N_9888,N_9725);
nor U10866 (N_10866,N_9427,N_9436);
nor U10867 (N_10867,N_9350,N_9214);
or U10868 (N_10868,N_9071,N_9563);
nor U10869 (N_10869,N_9584,N_9284);
nand U10870 (N_10870,N_9149,N_9272);
or U10871 (N_10871,N_9247,N_9463);
nand U10872 (N_10872,N_9614,N_9773);
or U10873 (N_10873,N_9899,N_9520);
nor U10874 (N_10874,N_9141,N_9357);
or U10875 (N_10875,N_9328,N_9215);
nor U10876 (N_10876,N_9459,N_9559);
nand U10877 (N_10877,N_9422,N_9660);
nor U10878 (N_10878,N_9112,N_9605);
or U10879 (N_10879,N_9054,N_9638);
nand U10880 (N_10880,N_9383,N_9200);
nand U10881 (N_10881,N_9472,N_9304);
xnor U10882 (N_10882,N_9666,N_9931);
nand U10883 (N_10883,N_9641,N_9676);
xor U10884 (N_10884,N_9333,N_9297);
xnor U10885 (N_10885,N_9606,N_9849);
and U10886 (N_10886,N_9532,N_9685);
xor U10887 (N_10887,N_9166,N_9057);
xor U10888 (N_10888,N_9008,N_9249);
nand U10889 (N_10889,N_9261,N_9937);
xor U10890 (N_10890,N_9596,N_9181);
nor U10891 (N_10891,N_9936,N_9630);
xor U10892 (N_10892,N_9734,N_9976);
nand U10893 (N_10893,N_9744,N_9369);
and U10894 (N_10894,N_9799,N_9912);
nor U10895 (N_10895,N_9472,N_9908);
and U10896 (N_10896,N_9200,N_9749);
nand U10897 (N_10897,N_9081,N_9461);
nor U10898 (N_10898,N_9796,N_9132);
nor U10899 (N_10899,N_9876,N_9144);
xnor U10900 (N_10900,N_9805,N_9344);
and U10901 (N_10901,N_9725,N_9554);
or U10902 (N_10902,N_9378,N_9050);
or U10903 (N_10903,N_9474,N_9889);
xor U10904 (N_10904,N_9663,N_9142);
xnor U10905 (N_10905,N_9611,N_9745);
xor U10906 (N_10906,N_9581,N_9505);
and U10907 (N_10907,N_9015,N_9563);
nor U10908 (N_10908,N_9297,N_9925);
and U10909 (N_10909,N_9613,N_9757);
nor U10910 (N_10910,N_9580,N_9195);
or U10911 (N_10911,N_9157,N_9094);
nand U10912 (N_10912,N_9230,N_9316);
nor U10913 (N_10913,N_9513,N_9240);
nor U10914 (N_10914,N_9045,N_9488);
or U10915 (N_10915,N_9174,N_9925);
nand U10916 (N_10916,N_9392,N_9329);
nand U10917 (N_10917,N_9854,N_9694);
xor U10918 (N_10918,N_9020,N_9081);
xor U10919 (N_10919,N_9953,N_9774);
nand U10920 (N_10920,N_9752,N_9222);
and U10921 (N_10921,N_9339,N_9277);
nand U10922 (N_10922,N_9034,N_9863);
nor U10923 (N_10923,N_9288,N_9499);
nand U10924 (N_10924,N_9004,N_9716);
nand U10925 (N_10925,N_9897,N_9620);
xnor U10926 (N_10926,N_9302,N_9421);
or U10927 (N_10927,N_9355,N_9930);
nor U10928 (N_10928,N_9357,N_9530);
and U10929 (N_10929,N_9660,N_9675);
nand U10930 (N_10930,N_9258,N_9976);
xnor U10931 (N_10931,N_9216,N_9176);
nand U10932 (N_10932,N_9631,N_9383);
xor U10933 (N_10933,N_9386,N_9915);
and U10934 (N_10934,N_9569,N_9841);
xnor U10935 (N_10935,N_9736,N_9132);
xnor U10936 (N_10936,N_9044,N_9989);
nand U10937 (N_10937,N_9725,N_9651);
nand U10938 (N_10938,N_9656,N_9366);
or U10939 (N_10939,N_9202,N_9559);
nand U10940 (N_10940,N_9340,N_9701);
xor U10941 (N_10941,N_9193,N_9993);
or U10942 (N_10942,N_9967,N_9712);
or U10943 (N_10943,N_9477,N_9572);
nand U10944 (N_10944,N_9135,N_9623);
xnor U10945 (N_10945,N_9107,N_9856);
xnor U10946 (N_10946,N_9147,N_9098);
and U10947 (N_10947,N_9914,N_9226);
or U10948 (N_10948,N_9007,N_9592);
and U10949 (N_10949,N_9984,N_9024);
and U10950 (N_10950,N_9410,N_9065);
xor U10951 (N_10951,N_9753,N_9589);
nand U10952 (N_10952,N_9258,N_9586);
or U10953 (N_10953,N_9026,N_9698);
nand U10954 (N_10954,N_9850,N_9822);
nor U10955 (N_10955,N_9593,N_9027);
nor U10956 (N_10956,N_9290,N_9462);
nand U10957 (N_10957,N_9302,N_9163);
nand U10958 (N_10958,N_9914,N_9924);
or U10959 (N_10959,N_9839,N_9747);
nand U10960 (N_10960,N_9294,N_9980);
and U10961 (N_10961,N_9288,N_9474);
nand U10962 (N_10962,N_9970,N_9672);
and U10963 (N_10963,N_9728,N_9666);
or U10964 (N_10964,N_9052,N_9802);
xnor U10965 (N_10965,N_9374,N_9872);
nor U10966 (N_10966,N_9077,N_9978);
and U10967 (N_10967,N_9842,N_9532);
nand U10968 (N_10968,N_9964,N_9408);
or U10969 (N_10969,N_9958,N_9285);
nand U10970 (N_10970,N_9570,N_9758);
nand U10971 (N_10971,N_9546,N_9388);
or U10972 (N_10972,N_9059,N_9545);
or U10973 (N_10973,N_9561,N_9711);
or U10974 (N_10974,N_9094,N_9664);
and U10975 (N_10975,N_9389,N_9149);
nor U10976 (N_10976,N_9051,N_9975);
or U10977 (N_10977,N_9253,N_9319);
xnor U10978 (N_10978,N_9447,N_9339);
and U10979 (N_10979,N_9056,N_9151);
and U10980 (N_10980,N_9091,N_9202);
xnor U10981 (N_10981,N_9668,N_9088);
nand U10982 (N_10982,N_9691,N_9462);
or U10983 (N_10983,N_9316,N_9686);
xnor U10984 (N_10984,N_9983,N_9681);
nand U10985 (N_10985,N_9916,N_9512);
and U10986 (N_10986,N_9890,N_9568);
xor U10987 (N_10987,N_9835,N_9366);
xor U10988 (N_10988,N_9088,N_9922);
or U10989 (N_10989,N_9949,N_9127);
xor U10990 (N_10990,N_9740,N_9295);
nor U10991 (N_10991,N_9103,N_9162);
nor U10992 (N_10992,N_9605,N_9552);
nor U10993 (N_10993,N_9878,N_9057);
xnor U10994 (N_10994,N_9117,N_9664);
xor U10995 (N_10995,N_9029,N_9490);
and U10996 (N_10996,N_9769,N_9246);
xnor U10997 (N_10997,N_9765,N_9424);
nor U10998 (N_10998,N_9052,N_9431);
or U10999 (N_10999,N_9911,N_9024);
and U11000 (N_11000,N_10736,N_10685);
and U11001 (N_11001,N_10236,N_10772);
or U11002 (N_11002,N_10264,N_10589);
nor U11003 (N_11003,N_10858,N_10691);
and U11004 (N_11004,N_10355,N_10136);
and U11005 (N_11005,N_10290,N_10612);
and U11006 (N_11006,N_10856,N_10559);
nand U11007 (N_11007,N_10238,N_10217);
xor U11008 (N_11008,N_10921,N_10545);
or U11009 (N_11009,N_10558,N_10582);
xnor U11010 (N_11010,N_10020,N_10498);
and U11011 (N_11011,N_10576,N_10251);
nand U11012 (N_11012,N_10587,N_10477);
or U11013 (N_11013,N_10322,N_10708);
and U11014 (N_11014,N_10200,N_10280);
or U11015 (N_11015,N_10653,N_10434);
xor U11016 (N_11016,N_10261,N_10276);
nand U11017 (N_11017,N_10321,N_10373);
nor U11018 (N_11018,N_10121,N_10744);
xor U11019 (N_11019,N_10777,N_10099);
or U11020 (N_11020,N_10516,N_10330);
or U11021 (N_11021,N_10523,N_10671);
xnor U11022 (N_11022,N_10996,N_10940);
or U11023 (N_11023,N_10230,N_10279);
nand U11024 (N_11024,N_10104,N_10959);
xnor U11025 (N_11025,N_10145,N_10155);
xor U11026 (N_11026,N_10323,N_10361);
nor U11027 (N_11027,N_10304,N_10511);
and U11028 (N_11028,N_10480,N_10388);
nand U11029 (N_11029,N_10985,N_10951);
nand U11030 (N_11030,N_10339,N_10014);
or U11031 (N_11031,N_10939,N_10897);
and U11032 (N_11032,N_10364,N_10920);
nand U11033 (N_11033,N_10118,N_10004);
xnor U11034 (N_11034,N_10332,N_10656);
and U11035 (N_11035,N_10954,N_10175);
nand U11036 (N_11036,N_10504,N_10342);
and U11037 (N_11037,N_10187,N_10196);
nor U11038 (N_11038,N_10611,N_10098);
or U11039 (N_11039,N_10271,N_10305);
and U11040 (N_11040,N_10444,N_10378);
xor U11041 (N_11041,N_10413,N_10181);
or U11042 (N_11042,N_10423,N_10336);
or U11043 (N_11043,N_10866,N_10536);
nand U11044 (N_11044,N_10282,N_10199);
xnor U11045 (N_11045,N_10811,N_10462);
xnor U11046 (N_11046,N_10335,N_10624);
or U11047 (N_11047,N_10619,N_10551);
xor U11048 (N_11048,N_10844,N_10605);
nand U11049 (N_11049,N_10763,N_10267);
or U11050 (N_11050,N_10519,N_10234);
and U11051 (N_11051,N_10334,N_10829);
or U11052 (N_11052,N_10971,N_10878);
nand U11053 (N_11053,N_10639,N_10302);
xor U11054 (N_11054,N_10179,N_10190);
nand U11055 (N_11055,N_10815,N_10184);
nor U11056 (N_11056,N_10781,N_10407);
or U11057 (N_11057,N_10202,N_10817);
and U11058 (N_11058,N_10703,N_10124);
and U11059 (N_11059,N_10440,N_10592);
nor U11060 (N_11060,N_10274,N_10901);
or U11061 (N_11061,N_10561,N_10354);
nand U11062 (N_11062,N_10823,N_10659);
nand U11063 (N_11063,N_10239,N_10418);
and U11064 (N_11064,N_10734,N_10151);
nand U11065 (N_11065,N_10879,N_10982);
nand U11066 (N_11066,N_10645,N_10320);
and U11067 (N_11067,N_10412,N_10924);
nand U11068 (N_11068,N_10648,N_10788);
or U11069 (N_11069,N_10032,N_10510);
nor U11070 (N_11070,N_10075,N_10748);
nand U11071 (N_11071,N_10052,N_10137);
and U11072 (N_11072,N_10689,N_10860);
xor U11073 (N_11073,N_10345,N_10735);
xnor U11074 (N_11074,N_10352,N_10380);
or U11075 (N_11075,N_10517,N_10713);
nand U11076 (N_11076,N_10430,N_10543);
nor U11077 (N_11077,N_10360,N_10168);
nor U11078 (N_11078,N_10021,N_10278);
or U11079 (N_11079,N_10984,N_10919);
or U11080 (N_11080,N_10556,N_10186);
xnor U11081 (N_11081,N_10188,N_10270);
and U11082 (N_11082,N_10716,N_10937);
and U11083 (N_11083,N_10141,N_10712);
nand U11084 (N_11084,N_10415,N_10376);
nor U11085 (N_11085,N_10068,N_10389);
nor U11086 (N_11086,N_10191,N_10180);
nor U11087 (N_11087,N_10701,N_10630);
xor U11088 (N_11088,N_10599,N_10318);
xor U11089 (N_11089,N_10262,N_10909);
or U11090 (N_11090,N_10309,N_10082);
or U11091 (N_11091,N_10833,N_10719);
or U11092 (N_11092,N_10529,N_10260);
nand U11093 (N_11093,N_10385,N_10852);
xnor U11094 (N_11094,N_10614,N_10315);
xnor U11095 (N_11095,N_10802,N_10353);
nor U11096 (N_11096,N_10953,N_10973);
xor U11097 (N_11097,N_10835,N_10720);
and U11098 (N_11098,N_10649,N_10492);
xor U11099 (N_11099,N_10818,N_10874);
xnor U11100 (N_11100,N_10692,N_10441);
or U11101 (N_11101,N_10314,N_10421);
nor U11102 (N_11102,N_10842,N_10864);
nor U11103 (N_11103,N_10483,N_10031);
nor U11104 (N_11104,N_10149,N_10058);
nand U11105 (N_11105,N_10227,N_10515);
and U11106 (N_11106,N_10346,N_10045);
or U11107 (N_11107,N_10896,N_10437);
and U11108 (N_11108,N_10950,N_10451);
nor U11109 (N_11109,N_10481,N_10681);
nor U11110 (N_11110,N_10790,N_10872);
nor U11111 (N_11111,N_10573,N_10550);
xor U11112 (N_11112,N_10016,N_10591);
and U11113 (N_11113,N_10223,N_10257);
xnor U11114 (N_11114,N_10123,N_10208);
and U11115 (N_11115,N_10733,N_10494);
xor U11116 (N_11116,N_10759,N_10524);
or U11117 (N_11117,N_10158,N_10508);
nand U11118 (N_11118,N_10647,N_10764);
and U11119 (N_11119,N_10646,N_10225);
nor U11120 (N_11120,N_10436,N_10221);
nor U11121 (N_11121,N_10269,N_10888);
or U11122 (N_11122,N_10870,N_10411);
xor U11123 (N_11123,N_10534,N_10918);
xor U11124 (N_11124,N_10846,N_10590);
nand U11125 (N_11125,N_10538,N_10869);
or U11126 (N_11126,N_10706,N_10432);
or U11127 (N_11127,N_10102,N_10549);
and U11128 (N_11128,N_10542,N_10891);
or U11129 (N_11129,N_10533,N_10029);
or U11130 (N_11130,N_10563,N_10015);
and U11131 (N_11131,N_10779,N_10938);
or U11132 (N_11132,N_10072,N_10443);
and U11133 (N_11133,N_10933,N_10327);
and U11134 (N_11134,N_10328,N_10969);
or U11135 (N_11135,N_10310,N_10008);
xor U11136 (N_11136,N_10452,N_10762);
nor U11137 (N_11137,N_10885,N_10643);
or U11138 (N_11138,N_10770,N_10402);
and U11139 (N_11139,N_10688,N_10193);
xor U11140 (N_11140,N_10146,N_10473);
nor U11141 (N_11141,N_10560,N_10999);
nor U11142 (N_11142,N_10140,N_10286);
and U11143 (N_11143,N_10166,N_10172);
or U11144 (N_11144,N_10489,N_10721);
nor U11145 (N_11145,N_10908,N_10571);
xnor U11146 (N_11146,N_10340,N_10800);
xnor U11147 (N_11147,N_10981,N_10666);
or U11148 (N_11148,N_10059,N_10727);
nand U11149 (N_11149,N_10034,N_10663);
and U11150 (N_11150,N_10917,N_10813);
nand U11151 (N_11151,N_10192,N_10085);
or U11152 (N_11152,N_10636,N_10952);
and U11153 (N_11153,N_10774,N_10690);
or U11154 (N_11154,N_10446,N_10326);
nor U11155 (N_11155,N_10694,N_10163);
nand U11156 (N_11156,N_10922,N_10367);
or U11157 (N_11157,N_10568,N_10297);
or U11158 (N_11158,N_10362,N_10396);
nor U11159 (N_11159,N_10975,N_10512);
nor U11160 (N_11160,N_10488,N_10993);
or U11161 (N_11161,N_10469,N_10760);
and U11162 (N_11162,N_10174,N_10111);
nand U11163 (N_11163,N_10555,N_10859);
and U11164 (N_11164,N_10294,N_10577);
nand U11165 (N_11165,N_10672,N_10078);
or U11166 (N_11166,N_10055,N_10638);
nand U11167 (N_11167,N_10868,N_10358);
and U11168 (N_11168,N_10097,N_10000);
nor U11169 (N_11169,N_10381,N_10509);
or U11170 (N_11170,N_10363,N_10377);
nor U11171 (N_11171,N_10350,N_10356);
nand U11172 (N_11172,N_10926,N_10383);
nor U11173 (N_11173,N_10417,N_10037);
and U11174 (N_11174,N_10070,N_10784);
and U11175 (N_11175,N_10329,N_10007);
or U11176 (N_11176,N_10718,N_10005);
or U11177 (N_11177,N_10684,N_10991);
nor U11178 (N_11178,N_10821,N_10203);
and U11179 (N_11179,N_10880,N_10847);
xnor U11180 (N_11180,N_10929,N_10107);
nor U11181 (N_11181,N_10226,N_10403);
nand U11182 (N_11182,N_10125,N_10303);
nand U11183 (N_11183,N_10678,N_10069);
nor U11184 (N_11184,N_10899,N_10414);
and U11185 (N_11185,N_10958,N_10903);
nand U11186 (N_11186,N_10080,N_10916);
or U11187 (N_11187,N_10170,N_10898);
or U11188 (N_11188,N_10925,N_10812);
and U11189 (N_11189,N_10114,N_10507);
nand U11190 (N_11190,N_10066,N_10033);
and U11191 (N_11191,N_10474,N_10240);
or U11192 (N_11192,N_10062,N_10743);
and U11193 (N_11193,N_10526,N_10017);
nor U11194 (N_11194,N_10698,N_10875);
or U11195 (N_11195,N_10990,N_10127);
nand U11196 (N_11196,N_10810,N_10795);
xnor U11197 (N_11197,N_10265,N_10243);
nand U11198 (N_11198,N_10466,N_10479);
nor U11199 (N_11199,N_10911,N_10369);
nand U11200 (N_11200,N_10861,N_10902);
and U11201 (N_11201,N_10038,N_10700);
nand U11202 (N_11202,N_10704,N_10094);
nand U11203 (N_11203,N_10333,N_10120);
xnor U11204 (N_11204,N_10801,N_10207);
xnor U11205 (N_11205,N_10397,N_10632);
or U11206 (N_11206,N_10325,N_10729);
and U11207 (N_11207,N_10886,N_10967);
or U11208 (N_11208,N_10955,N_10129);
nor U11209 (N_11209,N_10475,N_10600);
nor U11210 (N_11210,N_10862,N_10301);
and U11211 (N_11211,N_10883,N_10987);
nor U11212 (N_11212,N_10505,N_10461);
nor U11213 (N_11213,N_10637,N_10252);
or U11214 (N_11214,N_10424,N_10518);
nor U11215 (N_11215,N_10197,N_10608);
or U11216 (N_11216,N_10826,N_10827);
or U11217 (N_11217,N_10154,N_10410);
or U11218 (N_11218,N_10357,N_10831);
and U11219 (N_11219,N_10962,N_10845);
nor U11220 (N_11220,N_10914,N_10022);
nor U11221 (N_11221,N_10669,N_10843);
nor U11222 (N_11222,N_10983,N_10283);
nand U11223 (N_11223,N_10088,N_10351);
nor U11224 (N_11224,N_10131,N_10242);
nand U11225 (N_11225,N_10285,N_10687);
xor U11226 (N_11226,N_10408,N_10799);
xor U11227 (N_11227,N_10173,N_10287);
nor U11228 (N_11228,N_10693,N_10667);
nand U11229 (N_11229,N_10820,N_10347);
nand U11230 (N_11230,N_10616,N_10247);
nand U11231 (N_11231,N_10579,N_10384);
nand U11232 (N_11232,N_10416,N_10541);
or U11233 (N_11233,N_10433,N_10295);
xnor U11234 (N_11234,N_10528,N_10372);
nor U11235 (N_11235,N_10644,N_10994);
or U11236 (N_11236,N_10628,N_10949);
nand U11237 (N_11237,N_10502,N_10025);
nand U11238 (N_11238,N_10064,N_10460);
xor U11239 (N_11239,N_10039,N_10881);
or U11240 (N_11240,N_10676,N_10796);
or U11241 (N_11241,N_10439,N_10081);
and U11242 (N_11242,N_10482,N_10359);
nand U11243 (N_11243,N_10048,N_10521);
nor U11244 (N_11244,N_10893,N_10049);
xnor U11245 (N_11245,N_10171,N_10404);
nand U11246 (N_11246,N_10185,N_10050);
xnor U11247 (N_11247,N_10244,N_10613);
nor U11248 (N_11248,N_10241,N_10936);
nor U11249 (N_11249,N_10857,N_10450);
nand U11250 (N_11250,N_10544,N_10824);
nor U11251 (N_11251,N_10840,N_10670);
and U11252 (N_11252,N_10231,N_10379);
nor U11253 (N_11253,N_10819,N_10679);
or U11254 (N_11254,N_10915,N_10836);
and U11255 (N_11255,N_10183,N_10786);
xnor U11256 (N_11256,N_10699,N_10079);
xnor U11257 (N_11257,N_10177,N_10745);
nor U11258 (N_11258,N_10368,N_10514);
xnor U11259 (N_11259,N_10932,N_10957);
or U11260 (N_11260,N_10018,N_10793);
xor U11261 (N_11261,N_10012,N_10974);
and U11262 (N_11262,N_10998,N_10750);
nand U11263 (N_11263,N_10675,N_10426);
nor U11264 (N_11264,N_10814,N_10245);
and U11265 (N_11265,N_10453,N_10442);
or U11266 (N_11266,N_10429,N_10569);
nor U11267 (N_11267,N_10765,N_10660);
or U11268 (N_11268,N_10960,N_10895);
nor U11269 (N_11269,N_10393,N_10715);
nand U11270 (N_11270,N_10625,N_10749);
and U11271 (N_11271,N_10532,N_10520);
nor U11272 (N_11272,N_10597,N_10742);
xnor U11273 (N_11273,N_10618,N_10865);
xnor U11274 (N_11274,N_10476,N_10606);
nand U11275 (N_11275,N_10548,N_10463);
nand U11276 (N_11276,N_10074,N_10776);
and U11277 (N_11277,N_10740,N_10941);
or U11278 (N_11278,N_10527,N_10970);
nand U11279 (N_11279,N_10109,N_10317);
nor U11280 (N_11280,N_10757,N_10633);
nor U11281 (N_11281,N_10272,N_10602);
or U11282 (N_11282,N_10822,N_10714);
nor U11283 (N_11283,N_10841,N_10194);
nor U11284 (N_11284,N_10409,N_10258);
or U11285 (N_11285,N_10702,N_10060);
xor U11286 (N_11286,N_10850,N_10964);
xnor U11287 (N_11287,N_10448,N_10807);
nand U11288 (N_11288,N_10428,N_10495);
nand U11289 (N_11289,N_10567,N_10565);
xor U11290 (N_11290,N_10054,N_10112);
or U11291 (N_11291,N_10574,N_10837);
xor U11292 (N_11292,N_10655,N_10894);
and U11293 (N_11293,N_10246,N_10210);
xor U11294 (N_11294,N_10797,N_10047);
nor U11295 (N_11295,N_10108,N_10289);
xor U11296 (N_11296,N_10201,N_10890);
or U11297 (N_11297,N_10553,N_10027);
and U11298 (N_11298,N_10132,N_10405);
xor U11299 (N_11299,N_10316,N_10406);
and U11300 (N_11300,N_10882,N_10254);
nor U11301 (N_11301,N_10106,N_10293);
or U11302 (N_11302,N_10013,N_10988);
xor U11303 (N_11303,N_10500,N_10906);
nand U11304 (N_11304,N_10755,N_10089);
and U11305 (N_11305,N_10023,N_10552);
nand U11306 (N_11306,N_10931,N_10043);
nor U11307 (N_11307,N_10945,N_10601);
nor U11308 (N_11308,N_10782,N_10387);
xnor U11309 (N_11309,N_10913,N_10213);
and U11310 (N_11310,N_10621,N_10665);
or U11311 (N_11311,N_10593,N_10087);
xnor U11312 (N_11312,N_10848,N_10046);
nand U11313 (N_11313,N_10319,N_10311);
nand U11314 (N_11314,N_10067,N_10641);
and U11315 (N_11315,N_10738,N_10216);
nand U11316 (N_11316,N_10259,N_10133);
nand U11317 (N_11317,N_10499,N_10176);
nand U11318 (N_11318,N_10465,N_10178);
nor U11319 (N_11319,N_10609,N_10233);
and U11320 (N_11320,N_10491,N_10584);
xnor U11321 (N_11321,N_10224,N_10851);
xor U11322 (N_11322,N_10904,N_10161);
nor U11323 (N_11323,N_10229,N_10547);
nor U11324 (N_11324,N_10654,N_10657);
nand U11325 (N_11325,N_10871,N_10503);
and U11326 (N_11326,N_10331,N_10739);
and U11327 (N_11327,N_10530,N_10662);
nand U11328 (N_11328,N_10711,N_10255);
nor U11329 (N_11329,N_10496,N_10767);
xor U11330 (N_11330,N_10493,N_10091);
and U11331 (N_11331,N_10586,N_10296);
xnor U11332 (N_11332,N_10126,N_10658);
or U11333 (N_11333,N_10997,N_10972);
nor U11334 (N_11334,N_10741,N_10620);
xnor U11335 (N_11335,N_10263,N_10009);
nand U11336 (N_11336,N_10071,N_10930);
nor U11337 (N_11337,N_10884,N_10564);
nor U11338 (N_11338,N_10169,N_10751);
or U11339 (N_11339,N_10392,N_10768);
nand U11340 (N_11340,N_10731,N_10370);
and U11341 (N_11341,N_10337,N_10642);
xor U11342 (N_11342,N_10732,N_10531);
nand U11343 (N_11343,N_10454,N_10787);
nor U11344 (N_11344,N_10134,N_10113);
and U11345 (N_11345,N_10422,N_10809);
xnor U11346 (N_11346,N_10853,N_10273);
and U11347 (N_11347,N_10401,N_10617);
xnor U11348 (N_11348,N_10570,N_10391);
or U11349 (N_11349,N_10947,N_10250);
nand U11350 (N_11350,N_10956,N_10976);
or U11351 (N_11351,N_10035,N_10832);
nand U11352 (N_11352,N_10724,N_10537);
or U11353 (N_11353,N_10139,N_10209);
nand U11354 (N_11354,N_10595,N_10157);
nand U11355 (N_11355,N_10220,N_10980);
nand U11356 (N_11356,N_10603,N_10828);
xor U11357 (N_11357,N_10501,N_10943);
or U11358 (N_11358,N_10771,N_10298);
nand U11359 (N_11359,N_10472,N_10961);
or U11360 (N_11360,N_10816,N_10338);
or U11361 (N_11361,N_10773,N_10281);
xor U11362 (N_11362,N_10044,N_10578);
or U11363 (N_11363,N_10855,N_10839);
or U11364 (N_11364,N_10195,N_10420);
nor U11365 (N_11365,N_10651,N_10775);
xor U11366 (N_11366,N_10594,N_10825);
and U11367 (N_11367,N_10854,N_10892);
nor U11368 (N_11368,N_10723,N_10053);
xor U11369 (N_11369,N_10096,N_10977);
or U11370 (N_11370,N_10083,N_10717);
nor U11371 (N_11371,N_10623,N_10769);
and U11372 (N_11372,N_10927,N_10572);
and U11373 (N_11373,N_10095,N_10664);
and U11374 (N_11374,N_10513,N_10863);
nand U11375 (N_11375,N_10431,N_10093);
nand U11376 (N_11376,N_10794,N_10312);
nand U11377 (N_11377,N_10992,N_10061);
nand U11378 (N_11378,N_10497,N_10935);
or U11379 (N_11379,N_10348,N_10554);
nand U11380 (N_11380,N_10783,N_10728);
xor U11381 (N_11381,N_10838,N_10539);
xnor U11382 (N_11382,N_10143,N_10634);
and U11383 (N_11383,N_10707,N_10695);
nor U11384 (N_11384,N_10036,N_10056);
or U11385 (N_11385,N_10635,N_10291);
nor U11386 (N_11386,N_10458,N_10607);
xnor U11387 (N_11387,N_10588,N_10989);
nor U11388 (N_11388,N_10726,N_10910);
nor U11389 (N_11389,N_10737,N_10073);
xnor U11390 (N_11390,N_10117,N_10487);
or U11391 (N_11391,N_10366,N_10674);
xnor U11392 (N_11392,N_10065,N_10374);
and U11393 (N_11393,N_10456,N_10459);
and U11394 (N_11394,N_10248,N_10198);
nor U11395 (N_11395,N_10300,N_10341);
nand U11396 (N_11396,N_10907,N_10923);
nand U11397 (N_11397,N_10449,N_10631);
or U11398 (N_11398,N_10092,N_10214);
nand U11399 (N_11399,N_10110,N_10615);
or U11400 (N_11400,N_10995,N_10697);
nand U11401 (N_11401,N_10754,N_10668);
or U11402 (N_11402,N_10486,N_10467);
nand U11403 (N_11403,N_10232,N_10596);
nand U11404 (N_11404,N_10876,N_10400);
and U11405 (N_11405,N_10581,N_10164);
and U11406 (N_11406,N_10490,N_10028);
or U11407 (N_11407,N_10468,N_10162);
and U11408 (N_11408,N_10562,N_10806);
nand U11409 (N_11409,N_10979,N_10873);
and U11410 (N_11410,N_10566,N_10789);
nand U11411 (N_11411,N_10948,N_10535);
or U11412 (N_11412,N_10057,N_10661);
xor U11413 (N_11413,N_10966,N_10798);
nand U11414 (N_11414,N_10830,N_10152);
xnor U11415 (N_11415,N_10041,N_10159);
nand U11416 (N_11416,N_10447,N_10101);
or U11417 (N_11417,N_10306,N_10900);
nand U11418 (N_11418,N_10805,N_10455);
nor U11419 (N_11419,N_10610,N_10324);
nand U11420 (N_11420,N_10206,N_10382);
xor U11421 (N_11421,N_10212,N_10103);
and U11422 (N_11422,N_10189,N_10153);
and U11423 (N_11423,N_10024,N_10394);
nor U11424 (N_11424,N_10522,N_10766);
or U11425 (N_11425,N_10288,N_10485);
and U11426 (N_11426,N_10419,N_10144);
or U11427 (N_11427,N_10116,N_10780);
xnor U11428 (N_11428,N_10142,N_10343);
or U11429 (N_11429,N_10165,N_10877);
nand U11430 (N_11430,N_10710,N_10705);
xnor U11431 (N_11431,N_10084,N_10237);
xor U11432 (N_11432,N_10722,N_10575);
xor U11433 (N_11433,N_10235,N_10725);
and U11434 (N_11434,N_10756,N_10135);
xor U11435 (N_11435,N_10253,N_10580);
xnor U11436 (N_11436,N_10650,N_10138);
xnor U11437 (N_11437,N_10752,N_10399);
xor U11438 (N_11438,N_10889,N_10215);
or U11439 (N_11439,N_10292,N_10928);
nand U11440 (N_11440,N_10375,N_10156);
and U11441 (N_11441,N_10130,N_10791);
and U11442 (N_11442,N_10887,N_10944);
nand U11443 (N_11443,N_10299,N_10598);
xnor U11444 (N_11444,N_10167,N_10652);
xnor U11445 (N_11445,N_10160,N_10525);
or U11446 (N_11446,N_10585,N_10803);
nand U11447 (N_11447,N_10627,N_10804);
xnor U11448 (N_11448,N_10182,N_10640);
xor U11449 (N_11449,N_10673,N_10105);
and U11450 (N_11450,N_10968,N_10427);
nor U11451 (N_11451,N_10506,N_10963);
nor U11452 (N_11452,N_10119,N_10395);
xnor U11453 (N_11453,N_10077,N_10268);
nand U11454 (N_11454,N_10808,N_10934);
xnor U11455 (N_11455,N_10778,N_10148);
nor U11456 (N_11456,N_10150,N_10128);
or U11457 (N_11457,N_10115,N_10753);
or U11458 (N_11458,N_10284,N_10978);
nor U11459 (N_11459,N_10464,N_10746);
or U11460 (N_11460,N_10682,N_10344);
and U11461 (N_11461,N_10313,N_10002);
xnor U11462 (N_11462,N_10622,N_10557);
nand U11463 (N_11463,N_10942,N_10849);
or U11464 (N_11464,N_10277,N_10349);
nor U11465 (N_11465,N_10011,N_10398);
xor U11466 (N_11466,N_10090,N_10438);
nor U11467 (N_11467,N_10147,N_10478);
or U11468 (N_11468,N_10019,N_10761);
or U11469 (N_11469,N_10435,N_10604);
nor U11470 (N_11470,N_10063,N_10626);
or U11471 (N_11471,N_10470,N_10122);
and U11472 (N_11472,N_10030,N_10307);
or U11473 (N_11473,N_10696,N_10205);
nand U11474 (N_11474,N_10308,N_10086);
xnor U11475 (N_11475,N_10583,N_10228);
or U11476 (N_11476,N_10222,N_10946);
xor U11477 (N_11477,N_10484,N_10445);
or U11478 (N_11478,N_10629,N_10249);
nand U11479 (N_11479,N_10758,N_10792);
xnor U11480 (N_11480,N_10026,N_10986);
nor U11481 (N_11481,N_10686,N_10540);
and U11482 (N_11482,N_10218,N_10457);
nand U11483 (N_11483,N_10371,N_10785);
nand U11484 (N_11484,N_10042,N_10100);
nand U11485 (N_11485,N_10471,N_10040);
xnor U11486 (N_11486,N_10905,N_10256);
nor U11487 (N_11487,N_10867,N_10386);
xnor U11488 (N_11488,N_10425,N_10365);
or U11489 (N_11489,N_10834,N_10965);
and U11490 (N_11490,N_10076,N_10709);
or U11491 (N_11491,N_10677,N_10390);
nor U11492 (N_11492,N_10006,N_10266);
xnor U11493 (N_11493,N_10010,N_10546);
and U11494 (N_11494,N_10912,N_10275);
nor U11495 (N_11495,N_10211,N_10051);
and U11496 (N_11496,N_10680,N_10001);
nand U11497 (N_11497,N_10003,N_10747);
or U11498 (N_11498,N_10204,N_10730);
xnor U11499 (N_11499,N_10683,N_10219);
or U11500 (N_11500,N_10099,N_10749);
xor U11501 (N_11501,N_10991,N_10782);
or U11502 (N_11502,N_10480,N_10558);
and U11503 (N_11503,N_10631,N_10926);
nor U11504 (N_11504,N_10983,N_10497);
and U11505 (N_11505,N_10772,N_10494);
or U11506 (N_11506,N_10836,N_10807);
nand U11507 (N_11507,N_10786,N_10799);
nor U11508 (N_11508,N_10001,N_10317);
nor U11509 (N_11509,N_10323,N_10014);
nand U11510 (N_11510,N_10109,N_10594);
nor U11511 (N_11511,N_10055,N_10460);
or U11512 (N_11512,N_10768,N_10691);
xnor U11513 (N_11513,N_10129,N_10006);
nor U11514 (N_11514,N_10461,N_10886);
and U11515 (N_11515,N_10468,N_10362);
or U11516 (N_11516,N_10974,N_10047);
nor U11517 (N_11517,N_10225,N_10802);
nor U11518 (N_11518,N_10455,N_10551);
or U11519 (N_11519,N_10742,N_10602);
xor U11520 (N_11520,N_10414,N_10722);
nand U11521 (N_11521,N_10163,N_10958);
and U11522 (N_11522,N_10931,N_10562);
nand U11523 (N_11523,N_10107,N_10507);
xnor U11524 (N_11524,N_10173,N_10109);
xor U11525 (N_11525,N_10720,N_10985);
xor U11526 (N_11526,N_10192,N_10122);
or U11527 (N_11527,N_10353,N_10701);
xor U11528 (N_11528,N_10662,N_10126);
and U11529 (N_11529,N_10792,N_10628);
nand U11530 (N_11530,N_10620,N_10310);
or U11531 (N_11531,N_10147,N_10898);
or U11532 (N_11532,N_10478,N_10364);
and U11533 (N_11533,N_10289,N_10164);
xor U11534 (N_11534,N_10740,N_10580);
nor U11535 (N_11535,N_10730,N_10448);
or U11536 (N_11536,N_10522,N_10229);
xor U11537 (N_11537,N_10545,N_10383);
xor U11538 (N_11538,N_10756,N_10171);
xor U11539 (N_11539,N_10625,N_10827);
and U11540 (N_11540,N_10066,N_10334);
nor U11541 (N_11541,N_10296,N_10013);
and U11542 (N_11542,N_10308,N_10343);
xor U11543 (N_11543,N_10435,N_10788);
xor U11544 (N_11544,N_10154,N_10662);
or U11545 (N_11545,N_10596,N_10279);
or U11546 (N_11546,N_10385,N_10719);
nor U11547 (N_11547,N_10314,N_10718);
nor U11548 (N_11548,N_10370,N_10842);
and U11549 (N_11549,N_10764,N_10462);
and U11550 (N_11550,N_10314,N_10722);
or U11551 (N_11551,N_10906,N_10258);
nor U11552 (N_11552,N_10952,N_10313);
and U11553 (N_11553,N_10515,N_10140);
xnor U11554 (N_11554,N_10526,N_10581);
nand U11555 (N_11555,N_10299,N_10346);
nand U11556 (N_11556,N_10295,N_10364);
xnor U11557 (N_11557,N_10643,N_10652);
xor U11558 (N_11558,N_10580,N_10737);
nor U11559 (N_11559,N_10610,N_10075);
or U11560 (N_11560,N_10039,N_10468);
or U11561 (N_11561,N_10325,N_10631);
and U11562 (N_11562,N_10973,N_10803);
nand U11563 (N_11563,N_10964,N_10154);
nand U11564 (N_11564,N_10407,N_10928);
and U11565 (N_11565,N_10973,N_10852);
or U11566 (N_11566,N_10277,N_10211);
nor U11567 (N_11567,N_10864,N_10417);
or U11568 (N_11568,N_10603,N_10229);
or U11569 (N_11569,N_10207,N_10328);
and U11570 (N_11570,N_10427,N_10941);
nor U11571 (N_11571,N_10088,N_10829);
and U11572 (N_11572,N_10970,N_10048);
nand U11573 (N_11573,N_10516,N_10448);
and U11574 (N_11574,N_10435,N_10951);
nand U11575 (N_11575,N_10886,N_10531);
nand U11576 (N_11576,N_10206,N_10168);
nor U11577 (N_11577,N_10737,N_10550);
nor U11578 (N_11578,N_10397,N_10653);
xnor U11579 (N_11579,N_10006,N_10462);
or U11580 (N_11580,N_10153,N_10548);
xnor U11581 (N_11581,N_10544,N_10547);
nor U11582 (N_11582,N_10233,N_10763);
and U11583 (N_11583,N_10213,N_10016);
nand U11584 (N_11584,N_10211,N_10564);
nor U11585 (N_11585,N_10943,N_10048);
and U11586 (N_11586,N_10305,N_10333);
and U11587 (N_11587,N_10882,N_10472);
xor U11588 (N_11588,N_10644,N_10223);
nand U11589 (N_11589,N_10068,N_10623);
nand U11590 (N_11590,N_10497,N_10387);
xnor U11591 (N_11591,N_10528,N_10172);
nand U11592 (N_11592,N_10903,N_10997);
nor U11593 (N_11593,N_10188,N_10046);
or U11594 (N_11594,N_10109,N_10262);
or U11595 (N_11595,N_10397,N_10890);
or U11596 (N_11596,N_10737,N_10793);
nand U11597 (N_11597,N_10573,N_10327);
or U11598 (N_11598,N_10502,N_10782);
or U11599 (N_11599,N_10901,N_10384);
xnor U11600 (N_11600,N_10982,N_10183);
xnor U11601 (N_11601,N_10004,N_10185);
or U11602 (N_11602,N_10682,N_10989);
and U11603 (N_11603,N_10118,N_10424);
xnor U11604 (N_11604,N_10018,N_10799);
or U11605 (N_11605,N_10080,N_10235);
nor U11606 (N_11606,N_10945,N_10702);
nand U11607 (N_11607,N_10670,N_10425);
nor U11608 (N_11608,N_10821,N_10973);
xor U11609 (N_11609,N_10052,N_10641);
and U11610 (N_11610,N_10247,N_10647);
and U11611 (N_11611,N_10748,N_10422);
xor U11612 (N_11612,N_10883,N_10067);
nand U11613 (N_11613,N_10425,N_10988);
nand U11614 (N_11614,N_10062,N_10613);
or U11615 (N_11615,N_10616,N_10958);
nor U11616 (N_11616,N_10438,N_10254);
and U11617 (N_11617,N_10866,N_10284);
nand U11618 (N_11618,N_10826,N_10947);
and U11619 (N_11619,N_10509,N_10833);
or U11620 (N_11620,N_10964,N_10410);
nand U11621 (N_11621,N_10497,N_10704);
nand U11622 (N_11622,N_10944,N_10769);
nor U11623 (N_11623,N_10711,N_10409);
and U11624 (N_11624,N_10203,N_10794);
nor U11625 (N_11625,N_10927,N_10639);
xnor U11626 (N_11626,N_10957,N_10038);
and U11627 (N_11627,N_10609,N_10409);
and U11628 (N_11628,N_10106,N_10305);
nor U11629 (N_11629,N_10627,N_10439);
nor U11630 (N_11630,N_10883,N_10058);
and U11631 (N_11631,N_10354,N_10273);
and U11632 (N_11632,N_10243,N_10204);
and U11633 (N_11633,N_10038,N_10613);
nor U11634 (N_11634,N_10991,N_10860);
or U11635 (N_11635,N_10666,N_10000);
nand U11636 (N_11636,N_10893,N_10319);
or U11637 (N_11637,N_10805,N_10596);
and U11638 (N_11638,N_10074,N_10136);
and U11639 (N_11639,N_10807,N_10914);
and U11640 (N_11640,N_10890,N_10387);
nor U11641 (N_11641,N_10732,N_10896);
nor U11642 (N_11642,N_10120,N_10971);
nor U11643 (N_11643,N_10595,N_10222);
and U11644 (N_11644,N_10053,N_10074);
nand U11645 (N_11645,N_10922,N_10480);
nor U11646 (N_11646,N_10855,N_10732);
and U11647 (N_11647,N_10356,N_10601);
nor U11648 (N_11648,N_10549,N_10661);
and U11649 (N_11649,N_10169,N_10661);
and U11650 (N_11650,N_10439,N_10769);
or U11651 (N_11651,N_10931,N_10513);
or U11652 (N_11652,N_10053,N_10402);
and U11653 (N_11653,N_10577,N_10711);
and U11654 (N_11654,N_10803,N_10194);
or U11655 (N_11655,N_10743,N_10334);
and U11656 (N_11656,N_10032,N_10100);
or U11657 (N_11657,N_10373,N_10498);
nand U11658 (N_11658,N_10637,N_10058);
nand U11659 (N_11659,N_10472,N_10387);
and U11660 (N_11660,N_10641,N_10491);
or U11661 (N_11661,N_10252,N_10273);
nor U11662 (N_11662,N_10008,N_10536);
and U11663 (N_11663,N_10092,N_10078);
xor U11664 (N_11664,N_10365,N_10968);
xnor U11665 (N_11665,N_10962,N_10307);
nor U11666 (N_11666,N_10862,N_10744);
xor U11667 (N_11667,N_10365,N_10222);
xor U11668 (N_11668,N_10492,N_10968);
xor U11669 (N_11669,N_10597,N_10438);
xnor U11670 (N_11670,N_10428,N_10376);
or U11671 (N_11671,N_10717,N_10097);
nand U11672 (N_11672,N_10756,N_10862);
or U11673 (N_11673,N_10224,N_10202);
nor U11674 (N_11674,N_10435,N_10533);
nor U11675 (N_11675,N_10515,N_10207);
nand U11676 (N_11676,N_10959,N_10100);
or U11677 (N_11677,N_10341,N_10718);
or U11678 (N_11678,N_10236,N_10631);
nor U11679 (N_11679,N_10049,N_10363);
and U11680 (N_11680,N_10919,N_10399);
nor U11681 (N_11681,N_10519,N_10558);
and U11682 (N_11682,N_10755,N_10924);
nor U11683 (N_11683,N_10867,N_10046);
nor U11684 (N_11684,N_10895,N_10883);
and U11685 (N_11685,N_10806,N_10675);
and U11686 (N_11686,N_10158,N_10830);
or U11687 (N_11687,N_10628,N_10507);
xnor U11688 (N_11688,N_10084,N_10777);
xnor U11689 (N_11689,N_10131,N_10832);
xnor U11690 (N_11690,N_10403,N_10945);
xnor U11691 (N_11691,N_10288,N_10096);
or U11692 (N_11692,N_10129,N_10333);
and U11693 (N_11693,N_10500,N_10802);
nor U11694 (N_11694,N_10064,N_10556);
and U11695 (N_11695,N_10980,N_10362);
xnor U11696 (N_11696,N_10747,N_10422);
or U11697 (N_11697,N_10688,N_10827);
nand U11698 (N_11698,N_10283,N_10882);
or U11699 (N_11699,N_10870,N_10893);
or U11700 (N_11700,N_10394,N_10552);
nor U11701 (N_11701,N_10772,N_10770);
nor U11702 (N_11702,N_10415,N_10210);
xnor U11703 (N_11703,N_10495,N_10672);
or U11704 (N_11704,N_10385,N_10595);
nand U11705 (N_11705,N_10930,N_10038);
xnor U11706 (N_11706,N_10528,N_10494);
nand U11707 (N_11707,N_10361,N_10729);
nor U11708 (N_11708,N_10493,N_10986);
xnor U11709 (N_11709,N_10617,N_10605);
or U11710 (N_11710,N_10632,N_10590);
xor U11711 (N_11711,N_10836,N_10134);
and U11712 (N_11712,N_10654,N_10346);
nor U11713 (N_11713,N_10168,N_10942);
or U11714 (N_11714,N_10947,N_10870);
nand U11715 (N_11715,N_10574,N_10462);
nor U11716 (N_11716,N_10367,N_10441);
or U11717 (N_11717,N_10686,N_10025);
nand U11718 (N_11718,N_10165,N_10542);
nand U11719 (N_11719,N_10167,N_10089);
nor U11720 (N_11720,N_10796,N_10739);
nand U11721 (N_11721,N_10428,N_10261);
nand U11722 (N_11722,N_10066,N_10838);
and U11723 (N_11723,N_10732,N_10058);
nor U11724 (N_11724,N_10898,N_10294);
nor U11725 (N_11725,N_10997,N_10654);
or U11726 (N_11726,N_10922,N_10673);
xor U11727 (N_11727,N_10733,N_10214);
and U11728 (N_11728,N_10692,N_10580);
nand U11729 (N_11729,N_10887,N_10255);
or U11730 (N_11730,N_10879,N_10632);
and U11731 (N_11731,N_10819,N_10627);
nand U11732 (N_11732,N_10192,N_10955);
nor U11733 (N_11733,N_10596,N_10696);
and U11734 (N_11734,N_10011,N_10133);
or U11735 (N_11735,N_10897,N_10678);
nand U11736 (N_11736,N_10822,N_10638);
nor U11737 (N_11737,N_10136,N_10063);
nand U11738 (N_11738,N_10728,N_10033);
xor U11739 (N_11739,N_10342,N_10196);
xor U11740 (N_11740,N_10513,N_10446);
nor U11741 (N_11741,N_10506,N_10424);
and U11742 (N_11742,N_10846,N_10896);
and U11743 (N_11743,N_10738,N_10051);
nor U11744 (N_11744,N_10827,N_10049);
nor U11745 (N_11745,N_10796,N_10346);
nor U11746 (N_11746,N_10219,N_10053);
xnor U11747 (N_11747,N_10979,N_10566);
nand U11748 (N_11748,N_10515,N_10913);
or U11749 (N_11749,N_10955,N_10233);
or U11750 (N_11750,N_10988,N_10118);
nand U11751 (N_11751,N_10544,N_10959);
nor U11752 (N_11752,N_10915,N_10341);
or U11753 (N_11753,N_10332,N_10638);
nand U11754 (N_11754,N_10156,N_10832);
xor U11755 (N_11755,N_10600,N_10812);
or U11756 (N_11756,N_10464,N_10036);
nand U11757 (N_11757,N_10519,N_10979);
nor U11758 (N_11758,N_10889,N_10318);
xor U11759 (N_11759,N_10578,N_10910);
nor U11760 (N_11760,N_10336,N_10309);
nor U11761 (N_11761,N_10392,N_10511);
or U11762 (N_11762,N_10806,N_10195);
and U11763 (N_11763,N_10818,N_10035);
and U11764 (N_11764,N_10448,N_10351);
or U11765 (N_11765,N_10065,N_10246);
and U11766 (N_11766,N_10234,N_10528);
nand U11767 (N_11767,N_10159,N_10396);
and U11768 (N_11768,N_10184,N_10927);
nand U11769 (N_11769,N_10704,N_10346);
xor U11770 (N_11770,N_10330,N_10854);
and U11771 (N_11771,N_10300,N_10658);
xor U11772 (N_11772,N_10901,N_10781);
nor U11773 (N_11773,N_10339,N_10713);
nor U11774 (N_11774,N_10470,N_10637);
and U11775 (N_11775,N_10688,N_10796);
and U11776 (N_11776,N_10631,N_10235);
and U11777 (N_11777,N_10233,N_10878);
nor U11778 (N_11778,N_10417,N_10670);
nand U11779 (N_11779,N_10566,N_10549);
nor U11780 (N_11780,N_10335,N_10817);
nor U11781 (N_11781,N_10571,N_10854);
nor U11782 (N_11782,N_10695,N_10914);
and U11783 (N_11783,N_10976,N_10920);
nand U11784 (N_11784,N_10432,N_10202);
xor U11785 (N_11785,N_10226,N_10488);
xor U11786 (N_11786,N_10014,N_10442);
xnor U11787 (N_11787,N_10895,N_10990);
nor U11788 (N_11788,N_10121,N_10353);
nand U11789 (N_11789,N_10699,N_10074);
or U11790 (N_11790,N_10971,N_10022);
xnor U11791 (N_11791,N_10028,N_10391);
and U11792 (N_11792,N_10406,N_10029);
and U11793 (N_11793,N_10349,N_10480);
nand U11794 (N_11794,N_10407,N_10122);
xor U11795 (N_11795,N_10661,N_10769);
or U11796 (N_11796,N_10963,N_10916);
xor U11797 (N_11797,N_10582,N_10563);
and U11798 (N_11798,N_10334,N_10258);
and U11799 (N_11799,N_10438,N_10611);
or U11800 (N_11800,N_10412,N_10665);
nor U11801 (N_11801,N_10897,N_10966);
or U11802 (N_11802,N_10649,N_10662);
nand U11803 (N_11803,N_10297,N_10277);
xnor U11804 (N_11804,N_10784,N_10134);
and U11805 (N_11805,N_10306,N_10856);
or U11806 (N_11806,N_10432,N_10381);
nand U11807 (N_11807,N_10505,N_10173);
and U11808 (N_11808,N_10135,N_10854);
nand U11809 (N_11809,N_10453,N_10017);
or U11810 (N_11810,N_10178,N_10540);
xnor U11811 (N_11811,N_10613,N_10245);
nor U11812 (N_11812,N_10016,N_10388);
nand U11813 (N_11813,N_10082,N_10579);
xnor U11814 (N_11814,N_10848,N_10204);
nor U11815 (N_11815,N_10071,N_10341);
nand U11816 (N_11816,N_10016,N_10171);
nand U11817 (N_11817,N_10926,N_10103);
or U11818 (N_11818,N_10643,N_10059);
or U11819 (N_11819,N_10445,N_10229);
xnor U11820 (N_11820,N_10897,N_10956);
xnor U11821 (N_11821,N_10081,N_10213);
nand U11822 (N_11822,N_10939,N_10886);
nor U11823 (N_11823,N_10659,N_10778);
nand U11824 (N_11824,N_10600,N_10864);
or U11825 (N_11825,N_10619,N_10830);
and U11826 (N_11826,N_10629,N_10313);
and U11827 (N_11827,N_10412,N_10140);
nor U11828 (N_11828,N_10975,N_10773);
or U11829 (N_11829,N_10352,N_10018);
or U11830 (N_11830,N_10215,N_10385);
nand U11831 (N_11831,N_10681,N_10706);
xnor U11832 (N_11832,N_10971,N_10788);
nand U11833 (N_11833,N_10747,N_10525);
nand U11834 (N_11834,N_10208,N_10282);
or U11835 (N_11835,N_10177,N_10359);
nor U11836 (N_11836,N_10618,N_10289);
xnor U11837 (N_11837,N_10892,N_10949);
nand U11838 (N_11838,N_10007,N_10335);
xnor U11839 (N_11839,N_10109,N_10609);
nand U11840 (N_11840,N_10429,N_10995);
nor U11841 (N_11841,N_10385,N_10750);
xor U11842 (N_11842,N_10099,N_10128);
xnor U11843 (N_11843,N_10749,N_10715);
xnor U11844 (N_11844,N_10921,N_10908);
or U11845 (N_11845,N_10159,N_10767);
and U11846 (N_11846,N_10134,N_10224);
or U11847 (N_11847,N_10745,N_10890);
or U11848 (N_11848,N_10234,N_10600);
or U11849 (N_11849,N_10886,N_10505);
xnor U11850 (N_11850,N_10296,N_10505);
nor U11851 (N_11851,N_10018,N_10492);
or U11852 (N_11852,N_10180,N_10937);
and U11853 (N_11853,N_10329,N_10502);
xnor U11854 (N_11854,N_10604,N_10898);
nand U11855 (N_11855,N_10522,N_10241);
nor U11856 (N_11856,N_10120,N_10684);
xnor U11857 (N_11857,N_10378,N_10760);
nor U11858 (N_11858,N_10268,N_10419);
or U11859 (N_11859,N_10368,N_10723);
or U11860 (N_11860,N_10495,N_10039);
or U11861 (N_11861,N_10966,N_10910);
nand U11862 (N_11862,N_10777,N_10662);
and U11863 (N_11863,N_10836,N_10859);
and U11864 (N_11864,N_10554,N_10761);
and U11865 (N_11865,N_10570,N_10426);
xor U11866 (N_11866,N_10623,N_10151);
or U11867 (N_11867,N_10691,N_10336);
nor U11868 (N_11868,N_10019,N_10234);
and U11869 (N_11869,N_10271,N_10926);
nand U11870 (N_11870,N_10274,N_10975);
xnor U11871 (N_11871,N_10938,N_10934);
nor U11872 (N_11872,N_10132,N_10944);
or U11873 (N_11873,N_10469,N_10982);
or U11874 (N_11874,N_10907,N_10438);
nand U11875 (N_11875,N_10461,N_10462);
and U11876 (N_11876,N_10847,N_10751);
and U11877 (N_11877,N_10512,N_10232);
nor U11878 (N_11878,N_10615,N_10697);
or U11879 (N_11879,N_10453,N_10531);
xnor U11880 (N_11880,N_10098,N_10874);
nor U11881 (N_11881,N_10810,N_10741);
nand U11882 (N_11882,N_10538,N_10976);
and U11883 (N_11883,N_10809,N_10555);
nor U11884 (N_11884,N_10684,N_10482);
nand U11885 (N_11885,N_10888,N_10608);
xor U11886 (N_11886,N_10443,N_10804);
or U11887 (N_11887,N_10324,N_10199);
nand U11888 (N_11888,N_10540,N_10353);
and U11889 (N_11889,N_10455,N_10494);
xor U11890 (N_11890,N_10011,N_10016);
and U11891 (N_11891,N_10612,N_10846);
and U11892 (N_11892,N_10959,N_10467);
xor U11893 (N_11893,N_10735,N_10181);
xnor U11894 (N_11894,N_10495,N_10736);
or U11895 (N_11895,N_10472,N_10590);
or U11896 (N_11896,N_10780,N_10037);
nand U11897 (N_11897,N_10815,N_10691);
and U11898 (N_11898,N_10871,N_10866);
nor U11899 (N_11899,N_10074,N_10166);
nand U11900 (N_11900,N_10966,N_10436);
xnor U11901 (N_11901,N_10458,N_10897);
nand U11902 (N_11902,N_10974,N_10367);
or U11903 (N_11903,N_10413,N_10528);
xnor U11904 (N_11904,N_10320,N_10682);
or U11905 (N_11905,N_10413,N_10925);
xor U11906 (N_11906,N_10259,N_10873);
xnor U11907 (N_11907,N_10911,N_10479);
or U11908 (N_11908,N_10072,N_10205);
or U11909 (N_11909,N_10414,N_10363);
and U11910 (N_11910,N_10889,N_10061);
nand U11911 (N_11911,N_10614,N_10950);
xor U11912 (N_11912,N_10562,N_10561);
xnor U11913 (N_11913,N_10500,N_10974);
xnor U11914 (N_11914,N_10110,N_10795);
or U11915 (N_11915,N_10295,N_10722);
nor U11916 (N_11916,N_10340,N_10442);
or U11917 (N_11917,N_10722,N_10772);
and U11918 (N_11918,N_10408,N_10328);
or U11919 (N_11919,N_10040,N_10540);
or U11920 (N_11920,N_10250,N_10285);
xor U11921 (N_11921,N_10870,N_10898);
nor U11922 (N_11922,N_10178,N_10985);
and U11923 (N_11923,N_10203,N_10673);
or U11924 (N_11924,N_10778,N_10270);
nor U11925 (N_11925,N_10160,N_10424);
or U11926 (N_11926,N_10138,N_10991);
xor U11927 (N_11927,N_10443,N_10192);
nand U11928 (N_11928,N_10648,N_10625);
xnor U11929 (N_11929,N_10858,N_10355);
or U11930 (N_11930,N_10906,N_10766);
and U11931 (N_11931,N_10789,N_10140);
nor U11932 (N_11932,N_10987,N_10014);
and U11933 (N_11933,N_10912,N_10964);
and U11934 (N_11934,N_10029,N_10461);
and U11935 (N_11935,N_10206,N_10968);
or U11936 (N_11936,N_10568,N_10202);
nor U11937 (N_11937,N_10810,N_10728);
and U11938 (N_11938,N_10509,N_10345);
or U11939 (N_11939,N_10465,N_10417);
and U11940 (N_11940,N_10097,N_10104);
xor U11941 (N_11941,N_10005,N_10381);
nand U11942 (N_11942,N_10950,N_10779);
nor U11943 (N_11943,N_10878,N_10855);
nand U11944 (N_11944,N_10662,N_10274);
and U11945 (N_11945,N_10964,N_10893);
nand U11946 (N_11946,N_10567,N_10461);
nand U11947 (N_11947,N_10130,N_10009);
nor U11948 (N_11948,N_10322,N_10402);
xor U11949 (N_11949,N_10832,N_10317);
and U11950 (N_11950,N_10938,N_10388);
nor U11951 (N_11951,N_10501,N_10461);
or U11952 (N_11952,N_10214,N_10682);
xnor U11953 (N_11953,N_10322,N_10128);
nor U11954 (N_11954,N_10584,N_10674);
nand U11955 (N_11955,N_10014,N_10785);
xor U11956 (N_11956,N_10057,N_10255);
nor U11957 (N_11957,N_10103,N_10179);
nand U11958 (N_11958,N_10590,N_10271);
or U11959 (N_11959,N_10423,N_10925);
and U11960 (N_11960,N_10542,N_10229);
xnor U11961 (N_11961,N_10535,N_10581);
nand U11962 (N_11962,N_10580,N_10694);
nand U11963 (N_11963,N_10942,N_10493);
and U11964 (N_11964,N_10029,N_10882);
nor U11965 (N_11965,N_10050,N_10601);
and U11966 (N_11966,N_10662,N_10239);
nor U11967 (N_11967,N_10682,N_10445);
nor U11968 (N_11968,N_10629,N_10495);
nand U11969 (N_11969,N_10921,N_10540);
nand U11970 (N_11970,N_10784,N_10828);
nor U11971 (N_11971,N_10533,N_10178);
nor U11972 (N_11972,N_10175,N_10582);
xnor U11973 (N_11973,N_10689,N_10185);
and U11974 (N_11974,N_10460,N_10769);
xor U11975 (N_11975,N_10961,N_10227);
nand U11976 (N_11976,N_10719,N_10734);
xor U11977 (N_11977,N_10691,N_10007);
or U11978 (N_11978,N_10739,N_10564);
nor U11979 (N_11979,N_10671,N_10674);
nand U11980 (N_11980,N_10031,N_10595);
nor U11981 (N_11981,N_10435,N_10552);
and U11982 (N_11982,N_10269,N_10869);
nor U11983 (N_11983,N_10973,N_10392);
or U11984 (N_11984,N_10114,N_10118);
and U11985 (N_11985,N_10129,N_10641);
or U11986 (N_11986,N_10980,N_10004);
nand U11987 (N_11987,N_10191,N_10302);
or U11988 (N_11988,N_10159,N_10801);
or U11989 (N_11989,N_10179,N_10217);
nor U11990 (N_11990,N_10993,N_10638);
nand U11991 (N_11991,N_10958,N_10258);
xor U11992 (N_11992,N_10789,N_10183);
nor U11993 (N_11993,N_10880,N_10610);
nand U11994 (N_11994,N_10834,N_10710);
nand U11995 (N_11995,N_10234,N_10562);
and U11996 (N_11996,N_10375,N_10309);
nand U11997 (N_11997,N_10379,N_10252);
xnor U11998 (N_11998,N_10268,N_10870);
or U11999 (N_11999,N_10985,N_10762);
and U12000 (N_12000,N_11274,N_11528);
or U12001 (N_12001,N_11774,N_11604);
or U12002 (N_12002,N_11179,N_11969);
nor U12003 (N_12003,N_11278,N_11159);
or U12004 (N_12004,N_11875,N_11061);
xor U12005 (N_12005,N_11117,N_11699);
xor U12006 (N_12006,N_11230,N_11880);
and U12007 (N_12007,N_11867,N_11131);
or U12008 (N_12008,N_11817,N_11458);
nand U12009 (N_12009,N_11432,N_11563);
nor U12010 (N_12010,N_11657,N_11452);
and U12011 (N_12011,N_11894,N_11222);
nor U12012 (N_12012,N_11918,N_11929);
nand U12013 (N_12013,N_11508,N_11122);
nand U12014 (N_12014,N_11393,N_11441);
nand U12015 (N_12015,N_11749,N_11794);
nor U12016 (N_12016,N_11390,N_11013);
xor U12017 (N_12017,N_11654,N_11669);
or U12018 (N_12018,N_11414,N_11132);
or U12019 (N_12019,N_11134,N_11087);
nor U12020 (N_12020,N_11700,N_11833);
nand U12021 (N_12021,N_11124,N_11188);
xor U12022 (N_12022,N_11961,N_11262);
xor U12023 (N_12023,N_11693,N_11183);
or U12024 (N_12024,N_11944,N_11678);
nor U12025 (N_12025,N_11307,N_11440);
and U12026 (N_12026,N_11586,N_11849);
nor U12027 (N_12027,N_11315,N_11583);
nor U12028 (N_12028,N_11778,N_11896);
xor U12029 (N_12029,N_11351,N_11069);
nor U12030 (N_12030,N_11627,N_11852);
nor U12031 (N_12031,N_11858,N_11234);
or U12032 (N_12032,N_11769,N_11493);
nor U12033 (N_12033,N_11316,N_11513);
and U12034 (N_12034,N_11067,N_11265);
or U12035 (N_12035,N_11406,N_11320);
or U12036 (N_12036,N_11339,N_11031);
or U12037 (N_12037,N_11254,N_11088);
nor U12038 (N_12038,N_11812,N_11506);
or U12039 (N_12039,N_11281,N_11670);
or U12040 (N_12040,N_11890,N_11377);
xor U12041 (N_12041,N_11856,N_11287);
xnor U12042 (N_12042,N_11569,N_11327);
nand U12043 (N_12043,N_11156,N_11555);
nand U12044 (N_12044,N_11611,N_11802);
and U12045 (N_12045,N_11871,N_11859);
nand U12046 (N_12046,N_11803,N_11570);
and U12047 (N_12047,N_11063,N_11497);
xnor U12048 (N_12048,N_11838,N_11359);
and U12049 (N_12049,N_11261,N_11834);
or U12050 (N_12050,N_11799,N_11864);
xor U12051 (N_12051,N_11048,N_11394);
xor U12052 (N_12052,N_11863,N_11163);
nor U12053 (N_12053,N_11908,N_11939);
and U12054 (N_12054,N_11155,N_11781);
nand U12055 (N_12055,N_11387,N_11072);
and U12056 (N_12056,N_11362,N_11522);
nand U12057 (N_12057,N_11417,N_11358);
xnor U12058 (N_12058,N_11488,N_11957);
nor U12059 (N_12059,N_11715,N_11425);
xnor U12060 (N_12060,N_11285,N_11973);
nor U12061 (N_12061,N_11819,N_11951);
nor U12062 (N_12062,N_11956,N_11851);
nor U12063 (N_12063,N_11053,N_11972);
nand U12064 (N_12064,N_11845,N_11151);
nand U12065 (N_12065,N_11244,N_11797);
and U12066 (N_12066,N_11688,N_11275);
and U12067 (N_12067,N_11444,N_11930);
nand U12068 (N_12068,N_11130,N_11631);
or U12069 (N_12069,N_11109,N_11346);
xnor U12070 (N_12070,N_11223,N_11753);
nand U12071 (N_12071,N_11897,N_11696);
xor U12072 (N_12072,N_11750,N_11347);
or U12073 (N_12073,N_11104,N_11800);
and U12074 (N_12074,N_11581,N_11165);
nand U12075 (N_12075,N_11991,N_11399);
xor U12076 (N_12076,N_11364,N_11567);
xnor U12077 (N_12077,N_11577,N_11735);
nand U12078 (N_12078,N_11267,N_11883);
xnor U12079 (N_12079,N_11879,N_11355);
xnor U12080 (N_12080,N_11807,N_11202);
xor U12081 (N_12081,N_11143,N_11025);
nor U12082 (N_12082,N_11723,N_11614);
or U12083 (N_12083,N_11184,N_11256);
nand U12084 (N_12084,N_11617,N_11332);
xnor U12085 (N_12085,N_11129,N_11153);
nor U12086 (N_12086,N_11509,N_11588);
nand U12087 (N_12087,N_11822,N_11695);
and U12088 (N_12088,N_11469,N_11572);
xnor U12089 (N_12089,N_11564,N_11200);
nand U12090 (N_12090,N_11083,N_11643);
nor U12091 (N_12091,N_11292,N_11810);
nand U12092 (N_12092,N_11106,N_11176);
nand U12093 (N_12093,N_11645,N_11692);
nand U12094 (N_12094,N_11895,N_11502);
xnor U12095 (N_12095,N_11997,N_11659);
and U12096 (N_12096,N_11668,N_11789);
or U12097 (N_12097,N_11701,N_11684);
or U12098 (N_12098,N_11095,N_11848);
nor U12099 (N_12099,N_11873,N_11435);
and U12100 (N_12100,N_11021,N_11641);
nand U12101 (N_12101,N_11027,N_11099);
xnor U12102 (N_12102,N_11911,N_11376);
or U12103 (N_12103,N_11736,N_11028);
nor U12104 (N_12104,N_11751,N_11714);
or U12105 (N_12105,N_11058,N_11658);
and U12106 (N_12106,N_11827,N_11330);
nand U12107 (N_12107,N_11809,N_11100);
and U12108 (N_12108,N_11537,N_11640);
xor U12109 (N_12109,N_11733,N_11790);
xnor U12110 (N_12110,N_11514,N_11891);
nor U12111 (N_12111,N_11585,N_11804);
nand U12112 (N_12112,N_11225,N_11589);
and U12113 (N_12113,N_11243,N_11405);
or U12114 (N_12114,N_11385,N_11717);
nand U12115 (N_12115,N_11447,N_11648);
nor U12116 (N_12116,N_11077,N_11326);
and U12117 (N_12117,N_11408,N_11269);
xnor U12118 (N_12118,N_11811,N_11328);
xnor U12119 (N_12119,N_11898,N_11483);
nand U12120 (N_12120,N_11638,N_11599);
nand U12121 (N_12121,N_11980,N_11191);
xor U12122 (N_12122,N_11742,N_11986);
and U12123 (N_12123,N_11372,N_11177);
or U12124 (N_12124,N_11224,N_11283);
nand U12125 (N_12125,N_11312,N_11089);
nand U12126 (N_12126,N_11877,N_11368);
nand U12127 (N_12127,N_11801,N_11665);
and U12128 (N_12128,N_11460,N_11498);
xor U12129 (N_12129,N_11097,N_11039);
and U12130 (N_12130,N_11420,N_11874);
xor U12131 (N_12131,N_11219,N_11722);
or U12132 (N_12132,N_11732,N_11968);
nor U12133 (N_12133,N_11306,N_11207);
or U12134 (N_12134,N_11584,N_11270);
or U12135 (N_12135,N_11002,N_11642);
or U12136 (N_12136,N_11610,N_11870);
or U12137 (N_12137,N_11575,N_11091);
or U12138 (N_12138,N_11015,N_11016);
nand U12139 (N_12139,N_11369,N_11352);
nor U12140 (N_12140,N_11535,N_11562);
xor U12141 (N_12141,N_11724,N_11383);
xnor U12142 (N_12142,N_11304,N_11990);
nand U12143 (N_12143,N_11418,N_11975);
xor U12144 (N_12144,N_11906,N_11303);
nor U12145 (N_12145,N_11996,N_11615);
nor U12146 (N_12146,N_11865,N_11633);
nand U12147 (N_12147,N_11515,N_11853);
and U12148 (N_12148,N_11820,N_11538);
or U12149 (N_12149,N_11152,N_11526);
or U12150 (N_12150,N_11246,N_11211);
nor U12151 (N_12151,N_11671,N_11532);
nand U12152 (N_12152,N_11296,N_11194);
nor U12153 (N_12153,N_11135,N_11938);
nand U12154 (N_12154,N_11601,N_11900);
nand U12155 (N_12155,N_11829,N_11725);
nand U12156 (N_12156,N_11470,N_11210);
nand U12157 (N_12157,N_11030,N_11412);
xnor U12158 (N_12158,N_11279,N_11398);
nor U12159 (N_12159,N_11793,N_11170);
and U12160 (N_12160,N_11719,N_11756);
nand U12161 (N_12161,N_11505,N_11161);
xor U12162 (N_12162,N_11319,N_11338);
or U12163 (N_12163,N_11830,N_11886);
and U12164 (N_12164,N_11913,N_11466);
nor U12165 (N_12165,N_11235,N_11912);
nor U12166 (N_12166,N_11743,N_11345);
or U12167 (N_12167,N_11245,N_11311);
and U12168 (N_12168,N_11689,N_11241);
nand U12169 (N_12169,N_11680,N_11003);
nor U12170 (N_12170,N_11844,N_11098);
nor U12171 (N_12171,N_11409,N_11144);
or U12172 (N_12172,N_11059,N_11545);
xnor U12173 (N_12173,N_11022,N_11373);
nand U12174 (N_12174,N_11836,N_11258);
or U12175 (N_12175,N_11632,N_11998);
nand U12176 (N_12176,N_11828,N_11438);
and U12177 (N_12177,N_11783,N_11560);
and U12178 (N_12178,N_11655,N_11228);
or U12179 (N_12179,N_11374,N_11754);
xnor U12180 (N_12180,N_11321,N_11835);
and U12181 (N_12181,N_11110,N_11388);
or U12182 (N_12182,N_11983,N_11299);
or U12183 (N_12183,N_11363,N_11033);
xor U12184 (N_12184,N_11571,N_11504);
and U12185 (N_12185,N_11391,N_11038);
nand U12186 (N_12186,N_11662,N_11966);
and U12187 (N_12187,N_11952,N_11443);
and U12188 (N_12188,N_11941,N_11901);
xor U12189 (N_12189,N_11251,N_11579);
and U12190 (N_12190,N_11079,N_11909);
nand U12191 (N_12191,N_11381,N_11694);
nand U12192 (N_12192,N_11136,N_11726);
nor U12193 (N_12193,N_11839,N_11910);
nand U12194 (N_12194,N_11557,N_11737);
nor U12195 (N_12195,N_11476,N_11150);
nand U12196 (N_12196,N_11081,N_11185);
xnor U12197 (N_12197,N_11806,N_11268);
nand U12198 (N_12198,N_11960,N_11430);
or U12199 (N_12199,N_11962,N_11550);
and U12200 (N_12200,N_11066,N_11423);
nor U12201 (N_12201,N_11041,N_11313);
and U12202 (N_12202,N_11380,N_11056);
nor U12203 (N_12203,N_11702,N_11011);
or U12204 (N_12204,N_11795,N_11431);
xor U12205 (N_12205,N_11914,N_11217);
nor U12206 (N_12206,N_11593,N_11300);
and U12207 (N_12207,N_11349,N_11672);
or U12208 (N_12208,N_11704,N_11995);
or U12209 (N_12209,N_11178,N_11289);
nand U12210 (N_12210,N_11455,N_11040);
nor U12211 (N_12211,N_11477,N_11093);
and U12212 (N_12212,N_11147,N_11925);
or U12213 (N_12213,N_11650,N_11543);
or U12214 (N_12214,N_11644,N_11442);
and U12215 (N_12215,N_11457,N_11548);
nor U12216 (N_12216,N_11356,N_11796);
nand U12217 (N_12217,N_11158,N_11318);
nor U12218 (N_12218,N_11322,N_11653);
nor U12219 (N_12219,N_11675,N_11857);
and U12220 (N_12220,N_11213,N_11784);
and U12221 (N_12221,N_11965,N_11463);
and U12222 (N_12222,N_11342,N_11798);
or U12223 (N_12223,N_11832,N_11646);
and U12224 (N_12224,N_11102,N_11231);
and U12225 (N_12225,N_11167,N_11782);
nand U12226 (N_12226,N_11727,N_11936);
and U12227 (N_12227,N_11331,N_11761);
nand U12228 (N_12228,N_11023,N_11334);
and U12229 (N_12229,N_11065,N_11825);
or U12230 (N_12230,N_11721,N_11716);
nand U12231 (N_12231,N_11366,N_11578);
and U12232 (N_12232,N_11000,N_11510);
and U12233 (N_12233,N_11392,N_11402);
nand U12234 (N_12234,N_11220,N_11597);
and U12235 (N_12235,N_11872,N_11888);
nand U12236 (N_12236,N_11758,N_11453);
and U12237 (N_12237,N_11964,N_11297);
or U12238 (N_12238,N_11101,N_11826);
xnor U12239 (N_12239,N_11903,N_11421);
nor U12240 (N_12240,N_11924,N_11467);
and U12241 (N_12241,N_11049,N_11892);
xnor U12242 (N_12242,N_11933,N_11242);
and U12243 (N_12243,N_11765,N_11272);
nand U12244 (N_12244,N_11608,N_11950);
nand U12245 (N_12245,N_11146,N_11454);
nand U12246 (N_12246,N_11233,N_11456);
nand U12247 (N_12247,N_11187,N_11847);
nand U12248 (N_12248,N_11541,N_11255);
nor U12249 (N_12249,N_11410,N_11172);
nor U12250 (N_12250,N_11620,N_11547);
nor U12251 (N_12251,N_11293,N_11573);
xor U12252 (N_12252,N_11630,N_11978);
xnor U12253 (N_12253,N_11916,N_11173);
and U12254 (N_12254,N_11232,N_11019);
or U12255 (N_12255,N_11698,N_11127);
and U12256 (N_12256,N_11057,N_11926);
and U12257 (N_12257,N_11487,N_11486);
nor U12258 (N_12258,N_11196,N_11111);
or U12259 (N_12259,N_11862,N_11495);
nor U12260 (N_12260,N_11214,N_11193);
nand U12261 (N_12261,N_11705,N_11182);
nor U12262 (N_12262,N_11419,N_11481);
or U12263 (N_12263,N_11728,N_11426);
or U12264 (N_12264,N_11959,N_11866);
xor U12265 (N_12265,N_11841,N_11780);
and U12266 (N_12266,N_11309,N_11375);
nor U12267 (N_12267,N_11623,N_11468);
nand U12268 (N_12268,N_11496,N_11325);
and U12269 (N_12269,N_11353,N_11501);
and U12270 (N_12270,N_11461,N_11730);
or U12271 (N_12271,N_11428,N_11120);
nor U12272 (N_12272,N_11096,N_11625);
nor U12273 (N_12273,N_11465,N_11180);
or U12274 (N_12274,N_11777,N_11651);
xor U12275 (N_12275,N_11478,N_11071);
and U12276 (N_12276,N_11937,N_11762);
nor U12277 (N_12277,N_11073,N_11133);
nand U12278 (N_12278,N_11955,N_11710);
nor U12279 (N_12279,N_11922,N_11471);
xnor U12280 (N_12280,N_11017,N_11094);
xnor U12281 (N_12281,N_11343,N_11404);
or U12282 (N_12282,N_11215,N_11086);
xnor U12283 (N_12283,N_11881,N_11168);
and U12284 (N_12284,N_11250,N_11062);
nor U12285 (N_12285,N_11212,N_11624);
nand U12286 (N_12286,N_11947,N_11533);
nand U12287 (N_12287,N_11475,N_11954);
or U12288 (N_12288,N_11169,N_11229);
xnor U12289 (N_12289,N_11080,N_11882);
nor U12290 (N_12290,N_11854,N_11904);
nand U12291 (N_12291,N_11186,N_11718);
and U12292 (N_12292,N_11531,N_11484);
xnor U12293 (N_12293,N_11503,N_11189);
nand U12294 (N_12294,N_11667,N_11218);
nand U12295 (N_12295,N_11606,N_11576);
nor U12296 (N_12296,N_11472,N_11915);
xnor U12297 (N_12297,N_11539,N_11450);
xor U12298 (N_12298,N_11860,N_11149);
xnor U12299 (N_12299,N_11192,N_11755);
or U12300 (N_12300,N_11181,N_11823);
nand U12301 (N_12301,N_11263,N_11740);
xnor U12302 (N_12302,N_11677,N_11491);
xor U12303 (N_12303,N_11734,N_11963);
nand U12304 (N_12304,N_11205,N_11448);
xnor U12305 (N_12305,N_11824,N_11666);
nand U12306 (N_12306,N_11084,N_11103);
nand U12307 (N_12307,N_11489,N_11775);
nor U12308 (N_12308,N_11565,N_11816);
nand U12309 (N_12309,N_11125,N_11350);
nand U12310 (N_12310,N_11618,N_11395);
nor U12311 (N_12311,N_11766,N_11208);
or U12312 (N_12312,N_11923,N_11273);
xor U12313 (N_12313,N_11164,N_11686);
and U12314 (N_12314,N_11075,N_11970);
nor U12315 (N_12315,N_11107,N_11741);
and U12316 (N_12316,N_11940,N_11869);
or U12317 (N_12317,N_11195,N_11767);
and U12318 (N_12318,N_11494,N_11047);
xor U12319 (N_12319,N_11291,N_11818);
nand U12320 (N_12320,N_11026,N_11747);
and U12321 (N_12321,N_11121,N_11445);
and U12322 (N_12322,N_11382,N_11266);
and U12323 (N_12323,N_11529,N_11814);
xor U12324 (N_12324,N_11074,N_11157);
xnor U12325 (N_12325,N_11523,N_11674);
nor U12326 (N_12326,N_11948,N_11413);
xor U12327 (N_12327,N_11070,N_11396);
or U12328 (N_12328,N_11427,N_11174);
nand U12329 (N_12329,N_11434,N_11889);
xnor U12330 (N_12330,N_11551,N_11596);
or U12331 (N_12331,N_11060,N_11805);
nand U12332 (N_12332,N_11935,N_11525);
or U12333 (N_12333,N_11984,N_11282);
or U12334 (N_12334,N_11681,N_11227);
or U12335 (N_12335,N_11788,N_11943);
xor U12336 (N_12336,N_11294,N_11899);
or U12337 (N_12337,N_11190,N_11534);
or U12338 (N_12338,N_11549,N_11113);
or U12339 (N_12339,N_11687,N_11198);
nor U12340 (N_12340,N_11462,N_11042);
nand U12341 (N_12341,N_11365,N_11237);
xnor U12342 (N_12342,N_11616,N_11401);
nor U12343 (N_12343,N_11840,N_11785);
and U12344 (N_12344,N_11971,N_11932);
nand U12345 (N_12345,N_11018,N_11540);
or U12346 (N_12346,N_11249,N_11012);
and U12347 (N_12347,N_11407,N_11574);
nand U12348 (N_12348,N_11361,N_11976);
nand U12349 (N_12349,N_11123,N_11206);
xnor U12350 (N_12350,N_11760,N_11386);
and U12351 (N_12351,N_11302,N_11776);
nand U12352 (N_12352,N_11240,N_11787);
and U12353 (N_12353,N_11595,N_11931);
and U12354 (N_12354,N_11763,N_11709);
nor U12355 (N_12355,N_11141,N_11051);
or U12356 (N_12356,N_11942,N_11424);
xor U12357 (N_12357,N_11295,N_11511);
or U12358 (N_12358,N_11336,N_11055);
nor U12359 (N_12359,N_11636,N_11813);
or U12360 (N_12360,N_11546,N_11329);
xnor U12361 (N_12361,N_11451,N_11010);
nor U12362 (N_12362,N_11119,N_11140);
or U12363 (N_12363,N_11945,N_11974);
xnor U12364 (N_12364,N_11009,N_11112);
or U12365 (N_12365,N_11415,N_11988);
or U12366 (N_12366,N_11609,N_11354);
or U12367 (N_12367,N_11639,N_11115);
and U12368 (N_12368,N_11707,N_11459);
nor U12369 (N_12369,N_11379,N_11928);
and U12370 (N_12370,N_11661,N_11808);
nor U12371 (N_12371,N_11226,N_11967);
xor U12372 (N_12372,N_11199,N_11559);
xnor U12373 (N_12373,N_11979,N_11148);
nand U12374 (N_12374,N_11744,N_11046);
or U12375 (N_12375,N_11260,N_11902);
nor U12376 (N_12376,N_11536,N_11982);
xnor U12377 (N_12377,N_11868,N_11757);
xnor U12378 (N_12378,N_11137,N_11580);
or U12379 (N_12379,N_11082,N_11020);
nor U12380 (N_12380,N_11305,N_11078);
nor U12381 (N_12381,N_11517,N_11310);
xor U12382 (N_12382,N_11197,N_11344);
nor U12383 (N_12383,N_11516,N_11341);
xor U12384 (N_12384,N_11280,N_11568);
xor U12385 (N_12385,N_11992,N_11064);
xor U12386 (N_12386,N_11276,N_11770);
and U12387 (N_12387,N_11092,N_11587);
and U12388 (N_12388,N_11034,N_11474);
and U12389 (N_12389,N_11768,N_11422);
xor U12390 (N_12390,N_11771,N_11773);
and U12391 (N_12391,N_11236,N_11397);
nor U12392 (N_12392,N_11706,N_11544);
and U12393 (N_12393,N_11052,N_11142);
and U12394 (N_12394,N_11958,N_11602);
nor U12395 (N_12395,N_11542,N_11720);
xnor U12396 (N_12396,N_11288,N_11977);
nor U12397 (N_12397,N_11518,N_11842);
nand U12398 (N_12398,N_11389,N_11558);
xor U12399 (N_12399,N_11277,N_11713);
xor U12400 (N_12400,N_11748,N_11919);
or U12401 (N_12401,N_11128,N_11492);
or U12402 (N_12402,N_11439,N_11286);
or U12403 (N_12403,N_11690,N_11203);
or U12404 (N_12404,N_11248,N_11553);
or U12405 (N_12405,N_11711,N_11238);
nor U12406 (N_12406,N_11360,N_11682);
nor U12407 (N_12407,N_11647,N_11482);
or U12408 (N_12408,N_11626,N_11166);
nor U12409 (N_12409,N_11521,N_11685);
nor U12410 (N_12410,N_11855,N_11171);
and U12411 (N_12411,N_11815,N_11676);
nand U12412 (N_12412,N_11729,N_11552);
xor U12413 (N_12413,N_11449,N_11605);
xor U12414 (N_12414,N_11500,N_11566);
and U12415 (N_12415,N_11861,N_11036);
xnor U12416 (N_12416,N_11663,N_11634);
or U12417 (N_12417,N_11985,N_11561);
nor U12418 (N_12418,N_11008,N_11953);
nand U12419 (N_12419,N_11490,N_11160);
nor U12420 (N_12420,N_11298,N_11239);
nand U12421 (N_12421,N_11876,N_11987);
or U12422 (N_12422,N_11257,N_11337);
and U12423 (N_12423,N_11981,N_11907);
xor U12424 (N_12424,N_11507,N_11917);
nand U12425 (N_12425,N_11400,N_11271);
nand U12426 (N_12426,N_11001,N_11485);
and U12427 (N_12427,N_11739,N_11348);
or U12428 (N_12428,N_11004,N_11411);
nor U12429 (N_12429,N_11554,N_11367);
xnor U12430 (N_12430,N_11499,N_11126);
xnor U12431 (N_12431,N_11999,N_11085);
nand U12432 (N_12432,N_11878,N_11139);
nand U12433 (N_12433,N_11317,N_11403);
and U12434 (N_12434,N_11044,N_11921);
nand U12435 (N_12435,N_11683,N_11247);
nand U12436 (N_12436,N_11433,N_11384);
nor U12437 (N_12437,N_11590,N_11530);
or U12438 (N_12438,N_11138,N_11024);
nor U12439 (N_12439,N_11837,N_11786);
nor U12440 (N_12440,N_11591,N_11259);
and U12441 (N_12441,N_11284,N_11446);
nand U12442 (N_12442,N_11738,N_11556);
or U12443 (N_12443,N_11594,N_11037);
nor U12444 (N_12444,N_11946,N_11821);
xnor U12445 (N_12445,N_11598,N_11592);
or U12446 (N_12446,N_11612,N_11779);
xnor U12447 (N_12447,N_11691,N_11480);
and U12448 (N_12448,N_11893,N_11949);
nor U12449 (N_12449,N_11429,N_11301);
xnor U12450 (N_12450,N_11656,N_11887);
and U12451 (N_12451,N_11619,N_11340);
xnor U12452 (N_12452,N_11324,N_11108);
nor U12453 (N_12453,N_11520,N_11512);
or U12454 (N_12454,N_11005,N_11378);
nand U12455 (N_12455,N_11524,N_11252);
nand U12456 (N_12456,N_11209,N_11308);
nand U12457 (N_12457,N_11831,N_11731);
xor U12458 (N_12458,N_11416,N_11437);
xor U12459 (N_12459,N_11628,N_11519);
or U12460 (N_12460,N_11076,N_11772);
nor U12461 (N_12461,N_11175,N_11603);
nor U12462 (N_12462,N_11649,N_11989);
nand U12463 (N_12463,N_11607,N_11745);
nor U12464 (N_12464,N_11357,N_11145);
and U12465 (N_12465,N_11314,N_11464);
xor U12466 (N_12466,N_11843,N_11253);
and U12467 (N_12467,N_11673,N_11007);
nand U12468 (N_12468,N_11221,N_11479);
and U12469 (N_12469,N_11746,N_11335);
or U12470 (N_12470,N_11708,N_11697);
nand U12471 (N_12471,N_11752,N_11154);
nor U12472 (N_12472,N_11885,N_11436);
and U12473 (N_12473,N_11162,N_11582);
nand U12474 (N_12474,N_11029,N_11290);
and U12475 (N_12475,N_11323,N_11759);
and U12476 (N_12476,N_11629,N_11054);
nor U12477 (N_12477,N_11764,N_11118);
xor U12478 (N_12478,N_11204,N_11050);
nand U12479 (N_12479,N_11114,N_11090);
xnor U12480 (N_12480,N_11927,N_11905);
or U12481 (N_12481,N_11035,N_11116);
nand U12482 (N_12482,N_11703,N_11371);
nand U12483 (N_12483,N_11264,N_11527);
nand U12484 (N_12484,N_11600,N_11105);
and U12485 (N_12485,N_11791,N_11032);
and U12486 (N_12486,N_11660,N_11664);
and U12487 (N_12487,N_11068,N_11792);
and U12488 (N_12488,N_11613,N_11934);
xor U12489 (N_12489,N_11846,N_11884);
nand U12490 (N_12490,N_11622,N_11920);
xnor U12491 (N_12491,N_11216,N_11014);
xnor U12492 (N_12492,N_11045,N_11637);
and U12493 (N_12493,N_11994,N_11850);
and U12494 (N_12494,N_11712,N_11201);
xor U12495 (N_12495,N_11006,N_11043);
and U12496 (N_12496,N_11635,N_11679);
xnor U12497 (N_12497,N_11473,N_11621);
nor U12498 (N_12498,N_11370,N_11993);
or U12499 (N_12499,N_11652,N_11333);
and U12500 (N_12500,N_11724,N_11070);
or U12501 (N_12501,N_11385,N_11721);
and U12502 (N_12502,N_11292,N_11662);
nor U12503 (N_12503,N_11843,N_11662);
or U12504 (N_12504,N_11567,N_11202);
xnor U12505 (N_12505,N_11272,N_11857);
nor U12506 (N_12506,N_11086,N_11057);
nor U12507 (N_12507,N_11723,N_11013);
nand U12508 (N_12508,N_11185,N_11003);
nor U12509 (N_12509,N_11786,N_11098);
or U12510 (N_12510,N_11448,N_11660);
or U12511 (N_12511,N_11690,N_11067);
or U12512 (N_12512,N_11514,N_11250);
nor U12513 (N_12513,N_11390,N_11955);
nor U12514 (N_12514,N_11044,N_11432);
or U12515 (N_12515,N_11079,N_11689);
xnor U12516 (N_12516,N_11906,N_11218);
nand U12517 (N_12517,N_11047,N_11376);
nor U12518 (N_12518,N_11408,N_11372);
or U12519 (N_12519,N_11468,N_11950);
nand U12520 (N_12520,N_11603,N_11413);
nor U12521 (N_12521,N_11079,N_11453);
or U12522 (N_12522,N_11957,N_11673);
nor U12523 (N_12523,N_11975,N_11324);
nand U12524 (N_12524,N_11944,N_11229);
nor U12525 (N_12525,N_11214,N_11719);
nor U12526 (N_12526,N_11675,N_11874);
and U12527 (N_12527,N_11250,N_11776);
nand U12528 (N_12528,N_11069,N_11514);
or U12529 (N_12529,N_11768,N_11410);
and U12530 (N_12530,N_11292,N_11314);
and U12531 (N_12531,N_11773,N_11167);
nor U12532 (N_12532,N_11628,N_11612);
xor U12533 (N_12533,N_11670,N_11366);
or U12534 (N_12534,N_11925,N_11613);
and U12535 (N_12535,N_11991,N_11891);
nand U12536 (N_12536,N_11100,N_11072);
nor U12537 (N_12537,N_11334,N_11854);
nor U12538 (N_12538,N_11251,N_11629);
and U12539 (N_12539,N_11832,N_11032);
nor U12540 (N_12540,N_11907,N_11560);
nand U12541 (N_12541,N_11262,N_11422);
or U12542 (N_12542,N_11518,N_11522);
nor U12543 (N_12543,N_11404,N_11540);
or U12544 (N_12544,N_11634,N_11390);
nand U12545 (N_12545,N_11303,N_11863);
xnor U12546 (N_12546,N_11307,N_11473);
nor U12547 (N_12547,N_11166,N_11333);
xnor U12548 (N_12548,N_11425,N_11440);
xor U12549 (N_12549,N_11842,N_11035);
nand U12550 (N_12550,N_11372,N_11513);
nor U12551 (N_12551,N_11960,N_11168);
or U12552 (N_12552,N_11278,N_11435);
nand U12553 (N_12553,N_11825,N_11010);
nand U12554 (N_12554,N_11604,N_11314);
and U12555 (N_12555,N_11943,N_11830);
nor U12556 (N_12556,N_11242,N_11113);
or U12557 (N_12557,N_11221,N_11024);
xnor U12558 (N_12558,N_11862,N_11693);
nand U12559 (N_12559,N_11570,N_11213);
xnor U12560 (N_12560,N_11105,N_11274);
nand U12561 (N_12561,N_11225,N_11042);
nor U12562 (N_12562,N_11678,N_11331);
xnor U12563 (N_12563,N_11174,N_11956);
xnor U12564 (N_12564,N_11417,N_11534);
or U12565 (N_12565,N_11228,N_11396);
and U12566 (N_12566,N_11706,N_11273);
and U12567 (N_12567,N_11132,N_11351);
nor U12568 (N_12568,N_11140,N_11643);
nand U12569 (N_12569,N_11370,N_11499);
nor U12570 (N_12570,N_11169,N_11881);
xnor U12571 (N_12571,N_11405,N_11541);
or U12572 (N_12572,N_11037,N_11185);
xnor U12573 (N_12573,N_11419,N_11296);
and U12574 (N_12574,N_11822,N_11309);
or U12575 (N_12575,N_11252,N_11169);
nand U12576 (N_12576,N_11720,N_11255);
nor U12577 (N_12577,N_11929,N_11111);
or U12578 (N_12578,N_11343,N_11930);
nor U12579 (N_12579,N_11529,N_11460);
nor U12580 (N_12580,N_11192,N_11206);
nor U12581 (N_12581,N_11565,N_11365);
or U12582 (N_12582,N_11264,N_11721);
xor U12583 (N_12583,N_11268,N_11049);
or U12584 (N_12584,N_11063,N_11716);
xnor U12585 (N_12585,N_11755,N_11131);
or U12586 (N_12586,N_11952,N_11384);
nor U12587 (N_12587,N_11410,N_11464);
nand U12588 (N_12588,N_11829,N_11201);
nand U12589 (N_12589,N_11400,N_11059);
and U12590 (N_12590,N_11969,N_11120);
xnor U12591 (N_12591,N_11354,N_11758);
nor U12592 (N_12592,N_11062,N_11375);
xor U12593 (N_12593,N_11743,N_11695);
and U12594 (N_12594,N_11342,N_11579);
and U12595 (N_12595,N_11513,N_11936);
xor U12596 (N_12596,N_11319,N_11600);
and U12597 (N_12597,N_11434,N_11887);
nor U12598 (N_12598,N_11935,N_11069);
nor U12599 (N_12599,N_11627,N_11866);
nand U12600 (N_12600,N_11936,N_11890);
or U12601 (N_12601,N_11173,N_11330);
nor U12602 (N_12602,N_11839,N_11368);
nand U12603 (N_12603,N_11580,N_11869);
nor U12604 (N_12604,N_11231,N_11052);
xor U12605 (N_12605,N_11244,N_11842);
or U12606 (N_12606,N_11550,N_11970);
xnor U12607 (N_12607,N_11346,N_11534);
nand U12608 (N_12608,N_11628,N_11212);
and U12609 (N_12609,N_11054,N_11591);
nand U12610 (N_12610,N_11255,N_11635);
xnor U12611 (N_12611,N_11560,N_11982);
nand U12612 (N_12612,N_11424,N_11884);
or U12613 (N_12613,N_11360,N_11328);
nand U12614 (N_12614,N_11201,N_11747);
and U12615 (N_12615,N_11894,N_11324);
xor U12616 (N_12616,N_11407,N_11265);
nor U12617 (N_12617,N_11437,N_11940);
and U12618 (N_12618,N_11714,N_11119);
and U12619 (N_12619,N_11931,N_11002);
nand U12620 (N_12620,N_11969,N_11156);
and U12621 (N_12621,N_11917,N_11156);
and U12622 (N_12622,N_11022,N_11403);
or U12623 (N_12623,N_11216,N_11078);
or U12624 (N_12624,N_11804,N_11658);
xor U12625 (N_12625,N_11056,N_11876);
nand U12626 (N_12626,N_11912,N_11224);
and U12627 (N_12627,N_11597,N_11321);
nand U12628 (N_12628,N_11530,N_11339);
or U12629 (N_12629,N_11083,N_11753);
nand U12630 (N_12630,N_11724,N_11762);
nor U12631 (N_12631,N_11861,N_11695);
xor U12632 (N_12632,N_11645,N_11891);
xnor U12633 (N_12633,N_11285,N_11855);
nor U12634 (N_12634,N_11113,N_11460);
nand U12635 (N_12635,N_11359,N_11864);
xnor U12636 (N_12636,N_11139,N_11563);
or U12637 (N_12637,N_11040,N_11112);
nor U12638 (N_12638,N_11654,N_11396);
nand U12639 (N_12639,N_11399,N_11269);
and U12640 (N_12640,N_11644,N_11335);
nand U12641 (N_12641,N_11388,N_11705);
xnor U12642 (N_12642,N_11756,N_11650);
xnor U12643 (N_12643,N_11937,N_11010);
or U12644 (N_12644,N_11291,N_11334);
and U12645 (N_12645,N_11299,N_11755);
or U12646 (N_12646,N_11159,N_11148);
xnor U12647 (N_12647,N_11337,N_11204);
and U12648 (N_12648,N_11963,N_11812);
or U12649 (N_12649,N_11488,N_11844);
and U12650 (N_12650,N_11624,N_11593);
nand U12651 (N_12651,N_11989,N_11950);
or U12652 (N_12652,N_11881,N_11182);
nand U12653 (N_12653,N_11073,N_11419);
nand U12654 (N_12654,N_11720,N_11595);
nand U12655 (N_12655,N_11757,N_11750);
nand U12656 (N_12656,N_11746,N_11392);
and U12657 (N_12657,N_11219,N_11999);
and U12658 (N_12658,N_11210,N_11694);
nand U12659 (N_12659,N_11383,N_11050);
xnor U12660 (N_12660,N_11863,N_11376);
and U12661 (N_12661,N_11256,N_11363);
nand U12662 (N_12662,N_11392,N_11730);
nand U12663 (N_12663,N_11203,N_11211);
nor U12664 (N_12664,N_11620,N_11831);
or U12665 (N_12665,N_11290,N_11088);
or U12666 (N_12666,N_11363,N_11911);
nor U12667 (N_12667,N_11783,N_11242);
xor U12668 (N_12668,N_11590,N_11797);
nand U12669 (N_12669,N_11559,N_11013);
or U12670 (N_12670,N_11892,N_11777);
nor U12671 (N_12671,N_11792,N_11800);
xnor U12672 (N_12672,N_11378,N_11347);
nor U12673 (N_12673,N_11725,N_11545);
xnor U12674 (N_12674,N_11054,N_11424);
nand U12675 (N_12675,N_11951,N_11517);
xnor U12676 (N_12676,N_11654,N_11944);
and U12677 (N_12677,N_11984,N_11884);
or U12678 (N_12678,N_11155,N_11502);
or U12679 (N_12679,N_11360,N_11934);
nand U12680 (N_12680,N_11177,N_11959);
nor U12681 (N_12681,N_11816,N_11680);
and U12682 (N_12682,N_11502,N_11481);
nand U12683 (N_12683,N_11754,N_11581);
and U12684 (N_12684,N_11395,N_11621);
nor U12685 (N_12685,N_11066,N_11466);
nand U12686 (N_12686,N_11123,N_11921);
nor U12687 (N_12687,N_11757,N_11001);
and U12688 (N_12688,N_11515,N_11411);
and U12689 (N_12689,N_11137,N_11437);
and U12690 (N_12690,N_11578,N_11184);
xor U12691 (N_12691,N_11115,N_11084);
nand U12692 (N_12692,N_11632,N_11972);
and U12693 (N_12693,N_11155,N_11617);
xnor U12694 (N_12694,N_11519,N_11052);
or U12695 (N_12695,N_11705,N_11526);
or U12696 (N_12696,N_11839,N_11918);
nand U12697 (N_12697,N_11702,N_11963);
xor U12698 (N_12698,N_11824,N_11538);
or U12699 (N_12699,N_11184,N_11969);
nor U12700 (N_12700,N_11983,N_11981);
and U12701 (N_12701,N_11402,N_11332);
or U12702 (N_12702,N_11295,N_11348);
or U12703 (N_12703,N_11427,N_11249);
nand U12704 (N_12704,N_11448,N_11973);
nand U12705 (N_12705,N_11263,N_11451);
xor U12706 (N_12706,N_11621,N_11141);
xor U12707 (N_12707,N_11747,N_11208);
nand U12708 (N_12708,N_11703,N_11174);
nand U12709 (N_12709,N_11392,N_11779);
xnor U12710 (N_12710,N_11497,N_11791);
and U12711 (N_12711,N_11763,N_11380);
nor U12712 (N_12712,N_11005,N_11504);
nor U12713 (N_12713,N_11846,N_11473);
nand U12714 (N_12714,N_11889,N_11065);
and U12715 (N_12715,N_11723,N_11539);
nand U12716 (N_12716,N_11336,N_11881);
or U12717 (N_12717,N_11940,N_11561);
and U12718 (N_12718,N_11011,N_11198);
nor U12719 (N_12719,N_11644,N_11163);
or U12720 (N_12720,N_11171,N_11994);
nand U12721 (N_12721,N_11172,N_11632);
xnor U12722 (N_12722,N_11209,N_11362);
or U12723 (N_12723,N_11474,N_11308);
or U12724 (N_12724,N_11424,N_11604);
nand U12725 (N_12725,N_11283,N_11707);
nor U12726 (N_12726,N_11817,N_11045);
nand U12727 (N_12727,N_11833,N_11441);
nand U12728 (N_12728,N_11244,N_11372);
nand U12729 (N_12729,N_11745,N_11305);
xnor U12730 (N_12730,N_11379,N_11397);
and U12731 (N_12731,N_11559,N_11879);
or U12732 (N_12732,N_11595,N_11118);
xor U12733 (N_12733,N_11666,N_11854);
nor U12734 (N_12734,N_11847,N_11780);
and U12735 (N_12735,N_11056,N_11425);
or U12736 (N_12736,N_11094,N_11723);
nand U12737 (N_12737,N_11724,N_11845);
nor U12738 (N_12738,N_11849,N_11787);
xor U12739 (N_12739,N_11080,N_11754);
nand U12740 (N_12740,N_11389,N_11044);
nor U12741 (N_12741,N_11527,N_11011);
or U12742 (N_12742,N_11103,N_11453);
xor U12743 (N_12743,N_11510,N_11515);
nand U12744 (N_12744,N_11832,N_11315);
and U12745 (N_12745,N_11879,N_11944);
nand U12746 (N_12746,N_11343,N_11797);
and U12747 (N_12747,N_11037,N_11274);
nor U12748 (N_12748,N_11510,N_11201);
nand U12749 (N_12749,N_11113,N_11689);
or U12750 (N_12750,N_11444,N_11249);
or U12751 (N_12751,N_11704,N_11792);
or U12752 (N_12752,N_11400,N_11810);
and U12753 (N_12753,N_11604,N_11563);
nor U12754 (N_12754,N_11341,N_11861);
xnor U12755 (N_12755,N_11101,N_11815);
xnor U12756 (N_12756,N_11482,N_11619);
nand U12757 (N_12757,N_11291,N_11270);
xor U12758 (N_12758,N_11835,N_11222);
and U12759 (N_12759,N_11697,N_11815);
or U12760 (N_12760,N_11152,N_11035);
and U12761 (N_12761,N_11402,N_11139);
nor U12762 (N_12762,N_11805,N_11849);
nor U12763 (N_12763,N_11958,N_11727);
or U12764 (N_12764,N_11318,N_11960);
nand U12765 (N_12765,N_11395,N_11786);
xnor U12766 (N_12766,N_11221,N_11351);
nor U12767 (N_12767,N_11031,N_11898);
nor U12768 (N_12768,N_11398,N_11475);
xor U12769 (N_12769,N_11431,N_11383);
nand U12770 (N_12770,N_11523,N_11347);
nand U12771 (N_12771,N_11664,N_11363);
nor U12772 (N_12772,N_11326,N_11696);
or U12773 (N_12773,N_11714,N_11225);
nand U12774 (N_12774,N_11243,N_11945);
or U12775 (N_12775,N_11693,N_11739);
and U12776 (N_12776,N_11866,N_11569);
nand U12777 (N_12777,N_11537,N_11248);
and U12778 (N_12778,N_11617,N_11549);
xor U12779 (N_12779,N_11719,N_11317);
xor U12780 (N_12780,N_11020,N_11378);
or U12781 (N_12781,N_11634,N_11132);
or U12782 (N_12782,N_11332,N_11898);
xor U12783 (N_12783,N_11380,N_11083);
nor U12784 (N_12784,N_11451,N_11093);
and U12785 (N_12785,N_11634,N_11838);
nor U12786 (N_12786,N_11171,N_11073);
or U12787 (N_12787,N_11795,N_11962);
nand U12788 (N_12788,N_11912,N_11577);
or U12789 (N_12789,N_11032,N_11252);
or U12790 (N_12790,N_11110,N_11645);
nand U12791 (N_12791,N_11221,N_11517);
nor U12792 (N_12792,N_11518,N_11389);
nand U12793 (N_12793,N_11572,N_11439);
or U12794 (N_12794,N_11666,N_11503);
xnor U12795 (N_12795,N_11856,N_11848);
nand U12796 (N_12796,N_11513,N_11208);
or U12797 (N_12797,N_11994,N_11639);
xor U12798 (N_12798,N_11456,N_11380);
nand U12799 (N_12799,N_11613,N_11025);
or U12800 (N_12800,N_11433,N_11137);
nand U12801 (N_12801,N_11283,N_11067);
nand U12802 (N_12802,N_11525,N_11056);
nor U12803 (N_12803,N_11899,N_11139);
xor U12804 (N_12804,N_11786,N_11856);
nand U12805 (N_12805,N_11564,N_11875);
nand U12806 (N_12806,N_11600,N_11516);
nor U12807 (N_12807,N_11047,N_11222);
nand U12808 (N_12808,N_11772,N_11715);
nor U12809 (N_12809,N_11116,N_11973);
and U12810 (N_12810,N_11346,N_11668);
or U12811 (N_12811,N_11580,N_11491);
xnor U12812 (N_12812,N_11071,N_11179);
nand U12813 (N_12813,N_11880,N_11722);
nor U12814 (N_12814,N_11458,N_11561);
nand U12815 (N_12815,N_11448,N_11422);
and U12816 (N_12816,N_11139,N_11429);
nand U12817 (N_12817,N_11924,N_11480);
or U12818 (N_12818,N_11388,N_11148);
nor U12819 (N_12819,N_11897,N_11650);
nand U12820 (N_12820,N_11105,N_11607);
xor U12821 (N_12821,N_11822,N_11623);
xor U12822 (N_12822,N_11315,N_11622);
nor U12823 (N_12823,N_11256,N_11317);
or U12824 (N_12824,N_11273,N_11365);
xor U12825 (N_12825,N_11073,N_11622);
xnor U12826 (N_12826,N_11701,N_11211);
nand U12827 (N_12827,N_11735,N_11755);
or U12828 (N_12828,N_11733,N_11179);
or U12829 (N_12829,N_11395,N_11753);
or U12830 (N_12830,N_11404,N_11976);
nor U12831 (N_12831,N_11193,N_11195);
xnor U12832 (N_12832,N_11893,N_11003);
or U12833 (N_12833,N_11898,N_11918);
nor U12834 (N_12834,N_11751,N_11832);
or U12835 (N_12835,N_11478,N_11504);
and U12836 (N_12836,N_11385,N_11928);
nor U12837 (N_12837,N_11074,N_11695);
nand U12838 (N_12838,N_11653,N_11011);
nand U12839 (N_12839,N_11452,N_11555);
nand U12840 (N_12840,N_11354,N_11613);
nand U12841 (N_12841,N_11167,N_11566);
nor U12842 (N_12842,N_11290,N_11441);
nand U12843 (N_12843,N_11910,N_11252);
nand U12844 (N_12844,N_11857,N_11107);
or U12845 (N_12845,N_11379,N_11365);
xor U12846 (N_12846,N_11453,N_11093);
or U12847 (N_12847,N_11441,N_11621);
and U12848 (N_12848,N_11346,N_11607);
and U12849 (N_12849,N_11874,N_11681);
nand U12850 (N_12850,N_11902,N_11818);
nor U12851 (N_12851,N_11228,N_11049);
or U12852 (N_12852,N_11651,N_11773);
and U12853 (N_12853,N_11492,N_11039);
nor U12854 (N_12854,N_11447,N_11639);
and U12855 (N_12855,N_11135,N_11451);
or U12856 (N_12856,N_11856,N_11799);
xor U12857 (N_12857,N_11698,N_11145);
and U12858 (N_12858,N_11966,N_11870);
and U12859 (N_12859,N_11806,N_11339);
nor U12860 (N_12860,N_11365,N_11282);
and U12861 (N_12861,N_11703,N_11787);
xor U12862 (N_12862,N_11964,N_11270);
or U12863 (N_12863,N_11236,N_11823);
xnor U12864 (N_12864,N_11075,N_11334);
nor U12865 (N_12865,N_11544,N_11125);
nand U12866 (N_12866,N_11533,N_11367);
or U12867 (N_12867,N_11891,N_11667);
or U12868 (N_12868,N_11458,N_11385);
and U12869 (N_12869,N_11437,N_11765);
nor U12870 (N_12870,N_11319,N_11947);
or U12871 (N_12871,N_11016,N_11264);
nor U12872 (N_12872,N_11137,N_11728);
nor U12873 (N_12873,N_11831,N_11638);
or U12874 (N_12874,N_11621,N_11711);
nand U12875 (N_12875,N_11218,N_11774);
nor U12876 (N_12876,N_11864,N_11879);
xor U12877 (N_12877,N_11812,N_11150);
nor U12878 (N_12878,N_11660,N_11437);
nand U12879 (N_12879,N_11904,N_11267);
or U12880 (N_12880,N_11756,N_11424);
and U12881 (N_12881,N_11665,N_11512);
nand U12882 (N_12882,N_11795,N_11422);
nor U12883 (N_12883,N_11453,N_11712);
xnor U12884 (N_12884,N_11608,N_11031);
nand U12885 (N_12885,N_11664,N_11701);
and U12886 (N_12886,N_11476,N_11924);
or U12887 (N_12887,N_11931,N_11757);
and U12888 (N_12888,N_11854,N_11036);
nand U12889 (N_12889,N_11671,N_11913);
xor U12890 (N_12890,N_11778,N_11743);
nor U12891 (N_12891,N_11151,N_11238);
and U12892 (N_12892,N_11503,N_11054);
and U12893 (N_12893,N_11560,N_11208);
xnor U12894 (N_12894,N_11434,N_11358);
or U12895 (N_12895,N_11988,N_11222);
nor U12896 (N_12896,N_11735,N_11723);
or U12897 (N_12897,N_11609,N_11046);
nand U12898 (N_12898,N_11286,N_11129);
or U12899 (N_12899,N_11340,N_11465);
xor U12900 (N_12900,N_11744,N_11355);
xnor U12901 (N_12901,N_11025,N_11882);
nand U12902 (N_12902,N_11888,N_11638);
xnor U12903 (N_12903,N_11252,N_11605);
and U12904 (N_12904,N_11019,N_11955);
nand U12905 (N_12905,N_11914,N_11497);
or U12906 (N_12906,N_11213,N_11781);
and U12907 (N_12907,N_11925,N_11094);
and U12908 (N_12908,N_11572,N_11222);
nor U12909 (N_12909,N_11162,N_11876);
nand U12910 (N_12910,N_11667,N_11402);
nand U12911 (N_12911,N_11029,N_11469);
and U12912 (N_12912,N_11008,N_11097);
or U12913 (N_12913,N_11674,N_11468);
and U12914 (N_12914,N_11237,N_11651);
or U12915 (N_12915,N_11714,N_11287);
and U12916 (N_12916,N_11142,N_11731);
nor U12917 (N_12917,N_11947,N_11353);
nor U12918 (N_12918,N_11878,N_11874);
nor U12919 (N_12919,N_11669,N_11113);
xnor U12920 (N_12920,N_11415,N_11280);
nor U12921 (N_12921,N_11019,N_11853);
and U12922 (N_12922,N_11255,N_11908);
nand U12923 (N_12923,N_11781,N_11116);
or U12924 (N_12924,N_11901,N_11880);
nand U12925 (N_12925,N_11216,N_11542);
or U12926 (N_12926,N_11477,N_11266);
and U12927 (N_12927,N_11268,N_11244);
xor U12928 (N_12928,N_11154,N_11050);
xnor U12929 (N_12929,N_11702,N_11978);
or U12930 (N_12930,N_11131,N_11624);
nand U12931 (N_12931,N_11252,N_11904);
xor U12932 (N_12932,N_11368,N_11708);
nand U12933 (N_12933,N_11171,N_11776);
nand U12934 (N_12934,N_11110,N_11304);
xnor U12935 (N_12935,N_11305,N_11777);
nand U12936 (N_12936,N_11590,N_11071);
or U12937 (N_12937,N_11779,N_11859);
xor U12938 (N_12938,N_11742,N_11629);
or U12939 (N_12939,N_11470,N_11331);
or U12940 (N_12940,N_11058,N_11648);
xor U12941 (N_12941,N_11154,N_11375);
nand U12942 (N_12942,N_11982,N_11948);
xor U12943 (N_12943,N_11297,N_11111);
nand U12944 (N_12944,N_11757,N_11771);
nand U12945 (N_12945,N_11721,N_11713);
nor U12946 (N_12946,N_11933,N_11031);
or U12947 (N_12947,N_11731,N_11480);
and U12948 (N_12948,N_11101,N_11788);
or U12949 (N_12949,N_11327,N_11849);
nor U12950 (N_12950,N_11302,N_11167);
nand U12951 (N_12951,N_11533,N_11096);
nor U12952 (N_12952,N_11181,N_11328);
nand U12953 (N_12953,N_11096,N_11364);
nor U12954 (N_12954,N_11367,N_11543);
xnor U12955 (N_12955,N_11690,N_11844);
nand U12956 (N_12956,N_11968,N_11239);
or U12957 (N_12957,N_11275,N_11215);
xor U12958 (N_12958,N_11081,N_11404);
nand U12959 (N_12959,N_11110,N_11345);
and U12960 (N_12960,N_11105,N_11116);
and U12961 (N_12961,N_11145,N_11294);
xnor U12962 (N_12962,N_11514,N_11570);
nor U12963 (N_12963,N_11707,N_11277);
nand U12964 (N_12964,N_11718,N_11455);
nor U12965 (N_12965,N_11257,N_11250);
and U12966 (N_12966,N_11215,N_11411);
and U12967 (N_12967,N_11122,N_11924);
or U12968 (N_12968,N_11883,N_11754);
nand U12969 (N_12969,N_11861,N_11972);
and U12970 (N_12970,N_11237,N_11131);
xor U12971 (N_12971,N_11563,N_11660);
or U12972 (N_12972,N_11671,N_11239);
nor U12973 (N_12973,N_11491,N_11409);
nand U12974 (N_12974,N_11602,N_11456);
nor U12975 (N_12975,N_11949,N_11640);
and U12976 (N_12976,N_11736,N_11957);
xnor U12977 (N_12977,N_11368,N_11710);
xnor U12978 (N_12978,N_11671,N_11311);
and U12979 (N_12979,N_11610,N_11964);
and U12980 (N_12980,N_11136,N_11163);
and U12981 (N_12981,N_11196,N_11698);
and U12982 (N_12982,N_11702,N_11472);
and U12983 (N_12983,N_11849,N_11519);
nand U12984 (N_12984,N_11810,N_11854);
and U12985 (N_12985,N_11227,N_11392);
nand U12986 (N_12986,N_11643,N_11587);
and U12987 (N_12987,N_11026,N_11437);
nor U12988 (N_12988,N_11777,N_11555);
nand U12989 (N_12989,N_11959,N_11472);
nor U12990 (N_12990,N_11369,N_11440);
nor U12991 (N_12991,N_11901,N_11182);
nor U12992 (N_12992,N_11676,N_11423);
and U12993 (N_12993,N_11959,N_11794);
xnor U12994 (N_12994,N_11711,N_11261);
and U12995 (N_12995,N_11240,N_11007);
and U12996 (N_12996,N_11170,N_11507);
nand U12997 (N_12997,N_11668,N_11107);
nand U12998 (N_12998,N_11984,N_11442);
and U12999 (N_12999,N_11353,N_11551);
nor U13000 (N_13000,N_12784,N_12065);
or U13001 (N_13001,N_12719,N_12907);
nand U13002 (N_13002,N_12400,N_12139);
or U13003 (N_13003,N_12180,N_12676);
nor U13004 (N_13004,N_12957,N_12373);
nor U13005 (N_13005,N_12260,N_12145);
xnor U13006 (N_13006,N_12130,N_12293);
or U13007 (N_13007,N_12518,N_12868);
or U13008 (N_13008,N_12574,N_12126);
nor U13009 (N_13009,N_12999,N_12779);
nand U13010 (N_13010,N_12242,N_12668);
and U13011 (N_13011,N_12950,N_12646);
nand U13012 (N_13012,N_12214,N_12072);
nand U13013 (N_13013,N_12577,N_12044);
or U13014 (N_13014,N_12187,N_12621);
nor U13015 (N_13015,N_12171,N_12054);
xor U13016 (N_13016,N_12360,N_12745);
and U13017 (N_13017,N_12380,N_12462);
nand U13018 (N_13018,N_12367,N_12693);
nand U13019 (N_13019,N_12204,N_12250);
nor U13020 (N_13020,N_12697,N_12437);
nor U13021 (N_13021,N_12424,N_12759);
or U13022 (N_13022,N_12528,N_12468);
nand U13023 (N_13023,N_12743,N_12164);
or U13024 (N_13024,N_12057,N_12262);
nor U13025 (N_13025,N_12484,N_12202);
nand U13026 (N_13026,N_12850,N_12459);
nand U13027 (N_13027,N_12622,N_12964);
xor U13028 (N_13028,N_12182,N_12946);
and U13029 (N_13029,N_12474,N_12819);
nand U13030 (N_13030,N_12525,N_12822);
nor U13031 (N_13031,N_12485,N_12448);
xnor U13032 (N_13032,N_12547,N_12857);
or U13033 (N_13033,N_12770,N_12690);
and U13034 (N_13034,N_12852,N_12123);
nor U13035 (N_13035,N_12099,N_12159);
nand U13036 (N_13036,N_12633,N_12737);
xnor U13037 (N_13037,N_12575,N_12364);
and U13038 (N_13038,N_12684,N_12884);
nand U13039 (N_13039,N_12751,N_12592);
nor U13040 (N_13040,N_12681,N_12166);
nand U13041 (N_13041,N_12301,N_12457);
xnor U13042 (N_13042,N_12285,N_12168);
nand U13043 (N_13043,N_12553,N_12025);
or U13044 (N_13044,N_12066,N_12625);
xor U13045 (N_13045,N_12004,N_12512);
nand U13046 (N_13046,N_12791,N_12515);
nor U13047 (N_13047,N_12392,N_12692);
xor U13048 (N_13048,N_12943,N_12877);
xnor U13049 (N_13049,N_12189,N_12607);
or U13050 (N_13050,N_12090,N_12605);
and U13051 (N_13051,N_12479,N_12221);
nor U13052 (N_13052,N_12270,N_12100);
nand U13053 (N_13053,N_12982,N_12344);
or U13054 (N_13054,N_12069,N_12033);
xnor U13055 (N_13055,N_12273,N_12452);
and U13056 (N_13056,N_12427,N_12703);
nor U13057 (N_13057,N_12489,N_12073);
nand U13058 (N_13058,N_12629,N_12352);
nor U13059 (N_13059,N_12193,N_12058);
nand U13060 (N_13060,N_12312,N_12430);
or U13061 (N_13061,N_12695,N_12807);
or U13062 (N_13062,N_12562,N_12021);
nor U13063 (N_13063,N_12175,N_12153);
and U13064 (N_13064,N_12141,N_12418);
and U13065 (N_13065,N_12490,N_12009);
nor U13066 (N_13066,N_12840,N_12998);
nor U13067 (N_13067,N_12778,N_12029);
nor U13068 (N_13068,N_12304,N_12048);
nand U13069 (N_13069,N_12002,N_12776);
or U13070 (N_13070,N_12238,N_12319);
and U13071 (N_13071,N_12989,N_12197);
and U13072 (N_13072,N_12353,N_12632);
nand U13073 (N_13073,N_12675,N_12067);
xnor U13074 (N_13074,N_12519,N_12712);
nor U13075 (N_13075,N_12649,N_12348);
nand U13076 (N_13076,N_12031,N_12381);
and U13077 (N_13077,N_12915,N_12134);
nor U13078 (N_13078,N_12597,N_12912);
xnor U13079 (N_13079,N_12713,N_12920);
or U13080 (N_13080,N_12150,N_12074);
or U13081 (N_13081,N_12570,N_12094);
nor U13082 (N_13082,N_12885,N_12615);
or U13083 (N_13083,N_12325,N_12390);
and U13084 (N_13084,N_12120,N_12599);
or U13085 (N_13085,N_12201,N_12787);
xnor U13086 (N_13086,N_12942,N_12103);
and U13087 (N_13087,N_12742,N_12538);
nor U13088 (N_13088,N_12642,N_12389);
nand U13089 (N_13089,N_12661,N_12112);
xor U13090 (N_13090,N_12415,N_12209);
xor U13091 (N_13091,N_12556,N_12508);
xnor U13092 (N_13092,N_12612,N_12454);
nor U13093 (N_13093,N_12289,N_12053);
or U13094 (N_13094,N_12035,N_12410);
nand U13095 (N_13095,N_12143,N_12817);
nand U13096 (N_13096,N_12958,N_12557);
nor U13097 (N_13097,N_12305,N_12917);
xnor U13098 (N_13098,N_12488,N_12287);
and U13099 (N_13099,N_12905,N_12192);
xor U13100 (N_13100,N_12555,N_12284);
xor U13101 (N_13101,N_12500,N_12248);
or U13102 (N_13102,N_12540,N_12186);
nand U13103 (N_13103,N_12520,N_12683);
or U13104 (N_13104,N_12084,N_12335);
nand U13105 (N_13105,N_12409,N_12816);
or U13106 (N_13106,N_12256,N_12155);
nor U13107 (N_13107,N_12384,N_12315);
nand U13108 (N_13108,N_12342,N_12620);
xnor U13109 (N_13109,N_12937,N_12952);
or U13110 (N_13110,N_12331,N_12487);
nand U13111 (N_13111,N_12366,N_12533);
nand U13112 (N_13112,N_12199,N_12224);
or U13113 (N_13113,N_12036,N_12503);
or U13114 (N_13114,N_12679,N_12723);
xor U13115 (N_13115,N_12636,N_12516);
or U13116 (N_13116,N_12541,N_12812);
nor U13117 (N_13117,N_12077,N_12865);
xor U13118 (N_13118,N_12652,N_12461);
nand U13119 (N_13119,N_12083,N_12370);
nand U13120 (N_13120,N_12463,N_12873);
xnor U13121 (N_13121,N_12551,N_12135);
xor U13122 (N_13122,N_12229,N_12295);
xnor U13123 (N_13123,N_12530,N_12206);
nor U13124 (N_13124,N_12825,N_12420);
nor U13125 (N_13125,N_12746,N_12583);
and U13126 (N_13126,N_12429,N_12008);
xor U13127 (N_13127,N_12213,N_12061);
and U13128 (N_13128,N_12235,N_12866);
xnor U13129 (N_13129,N_12445,N_12827);
nor U13130 (N_13130,N_12404,N_12888);
xnor U13131 (N_13131,N_12896,N_12241);
xnor U13132 (N_13132,N_12948,N_12718);
and U13133 (N_13133,N_12212,N_12945);
or U13134 (N_13134,N_12593,N_12830);
nand U13135 (N_13135,N_12983,N_12910);
nand U13136 (N_13136,N_12811,N_12715);
and U13137 (N_13137,N_12858,N_12223);
and U13138 (N_13138,N_12041,N_12147);
or U13139 (N_13139,N_12694,N_12271);
or U13140 (N_13140,N_12849,N_12643);
and U13141 (N_13141,N_12124,N_12875);
xnor U13142 (N_13142,N_12176,N_12527);
and U13143 (N_13143,N_12097,N_12215);
or U13144 (N_13144,N_12396,N_12296);
and U13145 (N_13145,N_12908,N_12470);
or U13146 (N_13146,N_12919,N_12792);
or U13147 (N_13147,N_12671,N_12231);
nand U13148 (N_13148,N_12356,N_12934);
nand U13149 (N_13149,N_12309,N_12843);
and U13150 (N_13150,N_12521,N_12783);
and U13151 (N_13151,N_12980,N_12890);
or U13152 (N_13152,N_12641,N_12290);
xnor U13153 (N_13153,N_12511,N_12345);
nor U13154 (N_13154,N_12173,N_12600);
or U13155 (N_13155,N_12504,N_12631);
xnor U13156 (N_13156,N_12027,N_12738);
xor U13157 (N_13157,N_12432,N_12855);
and U13158 (N_13158,N_12374,N_12423);
or U13159 (N_13159,N_12050,N_12286);
nor U13160 (N_13160,N_12730,N_12225);
and U13161 (N_13161,N_12647,N_12482);
nor U13162 (N_13162,N_12497,N_12656);
or U13163 (N_13163,N_12846,N_12351);
xor U13164 (N_13164,N_12379,N_12341);
or U13165 (N_13165,N_12988,N_12434);
nor U13166 (N_13166,N_12786,N_12024);
nor U13167 (N_13167,N_12648,N_12623);
or U13168 (N_13168,N_12771,N_12034);
and U13169 (N_13169,N_12191,N_12507);
or U13170 (N_13170,N_12372,N_12757);
xor U13171 (N_13171,N_12350,N_12226);
or U13172 (N_13172,N_12116,N_12052);
or U13173 (N_13173,N_12914,N_12701);
or U13174 (N_13174,N_12450,N_12458);
xnor U13175 (N_13175,N_12524,N_12844);
nand U13176 (N_13176,N_12940,N_12276);
nor U13177 (N_13177,N_12117,N_12687);
xnor U13178 (N_13178,N_12906,N_12925);
nor U13179 (N_13179,N_12015,N_12968);
nand U13180 (N_13180,N_12685,N_12108);
nand U13181 (N_13181,N_12616,N_12725);
or U13182 (N_13182,N_12740,N_12358);
xnor U13183 (N_13183,N_12727,N_12330);
and U13184 (N_13184,N_12814,N_12337);
xor U13185 (N_13185,N_12086,N_12582);
and U13186 (N_13186,N_12469,N_12377);
or U13187 (N_13187,N_12265,N_12359);
xor U13188 (N_13188,N_12526,N_12078);
and U13189 (N_13189,N_12602,N_12585);
nor U13190 (N_13190,N_12010,N_12502);
xnor U13191 (N_13191,N_12431,N_12056);
and U13192 (N_13192,N_12523,N_12928);
nor U13193 (N_13193,N_12595,N_12198);
nor U13194 (N_13194,N_12466,N_12788);
nand U13195 (N_13195,N_12261,N_12651);
or U13196 (N_13196,N_12997,N_12971);
nor U13197 (N_13197,N_12218,N_12796);
xor U13198 (N_13198,N_12001,N_12017);
nand U13199 (N_13199,N_12203,N_12617);
or U13200 (N_13200,N_12278,N_12005);
or U13201 (N_13201,N_12926,N_12571);
and U13202 (N_13202,N_12068,N_12809);
or U13203 (N_13203,N_12748,N_12307);
and U13204 (N_13204,N_12087,N_12672);
or U13205 (N_13205,N_12161,N_12070);
and U13206 (N_13206,N_12333,N_12961);
xnor U13207 (N_13207,N_12102,N_12773);
nor U13208 (N_13208,N_12160,N_12550);
nand U13209 (N_13209,N_12493,N_12513);
and U13210 (N_13210,N_12279,N_12800);
and U13211 (N_13211,N_12837,N_12382);
or U13212 (N_13212,N_12177,N_12572);
nand U13213 (N_13213,N_12949,N_12918);
xor U13214 (N_13214,N_12096,N_12883);
nand U13215 (N_13215,N_12085,N_12408);
and U13216 (N_13216,N_12898,N_12165);
xor U13217 (N_13217,N_12799,N_12438);
xnor U13218 (N_13218,N_12760,N_12728);
xnor U13219 (N_13219,N_12088,N_12764);
nand U13220 (N_13220,N_12343,N_12882);
nor U13221 (N_13221,N_12022,N_12777);
nand U13222 (N_13222,N_12698,N_12184);
nor U13223 (N_13223,N_12498,N_12146);
or U13224 (N_13224,N_12972,N_12303);
nor U13225 (N_13225,N_12413,N_12332);
or U13226 (N_13226,N_12828,N_12831);
nor U13227 (N_13227,N_12752,N_12334);
xor U13228 (N_13228,N_12492,N_12970);
nand U13229 (N_13229,N_12900,N_12804);
nor U13230 (N_13230,N_12886,N_12051);
nand U13231 (N_13231,N_12422,N_12584);
nor U13232 (N_13232,N_12721,N_12974);
nand U13233 (N_13233,N_12297,N_12109);
nor U13234 (N_13234,N_12864,N_12499);
xor U13235 (N_13235,N_12781,N_12870);
nand U13236 (N_13236,N_12838,N_12591);
xnor U13237 (N_13237,N_12892,N_12986);
or U13238 (N_13238,N_12514,N_12722);
and U13239 (N_13239,N_12440,N_12994);
or U13240 (N_13240,N_12901,N_12491);
nand U13241 (N_13241,N_12909,N_12711);
xor U13242 (N_13242,N_12232,N_12251);
nand U13243 (N_13243,N_12222,N_12594);
nor U13244 (N_13244,N_12378,N_12963);
nand U13245 (N_13245,N_12939,N_12750);
xor U13246 (N_13246,N_12893,N_12729);
xnor U13247 (N_13247,N_12302,N_12254);
nor U13248 (N_13248,N_12259,N_12196);
nand U13249 (N_13249,N_12327,N_12030);
nor U13250 (N_13250,N_12996,N_12467);
and U13251 (N_13251,N_12969,N_12696);
or U13252 (N_13252,N_12634,N_12565);
xor U13253 (N_13253,N_12115,N_12253);
and U13254 (N_13254,N_12689,N_12876);
or U13255 (N_13255,N_12707,N_12821);
or U13256 (N_13256,N_12043,N_12243);
or U13257 (N_13257,N_12111,N_12042);
nand U13258 (N_13258,N_12589,N_12581);
xor U13259 (N_13259,N_12233,N_12393);
nor U13260 (N_13260,N_12405,N_12023);
nand U13261 (N_13261,N_12978,N_12923);
nand U13262 (N_13262,N_12075,N_12753);
and U13263 (N_13263,N_12011,N_12269);
xnor U13264 (N_13264,N_12006,N_12455);
and U13265 (N_13265,N_12425,N_12158);
or U13266 (N_13266,N_12249,N_12483);
nand U13267 (N_13267,N_12299,N_12931);
xnor U13268 (N_13268,N_12114,N_12014);
or U13269 (N_13269,N_12941,N_12105);
xnor U13270 (N_13270,N_12283,N_12446);
or U13271 (N_13271,N_12732,N_12219);
nand U13272 (N_13272,N_12878,N_12183);
xor U13273 (N_13273,N_12793,N_12720);
or U13274 (N_13274,N_12549,N_12336);
xor U13275 (N_13275,N_12579,N_12806);
or U13276 (N_13276,N_12839,N_12151);
nand U13277 (N_13277,N_12272,N_12121);
nor U13278 (N_13278,N_12954,N_12780);
and U13279 (N_13279,N_12349,N_12355);
nand U13280 (N_13280,N_12110,N_12558);
nor U13281 (N_13281,N_12944,N_12619);
and U13282 (N_13282,N_12604,N_12590);
nand U13283 (N_13283,N_12460,N_12294);
or U13284 (N_13284,N_12339,N_12559);
xnor U13285 (N_13285,N_12673,N_12845);
nand U13286 (N_13286,N_12606,N_12125);
nor U13287 (N_13287,N_12699,N_12929);
nor U13288 (N_13288,N_12956,N_12026);
or U13289 (N_13289,N_12824,N_12536);
and U13290 (N_13290,N_12797,N_12618);
and U13291 (N_13291,N_12869,N_12388);
or U13292 (N_13292,N_12862,N_12790);
nor U13293 (N_13293,N_12216,N_12635);
or U13294 (N_13294,N_12419,N_12059);
nor U13295 (N_13295,N_12714,N_12509);
nor U13296 (N_13296,N_12993,N_12003);
xnor U13297 (N_13297,N_12767,N_12104);
and U13298 (N_13298,N_12140,N_12789);
and U13299 (N_13299,N_12414,N_12539);
or U13300 (N_13300,N_12435,N_12433);
nor U13301 (N_13301,N_12246,N_12028);
nand U13302 (N_13302,N_12586,N_12324);
xor U13303 (N_13303,N_12670,N_12237);
nand U13304 (N_13304,N_12368,N_12152);
and U13305 (N_13305,N_12924,N_12129);
nand U13306 (N_13306,N_12667,N_12567);
nor U13307 (N_13307,N_12535,N_12735);
and U13308 (N_13308,N_12476,N_12480);
nor U13309 (N_13309,N_12190,N_12992);
nand U13310 (N_13310,N_12205,N_12040);
xnor U13311 (N_13311,N_12239,N_12210);
or U13312 (N_13312,N_12383,N_12132);
nand U13313 (N_13313,N_12032,N_12802);
and U13314 (N_13314,N_12637,N_12960);
nor U13315 (N_13315,N_12805,N_12990);
nor U13316 (N_13316,N_12913,N_12363);
xor U13317 (N_13317,N_12847,N_12856);
or U13318 (N_13318,N_12188,N_12659);
xnor U13319 (N_13319,N_12543,N_12962);
and U13320 (N_13320,N_12236,N_12119);
nand U13321 (N_13321,N_12578,N_12037);
nor U13322 (N_13322,N_12947,N_12149);
xor U13323 (N_13323,N_12871,N_12660);
nor U13324 (N_13324,N_12977,N_12609);
xor U13325 (N_13325,N_12417,N_12568);
and U13326 (N_13326,N_12311,N_12306);
nand U13327 (N_13327,N_12495,N_12081);
and U13328 (N_13328,N_12756,N_12747);
and U13329 (N_13329,N_12922,N_12818);
xnor U13330 (N_13330,N_12772,N_12494);
nand U13331 (N_13331,N_12863,N_12247);
nand U13332 (N_13332,N_12984,N_12724);
nand U13333 (N_13333,N_12257,N_12853);
nor U13334 (N_13334,N_12542,N_12049);
xor U13335 (N_13335,N_12338,N_12282);
nand U13336 (N_13336,N_12563,N_12510);
nor U13337 (N_13337,N_12785,N_12669);
nor U13338 (N_13338,N_12608,N_12826);
nor U13339 (N_13339,N_12981,N_12441);
xor U13340 (N_13340,N_12758,N_12854);
xnor U13341 (N_13341,N_12552,N_12064);
nor U13342 (N_13342,N_12880,N_12411);
or U13343 (N_13343,N_12587,N_12680);
and U13344 (N_13344,N_12442,N_12318);
nor U13345 (N_13345,N_12464,N_12733);
nor U13346 (N_13346,N_12775,N_12228);
nor U13347 (N_13347,N_12456,N_12137);
and U13348 (N_13348,N_12761,N_12537);
nor U13349 (N_13349,N_12453,N_12505);
or U13350 (N_13350,N_12995,N_12071);
nand U13351 (N_13351,N_12038,N_12874);
xnor U13352 (N_13352,N_12554,N_12953);
or U13353 (N_13353,N_12674,N_12106);
nand U13354 (N_13354,N_12169,N_12653);
nand U13355 (N_13355,N_12895,N_12385);
nand U13356 (N_13356,N_12588,N_12200);
nand U13357 (N_13357,N_12107,N_12207);
and U13358 (N_13358,N_12428,N_12162);
xor U13359 (N_13359,N_12832,N_12478);
or U13360 (N_13360,N_12976,N_12397);
nand U13361 (N_13361,N_12300,N_12128);
nand U13362 (N_13362,N_12181,N_12047);
nand U13363 (N_13363,N_12650,N_12314);
nand U13364 (N_13364,N_12517,N_12798);
xnor U13365 (N_13365,N_12501,N_12291);
and U13366 (N_13366,N_12227,N_12255);
or U13367 (N_13367,N_12664,N_12702);
nor U13368 (N_13368,N_12020,N_12532);
or U13369 (N_13369,N_12529,N_12375);
nand U13370 (N_13370,N_12091,N_12308);
or U13371 (N_13371,N_12902,N_12930);
nand U13372 (N_13372,N_12407,N_12347);
nor U13373 (N_13373,N_12704,N_12700);
nand U13374 (N_13374,N_12185,N_12938);
or U13375 (N_13375,N_12369,N_12079);
and U13376 (N_13376,N_12769,N_12403);
and U13377 (N_13377,N_12645,N_12613);
xor U13378 (N_13378,N_12018,N_12973);
nand U13379 (N_13379,N_12851,N_12566);
and U13380 (N_13380,N_12402,N_12967);
nor U13381 (N_13381,N_12486,N_12127);
nand U13382 (N_13382,N_12118,N_12544);
and U13383 (N_13383,N_12245,N_12095);
or U13384 (N_13384,N_12039,N_12810);
nand U13385 (N_13385,N_12230,N_12734);
nor U13386 (N_13386,N_12763,N_12481);
nor U13387 (N_13387,N_12640,N_12598);
and U13388 (N_13388,N_12471,N_12401);
or U13389 (N_13389,N_12959,N_12007);
and U13390 (N_13390,N_12921,N_12813);
nor U13391 (N_13391,N_12365,N_12841);
and U13392 (N_13392,N_12891,N_12546);
nor U13393 (N_13393,N_12275,N_12731);
nor U13394 (N_13394,N_12774,N_12782);
nand U13395 (N_13395,N_12795,N_12710);
or U13396 (N_13396,N_12046,N_12658);
nor U13397 (N_13397,N_12688,N_12709);
or U13398 (N_13398,N_12274,N_12705);
nor U13399 (N_13399,N_12013,N_12157);
and U13400 (N_13400,N_12576,N_12823);
and U13401 (N_13401,N_12174,N_12156);
nor U13402 (N_13402,N_12394,N_12765);
nor U13403 (N_13403,N_12465,N_12596);
and U13404 (N_13404,N_12911,N_12678);
or U13405 (N_13405,N_12630,N_12665);
or U13406 (N_13406,N_12317,N_12447);
and U13407 (N_13407,N_12879,N_12406);
or U13408 (N_13408,N_12655,N_12416);
xnor U13409 (N_13409,N_12496,N_12894);
nand U13410 (N_13410,N_12234,N_12063);
nor U13411 (N_13411,N_12754,N_12449);
or U13412 (N_13412,N_12644,N_12889);
nand U13413 (N_13413,N_12749,N_12534);
and U13414 (N_13414,N_12019,N_12264);
and U13415 (N_13415,N_12985,N_12951);
xor U13416 (N_13416,N_12421,N_12292);
nand U13417 (N_13417,N_12603,N_12657);
or U13418 (N_13418,N_12545,N_12477);
xor U13419 (N_13419,N_12881,N_12611);
nor U13420 (N_13420,N_12277,N_12101);
and U13421 (N_13421,N_12561,N_12627);
xor U13422 (N_13422,N_12473,N_12113);
or U13423 (N_13423,N_12897,N_12144);
nor U13424 (N_13424,N_12055,N_12472);
nor U13425 (N_13425,N_12736,N_12768);
nand U13426 (N_13426,N_12076,N_12211);
xor U13427 (N_13427,N_12580,N_12170);
and U13428 (N_13428,N_12975,N_12933);
nand U13429 (N_13429,N_12391,N_12252);
nand U13430 (N_13430,N_12935,N_12717);
nand U13431 (N_13431,N_12268,N_12080);
nand U13432 (N_13432,N_12340,N_12320);
xor U13433 (N_13433,N_12475,N_12267);
and U13434 (N_13434,N_12662,N_12899);
xnor U13435 (N_13435,N_12323,N_12258);
nand U13436 (N_13436,N_12439,N_12298);
nand U13437 (N_13437,N_12266,N_12601);
nor U13438 (N_13438,N_12386,N_12638);
and U13439 (N_13439,N_12726,N_12691);
or U13440 (N_13440,N_12829,N_12133);
nor U13441 (N_13441,N_12744,N_12361);
nand U13442 (N_13442,N_12179,N_12328);
and U13443 (N_13443,N_12965,N_12706);
nor U13444 (N_13444,N_12820,N_12354);
or U13445 (N_13445,N_12217,N_12614);
nand U13446 (N_13446,N_12244,N_12936);
nand U13447 (N_13447,N_12167,N_12966);
nor U13448 (N_13448,N_12716,N_12834);
xor U13449 (N_13449,N_12194,N_12062);
and U13450 (N_13450,N_12979,N_12412);
and U13451 (N_13451,N_12803,N_12093);
xor U13452 (N_13452,N_12346,N_12000);
and U13453 (N_13453,N_12808,N_12569);
nor U13454 (N_13454,N_12313,N_12195);
nor U13455 (N_13455,N_12288,N_12451);
or U13456 (N_13456,N_12060,N_12122);
xor U13457 (N_13457,N_12426,N_12955);
xor U13458 (N_13458,N_12741,N_12281);
and U13459 (N_13459,N_12560,N_12836);
nor U13460 (N_13460,N_12148,N_12860);
or U13461 (N_13461,N_12163,N_12531);
xor U13462 (N_13462,N_12927,N_12138);
and U13463 (N_13463,N_12321,N_12573);
nand U13464 (N_13464,N_12371,N_12436);
nor U13465 (N_13465,N_12208,N_12835);
or U13466 (N_13466,N_12016,N_12639);
nor U13467 (N_13467,N_12329,N_12867);
nand U13468 (N_13468,N_12932,N_12666);
and U13469 (N_13469,N_12089,N_12861);
or U13470 (N_13470,N_12387,N_12316);
xnor U13471 (N_13471,N_12362,N_12987);
and U13472 (N_13472,N_12136,N_12755);
nand U13473 (N_13473,N_12762,N_12443);
nor U13474 (N_13474,N_12172,N_12263);
nor U13475 (N_13475,N_12991,N_12682);
or U13476 (N_13476,N_12376,N_12663);
or U13477 (N_13477,N_12240,N_12506);
nand U13478 (N_13478,N_12766,N_12564);
nand U13479 (N_13479,N_12399,N_12624);
or U13480 (N_13480,N_12357,N_12903);
nand U13481 (N_13481,N_12904,N_12178);
or U13482 (N_13482,N_12045,N_12444);
or U13483 (N_13483,N_12154,N_12815);
xnor U13484 (N_13484,N_12708,N_12859);
xnor U13485 (N_13485,N_12082,N_12142);
nand U13486 (N_13486,N_12677,N_12522);
nor U13487 (N_13487,N_12548,N_12848);
nor U13488 (N_13488,N_12610,N_12322);
or U13489 (N_13489,N_12395,N_12310);
nor U13490 (N_13490,N_12220,N_12326);
or U13491 (N_13491,N_12842,N_12098);
xor U13492 (N_13492,N_12012,N_12626);
and U13493 (N_13493,N_12801,N_12872);
nor U13494 (N_13494,N_12833,N_12092);
xnor U13495 (N_13495,N_12628,N_12739);
nor U13496 (N_13496,N_12398,N_12280);
nor U13497 (N_13497,N_12887,N_12794);
and U13498 (N_13498,N_12916,N_12686);
nor U13499 (N_13499,N_12654,N_12131);
nand U13500 (N_13500,N_12689,N_12594);
nand U13501 (N_13501,N_12897,N_12938);
and U13502 (N_13502,N_12031,N_12566);
nand U13503 (N_13503,N_12948,N_12482);
and U13504 (N_13504,N_12930,N_12449);
nand U13505 (N_13505,N_12274,N_12201);
xor U13506 (N_13506,N_12835,N_12961);
nor U13507 (N_13507,N_12616,N_12214);
and U13508 (N_13508,N_12853,N_12998);
or U13509 (N_13509,N_12965,N_12078);
and U13510 (N_13510,N_12258,N_12776);
xnor U13511 (N_13511,N_12825,N_12871);
and U13512 (N_13512,N_12928,N_12004);
or U13513 (N_13513,N_12020,N_12678);
nand U13514 (N_13514,N_12775,N_12982);
nor U13515 (N_13515,N_12779,N_12793);
and U13516 (N_13516,N_12687,N_12122);
and U13517 (N_13517,N_12072,N_12035);
nand U13518 (N_13518,N_12303,N_12578);
xnor U13519 (N_13519,N_12678,N_12627);
xnor U13520 (N_13520,N_12946,N_12373);
xnor U13521 (N_13521,N_12203,N_12785);
nand U13522 (N_13522,N_12991,N_12327);
xor U13523 (N_13523,N_12230,N_12251);
or U13524 (N_13524,N_12310,N_12867);
nand U13525 (N_13525,N_12619,N_12324);
or U13526 (N_13526,N_12485,N_12964);
nand U13527 (N_13527,N_12105,N_12108);
xnor U13528 (N_13528,N_12674,N_12335);
xor U13529 (N_13529,N_12179,N_12625);
and U13530 (N_13530,N_12695,N_12329);
and U13531 (N_13531,N_12673,N_12343);
xor U13532 (N_13532,N_12475,N_12509);
or U13533 (N_13533,N_12750,N_12214);
and U13534 (N_13534,N_12195,N_12474);
or U13535 (N_13535,N_12097,N_12818);
nor U13536 (N_13536,N_12036,N_12006);
xor U13537 (N_13537,N_12326,N_12076);
xnor U13538 (N_13538,N_12123,N_12708);
and U13539 (N_13539,N_12768,N_12093);
or U13540 (N_13540,N_12571,N_12561);
xor U13541 (N_13541,N_12046,N_12375);
xnor U13542 (N_13542,N_12769,N_12880);
xor U13543 (N_13543,N_12201,N_12684);
nand U13544 (N_13544,N_12070,N_12207);
nor U13545 (N_13545,N_12071,N_12270);
and U13546 (N_13546,N_12271,N_12792);
or U13547 (N_13547,N_12039,N_12798);
nand U13548 (N_13548,N_12411,N_12682);
or U13549 (N_13549,N_12925,N_12810);
nand U13550 (N_13550,N_12235,N_12528);
xor U13551 (N_13551,N_12385,N_12553);
and U13552 (N_13552,N_12635,N_12275);
nor U13553 (N_13553,N_12893,N_12259);
or U13554 (N_13554,N_12345,N_12123);
nand U13555 (N_13555,N_12491,N_12451);
nand U13556 (N_13556,N_12024,N_12555);
and U13557 (N_13557,N_12658,N_12966);
or U13558 (N_13558,N_12528,N_12304);
nand U13559 (N_13559,N_12693,N_12055);
nor U13560 (N_13560,N_12759,N_12153);
xor U13561 (N_13561,N_12068,N_12299);
or U13562 (N_13562,N_12021,N_12119);
nor U13563 (N_13563,N_12202,N_12733);
or U13564 (N_13564,N_12223,N_12802);
xnor U13565 (N_13565,N_12083,N_12448);
and U13566 (N_13566,N_12893,N_12056);
or U13567 (N_13567,N_12726,N_12722);
xnor U13568 (N_13568,N_12536,N_12488);
xnor U13569 (N_13569,N_12591,N_12624);
and U13570 (N_13570,N_12872,N_12899);
nor U13571 (N_13571,N_12074,N_12594);
or U13572 (N_13572,N_12226,N_12320);
and U13573 (N_13573,N_12207,N_12047);
nor U13574 (N_13574,N_12461,N_12936);
nor U13575 (N_13575,N_12874,N_12351);
nor U13576 (N_13576,N_12845,N_12025);
and U13577 (N_13577,N_12423,N_12092);
nand U13578 (N_13578,N_12946,N_12144);
or U13579 (N_13579,N_12345,N_12809);
or U13580 (N_13580,N_12018,N_12050);
and U13581 (N_13581,N_12092,N_12179);
xor U13582 (N_13582,N_12494,N_12373);
or U13583 (N_13583,N_12595,N_12457);
or U13584 (N_13584,N_12739,N_12660);
xnor U13585 (N_13585,N_12169,N_12905);
nand U13586 (N_13586,N_12372,N_12245);
nand U13587 (N_13587,N_12630,N_12010);
xnor U13588 (N_13588,N_12806,N_12351);
xnor U13589 (N_13589,N_12383,N_12709);
xnor U13590 (N_13590,N_12381,N_12780);
or U13591 (N_13591,N_12119,N_12332);
xor U13592 (N_13592,N_12568,N_12709);
nand U13593 (N_13593,N_12268,N_12605);
or U13594 (N_13594,N_12246,N_12539);
xnor U13595 (N_13595,N_12482,N_12257);
and U13596 (N_13596,N_12003,N_12685);
or U13597 (N_13597,N_12641,N_12766);
xor U13598 (N_13598,N_12595,N_12688);
nand U13599 (N_13599,N_12206,N_12356);
xnor U13600 (N_13600,N_12844,N_12166);
nand U13601 (N_13601,N_12127,N_12762);
or U13602 (N_13602,N_12074,N_12193);
and U13603 (N_13603,N_12309,N_12961);
xnor U13604 (N_13604,N_12385,N_12548);
nor U13605 (N_13605,N_12560,N_12199);
nor U13606 (N_13606,N_12081,N_12942);
nand U13607 (N_13607,N_12608,N_12148);
xor U13608 (N_13608,N_12300,N_12307);
nand U13609 (N_13609,N_12847,N_12745);
or U13610 (N_13610,N_12629,N_12156);
nor U13611 (N_13611,N_12079,N_12247);
nand U13612 (N_13612,N_12792,N_12313);
or U13613 (N_13613,N_12955,N_12509);
xor U13614 (N_13614,N_12817,N_12601);
xnor U13615 (N_13615,N_12223,N_12850);
nor U13616 (N_13616,N_12596,N_12161);
xor U13617 (N_13617,N_12091,N_12297);
and U13618 (N_13618,N_12039,N_12409);
nor U13619 (N_13619,N_12468,N_12384);
nand U13620 (N_13620,N_12320,N_12323);
nand U13621 (N_13621,N_12978,N_12885);
nor U13622 (N_13622,N_12091,N_12901);
xnor U13623 (N_13623,N_12007,N_12421);
or U13624 (N_13624,N_12427,N_12886);
and U13625 (N_13625,N_12592,N_12892);
and U13626 (N_13626,N_12871,N_12700);
nand U13627 (N_13627,N_12349,N_12847);
nand U13628 (N_13628,N_12389,N_12776);
or U13629 (N_13629,N_12622,N_12010);
nor U13630 (N_13630,N_12720,N_12301);
and U13631 (N_13631,N_12194,N_12014);
or U13632 (N_13632,N_12188,N_12204);
xnor U13633 (N_13633,N_12784,N_12184);
and U13634 (N_13634,N_12773,N_12160);
nor U13635 (N_13635,N_12170,N_12512);
and U13636 (N_13636,N_12500,N_12809);
nand U13637 (N_13637,N_12836,N_12464);
nor U13638 (N_13638,N_12216,N_12211);
or U13639 (N_13639,N_12023,N_12940);
and U13640 (N_13640,N_12811,N_12630);
and U13641 (N_13641,N_12739,N_12280);
xnor U13642 (N_13642,N_12046,N_12393);
nor U13643 (N_13643,N_12878,N_12093);
nor U13644 (N_13644,N_12581,N_12619);
and U13645 (N_13645,N_12743,N_12829);
and U13646 (N_13646,N_12967,N_12021);
and U13647 (N_13647,N_12816,N_12207);
nor U13648 (N_13648,N_12060,N_12130);
nor U13649 (N_13649,N_12991,N_12126);
nor U13650 (N_13650,N_12606,N_12447);
nand U13651 (N_13651,N_12273,N_12066);
and U13652 (N_13652,N_12591,N_12584);
nand U13653 (N_13653,N_12821,N_12891);
xnor U13654 (N_13654,N_12837,N_12595);
nor U13655 (N_13655,N_12529,N_12838);
nand U13656 (N_13656,N_12760,N_12732);
xnor U13657 (N_13657,N_12273,N_12209);
or U13658 (N_13658,N_12622,N_12521);
nor U13659 (N_13659,N_12916,N_12312);
nor U13660 (N_13660,N_12054,N_12258);
xor U13661 (N_13661,N_12711,N_12537);
nand U13662 (N_13662,N_12081,N_12304);
xnor U13663 (N_13663,N_12424,N_12723);
xor U13664 (N_13664,N_12511,N_12410);
nand U13665 (N_13665,N_12650,N_12909);
and U13666 (N_13666,N_12888,N_12811);
xor U13667 (N_13667,N_12891,N_12429);
or U13668 (N_13668,N_12698,N_12243);
or U13669 (N_13669,N_12459,N_12040);
and U13670 (N_13670,N_12662,N_12004);
nor U13671 (N_13671,N_12697,N_12520);
xor U13672 (N_13672,N_12351,N_12559);
or U13673 (N_13673,N_12018,N_12535);
nor U13674 (N_13674,N_12849,N_12996);
and U13675 (N_13675,N_12829,N_12430);
nand U13676 (N_13676,N_12879,N_12921);
nor U13677 (N_13677,N_12409,N_12555);
and U13678 (N_13678,N_12875,N_12084);
or U13679 (N_13679,N_12400,N_12518);
nor U13680 (N_13680,N_12268,N_12288);
and U13681 (N_13681,N_12958,N_12164);
and U13682 (N_13682,N_12828,N_12283);
and U13683 (N_13683,N_12093,N_12640);
nand U13684 (N_13684,N_12177,N_12513);
and U13685 (N_13685,N_12066,N_12871);
nor U13686 (N_13686,N_12382,N_12773);
xnor U13687 (N_13687,N_12032,N_12654);
nand U13688 (N_13688,N_12351,N_12386);
xor U13689 (N_13689,N_12878,N_12577);
or U13690 (N_13690,N_12230,N_12585);
and U13691 (N_13691,N_12754,N_12334);
nand U13692 (N_13692,N_12773,N_12928);
nor U13693 (N_13693,N_12725,N_12274);
nand U13694 (N_13694,N_12304,N_12992);
or U13695 (N_13695,N_12309,N_12789);
and U13696 (N_13696,N_12563,N_12719);
nand U13697 (N_13697,N_12191,N_12114);
nand U13698 (N_13698,N_12742,N_12715);
xnor U13699 (N_13699,N_12641,N_12604);
nor U13700 (N_13700,N_12238,N_12449);
xnor U13701 (N_13701,N_12801,N_12693);
xor U13702 (N_13702,N_12203,N_12882);
and U13703 (N_13703,N_12849,N_12787);
xor U13704 (N_13704,N_12754,N_12189);
xnor U13705 (N_13705,N_12887,N_12752);
and U13706 (N_13706,N_12236,N_12170);
and U13707 (N_13707,N_12136,N_12451);
or U13708 (N_13708,N_12143,N_12839);
xnor U13709 (N_13709,N_12773,N_12220);
and U13710 (N_13710,N_12953,N_12012);
xor U13711 (N_13711,N_12862,N_12257);
nand U13712 (N_13712,N_12511,N_12532);
nand U13713 (N_13713,N_12879,N_12789);
xor U13714 (N_13714,N_12832,N_12066);
or U13715 (N_13715,N_12394,N_12446);
nor U13716 (N_13716,N_12874,N_12291);
or U13717 (N_13717,N_12583,N_12071);
xnor U13718 (N_13718,N_12494,N_12827);
xor U13719 (N_13719,N_12942,N_12857);
or U13720 (N_13720,N_12452,N_12816);
nand U13721 (N_13721,N_12920,N_12577);
or U13722 (N_13722,N_12083,N_12434);
xnor U13723 (N_13723,N_12956,N_12397);
nand U13724 (N_13724,N_12108,N_12765);
nor U13725 (N_13725,N_12290,N_12465);
or U13726 (N_13726,N_12326,N_12565);
nand U13727 (N_13727,N_12869,N_12684);
and U13728 (N_13728,N_12886,N_12598);
nand U13729 (N_13729,N_12324,N_12769);
nand U13730 (N_13730,N_12948,N_12121);
and U13731 (N_13731,N_12727,N_12490);
nand U13732 (N_13732,N_12024,N_12046);
xor U13733 (N_13733,N_12301,N_12330);
xnor U13734 (N_13734,N_12891,N_12726);
and U13735 (N_13735,N_12804,N_12449);
and U13736 (N_13736,N_12560,N_12548);
and U13737 (N_13737,N_12825,N_12750);
and U13738 (N_13738,N_12093,N_12398);
or U13739 (N_13739,N_12927,N_12624);
or U13740 (N_13740,N_12363,N_12851);
xnor U13741 (N_13741,N_12529,N_12129);
xor U13742 (N_13742,N_12856,N_12990);
xor U13743 (N_13743,N_12303,N_12374);
and U13744 (N_13744,N_12595,N_12854);
nor U13745 (N_13745,N_12630,N_12900);
nand U13746 (N_13746,N_12342,N_12789);
nand U13747 (N_13747,N_12525,N_12441);
and U13748 (N_13748,N_12193,N_12987);
or U13749 (N_13749,N_12313,N_12444);
nor U13750 (N_13750,N_12193,N_12069);
nor U13751 (N_13751,N_12692,N_12646);
nor U13752 (N_13752,N_12878,N_12394);
and U13753 (N_13753,N_12164,N_12702);
nor U13754 (N_13754,N_12136,N_12719);
nor U13755 (N_13755,N_12659,N_12558);
xnor U13756 (N_13756,N_12608,N_12330);
nor U13757 (N_13757,N_12235,N_12681);
nand U13758 (N_13758,N_12294,N_12363);
xor U13759 (N_13759,N_12907,N_12535);
or U13760 (N_13760,N_12607,N_12052);
xnor U13761 (N_13761,N_12654,N_12177);
nand U13762 (N_13762,N_12183,N_12517);
nand U13763 (N_13763,N_12820,N_12043);
or U13764 (N_13764,N_12872,N_12295);
xnor U13765 (N_13765,N_12179,N_12297);
xnor U13766 (N_13766,N_12723,N_12874);
nand U13767 (N_13767,N_12878,N_12008);
or U13768 (N_13768,N_12996,N_12990);
nor U13769 (N_13769,N_12450,N_12436);
and U13770 (N_13770,N_12654,N_12663);
xor U13771 (N_13771,N_12741,N_12129);
and U13772 (N_13772,N_12760,N_12272);
and U13773 (N_13773,N_12094,N_12663);
nor U13774 (N_13774,N_12714,N_12366);
nor U13775 (N_13775,N_12315,N_12400);
nor U13776 (N_13776,N_12565,N_12891);
nand U13777 (N_13777,N_12435,N_12008);
nor U13778 (N_13778,N_12542,N_12260);
or U13779 (N_13779,N_12098,N_12417);
and U13780 (N_13780,N_12501,N_12899);
and U13781 (N_13781,N_12990,N_12304);
and U13782 (N_13782,N_12230,N_12133);
xnor U13783 (N_13783,N_12331,N_12187);
nor U13784 (N_13784,N_12758,N_12328);
and U13785 (N_13785,N_12436,N_12570);
and U13786 (N_13786,N_12101,N_12340);
xnor U13787 (N_13787,N_12071,N_12142);
nand U13788 (N_13788,N_12397,N_12351);
nand U13789 (N_13789,N_12240,N_12457);
nor U13790 (N_13790,N_12592,N_12633);
or U13791 (N_13791,N_12119,N_12719);
nor U13792 (N_13792,N_12485,N_12778);
nand U13793 (N_13793,N_12473,N_12659);
nor U13794 (N_13794,N_12157,N_12325);
nand U13795 (N_13795,N_12617,N_12963);
nor U13796 (N_13796,N_12121,N_12330);
nor U13797 (N_13797,N_12281,N_12197);
nand U13798 (N_13798,N_12556,N_12994);
and U13799 (N_13799,N_12677,N_12251);
nand U13800 (N_13800,N_12967,N_12479);
xnor U13801 (N_13801,N_12955,N_12750);
nor U13802 (N_13802,N_12103,N_12276);
or U13803 (N_13803,N_12360,N_12720);
nor U13804 (N_13804,N_12165,N_12455);
nor U13805 (N_13805,N_12731,N_12988);
nor U13806 (N_13806,N_12864,N_12949);
xnor U13807 (N_13807,N_12866,N_12032);
and U13808 (N_13808,N_12818,N_12714);
nor U13809 (N_13809,N_12766,N_12674);
nand U13810 (N_13810,N_12017,N_12577);
or U13811 (N_13811,N_12974,N_12518);
or U13812 (N_13812,N_12886,N_12358);
and U13813 (N_13813,N_12244,N_12721);
nor U13814 (N_13814,N_12216,N_12177);
xnor U13815 (N_13815,N_12670,N_12651);
xnor U13816 (N_13816,N_12181,N_12756);
nor U13817 (N_13817,N_12132,N_12080);
and U13818 (N_13818,N_12704,N_12204);
nand U13819 (N_13819,N_12471,N_12015);
xnor U13820 (N_13820,N_12276,N_12005);
or U13821 (N_13821,N_12666,N_12489);
and U13822 (N_13822,N_12537,N_12400);
or U13823 (N_13823,N_12514,N_12578);
nand U13824 (N_13824,N_12199,N_12693);
nand U13825 (N_13825,N_12001,N_12454);
or U13826 (N_13826,N_12451,N_12240);
nand U13827 (N_13827,N_12635,N_12287);
nand U13828 (N_13828,N_12556,N_12905);
xnor U13829 (N_13829,N_12164,N_12301);
or U13830 (N_13830,N_12292,N_12636);
or U13831 (N_13831,N_12268,N_12067);
nor U13832 (N_13832,N_12559,N_12018);
nor U13833 (N_13833,N_12934,N_12939);
nand U13834 (N_13834,N_12349,N_12078);
and U13835 (N_13835,N_12266,N_12134);
nand U13836 (N_13836,N_12773,N_12499);
nor U13837 (N_13837,N_12233,N_12343);
nor U13838 (N_13838,N_12381,N_12202);
and U13839 (N_13839,N_12075,N_12213);
nor U13840 (N_13840,N_12589,N_12283);
xor U13841 (N_13841,N_12697,N_12237);
xor U13842 (N_13842,N_12868,N_12602);
or U13843 (N_13843,N_12033,N_12172);
or U13844 (N_13844,N_12269,N_12055);
xnor U13845 (N_13845,N_12633,N_12312);
nand U13846 (N_13846,N_12349,N_12751);
or U13847 (N_13847,N_12160,N_12417);
xor U13848 (N_13848,N_12974,N_12604);
nand U13849 (N_13849,N_12103,N_12804);
and U13850 (N_13850,N_12252,N_12866);
and U13851 (N_13851,N_12492,N_12546);
and U13852 (N_13852,N_12756,N_12642);
xnor U13853 (N_13853,N_12778,N_12374);
xor U13854 (N_13854,N_12268,N_12892);
nor U13855 (N_13855,N_12568,N_12380);
and U13856 (N_13856,N_12360,N_12079);
xnor U13857 (N_13857,N_12361,N_12958);
nand U13858 (N_13858,N_12084,N_12870);
nand U13859 (N_13859,N_12258,N_12787);
nor U13860 (N_13860,N_12605,N_12703);
nor U13861 (N_13861,N_12430,N_12295);
xnor U13862 (N_13862,N_12247,N_12928);
or U13863 (N_13863,N_12164,N_12816);
or U13864 (N_13864,N_12584,N_12020);
and U13865 (N_13865,N_12807,N_12456);
nor U13866 (N_13866,N_12854,N_12674);
or U13867 (N_13867,N_12433,N_12417);
or U13868 (N_13868,N_12803,N_12799);
and U13869 (N_13869,N_12132,N_12796);
nor U13870 (N_13870,N_12636,N_12370);
nor U13871 (N_13871,N_12511,N_12255);
nand U13872 (N_13872,N_12633,N_12942);
xor U13873 (N_13873,N_12445,N_12870);
nor U13874 (N_13874,N_12247,N_12644);
nor U13875 (N_13875,N_12984,N_12601);
or U13876 (N_13876,N_12957,N_12946);
xor U13877 (N_13877,N_12294,N_12897);
nor U13878 (N_13878,N_12158,N_12122);
nor U13879 (N_13879,N_12057,N_12883);
nand U13880 (N_13880,N_12284,N_12344);
and U13881 (N_13881,N_12122,N_12696);
and U13882 (N_13882,N_12209,N_12253);
or U13883 (N_13883,N_12800,N_12896);
nor U13884 (N_13884,N_12159,N_12873);
and U13885 (N_13885,N_12215,N_12419);
or U13886 (N_13886,N_12276,N_12230);
nand U13887 (N_13887,N_12756,N_12530);
and U13888 (N_13888,N_12932,N_12981);
nor U13889 (N_13889,N_12617,N_12313);
nand U13890 (N_13890,N_12765,N_12189);
or U13891 (N_13891,N_12579,N_12241);
nand U13892 (N_13892,N_12419,N_12407);
and U13893 (N_13893,N_12724,N_12331);
xnor U13894 (N_13894,N_12554,N_12328);
and U13895 (N_13895,N_12901,N_12354);
nand U13896 (N_13896,N_12200,N_12105);
or U13897 (N_13897,N_12798,N_12590);
xnor U13898 (N_13898,N_12789,N_12487);
or U13899 (N_13899,N_12473,N_12414);
or U13900 (N_13900,N_12536,N_12474);
xor U13901 (N_13901,N_12894,N_12852);
and U13902 (N_13902,N_12453,N_12020);
nand U13903 (N_13903,N_12919,N_12215);
or U13904 (N_13904,N_12403,N_12475);
xor U13905 (N_13905,N_12184,N_12357);
nand U13906 (N_13906,N_12748,N_12911);
xnor U13907 (N_13907,N_12314,N_12265);
nand U13908 (N_13908,N_12798,N_12885);
and U13909 (N_13909,N_12210,N_12221);
xor U13910 (N_13910,N_12433,N_12752);
or U13911 (N_13911,N_12990,N_12932);
or U13912 (N_13912,N_12328,N_12211);
nand U13913 (N_13913,N_12161,N_12350);
nor U13914 (N_13914,N_12503,N_12106);
and U13915 (N_13915,N_12845,N_12498);
nand U13916 (N_13916,N_12531,N_12812);
and U13917 (N_13917,N_12667,N_12146);
and U13918 (N_13918,N_12011,N_12231);
nor U13919 (N_13919,N_12206,N_12875);
or U13920 (N_13920,N_12119,N_12927);
nor U13921 (N_13921,N_12831,N_12000);
or U13922 (N_13922,N_12359,N_12066);
nor U13923 (N_13923,N_12834,N_12457);
and U13924 (N_13924,N_12237,N_12962);
or U13925 (N_13925,N_12189,N_12543);
nand U13926 (N_13926,N_12996,N_12279);
nor U13927 (N_13927,N_12873,N_12683);
and U13928 (N_13928,N_12158,N_12236);
or U13929 (N_13929,N_12562,N_12438);
or U13930 (N_13930,N_12373,N_12824);
xnor U13931 (N_13931,N_12535,N_12380);
and U13932 (N_13932,N_12134,N_12651);
nand U13933 (N_13933,N_12753,N_12758);
and U13934 (N_13934,N_12368,N_12055);
nand U13935 (N_13935,N_12001,N_12943);
nand U13936 (N_13936,N_12950,N_12471);
xor U13937 (N_13937,N_12503,N_12982);
nand U13938 (N_13938,N_12844,N_12510);
nand U13939 (N_13939,N_12206,N_12181);
xor U13940 (N_13940,N_12617,N_12138);
nor U13941 (N_13941,N_12542,N_12728);
nand U13942 (N_13942,N_12899,N_12983);
xor U13943 (N_13943,N_12681,N_12851);
or U13944 (N_13944,N_12035,N_12389);
or U13945 (N_13945,N_12410,N_12418);
nand U13946 (N_13946,N_12774,N_12130);
and U13947 (N_13947,N_12080,N_12154);
nand U13948 (N_13948,N_12864,N_12915);
nand U13949 (N_13949,N_12959,N_12868);
and U13950 (N_13950,N_12265,N_12113);
xnor U13951 (N_13951,N_12223,N_12785);
nor U13952 (N_13952,N_12960,N_12566);
xnor U13953 (N_13953,N_12776,N_12441);
nor U13954 (N_13954,N_12165,N_12891);
and U13955 (N_13955,N_12066,N_12416);
nor U13956 (N_13956,N_12743,N_12272);
nor U13957 (N_13957,N_12602,N_12543);
nand U13958 (N_13958,N_12216,N_12731);
nor U13959 (N_13959,N_12952,N_12105);
and U13960 (N_13960,N_12162,N_12115);
nand U13961 (N_13961,N_12114,N_12381);
xnor U13962 (N_13962,N_12773,N_12197);
nand U13963 (N_13963,N_12543,N_12277);
nand U13964 (N_13964,N_12104,N_12123);
nand U13965 (N_13965,N_12721,N_12336);
or U13966 (N_13966,N_12200,N_12747);
or U13967 (N_13967,N_12778,N_12605);
or U13968 (N_13968,N_12862,N_12564);
and U13969 (N_13969,N_12267,N_12121);
and U13970 (N_13970,N_12702,N_12905);
xor U13971 (N_13971,N_12324,N_12144);
or U13972 (N_13972,N_12788,N_12794);
xor U13973 (N_13973,N_12536,N_12435);
nand U13974 (N_13974,N_12031,N_12573);
nor U13975 (N_13975,N_12162,N_12993);
xor U13976 (N_13976,N_12905,N_12837);
and U13977 (N_13977,N_12779,N_12314);
nand U13978 (N_13978,N_12882,N_12028);
nor U13979 (N_13979,N_12469,N_12536);
nand U13980 (N_13980,N_12109,N_12117);
and U13981 (N_13981,N_12370,N_12675);
or U13982 (N_13982,N_12392,N_12089);
nand U13983 (N_13983,N_12217,N_12808);
and U13984 (N_13984,N_12483,N_12932);
xnor U13985 (N_13985,N_12467,N_12226);
xor U13986 (N_13986,N_12208,N_12291);
and U13987 (N_13987,N_12832,N_12216);
nand U13988 (N_13988,N_12743,N_12726);
nand U13989 (N_13989,N_12486,N_12740);
or U13990 (N_13990,N_12663,N_12133);
or U13991 (N_13991,N_12568,N_12276);
nand U13992 (N_13992,N_12834,N_12459);
or U13993 (N_13993,N_12195,N_12424);
nor U13994 (N_13994,N_12380,N_12614);
nor U13995 (N_13995,N_12690,N_12403);
or U13996 (N_13996,N_12024,N_12067);
or U13997 (N_13997,N_12488,N_12220);
nor U13998 (N_13998,N_12688,N_12757);
or U13999 (N_13999,N_12434,N_12822);
nand U14000 (N_14000,N_13049,N_13184);
nand U14001 (N_14001,N_13248,N_13658);
xor U14002 (N_14002,N_13554,N_13315);
nand U14003 (N_14003,N_13696,N_13317);
or U14004 (N_14004,N_13560,N_13744);
xor U14005 (N_14005,N_13760,N_13603);
and U14006 (N_14006,N_13091,N_13322);
xor U14007 (N_14007,N_13319,N_13213);
or U14008 (N_14008,N_13572,N_13855);
and U14009 (N_14009,N_13454,N_13134);
or U14010 (N_14010,N_13095,N_13373);
or U14011 (N_14011,N_13178,N_13848);
xor U14012 (N_14012,N_13298,N_13456);
or U14013 (N_14013,N_13871,N_13720);
or U14014 (N_14014,N_13902,N_13507);
or U14015 (N_14015,N_13958,N_13064);
or U14016 (N_14016,N_13736,N_13039);
nand U14017 (N_14017,N_13909,N_13020);
nand U14018 (N_14018,N_13687,N_13003);
or U14019 (N_14019,N_13180,N_13277);
xor U14020 (N_14020,N_13547,N_13903);
nand U14021 (N_14021,N_13432,N_13475);
or U14022 (N_14022,N_13441,N_13154);
xnor U14023 (N_14023,N_13991,N_13998);
and U14024 (N_14024,N_13098,N_13934);
xnor U14025 (N_14025,N_13664,N_13831);
and U14026 (N_14026,N_13022,N_13127);
xnor U14027 (N_14027,N_13961,N_13829);
and U14028 (N_14028,N_13533,N_13637);
or U14029 (N_14029,N_13989,N_13173);
and U14030 (N_14030,N_13258,N_13847);
or U14031 (N_14031,N_13113,N_13701);
and U14032 (N_14032,N_13549,N_13573);
or U14033 (N_14033,N_13659,N_13815);
nand U14034 (N_14034,N_13785,N_13191);
nor U14035 (N_14035,N_13527,N_13017);
or U14036 (N_14036,N_13399,N_13293);
or U14037 (N_14037,N_13587,N_13806);
and U14038 (N_14038,N_13811,N_13202);
nor U14039 (N_14039,N_13254,N_13510);
nand U14040 (N_14040,N_13261,N_13114);
and U14041 (N_14041,N_13329,N_13429);
nor U14042 (N_14042,N_13296,N_13633);
xor U14043 (N_14043,N_13438,N_13155);
or U14044 (N_14044,N_13337,N_13892);
xnor U14045 (N_14045,N_13595,N_13713);
and U14046 (N_14046,N_13052,N_13339);
nor U14047 (N_14047,N_13000,N_13336);
or U14048 (N_14048,N_13644,N_13634);
and U14049 (N_14049,N_13009,N_13354);
nand U14050 (N_14050,N_13726,N_13236);
nor U14051 (N_14051,N_13818,N_13118);
xor U14052 (N_14052,N_13038,N_13823);
or U14053 (N_14053,N_13982,N_13085);
nor U14054 (N_14054,N_13410,N_13120);
xnor U14055 (N_14055,N_13156,N_13538);
and U14056 (N_14056,N_13645,N_13467);
or U14057 (N_14057,N_13711,N_13469);
or U14058 (N_14058,N_13259,N_13376);
xor U14059 (N_14059,N_13845,N_13166);
nand U14060 (N_14060,N_13981,N_13087);
xor U14061 (N_14061,N_13448,N_13552);
xor U14062 (N_14062,N_13840,N_13241);
and U14063 (N_14063,N_13660,N_13514);
nand U14064 (N_14064,N_13382,N_13649);
or U14065 (N_14065,N_13655,N_13117);
and U14066 (N_14066,N_13235,N_13297);
xnor U14067 (N_14067,N_13986,N_13607);
nor U14068 (N_14068,N_13027,N_13500);
nand U14069 (N_14069,N_13068,N_13995);
xor U14070 (N_14070,N_13691,N_13486);
nand U14071 (N_14071,N_13937,N_13632);
nand U14072 (N_14072,N_13016,N_13598);
or U14073 (N_14073,N_13985,N_13565);
nand U14074 (N_14074,N_13733,N_13051);
xnor U14075 (N_14075,N_13627,N_13749);
nor U14076 (N_14076,N_13047,N_13103);
and U14077 (N_14077,N_13819,N_13199);
and U14078 (N_14078,N_13451,N_13046);
and U14079 (N_14079,N_13057,N_13231);
or U14080 (N_14080,N_13245,N_13251);
xor U14081 (N_14081,N_13616,N_13563);
or U14082 (N_14082,N_13576,N_13387);
nor U14083 (N_14083,N_13792,N_13423);
xor U14084 (N_14084,N_13752,N_13705);
nor U14085 (N_14085,N_13066,N_13888);
nand U14086 (N_14086,N_13464,N_13877);
nor U14087 (N_14087,N_13583,N_13667);
or U14088 (N_14088,N_13569,N_13625);
and U14089 (N_14089,N_13025,N_13215);
nand U14090 (N_14090,N_13710,N_13082);
xnor U14091 (N_14091,N_13544,N_13990);
nand U14092 (N_14092,N_13161,N_13348);
nand U14093 (N_14093,N_13663,N_13487);
nor U14094 (N_14094,N_13176,N_13287);
xnor U14095 (N_14095,N_13882,N_13345);
and U14096 (N_14096,N_13588,N_13568);
or U14097 (N_14097,N_13474,N_13775);
and U14098 (N_14098,N_13683,N_13124);
nor U14099 (N_14099,N_13478,N_13876);
nand U14100 (N_14100,N_13657,N_13431);
or U14101 (N_14101,N_13362,N_13269);
nand U14102 (N_14102,N_13366,N_13030);
and U14103 (N_14103,N_13965,N_13401);
or U14104 (N_14104,N_13940,N_13735);
nor U14105 (N_14105,N_13837,N_13140);
xor U14106 (N_14106,N_13642,N_13971);
xnor U14107 (N_14107,N_13872,N_13135);
nand U14108 (N_14108,N_13650,N_13255);
nor U14109 (N_14109,N_13923,N_13916);
xor U14110 (N_14110,N_13243,N_13369);
nand U14111 (N_14111,N_13935,N_13518);
or U14112 (N_14112,N_13630,N_13945);
or U14113 (N_14113,N_13090,N_13280);
xor U14114 (N_14114,N_13232,N_13508);
nand U14115 (N_14115,N_13577,N_13059);
or U14116 (N_14116,N_13150,N_13954);
nand U14117 (N_14117,N_13446,N_13273);
nand U14118 (N_14118,N_13955,N_13521);
nand U14119 (N_14119,N_13162,N_13686);
or U14120 (N_14120,N_13706,N_13968);
nand U14121 (N_14121,N_13602,N_13417);
and U14122 (N_14122,N_13962,N_13946);
nand U14123 (N_14123,N_13033,N_13424);
xnor U14124 (N_14124,N_13041,N_13788);
and U14125 (N_14125,N_13580,N_13026);
nor U14126 (N_14126,N_13942,N_13192);
and U14127 (N_14127,N_13647,N_13160);
nand U14128 (N_14128,N_13987,N_13597);
nor U14129 (N_14129,N_13719,N_13921);
nand U14130 (N_14130,N_13931,N_13964);
nor U14131 (N_14131,N_13874,N_13693);
nor U14132 (N_14132,N_13485,N_13895);
xnor U14133 (N_14133,N_13730,N_13018);
xor U14134 (N_14134,N_13707,N_13671);
nand U14135 (N_14135,N_13759,N_13128);
xor U14136 (N_14136,N_13624,N_13629);
nor U14137 (N_14137,N_13949,N_13996);
or U14138 (N_14138,N_13307,N_13078);
nor U14139 (N_14139,N_13428,N_13434);
xnor U14140 (N_14140,N_13757,N_13409);
or U14141 (N_14141,N_13076,N_13218);
nand U14142 (N_14142,N_13321,N_13360);
and U14143 (N_14143,N_13539,N_13926);
or U14144 (N_14144,N_13503,N_13787);
and U14145 (N_14145,N_13543,N_13195);
nor U14146 (N_14146,N_13004,N_13656);
and U14147 (N_14147,N_13661,N_13748);
or U14148 (N_14148,N_13574,N_13139);
or U14149 (N_14149,N_13217,N_13562);
and U14150 (N_14150,N_13021,N_13072);
or U14151 (N_14151,N_13074,N_13152);
or U14152 (N_14152,N_13688,N_13812);
or U14153 (N_14153,N_13918,N_13083);
xnor U14154 (N_14154,N_13879,N_13679);
nand U14155 (N_14155,N_13861,N_13612);
nand U14156 (N_14156,N_13917,N_13179);
and U14157 (N_14157,N_13252,N_13782);
nor U14158 (N_14158,N_13641,N_13024);
and U14159 (N_14159,N_13698,N_13993);
xnor U14160 (N_14160,N_13692,N_13053);
or U14161 (N_14161,N_13164,N_13770);
nor U14162 (N_14162,N_13673,N_13535);
xor U14163 (N_14163,N_13073,N_13700);
xnor U14164 (N_14164,N_13129,N_13188);
nand U14165 (N_14165,N_13286,N_13584);
xnor U14166 (N_14166,N_13662,N_13359);
or U14167 (N_14167,N_13061,N_13609);
and U14168 (N_14168,N_13941,N_13765);
xor U14169 (N_14169,N_13276,N_13593);
or U14170 (N_14170,N_13623,N_13318);
and U14171 (N_14171,N_13183,N_13002);
and U14172 (N_14172,N_13900,N_13517);
or U14173 (N_14173,N_13100,N_13894);
nor U14174 (N_14174,N_13794,N_13011);
xor U14175 (N_14175,N_13718,N_13732);
nand U14176 (N_14176,N_13738,N_13175);
nor U14177 (N_14177,N_13695,N_13393);
nor U14178 (N_14178,N_13800,N_13141);
and U14179 (N_14179,N_13289,N_13567);
xor U14180 (N_14180,N_13558,N_13948);
or U14181 (N_14181,N_13167,N_13797);
and U14182 (N_14182,N_13005,N_13372);
and U14183 (N_14183,N_13126,N_13887);
or U14184 (N_14184,N_13460,N_13751);
nor U14185 (N_14185,N_13553,N_13343);
xor U14186 (N_14186,N_13324,N_13802);
and U14187 (N_14187,N_13906,N_13414);
nand U14188 (N_14188,N_13309,N_13099);
and U14189 (N_14189,N_13356,N_13405);
and U14190 (N_14190,N_13530,N_13911);
or U14191 (N_14191,N_13970,N_13461);
nor U14192 (N_14192,N_13817,N_13672);
or U14193 (N_14193,N_13353,N_13153);
nand U14194 (N_14194,N_13924,N_13209);
or U14195 (N_14195,N_13189,N_13086);
xor U14196 (N_14196,N_13684,N_13230);
nor U14197 (N_14197,N_13610,N_13699);
or U14198 (N_14198,N_13756,N_13867);
nand U14199 (N_14199,N_13639,N_13858);
xnor U14200 (N_14200,N_13846,N_13793);
and U14201 (N_14201,N_13395,N_13626);
or U14202 (N_14202,N_13651,N_13575);
or U14203 (N_14203,N_13959,N_13292);
and U14204 (N_14204,N_13422,N_13224);
nand U14205 (N_14205,N_13884,N_13810);
nor U14206 (N_14206,N_13151,N_13044);
nand U14207 (N_14207,N_13925,N_13420);
nor U14208 (N_14208,N_13772,N_13983);
nand U14209 (N_14209,N_13769,N_13541);
and U14210 (N_14210,N_13512,N_13449);
and U14211 (N_14211,N_13766,N_13403);
xnor U14212 (N_14212,N_13375,N_13358);
nor U14213 (N_14213,N_13445,N_13621);
nor U14214 (N_14214,N_13972,N_13455);
xnor U14215 (N_14215,N_13640,N_13476);
nand U14216 (N_14216,N_13037,N_13863);
or U14217 (N_14217,N_13186,N_13170);
nand U14218 (N_14218,N_13893,N_13520);
and U14219 (N_14219,N_13392,N_13466);
and U14220 (N_14220,N_13056,N_13440);
xnor U14221 (N_14221,N_13680,N_13123);
xnor U14222 (N_14222,N_13783,N_13506);
nand U14223 (N_14223,N_13212,N_13807);
xor U14224 (N_14224,N_13029,N_13537);
nor U14225 (N_14225,N_13132,N_13550);
and U14226 (N_14226,N_13979,N_13670);
nand U14227 (N_14227,N_13808,N_13731);
nand U14228 (N_14228,N_13346,N_13891);
nand U14229 (N_14229,N_13851,N_13328);
or U14230 (N_14230,N_13338,N_13201);
xor U14231 (N_14231,N_13274,N_13685);
xor U14232 (N_14232,N_13784,N_13190);
xor U14233 (N_14233,N_13873,N_13249);
nor U14234 (N_14234,N_13885,N_13206);
nor U14235 (N_14235,N_13435,N_13516);
nand U14236 (N_14236,N_13219,N_13147);
xnor U14237 (N_14237,N_13652,N_13601);
and U14238 (N_14238,N_13531,N_13984);
nor U14239 (N_14239,N_13092,N_13635);
or U14240 (N_14240,N_13638,N_13394);
nor U14241 (N_14241,N_13268,N_13529);
nor U14242 (N_14242,N_13850,N_13115);
nor U14243 (N_14243,N_13270,N_13250);
or U14244 (N_14244,N_13484,N_13622);
nor U14245 (N_14245,N_13244,N_13725);
xor U14246 (N_14246,N_13480,N_13400);
xnor U14247 (N_14247,N_13246,N_13967);
or U14248 (N_14248,N_13015,N_13226);
nor U14249 (N_14249,N_13384,N_13330);
nand U14250 (N_14250,N_13834,N_13830);
or U14251 (N_14251,N_13795,N_13743);
and U14252 (N_14252,N_13704,N_13585);
and U14253 (N_14253,N_13511,N_13299);
nor U14254 (N_14254,N_13798,N_13106);
and U14255 (N_14255,N_13238,N_13697);
xnor U14256 (N_14256,N_13077,N_13444);
nor U14257 (N_14257,N_13799,N_13524);
nor U14258 (N_14258,N_13963,N_13494);
and U14259 (N_14259,N_13388,N_13590);
or U14260 (N_14260,N_13145,N_13540);
nor U14261 (N_14261,N_13854,N_13723);
and U14262 (N_14262,N_13674,N_13690);
xnor U14263 (N_14263,N_13589,N_13227);
nor U14264 (N_14264,N_13960,N_13897);
nor U14265 (N_14265,N_13363,N_13304);
xor U14266 (N_14266,N_13805,N_13826);
xor U14267 (N_14267,N_13492,N_13331);
or U14268 (N_14268,N_13223,N_13952);
nand U14269 (N_14269,N_13426,N_13496);
nand U14270 (N_14270,N_13714,N_13839);
nor U14271 (N_14271,N_13755,N_13028);
and U14272 (N_14272,N_13221,N_13216);
nand U14273 (N_14273,N_13515,N_13758);
nor U14274 (N_14274,N_13764,N_13427);
nand U14275 (N_14275,N_13742,N_13592);
xor U14276 (N_14276,N_13386,N_13396);
xor U14277 (N_14277,N_13036,N_13089);
nand U14278 (N_14278,N_13646,N_13605);
and U14279 (N_14279,N_13442,N_13408);
nand U14280 (N_14280,N_13168,N_13578);
nor U14281 (N_14281,N_13165,N_13545);
or U14282 (N_14282,N_13010,N_13007);
and U14283 (N_14283,N_13896,N_13341);
nor U14284 (N_14284,N_13171,N_13803);
or U14285 (N_14285,N_13367,N_13148);
or U14286 (N_14286,N_13617,N_13869);
and U14287 (N_14287,N_13210,N_13125);
nand U14288 (N_14288,N_13822,N_13801);
nand U14289 (N_14289,N_13768,N_13551);
nor U14290 (N_14290,N_13247,N_13116);
xnor U14291 (N_14291,N_13097,N_13283);
xor U14292 (N_14292,N_13240,N_13907);
nor U14293 (N_14293,N_13901,N_13109);
nand U14294 (N_14294,N_13111,N_13717);
or U14295 (N_14295,N_13702,N_13075);
nand U14296 (N_14296,N_13481,N_13814);
or U14297 (N_14297,N_13204,N_13266);
and U14298 (N_14298,N_13316,N_13045);
xor U14299 (N_14299,N_13586,N_13404);
nand U14300 (N_14300,N_13648,N_13501);
nand U14301 (N_14301,N_13381,N_13205);
nor U14302 (N_14302,N_13746,N_13675);
xnor U14303 (N_14303,N_13470,N_13069);
xnor U14304 (N_14304,N_13929,N_13922);
nor U14305 (N_14305,N_13490,N_13306);
nor U14306 (N_14306,N_13729,N_13012);
or U14307 (N_14307,N_13842,N_13526);
nor U14308 (N_14308,N_13878,N_13880);
and U14309 (N_14309,N_13868,N_13267);
and U14310 (N_14310,N_13912,N_13402);
nand U14311 (N_14311,N_13043,N_13859);
and U14312 (N_14312,N_13001,N_13890);
xor U14313 (N_14313,N_13110,N_13080);
and U14314 (N_14314,N_13313,N_13786);
nor U14315 (N_14315,N_13262,N_13253);
nor U14316 (N_14316,N_13112,N_13750);
or U14317 (N_14317,N_13157,N_13532);
nor U14318 (N_14318,N_13745,N_13913);
nor U14319 (N_14319,N_13325,N_13344);
or U14320 (N_14320,N_13643,N_13491);
xor U14321 (N_14321,N_13181,N_13519);
or U14322 (N_14322,N_13727,N_13489);
or U14323 (N_14323,N_13067,N_13105);
nand U14324 (N_14324,N_13121,N_13459);
or U14325 (N_14325,N_13498,N_13006);
nand U14326 (N_14326,N_13620,N_13944);
xnor U14327 (N_14327,N_13196,N_13291);
xnor U14328 (N_14328,N_13796,N_13919);
nand U14329 (N_14329,N_13557,N_13774);
and U14330 (N_14330,N_13482,N_13477);
nand U14331 (N_14331,N_13809,N_13054);
or U14332 (N_14332,N_13055,N_13488);
or U14333 (N_14333,N_13728,N_13294);
xor U14334 (N_14334,N_13312,N_13841);
or U14335 (N_14335,N_13463,N_13581);
nor U14336 (N_14336,N_13957,N_13523);
and U14337 (N_14337,N_13347,N_13013);
xor U14338 (N_14338,N_13263,N_13256);
or U14339 (N_14339,N_13682,N_13421);
nand U14340 (N_14340,N_13174,N_13042);
and U14341 (N_14341,N_13579,N_13899);
or U14342 (N_14342,N_13285,N_13666);
nand U14343 (N_14343,N_13357,N_13951);
nand U14344 (N_14344,N_13398,N_13452);
xor U14345 (N_14345,N_13992,N_13789);
nand U14346 (N_14346,N_13914,N_13864);
or U14347 (N_14347,N_13497,N_13977);
or U14348 (N_14348,N_13088,N_13712);
and U14349 (N_14349,N_13133,N_13014);
nand U14350 (N_14350,N_13406,N_13504);
nor U14351 (N_14351,N_13365,N_13234);
and U14352 (N_14352,N_13272,N_13479);
nor U14353 (N_14353,N_13193,N_13462);
or U14354 (N_14354,N_13776,N_13198);
or U14355 (N_14355,N_13857,N_13668);
xnor U14356 (N_14356,N_13827,N_13048);
and U14357 (N_14357,N_13976,N_13327);
nor U14358 (N_14358,N_13938,N_13820);
nand U14359 (N_14359,N_13556,N_13374);
and U14360 (N_14360,N_13265,N_13665);
nand U14361 (N_14361,N_13342,N_13582);
nand U14362 (N_14362,N_13468,N_13762);
nor U14363 (N_14363,N_13211,N_13821);
nand U14364 (N_14364,N_13716,N_13791);
and U14365 (N_14365,N_13943,N_13450);
or U14366 (N_14366,N_13611,N_13988);
nand U14367 (N_14367,N_13185,N_13828);
xnor U14368 (N_14368,N_13065,N_13860);
nor U14369 (N_14369,N_13314,N_13999);
nor U14370 (N_14370,N_13471,N_13910);
nor U14371 (N_14371,N_13302,N_13040);
or U14372 (N_14372,N_13915,N_13505);
or U14373 (N_14373,N_13947,N_13631);
xnor U14374 (N_14374,N_13239,N_13499);
xnor U14375 (N_14375,N_13950,N_13453);
nor U14376 (N_14376,N_13870,N_13093);
and U14377 (N_14377,N_13559,N_13301);
nor U14378 (N_14378,N_13920,N_13371);
or U14379 (N_14379,N_13229,N_13131);
nor U14380 (N_14380,N_13233,N_13495);
nor U14381 (N_14381,N_13439,N_13865);
and U14382 (N_14382,N_13678,N_13875);
and U14383 (N_14383,N_13740,N_13599);
or U14384 (N_14384,N_13534,N_13721);
xor U14385 (N_14385,N_13548,N_13737);
or U14386 (N_14386,N_13295,N_13351);
and U14387 (N_14387,N_13613,N_13385);
or U14388 (N_14388,N_13994,N_13334);
nand U14389 (N_14389,N_13654,N_13208);
xor U14390 (N_14390,N_13242,N_13288);
nor U14391 (N_14391,N_13411,N_13604);
or U14392 (N_14392,N_13320,N_13836);
nor U14393 (N_14393,N_13619,N_13419);
and U14394 (N_14394,N_13119,N_13169);
nand U14395 (N_14395,N_13889,N_13866);
xor U14396 (N_14396,N_13407,N_13323);
and U14397 (N_14397,N_13031,N_13816);
xnor U14398 (N_14398,N_13023,N_13669);
nand U14399 (N_14399,N_13614,N_13724);
or U14400 (N_14400,N_13340,N_13397);
xor U14401 (N_14401,N_13997,N_13350);
nor U14402 (N_14402,N_13636,N_13364);
xor U14403 (N_14403,N_13264,N_13773);
xor U14404 (N_14404,N_13197,N_13102);
xor U14405 (N_14405,N_13536,N_13146);
nand U14406 (N_14406,N_13886,N_13222);
or U14407 (N_14407,N_13465,N_13856);
nand U14408 (N_14408,N_13416,N_13677);
or U14409 (N_14409,N_13502,N_13600);
or U14410 (N_14410,N_13975,N_13443);
or U14411 (N_14411,N_13493,N_13458);
or U14412 (N_14412,N_13653,N_13413);
nor U14413 (N_14413,N_13143,N_13130);
and U14414 (N_14414,N_13415,N_13849);
nand U14415 (N_14415,N_13980,N_13063);
or U14416 (N_14416,N_13564,N_13305);
xor U14417 (N_14417,N_13271,N_13969);
xnor U14418 (N_14418,N_13070,N_13333);
xor U14419 (N_14419,N_13300,N_13528);
nor U14420 (N_14420,N_13311,N_13835);
xor U14421 (N_14421,N_13905,N_13084);
or U14422 (N_14422,N_13290,N_13606);
and U14423 (N_14423,N_13081,N_13844);
and U14424 (N_14424,N_13335,N_13862);
nor U14425 (N_14425,N_13883,N_13904);
nand U14426 (N_14426,N_13019,N_13833);
xor U14427 (N_14427,N_13615,N_13260);
or U14428 (N_14428,N_13608,N_13852);
nand U14429 (N_14429,N_13380,N_13703);
xnor U14430 (N_14430,N_13881,N_13207);
or U14431 (N_14431,N_13898,N_13930);
and U14432 (N_14432,N_13966,N_13570);
nor U14433 (N_14433,N_13237,N_13594);
nand U14434 (N_14434,N_13928,N_13447);
or U14435 (N_14435,N_13225,N_13060);
nand U14436 (N_14436,N_13182,N_13149);
nand U14437 (N_14437,N_13689,N_13163);
or U14438 (N_14438,N_13108,N_13071);
nand U14439 (N_14439,N_13284,N_13332);
nand U14440 (N_14440,N_13741,N_13107);
and U14441 (N_14441,N_13257,N_13566);
nor U14442 (N_14442,N_13389,N_13804);
nand U14443 (N_14443,N_13676,N_13058);
nor U14444 (N_14444,N_13136,N_13008);
or U14445 (N_14445,N_13546,N_13747);
xor U14446 (N_14446,N_13187,N_13555);
and U14447 (N_14447,N_13172,N_13159);
and U14448 (N_14448,N_13079,N_13779);
nor U14449 (N_14449,N_13412,N_13383);
or U14450 (N_14450,N_13780,N_13932);
xnor U14451 (N_14451,N_13596,N_13457);
or U14452 (N_14452,N_13137,N_13939);
nor U14453 (N_14453,N_13050,N_13279);
and U14454 (N_14454,N_13763,N_13956);
xor U14455 (N_14455,N_13035,N_13418);
nand U14456 (N_14456,N_13767,N_13391);
nor U14457 (N_14457,N_13096,N_13473);
and U14458 (N_14458,N_13032,N_13739);
or U14459 (N_14459,N_13472,N_13361);
nor U14460 (N_14460,N_13158,N_13754);
nand U14461 (N_14461,N_13303,N_13142);
nor U14462 (N_14462,N_13708,N_13349);
nor U14463 (N_14463,N_13525,N_13275);
nor U14464 (N_14464,N_13832,N_13973);
nor U14465 (N_14465,N_13220,N_13927);
xnor U14466 (N_14466,N_13709,N_13781);
nand U14467 (N_14467,N_13513,N_13433);
nand U14468 (N_14468,N_13618,N_13771);
or U14469 (N_14469,N_13790,N_13308);
nand U14470 (N_14470,N_13722,N_13933);
nand U14471 (N_14471,N_13368,N_13278);
nor U14472 (N_14472,N_13379,N_13101);
nand U14473 (N_14473,N_13974,N_13194);
nor U14474 (N_14474,N_13177,N_13214);
nand U14475 (N_14475,N_13778,N_13908);
or U14476 (N_14476,N_13825,N_13228);
and U14477 (N_14477,N_13122,N_13681);
xor U14478 (N_14478,N_13561,N_13838);
and U14479 (N_14479,N_13326,N_13104);
nor U14480 (N_14480,N_13509,N_13761);
nor U14481 (N_14481,N_13437,N_13571);
nor U14482 (N_14482,N_13824,N_13628);
nand U14483 (N_14483,N_13282,N_13425);
or U14484 (N_14484,N_13542,N_13853);
nor U14485 (N_14485,N_13144,N_13390);
nand U14486 (N_14486,N_13777,N_13094);
or U14487 (N_14487,N_13522,N_13715);
xor U14488 (N_14488,N_13378,N_13377);
or U14489 (N_14489,N_13734,N_13813);
or U14490 (N_14490,N_13370,N_13978);
nand U14491 (N_14491,N_13310,N_13953);
nor U14492 (N_14492,N_13430,N_13591);
nand U14493 (N_14493,N_13281,N_13034);
nor U14494 (N_14494,N_13200,N_13062);
and U14495 (N_14495,N_13436,N_13355);
xor U14496 (N_14496,N_13694,N_13138);
or U14497 (N_14497,N_13843,N_13483);
or U14498 (N_14498,N_13352,N_13753);
and U14499 (N_14499,N_13203,N_13936);
and U14500 (N_14500,N_13783,N_13345);
nor U14501 (N_14501,N_13449,N_13387);
xor U14502 (N_14502,N_13355,N_13090);
nand U14503 (N_14503,N_13649,N_13247);
nor U14504 (N_14504,N_13121,N_13842);
or U14505 (N_14505,N_13245,N_13061);
or U14506 (N_14506,N_13258,N_13774);
and U14507 (N_14507,N_13337,N_13440);
nand U14508 (N_14508,N_13950,N_13750);
xnor U14509 (N_14509,N_13982,N_13294);
nor U14510 (N_14510,N_13288,N_13642);
and U14511 (N_14511,N_13125,N_13634);
nor U14512 (N_14512,N_13510,N_13143);
xnor U14513 (N_14513,N_13756,N_13281);
nor U14514 (N_14514,N_13235,N_13239);
xnor U14515 (N_14515,N_13550,N_13131);
nor U14516 (N_14516,N_13001,N_13546);
and U14517 (N_14517,N_13379,N_13902);
and U14518 (N_14518,N_13814,N_13062);
and U14519 (N_14519,N_13246,N_13780);
nand U14520 (N_14520,N_13096,N_13181);
xor U14521 (N_14521,N_13764,N_13531);
nor U14522 (N_14522,N_13645,N_13583);
or U14523 (N_14523,N_13526,N_13497);
xor U14524 (N_14524,N_13820,N_13173);
nand U14525 (N_14525,N_13528,N_13131);
nand U14526 (N_14526,N_13585,N_13258);
nor U14527 (N_14527,N_13864,N_13418);
nand U14528 (N_14528,N_13545,N_13472);
nand U14529 (N_14529,N_13968,N_13598);
xor U14530 (N_14530,N_13510,N_13012);
or U14531 (N_14531,N_13949,N_13764);
xnor U14532 (N_14532,N_13803,N_13696);
nor U14533 (N_14533,N_13280,N_13651);
or U14534 (N_14534,N_13168,N_13492);
nand U14535 (N_14535,N_13299,N_13682);
or U14536 (N_14536,N_13566,N_13111);
or U14537 (N_14537,N_13556,N_13346);
nor U14538 (N_14538,N_13468,N_13699);
nor U14539 (N_14539,N_13780,N_13243);
xor U14540 (N_14540,N_13437,N_13688);
or U14541 (N_14541,N_13624,N_13473);
and U14542 (N_14542,N_13160,N_13915);
nand U14543 (N_14543,N_13553,N_13236);
nand U14544 (N_14544,N_13422,N_13806);
nor U14545 (N_14545,N_13761,N_13678);
nor U14546 (N_14546,N_13644,N_13041);
xnor U14547 (N_14547,N_13360,N_13338);
and U14548 (N_14548,N_13147,N_13182);
and U14549 (N_14549,N_13978,N_13190);
xor U14550 (N_14550,N_13518,N_13511);
and U14551 (N_14551,N_13535,N_13630);
xor U14552 (N_14552,N_13569,N_13539);
xnor U14553 (N_14553,N_13769,N_13534);
nor U14554 (N_14554,N_13339,N_13763);
and U14555 (N_14555,N_13104,N_13577);
or U14556 (N_14556,N_13694,N_13827);
and U14557 (N_14557,N_13365,N_13671);
nand U14558 (N_14558,N_13966,N_13828);
or U14559 (N_14559,N_13492,N_13349);
xnor U14560 (N_14560,N_13599,N_13938);
nand U14561 (N_14561,N_13963,N_13618);
and U14562 (N_14562,N_13830,N_13237);
or U14563 (N_14563,N_13639,N_13242);
or U14564 (N_14564,N_13624,N_13545);
and U14565 (N_14565,N_13483,N_13756);
or U14566 (N_14566,N_13285,N_13152);
xor U14567 (N_14567,N_13164,N_13631);
and U14568 (N_14568,N_13708,N_13569);
and U14569 (N_14569,N_13432,N_13857);
nand U14570 (N_14570,N_13166,N_13459);
or U14571 (N_14571,N_13798,N_13800);
nor U14572 (N_14572,N_13330,N_13129);
xnor U14573 (N_14573,N_13095,N_13686);
nand U14574 (N_14574,N_13530,N_13961);
or U14575 (N_14575,N_13467,N_13417);
or U14576 (N_14576,N_13119,N_13587);
xor U14577 (N_14577,N_13088,N_13157);
xnor U14578 (N_14578,N_13354,N_13325);
nand U14579 (N_14579,N_13105,N_13987);
and U14580 (N_14580,N_13353,N_13252);
and U14581 (N_14581,N_13454,N_13916);
nand U14582 (N_14582,N_13456,N_13524);
and U14583 (N_14583,N_13543,N_13618);
xnor U14584 (N_14584,N_13602,N_13271);
nand U14585 (N_14585,N_13475,N_13893);
and U14586 (N_14586,N_13675,N_13031);
and U14587 (N_14587,N_13805,N_13603);
nand U14588 (N_14588,N_13537,N_13471);
and U14589 (N_14589,N_13574,N_13208);
nand U14590 (N_14590,N_13473,N_13579);
nor U14591 (N_14591,N_13709,N_13229);
xor U14592 (N_14592,N_13785,N_13015);
or U14593 (N_14593,N_13246,N_13752);
and U14594 (N_14594,N_13247,N_13381);
and U14595 (N_14595,N_13270,N_13253);
nand U14596 (N_14596,N_13245,N_13969);
xnor U14597 (N_14597,N_13753,N_13854);
nor U14598 (N_14598,N_13788,N_13216);
xnor U14599 (N_14599,N_13516,N_13982);
nand U14600 (N_14600,N_13706,N_13526);
or U14601 (N_14601,N_13915,N_13444);
nor U14602 (N_14602,N_13089,N_13457);
nor U14603 (N_14603,N_13345,N_13681);
nor U14604 (N_14604,N_13256,N_13594);
nor U14605 (N_14605,N_13654,N_13330);
nand U14606 (N_14606,N_13819,N_13514);
and U14607 (N_14607,N_13174,N_13632);
nor U14608 (N_14608,N_13879,N_13070);
or U14609 (N_14609,N_13877,N_13076);
and U14610 (N_14610,N_13260,N_13461);
nor U14611 (N_14611,N_13111,N_13858);
nand U14612 (N_14612,N_13851,N_13815);
nor U14613 (N_14613,N_13115,N_13327);
or U14614 (N_14614,N_13521,N_13780);
xor U14615 (N_14615,N_13433,N_13657);
nor U14616 (N_14616,N_13676,N_13489);
xnor U14617 (N_14617,N_13215,N_13172);
and U14618 (N_14618,N_13444,N_13206);
nor U14619 (N_14619,N_13691,N_13115);
nor U14620 (N_14620,N_13688,N_13645);
xnor U14621 (N_14621,N_13082,N_13652);
nand U14622 (N_14622,N_13091,N_13269);
xor U14623 (N_14623,N_13618,N_13792);
or U14624 (N_14624,N_13116,N_13417);
nand U14625 (N_14625,N_13868,N_13812);
nor U14626 (N_14626,N_13415,N_13293);
nor U14627 (N_14627,N_13910,N_13272);
or U14628 (N_14628,N_13836,N_13630);
nand U14629 (N_14629,N_13397,N_13833);
or U14630 (N_14630,N_13906,N_13128);
xor U14631 (N_14631,N_13365,N_13484);
xor U14632 (N_14632,N_13138,N_13902);
nor U14633 (N_14633,N_13092,N_13552);
and U14634 (N_14634,N_13792,N_13879);
or U14635 (N_14635,N_13068,N_13023);
and U14636 (N_14636,N_13732,N_13738);
nor U14637 (N_14637,N_13965,N_13962);
nor U14638 (N_14638,N_13285,N_13689);
nand U14639 (N_14639,N_13861,N_13664);
nor U14640 (N_14640,N_13339,N_13099);
or U14641 (N_14641,N_13633,N_13560);
nor U14642 (N_14642,N_13886,N_13771);
or U14643 (N_14643,N_13691,N_13199);
or U14644 (N_14644,N_13645,N_13167);
nand U14645 (N_14645,N_13637,N_13096);
and U14646 (N_14646,N_13812,N_13272);
or U14647 (N_14647,N_13919,N_13334);
nand U14648 (N_14648,N_13225,N_13886);
nand U14649 (N_14649,N_13190,N_13487);
nor U14650 (N_14650,N_13065,N_13938);
or U14651 (N_14651,N_13380,N_13965);
nand U14652 (N_14652,N_13921,N_13048);
nand U14653 (N_14653,N_13862,N_13430);
nor U14654 (N_14654,N_13748,N_13443);
nand U14655 (N_14655,N_13570,N_13707);
nand U14656 (N_14656,N_13270,N_13979);
nor U14657 (N_14657,N_13231,N_13733);
nand U14658 (N_14658,N_13827,N_13766);
and U14659 (N_14659,N_13133,N_13495);
and U14660 (N_14660,N_13259,N_13791);
nand U14661 (N_14661,N_13700,N_13203);
nand U14662 (N_14662,N_13086,N_13336);
or U14663 (N_14663,N_13219,N_13361);
or U14664 (N_14664,N_13286,N_13021);
or U14665 (N_14665,N_13252,N_13753);
nand U14666 (N_14666,N_13319,N_13964);
xnor U14667 (N_14667,N_13300,N_13476);
nor U14668 (N_14668,N_13678,N_13959);
and U14669 (N_14669,N_13872,N_13157);
and U14670 (N_14670,N_13986,N_13037);
nand U14671 (N_14671,N_13067,N_13308);
and U14672 (N_14672,N_13446,N_13659);
or U14673 (N_14673,N_13623,N_13036);
nor U14674 (N_14674,N_13401,N_13420);
nand U14675 (N_14675,N_13590,N_13392);
or U14676 (N_14676,N_13370,N_13259);
nand U14677 (N_14677,N_13883,N_13554);
and U14678 (N_14678,N_13315,N_13866);
xor U14679 (N_14679,N_13333,N_13818);
or U14680 (N_14680,N_13125,N_13105);
xnor U14681 (N_14681,N_13516,N_13680);
xnor U14682 (N_14682,N_13448,N_13338);
nor U14683 (N_14683,N_13003,N_13324);
or U14684 (N_14684,N_13832,N_13153);
or U14685 (N_14685,N_13784,N_13896);
xnor U14686 (N_14686,N_13822,N_13960);
nand U14687 (N_14687,N_13289,N_13505);
or U14688 (N_14688,N_13841,N_13033);
and U14689 (N_14689,N_13319,N_13685);
xnor U14690 (N_14690,N_13545,N_13171);
and U14691 (N_14691,N_13033,N_13241);
xnor U14692 (N_14692,N_13671,N_13186);
and U14693 (N_14693,N_13699,N_13455);
or U14694 (N_14694,N_13915,N_13510);
and U14695 (N_14695,N_13001,N_13570);
and U14696 (N_14696,N_13541,N_13034);
nand U14697 (N_14697,N_13099,N_13895);
nand U14698 (N_14698,N_13847,N_13749);
or U14699 (N_14699,N_13858,N_13745);
xor U14700 (N_14700,N_13065,N_13269);
nor U14701 (N_14701,N_13427,N_13748);
or U14702 (N_14702,N_13005,N_13334);
xnor U14703 (N_14703,N_13811,N_13341);
xor U14704 (N_14704,N_13541,N_13620);
or U14705 (N_14705,N_13911,N_13425);
nor U14706 (N_14706,N_13904,N_13528);
and U14707 (N_14707,N_13298,N_13131);
nand U14708 (N_14708,N_13997,N_13607);
and U14709 (N_14709,N_13302,N_13383);
or U14710 (N_14710,N_13354,N_13032);
or U14711 (N_14711,N_13612,N_13950);
xnor U14712 (N_14712,N_13197,N_13214);
and U14713 (N_14713,N_13409,N_13108);
nor U14714 (N_14714,N_13144,N_13694);
xor U14715 (N_14715,N_13618,N_13830);
nor U14716 (N_14716,N_13834,N_13148);
nor U14717 (N_14717,N_13265,N_13535);
xnor U14718 (N_14718,N_13471,N_13238);
nor U14719 (N_14719,N_13703,N_13350);
nand U14720 (N_14720,N_13013,N_13445);
nor U14721 (N_14721,N_13276,N_13590);
or U14722 (N_14722,N_13858,N_13448);
or U14723 (N_14723,N_13440,N_13772);
xor U14724 (N_14724,N_13135,N_13133);
nand U14725 (N_14725,N_13013,N_13509);
nor U14726 (N_14726,N_13933,N_13573);
xor U14727 (N_14727,N_13210,N_13015);
nor U14728 (N_14728,N_13610,N_13222);
and U14729 (N_14729,N_13168,N_13046);
and U14730 (N_14730,N_13287,N_13076);
and U14731 (N_14731,N_13413,N_13787);
nand U14732 (N_14732,N_13848,N_13734);
xor U14733 (N_14733,N_13285,N_13002);
xnor U14734 (N_14734,N_13429,N_13991);
xnor U14735 (N_14735,N_13923,N_13795);
and U14736 (N_14736,N_13094,N_13807);
xnor U14737 (N_14737,N_13925,N_13592);
nand U14738 (N_14738,N_13722,N_13165);
xnor U14739 (N_14739,N_13676,N_13513);
nor U14740 (N_14740,N_13838,N_13038);
or U14741 (N_14741,N_13551,N_13681);
and U14742 (N_14742,N_13678,N_13945);
nor U14743 (N_14743,N_13311,N_13083);
nand U14744 (N_14744,N_13480,N_13828);
and U14745 (N_14745,N_13183,N_13472);
nand U14746 (N_14746,N_13334,N_13445);
nand U14747 (N_14747,N_13462,N_13887);
xor U14748 (N_14748,N_13246,N_13675);
xnor U14749 (N_14749,N_13787,N_13647);
nor U14750 (N_14750,N_13497,N_13577);
nor U14751 (N_14751,N_13363,N_13896);
or U14752 (N_14752,N_13659,N_13100);
or U14753 (N_14753,N_13475,N_13677);
nor U14754 (N_14754,N_13617,N_13204);
and U14755 (N_14755,N_13872,N_13732);
nand U14756 (N_14756,N_13887,N_13951);
nand U14757 (N_14757,N_13962,N_13029);
or U14758 (N_14758,N_13731,N_13832);
nor U14759 (N_14759,N_13289,N_13944);
or U14760 (N_14760,N_13984,N_13513);
xnor U14761 (N_14761,N_13938,N_13660);
or U14762 (N_14762,N_13710,N_13724);
nand U14763 (N_14763,N_13630,N_13923);
or U14764 (N_14764,N_13436,N_13907);
nor U14765 (N_14765,N_13282,N_13116);
xnor U14766 (N_14766,N_13408,N_13122);
nor U14767 (N_14767,N_13987,N_13611);
and U14768 (N_14768,N_13872,N_13282);
or U14769 (N_14769,N_13185,N_13340);
or U14770 (N_14770,N_13470,N_13144);
or U14771 (N_14771,N_13678,N_13194);
or U14772 (N_14772,N_13956,N_13227);
nor U14773 (N_14773,N_13857,N_13353);
nor U14774 (N_14774,N_13362,N_13899);
nand U14775 (N_14775,N_13328,N_13890);
or U14776 (N_14776,N_13451,N_13365);
and U14777 (N_14777,N_13201,N_13737);
or U14778 (N_14778,N_13974,N_13473);
nor U14779 (N_14779,N_13110,N_13067);
or U14780 (N_14780,N_13824,N_13006);
xor U14781 (N_14781,N_13556,N_13533);
or U14782 (N_14782,N_13137,N_13019);
xnor U14783 (N_14783,N_13836,N_13433);
and U14784 (N_14784,N_13228,N_13465);
nor U14785 (N_14785,N_13018,N_13104);
or U14786 (N_14786,N_13223,N_13226);
nor U14787 (N_14787,N_13333,N_13289);
nand U14788 (N_14788,N_13813,N_13140);
nand U14789 (N_14789,N_13903,N_13401);
and U14790 (N_14790,N_13454,N_13908);
and U14791 (N_14791,N_13877,N_13352);
xor U14792 (N_14792,N_13498,N_13126);
and U14793 (N_14793,N_13612,N_13806);
nand U14794 (N_14794,N_13109,N_13609);
nand U14795 (N_14795,N_13347,N_13323);
or U14796 (N_14796,N_13281,N_13402);
xor U14797 (N_14797,N_13724,N_13140);
nand U14798 (N_14798,N_13694,N_13663);
nor U14799 (N_14799,N_13920,N_13394);
xnor U14800 (N_14800,N_13187,N_13004);
and U14801 (N_14801,N_13446,N_13800);
or U14802 (N_14802,N_13507,N_13604);
or U14803 (N_14803,N_13216,N_13354);
or U14804 (N_14804,N_13010,N_13126);
or U14805 (N_14805,N_13622,N_13150);
xor U14806 (N_14806,N_13307,N_13270);
nand U14807 (N_14807,N_13069,N_13873);
nor U14808 (N_14808,N_13939,N_13898);
or U14809 (N_14809,N_13874,N_13981);
xnor U14810 (N_14810,N_13413,N_13959);
or U14811 (N_14811,N_13897,N_13259);
nand U14812 (N_14812,N_13573,N_13894);
or U14813 (N_14813,N_13126,N_13678);
or U14814 (N_14814,N_13259,N_13419);
xor U14815 (N_14815,N_13041,N_13380);
xor U14816 (N_14816,N_13125,N_13065);
nor U14817 (N_14817,N_13873,N_13791);
and U14818 (N_14818,N_13130,N_13906);
and U14819 (N_14819,N_13472,N_13904);
and U14820 (N_14820,N_13299,N_13284);
and U14821 (N_14821,N_13676,N_13341);
nor U14822 (N_14822,N_13011,N_13114);
xor U14823 (N_14823,N_13095,N_13557);
and U14824 (N_14824,N_13706,N_13236);
xor U14825 (N_14825,N_13512,N_13072);
or U14826 (N_14826,N_13391,N_13433);
xor U14827 (N_14827,N_13301,N_13632);
xnor U14828 (N_14828,N_13128,N_13874);
nor U14829 (N_14829,N_13803,N_13890);
nor U14830 (N_14830,N_13835,N_13768);
or U14831 (N_14831,N_13868,N_13012);
xnor U14832 (N_14832,N_13408,N_13843);
nor U14833 (N_14833,N_13200,N_13093);
nand U14834 (N_14834,N_13683,N_13366);
nor U14835 (N_14835,N_13686,N_13662);
nand U14836 (N_14836,N_13213,N_13331);
xor U14837 (N_14837,N_13747,N_13462);
nor U14838 (N_14838,N_13444,N_13875);
nand U14839 (N_14839,N_13703,N_13004);
nor U14840 (N_14840,N_13548,N_13078);
and U14841 (N_14841,N_13877,N_13339);
xor U14842 (N_14842,N_13251,N_13082);
or U14843 (N_14843,N_13932,N_13735);
nor U14844 (N_14844,N_13107,N_13701);
and U14845 (N_14845,N_13283,N_13212);
or U14846 (N_14846,N_13358,N_13432);
nor U14847 (N_14847,N_13514,N_13499);
or U14848 (N_14848,N_13748,N_13481);
nor U14849 (N_14849,N_13257,N_13830);
or U14850 (N_14850,N_13217,N_13719);
nor U14851 (N_14851,N_13563,N_13081);
or U14852 (N_14852,N_13139,N_13230);
nor U14853 (N_14853,N_13223,N_13097);
or U14854 (N_14854,N_13482,N_13245);
nor U14855 (N_14855,N_13743,N_13281);
and U14856 (N_14856,N_13881,N_13841);
or U14857 (N_14857,N_13951,N_13762);
xnor U14858 (N_14858,N_13660,N_13476);
nand U14859 (N_14859,N_13427,N_13038);
nand U14860 (N_14860,N_13377,N_13960);
and U14861 (N_14861,N_13164,N_13515);
xor U14862 (N_14862,N_13445,N_13109);
and U14863 (N_14863,N_13983,N_13822);
and U14864 (N_14864,N_13357,N_13537);
and U14865 (N_14865,N_13224,N_13939);
nor U14866 (N_14866,N_13093,N_13204);
or U14867 (N_14867,N_13843,N_13773);
or U14868 (N_14868,N_13053,N_13947);
nor U14869 (N_14869,N_13868,N_13389);
or U14870 (N_14870,N_13009,N_13919);
or U14871 (N_14871,N_13640,N_13128);
xnor U14872 (N_14872,N_13061,N_13646);
and U14873 (N_14873,N_13921,N_13727);
nor U14874 (N_14874,N_13910,N_13433);
nand U14875 (N_14875,N_13498,N_13114);
and U14876 (N_14876,N_13767,N_13228);
nand U14877 (N_14877,N_13638,N_13615);
or U14878 (N_14878,N_13566,N_13485);
and U14879 (N_14879,N_13649,N_13810);
nand U14880 (N_14880,N_13990,N_13094);
and U14881 (N_14881,N_13435,N_13898);
or U14882 (N_14882,N_13867,N_13175);
nand U14883 (N_14883,N_13714,N_13569);
nor U14884 (N_14884,N_13237,N_13197);
xor U14885 (N_14885,N_13188,N_13370);
or U14886 (N_14886,N_13435,N_13971);
and U14887 (N_14887,N_13515,N_13580);
xor U14888 (N_14888,N_13591,N_13033);
nor U14889 (N_14889,N_13184,N_13363);
nand U14890 (N_14890,N_13680,N_13683);
xnor U14891 (N_14891,N_13710,N_13236);
nand U14892 (N_14892,N_13713,N_13343);
nor U14893 (N_14893,N_13024,N_13005);
nor U14894 (N_14894,N_13969,N_13793);
or U14895 (N_14895,N_13699,N_13369);
nand U14896 (N_14896,N_13810,N_13295);
or U14897 (N_14897,N_13971,N_13583);
or U14898 (N_14898,N_13259,N_13069);
xnor U14899 (N_14899,N_13596,N_13370);
or U14900 (N_14900,N_13304,N_13334);
nand U14901 (N_14901,N_13372,N_13349);
and U14902 (N_14902,N_13751,N_13139);
or U14903 (N_14903,N_13621,N_13973);
and U14904 (N_14904,N_13602,N_13706);
nor U14905 (N_14905,N_13798,N_13721);
nand U14906 (N_14906,N_13512,N_13727);
or U14907 (N_14907,N_13802,N_13916);
and U14908 (N_14908,N_13630,N_13048);
and U14909 (N_14909,N_13453,N_13426);
and U14910 (N_14910,N_13754,N_13547);
xor U14911 (N_14911,N_13156,N_13259);
and U14912 (N_14912,N_13129,N_13208);
or U14913 (N_14913,N_13427,N_13883);
nand U14914 (N_14914,N_13092,N_13211);
nand U14915 (N_14915,N_13977,N_13709);
nand U14916 (N_14916,N_13960,N_13188);
nor U14917 (N_14917,N_13200,N_13897);
nor U14918 (N_14918,N_13332,N_13181);
xnor U14919 (N_14919,N_13319,N_13765);
or U14920 (N_14920,N_13859,N_13255);
or U14921 (N_14921,N_13787,N_13985);
nor U14922 (N_14922,N_13741,N_13045);
nor U14923 (N_14923,N_13040,N_13108);
xnor U14924 (N_14924,N_13378,N_13348);
and U14925 (N_14925,N_13463,N_13722);
or U14926 (N_14926,N_13203,N_13145);
xnor U14927 (N_14927,N_13140,N_13126);
nor U14928 (N_14928,N_13977,N_13840);
or U14929 (N_14929,N_13179,N_13352);
and U14930 (N_14930,N_13680,N_13083);
nor U14931 (N_14931,N_13601,N_13907);
xor U14932 (N_14932,N_13681,N_13615);
nor U14933 (N_14933,N_13797,N_13048);
nor U14934 (N_14934,N_13088,N_13295);
xor U14935 (N_14935,N_13659,N_13708);
nand U14936 (N_14936,N_13263,N_13858);
nand U14937 (N_14937,N_13275,N_13172);
and U14938 (N_14938,N_13020,N_13918);
or U14939 (N_14939,N_13572,N_13760);
nand U14940 (N_14940,N_13503,N_13738);
and U14941 (N_14941,N_13068,N_13650);
xnor U14942 (N_14942,N_13420,N_13922);
nand U14943 (N_14943,N_13492,N_13023);
nor U14944 (N_14944,N_13441,N_13387);
xor U14945 (N_14945,N_13096,N_13686);
nand U14946 (N_14946,N_13151,N_13340);
xor U14947 (N_14947,N_13232,N_13422);
nor U14948 (N_14948,N_13593,N_13138);
nor U14949 (N_14949,N_13591,N_13289);
or U14950 (N_14950,N_13748,N_13886);
xor U14951 (N_14951,N_13802,N_13669);
and U14952 (N_14952,N_13610,N_13445);
nor U14953 (N_14953,N_13713,N_13031);
nor U14954 (N_14954,N_13401,N_13253);
or U14955 (N_14955,N_13352,N_13568);
xnor U14956 (N_14956,N_13233,N_13003);
and U14957 (N_14957,N_13909,N_13441);
xor U14958 (N_14958,N_13980,N_13818);
nor U14959 (N_14959,N_13744,N_13687);
or U14960 (N_14960,N_13439,N_13578);
nand U14961 (N_14961,N_13648,N_13937);
or U14962 (N_14962,N_13927,N_13174);
xnor U14963 (N_14963,N_13091,N_13785);
xnor U14964 (N_14964,N_13795,N_13304);
xnor U14965 (N_14965,N_13024,N_13980);
nand U14966 (N_14966,N_13738,N_13071);
and U14967 (N_14967,N_13077,N_13103);
nand U14968 (N_14968,N_13964,N_13761);
or U14969 (N_14969,N_13102,N_13239);
nand U14970 (N_14970,N_13160,N_13347);
nor U14971 (N_14971,N_13793,N_13856);
nand U14972 (N_14972,N_13257,N_13331);
nor U14973 (N_14973,N_13450,N_13860);
or U14974 (N_14974,N_13344,N_13639);
and U14975 (N_14975,N_13898,N_13382);
nand U14976 (N_14976,N_13134,N_13462);
or U14977 (N_14977,N_13517,N_13238);
and U14978 (N_14978,N_13553,N_13361);
xnor U14979 (N_14979,N_13243,N_13675);
nand U14980 (N_14980,N_13322,N_13673);
or U14981 (N_14981,N_13286,N_13984);
nand U14982 (N_14982,N_13883,N_13453);
or U14983 (N_14983,N_13501,N_13202);
xnor U14984 (N_14984,N_13126,N_13905);
nor U14985 (N_14985,N_13345,N_13984);
nor U14986 (N_14986,N_13147,N_13455);
or U14987 (N_14987,N_13334,N_13389);
nand U14988 (N_14988,N_13841,N_13450);
and U14989 (N_14989,N_13554,N_13956);
nand U14990 (N_14990,N_13129,N_13605);
nand U14991 (N_14991,N_13495,N_13045);
xor U14992 (N_14992,N_13661,N_13880);
xnor U14993 (N_14993,N_13078,N_13092);
xor U14994 (N_14994,N_13430,N_13811);
or U14995 (N_14995,N_13930,N_13653);
xor U14996 (N_14996,N_13098,N_13853);
or U14997 (N_14997,N_13238,N_13352);
or U14998 (N_14998,N_13678,N_13112);
nand U14999 (N_14999,N_13581,N_13337);
nand U15000 (N_15000,N_14525,N_14283);
nor U15001 (N_15001,N_14929,N_14098);
nor U15002 (N_15002,N_14248,N_14056);
nand U15003 (N_15003,N_14013,N_14369);
xnor U15004 (N_15004,N_14635,N_14552);
nand U15005 (N_15005,N_14387,N_14923);
nor U15006 (N_15006,N_14993,N_14595);
nand U15007 (N_15007,N_14408,N_14543);
and U15008 (N_15008,N_14023,N_14512);
and U15009 (N_15009,N_14809,N_14094);
and U15010 (N_15010,N_14535,N_14076);
or U15011 (N_15011,N_14955,N_14601);
nor U15012 (N_15012,N_14950,N_14902);
and U15013 (N_15013,N_14703,N_14747);
xnor U15014 (N_15014,N_14879,N_14174);
nor U15015 (N_15015,N_14011,N_14469);
or U15016 (N_15016,N_14611,N_14969);
nor U15017 (N_15017,N_14700,N_14613);
or U15018 (N_15018,N_14072,N_14466);
xor U15019 (N_15019,N_14158,N_14890);
nand U15020 (N_15020,N_14610,N_14351);
xnor U15021 (N_15021,N_14041,N_14003);
xor U15022 (N_15022,N_14465,N_14200);
nand U15023 (N_15023,N_14160,N_14756);
nor U15024 (N_15024,N_14165,N_14529);
nand U15025 (N_15025,N_14889,N_14823);
and U15026 (N_15026,N_14623,N_14679);
xor U15027 (N_15027,N_14268,N_14640);
xnor U15028 (N_15028,N_14990,N_14253);
xor U15029 (N_15029,N_14767,N_14453);
xor U15030 (N_15030,N_14571,N_14524);
nor U15031 (N_15031,N_14562,N_14522);
nand U15032 (N_15032,N_14191,N_14102);
xnor U15033 (N_15033,N_14356,N_14954);
or U15034 (N_15034,N_14557,N_14170);
or U15035 (N_15035,N_14006,N_14898);
nand U15036 (N_15036,N_14289,N_14398);
xnor U15037 (N_15037,N_14667,N_14963);
xor U15038 (N_15038,N_14657,N_14718);
or U15039 (N_15039,N_14149,N_14295);
and U15040 (N_15040,N_14516,N_14928);
and U15041 (N_15041,N_14821,N_14900);
xnor U15042 (N_15042,N_14340,N_14674);
and U15043 (N_15043,N_14213,N_14171);
nor U15044 (N_15044,N_14463,N_14561);
nor U15045 (N_15045,N_14989,N_14856);
or U15046 (N_15046,N_14329,N_14089);
xor U15047 (N_15047,N_14447,N_14456);
nor U15048 (N_15048,N_14786,N_14723);
or U15049 (N_15049,N_14096,N_14620);
or U15050 (N_15050,N_14942,N_14047);
xnor U15051 (N_15051,N_14816,N_14793);
nor U15052 (N_15052,N_14842,N_14943);
or U15053 (N_15053,N_14684,N_14261);
nand U15054 (N_15054,N_14488,N_14251);
xnor U15055 (N_15055,N_14282,N_14030);
nand U15056 (N_15056,N_14332,N_14903);
nor U15057 (N_15057,N_14231,N_14361);
nor U15058 (N_15058,N_14537,N_14281);
and U15059 (N_15059,N_14000,N_14145);
xor U15060 (N_15060,N_14059,N_14719);
nand U15061 (N_15061,N_14214,N_14300);
nor U15062 (N_15062,N_14685,N_14808);
nor U15063 (N_15063,N_14945,N_14227);
or U15064 (N_15064,N_14142,N_14125);
or U15065 (N_15065,N_14711,N_14585);
xor U15066 (N_15066,N_14492,N_14454);
nand U15067 (N_15067,N_14401,N_14947);
xnor U15068 (N_15068,N_14185,N_14377);
nor U15069 (N_15069,N_14830,N_14549);
or U15070 (N_15070,N_14598,N_14020);
xnor U15071 (N_15071,N_14441,N_14275);
nand U15072 (N_15072,N_14981,N_14479);
nand U15073 (N_15073,N_14655,N_14960);
nor U15074 (N_15074,N_14997,N_14068);
xor U15075 (N_15075,N_14860,N_14314);
or U15076 (N_15076,N_14720,N_14690);
nor U15077 (N_15077,N_14825,N_14473);
nor U15078 (N_15078,N_14426,N_14504);
or U15079 (N_15079,N_14192,N_14725);
nand U15080 (N_15080,N_14163,N_14382);
or U15081 (N_15081,N_14858,N_14226);
nand U15082 (N_15082,N_14877,N_14910);
nand U15083 (N_15083,N_14977,N_14153);
or U15084 (N_15084,N_14864,N_14166);
and U15085 (N_15085,N_14276,N_14054);
nand U15086 (N_15086,N_14882,N_14381);
and U15087 (N_15087,N_14603,N_14859);
nand U15088 (N_15088,N_14616,N_14560);
or U15089 (N_15089,N_14622,N_14052);
xnor U15090 (N_15090,N_14451,N_14578);
or U15091 (N_15091,N_14907,N_14061);
and U15092 (N_15092,N_14057,N_14067);
or U15093 (N_15093,N_14333,N_14090);
and U15094 (N_15094,N_14671,N_14895);
nand U15095 (N_15095,N_14146,N_14007);
nand U15096 (N_15096,N_14217,N_14548);
nand U15097 (N_15097,N_14505,N_14404);
and U15098 (N_15098,N_14687,N_14341);
or U15099 (N_15099,N_14273,N_14737);
and U15100 (N_15100,N_14254,N_14366);
or U15101 (N_15101,N_14748,N_14405);
nor U15102 (N_15102,N_14932,N_14117);
and U15103 (N_15103,N_14209,N_14501);
and U15104 (N_15104,N_14223,N_14956);
and U15105 (N_15105,N_14834,N_14316);
nand U15106 (N_15106,N_14123,N_14312);
nor U15107 (N_15107,N_14712,N_14503);
nand U15108 (N_15108,N_14139,N_14857);
and U15109 (N_15109,N_14471,N_14869);
or U15110 (N_15110,N_14544,N_14205);
and U15111 (N_15111,N_14033,N_14754);
and U15112 (N_15112,N_14347,N_14461);
nand U15113 (N_15113,N_14490,N_14964);
xnor U15114 (N_15114,N_14713,N_14063);
and U15115 (N_15115,N_14403,N_14339);
and U15116 (N_15116,N_14978,N_14733);
nand U15117 (N_15117,N_14394,N_14155);
xnor U15118 (N_15118,N_14257,N_14681);
or U15119 (N_15119,N_14129,N_14293);
and U15120 (N_15120,N_14468,N_14927);
and U15121 (N_15121,N_14818,N_14965);
and U15122 (N_15122,N_14497,N_14573);
or U15123 (N_15123,N_14495,N_14175);
xnor U15124 (N_15124,N_14088,N_14766);
and U15125 (N_15125,N_14764,N_14176);
nand U15126 (N_15126,N_14844,N_14705);
or U15127 (N_15127,N_14092,N_14122);
xor U15128 (N_15128,N_14986,N_14106);
and U15129 (N_15129,N_14034,N_14686);
or U15130 (N_15130,N_14082,N_14435);
and U15131 (N_15131,N_14198,N_14169);
or U15132 (N_15132,N_14788,N_14630);
and U15133 (N_15133,N_14768,N_14364);
or U15134 (N_15134,N_14936,N_14527);
or U15135 (N_15135,N_14514,N_14645);
nor U15136 (N_15136,N_14915,N_14948);
and U15137 (N_15137,N_14589,N_14644);
or U15138 (N_15138,N_14670,N_14776);
nand U15139 (N_15139,N_14855,N_14588);
and U15140 (N_15140,N_14049,N_14559);
and U15141 (N_15141,N_14846,N_14672);
xnor U15142 (N_15142,N_14500,N_14836);
xor U15143 (N_15143,N_14162,N_14320);
nor U15144 (N_15144,N_14722,N_14147);
or U15145 (N_15145,N_14246,N_14968);
and U15146 (N_15146,N_14012,N_14868);
and U15147 (N_15147,N_14288,N_14753);
and U15148 (N_15148,N_14309,N_14563);
and U15149 (N_15149,N_14400,N_14941);
and U15150 (N_15150,N_14570,N_14871);
xnor U15151 (N_15151,N_14653,N_14569);
and U15152 (N_15152,N_14091,N_14532);
or U15153 (N_15153,N_14621,N_14840);
and U15154 (N_15154,N_14474,N_14373);
nor U15155 (N_15155,N_14513,N_14795);
nand U15156 (N_15156,N_14799,N_14673);
and U15157 (N_15157,N_14342,N_14785);
nand U15158 (N_15158,N_14521,N_14368);
or U15159 (N_15159,N_14779,N_14999);
nand U15160 (N_15160,N_14913,N_14971);
or U15161 (N_15161,N_14104,N_14380);
xnor U15162 (N_15162,N_14250,N_14609);
nand U15163 (N_15163,N_14832,N_14229);
or U15164 (N_15164,N_14996,N_14040);
or U15165 (N_15165,N_14010,N_14534);
nand U15166 (N_15166,N_14695,N_14113);
nand U15167 (N_15167,N_14424,N_14930);
xnor U15168 (N_15168,N_14439,N_14038);
nand U15169 (N_15169,N_14310,N_14597);
xor U15170 (N_15170,N_14908,N_14749);
nand U15171 (N_15171,N_14888,N_14416);
and U15172 (N_15172,N_14498,N_14018);
nand U15173 (N_15173,N_14899,N_14920);
nand U15174 (N_15174,N_14724,N_14266);
xor U15175 (N_15175,N_14262,N_14843);
nor U15176 (N_15176,N_14014,N_14952);
xor U15177 (N_15177,N_14388,N_14304);
and U15178 (N_15178,N_14225,N_14957);
and U15179 (N_15179,N_14233,N_14350);
nand U15180 (N_15180,N_14193,N_14692);
nor U15181 (N_15181,N_14547,N_14390);
or U15182 (N_15182,N_14208,N_14420);
and U15183 (N_15183,N_14070,N_14272);
nor U15184 (N_15184,N_14639,N_14376);
and U15185 (N_15185,N_14087,N_14448);
nand U15186 (N_15186,N_14182,N_14274);
nor U15187 (N_15187,N_14873,N_14241);
nor U15188 (N_15188,N_14105,N_14084);
or U15189 (N_15189,N_14696,N_14704);
and U15190 (N_15190,N_14140,N_14240);
nor U15191 (N_15191,N_14650,N_14277);
and U15192 (N_15192,N_14717,N_14103);
nand U15193 (N_15193,N_14729,N_14884);
or U15194 (N_15194,N_14829,N_14750);
nor U15195 (N_15195,N_14736,N_14446);
and U15196 (N_15196,N_14666,N_14502);
xnor U15197 (N_15197,N_14581,N_14156);
xor U15198 (N_15198,N_14083,N_14702);
nor U15199 (N_15199,N_14852,N_14554);
xor U15200 (N_15200,N_14551,N_14530);
nand U15201 (N_15201,N_14385,N_14462);
nor U15202 (N_15202,N_14819,N_14677);
xor U15203 (N_15203,N_14894,N_14431);
and U15204 (N_15204,N_14983,N_14697);
and U15205 (N_15205,N_14693,N_14769);
and U15206 (N_15206,N_14837,N_14402);
nor U15207 (N_15207,N_14592,N_14797);
nand U15208 (N_15208,N_14510,N_14450);
or U15209 (N_15209,N_14574,N_14780);
and U15210 (N_15210,N_14337,N_14976);
nand U15211 (N_15211,N_14567,N_14912);
or U15212 (N_15212,N_14520,N_14765);
nand U15213 (N_15213,N_14746,N_14699);
or U15214 (N_15214,N_14953,N_14949);
and U15215 (N_15215,N_14594,N_14706);
nand U15216 (N_15216,N_14331,N_14303);
nand U15217 (N_15217,N_14016,N_14614);
nand U15218 (N_15218,N_14157,N_14599);
or U15219 (N_15219,N_14627,N_14414);
xor U15220 (N_15220,N_14099,N_14833);
nand U15221 (N_15221,N_14258,N_14338);
xor U15222 (N_15222,N_14798,N_14587);
nor U15223 (N_15223,N_14961,N_14045);
nand U15224 (N_15224,N_14878,N_14035);
nor U15225 (N_15225,N_14349,N_14861);
nor U15226 (N_15226,N_14423,N_14847);
xor U15227 (N_15227,N_14773,N_14159);
xor U15228 (N_15228,N_14352,N_14234);
or U15229 (N_15229,N_14641,N_14443);
xor U15230 (N_15230,N_14606,N_14874);
nand U15231 (N_15231,N_14896,N_14178);
nand U15232 (N_15232,N_14714,N_14464);
xor U15233 (N_15233,N_14814,N_14663);
nor U15234 (N_15234,N_14384,N_14519);
xnor U15235 (N_15235,N_14154,N_14112);
xor U15236 (N_15236,N_14228,N_14039);
nor U15237 (N_15237,N_14716,N_14991);
or U15238 (N_15238,N_14583,N_14726);
xnor U15239 (N_15239,N_14743,N_14985);
and U15240 (N_15240,N_14301,N_14467);
xor U15241 (N_15241,N_14807,N_14883);
or U15242 (N_15242,N_14988,N_14212);
and U15243 (N_15243,N_14710,N_14811);
nand U15244 (N_15244,N_14238,N_14418);
nand U15245 (N_15245,N_14410,N_14186);
xor U15246 (N_15246,N_14744,N_14181);
nor U15247 (N_15247,N_14741,N_14161);
and U15248 (N_15248,N_14870,N_14546);
nor U15249 (N_15249,N_14242,N_14457);
nand U15250 (N_15250,N_14375,N_14688);
and U15251 (N_15251,N_14066,N_14108);
xnor U15252 (N_15252,N_14781,N_14515);
and U15253 (N_15253,N_14021,N_14721);
nand U15254 (N_15254,N_14399,N_14862);
or U15255 (N_15255,N_14101,N_14239);
or U15256 (N_15256,N_14334,N_14081);
nand U15257 (N_15257,N_14701,N_14572);
and U15258 (N_15258,N_14211,N_14069);
and U15259 (N_15259,N_14917,N_14493);
xnor U15260 (N_15260,N_14576,N_14734);
xor U15261 (N_15261,N_14951,N_14188);
nand U15262 (N_15262,N_14762,N_14732);
xor U15263 (N_15263,N_14236,N_14370);
nor U15264 (N_15264,N_14187,N_14132);
nand U15265 (N_15265,N_14220,N_14805);
and U15266 (N_15266,N_14128,N_14680);
xnor U15267 (N_15267,N_14260,N_14801);
nand U15268 (N_15268,N_14026,N_14249);
nor U15269 (N_15269,N_14100,N_14566);
nor U15270 (N_15270,N_14015,N_14302);
and U15271 (N_15271,N_14817,N_14053);
or U15272 (N_15272,N_14201,N_14343);
or U15273 (N_15273,N_14517,N_14429);
nand U15274 (N_15274,N_14914,N_14319);
or U15275 (N_15275,N_14586,N_14777);
or U15276 (N_15276,N_14458,N_14642);
and U15277 (N_15277,N_14631,N_14851);
or U15278 (N_15278,N_14810,N_14675);
and U15279 (N_15279,N_14298,N_14555);
nand U15280 (N_15280,N_14255,N_14327);
nand U15281 (N_15281,N_14742,N_14848);
xor U15282 (N_15282,N_14050,N_14784);
and U15283 (N_15283,N_14865,N_14975);
and U15284 (N_15284,N_14982,N_14481);
and U15285 (N_15285,N_14728,N_14305);
and U15286 (N_15286,N_14905,N_14958);
xnor U15287 (N_15287,N_14796,N_14152);
nand U15288 (N_15288,N_14425,N_14531);
nor U15289 (N_15289,N_14126,N_14218);
and U15290 (N_15290,N_14691,N_14173);
and U15291 (N_15291,N_14523,N_14660);
nand U15292 (N_15292,N_14665,N_14017);
xnor U15293 (N_15293,N_14179,N_14538);
nor U15294 (N_15294,N_14646,N_14036);
nand U15295 (N_15295,N_14417,N_14078);
xnor U15296 (N_15296,N_14540,N_14134);
xnor U15297 (N_15297,N_14872,N_14137);
and U15298 (N_15298,N_14393,N_14564);
and U15299 (N_15299,N_14438,N_14037);
nand U15300 (N_15300,N_14863,N_14921);
nand U15301 (N_15301,N_14328,N_14542);
and U15302 (N_15302,N_14919,N_14866);
nor U15303 (N_15303,N_14051,N_14323);
nand U15304 (N_15304,N_14783,N_14436);
nor U15305 (N_15305,N_14636,N_14355);
and U15306 (N_15306,N_14664,N_14189);
and U15307 (N_15307,N_14372,N_14415);
or U15308 (N_15308,N_14483,N_14841);
or U15309 (N_15309,N_14709,N_14306);
and U15310 (N_15310,N_14144,N_14354);
or U15311 (N_15311,N_14259,N_14615);
or U15312 (N_15312,N_14299,N_14730);
or U15313 (N_15313,N_14321,N_14740);
and U15314 (N_15314,N_14118,N_14264);
nand U15315 (N_15315,N_14835,N_14934);
or U15316 (N_15316,N_14926,N_14203);
or U15317 (N_15317,N_14210,N_14389);
nor U15318 (N_15318,N_14545,N_14489);
or U15319 (N_15319,N_14318,N_14267);
nor U15320 (N_15320,N_14419,N_14669);
xor U15321 (N_15321,N_14838,N_14433);
nand U15322 (N_15322,N_14933,N_14484);
nor U15323 (N_15323,N_14694,N_14031);
nor U15324 (N_15324,N_14880,N_14107);
or U15325 (N_15325,N_14120,N_14345);
or U15326 (N_15326,N_14245,N_14138);
nand U15327 (N_15327,N_14628,N_14661);
nand U15328 (N_15328,N_14715,N_14449);
nor U15329 (N_15329,N_14284,N_14886);
xor U15330 (N_15330,N_14761,N_14875);
or U15331 (N_15331,N_14649,N_14792);
xor U15332 (N_15332,N_14075,N_14853);
nor U15333 (N_15333,N_14850,N_14682);
xor U15334 (N_15334,N_14891,N_14541);
nand U15335 (N_15335,N_14656,N_14618);
nor U15336 (N_15336,N_14658,N_14365);
and U15337 (N_15337,N_14800,N_14787);
nand U15338 (N_15338,N_14279,N_14028);
or U15339 (N_15339,N_14499,N_14042);
or U15340 (N_15340,N_14358,N_14317);
or U15341 (N_15341,N_14487,N_14190);
xor U15342 (N_15342,N_14931,N_14475);
and U15343 (N_15343,N_14591,N_14739);
and U15344 (N_15344,N_14803,N_14826);
nor U15345 (N_15345,N_14348,N_14791);
nand U15346 (N_15346,N_14604,N_14839);
and U15347 (N_15347,N_14378,N_14244);
nand U15348 (N_15348,N_14772,N_14593);
or U15349 (N_15349,N_14285,N_14206);
nor U15350 (N_15350,N_14197,N_14392);
nand U15351 (N_15351,N_14172,N_14528);
or U15352 (N_15352,N_14130,N_14918);
or U15353 (N_15353,N_14216,N_14533);
and U15354 (N_15354,N_14442,N_14944);
xnor U15355 (N_15355,N_14617,N_14526);
or U15356 (N_15356,N_14782,N_14110);
nand U15357 (N_15357,N_14291,N_14055);
or U15358 (N_15358,N_14980,N_14270);
or U15359 (N_15359,N_14353,N_14491);
and U15360 (N_15360,N_14536,N_14071);
nor U15361 (N_15361,N_14459,N_14127);
xor U15362 (N_15362,N_14287,N_14252);
xor U15363 (N_15363,N_14608,N_14095);
nand U15364 (N_15364,N_14897,N_14150);
or U15365 (N_15365,N_14979,N_14177);
nor U15366 (N_15366,N_14024,N_14432);
nand U15367 (N_15367,N_14079,N_14738);
nor U15368 (N_15368,N_14962,N_14938);
nor U15369 (N_15369,N_14984,N_14445);
or U15370 (N_15370,N_14064,N_14815);
or U15371 (N_15371,N_14472,N_14428);
nor U15372 (N_15372,N_14427,N_14727);
nor U15373 (N_15373,N_14001,N_14025);
nand U15374 (N_15374,N_14085,N_14643);
and U15375 (N_15375,N_14027,N_14794);
nor U15376 (N_15376,N_14115,N_14970);
nand U15377 (N_15377,N_14676,N_14440);
xor U15378 (N_15378,N_14396,N_14509);
or U15379 (N_15379,N_14887,N_14019);
nor U15380 (N_15380,N_14151,N_14731);
and U15381 (N_15381,N_14297,N_14974);
xnor U15382 (N_15382,N_14596,N_14575);
nand U15383 (N_15383,N_14906,N_14619);
or U15384 (N_15384,N_14383,N_14924);
or U15385 (N_15385,N_14386,N_14959);
nand U15386 (N_15386,N_14632,N_14046);
nand U15387 (N_15387,N_14987,N_14232);
and U15388 (N_15388,N_14397,N_14651);
and U15389 (N_15389,N_14496,N_14080);
and U15390 (N_15390,N_14757,N_14995);
nor U15391 (N_15391,N_14922,N_14998);
nor U15392 (N_15392,N_14135,N_14494);
and U15393 (N_15393,N_14476,N_14195);
xor U15394 (N_15394,N_14395,N_14939);
and U15395 (N_15395,N_14235,N_14607);
xnor U15396 (N_15396,N_14760,N_14256);
nor U15397 (N_15397,N_14265,N_14478);
or U15398 (N_15398,N_14972,N_14048);
and U15399 (N_15399,N_14452,N_14633);
or U15400 (N_15400,N_14335,N_14827);
nor U15401 (N_15401,N_14849,N_14344);
nand U15402 (N_15402,N_14029,N_14164);
nand U15403 (N_15403,N_14243,N_14371);
or U15404 (N_15404,N_14937,N_14925);
nor U15405 (N_15405,N_14324,N_14707);
and U15406 (N_15406,N_14828,N_14508);
or U15407 (N_15407,N_14477,N_14168);
nand U15408 (N_15408,N_14708,N_14148);
or U15409 (N_15409,N_14579,N_14820);
nor U15410 (N_15410,N_14434,N_14745);
xor U15411 (N_15411,N_14752,N_14539);
nor U15412 (N_15412,N_14577,N_14946);
and U15413 (N_15413,N_14136,N_14876);
xnor U15414 (N_15414,N_14916,N_14359);
nand U15415 (N_15415,N_14698,N_14652);
and U15416 (N_15416,N_14507,N_14221);
nand U15417 (N_15417,N_14065,N_14867);
nand U15418 (N_15418,N_14582,N_14360);
nor U15419 (N_15419,N_14062,N_14437);
nor U15420 (N_15420,N_14271,N_14294);
nor U15421 (N_15421,N_14689,N_14812);
and U15422 (N_15422,N_14824,N_14480);
nor U15423 (N_15423,N_14612,N_14940);
and U15424 (N_15424,N_14357,N_14755);
nor U15425 (N_15425,N_14775,N_14584);
and U15426 (N_15426,N_14763,N_14073);
xnor U15427 (N_15427,N_14077,N_14881);
nand U15428 (N_15428,N_14470,N_14624);
nand U15429 (N_15429,N_14124,N_14774);
nand U15430 (N_15430,N_14322,N_14313);
xnor U15431 (N_15431,N_14058,N_14994);
nand U15432 (N_15432,N_14407,N_14901);
and U15433 (N_15433,N_14280,N_14659);
nor U15434 (N_15434,N_14086,N_14060);
and U15435 (N_15435,N_14813,N_14506);
or U15436 (N_15436,N_14336,N_14247);
xor U15437 (N_15437,N_14911,N_14485);
and U15438 (N_15438,N_14556,N_14290);
xor U15439 (N_15439,N_14600,N_14413);
xnor U15440 (N_15440,N_14421,N_14074);
nor U15441 (N_15441,N_14215,N_14683);
or U15442 (N_15442,N_14778,N_14009);
xnor U15443 (N_15443,N_14967,N_14111);
or U15444 (N_15444,N_14790,N_14362);
or U15445 (N_15445,N_14893,N_14263);
nor U15446 (N_15446,N_14196,N_14222);
nor U15447 (N_15447,N_14580,N_14626);
and U15448 (N_15448,N_14892,N_14296);
or U15449 (N_15449,N_14992,N_14292);
nand U15450 (N_15450,N_14199,N_14804);
or U15451 (N_15451,N_14822,N_14966);
or U15452 (N_15452,N_14219,N_14637);
or U15453 (N_15453,N_14648,N_14374);
or U15454 (N_15454,N_14422,N_14662);
or U15455 (N_15455,N_14194,N_14553);
nor U15456 (N_15456,N_14330,N_14224);
and U15457 (N_15457,N_14759,N_14307);
nand U15458 (N_15458,N_14207,N_14806);
or U15459 (N_15459,N_14269,N_14121);
and U15460 (N_15460,N_14043,N_14119);
xor U15461 (N_15461,N_14363,N_14771);
xor U15462 (N_15462,N_14973,N_14602);
or U15463 (N_15463,N_14022,N_14346);
nor U15464 (N_15464,N_14167,N_14831);
or U15465 (N_15465,N_14131,N_14590);
xor U15466 (N_15466,N_14237,N_14654);
nor U15467 (N_15467,N_14180,N_14114);
nor U15468 (N_15468,N_14411,N_14486);
xor U15469 (N_15469,N_14629,N_14005);
or U15470 (N_15470,N_14455,N_14143);
or U15471 (N_15471,N_14230,N_14116);
and U15472 (N_15472,N_14668,N_14326);
nand U15473 (N_15473,N_14367,N_14568);
and U15474 (N_15474,N_14391,N_14638);
nor U15475 (N_15475,N_14909,N_14605);
nor U15476 (N_15476,N_14558,N_14315);
xnor U15477 (N_15477,N_14565,N_14412);
nor U15478 (N_15478,N_14802,N_14044);
nand U15479 (N_15479,N_14751,N_14885);
and U15480 (N_15480,N_14204,N_14184);
and U15481 (N_15481,N_14854,N_14202);
xnor U15482 (N_15482,N_14460,N_14735);
xor U15483 (N_15483,N_14904,N_14409);
nor U15484 (N_15484,N_14430,N_14183);
nor U15485 (N_15485,N_14845,N_14308);
and U15486 (N_15486,N_14789,N_14032);
nor U15487 (N_15487,N_14325,N_14444);
or U15488 (N_15488,N_14141,N_14286);
and U15489 (N_15489,N_14518,N_14935);
xor U15490 (N_15490,N_14625,N_14379);
or U15491 (N_15491,N_14002,N_14133);
or U15492 (N_15492,N_14758,N_14097);
xnor U15493 (N_15493,N_14093,N_14511);
nand U15494 (N_15494,N_14678,N_14550);
and U15495 (N_15495,N_14311,N_14634);
nand U15496 (N_15496,N_14278,N_14770);
nor U15497 (N_15497,N_14647,N_14109);
nor U15498 (N_15498,N_14004,N_14482);
nor U15499 (N_15499,N_14406,N_14008);
nand U15500 (N_15500,N_14560,N_14361);
nand U15501 (N_15501,N_14349,N_14561);
nor U15502 (N_15502,N_14434,N_14048);
or U15503 (N_15503,N_14808,N_14502);
xor U15504 (N_15504,N_14935,N_14130);
xor U15505 (N_15505,N_14562,N_14810);
nor U15506 (N_15506,N_14904,N_14672);
nand U15507 (N_15507,N_14485,N_14187);
xor U15508 (N_15508,N_14623,N_14115);
nand U15509 (N_15509,N_14444,N_14371);
xnor U15510 (N_15510,N_14589,N_14529);
xnor U15511 (N_15511,N_14395,N_14977);
nand U15512 (N_15512,N_14564,N_14853);
nor U15513 (N_15513,N_14494,N_14562);
and U15514 (N_15514,N_14575,N_14367);
nor U15515 (N_15515,N_14935,N_14635);
or U15516 (N_15516,N_14068,N_14910);
and U15517 (N_15517,N_14122,N_14863);
or U15518 (N_15518,N_14957,N_14454);
xor U15519 (N_15519,N_14736,N_14450);
xor U15520 (N_15520,N_14905,N_14890);
and U15521 (N_15521,N_14722,N_14551);
nand U15522 (N_15522,N_14089,N_14358);
nor U15523 (N_15523,N_14300,N_14899);
nor U15524 (N_15524,N_14183,N_14794);
nand U15525 (N_15525,N_14150,N_14662);
and U15526 (N_15526,N_14025,N_14716);
and U15527 (N_15527,N_14562,N_14673);
xor U15528 (N_15528,N_14587,N_14497);
nor U15529 (N_15529,N_14188,N_14128);
or U15530 (N_15530,N_14502,N_14806);
xnor U15531 (N_15531,N_14474,N_14804);
or U15532 (N_15532,N_14983,N_14370);
xnor U15533 (N_15533,N_14201,N_14104);
nand U15534 (N_15534,N_14542,N_14022);
nand U15535 (N_15535,N_14215,N_14476);
or U15536 (N_15536,N_14668,N_14543);
and U15537 (N_15537,N_14078,N_14926);
nand U15538 (N_15538,N_14065,N_14969);
xnor U15539 (N_15539,N_14982,N_14587);
and U15540 (N_15540,N_14458,N_14512);
xnor U15541 (N_15541,N_14273,N_14042);
xor U15542 (N_15542,N_14234,N_14777);
nor U15543 (N_15543,N_14879,N_14924);
or U15544 (N_15544,N_14821,N_14252);
xor U15545 (N_15545,N_14917,N_14620);
xnor U15546 (N_15546,N_14770,N_14102);
nand U15547 (N_15547,N_14357,N_14308);
xor U15548 (N_15548,N_14563,N_14720);
nor U15549 (N_15549,N_14339,N_14848);
or U15550 (N_15550,N_14742,N_14488);
xor U15551 (N_15551,N_14657,N_14132);
nor U15552 (N_15552,N_14655,N_14023);
and U15553 (N_15553,N_14538,N_14399);
nand U15554 (N_15554,N_14795,N_14090);
nand U15555 (N_15555,N_14239,N_14213);
nand U15556 (N_15556,N_14528,N_14245);
xor U15557 (N_15557,N_14922,N_14643);
nand U15558 (N_15558,N_14993,N_14833);
xnor U15559 (N_15559,N_14745,N_14149);
nand U15560 (N_15560,N_14142,N_14584);
nor U15561 (N_15561,N_14527,N_14777);
nor U15562 (N_15562,N_14468,N_14820);
nand U15563 (N_15563,N_14087,N_14453);
nand U15564 (N_15564,N_14525,N_14446);
nor U15565 (N_15565,N_14688,N_14759);
xor U15566 (N_15566,N_14836,N_14723);
and U15567 (N_15567,N_14197,N_14593);
nand U15568 (N_15568,N_14504,N_14663);
or U15569 (N_15569,N_14153,N_14423);
xor U15570 (N_15570,N_14620,N_14696);
and U15571 (N_15571,N_14570,N_14732);
nor U15572 (N_15572,N_14365,N_14505);
nand U15573 (N_15573,N_14501,N_14859);
nor U15574 (N_15574,N_14142,N_14633);
xor U15575 (N_15575,N_14937,N_14817);
xor U15576 (N_15576,N_14662,N_14790);
nor U15577 (N_15577,N_14943,N_14509);
nand U15578 (N_15578,N_14441,N_14014);
xor U15579 (N_15579,N_14341,N_14148);
xor U15580 (N_15580,N_14010,N_14150);
xnor U15581 (N_15581,N_14683,N_14928);
nor U15582 (N_15582,N_14412,N_14873);
nand U15583 (N_15583,N_14968,N_14408);
nand U15584 (N_15584,N_14389,N_14405);
or U15585 (N_15585,N_14558,N_14525);
xnor U15586 (N_15586,N_14326,N_14901);
nand U15587 (N_15587,N_14242,N_14548);
or U15588 (N_15588,N_14091,N_14677);
xor U15589 (N_15589,N_14076,N_14514);
xor U15590 (N_15590,N_14326,N_14953);
xnor U15591 (N_15591,N_14151,N_14586);
and U15592 (N_15592,N_14742,N_14674);
nand U15593 (N_15593,N_14770,N_14429);
nand U15594 (N_15594,N_14523,N_14809);
and U15595 (N_15595,N_14797,N_14835);
or U15596 (N_15596,N_14943,N_14112);
nor U15597 (N_15597,N_14556,N_14227);
nor U15598 (N_15598,N_14156,N_14478);
xnor U15599 (N_15599,N_14413,N_14318);
or U15600 (N_15600,N_14718,N_14263);
nor U15601 (N_15601,N_14352,N_14777);
xnor U15602 (N_15602,N_14535,N_14104);
xnor U15603 (N_15603,N_14158,N_14024);
and U15604 (N_15604,N_14488,N_14559);
nor U15605 (N_15605,N_14766,N_14856);
or U15606 (N_15606,N_14892,N_14658);
nand U15607 (N_15607,N_14265,N_14617);
nand U15608 (N_15608,N_14581,N_14286);
or U15609 (N_15609,N_14532,N_14725);
xnor U15610 (N_15610,N_14054,N_14612);
nor U15611 (N_15611,N_14679,N_14018);
or U15612 (N_15612,N_14671,N_14753);
xor U15613 (N_15613,N_14020,N_14682);
xnor U15614 (N_15614,N_14614,N_14354);
or U15615 (N_15615,N_14187,N_14628);
xor U15616 (N_15616,N_14350,N_14138);
and U15617 (N_15617,N_14296,N_14614);
nand U15618 (N_15618,N_14665,N_14503);
or U15619 (N_15619,N_14485,N_14216);
and U15620 (N_15620,N_14982,N_14428);
nand U15621 (N_15621,N_14651,N_14312);
and U15622 (N_15622,N_14655,N_14454);
nor U15623 (N_15623,N_14546,N_14048);
or U15624 (N_15624,N_14604,N_14895);
xor U15625 (N_15625,N_14439,N_14163);
nor U15626 (N_15626,N_14910,N_14902);
nand U15627 (N_15627,N_14878,N_14200);
or U15628 (N_15628,N_14520,N_14682);
nor U15629 (N_15629,N_14210,N_14447);
nor U15630 (N_15630,N_14055,N_14124);
and U15631 (N_15631,N_14009,N_14318);
and U15632 (N_15632,N_14659,N_14866);
or U15633 (N_15633,N_14803,N_14916);
xnor U15634 (N_15634,N_14822,N_14233);
or U15635 (N_15635,N_14537,N_14945);
nor U15636 (N_15636,N_14735,N_14167);
nor U15637 (N_15637,N_14660,N_14416);
and U15638 (N_15638,N_14509,N_14025);
and U15639 (N_15639,N_14985,N_14001);
nand U15640 (N_15640,N_14347,N_14852);
or U15641 (N_15641,N_14763,N_14384);
or U15642 (N_15642,N_14323,N_14377);
xnor U15643 (N_15643,N_14502,N_14513);
nand U15644 (N_15644,N_14787,N_14539);
nand U15645 (N_15645,N_14592,N_14301);
nor U15646 (N_15646,N_14503,N_14160);
nor U15647 (N_15647,N_14033,N_14757);
nor U15648 (N_15648,N_14806,N_14486);
xnor U15649 (N_15649,N_14112,N_14622);
or U15650 (N_15650,N_14600,N_14033);
or U15651 (N_15651,N_14977,N_14706);
nor U15652 (N_15652,N_14956,N_14179);
nand U15653 (N_15653,N_14381,N_14205);
xor U15654 (N_15654,N_14775,N_14694);
and U15655 (N_15655,N_14422,N_14646);
nor U15656 (N_15656,N_14005,N_14480);
nor U15657 (N_15657,N_14205,N_14497);
nand U15658 (N_15658,N_14632,N_14455);
or U15659 (N_15659,N_14072,N_14262);
or U15660 (N_15660,N_14717,N_14788);
nor U15661 (N_15661,N_14441,N_14224);
or U15662 (N_15662,N_14027,N_14502);
or U15663 (N_15663,N_14785,N_14788);
nor U15664 (N_15664,N_14349,N_14742);
nand U15665 (N_15665,N_14030,N_14974);
nand U15666 (N_15666,N_14501,N_14752);
xor U15667 (N_15667,N_14437,N_14518);
and U15668 (N_15668,N_14272,N_14166);
xnor U15669 (N_15669,N_14260,N_14543);
and U15670 (N_15670,N_14743,N_14830);
nor U15671 (N_15671,N_14814,N_14340);
xor U15672 (N_15672,N_14774,N_14757);
or U15673 (N_15673,N_14314,N_14480);
or U15674 (N_15674,N_14110,N_14568);
nand U15675 (N_15675,N_14513,N_14443);
or U15676 (N_15676,N_14632,N_14139);
or U15677 (N_15677,N_14950,N_14070);
nand U15678 (N_15678,N_14240,N_14869);
nor U15679 (N_15679,N_14082,N_14853);
or U15680 (N_15680,N_14977,N_14957);
xor U15681 (N_15681,N_14569,N_14022);
or U15682 (N_15682,N_14603,N_14373);
nor U15683 (N_15683,N_14395,N_14967);
and U15684 (N_15684,N_14086,N_14406);
and U15685 (N_15685,N_14318,N_14737);
nor U15686 (N_15686,N_14970,N_14604);
nor U15687 (N_15687,N_14288,N_14413);
or U15688 (N_15688,N_14957,N_14149);
xor U15689 (N_15689,N_14807,N_14122);
nor U15690 (N_15690,N_14237,N_14372);
xnor U15691 (N_15691,N_14537,N_14534);
nor U15692 (N_15692,N_14561,N_14958);
nand U15693 (N_15693,N_14644,N_14063);
or U15694 (N_15694,N_14185,N_14310);
xnor U15695 (N_15695,N_14798,N_14225);
and U15696 (N_15696,N_14480,N_14884);
or U15697 (N_15697,N_14711,N_14091);
and U15698 (N_15698,N_14017,N_14502);
or U15699 (N_15699,N_14468,N_14982);
xor U15700 (N_15700,N_14457,N_14185);
nand U15701 (N_15701,N_14057,N_14135);
xnor U15702 (N_15702,N_14462,N_14921);
nor U15703 (N_15703,N_14215,N_14058);
nand U15704 (N_15704,N_14453,N_14922);
or U15705 (N_15705,N_14280,N_14381);
and U15706 (N_15706,N_14130,N_14850);
xnor U15707 (N_15707,N_14604,N_14466);
nand U15708 (N_15708,N_14372,N_14775);
nor U15709 (N_15709,N_14400,N_14746);
and U15710 (N_15710,N_14469,N_14325);
xnor U15711 (N_15711,N_14253,N_14683);
nand U15712 (N_15712,N_14692,N_14201);
nor U15713 (N_15713,N_14265,N_14845);
xor U15714 (N_15714,N_14363,N_14545);
and U15715 (N_15715,N_14867,N_14342);
and U15716 (N_15716,N_14914,N_14132);
nor U15717 (N_15717,N_14849,N_14065);
xnor U15718 (N_15718,N_14572,N_14748);
nand U15719 (N_15719,N_14141,N_14250);
nand U15720 (N_15720,N_14976,N_14348);
and U15721 (N_15721,N_14492,N_14650);
nor U15722 (N_15722,N_14563,N_14215);
or U15723 (N_15723,N_14341,N_14964);
nand U15724 (N_15724,N_14891,N_14105);
and U15725 (N_15725,N_14733,N_14654);
nor U15726 (N_15726,N_14459,N_14359);
nand U15727 (N_15727,N_14492,N_14914);
xor U15728 (N_15728,N_14701,N_14259);
or U15729 (N_15729,N_14242,N_14397);
or U15730 (N_15730,N_14350,N_14752);
nor U15731 (N_15731,N_14568,N_14524);
nand U15732 (N_15732,N_14990,N_14710);
or U15733 (N_15733,N_14973,N_14976);
nor U15734 (N_15734,N_14343,N_14798);
or U15735 (N_15735,N_14056,N_14240);
or U15736 (N_15736,N_14033,N_14788);
xnor U15737 (N_15737,N_14108,N_14555);
nor U15738 (N_15738,N_14659,N_14454);
nand U15739 (N_15739,N_14968,N_14500);
nor U15740 (N_15740,N_14571,N_14110);
or U15741 (N_15741,N_14891,N_14946);
and U15742 (N_15742,N_14453,N_14886);
and U15743 (N_15743,N_14983,N_14860);
or U15744 (N_15744,N_14225,N_14296);
or U15745 (N_15745,N_14092,N_14394);
nor U15746 (N_15746,N_14882,N_14824);
and U15747 (N_15747,N_14651,N_14573);
nor U15748 (N_15748,N_14127,N_14465);
nand U15749 (N_15749,N_14247,N_14226);
nor U15750 (N_15750,N_14164,N_14973);
and U15751 (N_15751,N_14942,N_14773);
nand U15752 (N_15752,N_14264,N_14644);
or U15753 (N_15753,N_14514,N_14290);
xor U15754 (N_15754,N_14759,N_14044);
xor U15755 (N_15755,N_14649,N_14466);
and U15756 (N_15756,N_14736,N_14375);
xor U15757 (N_15757,N_14776,N_14821);
nand U15758 (N_15758,N_14770,N_14023);
xnor U15759 (N_15759,N_14105,N_14102);
xnor U15760 (N_15760,N_14428,N_14758);
nand U15761 (N_15761,N_14158,N_14253);
nor U15762 (N_15762,N_14922,N_14521);
nand U15763 (N_15763,N_14053,N_14453);
and U15764 (N_15764,N_14522,N_14788);
and U15765 (N_15765,N_14947,N_14075);
or U15766 (N_15766,N_14117,N_14342);
xnor U15767 (N_15767,N_14245,N_14155);
and U15768 (N_15768,N_14147,N_14369);
nor U15769 (N_15769,N_14290,N_14450);
xnor U15770 (N_15770,N_14437,N_14122);
nand U15771 (N_15771,N_14527,N_14824);
nand U15772 (N_15772,N_14852,N_14088);
nand U15773 (N_15773,N_14177,N_14688);
xnor U15774 (N_15774,N_14326,N_14300);
or U15775 (N_15775,N_14327,N_14961);
nor U15776 (N_15776,N_14360,N_14971);
xor U15777 (N_15777,N_14790,N_14335);
nand U15778 (N_15778,N_14981,N_14851);
nor U15779 (N_15779,N_14920,N_14872);
nand U15780 (N_15780,N_14726,N_14509);
nand U15781 (N_15781,N_14893,N_14361);
xor U15782 (N_15782,N_14184,N_14139);
and U15783 (N_15783,N_14308,N_14759);
nand U15784 (N_15784,N_14464,N_14268);
nand U15785 (N_15785,N_14382,N_14092);
nor U15786 (N_15786,N_14755,N_14989);
or U15787 (N_15787,N_14125,N_14959);
and U15788 (N_15788,N_14587,N_14806);
nor U15789 (N_15789,N_14817,N_14829);
nand U15790 (N_15790,N_14028,N_14415);
xnor U15791 (N_15791,N_14513,N_14511);
and U15792 (N_15792,N_14317,N_14551);
or U15793 (N_15793,N_14502,N_14923);
or U15794 (N_15794,N_14181,N_14466);
nor U15795 (N_15795,N_14608,N_14764);
and U15796 (N_15796,N_14146,N_14861);
nand U15797 (N_15797,N_14522,N_14604);
xor U15798 (N_15798,N_14510,N_14622);
and U15799 (N_15799,N_14897,N_14990);
nand U15800 (N_15800,N_14401,N_14927);
nor U15801 (N_15801,N_14269,N_14118);
nor U15802 (N_15802,N_14811,N_14127);
nand U15803 (N_15803,N_14338,N_14311);
nand U15804 (N_15804,N_14903,N_14860);
xnor U15805 (N_15805,N_14751,N_14924);
nor U15806 (N_15806,N_14507,N_14960);
and U15807 (N_15807,N_14095,N_14348);
nand U15808 (N_15808,N_14439,N_14155);
nand U15809 (N_15809,N_14665,N_14049);
nor U15810 (N_15810,N_14760,N_14600);
nand U15811 (N_15811,N_14418,N_14740);
or U15812 (N_15812,N_14155,N_14029);
and U15813 (N_15813,N_14910,N_14052);
and U15814 (N_15814,N_14663,N_14064);
and U15815 (N_15815,N_14631,N_14490);
xor U15816 (N_15816,N_14028,N_14302);
and U15817 (N_15817,N_14141,N_14710);
or U15818 (N_15818,N_14225,N_14740);
nor U15819 (N_15819,N_14202,N_14304);
xor U15820 (N_15820,N_14397,N_14998);
or U15821 (N_15821,N_14170,N_14064);
and U15822 (N_15822,N_14279,N_14821);
or U15823 (N_15823,N_14680,N_14321);
or U15824 (N_15824,N_14189,N_14225);
nand U15825 (N_15825,N_14503,N_14234);
nand U15826 (N_15826,N_14314,N_14286);
xor U15827 (N_15827,N_14436,N_14926);
xor U15828 (N_15828,N_14826,N_14160);
nor U15829 (N_15829,N_14407,N_14093);
xnor U15830 (N_15830,N_14108,N_14028);
nor U15831 (N_15831,N_14692,N_14728);
or U15832 (N_15832,N_14496,N_14449);
xor U15833 (N_15833,N_14132,N_14231);
nand U15834 (N_15834,N_14422,N_14512);
nand U15835 (N_15835,N_14425,N_14622);
nand U15836 (N_15836,N_14055,N_14130);
nor U15837 (N_15837,N_14280,N_14085);
nand U15838 (N_15838,N_14351,N_14176);
xor U15839 (N_15839,N_14812,N_14988);
nor U15840 (N_15840,N_14760,N_14219);
xor U15841 (N_15841,N_14759,N_14441);
nor U15842 (N_15842,N_14140,N_14983);
or U15843 (N_15843,N_14664,N_14486);
xnor U15844 (N_15844,N_14612,N_14378);
xor U15845 (N_15845,N_14176,N_14864);
xnor U15846 (N_15846,N_14769,N_14058);
nand U15847 (N_15847,N_14352,N_14532);
and U15848 (N_15848,N_14303,N_14530);
nand U15849 (N_15849,N_14937,N_14450);
nand U15850 (N_15850,N_14789,N_14397);
and U15851 (N_15851,N_14399,N_14679);
or U15852 (N_15852,N_14488,N_14580);
xnor U15853 (N_15853,N_14918,N_14290);
and U15854 (N_15854,N_14725,N_14878);
nand U15855 (N_15855,N_14038,N_14449);
and U15856 (N_15856,N_14467,N_14007);
nor U15857 (N_15857,N_14898,N_14829);
nand U15858 (N_15858,N_14598,N_14626);
nand U15859 (N_15859,N_14821,N_14484);
nand U15860 (N_15860,N_14768,N_14433);
and U15861 (N_15861,N_14293,N_14641);
or U15862 (N_15862,N_14590,N_14481);
and U15863 (N_15863,N_14461,N_14345);
nand U15864 (N_15864,N_14224,N_14877);
xnor U15865 (N_15865,N_14774,N_14313);
xnor U15866 (N_15866,N_14747,N_14000);
and U15867 (N_15867,N_14412,N_14209);
xnor U15868 (N_15868,N_14311,N_14655);
and U15869 (N_15869,N_14566,N_14765);
xnor U15870 (N_15870,N_14164,N_14064);
xnor U15871 (N_15871,N_14511,N_14909);
or U15872 (N_15872,N_14614,N_14972);
nand U15873 (N_15873,N_14545,N_14999);
and U15874 (N_15874,N_14895,N_14472);
and U15875 (N_15875,N_14337,N_14474);
nor U15876 (N_15876,N_14348,N_14606);
or U15877 (N_15877,N_14005,N_14150);
and U15878 (N_15878,N_14375,N_14246);
nand U15879 (N_15879,N_14186,N_14317);
and U15880 (N_15880,N_14426,N_14472);
and U15881 (N_15881,N_14932,N_14101);
nand U15882 (N_15882,N_14831,N_14209);
or U15883 (N_15883,N_14063,N_14485);
and U15884 (N_15884,N_14483,N_14605);
or U15885 (N_15885,N_14506,N_14814);
nor U15886 (N_15886,N_14591,N_14074);
nand U15887 (N_15887,N_14468,N_14508);
nor U15888 (N_15888,N_14630,N_14534);
and U15889 (N_15889,N_14091,N_14674);
or U15890 (N_15890,N_14176,N_14631);
nor U15891 (N_15891,N_14185,N_14660);
or U15892 (N_15892,N_14816,N_14648);
and U15893 (N_15893,N_14953,N_14713);
or U15894 (N_15894,N_14996,N_14076);
xnor U15895 (N_15895,N_14908,N_14279);
nand U15896 (N_15896,N_14190,N_14987);
nand U15897 (N_15897,N_14101,N_14926);
xnor U15898 (N_15898,N_14227,N_14935);
xnor U15899 (N_15899,N_14229,N_14863);
and U15900 (N_15900,N_14351,N_14823);
nor U15901 (N_15901,N_14267,N_14283);
or U15902 (N_15902,N_14095,N_14884);
nand U15903 (N_15903,N_14057,N_14291);
xor U15904 (N_15904,N_14146,N_14651);
and U15905 (N_15905,N_14936,N_14621);
nand U15906 (N_15906,N_14347,N_14861);
nor U15907 (N_15907,N_14159,N_14556);
xnor U15908 (N_15908,N_14978,N_14830);
or U15909 (N_15909,N_14453,N_14341);
or U15910 (N_15910,N_14477,N_14023);
nand U15911 (N_15911,N_14627,N_14005);
or U15912 (N_15912,N_14829,N_14274);
xor U15913 (N_15913,N_14511,N_14663);
nor U15914 (N_15914,N_14175,N_14688);
or U15915 (N_15915,N_14575,N_14855);
nand U15916 (N_15916,N_14104,N_14331);
and U15917 (N_15917,N_14837,N_14318);
nand U15918 (N_15918,N_14857,N_14149);
and U15919 (N_15919,N_14059,N_14693);
and U15920 (N_15920,N_14942,N_14438);
or U15921 (N_15921,N_14725,N_14207);
xor U15922 (N_15922,N_14853,N_14925);
and U15923 (N_15923,N_14445,N_14665);
nand U15924 (N_15924,N_14503,N_14370);
xor U15925 (N_15925,N_14826,N_14321);
or U15926 (N_15926,N_14454,N_14248);
nand U15927 (N_15927,N_14862,N_14433);
and U15928 (N_15928,N_14764,N_14416);
xnor U15929 (N_15929,N_14661,N_14577);
or U15930 (N_15930,N_14477,N_14595);
or U15931 (N_15931,N_14645,N_14037);
and U15932 (N_15932,N_14131,N_14462);
nor U15933 (N_15933,N_14295,N_14558);
or U15934 (N_15934,N_14572,N_14118);
xnor U15935 (N_15935,N_14398,N_14460);
and U15936 (N_15936,N_14616,N_14256);
nor U15937 (N_15937,N_14420,N_14307);
nand U15938 (N_15938,N_14829,N_14621);
xor U15939 (N_15939,N_14791,N_14575);
and U15940 (N_15940,N_14176,N_14088);
nor U15941 (N_15941,N_14454,N_14528);
xor U15942 (N_15942,N_14145,N_14790);
and U15943 (N_15943,N_14259,N_14156);
nand U15944 (N_15944,N_14395,N_14699);
nand U15945 (N_15945,N_14958,N_14580);
nand U15946 (N_15946,N_14429,N_14065);
and U15947 (N_15947,N_14901,N_14189);
nor U15948 (N_15948,N_14004,N_14783);
or U15949 (N_15949,N_14147,N_14890);
nor U15950 (N_15950,N_14555,N_14916);
and U15951 (N_15951,N_14837,N_14936);
nor U15952 (N_15952,N_14258,N_14304);
nand U15953 (N_15953,N_14259,N_14046);
nor U15954 (N_15954,N_14935,N_14639);
xnor U15955 (N_15955,N_14331,N_14447);
and U15956 (N_15956,N_14803,N_14417);
xor U15957 (N_15957,N_14591,N_14675);
and U15958 (N_15958,N_14257,N_14515);
nand U15959 (N_15959,N_14239,N_14435);
xnor U15960 (N_15960,N_14133,N_14260);
or U15961 (N_15961,N_14917,N_14857);
xor U15962 (N_15962,N_14792,N_14184);
and U15963 (N_15963,N_14330,N_14771);
xor U15964 (N_15964,N_14026,N_14324);
xor U15965 (N_15965,N_14029,N_14086);
or U15966 (N_15966,N_14426,N_14111);
or U15967 (N_15967,N_14952,N_14612);
nor U15968 (N_15968,N_14876,N_14491);
or U15969 (N_15969,N_14232,N_14444);
or U15970 (N_15970,N_14457,N_14838);
nor U15971 (N_15971,N_14680,N_14372);
xor U15972 (N_15972,N_14902,N_14737);
nand U15973 (N_15973,N_14083,N_14448);
and U15974 (N_15974,N_14971,N_14167);
xor U15975 (N_15975,N_14256,N_14201);
xor U15976 (N_15976,N_14777,N_14353);
or U15977 (N_15977,N_14865,N_14151);
nor U15978 (N_15978,N_14074,N_14726);
xor U15979 (N_15979,N_14306,N_14247);
or U15980 (N_15980,N_14810,N_14556);
nand U15981 (N_15981,N_14814,N_14969);
and U15982 (N_15982,N_14465,N_14057);
xor U15983 (N_15983,N_14457,N_14880);
xnor U15984 (N_15984,N_14300,N_14685);
and U15985 (N_15985,N_14821,N_14046);
nor U15986 (N_15986,N_14661,N_14758);
xor U15987 (N_15987,N_14970,N_14333);
or U15988 (N_15988,N_14103,N_14902);
nor U15989 (N_15989,N_14218,N_14080);
nand U15990 (N_15990,N_14335,N_14361);
and U15991 (N_15991,N_14429,N_14843);
xor U15992 (N_15992,N_14094,N_14377);
or U15993 (N_15993,N_14492,N_14098);
xnor U15994 (N_15994,N_14247,N_14492);
or U15995 (N_15995,N_14985,N_14152);
xnor U15996 (N_15996,N_14670,N_14291);
or U15997 (N_15997,N_14067,N_14582);
and U15998 (N_15998,N_14328,N_14731);
or U15999 (N_15999,N_14860,N_14258);
or U16000 (N_16000,N_15694,N_15868);
nand U16001 (N_16001,N_15909,N_15944);
nand U16002 (N_16002,N_15563,N_15369);
xor U16003 (N_16003,N_15424,N_15255);
nand U16004 (N_16004,N_15480,N_15198);
xor U16005 (N_16005,N_15608,N_15354);
nand U16006 (N_16006,N_15467,N_15123);
and U16007 (N_16007,N_15936,N_15578);
xor U16008 (N_16008,N_15698,N_15197);
nor U16009 (N_16009,N_15693,N_15590);
nor U16010 (N_16010,N_15705,N_15361);
nand U16011 (N_16011,N_15611,N_15171);
or U16012 (N_16012,N_15200,N_15027);
xor U16013 (N_16013,N_15904,N_15302);
xnor U16014 (N_16014,N_15525,N_15627);
nand U16015 (N_16015,N_15446,N_15718);
xnor U16016 (N_16016,N_15938,N_15143);
and U16017 (N_16017,N_15392,N_15675);
nand U16018 (N_16018,N_15210,N_15457);
xor U16019 (N_16019,N_15857,N_15914);
xnor U16020 (N_16020,N_15711,N_15798);
xor U16021 (N_16021,N_15336,N_15283);
nand U16022 (N_16022,N_15425,N_15107);
xor U16023 (N_16023,N_15257,N_15008);
xor U16024 (N_16024,N_15286,N_15014);
and U16025 (N_16025,N_15539,N_15845);
nor U16026 (N_16026,N_15137,N_15090);
or U16027 (N_16027,N_15294,N_15267);
nand U16028 (N_16028,N_15109,N_15524);
nor U16029 (N_16029,N_15814,N_15553);
or U16030 (N_16030,N_15103,N_15493);
or U16031 (N_16031,N_15933,N_15818);
nand U16032 (N_16032,N_15466,N_15812);
nor U16033 (N_16033,N_15727,N_15229);
or U16034 (N_16034,N_15385,N_15511);
nand U16035 (N_16035,N_15783,N_15562);
or U16036 (N_16036,N_15013,N_15376);
and U16037 (N_16037,N_15745,N_15777);
and U16038 (N_16038,N_15737,N_15174);
and U16039 (N_16039,N_15079,N_15431);
or U16040 (N_16040,N_15688,N_15897);
and U16041 (N_16041,N_15037,N_15266);
or U16042 (N_16042,N_15854,N_15715);
nor U16043 (N_16043,N_15543,N_15327);
xor U16044 (N_16044,N_15568,N_15018);
xor U16045 (N_16045,N_15393,N_15864);
or U16046 (N_16046,N_15980,N_15499);
nand U16047 (N_16047,N_15348,N_15606);
and U16048 (N_16048,N_15020,N_15068);
nor U16049 (N_16049,N_15112,N_15146);
and U16050 (N_16050,N_15333,N_15155);
or U16051 (N_16051,N_15894,N_15866);
xor U16052 (N_16052,N_15755,N_15587);
and U16053 (N_16053,N_15199,N_15922);
xor U16054 (N_16054,N_15303,N_15411);
or U16055 (N_16055,N_15192,N_15622);
or U16056 (N_16056,N_15040,N_15416);
and U16057 (N_16057,N_15988,N_15961);
xnor U16058 (N_16058,N_15477,N_15990);
xnor U16059 (N_16059,N_15338,N_15643);
or U16060 (N_16060,N_15397,N_15722);
nor U16061 (N_16061,N_15029,N_15637);
and U16062 (N_16062,N_15714,N_15928);
nand U16063 (N_16063,N_15053,N_15374);
or U16064 (N_16064,N_15902,N_15599);
xnor U16065 (N_16065,N_15005,N_15516);
or U16066 (N_16066,N_15849,N_15832);
or U16067 (N_16067,N_15660,N_15263);
xnor U16068 (N_16068,N_15311,N_15567);
nor U16069 (N_16069,N_15597,N_15676);
nand U16070 (N_16070,N_15974,N_15158);
xnor U16071 (N_16071,N_15180,N_15323);
nand U16072 (N_16072,N_15825,N_15918);
or U16073 (N_16073,N_15696,N_15657);
nand U16074 (N_16074,N_15681,N_15373);
nand U16075 (N_16075,N_15246,N_15547);
nand U16076 (N_16076,N_15429,N_15955);
xor U16077 (N_16077,N_15679,N_15650);
nand U16078 (N_16078,N_15991,N_15639);
nand U16079 (N_16079,N_15796,N_15205);
nor U16080 (N_16080,N_15548,N_15498);
xor U16081 (N_16081,N_15830,N_15596);
xor U16082 (N_16082,N_15025,N_15779);
nand U16083 (N_16083,N_15189,N_15245);
and U16084 (N_16084,N_15757,N_15566);
xnor U16085 (N_16085,N_15736,N_15747);
nand U16086 (N_16086,N_15748,N_15207);
or U16087 (N_16087,N_15546,N_15196);
or U16088 (N_16088,N_15811,N_15447);
or U16089 (N_16089,N_15863,N_15708);
and U16090 (N_16090,N_15906,N_15970);
or U16091 (N_16091,N_15276,N_15649);
nor U16092 (N_16092,N_15867,N_15326);
or U16093 (N_16093,N_15038,N_15950);
and U16094 (N_16094,N_15407,N_15600);
and U16095 (N_16095,N_15529,N_15069);
xor U16096 (N_16096,N_15317,N_15280);
and U16097 (N_16097,N_15182,N_15664);
and U16098 (N_16098,N_15042,N_15172);
nor U16099 (N_16099,N_15278,N_15084);
nor U16100 (N_16100,N_15176,N_15709);
nand U16101 (N_16101,N_15169,N_15793);
xor U16102 (N_16102,N_15764,N_15775);
nand U16103 (N_16103,N_15206,N_15468);
or U16104 (N_16104,N_15828,N_15086);
nand U16105 (N_16105,N_15778,N_15758);
nor U16106 (N_16106,N_15035,N_15762);
nand U16107 (N_16107,N_15476,N_15532);
nand U16108 (N_16108,N_15183,N_15419);
or U16109 (N_16109,N_15337,N_15167);
nand U16110 (N_16110,N_15475,N_15380);
or U16111 (N_16111,N_15570,N_15931);
nor U16112 (N_16112,N_15929,N_15509);
nor U16113 (N_16113,N_15275,N_15114);
xnor U16114 (N_16114,N_15871,N_15417);
xnor U16115 (N_16115,N_15617,N_15594);
xnor U16116 (N_16116,N_15043,N_15973);
or U16117 (N_16117,N_15349,N_15690);
nand U16118 (N_16118,N_15619,N_15653);
xor U16119 (N_16119,N_15220,N_15557);
or U16120 (N_16120,N_15923,N_15471);
nand U16121 (N_16121,N_15707,N_15217);
nand U16122 (N_16122,N_15728,N_15223);
or U16123 (N_16123,N_15773,N_15844);
and U16124 (N_16124,N_15971,N_15989);
and U16125 (N_16125,N_15651,N_15683);
or U16126 (N_16126,N_15147,N_15833);
and U16127 (N_16127,N_15876,N_15921);
nor U16128 (N_16128,N_15249,N_15074);
and U16129 (N_16129,N_15256,N_15061);
or U16130 (N_16130,N_15451,N_15449);
or U16131 (N_16131,N_15315,N_15607);
or U16132 (N_16132,N_15692,N_15157);
or U16133 (N_16133,N_15238,N_15211);
and U16134 (N_16134,N_15487,N_15148);
nand U16135 (N_16135,N_15852,N_15356);
xnor U16136 (N_16136,N_15228,N_15436);
nor U16137 (N_16137,N_15910,N_15605);
xnor U16138 (N_16138,N_15873,N_15343);
xor U16139 (N_16139,N_15295,N_15995);
nor U16140 (N_16140,N_15463,N_15222);
or U16141 (N_16141,N_15292,N_15017);
nor U16142 (N_16142,N_15111,N_15335);
and U16143 (N_16143,N_15898,N_15352);
xnor U16144 (N_16144,N_15638,N_15884);
xnor U16145 (N_16145,N_15161,N_15413);
nor U16146 (N_16146,N_15368,N_15260);
or U16147 (N_16147,N_15485,N_15494);
xor U16148 (N_16148,N_15691,N_15791);
and U16149 (N_16149,N_15756,N_15846);
xor U16150 (N_16150,N_15241,N_15659);
nor U16151 (N_16151,N_15099,N_15306);
and U16152 (N_16152,N_15089,N_15345);
xor U16153 (N_16153,N_15666,N_15126);
xnor U16154 (N_16154,N_15558,N_15486);
or U16155 (N_16155,N_15689,N_15853);
xor U16156 (N_16156,N_15328,N_15110);
or U16157 (N_16157,N_15517,N_15507);
nor U16158 (N_16158,N_15877,N_15882);
and U16159 (N_16159,N_15244,N_15859);
and U16160 (N_16160,N_15193,N_15290);
or U16161 (N_16161,N_15802,N_15996);
nor U16162 (N_16162,N_15066,N_15184);
or U16163 (N_16163,N_15685,N_15761);
xnor U16164 (N_16164,N_15700,N_15998);
or U16165 (N_16165,N_15874,N_15542);
nor U16166 (N_16166,N_15734,N_15076);
or U16167 (N_16167,N_15564,N_15132);
or U16168 (N_16168,N_15344,N_15699);
or U16169 (N_16169,N_15975,N_15760);
nor U16170 (N_16170,N_15581,N_15746);
or U16171 (N_16171,N_15384,N_15834);
nor U16172 (N_16172,N_15496,N_15209);
xor U16173 (N_16173,N_15360,N_15396);
and U16174 (N_16174,N_15939,N_15686);
nand U16175 (N_16175,N_15536,N_15763);
and U16176 (N_16176,N_15404,N_15506);
nand U16177 (N_16177,N_15682,N_15164);
and U16178 (N_16178,N_15837,N_15963);
nor U16179 (N_16179,N_15582,N_15829);
or U16180 (N_16180,N_15883,N_15967);
or U16181 (N_16181,N_15258,N_15454);
xnor U16182 (N_16182,N_15966,N_15843);
nand U16183 (N_16183,N_15838,N_15461);
nand U16184 (N_16184,N_15815,N_15309);
or U16185 (N_16185,N_15034,N_15389);
and U16186 (N_16186,N_15819,N_15795);
nand U16187 (N_16187,N_15296,N_15119);
and U16188 (N_16188,N_15213,N_15505);
or U16189 (N_16189,N_15538,N_15554);
nor U16190 (N_16190,N_15372,N_15526);
nor U16191 (N_16191,N_15022,N_15887);
nand U16192 (N_16192,N_15273,N_15319);
nand U16193 (N_16193,N_15188,N_15628);
nor U16194 (N_16194,N_15999,N_15142);
nor U16195 (N_16195,N_15221,N_15515);
xor U16196 (N_16196,N_15813,N_15214);
xor U16197 (N_16197,N_15572,N_15836);
and U16198 (N_16198,N_15106,N_15635);
nor U16199 (N_16199,N_15121,N_15907);
nor U16200 (N_16200,N_15488,N_15865);
and U16201 (N_16201,N_15208,N_15321);
nand U16202 (N_16202,N_15674,N_15009);
or U16203 (N_16203,N_15264,N_15655);
nand U16204 (N_16204,N_15561,N_15924);
nand U16205 (N_16205,N_15300,N_15723);
and U16206 (N_16206,N_15115,N_15168);
nand U16207 (N_16207,N_15489,N_15672);
xor U16208 (N_16208,N_15589,N_15041);
or U16209 (N_16209,N_15891,N_15574);
or U16210 (N_16210,N_15093,N_15353);
and U16211 (N_16211,N_15301,N_15786);
nor U16212 (N_16212,N_15268,N_15194);
xor U16213 (N_16213,N_15972,N_15329);
and U16214 (N_16214,N_15004,N_15334);
and U16215 (N_16215,N_15410,N_15768);
xor U16216 (N_16216,N_15801,N_15265);
nand U16217 (N_16217,N_15156,N_15797);
xnor U16218 (N_16218,N_15781,N_15946);
nor U16219 (N_16219,N_15453,N_15144);
nand U16220 (N_16220,N_15339,N_15231);
nor U16221 (N_16221,N_15642,N_15550);
nor U16222 (N_16222,N_15519,N_15036);
nor U16223 (N_16223,N_15085,N_15776);
or U16224 (N_16224,N_15163,N_15378);
nand U16225 (N_16225,N_15418,N_15011);
and U16226 (N_16226,N_15512,N_15919);
and U16227 (N_16227,N_15633,N_15400);
and U16228 (N_16228,N_15710,N_15983);
nor U16229 (N_16229,N_15913,N_15624);
nor U16230 (N_16230,N_15997,N_15771);
nor U16231 (N_16231,N_15096,N_15740);
nand U16232 (N_16232,N_15847,N_15316);
xor U16233 (N_16233,N_15881,N_15872);
and U16234 (N_16234,N_15120,N_15433);
nor U16235 (N_16235,N_15347,N_15495);
nand U16236 (N_16236,N_15595,N_15888);
nor U16237 (N_16237,N_15088,N_15077);
xor U16238 (N_16238,N_15340,N_15289);
nor U16239 (N_16239,N_15861,N_15252);
or U16240 (N_16240,N_15405,N_15021);
or U16241 (N_16241,N_15960,N_15362);
nor U16242 (N_16242,N_15942,N_15926);
and U16243 (N_16243,N_15704,N_15769);
xnor U16244 (N_16244,N_15750,N_15363);
xor U16245 (N_16245,N_15911,N_15072);
nor U16246 (N_16246,N_15070,N_15226);
xnor U16247 (N_16247,N_15320,N_15994);
or U16248 (N_16248,N_15242,N_15313);
xnor U16249 (N_16249,N_15420,N_15903);
nand U16250 (N_16250,N_15139,N_15724);
and U16251 (N_16251,N_15437,N_15422);
or U16252 (N_16252,N_15145,N_15428);
nand U16253 (N_16253,N_15592,N_15917);
and U16254 (N_16254,N_15039,N_15219);
nor U16255 (N_16255,N_15695,N_15170);
nor U16256 (N_16256,N_15678,N_15807);
or U16257 (N_16257,N_15535,N_15002);
nor U16258 (N_16258,N_15359,N_15725);
xnor U16259 (N_16259,N_15782,N_15190);
xor U16260 (N_16260,N_15297,N_15717);
xor U16261 (N_16261,N_15993,N_15982);
and U16262 (N_16262,N_15181,N_15341);
xor U16263 (N_16263,N_15150,N_15886);
or U16264 (N_16264,N_15024,N_15408);
nor U16265 (N_16265,N_15518,N_15860);
or U16266 (N_16266,N_15810,N_15234);
or U16267 (N_16267,N_15443,N_15033);
xor U16268 (N_16268,N_15094,N_15987);
or U16269 (N_16269,N_15056,N_15288);
and U16270 (N_16270,N_15530,N_15159);
nand U16271 (N_16271,N_15965,N_15007);
and U16272 (N_16272,N_15920,N_15375);
nand U16273 (N_16273,N_15104,N_15136);
xnor U16274 (N_16274,N_15645,N_15279);
xnor U16275 (N_16275,N_15555,N_15230);
nor U16276 (N_16276,N_15383,N_15935);
nand U16277 (N_16277,N_15012,N_15464);
or U16278 (N_16278,N_15957,N_15116);
nand U16279 (N_16279,N_15441,N_15614);
nand U16280 (N_16280,N_15048,N_15804);
nor U16281 (N_16281,N_15522,N_15125);
nor U16282 (N_16282,N_15945,N_15665);
nor U16283 (N_16283,N_15749,N_15789);
and U16284 (N_16284,N_15177,N_15806);
nand U16285 (N_16285,N_15805,N_15367);
nand U16286 (N_16286,N_15049,N_15262);
xnor U16287 (N_16287,N_15565,N_15346);
or U16288 (N_16288,N_15430,N_15491);
or U16289 (N_16289,N_15379,N_15308);
nand U16290 (N_16290,N_15948,N_15059);
and U16291 (N_16291,N_15000,N_15968);
and U16292 (N_16292,N_15215,N_15365);
nand U16293 (N_16293,N_15803,N_15299);
xor U16294 (N_16294,N_15044,N_15272);
and U16295 (N_16295,N_15186,N_15500);
xnor U16296 (N_16296,N_15324,N_15479);
xor U16297 (N_16297,N_15701,N_15735);
nor U16298 (N_16298,N_15523,N_15890);
or U16299 (N_16299,N_15381,N_15458);
nor U16300 (N_16300,N_15473,N_15395);
nand U16301 (N_16301,N_15584,N_15744);
nor U16302 (N_16302,N_15490,N_15460);
nand U16303 (N_16303,N_15981,N_15527);
nor U16304 (N_16304,N_15827,N_15281);
nor U16305 (N_16305,N_15050,N_15482);
nor U16306 (N_16306,N_15001,N_15235);
xnor U16307 (N_16307,N_15092,N_15149);
xnor U16308 (N_16308,N_15179,N_15304);
or U16309 (N_16309,N_15175,N_15842);
or U16310 (N_16310,N_15733,N_15409);
nor U16311 (N_16311,N_15060,N_15604);
xnor U16312 (N_16312,N_15835,N_15661);
and U16313 (N_16313,N_15394,N_15081);
nand U16314 (N_16314,N_15218,N_15371);
or U16315 (N_16315,N_15616,N_15236);
xnor U16316 (N_16316,N_15387,N_15067);
nor U16317 (N_16317,N_15438,N_15969);
nand U16318 (N_16318,N_15954,N_15593);
nor U16319 (N_16319,N_15502,N_15648);
and U16320 (N_16320,N_15571,N_15366);
nor U16321 (N_16321,N_15481,N_15591);
or U16322 (N_16322,N_15652,N_15065);
nand U16323 (N_16323,N_15559,N_15951);
nor U16324 (N_16324,N_15195,N_15401);
nand U16325 (N_16325,N_15520,N_15253);
nand U16326 (N_16326,N_15702,N_15127);
and U16327 (N_16327,N_15122,N_15452);
or U16328 (N_16328,N_15588,N_15752);
nand U16329 (N_16329,N_15620,N_15545);
nand U16330 (N_16330,N_15899,N_15284);
and U16331 (N_16331,N_15091,N_15792);
and U16332 (N_16332,N_15046,N_15823);
and U16333 (N_16333,N_15869,N_15023);
nand U16334 (N_16334,N_15754,N_15154);
nor U16335 (N_16335,N_15006,N_15271);
nor U16336 (N_16336,N_15134,N_15809);
or U16337 (N_16337,N_15469,N_15817);
nor U16338 (N_16338,N_15851,N_15816);
xor U16339 (N_16339,N_15270,N_15730);
nand U16340 (N_16340,N_15108,N_15293);
nor U16341 (N_16341,N_15098,N_15626);
nand U16342 (N_16342,N_15448,N_15322);
nor U16343 (N_16343,N_15885,N_15259);
xor U16344 (N_16344,N_15130,N_15673);
xor U16345 (N_16345,N_15992,N_15738);
xor U16346 (N_16346,N_15332,N_15765);
and U16347 (N_16347,N_15185,N_15892);
xor U16348 (N_16348,N_15102,N_15483);
nand U16349 (N_16349,N_15569,N_15985);
and U16350 (N_16350,N_15455,N_15414);
nand U16351 (N_16351,N_15426,N_15028);
xnor U16352 (N_16352,N_15427,N_15759);
nor U16353 (N_16353,N_15741,N_15669);
xnor U16354 (N_16354,N_15943,N_15064);
xor U16355 (N_16355,N_15100,N_15585);
or U16356 (N_16356,N_15057,N_15583);
nand U16357 (N_16357,N_15879,N_15403);
nand U16358 (N_16358,N_15406,N_15351);
or U16359 (N_16359,N_15878,N_15031);
nor U16360 (N_16360,N_15124,N_15824);
nand U16361 (N_16361,N_15251,N_15916);
and U16362 (N_16362,N_15751,N_15537);
xor U16363 (N_16363,N_15634,N_15743);
nor U16364 (N_16364,N_15402,N_15610);
nand U16365 (N_16365,N_15784,N_15603);
and U16366 (N_16366,N_15831,N_15629);
and U16367 (N_16367,N_15510,N_15318);
or U16368 (N_16368,N_15905,N_15047);
nor U16369 (N_16369,N_15434,N_15254);
and U16370 (N_16370,N_15915,N_15656);
and U16371 (N_16371,N_15580,N_15984);
nand U16372 (N_16372,N_15342,N_15766);
nor U16373 (N_16373,N_15577,N_15941);
nand U16374 (N_16374,N_15662,N_15623);
and U16375 (N_16375,N_15331,N_15314);
or U16376 (N_16376,N_15613,N_15032);
xnor U16377 (N_16377,N_15250,N_15514);
nand U16378 (N_16378,N_15151,N_15128);
xor U16379 (N_16379,N_15390,N_15439);
or U16380 (N_16380,N_15528,N_15947);
nor U16381 (N_16381,N_15551,N_15855);
nand U16382 (N_16382,N_15140,N_15640);
nor U16383 (N_16383,N_15647,N_15932);
xor U16384 (N_16384,N_15513,N_15978);
and U16385 (N_16385,N_15556,N_15956);
nor U16386 (N_16386,N_15573,N_15117);
xnor U16387 (N_16387,N_15141,N_15977);
and U16388 (N_16388,N_15800,N_15310);
xor U16389 (N_16389,N_15080,N_15412);
and U16390 (N_16390,N_15398,N_15135);
and U16391 (N_16391,N_15073,N_15575);
and U16392 (N_16392,N_15325,N_15153);
or U16393 (N_16393,N_15636,N_15927);
or U16394 (N_16394,N_15051,N_15162);
xor U16395 (N_16395,N_15780,N_15612);
or U16396 (N_16396,N_15601,N_15560);
xor U16397 (N_16397,N_15875,N_15609);
and U16398 (N_16398,N_15986,N_15391);
xnor U16399 (N_16399,N_15357,N_15287);
xor U16400 (N_16400,N_15152,N_15671);
nor U16401 (N_16401,N_15083,N_15165);
xnor U16402 (N_16402,N_15787,N_15191);
nand U16403 (N_16403,N_15052,N_15531);
or U16404 (N_16404,N_15621,N_15456);
and U16405 (N_16405,N_15233,N_15243);
nand U16406 (N_16406,N_15201,N_15386);
or U16407 (N_16407,N_15484,N_15767);
and U16408 (N_16408,N_15862,N_15870);
and U16409 (N_16409,N_15474,N_15774);
xor U16410 (N_16410,N_15712,N_15719);
and U16411 (N_16411,N_15078,N_15858);
xnor U16412 (N_16412,N_15421,N_15742);
nor U16413 (N_16413,N_15912,N_15631);
xnor U16414 (N_16414,N_15677,N_15680);
or U16415 (N_16415,N_15358,N_15298);
nor U16416 (N_16416,N_15462,N_15937);
or U16417 (N_16417,N_15269,N_15504);
nor U16418 (N_16418,N_15839,N_15841);
or U16419 (N_16419,N_15015,N_15227);
nand U16420 (N_16420,N_15794,N_15544);
nand U16421 (N_16421,N_15703,N_15202);
and U16422 (N_16422,N_15895,N_15160);
nor U16423 (N_16423,N_15848,N_15350);
and U16424 (N_16424,N_15355,N_15055);
or U16425 (N_16425,N_15850,N_15440);
or U16426 (N_16426,N_15465,N_15247);
xnor U16427 (N_16427,N_15497,N_15618);
nor U16428 (N_16428,N_15670,N_15654);
nand U16429 (N_16429,N_15901,N_15896);
xor U16430 (N_16430,N_15641,N_15739);
xnor U16431 (N_16431,N_15203,N_15706);
nand U16432 (N_16432,N_15062,N_15131);
nor U16433 (N_16433,N_15178,N_15054);
or U16434 (N_16434,N_15840,N_15435);
nor U16435 (N_16435,N_15785,N_15101);
or U16436 (N_16436,N_15658,N_15097);
nor U16437 (N_16437,N_15503,N_15625);
nor U16438 (N_16438,N_15330,N_15713);
nor U16439 (N_16439,N_15095,N_15533);
or U16440 (N_16440,N_15964,N_15930);
and U16441 (N_16441,N_15808,N_15684);
nand U16442 (N_16442,N_15118,N_15889);
nand U16443 (N_16443,N_15312,N_15225);
or U16444 (N_16444,N_15377,N_15598);
or U16445 (N_16445,N_15644,N_15432);
nor U16446 (N_16446,N_15893,N_15285);
xnor U16447 (N_16447,N_15282,N_15138);
or U16448 (N_16448,N_15204,N_15307);
nor U16449 (N_16449,N_15716,N_15822);
or U16450 (N_16450,N_15113,N_15949);
xor U16451 (N_16451,N_15261,N_15364);
and U16452 (N_16452,N_15087,N_15444);
nand U16453 (N_16453,N_15212,N_15900);
and U16454 (N_16454,N_15472,N_15772);
xnor U16455 (N_16455,N_15521,N_15668);
nor U16456 (N_16456,N_15925,N_15576);
and U16457 (N_16457,N_15187,N_15075);
xnor U16458 (N_16458,N_15442,N_15237);
or U16459 (N_16459,N_15045,N_15697);
and U16460 (N_16460,N_15459,N_15277);
nand U16461 (N_16461,N_15908,N_15962);
or U16462 (N_16462,N_15770,N_15731);
xor U16463 (N_16463,N_15082,N_15720);
nand U16464 (N_16464,N_15370,N_15552);
nand U16465 (N_16465,N_15240,N_15940);
and U16466 (N_16466,N_15239,N_15173);
xor U16467 (N_16467,N_15615,N_15016);
and U16468 (N_16468,N_15415,N_15450);
xor U16469 (N_16469,N_15788,N_15726);
nand U16470 (N_16470,N_15216,N_15058);
nand U16471 (N_16471,N_15508,N_15790);
or U16472 (N_16472,N_15958,N_15541);
or U16473 (N_16473,N_15953,N_15382);
xor U16474 (N_16474,N_15071,N_15026);
xnor U16475 (N_16475,N_15630,N_15826);
nor U16476 (N_16476,N_15445,N_15721);
and U16477 (N_16477,N_15248,N_15534);
nand U16478 (N_16478,N_15667,N_15478);
xnor U16479 (N_16479,N_15952,N_15129);
or U16480 (N_16480,N_15019,N_15010);
nand U16481 (N_16481,N_15729,N_15003);
and U16482 (N_16482,N_15501,N_15232);
nand U16483 (N_16483,N_15540,N_15799);
nor U16484 (N_16484,N_15687,N_15291);
nor U16485 (N_16485,N_15105,N_15820);
or U16486 (N_16486,N_15166,N_15732);
and U16487 (N_16487,N_15470,N_15934);
xnor U16488 (N_16488,N_15959,N_15224);
nor U16489 (N_16489,N_15586,N_15979);
xnor U16490 (N_16490,N_15492,N_15305);
or U16491 (N_16491,N_15602,N_15663);
xnor U16492 (N_16492,N_15030,N_15753);
xnor U16493 (N_16493,N_15549,N_15133);
nor U16494 (N_16494,N_15579,N_15646);
or U16495 (N_16495,N_15856,N_15880);
nand U16496 (N_16496,N_15388,N_15976);
nor U16497 (N_16497,N_15063,N_15423);
or U16498 (N_16498,N_15821,N_15399);
nand U16499 (N_16499,N_15632,N_15274);
nor U16500 (N_16500,N_15389,N_15407);
and U16501 (N_16501,N_15474,N_15455);
and U16502 (N_16502,N_15574,N_15636);
and U16503 (N_16503,N_15503,N_15950);
nor U16504 (N_16504,N_15275,N_15782);
xor U16505 (N_16505,N_15132,N_15312);
nand U16506 (N_16506,N_15183,N_15941);
or U16507 (N_16507,N_15712,N_15094);
nand U16508 (N_16508,N_15348,N_15844);
and U16509 (N_16509,N_15771,N_15803);
nor U16510 (N_16510,N_15804,N_15401);
xnor U16511 (N_16511,N_15575,N_15016);
and U16512 (N_16512,N_15392,N_15513);
or U16513 (N_16513,N_15275,N_15547);
nor U16514 (N_16514,N_15990,N_15361);
and U16515 (N_16515,N_15889,N_15260);
or U16516 (N_16516,N_15952,N_15111);
nor U16517 (N_16517,N_15004,N_15702);
nand U16518 (N_16518,N_15820,N_15624);
nand U16519 (N_16519,N_15462,N_15140);
nand U16520 (N_16520,N_15372,N_15879);
nor U16521 (N_16521,N_15609,N_15438);
and U16522 (N_16522,N_15465,N_15774);
nor U16523 (N_16523,N_15958,N_15829);
xor U16524 (N_16524,N_15041,N_15194);
and U16525 (N_16525,N_15728,N_15617);
nor U16526 (N_16526,N_15471,N_15292);
nor U16527 (N_16527,N_15055,N_15777);
xnor U16528 (N_16528,N_15565,N_15223);
or U16529 (N_16529,N_15565,N_15097);
and U16530 (N_16530,N_15834,N_15750);
nand U16531 (N_16531,N_15012,N_15926);
or U16532 (N_16532,N_15303,N_15844);
nand U16533 (N_16533,N_15375,N_15221);
and U16534 (N_16534,N_15377,N_15986);
nor U16535 (N_16535,N_15987,N_15530);
nor U16536 (N_16536,N_15392,N_15255);
or U16537 (N_16537,N_15687,N_15068);
xor U16538 (N_16538,N_15009,N_15518);
xor U16539 (N_16539,N_15631,N_15502);
xor U16540 (N_16540,N_15990,N_15522);
nand U16541 (N_16541,N_15998,N_15264);
xnor U16542 (N_16542,N_15498,N_15299);
nand U16543 (N_16543,N_15015,N_15764);
xor U16544 (N_16544,N_15597,N_15912);
nand U16545 (N_16545,N_15030,N_15660);
xor U16546 (N_16546,N_15688,N_15521);
or U16547 (N_16547,N_15783,N_15266);
nand U16548 (N_16548,N_15865,N_15275);
and U16549 (N_16549,N_15019,N_15432);
nand U16550 (N_16550,N_15958,N_15372);
nor U16551 (N_16551,N_15359,N_15577);
xor U16552 (N_16552,N_15525,N_15959);
or U16553 (N_16553,N_15809,N_15748);
or U16554 (N_16554,N_15683,N_15176);
nand U16555 (N_16555,N_15685,N_15794);
and U16556 (N_16556,N_15316,N_15797);
nand U16557 (N_16557,N_15538,N_15325);
and U16558 (N_16558,N_15131,N_15469);
nor U16559 (N_16559,N_15800,N_15207);
or U16560 (N_16560,N_15800,N_15490);
nor U16561 (N_16561,N_15953,N_15872);
nor U16562 (N_16562,N_15612,N_15777);
nand U16563 (N_16563,N_15257,N_15846);
xnor U16564 (N_16564,N_15676,N_15064);
nor U16565 (N_16565,N_15396,N_15258);
or U16566 (N_16566,N_15429,N_15900);
nor U16567 (N_16567,N_15623,N_15825);
and U16568 (N_16568,N_15044,N_15163);
nor U16569 (N_16569,N_15540,N_15787);
and U16570 (N_16570,N_15373,N_15741);
and U16571 (N_16571,N_15043,N_15894);
and U16572 (N_16572,N_15501,N_15310);
or U16573 (N_16573,N_15036,N_15713);
nor U16574 (N_16574,N_15249,N_15509);
and U16575 (N_16575,N_15417,N_15650);
and U16576 (N_16576,N_15014,N_15438);
nand U16577 (N_16577,N_15731,N_15638);
nand U16578 (N_16578,N_15616,N_15218);
and U16579 (N_16579,N_15006,N_15056);
and U16580 (N_16580,N_15457,N_15381);
and U16581 (N_16581,N_15785,N_15798);
nand U16582 (N_16582,N_15461,N_15007);
and U16583 (N_16583,N_15105,N_15943);
and U16584 (N_16584,N_15340,N_15821);
and U16585 (N_16585,N_15400,N_15483);
or U16586 (N_16586,N_15298,N_15755);
xor U16587 (N_16587,N_15205,N_15711);
and U16588 (N_16588,N_15927,N_15748);
nand U16589 (N_16589,N_15981,N_15031);
nand U16590 (N_16590,N_15308,N_15171);
nand U16591 (N_16591,N_15992,N_15363);
or U16592 (N_16592,N_15847,N_15241);
or U16593 (N_16593,N_15783,N_15756);
or U16594 (N_16594,N_15860,N_15470);
xnor U16595 (N_16595,N_15171,N_15409);
nand U16596 (N_16596,N_15114,N_15592);
and U16597 (N_16597,N_15520,N_15061);
nor U16598 (N_16598,N_15199,N_15188);
and U16599 (N_16599,N_15637,N_15696);
or U16600 (N_16600,N_15211,N_15624);
nand U16601 (N_16601,N_15867,N_15796);
or U16602 (N_16602,N_15405,N_15553);
xor U16603 (N_16603,N_15690,N_15223);
nor U16604 (N_16604,N_15391,N_15358);
xnor U16605 (N_16605,N_15163,N_15430);
and U16606 (N_16606,N_15163,N_15264);
and U16607 (N_16607,N_15257,N_15325);
and U16608 (N_16608,N_15990,N_15705);
nand U16609 (N_16609,N_15950,N_15763);
xor U16610 (N_16610,N_15649,N_15430);
or U16611 (N_16611,N_15740,N_15115);
nand U16612 (N_16612,N_15441,N_15008);
or U16613 (N_16613,N_15488,N_15479);
or U16614 (N_16614,N_15429,N_15548);
or U16615 (N_16615,N_15662,N_15058);
nor U16616 (N_16616,N_15577,N_15220);
nor U16617 (N_16617,N_15439,N_15772);
xnor U16618 (N_16618,N_15896,N_15454);
and U16619 (N_16619,N_15573,N_15806);
nand U16620 (N_16620,N_15247,N_15714);
and U16621 (N_16621,N_15554,N_15851);
nor U16622 (N_16622,N_15016,N_15916);
or U16623 (N_16623,N_15964,N_15794);
or U16624 (N_16624,N_15561,N_15854);
xor U16625 (N_16625,N_15830,N_15912);
xnor U16626 (N_16626,N_15833,N_15037);
nor U16627 (N_16627,N_15855,N_15489);
xor U16628 (N_16628,N_15748,N_15233);
xor U16629 (N_16629,N_15795,N_15457);
nor U16630 (N_16630,N_15446,N_15155);
xor U16631 (N_16631,N_15436,N_15589);
and U16632 (N_16632,N_15475,N_15553);
and U16633 (N_16633,N_15336,N_15217);
xnor U16634 (N_16634,N_15407,N_15127);
or U16635 (N_16635,N_15157,N_15990);
or U16636 (N_16636,N_15801,N_15238);
xor U16637 (N_16637,N_15474,N_15075);
nor U16638 (N_16638,N_15968,N_15078);
xor U16639 (N_16639,N_15713,N_15270);
xor U16640 (N_16640,N_15518,N_15095);
nor U16641 (N_16641,N_15431,N_15844);
nand U16642 (N_16642,N_15700,N_15793);
nor U16643 (N_16643,N_15163,N_15507);
nor U16644 (N_16644,N_15235,N_15146);
nor U16645 (N_16645,N_15047,N_15614);
and U16646 (N_16646,N_15217,N_15874);
and U16647 (N_16647,N_15486,N_15750);
or U16648 (N_16648,N_15853,N_15517);
nand U16649 (N_16649,N_15112,N_15903);
or U16650 (N_16650,N_15720,N_15101);
xor U16651 (N_16651,N_15233,N_15989);
nor U16652 (N_16652,N_15612,N_15324);
nand U16653 (N_16653,N_15615,N_15198);
or U16654 (N_16654,N_15915,N_15781);
or U16655 (N_16655,N_15860,N_15193);
or U16656 (N_16656,N_15825,N_15482);
nand U16657 (N_16657,N_15367,N_15725);
xnor U16658 (N_16658,N_15072,N_15364);
or U16659 (N_16659,N_15667,N_15576);
xnor U16660 (N_16660,N_15625,N_15549);
nand U16661 (N_16661,N_15145,N_15860);
xnor U16662 (N_16662,N_15765,N_15335);
or U16663 (N_16663,N_15307,N_15400);
xnor U16664 (N_16664,N_15914,N_15514);
and U16665 (N_16665,N_15588,N_15395);
nand U16666 (N_16666,N_15141,N_15779);
and U16667 (N_16667,N_15623,N_15849);
xor U16668 (N_16668,N_15098,N_15767);
nor U16669 (N_16669,N_15254,N_15526);
or U16670 (N_16670,N_15279,N_15070);
xnor U16671 (N_16671,N_15214,N_15652);
nor U16672 (N_16672,N_15150,N_15758);
or U16673 (N_16673,N_15266,N_15898);
nand U16674 (N_16674,N_15381,N_15123);
and U16675 (N_16675,N_15253,N_15274);
or U16676 (N_16676,N_15360,N_15568);
nor U16677 (N_16677,N_15417,N_15973);
and U16678 (N_16678,N_15820,N_15942);
or U16679 (N_16679,N_15926,N_15082);
or U16680 (N_16680,N_15481,N_15489);
nand U16681 (N_16681,N_15963,N_15191);
nor U16682 (N_16682,N_15930,N_15688);
nor U16683 (N_16683,N_15069,N_15897);
or U16684 (N_16684,N_15316,N_15778);
and U16685 (N_16685,N_15052,N_15140);
and U16686 (N_16686,N_15249,N_15735);
and U16687 (N_16687,N_15228,N_15823);
xor U16688 (N_16688,N_15566,N_15236);
or U16689 (N_16689,N_15878,N_15192);
xnor U16690 (N_16690,N_15926,N_15977);
xnor U16691 (N_16691,N_15359,N_15901);
or U16692 (N_16692,N_15255,N_15836);
xnor U16693 (N_16693,N_15246,N_15171);
xor U16694 (N_16694,N_15273,N_15645);
or U16695 (N_16695,N_15707,N_15187);
and U16696 (N_16696,N_15142,N_15932);
nand U16697 (N_16697,N_15450,N_15667);
xnor U16698 (N_16698,N_15222,N_15550);
or U16699 (N_16699,N_15706,N_15830);
nand U16700 (N_16700,N_15614,N_15792);
xnor U16701 (N_16701,N_15237,N_15047);
xor U16702 (N_16702,N_15452,N_15032);
nand U16703 (N_16703,N_15314,N_15265);
and U16704 (N_16704,N_15365,N_15535);
nand U16705 (N_16705,N_15781,N_15323);
nand U16706 (N_16706,N_15740,N_15976);
or U16707 (N_16707,N_15274,N_15016);
and U16708 (N_16708,N_15867,N_15669);
xor U16709 (N_16709,N_15674,N_15657);
and U16710 (N_16710,N_15280,N_15077);
or U16711 (N_16711,N_15781,N_15356);
or U16712 (N_16712,N_15554,N_15453);
xor U16713 (N_16713,N_15330,N_15057);
nor U16714 (N_16714,N_15754,N_15334);
xnor U16715 (N_16715,N_15944,N_15715);
or U16716 (N_16716,N_15491,N_15358);
nor U16717 (N_16717,N_15441,N_15867);
nor U16718 (N_16718,N_15589,N_15794);
xor U16719 (N_16719,N_15892,N_15708);
and U16720 (N_16720,N_15163,N_15552);
nand U16721 (N_16721,N_15819,N_15814);
xor U16722 (N_16722,N_15948,N_15385);
nand U16723 (N_16723,N_15309,N_15776);
or U16724 (N_16724,N_15061,N_15590);
xnor U16725 (N_16725,N_15094,N_15547);
nand U16726 (N_16726,N_15792,N_15791);
or U16727 (N_16727,N_15150,N_15989);
nand U16728 (N_16728,N_15072,N_15583);
or U16729 (N_16729,N_15706,N_15316);
nor U16730 (N_16730,N_15601,N_15781);
and U16731 (N_16731,N_15475,N_15460);
nand U16732 (N_16732,N_15747,N_15621);
nor U16733 (N_16733,N_15136,N_15628);
or U16734 (N_16734,N_15647,N_15177);
xnor U16735 (N_16735,N_15540,N_15075);
or U16736 (N_16736,N_15531,N_15193);
or U16737 (N_16737,N_15503,N_15860);
nand U16738 (N_16738,N_15019,N_15478);
or U16739 (N_16739,N_15619,N_15970);
and U16740 (N_16740,N_15578,N_15024);
or U16741 (N_16741,N_15928,N_15568);
or U16742 (N_16742,N_15734,N_15394);
nand U16743 (N_16743,N_15134,N_15560);
nand U16744 (N_16744,N_15657,N_15846);
xor U16745 (N_16745,N_15889,N_15655);
nor U16746 (N_16746,N_15088,N_15173);
nand U16747 (N_16747,N_15092,N_15186);
nand U16748 (N_16748,N_15611,N_15127);
nor U16749 (N_16749,N_15585,N_15468);
nand U16750 (N_16750,N_15961,N_15918);
nand U16751 (N_16751,N_15149,N_15974);
xnor U16752 (N_16752,N_15493,N_15222);
nand U16753 (N_16753,N_15437,N_15480);
or U16754 (N_16754,N_15964,N_15475);
and U16755 (N_16755,N_15747,N_15817);
nor U16756 (N_16756,N_15580,N_15707);
and U16757 (N_16757,N_15503,N_15859);
xnor U16758 (N_16758,N_15780,N_15090);
nor U16759 (N_16759,N_15315,N_15005);
and U16760 (N_16760,N_15535,N_15417);
or U16761 (N_16761,N_15385,N_15774);
xor U16762 (N_16762,N_15100,N_15007);
nand U16763 (N_16763,N_15336,N_15308);
and U16764 (N_16764,N_15017,N_15185);
and U16765 (N_16765,N_15342,N_15549);
nand U16766 (N_16766,N_15183,N_15380);
nor U16767 (N_16767,N_15881,N_15905);
xnor U16768 (N_16768,N_15193,N_15753);
or U16769 (N_16769,N_15558,N_15123);
and U16770 (N_16770,N_15082,N_15017);
xor U16771 (N_16771,N_15093,N_15863);
nor U16772 (N_16772,N_15756,N_15340);
xnor U16773 (N_16773,N_15369,N_15033);
xor U16774 (N_16774,N_15134,N_15365);
nor U16775 (N_16775,N_15188,N_15762);
and U16776 (N_16776,N_15970,N_15259);
nor U16777 (N_16777,N_15964,N_15940);
nand U16778 (N_16778,N_15668,N_15262);
nand U16779 (N_16779,N_15111,N_15148);
xnor U16780 (N_16780,N_15995,N_15172);
and U16781 (N_16781,N_15291,N_15199);
xor U16782 (N_16782,N_15448,N_15422);
nor U16783 (N_16783,N_15983,N_15121);
nand U16784 (N_16784,N_15433,N_15921);
nand U16785 (N_16785,N_15076,N_15817);
nand U16786 (N_16786,N_15254,N_15255);
and U16787 (N_16787,N_15091,N_15640);
xor U16788 (N_16788,N_15200,N_15916);
or U16789 (N_16789,N_15284,N_15709);
xor U16790 (N_16790,N_15696,N_15203);
and U16791 (N_16791,N_15161,N_15620);
and U16792 (N_16792,N_15285,N_15681);
and U16793 (N_16793,N_15966,N_15302);
xnor U16794 (N_16794,N_15808,N_15626);
nor U16795 (N_16795,N_15569,N_15378);
and U16796 (N_16796,N_15332,N_15116);
xnor U16797 (N_16797,N_15516,N_15725);
or U16798 (N_16798,N_15456,N_15666);
nor U16799 (N_16799,N_15486,N_15759);
nor U16800 (N_16800,N_15017,N_15623);
nand U16801 (N_16801,N_15812,N_15702);
nand U16802 (N_16802,N_15924,N_15878);
nor U16803 (N_16803,N_15680,N_15545);
nor U16804 (N_16804,N_15539,N_15178);
nand U16805 (N_16805,N_15232,N_15867);
and U16806 (N_16806,N_15745,N_15652);
xor U16807 (N_16807,N_15823,N_15122);
xor U16808 (N_16808,N_15984,N_15761);
and U16809 (N_16809,N_15240,N_15638);
nand U16810 (N_16810,N_15429,N_15590);
nor U16811 (N_16811,N_15767,N_15941);
nor U16812 (N_16812,N_15690,N_15955);
nand U16813 (N_16813,N_15843,N_15385);
nor U16814 (N_16814,N_15896,N_15510);
nand U16815 (N_16815,N_15932,N_15496);
xor U16816 (N_16816,N_15022,N_15448);
or U16817 (N_16817,N_15996,N_15338);
nand U16818 (N_16818,N_15975,N_15904);
or U16819 (N_16819,N_15805,N_15034);
xor U16820 (N_16820,N_15752,N_15391);
nand U16821 (N_16821,N_15037,N_15360);
and U16822 (N_16822,N_15760,N_15220);
nor U16823 (N_16823,N_15845,N_15655);
xnor U16824 (N_16824,N_15085,N_15554);
xnor U16825 (N_16825,N_15718,N_15117);
nor U16826 (N_16826,N_15336,N_15216);
or U16827 (N_16827,N_15758,N_15352);
nand U16828 (N_16828,N_15435,N_15897);
nand U16829 (N_16829,N_15105,N_15591);
and U16830 (N_16830,N_15793,N_15464);
and U16831 (N_16831,N_15671,N_15567);
xor U16832 (N_16832,N_15000,N_15309);
and U16833 (N_16833,N_15261,N_15192);
nor U16834 (N_16834,N_15691,N_15574);
and U16835 (N_16835,N_15317,N_15400);
nor U16836 (N_16836,N_15017,N_15952);
nor U16837 (N_16837,N_15177,N_15200);
nand U16838 (N_16838,N_15965,N_15056);
and U16839 (N_16839,N_15168,N_15734);
and U16840 (N_16840,N_15842,N_15007);
nor U16841 (N_16841,N_15419,N_15906);
or U16842 (N_16842,N_15360,N_15428);
xor U16843 (N_16843,N_15736,N_15194);
nor U16844 (N_16844,N_15173,N_15255);
nand U16845 (N_16845,N_15093,N_15843);
xnor U16846 (N_16846,N_15687,N_15657);
nand U16847 (N_16847,N_15472,N_15257);
nor U16848 (N_16848,N_15647,N_15406);
nor U16849 (N_16849,N_15499,N_15206);
nand U16850 (N_16850,N_15196,N_15034);
and U16851 (N_16851,N_15128,N_15996);
and U16852 (N_16852,N_15688,N_15282);
or U16853 (N_16853,N_15683,N_15508);
and U16854 (N_16854,N_15825,N_15052);
xor U16855 (N_16855,N_15155,N_15180);
and U16856 (N_16856,N_15038,N_15134);
nor U16857 (N_16857,N_15066,N_15487);
and U16858 (N_16858,N_15591,N_15538);
and U16859 (N_16859,N_15727,N_15882);
or U16860 (N_16860,N_15966,N_15985);
or U16861 (N_16861,N_15563,N_15138);
or U16862 (N_16862,N_15039,N_15490);
nand U16863 (N_16863,N_15954,N_15197);
and U16864 (N_16864,N_15070,N_15199);
nand U16865 (N_16865,N_15916,N_15255);
or U16866 (N_16866,N_15045,N_15777);
nand U16867 (N_16867,N_15194,N_15652);
nor U16868 (N_16868,N_15416,N_15727);
xor U16869 (N_16869,N_15697,N_15565);
and U16870 (N_16870,N_15198,N_15271);
and U16871 (N_16871,N_15517,N_15315);
xnor U16872 (N_16872,N_15951,N_15768);
xnor U16873 (N_16873,N_15281,N_15168);
or U16874 (N_16874,N_15458,N_15724);
nand U16875 (N_16875,N_15807,N_15509);
xnor U16876 (N_16876,N_15023,N_15735);
nand U16877 (N_16877,N_15937,N_15354);
nor U16878 (N_16878,N_15996,N_15841);
or U16879 (N_16879,N_15423,N_15655);
or U16880 (N_16880,N_15586,N_15006);
nor U16881 (N_16881,N_15499,N_15465);
xnor U16882 (N_16882,N_15190,N_15841);
and U16883 (N_16883,N_15731,N_15323);
xor U16884 (N_16884,N_15047,N_15091);
nor U16885 (N_16885,N_15230,N_15301);
and U16886 (N_16886,N_15338,N_15079);
nor U16887 (N_16887,N_15821,N_15053);
or U16888 (N_16888,N_15448,N_15195);
or U16889 (N_16889,N_15033,N_15461);
or U16890 (N_16890,N_15101,N_15669);
nand U16891 (N_16891,N_15620,N_15879);
xor U16892 (N_16892,N_15613,N_15585);
nor U16893 (N_16893,N_15894,N_15163);
nor U16894 (N_16894,N_15661,N_15080);
nor U16895 (N_16895,N_15681,N_15253);
nand U16896 (N_16896,N_15294,N_15795);
and U16897 (N_16897,N_15346,N_15924);
and U16898 (N_16898,N_15337,N_15535);
or U16899 (N_16899,N_15060,N_15765);
nor U16900 (N_16900,N_15749,N_15255);
nand U16901 (N_16901,N_15688,N_15365);
or U16902 (N_16902,N_15596,N_15235);
nand U16903 (N_16903,N_15668,N_15882);
or U16904 (N_16904,N_15538,N_15068);
or U16905 (N_16905,N_15602,N_15092);
xnor U16906 (N_16906,N_15066,N_15466);
or U16907 (N_16907,N_15129,N_15934);
nand U16908 (N_16908,N_15872,N_15299);
or U16909 (N_16909,N_15511,N_15956);
nand U16910 (N_16910,N_15475,N_15774);
xnor U16911 (N_16911,N_15839,N_15366);
nand U16912 (N_16912,N_15741,N_15723);
xor U16913 (N_16913,N_15304,N_15836);
nand U16914 (N_16914,N_15984,N_15693);
nand U16915 (N_16915,N_15250,N_15899);
or U16916 (N_16916,N_15082,N_15855);
xnor U16917 (N_16917,N_15047,N_15846);
nor U16918 (N_16918,N_15251,N_15404);
or U16919 (N_16919,N_15356,N_15909);
or U16920 (N_16920,N_15917,N_15034);
or U16921 (N_16921,N_15679,N_15348);
nor U16922 (N_16922,N_15874,N_15868);
and U16923 (N_16923,N_15929,N_15852);
or U16924 (N_16924,N_15140,N_15074);
and U16925 (N_16925,N_15709,N_15184);
nand U16926 (N_16926,N_15143,N_15782);
and U16927 (N_16927,N_15951,N_15669);
xnor U16928 (N_16928,N_15708,N_15275);
or U16929 (N_16929,N_15901,N_15774);
or U16930 (N_16930,N_15759,N_15592);
and U16931 (N_16931,N_15810,N_15032);
and U16932 (N_16932,N_15440,N_15604);
nand U16933 (N_16933,N_15648,N_15881);
nand U16934 (N_16934,N_15821,N_15863);
nor U16935 (N_16935,N_15912,N_15803);
and U16936 (N_16936,N_15508,N_15457);
nor U16937 (N_16937,N_15009,N_15936);
nor U16938 (N_16938,N_15474,N_15777);
and U16939 (N_16939,N_15988,N_15483);
nand U16940 (N_16940,N_15144,N_15012);
or U16941 (N_16941,N_15533,N_15157);
nand U16942 (N_16942,N_15424,N_15973);
and U16943 (N_16943,N_15091,N_15578);
nor U16944 (N_16944,N_15361,N_15776);
and U16945 (N_16945,N_15302,N_15915);
or U16946 (N_16946,N_15943,N_15297);
nand U16947 (N_16947,N_15118,N_15135);
and U16948 (N_16948,N_15703,N_15443);
xor U16949 (N_16949,N_15072,N_15373);
nor U16950 (N_16950,N_15453,N_15416);
nor U16951 (N_16951,N_15064,N_15215);
or U16952 (N_16952,N_15172,N_15990);
nand U16953 (N_16953,N_15425,N_15400);
nand U16954 (N_16954,N_15921,N_15359);
nand U16955 (N_16955,N_15046,N_15399);
or U16956 (N_16956,N_15778,N_15344);
and U16957 (N_16957,N_15990,N_15253);
xnor U16958 (N_16958,N_15135,N_15307);
nor U16959 (N_16959,N_15838,N_15686);
xnor U16960 (N_16960,N_15099,N_15343);
xnor U16961 (N_16961,N_15770,N_15208);
and U16962 (N_16962,N_15806,N_15366);
and U16963 (N_16963,N_15137,N_15332);
or U16964 (N_16964,N_15197,N_15172);
or U16965 (N_16965,N_15614,N_15725);
nand U16966 (N_16966,N_15265,N_15136);
nand U16967 (N_16967,N_15213,N_15474);
nand U16968 (N_16968,N_15653,N_15342);
or U16969 (N_16969,N_15777,N_15627);
nand U16970 (N_16970,N_15981,N_15062);
or U16971 (N_16971,N_15993,N_15909);
nor U16972 (N_16972,N_15634,N_15379);
or U16973 (N_16973,N_15668,N_15905);
or U16974 (N_16974,N_15620,N_15818);
or U16975 (N_16975,N_15858,N_15623);
and U16976 (N_16976,N_15921,N_15089);
or U16977 (N_16977,N_15530,N_15963);
nor U16978 (N_16978,N_15307,N_15125);
nand U16979 (N_16979,N_15062,N_15074);
nor U16980 (N_16980,N_15902,N_15956);
nand U16981 (N_16981,N_15455,N_15831);
xor U16982 (N_16982,N_15297,N_15529);
xor U16983 (N_16983,N_15888,N_15311);
or U16984 (N_16984,N_15499,N_15637);
nor U16985 (N_16985,N_15488,N_15722);
nor U16986 (N_16986,N_15923,N_15460);
and U16987 (N_16987,N_15326,N_15590);
and U16988 (N_16988,N_15947,N_15410);
xor U16989 (N_16989,N_15238,N_15152);
xor U16990 (N_16990,N_15594,N_15589);
xnor U16991 (N_16991,N_15942,N_15526);
and U16992 (N_16992,N_15145,N_15510);
nand U16993 (N_16993,N_15511,N_15984);
nand U16994 (N_16994,N_15143,N_15529);
and U16995 (N_16995,N_15643,N_15506);
and U16996 (N_16996,N_15660,N_15789);
or U16997 (N_16997,N_15323,N_15245);
or U16998 (N_16998,N_15711,N_15844);
xor U16999 (N_16999,N_15251,N_15917);
and U17000 (N_17000,N_16392,N_16920);
and U17001 (N_17001,N_16004,N_16641);
nor U17002 (N_17002,N_16695,N_16944);
and U17003 (N_17003,N_16852,N_16908);
and U17004 (N_17004,N_16668,N_16999);
or U17005 (N_17005,N_16419,N_16138);
and U17006 (N_17006,N_16123,N_16888);
nand U17007 (N_17007,N_16163,N_16341);
nand U17008 (N_17008,N_16457,N_16555);
or U17009 (N_17009,N_16258,N_16070);
and U17010 (N_17010,N_16485,N_16318);
xor U17011 (N_17011,N_16152,N_16509);
and U17012 (N_17012,N_16882,N_16621);
nand U17013 (N_17013,N_16959,N_16887);
nor U17014 (N_17014,N_16569,N_16975);
or U17015 (N_17015,N_16722,N_16505);
nand U17016 (N_17016,N_16308,N_16415);
or U17017 (N_17017,N_16835,N_16907);
or U17018 (N_17018,N_16528,N_16733);
or U17019 (N_17019,N_16914,N_16370);
or U17020 (N_17020,N_16930,N_16469);
and U17021 (N_17021,N_16383,N_16616);
nand U17022 (N_17022,N_16105,N_16356);
or U17023 (N_17023,N_16165,N_16946);
and U17024 (N_17024,N_16497,N_16228);
xnor U17025 (N_17025,N_16149,N_16448);
xor U17026 (N_17026,N_16057,N_16359);
nor U17027 (N_17027,N_16285,N_16949);
or U17028 (N_17028,N_16250,N_16157);
xnor U17029 (N_17029,N_16752,N_16061);
xor U17030 (N_17030,N_16088,N_16186);
xnor U17031 (N_17031,N_16855,N_16310);
nand U17032 (N_17032,N_16282,N_16246);
and U17033 (N_17033,N_16340,N_16981);
nand U17034 (N_17034,N_16324,N_16515);
nor U17035 (N_17035,N_16588,N_16380);
nand U17036 (N_17036,N_16675,N_16235);
nor U17037 (N_17037,N_16772,N_16950);
xnor U17038 (N_17038,N_16169,N_16807);
xnor U17039 (N_17039,N_16886,N_16884);
nor U17040 (N_17040,N_16971,N_16982);
nand U17041 (N_17041,N_16510,N_16299);
nand U17042 (N_17042,N_16539,N_16756);
nand U17043 (N_17043,N_16550,N_16799);
and U17044 (N_17044,N_16312,N_16286);
or U17045 (N_17045,N_16470,N_16533);
nor U17046 (N_17046,N_16376,N_16050);
xnor U17047 (N_17047,N_16218,N_16594);
nor U17048 (N_17048,N_16990,N_16008);
nor U17049 (N_17049,N_16531,N_16630);
and U17050 (N_17050,N_16631,N_16798);
and U17051 (N_17051,N_16427,N_16435);
nand U17052 (N_17052,N_16489,N_16917);
or U17053 (N_17053,N_16601,N_16527);
xnor U17054 (N_17054,N_16034,N_16859);
nand U17055 (N_17055,N_16612,N_16922);
nor U17056 (N_17056,N_16552,N_16143);
and U17057 (N_17057,N_16978,N_16614);
nand U17058 (N_17058,N_16473,N_16900);
xor U17059 (N_17059,N_16877,N_16026);
nor U17060 (N_17060,N_16665,N_16049);
and U17061 (N_17061,N_16431,N_16170);
nand U17062 (N_17062,N_16710,N_16006);
xor U17063 (N_17063,N_16249,N_16248);
nand U17064 (N_17064,N_16503,N_16373);
and U17065 (N_17065,N_16844,N_16378);
xor U17066 (N_17066,N_16972,N_16754);
or U17067 (N_17067,N_16389,N_16232);
nor U17068 (N_17068,N_16110,N_16261);
or U17069 (N_17069,N_16629,N_16693);
and U17070 (N_17070,N_16150,N_16803);
nand U17071 (N_17071,N_16774,N_16748);
nor U17072 (N_17072,N_16192,N_16164);
or U17073 (N_17073,N_16092,N_16918);
or U17074 (N_17074,N_16116,N_16521);
or U17075 (N_17075,N_16390,N_16941);
or U17076 (N_17076,N_16176,N_16676);
or U17077 (N_17077,N_16739,N_16508);
or U17078 (N_17078,N_16610,N_16311);
and U17079 (N_17079,N_16190,N_16136);
nor U17080 (N_17080,N_16794,N_16266);
nor U17081 (N_17081,N_16534,N_16801);
nand U17082 (N_17082,N_16033,N_16275);
xor U17083 (N_17083,N_16649,N_16901);
nand U17084 (N_17084,N_16530,N_16768);
nor U17085 (N_17085,N_16016,N_16692);
and U17086 (N_17086,N_16837,N_16369);
xnor U17087 (N_17087,N_16706,N_16206);
nor U17088 (N_17088,N_16276,N_16828);
or U17089 (N_17089,N_16216,N_16051);
nor U17090 (N_17090,N_16581,N_16488);
nor U17091 (N_17091,N_16118,N_16065);
or U17092 (N_17092,N_16365,N_16921);
xnor U17093 (N_17093,N_16851,N_16055);
nand U17094 (N_17094,N_16411,N_16388);
xnor U17095 (N_17095,N_16556,N_16655);
or U17096 (N_17096,N_16000,N_16986);
nand U17097 (N_17097,N_16663,N_16291);
nand U17098 (N_17098,N_16168,N_16548);
xnor U17099 (N_17099,N_16547,N_16314);
nor U17100 (N_17100,N_16738,N_16181);
or U17101 (N_17101,N_16011,N_16934);
nand U17102 (N_17102,N_16073,N_16455);
nor U17103 (N_17103,N_16822,N_16728);
xor U17104 (N_17104,N_16862,N_16611);
and U17105 (N_17105,N_16545,N_16608);
nand U17106 (N_17106,N_16175,N_16333);
nand U17107 (N_17107,N_16513,N_16142);
nand U17108 (N_17108,N_16474,N_16234);
or U17109 (N_17109,N_16928,N_16028);
or U17110 (N_17110,N_16517,N_16148);
nand U17111 (N_17111,N_16074,N_16842);
and U17112 (N_17112,N_16865,N_16701);
nor U17113 (N_17113,N_16669,N_16770);
or U17114 (N_17114,N_16724,N_16736);
xor U17115 (N_17115,N_16323,N_16001);
nand U17116 (N_17116,N_16109,N_16410);
nand U17117 (N_17117,N_16654,N_16479);
and U17118 (N_17118,N_16953,N_16466);
and U17119 (N_17119,N_16656,N_16076);
or U17120 (N_17120,N_16082,N_16563);
nand U17121 (N_17121,N_16964,N_16054);
xnor U17122 (N_17122,N_16120,N_16788);
nand U17123 (N_17123,N_16367,N_16042);
and U17124 (N_17124,N_16281,N_16112);
nand U17125 (N_17125,N_16623,N_16477);
nand U17126 (N_17126,N_16989,N_16721);
or U17127 (N_17127,N_16607,N_16574);
or U17128 (N_17128,N_16771,N_16414);
nand U17129 (N_17129,N_16903,N_16155);
nor U17130 (N_17130,N_16892,N_16500);
and U17131 (N_17131,N_16624,N_16913);
xnor U17132 (N_17132,N_16845,N_16632);
nor U17133 (N_17133,N_16237,N_16178);
and U17134 (N_17134,N_16980,N_16832);
nand U17135 (N_17135,N_16587,N_16635);
nor U17136 (N_17136,N_16719,N_16296);
nor U17137 (N_17137,N_16287,N_16749);
or U17138 (N_17138,N_16328,N_16327);
and U17139 (N_17139,N_16247,N_16167);
and U17140 (N_17140,N_16685,N_16447);
nor U17141 (N_17141,N_16977,N_16151);
and U17142 (N_17142,N_16301,N_16452);
xnor U17143 (N_17143,N_16210,N_16336);
xor U17144 (N_17144,N_16751,N_16890);
nor U17145 (N_17145,N_16592,N_16189);
and U17146 (N_17146,N_16268,N_16344);
and U17147 (N_17147,N_16046,N_16360);
nor U17148 (N_17148,N_16429,N_16966);
nor U17149 (N_17149,N_16362,N_16478);
and U17150 (N_17150,N_16399,N_16915);
or U17151 (N_17151,N_16162,N_16638);
xor U17152 (N_17152,N_16764,N_16602);
nand U17153 (N_17153,N_16272,N_16127);
or U17154 (N_17154,N_16729,N_16916);
nand U17155 (N_17155,N_16860,N_16422);
or U17156 (N_17156,N_16948,N_16403);
xor U17157 (N_17157,N_16657,N_16830);
and U17158 (N_17158,N_16560,N_16716);
nand U17159 (N_17159,N_16677,N_16831);
nand U17160 (N_17160,N_16156,N_16577);
nand U17161 (N_17161,N_16511,N_16017);
or U17162 (N_17162,N_16240,N_16052);
nand U17163 (N_17163,N_16166,N_16618);
or U17164 (N_17164,N_16504,N_16955);
xnor U17165 (N_17165,N_16476,N_16124);
xnor U17166 (N_17166,N_16111,N_16827);
and U17167 (N_17167,N_16202,N_16086);
nor U17168 (N_17168,N_16361,N_16929);
nor U17169 (N_17169,N_16107,N_16651);
xnor U17170 (N_17170,N_16985,N_16071);
or U17171 (N_17171,N_16804,N_16967);
or U17172 (N_17172,N_16750,N_16535);
or U17173 (N_17173,N_16371,N_16699);
nor U17174 (N_17174,N_16861,N_16973);
xnor U17175 (N_17175,N_16122,N_16126);
and U17176 (N_17176,N_16713,N_16995);
nand U17177 (N_17177,N_16044,N_16209);
xor U17178 (N_17178,N_16683,N_16691);
nand U17179 (N_17179,N_16295,N_16544);
and U17180 (N_17180,N_16041,N_16348);
xor U17181 (N_17181,N_16108,N_16622);
nor U17182 (N_17182,N_16523,N_16096);
and U17183 (N_17183,N_16627,N_16245);
and U17184 (N_17184,N_16553,N_16117);
and U17185 (N_17185,N_16010,N_16613);
nand U17186 (N_17186,N_16334,N_16893);
xor U17187 (N_17187,N_16558,N_16666);
nor U17188 (N_17188,N_16525,N_16661);
nor U17189 (N_17189,N_16674,N_16141);
nor U17190 (N_17190,N_16696,N_16242);
xnor U17191 (N_17191,N_16625,N_16899);
nand U17192 (N_17192,N_16726,N_16889);
nand U17193 (N_17193,N_16895,N_16974);
xor U17194 (N_17194,N_16617,N_16251);
and U17195 (N_17195,N_16872,N_16075);
xor U17196 (N_17196,N_16820,N_16402);
xor U17197 (N_17197,N_16667,N_16300);
or U17198 (N_17198,N_16400,N_16912);
and U17199 (N_17199,N_16681,N_16717);
and U17200 (N_17200,N_16709,N_16450);
and U17201 (N_17201,N_16873,N_16896);
nand U17202 (N_17202,N_16812,N_16992);
xnor U17203 (N_17203,N_16220,N_16906);
nor U17204 (N_17204,N_16522,N_16227);
and U17205 (N_17205,N_16942,N_16321);
and U17206 (N_17206,N_16815,N_16083);
nor U17207 (N_17207,N_16064,N_16566);
nand U17208 (N_17208,N_16506,N_16104);
xnor U17209 (N_17209,N_16834,N_16923);
and U17210 (N_17210,N_16933,N_16062);
and U17211 (N_17211,N_16968,N_16306);
nand U17212 (N_17212,N_16174,N_16187);
or U17213 (N_17213,N_16097,N_16927);
nor U17214 (N_17214,N_16879,N_16813);
xor U17215 (N_17215,N_16711,N_16139);
and U17216 (N_17216,N_16874,N_16590);
and U17217 (N_17217,N_16221,N_16036);
xor U17218 (N_17218,N_16183,N_16605);
and U17219 (N_17219,N_16840,N_16956);
or U17220 (N_17220,N_16645,N_16686);
nand U17221 (N_17221,N_16542,N_16115);
nand U17222 (N_17222,N_16604,N_16319);
nor U17223 (N_17223,N_16012,N_16938);
xnor U17224 (N_17224,N_16351,N_16891);
xnor U17225 (N_17225,N_16332,N_16615);
and U17226 (N_17226,N_16278,N_16559);
nand U17227 (N_17227,N_16664,N_16003);
nor U17228 (N_17228,N_16264,N_16058);
nand U17229 (N_17229,N_16850,N_16983);
xnor U17230 (N_17230,N_16644,N_16829);
xnor U17231 (N_17231,N_16263,N_16121);
xnor U17232 (N_17232,N_16853,N_16407);
nor U17233 (N_17233,N_16072,N_16173);
nor U17234 (N_17234,N_16146,N_16129);
and U17235 (N_17235,N_16593,N_16269);
nand U17236 (N_17236,N_16442,N_16184);
nand U17237 (N_17237,N_16924,N_16274);
nor U17238 (N_17238,N_16459,N_16357);
and U17239 (N_17239,N_16628,N_16715);
or U17240 (N_17240,N_16180,N_16963);
nand U17241 (N_17241,N_16493,N_16087);
or U17242 (N_17242,N_16570,N_16395);
and U17243 (N_17243,N_16048,N_16401);
or U17244 (N_17244,N_16885,N_16626);
and U17245 (N_17245,N_16385,N_16440);
and U17246 (N_17246,N_16943,N_16773);
or U17247 (N_17247,N_16171,N_16763);
nor U17248 (N_17248,N_16598,N_16599);
or U17249 (N_17249,N_16067,N_16642);
nand U17250 (N_17250,N_16039,N_16222);
xor U17251 (N_17251,N_16498,N_16482);
and U17252 (N_17252,N_16991,N_16213);
or U17253 (N_17253,N_16894,N_16690);
and U17254 (N_17254,N_16355,N_16068);
nor U17255 (N_17255,N_16239,N_16059);
nand U17256 (N_17256,N_16911,N_16257);
or U17257 (N_17257,N_16185,N_16330);
xnor U17258 (N_17258,N_16468,N_16741);
nand U17259 (N_17259,N_16507,N_16653);
and U17260 (N_17260,N_16483,N_16066);
nor U17261 (N_17261,N_16433,N_16265);
and U17262 (N_17262,N_16791,N_16198);
nor U17263 (N_17263,N_16095,N_16684);
and U17264 (N_17264,N_16870,N_16304);
nor U17265 (N_17265,N_16494,N_16207);
xnor U17266 (N_17266,N_16743,N_16586);
or U17267 (N_17267,N_16777,N_16846);
xnor U17268 (N_17268,N_16810,N_16767);
or U17269 (N_17269,N_16014,N_16819);
nor U17270 (N_17270,N_16811,N_16796);
nor U17271 (N_17271,N_16514,N_16910);
xor U17272 (N_17272,N_16159,N_16761);
or U17273 (N_17273,N_16131,N_16776);
xor U17274 (N_17274,N_16343,N_16384);
xor U17275 (N_17275,N_16817,N_16765);
and U17276 (N_17276,N_16643,N_16406);
xor U17277 (N_17277,N_16769,N_16659);
xor U17278 (N_17278,N_16381,N_16289);
xor U17279 (N_17279,N_16345,N_16436);
and U17280 (N_17280,N_16808,N_16305);
nand U17281 (N_17281,N_16567,N_16783);
nor U17282 (N_17282,N_16905,N_16582);
nand U17283 (N_17283,N_16244,N_16600);
xor U17284 (N_17284,N_16718,N_16549);
nor U17285 (N_17285,N_16838,N_16491);
nand U17286 (N_17286,N_16680,N_16288);
nand U17287 (N_17287,N_16271,N_16571);
nor U17288 (N_17288,N_16465,N_16939);
nor U17289 (N_17289,N_16847,N_16866);
nor U17290 (N_17290,N_16671,N_16353);
and U17291 (N_17291,N_16596,N_16022);
nor U17292 (N_17292,N_16428,N_16597);
nor U17293 (N_17293,N_16572,N_16652);
xnor U17294 (N_17294,N_16080,N_16814);
or U17295 (N_17295,N_16755,N_16409);
nor U17296 (N_17296,N_16723,N_16426);
or U17297 (N_17297,N_16584,N_16694);
nor U17298 (N_17298,N_16009,N_16182);
nor U17299 (N_17299,N_16297,N_16194);
or U17300 (N_17300,N_16197,N_16160);
xnor U17301 (N_17301,N_16211,N_16416);
or U17302 (N_17302,N_16037,N_16988);
nor U17303 (N_17303,N_16688,N_16976);
nor U17304 (N_17304,N_16098,N_16637);
or U17305 (N_17305,N_16984,N_16200);
nor U17306 (N_17306,N_16658,N_16241);
nor U17307 (N_17307,N_16023,N_16077);
xnor U17308 (N_17308,N_16591,N_16703);
or U17309 (N_17309,N_16204,N_16698);
and U17310 (N_17310,N_16868,N_16821);
nand U17311 (N_17311,N_16780,N_16987);
and U17312 (N_17312,N_16425,N_16322);
nand U17313 (N_17313,N_16093,N_16382);
xor U17314 (N_17314,N_16205,N_16280);
nand U17315 (N_17315,N_16437,N_16573);
nand U17316 (N_17316,N_16565,N_16349);
xnor U17317 (N_17317,N_16779,N_16145);
and U17318 (N_17318,N_16329,N_16679);
nor U17319 (N_17319,N_16432,N_16284);
nand U17320 (N_17320,N_16737,N_16926);
xor U17321 (N_17321,N_16439,N_16270);
or U17322 (N_17322,N_16904,N_16201);
xor U17323 (N_17323,N_16960,N_16339);
or U17324 (N_17324,N_16215,N_16368);
or U17325 (N_17325,N_16824,N_16589);
xnor U17326 (N_17326,N_16687,N_16714);
and U17327 (N_17327,N_16226,N_16404);
and U17328 (N_17328,N_16255,N_16854);
nand U17329 (N_17329,N_16640,N_16826);
and U17330 (N_17330,N_16775,N_16208);
nand U17331 (N_17331,N_16759,N_16230);
nand U17332 (N_17332,N_16650,N_16158);
nand U17333 (N_17333,N_16540,N_16536);
or U17334 (N_17334,N_16229,N_16532);
nand U17335 (N_17335,N_16519,N_16945);
and U17336 (N_17336,N_16420,N_16753);
or U17337 (N_17337,N_16346,N_16467);
nor U17338 (N_17338,N_16393,N_16225);
and U17339 (N_17339,N_16848,N_16538);
and U17340 (N_17340,N_16841,N_16394);
or U17341 (N_17341,N_16858,N_16952);
and U17342 (N_17342,N_16518,N_16005);
xor U17343 (N_17343,N_16766,N_16697);
or U17344 (N_17344,N_16833,N_16546);
xor U17345 (N_17345,N_16620,N_16818);
nand U17346 (N_17346,N_16965,N_16994);
nand U17347 (N_17347,N_16372,N_16464);
nand U17348 (N_17348,N_16998,N_16609);
and U17349 (N_17349,N_16451,N_16352);
or U17350 (N_17350,N_16606,N_16704);
nand U17351 (N_17351,N_16418,N_16958);
nand U17352 (N_17352,N_16460,N_16293);
nor U17353 (N_17353,N_16458,N_16940);
and U17354 (N_17354,N_16326,N_16191);
nand U17355 (N_17355,N_16936,N_16662);
or U17356 (N_17356,N_16405,N_16454);
nor U17357 (N_17357,N_16516,N_16040);
nor U17358 (N_17358,N_16732,N_16060);
and U17359 (N_17359,N_16456,N_16475);
or U17360 (N_17360,N_16267,N_16734);
nand U17361 (N_17361,N_16782,N_16217);
nand U17362 (N_17362,N_16919,N_16744);
xnor U17363 (N_17363,N_16449,N_16670);
nor U17364 (N_17364,N_16849,N_16132);
and U17365 (N_17365,N_16702,N_16727);
and U17366 (N_17366,N_16233,N_16720);
nand U17367 (N_17367,N_16219,N_16196);
and U17368 (N_17368,N_16134,N_16747);
nand U17369 (N_17369,N_16883,N_16320);
nand U17370 (N_17370,N_16633,N_16678);
nand U17371 (N_17371,N_16337,N_16501);
or U17372 (N_17372,N_16094,N_16424);
nor U17373 (N_17373,N_16069,N_16199);
nand U17374 (N_17374,N_16954,N_16541);
and U17375 (N_17375,N_16292,N_16492);
and U17376 (N_17376,N_16935,N_16742);
and U17377 (N_17377,N_16932,N_16294);
nor U17378 (N_17378,N_16857,N_16133);
xnor U17379 (N_17379,N_16161,N_16091);
nand U17380 (N_17380,N_16785,N_16800);
xor U17381 (N_17381,N_16579,N_16839);
and U17382 (N_17382,N_16045,N_16583);
or U17383 (N_17383,N_16147,N_16979);
and U17384 (N_17384,N_16484,N_16135);
and U17385 (N_17385,N_16063,N_16902);
and U17386 (N_17386,N_16089,N_16002);
xnor U17387 (N_17387,N_16789,N_16363);
xor U17388 (N_17388,N_16947,N_16283);
and U17389 (N_17389,N_16490,N_16576);
or U17390 (N_17390,N_16561,N_16757);
or U17391 (N_17391,N_16792,N_16962);
nor U17392 (N_17392,N_16471,N_16793);
xor U17393 (N_17393,N_16195,N_16081);
or U17394 (N_17394,N_16997,N_16056);
nand U17395 (N_17395,N_16481,N_16636);
xor U17396 (N_17396,N_16880,N_16342);
nand U17397 (N_17397,N_16634,N_16347);
xor U17398 (N_17398,N_16412,N_16013);
nand U17399 (N_17399,N_16043,N_16580);
nor U17400 (N_17400,N_16961,N_16786);
nor U17401 (N_17401,N_16996,N_16103);
or U17402 (N_17402,N_16529,N_16931);
xor U17403 (N_17403,N_16438,N_16313);
or U17404 (N_17404,N_16027,N_16647);
or U17405 (N_17405,N_16787,N_16735);
nand U17406 (N_17406,N_16856,N_16188);
xnor U17407 (N_17407,N_16441,N_16878);
nor U17408 (N_17408,N_16020,N_16957);
nand U17409 (N_17409,N_16502,N_16795);
nand U17410 (N_17410,N_16863,N_16154);
or U17411 (N_17411,N_16397,N_16731);
nor U17412 (N_17412,N_16238,N_16700);
or U17413 (N_17413,N_16568,N_16252);
xnor U17414 (N_17414,N_16712,N_16867);
xor U17415 (N_17415,N_16038,N_16203);
or U17416 (N_17416,N_16937,N_16595);
or U17417 (N_17417,N_16524,N_16179);
and U17418 (N_17418,N_16350,N_16512);
nand U17419 (N_17419,N_16499,N_16639);
xnor U17420 (N_17420,N_16881,N_16090);
xor U17421 (N_17421,N_16708,N_16253);
nand U17422 (N_17422,N_16871,N_16100);
or U17423 (N_17423,N_16331,N_16029);
or U17424 (N_17424,N_16315,N_16256);
xor U17425 (N_17425,N_16030,N_16231);
nor U17426 (N_17426,N_16778,N_16366);
xor U17427 (N_17427,N_16487,N_16463);
xnor U17428 (N_17428,N_16797,N_16223);
xnor U17429 (N_17429,N_16021,N_16140);
and U17430 (N_17430,N_16836,N_16969);
nor U17431 (N_17431,N_16480,N_16543);
xnor U17432 (N_17432,N_16137,N_16085);
nand U17433 (N_17433,N_16106,N_16099);
or U17434 (N_17434,N_16254,N_16031);
nand U17435 (N_17435,N_16259,N_16303);
or U17436 (N_17436,N_16375,N_16018);
xor U17437 (N_17437,N_16307,N_16130);
nor U17438 (N_17438,N_16472,N_16078);
or U17439 (N_17439,N_16260,N_16575);
nor U17440 (N_17440,N_16102,N_16745);
nand U17441 (N_17441,N_16386,N_16354);
nand U17442 (N_17442,N_16379,N_16876);
and U17443 (N_17443,N_16809,N_16648);
or U17444 (N_17444,N_16781,N_16338);
nand U17445 (N_17445,N_16153,N_16423);
or U17446 (N_17446,N_16551,N_16740);
and U17447 (N_17447,N_16128,N_16843);
nand U17448 (N_17448,N_16298,N_16408);
and U17449 (N_17449,N_16125,N_16434);
nand U17450 (N_17450,N_16015,N_16790);
nand U17451 (N_17451,N_16290,N_16970);
nand U17452 (N_17452,N_16909,N_16316);
xnor U17453 (N_17453,N_16993,N_16461);
xnor U17454 (N_17454,N_16825,N_16214);
or U17455 (N_17455,N_16391,N_16746);
nand U17456 (N_17456,N_16619,N_16084);
or U17457 (N_17457,N_16398,N_16898);
or U17458 (N_17458,N_16725,N_16421);
nor U17459 (N_17459,N_16374,N_16212);
nand U17460 (N_17460,N_16025,N_16007);
xnor U17461 (N_17461,N_16453,N_16302);
xor U17462 (N_17462,N_16486,N_16557);
nor U17463 (N_17463,N_16672,N_16047);
nand U17464 (N_17464,N_16562,N_16177);
or U17465 (N_17465,N_16119,N_16114);
or U17466 (N_17466,N_16526,N_16364);
and U17467 (N_17467,N_16413,N_16762);
xor U17468 (N_17468,N_16279,N_16236);
nor U17469 (N_17469,N_16273,N_16032);
nand U17470 (N_17470,N_16446,N_16869);
nor U17471 (N_17471,N_16224,N_16578);
and U17472 (N_17472,N_16443,N_16806);
nor U17473 (N_17473,N_16660,N_16603);
and U17474 (N_17474,N_16358,N_16823);
nand U17475 (N_17475,N_16396,N_16193);
nor U17476 (N_17476,N_16730,N_16805);
or U17477 (N_17477,N_16113,N_16277);
or U17478 (N_17478,N_16325,N_16564);
and U17479 (N_17479,N_16335,N_16758);
xnor U17480 (N_17480,N_16784,N_16445);
or U17481 (N_17481,N_16144,N_16243);
or U17482 (N_17482,N_16520,N_16897);
or U17483 (N_17483,N_16689,N_16101);
nand U17484 (N_17484,N_16760,N_16554);
or U17485 (N_17485,N_16875,N_16705);
or U17486 (N_17486,N_16646,N_16462);
or U17487 (N_17487,N_16585,N_16673);
or U17488 (N_17488,N_16444,N_16802);
and U17489 (N_17489,N_16387,N_16707);
and U17490 (N_17490,N_16816,N_16925);
or U17491 (N_17491,N_16430,N_16537);
or U17492 (N_17492,N_16172,N_16079);
nand U17493 (N_17493,N_16262,N_16035);
and U17494 (N_17494,N_16864,N_16309);
nor U17495 (N_17495,N_16377,N_16682);
nor U17496 (N_17496,N_16024,N_16496);
nor U17497 (N_17497,N_16317,N_16951);
nor U17498 (N_17498,N_16053,N_16019);
nand U17499 (N_17499,N_16417,N_16495);
xor U17500 (N_17500,N_16622,N_16386);
xor U17501 (N_17501,N_16304,N_16840);
xor U17502 (N_17502,N_16759,N_16155);
nand U17503 (N_17503,N_16581,N_16105);
and U17504 (N_17504,N_16122,N_16098);
xor U17505 (N_17505,N_16962,N_16541);
and U17506 (N_17506,N_16826,N_16340);
and U17507 (N_17507,N_16519,N_16365);
nand U17508 (N_17508,N_16728,N_16422);
or U17509 (N_17509,N_16045,N_16085);
nor U17510 (N_17510,N_16366,N_16684);
and U17511 (N_17511,N_16948,N_16610);
nand U17512 (N_17512,N_16600,N_16314);
xor U17513 (N_17513,N_16569,N_16598);
xnor U17514 (N_17514,N_16540,N_16571);
nand U17515 (N_17515,N_16475,N_16767);
and U17516 (N_17516,N_16755,N_16186);
nor U17517 (N_17517,N_16413,N_16889);
nor U17518 (N_17518,N_16757,N_16766);
xor U17519 (N_17519,N_16238,N_16699);
xnor U17520 (N_17520,N_16272,N_16417);
and U17521 (N_17521,N_16608,N_16229);
nand U17522 (N_17522,N_16320,N_16835);
and U17523 (N_17523,N_16568,N_16576);
nand U17524 (N_17524,N_16305,N_16474);
nor U17525 (N_17525,N_16067,N_16428);
nor U17526 (N_17526,N_16481,N_16008);
nand U17527 (N_17527,N_16251,N_16161);
xnor U17528 (N_17528,N_16719,N_16304);
nand U17529 (N_17529,N_16582,N_16510);
or U17530 (N_17530,N_16893,N_16818);
nand U17531 (N_17531,N_16165,N_16155);
and U17532 (N_17532,N_16705,N_16057);
nor U17533 (N_17533,N_16631,N_16482);
nand U17534 (N_17534,N_16052,N_16537);
nand U17535 (N_17535,N_16047,N_16830);
nand U17536 (N_17536,N_16950,N_16842);
nand U17537 (N_17537,N_16302,N_16257);
and U17538 (N_17538,N_16429,N_16250);
or U17539 (N_17539,N_16735,N_16605);
or U17540 (N_17540,N_16527,N_16137);
nor U17541 (N_17541,N_16797,N_16241);
and U17542 (N_17542,N_16218,N_16758);
nand U17543 (N_17543,N_16508,N_16230);
or U17544 (N_17544,N_16048,N_16762);
xor U17545 (N_17545,N_16800,N_16313);
nand U17546 (N_17546,N_16851,N_16511);
or U17547 (N_17547,N_16799,N_16939);
nand U17548 (N_17548,N_16578,N_16044);
or U17549 (N_17549,N_16243,N_16792);
nor U17550 (N_17550,N_16441,N_16059);
nor U17551 (N_17551,N_16376,N_16553);
and U17552 (N_17552,N_16737,N_16413);
or U17553 (N_17553,N_16795,N_16586);
or U17554 (N_17554,N_16637,N_16163);
and U17555 (N_17555,N_16903,N_16168);
nand U17556 (N_17556,N_16452,N_16927);
nand U17557 (N_17557,N_16089,N_16618);
or U17558 (N_17558,N_16041,N_16872);
and U17559 (N_17559,N_16392,N_16223);
or U17560 (N_17560,N_16549,N_16958);
xnor U17561 (N_17561,N_16819,N_16896);
or U17562 (N_17562,N_16603,N_16938);
and U17563 (N_17563,N_16912,N_16225);
nor U17564 (N_17564,N_16382,N_16880);
nand U17565 (N_17565,N_16236,N_16764);
nand U17566 (N_17566,N_16217,N_16807);
nor U17567 (N_17567,N_16191,N_16134);
nand U17568 (N_17568,N_16596,N_16355);
or U17569 (N_17569,N_16406,N_16715);
xor U17570 (N_17570,N_16520,N_16926);
nand U17571 (N_17571,N_16220,N_16429);
nand U17572 (N_17572,N_16549,N_16910);
xnor U17573 (N_17573,N_16644,N_16134);
nor U17574 (N_17574,N_16750,N_16662);
or U17575 (N_17575,N_16375,N_16439);
or U17576 (N_17576,N_16807,N_16575);
nand U17577 (N_17577,N_16891,N_16504);
xnor U17578 (N_17578,N_16486,N_16564);
and U17579 (N_17579,N_16904,N_16736);
nor U17580 (N_17580,N_16635,N_16063);
nand U17581 (N_17581,N_16071,N_16061);
xnor U17582 (N_17582,N_16452,N_16273);
nor U17583 (N_17583,N_16673,N_16331);
or U17584 (N_17584,N_16845,N_16491);
xor U17585 (N_17585,N_16478,N_16253);
nor U17586 (N_17586,N_16891,N_16988);
and U17587 (N_17587,N_16338,N_16233);
and U17588 (N_17588,N_16334,N_16553);
and U17589 (N_17589,N_16385,N_16711);
xnor U17590 (N_17590,N_16465,N_16405);
xor U17591 (N_17591,N_16663,N_16596);
nor U17592 (N_17592,N_16333,N_16625);
or U17593 (N_17593,N_16944,N_16216);
or U17594 (N_17594,N_16271,N_16658);
nand U17595 (N_17595,N_16074,N_16966);
xor U17596 (N_17596,N_16408,N_16770);
nand U17597 (N_17597,N_16522,N_16966);
and U17598 (N_17598,N_16816,N_16860);
and U17599 (N_17599,N_16520,N_16332);
and U17600 (N_17600,N_16333,N_16543);
xor U17601 (N_17601,N_16516,N_16913);
nand U17602 (N_17602,N_16301,N_16767);
or U17603 (N_17603,N_16336,N_16207);
or U17604 (N_17604,N_16274,N_16392);
or U17605 (N_17605,N_16595,N_16699);
nand U17606 (N_17606,N_16306,N_16254);
and U17607 (N_17607,N_16824,N_16190);
nor U17608 (N_17608,N_16034,N_16750);
or U17609 (N_17609,N_16586,N_16702);
xnor U17610 (N_17610,N_16148,N_16357);
xnor U17611 (N_17611,N_16643,N_16020);
xnor U17612 (N_17612,N_16037,N_16917);
xnor U17613 (N_17613,N_16119,N_16664);
or U17614 (N_17614,N_16662,N_16370);
nand U17615 (N_17615,N_16046,N_16616);
and U17616 (N_17616,N_16466,N_16174);
or U17617 (N_17617,N_16209,N_16580);
xor U17618 (N_17618,N_16784,N_16980);
or U17619 (N_17619,N_16946,N_16261);
nor U17620 (N_17620,N_16540,N_16208);
or U17621 (N_17621,N_16976,N_16846);
nand U17622 (N_17622,N_16304,N_16369);
nand U17623 (N_17623,N_16092,N_16699);
or U17624 (N_17624,N_16154,N_16829);
or U17625 (N_17625,N_16134,N_16057);
and U17626 (N_17626,N_16493,N_16301);
nand U17627 (N_17627,N_16761,N_16645);
or U17628 (N_17628,N_16722,N_16970);
or U17629 (N_17629,N_16317,N_16514);
and U17630 (N_17630,N_16485,N_16330);
nor U17631 (N_17631,N_16706,N_16167);
and U17632 (N_17632,N_16484,N_16477);
nand U17633 (N_17633,N_16559,N_16522);
or U17634 (N_17634,N_16004,N_16326);
nand U17635 (N_17635,N_16768,N_16597);
xor U17636 (N_17636,N_16555,N_16915);
nor U17637 (N_17637,N_16847,N_16475);
nand U17638 (N_17638,N_16835,N_16986);
nor U17639 (N_17639,N_16713,N_16407);
or U17640 (N_17640,N_16456,N_16979);
or U17641 (N_17641,N_16090,N_16222);
and U17642 (N_17642,N_16658,N_16155);
nor U17643 (N_17643,N_16846,N_16212);
nor U17644 (N_17644,N_16022,N_16176);
and U17645 (N_17645,N_16646,N_16365);
nor U17646 (N_17646,N_16796,N_16849);
or U17647 (N_17647,N_16555,N_16381);
xnor U17648 (N_17648,N_16106,N_16782);
or U17649 (N_17649,N_16232,N_16618);
nand U17650 (N_17650,N_16405,N_16794);
nand U17651 (N_17651,N_16880,N_16114);
and U17652 (N_17652,N_16849,N_16664);
nor U17653 (N_17653,N_16112,N_16873);
or U17654 (N_17654,N_16065,N_16479);
xnor U17655 (N_17655,N_16257,N_16110);
nor U17656 (N_17656,N_16705,N_16213);
and U17657 (N_17657,N_16770,N_16170);
nor U17658 (N_17658,N_16395,N_16072);
nand U17659 (N_17659,N_16788,N_16093);
or U17660 (N_17660,N_16510,N_16883);
or U17661 (N_17661,N_16879,N_16618);
and U17662 (N_17662,N_16503,N_16434);
xnor U17663 (N_17663,N_16025,N_16050);
nor U17664 (N_17664,N_16713,N_16913);
xnor U17665 (N_17665,N_16758,N_16454);
or U17666 (N_17666,N_16168,N_16783);
xnor U17667 (N_17667,N_16722,N_16621);
or U17668 (N_17668,N_16673,N_16724);
and U17669 (N_17669,N_16109,N_16048);
xor U17670 (N_17670,N_16284,N_16057);
nor U17671 (N_17671,N_16512,N_16242);
or U17672 (N_17672,N_16461,N_16032);
nand U17673 (N_17673,N_16734,N_16477);
and U17674 (N_17674,N_16771,N_16755);
nand U17675 (N_17675,N_16471,N_16183);
xor U17676 (N_17676,N_16935,N_16462);
nand U17677 (N_17677,N_16784,N_16249);
nor U17678 (N_17678,N_16142,N_16100);
nor U17679 (N_17679,N_16408,N_16294);
and U17680 (N_17680,N_16705,N_16855);
xnor U17681 (N_17681,N_16548,N_16452);
xor U17682 (N_17682,N_16519,N_16093);
nand U17683 (N_17683,N_16344,N_16658);
nand U17684 (N_17684,N_16458,N_16948);
nand U17685 (N_17685,N_16503,N_16141);
and U17686 (N_17686,N_16624,N_16915);
nor U17687 (N_17687,N_16654,N_16275);
xnor U17688 (N_17688,N_16409,N_16797);
nand U17689 (N_17689,N_16765,N_16625);
xor U17690 (N_17690,N_16637,N_16310);
xnor U17691 (N_17691,N_16526,N_16389);
or U17692 (N_17692,N_16989,N_16052);
xor U17693 (N_17693,N_16716,N_16798);
nand U17694 (N_17694,N_16178,N_16442);
xnor U17695 (N_17695,N_16827,N_16727);
xor U17696 (N_17696,N_16668,N_16937);
nand U17697 (N_17697,N_16649,N_16436);
nand U17698 (N_17698,N_16884,N_16532);
nor U17699 (N_17699,N_16988,N_16527);
xor U17700 (N_17700,N_16133,N_16432);
xnor U17701 (N_17701,N_16827,N_16492);
nand U17702 (N_17702,N_16300,N_16355);
or U17703 (N_17703,N_16139,N_16082);
nand U17704 (N_17704,N_16399,N_16808);
nand U17705 (N_17705,N_16562,N_16694);
xnor U17706 (N_17706,N_16940,N_16530);
nand U17707 (N_17707,N_16622,N_16252);
nor U17708 (N_17708,N_16612,N_16204);
nand U17709 (N_17709,N_16560,N_16659);
nor U17710 (N_17710,N_16800,N_16346);
nor U17711 (N_17711,N_16514,N_16935);
and U17712 (N_17712,N_16542,N_16140);
nor U17713 (N_17713,N_16206,N_16109);
or U17714 (N_17714,N_16235,N_16880);
or U17715 (N_17715,N_16594,N_16724);
and U17716 (N_17716,N_16614,N_16608);
and U17717 (N_17717,N_16671,N_16134);
and U17718 (N_17718,N_16446,N_16738);
nand U17719 (N_17719,N_16854,N_16055);
and U17720 (N_17720,N_16297,N_16977);
and U17721 (N_17721,N_16189,N_16573);
xor U17722 (N_17722,N_16655,N_16981);
and U17723 (N_17723,N_16580,N_16587);
and U17724 (N_17724,N_16650,N_16135);
nand U17725 (N_17725,N_16321,N_16661);
or U17726 (N_17726,N_16951,N_16692);
nand U17727 (N_17727,N_16816,N_16650);
nand U17728 (N_17728,N_16764,N_16962);
nand U17729 (N_17729,N_16327,N_16057);
nor U17730 (N_17730,N_16929,N_16996);
or U17731 (N_17731,N_16082,N_16485);
nor U17732 (N_17732,N_16582,N_16406);
nor U17733 (N_17733,N_16471,N_16725);
xor U17734 (N_17734,N_16147,N_16380);
xnor U17735 (N_17735,N_16514,N_16594);
xor U17736 (N_17736,N_16359,N_16984);
xor U17737 (N_17737,N_16105,N_16656);
or U17738 (N_17738,N_16715,N_16268);
and U17739 (N_17739,N_16063,N_16908);
nor U17740 (N_17740,N_16529,N_16120);
nand U17741 (N_17741,N_16192,N_16298);
or U17742 (N_17742,N_16582,N_16010);
nor U17743 (N_17743,N_16049,N_16646);
nor U17744 (N_17744,N_16107,N_16611);
nand U17745 (N_17745,N_16076,N_16284);
or U17746 (N_17746,N_16334,N_16442);
nand U17747 (N_17747,N_16389,N_16572);
nor U17748 (N_17748,N_16612,N_16964);
nand U17749 (N_17749,N_16385,N_16175);
or U17750 (N_17750,N_16549,N_16231);
or U17751 (N_17751,N_16547,N_16470);
nand U17752 (N_17752,N_16527,N_16870);
or U17753 (N_17753,N_16637,N_16222);
and U17754 (N_17754,N_16763,N_16257);
xnor U17755 (N_17755,N_16995,N_16108);
nor U17756 (N_17756,N_16853,N_16446);
or U17757 (N_17757,N_16200,N_16433);
nand U17758 (N_17758,N_16161,N_16424);
xor U17759 (N_17759,N_16264,N_16518);
and U17760 (N_17760,N_16319,N_16536);
nor U17761 (N_17761,N_16055,N_16931);
nand U17762 (N_17762,N_16045,N_16366);
nand U17763 (N_17763,N_16162,N_16673);
nor U17764 (N_17764,N_16908,N_16596);
and U17765 (N_17765,N_16464,N_16701);
and U17766 (N_17766,N_16025,N_16435);
or U17767 (N_17767,N_16510,N_16974);
nand U17768 (N_17768,N_16486,N_16791);
nand U17769 (N_17769,N_16750,N_16475);
nor U17770 (N_17770,N_16130,N_16784);
nor U17771 (N_17771,N_16492,N_16945);
nand U17772 (N_17772,N_16557,N_16592);
xor U17773 (N_17773,N_16634,N_16197);
nor U17774 (N_17774,N_16433,N_16567);
or U17775 (N_17775,N_16501,N_16880);
nor U17776 (N_17776,N_16750,N_16098);
xnor U17777 (N_17777,N_16686,N_16613);
nor U17778 (N_17778,N_16882,N_16952);
xor U17779 (N_17779,N_16383,N_16805);
nor U17780 (N_17780,N_16207,N_16102);
nand U17781 (N_17781,N_16482,N_16355);
nand U17782 (N_17782,N_16087,N_16432);
or U17783 (N_17783,N_16638,N_16255);
xor U17784 (N_17784,N_16975,N_16748);
nand U17785 (N_17785,N_16365,N_16170);
and U17786 (N_17786,N_16421,N_16712);
or U17787 (N_17787,N_16083,N_16995);
and U17788 (N_17788,N_16402,N_16702);
or U17789 (N_17789,N_16590,N_16009);
nor U17790 (N_17790,N_16446,N_16384);
nor U17791 (N_17791,N_16970,N_16993);
and U17792 (N_17792,N_16932,N_16961);
and U17793 (N_17793,N_16292,N_16241);
xor U17794 (N_17794,N_16652,N_16171);
nor U17795 (N_17795,N_16584,N_16013);
xor U17796 (N_17796,N_16570,N_16782);
nor U17797 (N_17797,N_16248,N_16324);
nor U17798 (N_17798,N_16261,N_16183);
nor U17799 (N_17799,N_16834,N_16841);
xor U17800 (N_17800,N_16083,N_16525);
xnor U17801 (N_17801,N_16631,N_16057);
nor U17802 (N_17802,N_16739,N_16544);
nand U17803 (N_17803,N_16269,N_16678);
nand U17804 (N_17804,N_16223,N_16558);
nor U17805 (N_17805,N_16561,N_16688);
and U17806 (N_17806,N_16135,N_16162);
and U17807 (N_17807,N_16715,N_16174);
xor U17808 (N_17808,N_16257,N_16999);
nand U17809 (N_17809,N_16949,N_16092);
nor U17810 (N_17810,N_16497,N_16836);
or U17811 (N_17811,N_16516,N_16139);
xor U17812 (N_17812,N_16002,N_16583);
xnor U17813 (N_17813,N_16731,N_16349);
xnor U17814 (N_17814,N_16832,N_16611);
or U17815 (N_17815,N_16774,N_16131);
xnor U17816 (N_17816,N_16599,N_16221);
nor U17817 (N_17817,N_16118,N_16589);
xor U17818 (N_17818,N_16094,N_16456);
nand U17819 (N_17819,N_16165,N_16504);
nor U17820 (N_17820,N_16279,N_16030);
xor U17821 (N_17821,N_16641,N_16770);
and U17822 (N_17822,N_16617,N_16525);
xor U17823 (N_17823,N_16541,N_16130);
or U17824 (N_17824,N_16851,N_16380);
nor U17825 (N_17825,N_16607,N_16077);
and U17826 (N_17826,N_16248,N_16238);
nand U17827 (N_17827,N_16139,N_16653);
or U17828 (N_17828,N_16569,N_16682);
and U17829 (N_17829,N_16253,N_16385);
or U17830 (N_17830,N_16391,N_16563);
xnor U17831 (N_17831,N_16563,N_16777);
nand U17832 (N_17832,N_16845,N_16584);
xor U17833 (N_17833,N_16316,N_16346);
or U17834 (N_17834,N_16054,N_16265);
and U17835 (N_17835,N_16719,N_16503);
nor U17836 (N_17836,N_16689,N_16168);
xor U17837 (N_17837,N_16252,N_16197);
or U17838 (N_17838,N_16460,N_16410);
xnor U17839 (N_17839,N_16464,N_16271);
nor U17840 (N_17840,N_16411,N_16895);
nor U17841 (N_17841,N_16511,N_16991);
nor U17842 (N_17842,N_16851,N_16708);
or U17843 (N_17843,N_16342,N_16390);
or U17844 (N_17844,N_16616,N_16392);
nor U17845 (N_17845,N_16133,N_16990);
nor U17846 (N_17846,N_16464,N_16532);
and U17847 (N_17847,N_16000,N_16489);
nand U17848 (N_17848,N_16637,N_16192);
and U17849 (N_17849,N_16411,N_16119);
nand U17850 (N_17850,N_16631,N_16756);
nand U17851 (N_17851,N_16556,N_16758);
and U17852 (N_17852,N_16673,N_16276);
and U17853 (N_17853,N_16714,N_16832);
nand U17854 (N_17854,N_16640,N_16945);
xnor U17855 (N_17855,N_16545,N_16758);
or U17856 (N_17856,N_16331,N_16511);
and U17857 (N_17857,N_16065,N_16623);
nor U17858 (N_17858,N_16837,N_16157);
and U17859 (N_17859,N_16242,N_16594);
nor U17860 (N_17860,N_16361,N_16625);
nor U17861 (N_17861,N_16778,N_16176);
and U17862 (N_17862,N_16533,N_16365);
xnor U17863 (N_17863,N_16640,N_16064);
and U17864 (N_17864,N_16094,N_16239);
or U17865 (N_17865,N_16262,N_16419);
or U17866 (N_17866,N_16635,N_16607);
xnor U17867 (N_17867,N_16507,N_16099);
or U17868 (N_17868,N_16132,N_16261);
nor U17869 (N_17869,N_16471,N_16739);
or U17870 (N_17870,N_16223,N_16019);
and U17871 (N_17871,N_16541,N_16075);
nand U17872 (N_17872,N_16058,N_16190);
nand U17873 (N_17873,N_16700,N_16054);
and U17874 (N_17874,N_16571,N_16618);
or U17875 (N_17875,N_16270,N_16448);
and U17876 (N_17876,N_16993,N_16634);
and U17877 (N_17877,N_16609,N_16449);
or U17878 (N_17878,N_16591,N_16169);
and U17879 (N_17879,N_16969,N_16048);
xor U17880 (N_17880,N_16284,N_16105);
nand U17881 (N_17881,N_16473,N_16831);
nor U17882 (N_17882,N_16622,N_16681);
xor U17883 (N_17883,N_16707,N_16489);
xnor U17884 (N_17884,N_16807,N_16266);
xor U17885 (N_17885,N_16330,N_16044);
or U17886 (N_17886,N_16697,N_16738);
and U17887 (N_17887,N_16382,N_16516);
xor U17888 (N_17888,N_16487,N_16493);
xnor U17889 (N_17889,N_16847,N_16262);
nor U17890 (N_17890,N_16210,N_16872);
or U17891 (N_17891,N_16221,N_16391);
nand U17892 (N_17892,N_16382,N_16634);
xor U17893 (N_17893,N_16678,N_16331);
nor U17894 (N_17894,N_16811,N_16319);
nor U17895 (N_17895,N_16936,N_16294);
nand U17896 (N_17896,N_16387,N_16044);
and U17897 (N_17897,N_16738,N_16002);
nand U17898 (N_17898,N_16520,N_16477);
nor U17899 (N_17899,N_16585,N_16995);
nand U17900 (N_17900,N_16251,N_16126);
and U17901 (N_17901,N_16097,N_16461);
and U17902 (N_17902,N_16592,N_16864);
and U17903 (N_17903,N_16474,N_16650);
nand U17904 (N_17904,N_16395,N_16966);
nor U17905 (N_17905,N_16032,N_16745);
or U17906 (N_17906,N_16778,N_16812);
nand U17907 (N_17907,N_16087,N_16186);
xnor U17908 (N_17908,N_16176,N_16715);
or U17909 (N_17909,N_16356,N_16468);
nand U17910 (N_17910,N_16828,N_16809);
or U17911 (N_17911,N_16603,N_16908);
and U17912 (N_17912,N_16715,N_16769);
nand U17913 (N_17913,N_16825,N_16347);
and U17914 (N_17914,N_16708,N_16413);
nor U17915 (N_17915,N_16030,N_16260);
xnor U17916 (N_17916,N_16635,N_16313);
xor U17917 (N_17917,N_16083,N_16701);
or U17918 (N_17918,N_16741,N_16094);
nand U17919 (N_17919,N_16621,N_16659);
and U17920 (N_17920,N_16875,N_16151);
nand U17921 (N_17921,N_16315,N_16680);
xor U17922 (N_17922,N_16117,N_16445);
nand U17923 (N_17923,N_16344,N_16241);
nand U17924 (N_17924,N_16885,N_16406);
xor U17925 (N_17925,N_16870,N_16947);
nand U17926 (N_17926,N_16628,N_16165);
and U17927 (N_17927,N_16128,N_16493);
or U17928 (N_17928,N_16105,N_16802);
nand U17929 (N_17929,N_16686,N_16085);
nand U17930 (N_17930,N_16550,N_16978);
nor U17931 (N_17931,N_16370,N_16468);
nand U17932 (N_17932,N_16116,N_16761);
and U17933 (N_17933,N_16637,N_16154);
or U17934 (N_17934,N_16549,N_16921);
nand U17935 (N_17935,N_16184,N_16312);
xnor U17936 (N_17936,N_16951,N_16322);
and U17937 (N_17937,N_16341,N_16741);
xor U17938 (N_17938,N_16641,N_16389);
xor U17939 (N_17939,N_16291,N_16041);
xnor U17940 (N_17940,N_16278,N_16327);
nand U17941 (N_17941,N_16422,N_16867);
nand U17942 (N_17942,N_16271,N_16071);
or U17943 (N_17943,N_16797,N_16489);
nor U17944 (N_17944,N_16054,N_16306);
and U17945 (N_17945,N_16698,N_16315);
and U17946 (N_17946,N_16302,N_16128);
nand U17947 (N_17947,N_16029,N_16622);
or U17948 (N_17948,N_16130,N_16091);
and U17949 (N_17949,N_16223,N_16756);
nand U17950 (N_17950,N_16337,N_16454);
xnor U17951 (N_17951,N_16267,N_16843);
and U17952 (N_17952,N_16472,N_16503);
or U17953 (N_17953,N_16900,N_16555);
nand U17954 (N_17954,N_16502,N_16151);
or U17955 (N_17955,N_16465,N_16743);
and U17956 (N_17956,N_16139,N_16944);
and U17957 (N_17957,N_16159,N_16713);
nand U17958 (N_17958,N_16887,N_16061);
or U17959 (N_17959,N_16145,N_16974);
nor U17960 (N_17960,N_16912,N_16398);
nor U17961 (N_17961,N_16701,N_16871);
or U17962 (N_17962,N_16332,N_16553);
nor U17963 (N_17963,N_16942,N_16234);
and U17964 (N_17964,N_16411,N_16112);
nor U17965 (N_17965,N_16843,N_16528);
and U17966 (N_17966,N_16365,N_16689);
xor U17967 (N_17967,N_16003,N_16174);
xnor U17968 (N_17968,N_16574,N_16991);
nor U17969 (N_17969,N_16697,N_16080);
nor U17970 (N_17970,N_16835,N_16064);
and U17971 (N_17971,N_16784,N_16489);
and U17972 (N_17972,N_16167,N_16309);
and U17973 (N_17973,N_16344,N_16680);
or U17974 (N_17974,N_16994,N_16374);
nand U17975 (N_17975,N_16757,N_16493);
nor U17976 (N_17976,N_16449,N_16072);
nand U17977 (N_17977,N_16660,N_16334);
or U17978 (N_17978,N_16854,N_16597);
and U17979 (N_17979,N_16517,N_16418);
or U17980 (N_17980,N_16521,N_16537);
xnor U17981 (N_17981,N_16172,N_16397);
nor U17982 (N_17982,N_16840,N_16520);
xor U17983 (N_17983,N_16810,N_16610);
nand U17984 (N_17984,N_16780,N_16372);
or U17985 (N_17985,N_16022,N_16064);
or U17986 (N_17986,N_16832,N_16228);
and U17987 (N_17987,N_16032,N_16369);
nor U17988 (N_17988,N_16511,N_16829);
xnor U17989 (N_17989,N_16788,N_16782);
xor U17990 (N_17990,N_16994,N_16314);
nand U17991 (N_17991,N_16190,N_16152);
xnor U17992 (N_17992,N_16504,N_16795);
xnor U17993 (N_17993,N_16713,N_16458);
xnor U17994 (N_17994,N_16574,N_16942);
and U17995 (N_17995,N_16749,N_16548);
nor U17996 (N_17996,N_16031,N_16018);
nand U17997 (N_17997,N_16143,N_16712);
nand U17998 (N_17998,N_16161,N_16031);
nand U17999 (N_17999,N_16071,N_16156);
xor U18000 (N_18000,N_17937,N_17107);
or U18001 (N_18001,N_17499,N_17035);
and U18002 (N_18002,N_17422,N_17776);
nand U18003 (N_18003,N_17565,N_17369);
and U18004 (N_18004,N_17285,N_17350);
nand U18005 (N_18005,N_17971,N_17604);
and U18006 (N_18006,N_17779,N_17335);
and U18007 (N_18007,N_17274,N_17302);
and U18008 (N_18008,N_17169,N_17060);
nor U18009 (N_18009,N_17818,N_17367);
nor U18010 (N_18010,N_17943,N_17773);
xnor U18011 (N_18011,N_17252,N_17662);
nand U18012 (N_18012,N_17742,N_17944);
nand U18013 (N_18013,N_17714,N_17244);
nor U18014 (N_18014,N_17621,N_17466);
xor U18015 (N_18015,N_17082,N_17317);
xor U18016 (N_18016,N_17054,N_17484);
nand U18017 (N_18017,N_17343,N_17151);
or U18018 (N_18018,N_17724,N_17786);
nand U18019 (N_18019,N_17845,N_17235);
nand U18020 (N_18020,N_17100,N_17761);
or U18021 (N_18021,N_17827,N_17096);
nor U18022 (N_18022,N_17223,N_17051);
nor U18023 (N_18023,N_17814,N_17006);
xnor U18024 (N_18024,N_17311,N_17530);
xor U18025 (N_18025,N_17063,N_17140);
or U18026 (N_18026,N_17567,N_17044);
and U18027 (N_18027,N_17670,N_17455);
and U18028 (N_18028,N_17569,N_17372);
or U18029 (N_18029,N_17986,N_17284);
and U18030 (N_18030,N_17463,N_17009);
nand U18031 (N_18031,N_17889,N_17234);
or U18032 (N_18032,N_17848,N_17595);
nor U18033 (N_18033,N_17609,N_17646);
nand U18034 (N_18034,N_17475,N_17780);
nor U18035 (N_18035,N_17069,N_17798);
nor U18036 (N_18036,N_17440,N_17480);
or U18037 (N_18037,N_17053,N_17358);
nand U18038 (N_18038,N_17340,N_17197);
xnor U18039 (N_18039,N_17111,N_17913);
nand U18040 (N_18040,N_17675,N_17238);
xor U18041 (N_18041,N_17411,N_17696);
nor U18042 (N_18042,N_17478,N_17878);
nor U18043 (N_18043,N_17504,N_17263);
xor U18044 (N_18044,N_17697,N_17259);
or U18045 (N_18045,N_17799,N_17071);
xor U18046 (N_18046,N_17574,N_17453);
and U18047 (N_18047,N_17771,N_17007);
and U18048 (N_18048,N_17092,N_17099);
and U18049 (N_18049,N_17619,N_17547);
or U18050 (N_18050,N_17982,N_17147);
nand U18051 (N_18051,N_17948,N_17170);
nor U18052 (N_18052,N_17141,N_17860);
or U18053 (N_18053,N_17510,N_17528);
nand U18054 (N_18054,N_17325,N_17098);
xnor U18055 (N_18055,N_17308,N_17388);
xnor U18056 (N_18056,N_17294,N_17907);
nand U18057 (N_18057,N_17433,N_17571);
or U18058 (N_18058,N_17136,N_17130);
or U18059 (N_18059,N_17674,N_17166);
or U18060 (N_18060,N_17518,N_17239);
and U18061 (N_18061,N_17751,N_17313);
nand U18062 (N_18062,N_17614,N_17014);
nand U18063 (N_18063,N_17795,N_17602);
nor U18064 (N_18064,N_17182,N_17080);
or U18065 (N_18065,N_17836,N_17163);
nor U18066 (N_18066,N_17938,N_17373);
xor U18067 (N_18067,N_17318,N_17032);
nand U18068 (N_18068,N_17105,N_17536);
nor U18069 (N_18069,N_17355,N_17209);
nand U18070 (N_18070,N_17237,N_17002);
nand U18071 (N_18071,N_17632,N_17430);
nand U18072 (N_18072,N_17420,N_17462);
xnor U18073 (N_18073,N_17380,N_17921);
xor U18074 (N_18074,N_17406,N_17570);
or U18075 (N_18075,N_17428,N_17073);
nand U18076 (N_18076,N_17483,N_17923);
or U18077 (N_18077,N_17042,N_17431);
nand U18078 (N_18078,N_17931,N_17143);
or U18079 (N_18079,N_17061,N_17250);
or U18080 (N_18080,N_17660,N_17055);
xor U18081 (N_18081,N_17190,N_17895);
and U18082 (N_18082,N_17142,N_17506);
nand U18083 (N_18083,N_17957,N_17084);
nand U18084 (N_18084,N_17755,N_17286);
xnor U18085 (N_18085,N_17973,N_17908);
nor U18086 (N_18086,N_17535,N_17666);
or U18087 (N_18087,N_17959,N_17371);
and U18088 (N_18088,N_17892,N_17321);
or U18089 (N_18089,N_17902,N_17048);
nand U18090 (N_18090,N_17282,N_17970);
xor U18091 (N_18091,N_17187,N_17467);
and U18092 (N_18092,N_17052,N_17523);
nor U18093 (N_18093,N_17852,N_17503);
nor U18094 (N_18094,N_17337,N_17759);
or U18095 (N_18095,N_17121,N_17767);
or U18096 (N_18096,N_17165,N_17950);
and U18097 (N_18097,N_17947,N_17254);
xor U18098 (N_18098,N_17146,N_17010);
and U18099 (N_18099,N_17634,N_17249);
or U18100 (N_18100,N_17900,N_17904);
nand U18101 (N_18101,N_17323,N_17029);
and U18102 (N_18102,N_17213,N_17086);
nand U18103 (N_18103,N_17362,N_17977);
and U18104 (N_18104,N_17633,N_17550);
xor U18105 (N_18105,N_17514,N_17884);
nand U18106 (N_18106,N_17864,N_17587);
xor U18107 (N_18107,N_17497,N_17865);
and U18108 (N_18108,N_17496,N_17998);
nor U18109 (N_18109,N_17819,N_17677);
and U18110 (N_18110,N_17087,N_17334);
and U18111 (N_18111,N_17625,N_17232);
xor U18112 (N_18112,N_17588,N_17718);
and U18113 (N_18113,N_17058,N_17793);
nor U18114 (N_18114,N_17655,N_17426);
xor U18115 (N_18115,N_17331,N_17410);
nand U18116 (N_18116,N_17920,N_17131);
xnor U18117 (N_18117,N_17457,N_17226);
nor U18118 (N_18118,N_17370,N_17278);
nor U18119 (N_18119,N_17616,N_17749);
or U18120 (N_18120,N_17148,N_17966);
nand U18121 (N_18121,N_17622,N_17615);
or U18122 (N_18122,N_17090,N_17781);
and U18123 (N_18123,N_17137,N_17031);
nor U18124 (N_18124,N_17995,N_17607);
or U18125 (N_18125,N_17653,N_17488);
nand U18126 (N_18126,N_17231,N_17752);
and U18127 (N_18127,N_17418,N_17722);
nand U18128 (N_18128,N_17119,N_17206);
xnor U18129 (N_18129,N_17184,N_17139);
or U18130 (N_18130,N_17630,N_17753);
and U18131 (N_18131,N_17251,N_17482);
or U18132 (N_18132,N_17582,N_17954);
nor U18133 (N_18133,N_17933,N_17915);
xnor U18134 (N_18134,N_17705,N_17981);
or U18135 (N_18135,N_17850,N_17290);
and U18136 (N_18136,N_17415,N_17731);
and U18137 (N_18137,N_17785,N_17620);
xor U18138 (N_18138,N_17561,N_17867);
and U18139 (N_18139,N_17432,N_17922);
nor U18140 (N_18140,N_17091,N_17050);
or U18141 (N_18141,N_17702,N_17545);
nand U18142 (N_18142,N_17534,N_17078);
nand U18143 (N_18143,N_17603,N_17026);
xnor U18144 (N_18144,N_17955,N_17548);
nand U18145 (N_18145,N_17424,N_17964);
xnor U18146 (N_18146,N_17095,N_17610);
and U18147 (N_18147,N_17085,N_17553);
nor U18148 (N_18148,N_17345,N_17794);
or U18149 (N_18149,N_17840,N_17292);
or U18150 (N_18150,N_17332,N_17508);
nor U18151 (N_18151,N_17210,N_17917);
nand U18152 (N_18152,N_17382,N_17783);
nand U18153 (N_18153,N_17381,N_17038);
and U18154 (N_18154,N_17152,N_17713);
nand U18155 (N_18155,N_17024,N_17450);
xor U18156 (N_18156,N_17366,N_17576);
nand U18157 (N_18157,N_17558,N_17606);
nand U18158 (N_18158,N_17277,N_17460);
nor U18159 (N_18159,N_17300,N_17994);
and U18160 (N_18160,N_17649,N_17976);
xnor U18161 (N_18161,N_17474,N_17454);
and U18162 (N_18162,N_17017,N_17260);
or U18163 (N_18163,N_17062,N_17979);
nor U18164 (N_18164,N_17796,N_17368);
and U18165 (N_18165,N_17663,N_17189);
nand U18166 (N_18166,N_17229,N_17887);
and U18167 (N_18167,N_17305,N_17672);
or U18168 (N_18168,N_17703,N_17778);
or U18169 (N_18169,N_17314,N_17680);
or U18170 (N_18170,N_17270,N_17477);
nor U18171 (N_18171,N_17802,N_17888);
nor U18172 (N_18172,N_17132,N_17436);
and U18173 (N_18173,N_17160,N_17495);
and U18174 (N_18174,N_17935,N_17600);
nand U18175 (N_18175,N_17127,N_17122);
xor U18176 (N_18176,N_17135,N_17578);
xnor U18177 (N_18177,N_17806,N_17097);
or U18178 (N_18178,N_17880,N_17013);
nor U18179 (N_18179,N_17591,N_17765);
and U18180 (N_18180,N_17447,N_17364);
or U18181 (N_18181,N_17877,N_17809);
and U18182 (N_18182,N_17441,N_17461);
or U18183 (N_18183,N_17968,N_17790);
nor U18184 (N_18184,N_17732,N_17312);
xnor U18185 (N_18185,N_17280,N_17684);
nand U18186 (N_18186,N_17766,N_17719);
nor U18187 (N_18187,N_17064,N_17172);
xnor U18188 (N_18188,N_17081,N_17720);
nand U18189 (N_18189,N_17654,N_17631);
or U18190 (N_18190,N_17365,N_17228);
xnor U18191 (N_18191,N_17328,N_17936);
or U18192 (N_18192,N_17804,N_17517);
or U18193 (N_18193,N_17434,N_17458);
nor U18194 (N_18194,N_17640,N_17853);
or U18195 (N_18195,N_17671,N_17989);
and U18196 (N_18196,N_17425,N_17939);
or U18197 (N_18197,N_17109,N_17896);
nor U18198 (N_18198,N_17925,N_17188);
nand U18199 (N_18199,N_17124,N_17158);
nand U18200 (N_18200,N_17645,N_17327);
and U18201 (N_18201,N_17106,N_17808);
nand U18202 (N_18202,N_17018,N_17863);
nand U18203 (N_18203,N_17826,N_17505);
and U18204 (N_18204,N_17159,N_17849);
xor U18205 (N_18205,N_17324,N_17690);
xor U18206 (N_18206,N_17816,N_17033);
nor U18207 (N_18207,N_17427,N_17171);
xor U18208 (N_18208,N_17316,N_17906);
xnor U18209 (N_18209,N_17067,N_17423);
nand U18210 (N_18210,N_17201,N_17828);
xnor U18211 (N_18211,N_17643,N_17245);
nand U18212 (N_18212,N_17205,N_17928);
nor U18213 (N_18213,N_17813,N_17554);
and U18214 (N_18214,N_17162,N_17811);
nand U18215 (N_18215,N_17004,N_17685);
nand U18216 (N_18216,N_17624,N_17635);
nand U18217 (N_18217,N_17469,N_17834);
or U18218 (N_18218,N_17012,N_17176);
and U18219 (N_18219,N_17777,N_17575);
xor U18220 (N_18220,N_17193,N_17704);
xnor U18221 (N_18221,N_17695,N_17472);
and U18222 (N_18222,N_17586,N_17056);
nand U18223 (N_18223,N_17740,N_17339);
nand U18224 (N_18224,N_17583,N_17074);
and U18225 (N_18225,N_17637,N_17155);
nand U18226 (N_18226,N_17792,N_17304);
and U18227 (N_18227,N_17676,N_17596);
xnor U18228 (N_18228,N_17198,N_17295);
and U18229 (N_18229,N_17605,N_17248);
or U18230 (N_18230,N_17835,N_17760);
nor U18231 (N_18231,N_17651,N_17279);
or U18232 (N_18232,N_17089,N_17531);
or U18233 (N_18233,N_17627,N_17661);
nand U18234 (N_18234,N_17710,N_17479);
nand U18235 (N_18235,N_17844,N_17173);
xor U18236 (N_18236,N_17126,N_17299);
or U18237 (N_18237,N_17247,N_17094);
nor U18238 (N_18238,N_17273,N_17956);
or U18239 (N_18239,N_17526,N_17572);
and U18240 (N_18240,N_17218,N_17648);
nor U18241 (N_18241,N_17047,N_17214);
xor U18242 (N_18242,N_17784,N_17529);
or U18243 (N_18243,N_17893,N_17445);
and U18244 (N_18244,N_17599,N_17594);
nor U18245 (N_18245,N_17791,N_17065);
or U18246 (N_18246,N_17664,N_17725);
or U18247 (N_18247,N_17608,N_17439);
xnor U18248 (N_18248,N_17805,N_17133);
and U18249 (N_18249,N_17876,N_17629);
or U18250 (N_18250,N_17841,N_17379);
nand U18251 (N_18251,N_17230,N_17585);
and U18252 (N_18252,N_17150,N_17041);
and U18253 (N_18253,N_17438,N_17909);
xor U18254 (N_18254,N_17543,N_17110);
xor U18255 (N_18255,N_17405,N_17824);
or U18256 (N_18256,N_17952,N_17967);
nor U18257 (N_18257,N_17568,N_17872);
nand U18258 (N_18258,N_17102,N_17521);
nor U18259 (N_18259,N_17498,N_17224);
and U18260 (N_18260,N_17665,N_17177);
or U18261 (N_18261,N_17866,N_17289);
nand U18262 (N_18262,N_17402,N_17397);
xnor U18263 (N_18263,N_17984,N_17222);
and U18264 (N_18264,N_17003,N_17540);
and U18265 (N_18265,N_17386,N_17942);
and U18266 (N_18266,N_17961,N_17387);
nand U18267 (N_18267,N_17855,N_17233);
or U18268 (N_18268,N_17359,N_17659);
xor U18269 (N_18269,N_17638,N_17739);
or U18270 (N_18270,N_17825,N_17515);
nand U18271 (N_18271,N_17398,N_17999);
nand U18272 (N_18272,N_17590,N_17837);
nand U18273 (N_18273,N_17036,N_17885);
or U18274 (N_18274,N_17958,N_17291);
nand U18275 (N_18275,N_17138,N_17823);
or U18276 (N_18276,N_17847,N_17862);
or U18277 (N_18277,N_17527,N_17442);
xor U18278 (N_18278,N_17821,N_17829);
xor U18279 (N_18279,N_17396,N_17429);
nand U18280 (N_18280,N_17112,N_17326);
and U18281 (N_18281,N_17916,N_17212);
nor U18282 (N_18282,N_17987,N_17195);
xnor U18283 (N_18283,N_17501,N_17219);
or U18284 (N_18284,N_17113,N_17057);
nor U18285 (N_18285,N_17762,N_17348);
or U18286 (N_18286,N_17117,N_17891);
nor U18287 (N_18287,N_17644,N_17181);
xnor U18288 (N_18288,N_17681,N_17361);
xnor U18289 (N_18289,N_17417,N_17833);
nand U18290 (N_18290,N_17682,N_17227);
nand U18291 (N_18291,N_17859,N_17949);
or U18292 (N_18292,N_17800,N_17716);
nor U18293 (N_18293,N_17025,N_17019);
and U18294 (N_18294,N_17511,N_17465);
and U18295 (N_18295,N_17356,N_17268);
xor U18296 (N_18296,N_17493,N_17559);
and U18297 (N_18297,N_17349,N_17407);
nor U18298 (N_18298,N_17246,N_17544);
xor U18299 (N_18299,N_17838,N_17256);
or U18300 (N_18300,N_17437,N_17642);
xor U18301 (N_18301,N_17408,N_17487);
xnor U18302 (N_18302,N_17075,N_17673);
nor U18303 (N_18303,N_17975,N_17264);
nor U18304 (N_18304,N_17919,N_17581);
nor U18305 (N_18305,N_17211,N_17267);
nand U18306 (N_18306,N_17668,N_17392);
nor U18307 (N_18307,N_17691,N_17522);
and U18308 (N_18308,N_17555,N_17191);
nand U18309 (N_18309,N_17120,N_17161);
xor U18310 (N_18310,N_17903,N_17657);
xnor U18311 (N_18311,N_17101,N_17927);
nand U18312 (N_18312,N_17320,N_17403);
or U18313 (N_18313,N_17754,N_17960);
and U18314 (N_18314,N_17843,N_17686);
xor U18315 (N_18315,N_17721,N_17763);
nor U18316 (N_18316,N_17275,N_17192);
nor U18317 (N_18317,N_17129,N_17108);
xnor U18318 (N_18318,N_17932,N_17969);
and U18319 (N_18319,N_17490,N_17338);
or U18320 (N_18320,N_17329,N_17375);
and U18321 (N_18321,N_17728,N_17040);
and U18322 (N_18322,N_17393,N_17934);
or U18323 (N_18323,N_17027,N_17965);
nor U18324 (N_18324,N_17459,N_17687);
nand U18325 (N_18325,N_17116,N_17584);
nand U18326 (N_18326,N_17730,N_17046);
and U18327 (N_18327,N_17525,N_17541);
nor U18328 (N_18328,N_17079,N_17123);
nand U18329 (N_18329,N_17726,N_17283);
nand U18330 (N_18330,N_17412,N_17333);
nand U18331 (N_18331,N_17413,N_17839);
and U18332 (N_18332,N_17911,N_17991);
xnor U18333 (N_18333,N_17817,N_17881);
and U18334 (N_18334,N_17996,N_17168);
xnor U18335 (N_18335,N_17658,N_17030);
xor U18336 (N_18336,N_17118,N_17820);
nand U18337 (N_18337,N_17043,N_17985);
xor U18338 (N_18338,N_17953,N_17419);
xnor U18339 (N_18339,N_17788,N_17346);
or U18340 (N_18340,N_17281,N_17045);
or U18341 (N_18341,N_17993,N_17910);
or U18342 (N_18342,N_17008,N_17183);
and U18343 (N_18343,N_17683,N_17941);
and U18344 (N_18344,N_17551,N_17689);
and U18345 (N_18345,N_17088,N_17861);
nor U18346 (N_18346,N_17489,N_17924);
nand U18347 (N_18347,N_17549,N_17481);
xnor U18348 (N_18348,N_17186,N_17378);
xor U18349 (N_18349,N_17076,N_17879);
or U18350 (N_18350,N_17093,N_17342);
nor U18351 (N_18351,N_17049,N_17562);
nor U18352 (N_18352,N_17692,N_17034);
nand U18353 (N_18353,N_17476,N_17669);
and U18354 (N_18354,N_17978,N_17764);
or U18355 (N_18355,N_17322,N_17699);
nor U18356 (N_18356,N_17748,N_17694);
or U18357 (N_18357,N_17708,N_17072);
xor U18358 (N_18358,N_17733,N_17940);
nand U18359 (N_18359,N_17612,N_17203);
or U18360 (N_18360,N_17717,N_17390);
nor U18361 (N_18361,N_17734,N_17144);
nand U18362 (N_18362,N_17394,N_17180);
nor U18363 (N_18363,N_17507,N_17712);
or U18364 (N_18364,N_17023,N_17451);
nand U18365 (N_18365,N_17443,N_17471);
nand U18366 (N_18366,N_17217,N_17178);
xor U18367 (N_18367,N_17456,N_17898);
nor U18368 (N_18368,N_17240,N_17512);
xnor U18369 (N_18369,N_17128,N_17854);
or U18370 (N_18370,N_17736,N_17846);
or U18371 (N_18371,N_17770,N_17021);
or U18372 (N_18372,N_17974,N_17028);
nor U18373 (N_18373,N_17391,N_17963);
nand U18374 (N_18374,N_17347,N_17901);
nor U18375 (N_18375,N_17039,N_17711);
nor U18376 (N_18376,N_17868,N_17265);
nand U18377 (N_18377,N_17789,N_17988);
or U18378 (N_18378,N_17628,N_17352);
nor U18379 (N_18379,N_17374,N_17464);
xor U18380 (N_18380,N_17194,N_17377);
and U18381 (N_18381,N_17315,N_17639);
or U18382 (N_18382,N_17258,N_17611);
or U18383 (N_18383,N_17276,N_17395);
nand U18384 (N_18384,N_17983,N_17972);
and U18385 (N_18385,N_17491,N_17723);
and U18386 (N_18386,N_17513,N_17566);
nand U18387 (N_18387,N_17115,N_17001);
nor U18388 (N_18388,N_17414,N_17296);
and U18389 (N_18389,N_17797,N_17399);
or U18390 (N_18390,N_17444,N_17700);
nor U18391 (N_18391,N_17874,N_17533);
or U18392 (N_18392,N_17336,N_17351);
or U18393 (N_18393,N_17037,N_17563);
xnor U18394 (N_18394,N_17341,N_17914);
nand U18395 (N_18395,N_17842,N_17494);
nor U18396 (N_18396,N_17579,N_17743);
or U18397 (N_18397,N_17077,N_17747);
and U18398 (N_18398,N_17539,N_17667);
or U18399 (N_18399,N_17500,N_17207);
and U18400 (N_18400,N_17727,N_17946);
or U18401 (N_18401,N_17204,N_17560);
nor U18402 (N_18402,N_17552,N_17875);
nand U18403 (N_18403,N_17509,N_17890);
nand U18404 (N_18404,N_17384,N_17918);
or U18405 (N_18405,N_17871,N_17532);
or U18406 (N_18406,N_17185,N_17452);
xor U18407 (N_18407,N_17992,N_17678);
xnor U18408 (N_18408,N_17376,N_17470);
or U18409 (N_18409,N_17255,N_17011);
or U18410 (N_18410,N_17446,N_17520);
xnor U18411 (N_18411,N_17261,N_17744);
and U18412 (N_18412,N_17242,N_17962);
nand U18413 (N_18413,N_17729,N_17330);
nor U18414 (N_18414,N_17772,N_17899);
nand U18415 (N_18415,N_17400,N_17869);
nand U18416 (N_18416,N_17241,N_17449);
and U18417 (N_18417,N_17641,N_17709);
nor U18418 (N_18418,N_17750,N_17873);
xor U18419 (N_18419,N_17652,N_17134);
nand U18420 (N_18420,N_17179,N_17303);
nand U18421 (N_18421,N_17020,N_17757);
and U18422 (N_18422,N_17894,N_17524);
and U18423 (N_18423,N_17383,N_17758);
or U18424 (N_18424,N_17735,N_17679);
nor U18425 (N_18425,N_17769,N_17016);
and U18426 (N_18426,N_17882,N_17945);
and U18427 (N_18427,N_17309,N_17000);
and U18428 (N_18428,N_17775,N_17262);
nand U18429 (N_18429,N_17537,N_17409);
nor U18430 (N_18430,N_17617,N_17592);
and U18431 (N_18431,N_17266,N_17216);
nand U18432 (N_18432,N_17831,N_17149);
nand U18433 (N_18433,N_17856,N_17636);
and U18434 (N_18434,N_17650,N_17070);
nor U18435 (N_18435,N_17990,N_17492);
xor U18436 (N_18436,N_17404,N_17580);
xor U18437 (N_18437,N_17220,N_17626);
xor U18438 (N_18438,N_17803,N_17221);
xor U18439 (N_18439,N_17801,N_17353);
or U18440 (N_18440,N_17656,N_17215);
nand U18441 (N_18441,N_17756,N_17435);
and U18442 (N_18442,N_17929,N_17741);
or U18443 (N_18443,N_17005,N_17519);
or U18444 (N_18444,N_17167,N_17577);
xor U18445 (N_18445,N_17768,N_17597);
or U18446 (N_18446,N_17589,N_17156);
xnor U18447 (N_18447,N_17059,N_17022);
or U18448 (N_18448,N_17473,N_17287);
xnor U18449 (N_18449,N_17253,N_17306);
nand U18450 (N_18450,N_17068,N_17389);
xnor U18451 (N_18451,N_17557,N_17715);
or U18452 (N_18452,N_17883,N_17707);
xor U18453 (N_18453,N_17357,N_17857);
nand U18454 (N_18454,N_17926,N_17997);
xor U18455 (N_18455,N_17174,N_17502);
xnor U18456 (N_18456,N_17114,N_17243);
nor U18457 (N_18457,N_17870,N_17774);
nor U18458 (N_18458,N_17688,N_17153);
nand U18459 (N_18459,N_17297,N_17421);
and U18460 (N_18460,N_17897,N_17363);
and U18461 (N_18461,N_17613,N_17066);
nor U18462 (N_18462,N_17344,N_17787);
xnor U18463 (N_18463,N_17807,N_17542);
or U18464 (N_18464,N_17546,N_17269);
nand U18465 (N_18465,N_17385,N_17225);
or U18466 (N_18466,N_17701,N_17236);
or U18467 (N_18467,N_17125,N_17486);
or U18468 (N_18468,N_17593,N_17905);
nor U18469 (N_18469,N_17930,N_17401);
nor U18470 (N_18470,N_17737,N_17980);
and U18471 (N_18471,N_17516,N_17145);
nor U18472 (N_18472,N_17175,N_17468);
xor U18473 (N_18473,N_17886,N_17951);
xnor U18474 (N_18474,N_17815,N_17598);
xor U18475 (N_18475,N_17618,N_17782);
xor U18476 (N_18476,N_17199,N_17738);
xor U18477 (N_18477,N_17706,N_17272);
nand U18478 (N_18478,N_17693,N_17154);
nand U18479 (N_18479,N_17822,N_17485);
nand U18480 (N_18480,N_17810,N_17745);
and U18481 (N_18481,N_17912,N_17360);
and U18482 (N_18482,N_17208,N_17298);
and U18483 (N_18483,N_17200,N_17812);
xor U18484 (N_18484,N_17015,N_17698);
and U18485 (N_18485,N_17157,N_17830);
xnor U18486 (N_18486,N_17556,N_17354);
and U18487 (N_18487,N_17448,N_17647);
xnor U18488 (N_18488,N_17307,N_17196);
nor U18489 (N_18489,N_17257,N_17202);
nor U18490 (N_18490,N_17104,N_17746);
nand U18491 (N_18491,N_17573,N_17288);
nand U18492 (N_18492,N_17301,N_17832);
or U18493 (N_18493,N_17164,N_17851);
xor U18494 (N_18494,N_17271,N_17416);
and U18495 (N_18495,N_17319,N_17564);
nor U18496 (N_18496,N_17623,N_17083);
or U18497 (N_18497,N_17103,N_17538);
xor U18498 (N_18498,N_17293,N_17601);
nand U18499 (N_18499,N_17858,N_17310);
nor U18500 (N_18500,N_17473,N_17161);
nand U18501 (N_18501,N_17683,N_17739);
nand U18502 (N_18502,N_17995,N_17696);
nand U18503 (N_18503,N_17273,N_17290);
or U18504 (N_18504,N_17708,N_17214);
xor U18505 (N_18505,N_17312,N_17458);
nand U18506 (N_18506,N_17814,N_17713);
nand U18507 (N_18507,N_17970,N_17846);
and U18508 (N_18508,N_17998,N_17507);
nand U18509 (N_18509,N_17647,N_17653);
and U18510 (N_18510,N_17623,N_17331);
and U18511 (N_18511,N_17396,N_17700);
nand U18512 (N_18512,N_17605,N_17523);
xnor U18513 (N_18513,N_17917,N_17972);
nor U18514 (N_18514,N_17140,N_17573);
nand U18515 (N_18515,N_17440,N_17396);
and U18516 (N_18516,N_17843,N_17372);
and U18517 (N_18517,N_17256,N_17574);
nand U18518 (N_18518,N_17946,N_17438);
or U18519 (N_18519,N_17476,N_17650);
nand U18520 (N_18520,N_17917,N_17832);
nor U18521 (N_18521,N_17768,N_17618);
nand U18522 (N_18522,N_17771,N_17504);
nand U18523 (N_18523,N_17879,N_17436);
xor U18524 (N_18524,N_17885,N_17285);
xor U18525 (N_18525,N_17595,N_17978);
or U18526 (N_18526,N_17300,N_17284);
and U18527 (N_18527,N_17177,N_17583);
nor U18528 (N_18528,N_17145,N_17501);
or U18529 (N_18529,N_17237,N_17614);
xnor U18530 (N_18530,N_17698,N_17467);
xnor U18531 (N_18531,N_17305,N_17443);
xnor U18532 (N_18532,N_17919,N_17798);
or U18533 (N_18533,N_17222,N_17023);
and U18534 (N_18534,N_17746,N_17209);
xnor U18535 (N_18535,N_17903,N_17405);
or U18536 (N_18536,N_17461,N_17628);
nand U18537 (N_18537,N_17457,N_17268);
nor U18538 (N_18538,N_17961,N_17144);
and U18539 (N_18539,N_17897,N_17837);
xnor U18540 (N_18540,N_17301,N_17873);
nor U18541 (N_18541,N_17958,N_17143);
or U18542 (N_18542,N_17410,N_17765);
or U18543 (N_18543,N_17629,N_17660);
nand U18544 (N_18544,N_17205,N_17657);
nor U18545 (N_18545,N_17031,N_17438);
or U18546 (N_18546,N_17105,N_17303);
and U18547 (N_18547,N_17566,N_17756);
nand U18548 (N_18548,N_17161,N_17363);
or U18549 (N_18549,N_17433,N_17396);
or U18550 (N_18550,N_17423,N_17800);
nand U18551 (N_18551,N_17672,N_17678);
and U18552 (N_18552,N_17643,N_17285);
and U18553 (N_18553,N_17273,N_17645);
nand U18554 (N_18554,N_17788,N_17799);
and U18555 (N_18555,N_17211,N_17263);
nor U18556 (N_18556,N_17451,N_17838);
nand U18557 (N_18557,N_17386,N_17334);
or U18558 (N_18558,N_17488,N_17834);
nand U18559 (N_18559,N_17993,N_17120);
and U18560 (N_18560,N_17932,N_17126);
nor U18561 (N_18561,N_17779,N_17498);
nand U18562 (N_18562,N_17367,N_17251);
nor U18563 (N_18563,N_17986,N_17989);
and U18564 (N_18564,N_17234,N_17999);
and U18565 (N_18565,N_17817,N_17823);
nor U18566 (N_18566,N_17548,N_17985);
and U18567 (N_18567,N_17717,N_17152);
nor U18568 (N_18568,N_17705,N_17371);
and U18569 (N_18569,N_17779,N_17696);
nor U18570 (N_18570,N_17031,N_17002);
or U18571 (N_18571,N_17913,N_17570);
xnor U18572 (N_18572,N_17095,N_17496);
nand U18573 (N_18573,N_17602,N_17593);
or U18574 (N_18574,N_17095,N_17709);
nand U18575 (N_18575,N_17974,N_17654);
and U18576 (N_18576,N_17112,N_17627);
nand U18577 (N_18577,N_17328,N_17985);
nand U18578 (N_18578,N_17421,N_17051);
xnor U18579 (N_18579,N_17261,N_17009);
xnor U18580 (N_18580,N_17305,N_17279);
and U18581 (N_18581,N_17342,N_17780);
nand U18582 (N_18582,N_17009,N_17436);
nor U18583 (N_18583,N_17194,N_17668);
and U18584 (N_18584,N_17320,N_17349);
or U18585 (N_18585,N_17529,N_17843);
xnor U18586 (N_18586,N_17818,N_17469);
nand U18587 (N_18587,N_17299,N_17707);
nand U18588 (N_18588,N_17501,N_17766);
and U18589 (N_18589,N_17304,N_17066);
or U18590 (N_18590,N_17866,N_17308);
and U18591 (N_18591,N_17259,N_17199);
nor U18592 (N_18592,N_17390,N_17508);
nor U18593 (N_18593,N_17580,N_17481);
nor U18594 (N_18594,N_17785,N_17782);
or U18595 (N_18595,N_17689,N_17166);
and U18596 (N_18596,N_17924,N_17509);
nor U18597 (N_18597,N_17671,N_17408);
and U18598 (N_18598,N_17653,N_17287);
nor U18599 (N_18599,N_17586,N_17234);
xor U18600 (N_18600,N_17401,N_17165);
or U18601 (N_18601,N_17152,N_17333);
or U18602 (N_18602,N_17240,N_17315);
or U18603 (N_18603,N_17141,N_17036);
or U18604 (N_18604,N_17614,N_17198);
and U18605 (N_18605,N_17604,N_17570);
nor U18606 (N_18606,N_17790,N_17683);
or U18607 (N_18607,N_17147,N_17117);
nand U18608 (N_18608,N_17406,N_17587);
nand U18609 (N_18609,N_17594,N_17428);
and U18610 (N_18610,N_17696,N_17716);
nand U18611 (N_18611,N_17253,N_17456);
xnor U18612 (N_18612,N_17688,N_17083);
nor U18613 (N_18613,N_17867,N_17501);
or U18614 (N_18614,N_17101,N_17091);
nand U18615 (N_18615,N_17879,N_17105);
or U18616 (N_18616,N_17779,N_17939);
and U18617 (N_18617,N_17465,N_17351);
nor U18618 (N_18618,N_17298,N_17853);
nor U18619 (N_18619,N_17926,N_17019);
or U18620 (N_18620,N_17563,N_17968);
and U18621 (N_18621,N_17968,N_17796);
or U18622 (N_18622,N_17805,N_17551);
and U18623 (N_18623,N_17624,N_17373);
nand U18624 (N_18624,N_17073,N_17827);
or U18625 (N_18625,N_17042,N_17169);
or U18626 (N_18626,N_17782,N_17373);
nor U18627 (N_18627,N_17314,N_17151);
and U18628 (N_18628,N_17204,N_17859);
nor U18629 (N_18629,N_17677,N_17527);
nand U18630 (N_18630,N_17174,N_17995);
nand U18631 (N_18631,N_17490,N_17018);
nand U18632 (N_18632,N_17219,N_17662);
nand U18633 (N_18633,N_17854,N_17585);
or U18634 (N_18634,N_17593,N_17552);
nor U18635 (N_18635,N_17966,N_17432);
xnor U18636 (N_18636,N_17223,N_17812);
and U18637 (N_18637,N_17339,N_17550);
xnor U18638 (N_18638,N_17071,N_17361);
nor U18639 (N_18639,N_17534,N_17410);
xnor U18640 (N_18640,N_17387,N_17580);
or U18641 (N_18641,N_17820,N_17991);
xnor U18642 (N_18642,N_17663,N_17216);
nand U18643 (N_18643,N_17666,N_17835);
nor U18644 (N_18644,N_17943,N_17539);
nor U18645 (N_18645,N_17837,N_17137);
nand U18646 (N_18646,N_17127,N_17428);
nor U18647 (N_18647,N_17612,N_17706);
or U18648 (N_18648,N_17477,N_17968);
or U18649 (N_18649,N_17496,N_17945);
xnor U18650 (N_18650,N_17972,N_17605);
xor U18651 (N_18651,N_17298,N_17740);
xnor U18652 (N_18652,N_17627,N_17208);
or U18653 (N_18653,N_17670,N_17443);
nand U18654 (N_18654,N_17925,N_17537);
xnor U18655 (N_18655,N_17986,N_17930);
nand U18656 (N_18656,N_17970,N_17386);
xor U18657 (N_18657,N_17385,N_17812);
xnor U18658 (N_18658,N_17468,N_17008);
nor U18659 (N_18659,N_17153,N_17082);
xor U18660 (N_18660,N_17578,N_17615);
xor U18661 (N_18661,N_17472,N_17088);
nor U18662 (N_18662,N_17217,N_17056);
or U18663 (N_18663,N_17543,N_17596);
and U18664 (N_18664,N_17789,N_17828);
nand U18665 (N_18665,N_17946,N_17100);
xnor U18666 (N_18666,N_17896,N_17781);
nor U18667 (N_18667,N_17473,N_17601);
nor U18668 (N_18668,N_17760,N_17284);
nor U18669 (N_18669,N_17408,N_17810);
xnor U18670 (N_18670,N_17019,N_17432);
xnor U18671 (N_18671,N_17235,N_17874);
or U18672 (N_18672,N_17859,N_17982);
nand U18673 (N_18673,N_17267,N_17370);
or U18674 (N_18674,N_17081,N_17178);
nand U18675 (N_18675,N_17966,N_17265);
nand U18676 (N_18676,N_17564,N_17984);
and U18677 (N_18677,N_17704,N_17699);
xnor U18678 (N_18678,N_17471,N_17727);
nand U18679 (N_18679,N_17241,N_17060);
nand U18680 (N_18680,N_17617,N_17390);
nor U18681 (N_18681,N_17656,N_17384);
nand U18682 (N_18682,N_17099,N_17251);
nand U18683 (N_18683,N_17520,N_17481);
xor U18684 (N_18684,N_17928,N_17906);
xor U18685 (N_18685,N_17634,N_17281);
or U18686 (N_18686,N_17818,N_17211);
nor U18687 (N_18687,N_17878,N_17935);
or U18688 (N_18688,N_17532,N_17307);
and U18689 (N_18689,N_17034,N_17007);
and U18690 (N_18690,N_17573,N_17066);
xnor U18691 (N_18691,N_17550,N_17040);
nand U18692 (N_18692,N_17209,N_17548);
nand U18693 (N_18693,N_17102,N_17704);
or U18694 (N_18694,N_17170,N_17205);
and U18695 (N_18695,N_17919,N_17042);
nor U18696 (N_18696,N_17572,N_17554);
and U18697 (N_18697,N_17615,N_17868);
and U18698 (N_18698,N_17974,N_17945);
nor U18699 (N_18699,N_17972,N_17511);
and U18700 (N_18700,N_17184,N_17293);
or U18701 (N_18701,N_17433,N_17481);
nand U18702 (N_18702,N_17646,N_17846);
and U18703 (N_18703,N_17645,N_17898);
and U18704 (N_18704,N_17356,N_17017);
nor U18705 (N_18705,N_17096,N_17372);
and U18706 (N_18706,N_17624,N_17663);
and U18707 (N_18707,N_17489,N_17482);
xnor U18708 (N_18708,N_17050,N_17714);
xor U18709 (N_18709,N_17904,N_17578);
nor U18710 (N_18710,N_17203,N_17674);
nor U18711 (N_18711,N_17325,N_17478);
nand U18712 (N_18712,N_17241,N_17063);
nand U18713 (N_18713,N_17667,N_17106);
xor U18714 (N_18714,N_17902,N_17533);
nor U18715 (N_18715,N_17340,N_17188);
nand U18716 (N_18716,N_17301,N_17116);
or U18717 (N_18717,N_17026,N_17555);
nand U18718 (N_18718,N_17710,N_17876);
nor U18719 (N_18719,N_17313,N_17726);
nand U18720 (N_18720,N_17243,N_17227);
and U18721 (N_18721,N_17927,N_17870);
and U18722 (N_18722,N_17488,N_17913);
nand U18723 (N_18723,N_17663,N_17567);
xnor U18724 (N_18724,N_17084,N_17843);
and U18725 (N_18725,N_17073,N_17027);
nor U18726 (N_18726,N_17359,N_17499);
and U18727 (N_18727,N_17630,N_17294);
and U18728 (N_18728,N_17874,N_17771);
nand U18729 (N_18729,N_17751,N_17724);
xnor U18730 (N_18730,N_17908,N_17076);
xnor U18731 (N_18731,N_17446,N_17377);
xnor U18732 (N_18732,N_17659,N_17505);
or U18733 (N_18733,N_17917,N_17735);
or U18734 (N_18734,N_17158,N_17620);
nand U18735 (N_18735,N_17486,N_17133);
nor U18736 (N_18736,N_17553,N_17866);
and U18737 (N_18737,N_17237,N_17648);
or U18738 (N_18738,N_17815,N_17547);
nor U18739 (N_18739,N_17506,N_17716);
nand U18740 (N_18740,N_17303,N_17314);
or U18741 (N_18741,N_17510,N_17261);
nor U18742 (N_18742,N_17068,N_17145);
nand U18743 (N_18743,N_17640,N_17268);
nor U18744 (N_18744,N_17614,N_17625);
nor U18745 (N_18745,N_17300,N_17107);
nand U18746 (N_18746,N_17293,N_17759);
nand U18747 (N_18747,N_17544,N_17349);
and U18748 (N_18748,N_17918,N_17400);
xnor U18749 (N_18749,N_17976,N_17027);
nand U18750 (N_18750,N_17992,N_17995);
or U18751 (N_18751,N_17305,N_17102);
nor U18752 (N_18752,N_17970,N_17039);
nand U18753 (N_18753,N_17276,N_17300);
nand U18754 (N_18754,N_17492,N_17416);
nor U18755 (N_18755,N_17439,N_17851);
nand U18756 (N_18756,N_17613,N_17531);
or U18757 (N_18757,N_17082,N_17319);
nor U18758 (N_18758,N_17406,N_17356);
nand U18759 (N_18759,N_17910,N_17283);
or U18760 (N_18760,N_17126,N_17182);
nand U18761 (N_18761,N_17312,N_17547);
nor U18762 (N_18762,N_17140,N_17321);
nand U18763 (N_18763,N_17686,N_17739);
nor U18764 (N_18764,N_17514,N_17999);
and U18765 (N_18765,N_17512,N_17255);
nand U18766 (N_18766,N_17064,N_17711);
nand U18767 (N_18767,N_17580,N_17760);
nand U18768 (N_18768,N_17280,N_17629);
xnor U18769 (N_18769,N_17401,N_17738);
or U18770 (N_18770,N_17697,N_17285);
nand U18771 (N_18771,N_17694,N_17251);
nor U18772 (N_18772,N_17451,N_17605);
nor U18773 (N_18773,N_17602,N_17466);
xnor U18774 (N_18774,N_17021,N_17236);
nor U18775 (N_18775,N_17770,N_17049);
xnor U18776 (N_18776,N_17776,N_17354);
xnor U18777 (N_18777,N_17663,N_17095);
nor U18778 (N_18778,N_17182,N_17597);
or U18779 (N_18779,N_17339,N_17830);
and U18780 (N_18780,N_17405,N_17861);
and U18781 (N_18781,N_17045,N_17799);
xnor U18782 (N_18782,N_17504,N_17078);
xnor U18783 (N_18783,N_17851,N_17700);
xnor U18784 (N_18784,N_17739,N_17046);
or U18785 (N_18785,N_17233,N_17791);
nand U18786 (N_18786,N_17183,N_17748);
xor U18787 (N_18787,N_17222,N_17650);
nand U18788 (N_18788,N_17828,N_17317);
and U18789 (N_18789,N_17319,N_17207);
xnor U18790 (N_18790,N_17259,N_17892);
or U18791 (N_18791,N_17073,N_17683);
and U18792 (N_18792,N_17206,N_17783);
nand U18793 (N_18793,N_17189,N_17187);
nor U18794 (N_18794,N_17598,N_17380);
or U18795 (N_18795,N_17757,N_17089);
nand U18796 (N_18796,N_17132,N_17997);
and U18797 (N_18797,N_17475,N_17147);
nor U18798 (N_18798,N_17936,N_17939);
or U18799 (N_18799,N_17138,N_17535);
xnor U18800 (N_18800,N_17139,N_17804);
nand U18801 (N_18801,N_17352,N_17184);
and U18802 (N_18802,N_17713,N_17026);
nor U18803 (N_18803,N_17989,N_17517);
and U18804 (N_18804,N_17092,N_17714);
or U18805 (N_18805,N_17795,N_17660);
and U18806 (N_18806,N_17204,N_17707);
nor U18807 (N_18807,N_17298,N_17385);
nand U18808 (N_18808,N_17909,N_17204);
xnor U18809 (N_18809,N_17075,N_17608);
or U18810 (N_18810,N_17784,N_17801);
and U18811 (N_18811,N_17124,N_17118);
or U18812 (N_18812,N_17733,N_17708);
nand U18813 (N_18813,N_17200,N_17448);
nor U18814 (N_18814,N_17714,N_17001);
and U18815 (N_18815,N_17976,N_17314);
or U18816 (N_18816,N_17738,N_17809);
or U18817 (N_18817,N_17771,N_17971);
nand U18818 (N_18818,N_17007,N_17265);
nor U18819 (N_18819,N_17413,N_17391);
nor U18820 (N_18820,N_17499,N_17225);
xor U18821 (N_18821,N_17311,N_17365);
nor U18822 (N_18822,N_17812,N_17026);
or U18823 (N_18823,N_17098,N_17838);
and U18824 (N_18824,N_17771,N_17563);
or U18825 (N_18825,N_17936,N_17127);
or U18826 (N_18826,N_17118,N_17119);
nor U18827 (N_18827,N_17833,N_17772);
nand U18828 (N_18828,N_17347,N_17683);
nor U18829 (N_18829,N_17424,N_17331);
nand U18830 (N_18830,N_17754,N_17879);
nand U18831 (N_18831,N_17004,N_17487);
and U18832 (N_18832,N_17839,N_17712);
or U18833 (N_18833,N_17087,N_17562);
nand U18834 (N_18834,N_17754,N_17805);
nand U18835 (N_18835,N_17766,N_17291);
or U18836 (N_18836,N_17784,N_17561);
and U18837 (N_18837,N_17284,N_17878);
or U18838 (N_18838,N_17358,N_17249);
or U18839 (N_18839,N_17618,N_17455);
and U18840 (N_18840,N_17818,N_17264);
xnor U18841 (N_18841,N_17364,N_17365);
or U18842 (N_18842,N_17831,N_17421);
nand U18843 (N_18843,N_17740,N_17963);
xnor U18844 (N_18844,N_17434,N_17920);
nand U18845 (N_18845,N_17949,N_17056);
nand U18846 (N_18846,N_17425,N_17445);
or U18847 (N_18847,N_17194,N_17589);
nor U18848 (N_18848,N_17096,N_17364);
or U18849 (N_18849,N_17474,N_17562);
and U18850 (N_18850,N_17881,N_17073);
or U18851 (N_18851,N_17939,N_17079);
nand U18852 (N_18852,N_17351,N_17600);
nand U18853 (N_18853,N_17877,N_17311);
nor U18854 (N_18854,N_17396,N_17483);
xor U18855 (N_18855,N_17149,N_17855);
xnor U18856 (N_18856,N_17932,N_17206);
nand U18857 (N_18857,N_17936,N_17405);
nand U18858 (N_18858,N_17712,N_17982);
nor U18859 (N_18859,N_17810,N_17531);
nand U18860 (N_18860,N_17855,N_17991);
and U18861 (N_18861,N_17435,N_17789);
nand U18862 (N_18862,N_17325,N_17936);
nand U18863 (N_18863,N_17367,N_17565);
or U18864 (N_18864,N_17467,N_17345);
xnor U18865 (N_18865,N_17493,N_17032);
and U18866 (N_18866,N_17397,N_17820);
nand U18867 (N_18867,N_17601,N_17354);
nand U18868 (N_18868,N_17756,N_17633);
or U18869 (N_18869,N_17910,N_17172);
nand U18870 (N_18870,N_17964,N_17266);
and U18871 (N_18871,N_17212,N_17302);
nor U18872 (N_18872,N_17618,N_17201);
nor U18873 (N_18873,N_17374,N_17801);
nand U18874 (N_18874,N_17698,N_17882);
nor U18875 (N_18875,N_17514,N_17448);
nor U18876 (N_18876,N_17965,N_17057);
and U18877 (N_18877,N_17719,N_17763);
or U18878 (N_18878,N_17890,N_17988);
xnor U18879 (N_18879,N_17468,N_17754);
xnor U18880 (N_18880,N_17640,N_17472);
xnor U18881 (N_18881,N_17307,N_17289);
or U18882 (N_18882,N_17295,N_17945);
nand U18883 (N_18883,N_17217,N_17846);
nand U18884 (N_18884,N_17730,N_17776);
or U18885 (N_18885,N_17313,N_17646);
or U18886 (N_18886,N_17724,N_17970);
nor U18887 (N_18887,N_17681,N_17004);
nand U18888 (N_18888,N_17215,N_17747);
nor U18889 (N_18889,N_17037,N_17437);
and U18890 (N_18890,N_17853,N_17452);
xnor U18891 (N_18891,N_17216,N_17731);
nand U18892 (N_18892,N_17010,N_17375);
nand U18893 (N_18893,N_17626,N_17709);
and U18894 (N_18894,N_17112,N_17880);
xnor U18895 (N_18895,N_17367,N_17444);
nand U18896 (N_18896,N_17858,N_17417);
nand U18897 (N_18897,N_17817,N_17159);
and U18898 (N_18898,N_17008,N_17324);
xnor U18899 (N_18899,N_17903,N_17246);
or U18900 (N_18900,N_17776,N_17291);
nand U18901 (N_18901,N_17101,N_17840);
or U18902 (N_18902,N_17269,N_17843);
and U18903 (N_18903,N_17663,N_17290);
nor U18904 (N_18904,N_17851,N_17841);
xnor U18905 (N_18905,N_17630,N_17830);
or U18906 (N_18906,N_17099,N_17172);
or U18907 (N_18907,N_17029,N_17093);
and U18908 (N_18908,N_17044,N_17369);
nor U18909 (N_18909,N_17250,N_17955);
or U18910 (N_18910,N_17818,N_17234);
and U18911 (N_18911,N_17228,N_17645);
and U18912 (N_18912,N_17099,N_17713);
xnor U18913 (N_18913,N_17769,N_17298);
or U18914 (N_18914,N_17453,N_17658);
or U18915 (N_18915,N_17211,N_17005);
or U18916 (N_18916,N_17685,N_17755);
and U18917 (N_18917,N_17590,N_17028);
xor U18918 (N_18918,N_17428,N_17332);
xor U18919 (N_18919,N_17995,N_17046);
xor U18920 (N_18920,N_17189,N_17885);
nor U18921 (N_18921,N_17649,N_17412);
nor U18922 (N_18922,N_17586,N_17779);
and U18923 (N_18923,N_17836,N_17901);
nor U18924 (N_18924,N_17832,N_17972);
nor U18925 (N_18925,N_17391,N_17517);
and U18926 (N_18926,N_17947,N_17509);
xor U18927 (N_18927,N_17769,N_17624);
nor U18928 (N_18928,N_17243,N_17354);
nor U18929 (N_18929,N_17918,N_17531);
nand U18930 (N_18930,N_17325,N_17304);
nand U18931 (N_18931,N_17052,N_17348);
xor U18932 (N_18932,N_17628,N_17704);
nand U18933 (N_18933,N_17658,N_17873);
or U18934 (N_18934,N_17252,N_17947);
and U18935 (N_18935,N_17921,N_17676);
xor U18936 (N_18936,N_17408,N_17914);
nand U18937 (N_18937,N_17976,N_17999);
xor U18938 (N_18938,N_17171,N_17179);
xnor U18939 (N_18939,N_17327,N_17376);
nand U18940 (N_18940,N_17545,N_17138);
or U18941 (N_18941,N_17225,N_17612);
nor U18942 (N_18942,N_17063,N_17816);
nor U18943 (N_18943,N_17463,N_17810);
nor U18944 (N_18944,N_17958,N_17626);
xor U18945 (N_18945,N_17941,N_17922);
xor U18946 (N_18946,N_17506,N_17787);
nor U18947 (N_18947,N_17094,N_17113);
or U18948 (N_18948,N_17886,N_17182);
and U18949 (N_18949,N_17397,N_17575);
nand U18950 (N_18950,N_17905,N_17480);
nor U18951 (N_18951,N_17561,N_17157);
xor U18952 (N_18952,N_17496,N_17292);
and U18953 (N_18953,N_17090,N_17793);
or U18954 (N_18954,N_17236,N_17845);
nand U18955 (N_18955,N_17044,N_17556);
or U18956 (N_18956,N_17663,N_17150);
nand U18957 (N_18957,N_17522,N_17784);
xnor U18958 (N_18958,N_17543,N_17804);
and U18959 (N_18959,N_17757,N_17684);
nor U18960 (N_18960,N_17596,N_17154);
and U18961 (N_18961,N_17291,N_17070);
nor U18962 (N_18962,N_17642,N_17376);
nor U18963 (N_18963,N_17861,N_17940);
xnor U18964 (N_18964,N_17258,N_17536);
xnor U18965 (N_18965,N_17545,N_17652);
and U18966 (N_18966,N_17538,N_17781);
nand U18967 (N_18967,N_17035,N_17929);
nor U18968 (N_18968,N_17622,N_17203);
nand U18969 (N_18969,N_17789,N_17544);
or U18970 (N_18970,N_17330,N_17341);
nand U18971 (N_18971,N_17316,N_17266);
nand U18972 (N_18972,N_17441,N_17021);
nor U18973 (N_18973,N_17819,N_17330);
nand U18974 (N_18974,N_17739,N_17640);
and U18975 (N_18975,N_17777,N_17591);
xor U18976 (N_18976,N_17918,N_17785);
and U18977 (N_18977,N_17320,N_17091);
and U18978 (N_18978,N_17751,N_17610);
and U18979 (N_18979,N_17651,N_17275);
xor U18980 (N_18980,N_17099,N_17216);
and U18981 (N_18981,N_17256,N_17664);
xor U18982 (N_18982,N_17701,N_17758);
nand U18983 (N_18983,N_17257,N_17831);
and U18984 (N_18984,N_17395,N_17501);
or U18985 (N_18985,N_17024,N_17131);
xnor U18986 (N_18986,N_17629,N_17524);
xor U18987 (N_18987,N_17968,N_17658);
nand U18988 (N_18988,N_17844,N_17750);
xor U18989 (N_18989,N_17656,N_17176);
nor U18990 (N_18990,N_17660,N_17711);
nand U18991 (N_18991,N_17963,N_17299);
nand U18992 (N_18992,N_17370,N_17255);
nand U18993 (N_18993,N_17673,N_17559);
and U18994 (N_18994,N_17775,N_17904);
nand U18995 (N_18995,N_17134,N_17584);
and U18996 (N_18996,N_17709,N_17768);
or U18997 (N_18997,N_17028,N_17129);
or U18998 (N_18998,N_17465,N_17023);
and U18999 (N_18999,N_17188,N_17751);
or U19000 (N_19000,N_18108,N_18688);
and U19001 (N_19001,N_18578,N_18041);
nor U19002 (N_19002,N_18243,N_18565);
or U19003 (N_19003,N_18839,N_18026);
xor U19004 (N_19004,N_18826,N_18723);
xnor U19005 (N_19005,N_18403,N_18802);
or U19006 (N_19006,N_18725,N_18122);
or U19007 (N_19007,N_18359,N_18046);
and U19008 (N_19008,N_18406,N_18677);
xnor U19009 (N_19009,N_18297,N_18394);
and U19010 (N_19010,N_18402,N_18271);
nor U19011 (N_19011,N_18023,N_18196);
nand U19012 (N_19012,N_18367,N_18842);
and U19013 (N_19013,N_18903,N_18880);
and U19014 (N_19014,N_18669,N_18632);
nor U19015 (N_19015,N_18291,N_18020);
and U19016 (N_19016,N_18687,N_18404);
nor U19017 (N_19017,N_18222,N_18541);
and U19018 (N_19018,N_18408,N_18992);
xor U19019 (N_19019,N_18327,N_18328);
nor U19020 (N_19020,N_18888,N_18837);
and U19021 (N_19021,N_18814,N_18320);
and U19022 (N_19022,N_18765,N_18214);
nor U19023 (N_19023,N_18508,N_18847);
and U19024 (N_19024,N_18340,N_18832);
and U19025 (N_19025,N_18848,N_18973);
nand U19026 (N_19026,N_18345,N_18568);
and U19027 (N_19027,N_18716,N_18326);
xnor U19028 (N_19028,N_18812,N_18618);
and U19029 (N_19029,N_18061,N_18639);
or U19030 (N_19030,N_18646,N_18675);
xor U19031 (N_19031,N_18940,N_18948);
nand U19032 (N_19032,N_18799,N_18463);
or U19033 (N_19033,N_18014,N_18794);
or U19034 (N_19034,N_18392,N_18656);
xor U19035 (N_19035,N_18048,N_18130);
nor U19036 (N_19036,N_18754,N_18479);
nor U19037 (N_19037,N_18579,N_18595);
nor U19038 (N_19038,N_18528,N_18845);
and U19039 (N_19039,N_18892,N_18702);
and U19040 (N_19040,N_18501,N_18476);
nor U19041 (N_19041,N_18625,N_18849);
and U19042 (N_19042,N_18171,N_18721);
or U19043 (N_19043,N_18180,N_18818);
and U19044 (N_19044,N_18633,N_18853);
or U19045 (N_19045,N_18575,N_18066);
nand U19046 (N_19046,N_18651,N_18229);
nor U19047 (N_19047,N_18925,N_18142);
or U19048 (N_19048,N_18136,N_18741);
or U19049 (N_19049,N_18365,N_18195);
or U19050 (N_19050,N_18636,N_18768);
nor U19051 (N_19051,N_18265,N_18311);
or U19052 (N_19052,N_18961,N_18844);
nor U19053 (N_19053,N_18609,N_18366);
nor U19054 (N_19054,N_18509,N_18654);
nor U19055 (N_19055,N_18034,N_18589);
nor U19056 (N_19056,N_18024,N_18980);
or U19057 (N_19057,N_18671,N_18640);
or U19058 (N_19058,N_18277,N_18204);
and U19059 (N_19059,N_18088,N_18898);
or U19060 (N_19060,N_18772,N_18036);
nor U19061 (N_19061,N_18005,N_18119);
and U19062 (N_19062,N_18413,N_18986);
nand U19063 (N_19063,N_18432,N_18044);
xnor U19064 (N_19064,N_18778,N_18273);
and U19065 (N_19065,N_18283,N_18092);
or U19066 (N_19066,N_18132,N_18067);
nand U19067 (N_19067,N_18289,N_18648);
and U19068 (N_19068,N_18913,N_18140);
xnor U19069 (N_19069,N_18045,N_18444);
or U19070 (N_19070,N_18596,N_18093);
or U19071 (N_19071,N_18047,N_18909);
nand U19072 (N_19072,N_18105,N_18932);
nand U19073 (N_19073,N_18535,N_18660);
or U19074 (N_19074,N_18001,N_18022);
nand U19075 (N_19075,N_18025,N_18033);
nand U19076 (N_19076,N_18629,N_18858);
nand U19077 (N_19077,N_18550,N_18572);
nand U19078 (N_19078,N_18491,N_18551);
and U19079 (N_19079,N_18164,N_18492);
or U19080 (N_19080,N_18959,N_18415);
or U19081 (N_19081,N_18121,N_18593);
nor U19082 (N_19082,N_18907,N_18447);
and U19083 (N_19083,N_18598,N_18495);
and U19084 (N_19084,N_18835,N_18643);
or U19085 (N_19085,N_18664,N_18101);
or U19086 (N_19086,N_18729,N_18466);
and U19087 (N_19087,N_18743,N_18546);
nor U19088 (N_19088,N_18079,N_18834);
and U19089 (N_19089,N_18621,N_18674);
xor U19090 (N_19090,N_18324,N_18810);
nand U19091 (N_19091,N_18703,N_18599);
nor U19092 (N_19092,N_18971,N_18960);
or U19093 (N_19093,N_18889,N_18638);
xor U19094 (N_19094,N_18526,N_18054);
nor U19095 (N_19095,N_18351,N_18811);
or U19096 (N_19096,N_18538,N_18152);
nand U19097 (N_19097,N_18050,N_18352);
nand U19098 (N_19098,N_18915,N_18659);
or U19099 (N_19099,N_18472,N_18821);
xor U19100 (N_19100,N_18977,N_18698);
nor U19101 (N_19101,N_18544,N_18626);
nor U19102 (N_19102,N_18461,N_18559);
or U19103 (N_19103,N_18037,N_18264);
and U19104 (N_19104,N_18042,N_18715);
xnor U19105 (N_19105,N_18055,N_18653);
xnor U19106 (N_19106,N_18896,N_18694);
xor U19107 (N_19107,N_18013,N_18678);
and U19108 (N_19108,N_18594,N_18474);
nand U19109 (N_19109,N_18440,N_18699);
nand U19110 (N_19110,N_18086,N_18455);
xnor U19111 (N_19111,N_18877,N_18731);
and U19112 (N_19112,N_18337,N_18689);
nand U19113 (N_19113,N_18419,N_18829);
or U19114 (N_19114,N_18049,N_18943);
xnor U19115 (N_19115,N_18906,N_18155);
and U19116 (N_19116,N_18582,N_18970);
nand U19117 (N_19117,N_18983,N_18567);
nand U19118 (N_19118,N_18697,N_18790);
xnor U19119 (N_19119,N_18177,N_18543);
xnor U19120 (N_19120,N_18780,N_18900);
nor U19121 (N_19121,N_18241,N_18695);
nor U19122 (N_19122,N_18756,N_18602);
nor U19123 (N_19123,N_18512,N_18299);
and U19124 (N_19124,N_18872,N_18244);
or U19125 (N_19125,N_18564,N_18963);
nand U19126 (N_19126,N_18902,N_18300);
nand U19127 (N_19127,N_18205,N_18797);
or U19128 (N_19128,N_18255,N_18555);
nand U19129 (N_19129,N_18379,N_18708);
xnor U19130 (N_19130,N_18770,N_18720);
xor U19131 (N_19131,N_18315,N_18262);
nor U19132 (N_19132,N_18422,N_18998);
or U19133 (N_19133,N_18477,N_18323);
or U19134 (N_19134,N_18808,N_18257);
or U19135 (N_19135,N_18249,N_18782);
nand U19136 (N_19136,N_18165,N_18377);
and U19137 (N_19137,N_18893,N_18679);
nand U19138 (N_19138,N_18038,N_18803);
or U19139 (N_19139,N_18336,N_18967);
nand U19140 (N_19140,N_18159,N_18384);
nand U19141 (N_19141,N_18733,N_18712);
and U19142 (N_19142,N_18901,N_18557);
or U19143 (N_19143,N_18601,N_18994);
nor U19144 (N_19144,N_18278,N_18426);
and U19145 (N_19145,N_18836,N_18469);
and U19146 (N_19146,N_18717,N_18975);
xnor U19147 (N_19147,N_18414,N_18775);
nand U19148 (N_19148,N_18822,N_18104);
xnor U19149 (N_19149,N_18891,N_18087);
and U19150 (N_19150,N_18997,N_18350);
nand U19151 (N_19151,N_18928,N_18833);
or U19152 (N_19152,N_18870,N_18873);
or U19153 (N_19153,N_18287,N_18007);
nand U19154 (N_19154,N_18757,N_18825);
xor U19155 (N_19155,N_18939,N_18094);
and U19156 (N_19156,N_18245,N_18224);
nand U19157 (N_19157,N_18059,N_18655);
or U19158 (N_19158,N_18927,N_18886);
xor U19159 (N_19159,N_18129,N_18161);
nand U19160 (N_19160,N_18935,N_18857);
and U19161 (N_19161,N_18711,N_18773);
and U19162 (N_19162,N_18968,N_18192);
xor U19163 (N_19163,N_18138,N_18313);
or U19164 (N_19164,N_18309,N_18506);
and U19165 (N_19165,N_18281,N_18606);
xnor U19166 (N_19166,N_18577,N_18433);
nand U19167 (N_19167,N_18991,N_18393);
nand U19168 (N_19168,N_18126,N_18747);
or U19169 (N_19169,N_18391,N_18923);
and U19170 (N_19170,N_18964,N_18786);
or U19171 (N_19171,N_18396,N_18914);
nor U19172 (N_19172,N_18670,N_18332);
nor U19173 (N_19173,N_18256,N_18389);
or U19174 (N_19174,N_18360,N_18722);
or U19175 (N_19175,N_18742,N_18381);
or U19176 (N_19176,N_18623,N_18533);
or U19177 (N_19177,N_18681,N_18475);
nand U19178 (N_19178,N_18987,N_18356);
xor U19179 (N_19179,N_18074,N_18363);
nor U19180 (N_19180,N_18075,N_18260);
or U19181 (N_19181,N_18172,N_18482);
and U19182 (N_19182,N_18343,N_18372);
and U19183 (N_19183,N_18869,N_18330);
nand U19184 (N_19184,N_18062,N_18227);
xor U19185 (N_19185,N_18931,N_18739);
and U19186 (N_19186,N_18458,N_18247);
nor U19187 (N_19187,N_18220,N_18098);
or U19188 (N_19188,N_18591,N_18894);
xnor U19189 (N_19189,N_18107,N_18792);
nor U19190 (N_19190,N_18603,N_18258);
or U19191 (N_19191,N_18370,N_18411);
xor U19192 (N_19192,N_18056,N_18057);
and U19193 (N_19193,N_18573,N_18950);
nor U19194 (N_19194,N_18724,N_18652);
xnor U19195 (N_19195,N_18106,N_18198);
nor U19196 (N_19196,N_18123,N_18993);
or U19197 (N_19197,N_18542,N_18103);
and U19198 (N_19198,N_18769,N_18282);
xnor U19199 (N_19199,N_18497,N_18462);
or U19200 (N_19200,N_18125,N_18409);
nand U19201 (N_19201,N_18147,N_18860);
xor U19202 (N_19202,N_18060,N_18371);
nor U19203 (N_19203,N_18868,N_18956);
xor U19204 (N_19204,N_18700,N_18916);
nand U19205 (N_19205,N_18583,N_18390);
and U19206 (N_19206,N_18451,N_18270);
and U19207 (N_19207,N_18436,N_18460);
nor U19208 (N_19208,N_18331,N_18232);
nand U19209 (N_19209,N_18976,N_18128);
and U19210 (N_19210,N_18637,N_18912);
or U19211 (N_19211,N_18316,N_18069);
xor U19212 (N_19212,N_18070,N_18718);
nand U19213 (N_19213,N_18563,N_18684);
and U19214 (N_19214,N_18358,N_18425);
or U19215 (N_19215,N_18017,N_18251);
nand U19216 (N_19216,N_18111,N_18134);
or U19217 (N_19217,N_18325,N_18665);
xnor U19218 (N_19218,N_18569,N_18515);
and U19219 (N_19219,N_18974,N_18112);
or U19220 (N_19220,N_18073,N_18303);
and U19221 (N_19221,N_18401,N_18011);
xnor U19222 (N_19222,N_18503,N_18319);
nor U19223 (N_19223,N_18958,N_18614);
nand U19224 (N_19224,N_18824,N_18179);
nand U19225 (N_19225,N_18597,N_18223);
and U19226 (N_19226,N_18984,N_18003);
and U19227 (N_19227,N_18480,N_18875);
xor U19228 (N_19228,N_18449,N_18453);
xnor U19229 (N_19229,N_18235,N_18558);
nor U19230 (N_19230,N_18936,N_18882);
nand U19231 (N_19231,N_18275,N_18354);
or U19232 (N_19232,N_18279,N_18485);
xor U19233 (N_19233,N_18562,N_18375);
nand U19234 (N_19234,N_18946,N_18787);
nor U19235 (N_19235,N_18053,N_18237);
nor U19236 (N_19236,N_18793,N_18815);
nor U19237 (N_19237,N_18254,N_18890);
or U19238 (N_19238,N_18704,N_18955);
nor U19239 (N_19239,N_18314,N_18604);
nor U19240 (N_19240,N_18019,N_18441);
xnor U19241 (N_19241,N_18552,N_18090);
or U19242 (N_19242,N_18211,N_18201);
xnor U19243 (N_19243,N_18318,N_18800);
nand U19244 (N_19244,N_18376,N_18173);
and U19245 (N_19245,N_18981,N_18002);
xor U19246 (N_19246,N_18897,N_18216);
nor U19247 (N_19247,N_18008,N_18420);
nand U19248 (N_19248,N_18952,N_18197);
and U19249 (N_19249,N_18846,N_18428);
or U19250 (N_19250,N_18758,N_18862);
nor U19251 (N_19251,N_18553,N_18921);
xor U19252 (N_19252,N_18911,N_18728);
or U19253 (N_19253,N_18310,N_18286);
or U19254 (N_19254,N_18761,N_18215);
xnor U19255 (N_19255,N_18346,N_18517);
or U19256 (N_19256,N_18631,N_18202);
nand U19257 (N_19257,N_18368,N_18124);
nor U19258 (N_19258,N_18749,N_18693);
nor U19259 (N_19259,N_18524,N_18369);
and U19260 (N_19260,N_18184,N_18183);
nor U19261 (N_19261,N_18727,N_18021);
or U19262 (N_19262,N_18774,N_18305);
nand U19263 (N_19263,N_18341,N_18231);
or U19264 (N_19264,N_18942,N_18879);
nand U19265 (N_19265,N_18511,N_18957);
or U19266 (N_19266,N_18039,N_18321);
and U19267 (N_19267,N_18110,N_18004);
and U19268 (N_19268,N_18269,N_18416);
nor U19269 (N_19269,N_18851,N_18922);
nor U19270 (N_19270,N_18006,N_18854);
xnor U19271 (N_19271,N_18141,N_18445);
or U19272 (N_19272,N_18692,N_18487);
nand U19273 (N_19273,N_18096,N_18924);
xnor U19274 (N_19274,N_18624,N_18236);
or U19275 (N_19275,N_18176,N_18493);
or U19276 (N_19276,N_18185,N_18820);
xor U19277 (N_19277,N_18146,N_18581);
nor U19278 (N_19278,N_18755,N_18471);
nor U19279 (N_19279,N_18212,N_18418);
and U19280 (N_19280,N_18200,N_18884);
nand U19281 (N_19281,N_18540,N_18031);
or U19282 (N_19282,N_18355,N_18856);
nor U19283 (N_19283,N_18263,N_18947);
xnor U19284 (N_19284,N_18502,N_18828);
and U19285 (N_19285,N_18691,N_18522);
or U19286 (N_19286,N_18429,N_18488);
or U19287 (N_19287,N_18899,N_18657);
and U19288 (N_19288,N_18261,N_18918);
xnor U19289 (N_19289,N_18242,N_18949);
or U19290 (N_19290,N_18478,N_18250);
or U19291 (N_19291,N_18139,N_18430);
xor U19292 (N_19292,N_18089,N_18634);
and U19293 (N_19293,N_18586,N_18170);
and U19294 (N_19294,N_18798,N_18437);
or U19295 (N_19295,N_18989,N_18527);
xnor U19296 (N_19296,N_18954,N_18380);
or U19297 (N_19297,N_18118,N_18353);
nor U19298 (N_19298,N_18666,N_18292);
xor U19299 (N_19299,N_18945,N_18904);
nand U19300 (N_19300,N_18951,N_18154);
or U19301 (N_19301,N_18855,N_18068);
and U19302 (N_19302,N_18334,N_18871);
nand U19303 (N_19303,N_18199,N_18560);
xor U19304 (N_19304,N_18435,N_18645);
or U19305 (N_19305,N_18628,N_18113);
xor U19306 (N_19306,N_18117,N_18168);
nand U19307 (N_19307,N_18308,N_18417);
and U19308 (N_19308,N_18431,N_18744);
nor U19309 (N_19309,N_18745,N_18407);
xnor U19310 (N_19310,N_18162,N_18673);
xnor U19311 (N_19311,N_18468,N_18887);
nand U19312 (N_19312,N_18153,N_18737);
and U19313 (N_19313,N_18878,N_18317);
nor U19314 (N_19314,N_18467,N_18298);
or U19315 (N_19315,N_18966,N_18496);
and U19316 (N_19316,N_18133,N_18819);
nand U19317 (N_19317,N_18547,N_18807);
and U19318 (N_19318,N_18539,N_18293);
nor U19319 (N_19319,N_18446,N_18937);
nor U19320 (N_19320,N_18686,N_18169);
nand U19321 (N_19321,N_18226,N_18217);
xor U19322 (N_19322,N_18203,N_18521);
or U19323 (N_19323,N_18210,N_18908);
or U19324 (N_19324,N_18166,N_18080);
nand U19325 (N_19325,N_18919,N_18206);
nand U19326 (N_19326,N_18213,N_18456);
nor U19327 (N_19327,N_18574,N_18443);
nor U19328 (N_19328,N_18099,N_18160);
xnor U19329 (N_19329,N_18347,N_18690);
and U19330 (N_19330,N_18783,N_18619);
or U19331 (N_19331,N_18424,N_18018);
nand U19332 (N_19332,N_18612,N_18649);
nand U19333 (N_19333,N_18709,N_18710);
xor U19334 (N_19334,N_18804,N_18063);
xor U19335 (N_19335,N_18100,N_18536);
nand U19336 (N_19336,N_18627,N_18953);
xnor U19337 (N_19337,N_18191,N_18838);
xnor U19338 (N_19338,N_18187,N_18076);
nor U19339 (N_19339,N_18504,N_18373);
xor U19340 (N_19340,N_18454,N_18450);
nand U19341 (N_19341,N_18611,N_18398);
nand U19342 (N_19342,N_18995,N_18499);
and U19343 (N_19343,N_18081,N_18841);
nor U19344 (N_19344,N_18374,N_18442);
and U19345 (N_19345,N_18246,N_18072);
nor U19346 (N_19346,N_18507,N_18427);
and U19347 (N_19347,N_18040,N_18516);
nand U19348 (N_19348,N_18605,N_18127);
xor U19349 (N_19349,N_18190,N_18642);
nand U19350 (N_19350,N_18933,N_18620);
xnor U19351 (N_19351,N_18012,N_18534);
nand U19352 (N_19352,N_18616,N_18266);
xnor U19353 (N_19353,N_18484,N_18990);
and U19354 (N_19354,N_18344,N_18867);
nor U19355 (N_19355,N_18043,N_18883);
xnor U19356 (N_19356,N_18158,N_18561);
nand U19357 (N_19357,N_18505,N_18486);
xor U19358 (N_19358,N_18145,N_18570);
nand U19359 (N_19359,N_18208,N_18766);
nand U19360 (N_19360,N_18713,N_18143);
and U19361 (N_19361,N_18771,N_18464);
nand U19362 (N_19362,N_18051,N_18630);
or U19363 (N_19363,N_18186,N_18682);
nand U19364 (N_19364,N_18077,N_18816);
or U19365 (N_19365,N_18549,N_18592);
and U19366 (N_19366,N_18233,N_18500);
and U19367 (N_19367,N_18452,N_18996);
nand U19368 (N_19368,N_18661,N_18796);
nor U19369 (N_19369,N_18301,N_18296);
or U19370 (N_19370,N_18091,N_18514);
and U19371 (N_19371,N_18658,N_18362);
nand U19372 (N_19372,N_18157,N_18181);
nor U19373 (N_19373,N_18760,N_18707);
nor U19374 (N_19374,N_18714,N_18972);
xnor U19375 (N_19375,N_18483,N_18131);
nor U19376 (N_19376,N_18830,N_18342);
or U19377 (N_19377,N_18175,N_18732);
or U19378 (N_19378,N_18676,N_18459);
and U19379 (N_19379,N_18580,N_18763);
xor U19380 (N_19380,N_18641,N_18525);
xnor U19381 (N_19381,N_18530,N_18357);
nand U19382 (N_19382,N_18817,N_18163);
and U19383 (N_19383,N_18701,N_18751);
or U19384 (N_19384,N_18189,N_18777);
nand U19385 (N_19385,N_18934,N_18082);
nand U19386 (N_19386,N_18193,N_18000);
nor U19387 (N_19387,N_18498,N_18364);
and U19388 (N_19388,N_18400,N_18225);
nor U19389 (N_19389,N_18985,N_18663);
or U19390 (N_19390,N_18071,N_18457);
xnor U19391 (N_19391,N_18284,N_18329);
nand U19392 (N_19392,N_18135,N_18622);
and U19393 (N_19393,N_18150,N_18102);
and U19394 (N_19394,N_18779,N_18672);
xnor U19395 (N_19395,N_18294,N_18388);
or U19396 (N_19396,N_18613,N_18188);
nand U19397 (N_19397,N_18410,N_18979);
and U19398 (N_19398,N_18259,N_18009);
or U19399 (N_19399,N_18905,N_18685);
nor U19400 (N_19400,N_18537,N_18750);
and U19401 (N_19401,N_18863,N_18065);
nand U19402 (N_19402,N_18748,N_18576);
xnor U19403 (N_19403,N_18831,N_18209);
nand U19404 (N_19404,N_18349,N_18806);
and U19405 (N_19405,N_18240,N_18338);
or U19406 (N_19406,N_18412,N_18030);
and U19407 (N_19407,N_18885,N_18207);
nand U19408 (N_19408,N_18929,N_18584);
nand U19409 (N_19409,N_18650,N_18285);
nand U19410 (N_19410,N_18267,N_18590);
and U19411 (N_19411,N_18052,N_18753);
nor U19412 (N_19412,N_18941,N_18386);
nor U19413 (N_19413,N_18084,N_18156);
or U19414 (N_19414,N_18383,N_18813);
xor U19415 (N_19415,N_18668,N_18827);
nand U19416 (N_19416,N_18764,N_18439);
nand U19417 (N_19417,N_18859,N_18115);
nor U19418 (N_19418,N_18809,N_18607);
nor U19419 (N_19419,N_18805,N_18520);
nand U19420 (N_19420,N_18519,N_18734);
nand U19421 (N_19421,N_18571,N_18738);
xor U19422 (N_19422,N_18978,N_18144);
xnor U19423 (N_19423,N_18312,N_18322);
nand U19424 (N_19424,N_18554,N_18015);
nor U19425 (N_19425,N_18999,N_18969);
and U19426 (N_19426,N_18035,N_18680);
xnor U19427 (N_19427,N_18843,N_18610);
and U19428 (N_19428,N_18608,N_18348);
nand U19429 (N_19429,N_18290,N_18029);
xnor U19430 (N_19430,N_18776,N_18881);
nor U19431 (N_19431,N_18523,N_18234);
or U19432 (N_19432,N_18531,N_18962);
xnor U19433 (N_19433,N_18280,N_18114);
nor U19434 (N_19434,N_18735,N_18385);
xor U19435 (N_19435,N_18740,N_18274);
and U19436 (N_19436,N_18239,N_18635);
nor U19437 (N_19437,N_18781,N_18295);
nor U19438 (N_19438,N_18789,N_18784);
and U19439 (N_19439,N_18861,N_18615);
or U19440 (N_19440,N_18865,N_18490);
xor U19441 (N_19441,N_18470,N_18926);
or U19442 (N_19442,N_18016,N_18137);
or U19443 (N_19443,N_18438,N_18307);
nand U19444 (N_19444,N_18058,N_18706);
and U19445 (N_19445,N_18288,N_18852);
nor U19446 (N_19446,N_18333,N_18064);
and U19447 (N_19447,N_18248,N_18752);
nor U19448 (N_19448,N_18465,N_18335);
and U19449 (N_19449,N_18788,N_18667);
nor U19450 (N_19450,N_18481,N_18864);
and U19451 (N_19451,N_18545,N_18489);
xor U19452 (N_19452,N_18405,N_18795);
and U19453 (N_19453,N_18518,N_18399);
nor U19454 (N_19454,N_18736,N_18228);
nor U19455 (N_19455,N_18494,N_18548);
nand U19456 (N_19456,N_18920,N_18032);
or U19457 (N_19457,N_18759,N_18588);
nand U19458 (N_19458,N_18010,N_18378);
nor U19459 (N_19459,N_18178,N_18917);
nand U19460 (N_19460,N_18339,N_18302);
nand U19461 (N_19461,N_18696,N_18423);
nor U19462 (N_19462,N_18617,N_18938);
and U19463 (N_19463,N_18397,N_18473);
nand U19464 (N_19464,N_18874,N_18361);
nand U19465 (N_19465,N_18510,N_18532);
xor U19466 (N_19466,N_18421,N_18182);
and U19467 (N_19467,N_18600,N_18448);
nor U19468 (N_19468,N_18767,N_18167);
nor U19469 (N_19469,N_18194,N_18095);
xor U19470 (N_19470,N_18276,N_18116);
nor U19471 (N_19471,N_18585,N_18746);
xor U19472 (N_19472,N_18944,N_18078);
xnor U19473 (N_19473,N_18097,N_18382);
nand U19474 (N_19474,N_18218,N_18823);
nand U19475 (N_19475,N_18272,N_18529);
xnor U19476 (N_19476,N_18566,N_18785);
xor U19477 (N_19477,N_18148,N_18587);
nor U19478 (N_19478,N_18083,N_18230);
or U19479 (N_19479,N_18801,N_18306);
or U19480 (N_19480,N_18726,N_18174);
xor U19481 (N_19481,N_18151,N_18850);
nand U19482 (N_19482,N_18840,N_18219);
and U19483 (N_19483,N_18662,N_18930);
and U19484 (N_19484,N_18268,N_18085);
nand U19485 (N_19485,N_18120,N_18253);
nand U19486 (N_19486,N_18719,N_18149);
or U19487 (N_19487,N_18109,N_18762);
and U19488 (N_19488,N_18434,N_18238);
or U19489 (N_19489,N_18387,N_18683);
nand U19490 (N_19490,N_18395,N_18982);
nor U19491 (N_19491,N_18965,N_18988);
and U19492 (N_19492,N_18513,N_18866);
xnor U19493 (N_19493,N_18304,N_18221);
and U19494 (N_19494,N_18027,N_18791);
xnor U19495 (N_19495,N_18910,N_18705);
and U19496 (N_19496,N_18644,N_18028);
or U19497 (N_19497,N_18730,N_18647);
nand U19498 (N_19498,N_18895,N_18556);
nand U19499 (N_19499,N_18876,N_18252);
nor U19500 (N_19500,N_18446,N_18066);
nor U19501 (N_19501,N_18837,N_18769);
nand U19502 (N_19502,N_18143,N_18103);
xor U19503 (N_19503,N_18607,N_18326);
nand U19504 (N_19504,N_18647,N_18318);
and U19505 (N_19505,N_18914,N_18410);
or U19506 (N_19506,N_18602,N_18585);
and U19507 (N_19507,N_18627,N_18687);
nand U19508 (N_19508,N_18343,N_18819);
xnor U19509 (N_19509,N_18454,N_18106);
or U19510 (N_19510,N_18311,N_18842);
or U19511 (N_19511,N_18069,N_18604);
and U19512 (N_19512,N_18356,N_18795);
nand U19513 (N_19513,N_18637,N_18828);
or U19514 (N_19514,N_18916,N_18925);
xor U19515 (N_19515,N_18562,N_18939);
xnor U19516 (N_19516,N_18848,N_18977);
nand U19517 (N_19517,N_18794,N_18027);
nor U19518 (N_19518,N_18509,N_18900);
nor U19519 (N_19519,N_18386,N_18591);
or U19520 (N_19520,N_18428,N_18912);
nand U19521 (N_19521,N_18346,N_18528);
nand U19522 (N_19522,N_18526,N_18170);
or U19523 (N_19523,N_18642,N_18808);
nand U19524 (N_19524,N_18518,N_18107);
nand U19525 (N_19525,N_18687,N_18243);
nand U19526 (N_19526,N_18998,N_18290);
nand U19527 (N_19527,N_18195,N_18251);
nand U19528 (N_19528,N_18710,N_18744);
nand U19529 (N_19529,N_18814,N_18197);
nor U19530 (N_19530,N_18948,N_18419);
nand U19531 (N_19531,N_18633,N_18983);
or U19532 (N_19532,N_18474,N_18612);
and U19533 (N_19533,N_18168,N_18077);
nand U19534 (N_19534,N_18615,N_18028);
or U19535 (N_19535,N_18809,N_18875);
xnor U19536 (N_19536,N_18225,N_18894);
xnor U19537 (N_19537,N_18099,N_18794);
nand U19538 (N_19538,N_18652,N_18421);
or U19539 (N_19539,N_18812,N_18075);
nor U19540 (N_19540,N_18002,N_18270);
or U19541 (N_19541,N_18099,N_18669);
nor U19542 (N_19542,N_18853,N_18561);
and U19543 (N_19543,N_18176,N_18669);
xnor U19544 (N_19544,N_18989,N_18706);
xnor U19545 (N_19545,N_18598,N_18028);
nor U19546 (N_19546,N_18053,N_18082);
and U19547 (N_19547,N_18426,N_18178);
xnor U19548 (N_19548,N_18547,N_18459);
xor U19549 (N_19549,N_18323,N_18713);
and U19550 (N_19550,N_18258,N_18154);
xor U19551 (N_19551,N_18260,N_18553);
or U19552 (N_19552,N_18682,N_18197);
xor U19553 (N_19553,N_18730,N_18867);
or U19554 (N_19554,N_18198,N_18503);
or U19555 (N_19555,N_18678,N_18077);
or U19556 (N_19556,N_18006,N_18233);
nand U19557 (N_19557,N_18357,N_18646);
nor U19558 (N_19558,N_18181,N_18407);
nor U19559 (N_19559,N_18418,N_18918);
and U19560 (N_19560,N_18758,N_18470);
xor U19561 (N_19561,N_18605,N_18001);
or U19562 (N_19562,N_18746,N_18279);
and U19563 (N_19563,N_18322,N_18919);
and U19564 (N_19564,N_18081,N_18809);
xnor U19565 (N_19565,N_18116,N_18036);
or U19566 (N_19566,N_18737,N_18446);
or U19567 (N_19567,N_18226,N_18803);
and U19568 (N_19568,N_18558,N_18553);
or U19569 (N_19569,N_18032,N_18276);
xnor U19570 (N_19570,N_18585,N_18436);
xor U19571 (N_19571,N_18821,N_18180);
nor U19572 (N_19572,N_18083,N_18369);
or U19573 (N_19573,N_18735,N_18045);
and U19574 (N_19574,N_18689,N_18967);
xor U19575 (N_19575,N_18906,N_18573);
and U19576 (N_19576,N_18058,N_18717);
xnor U19577 (N_19577,N_18372,N_18437);
nor U19578 (N_19578,N_18588,N_18157);
xnor U19579 (N_19579,N_18052,N_18097);
nor U19580 (N_19580,N_18062,N_18059);
xnor U19581 (N_19581,N_18686,N_18336);
nor U19582 (N_19582,N_18302,N_18423);
xor U19583 (N_19583,N_18229,N_18795);
nand U19584 (N_19584,N_18028,N_18082);
and U19585 (N_19585,N_18777,N_18840);
nand U19586 (N_19586,N_18939,N_18420);
and U19587 (N_19587,N_18192,N_18122);
nor U19588 (N_19588,N_18871,N_18666);
nor U19589 (N_19589,N_18603,N_18217);
or U19590 (N_19590,N_18936,N_18316);
xor U19591 (N_19591,N_18264,N_18428);
xnor U19592 (N_19592,N_18788,N_18671);
and U19593 (N_19593,N_18516,N_18442);
and U19594 (N_19594,N_18079,N_18263);
nand U19595 (N_19595,N_18112,N_18172);
nand U19596 (N_19596,N_18460,N_18427);
and U19597 (N_19597,N_18443,N_18861);
and U19598 (N_19598,N_18780,N_18318);
xor U19599 (N_19599,N_18658,N_18547);
or U19600 (N_19600,N_18513,N_18511);
nor U19601 (N_19601,N_18571,N_18925);
and U19602 (N_19602,N_18022,N_18789);
and U19603 (N_19603,N_18953,N_18653);
and U19604 (N_19604,N_18627,N_18118);
and U19605 (N_19605,N_18273,N_18190);
nor U19606 (N_19606,N_18158,N_18649);
or U19607 (N_19607,N_18433,N_18140);
and U19608 (N_19608,N_18581,N_18552);
or U19609 (N_19609,N_18311,N_18600);
and U19610 (N_19610,N_18771,N_18887);
or U19611 (N_19611,N_18493,N_18661);
and U19612 (N_19612,N_18086,N_18649);
nor U19613 (N_19613,N_18729,N_18764);
or U19614 (N_19614,N_18973,N_18752);
or U19615 (N_19615,N_18127,N_18755);
xnor U19616 (N_19616,N_18265,N_18476);
or U19617 (N_19617,N_18501,N_18435);
or U19618 (N_19618,N_18114,N_18166);
or U19619 (N_19619,N_18497,N_18769);
xnor U19620 (N_19620,N_18352,N_18045);
nand U19621 (N_19621,N_18805,N_18892);
nor U19622 (N_19622,N_18236,N_18296);
nor U19623 (N_19623,N_18113,N_18918);
xnor U19624 (N_19624,N_18346,N_18866);
xnor U19625 (N_19625,N_18521,N_18617);
and U19626 (N_19626,N_18209,N_18039);
or U19627 (N_19627,N_18156,N_18470);
xor U19628 (N_19628,N_18038,N_18202);
or U19629 (N_19629,N_18001,N_18656);
or U19630 (N_19630,N_18749,N_18459);
nor U19631 (N_19631,N_18087,N_18140);
nor U19632 (N_19632,N_18463,N_18934);
xnor U19633 (N_19633,N_18177,N_18184);
nor U19634 (N_19634,N_18625,N_18730);
and U19635 (N_19635,N_18519,N_18081);
xnor U19636 (N_19636,N_18209,N_18776);
nand U19637 (N_19637,N_18661,N_18586);
nand U19638 (N_19638,N_18449,N_18956);
or U19639 (N_19639,N_18292,N_18827);
or U19640 (N_19640,N_18766,N_18421);
xnor U19641 (N_19641,N_18514,N_18935);
xor U19642 (N_19642,N_18679,N_18147);
or U19643 (N_19643,N_18935,N_18359);
or U19644 (N_19644,N_18894,N_18153);
or U19645 (N_19645,N_18469,N_18307);
nor U19646 (N_19646,N_18434,N_18351);
or U19647 (N_19647,N_18680,N_18836);
xor U19648 (N_19648,N_18387,N_18272);
xor U19649 (N_19649,N_18218,N_18084);
nor U19650 (N_19650,N_18480,N_18473);
nor U19651 (N_19651,N_18377,N_18780);
nand U19652 (N_19652,N_18941,N_18353);
or U19653 (N_19653,N_18095,N_18092);
xnor U19654 (N_19654,N_18054,N_18715);
nor U19655 (N_19655,N_18953,N_18450);
and U19656 (N_19656,N_18417,N_18064);
nand U19657 (N_19657,N_18684,N_18609);
nand U19658 (N_19658,N_18047,N_18368);
nand U19659 (N_19659,N_18175,N_18222);
and U19660 (N_19660,N_18904,N_18929);
xor U19661 (N_19661,N_18318,N_18813);
xnor U19662 (N_19662,N_18501,N_18070);
or U19663 (N_19663,N_18200,N_18264);
xnor U19664 (N_19664,N_18648,N_18767);
xor U19665 (N_19665,N_18587,N_18714);
nand U19666 (N_19666,N_18739,N_18412);
or U19667 (N_19667,N_18588,N_18204);
and U19668 (N_19668,N_18032,N_18533);
nor U19669 (N_19669,N_18549,N_18218);
or U19670 (N_19670,N_18108,N_18155);
nor U19671 (N_19671,N_18916,N_18024);
and U19672 (N_19672,N_18679,N_18012);
nand U19673 (N_19673,N_18709,N_18176);
nor U19674 (N_19674,N_18536,N_18706);
xnor U19675 (N_19675,N_18787,N_18664);
and U19676 (N_19676,N_18823,N_18278);
nand U19677 (N_19677,N_18278,N_18545);
and U19678 (N_19678,N_18632,N_18468);
or U19679 (N_19679,N_18182,N_18107);
or U19680 (N_19680,N_18598,N_18297);
nand U19681 (N_19681,N_18831,N_18120);
nand U19682 (N_19682,N_18933,N_18670);
nand U19683 (N_19683,N_18247,N_18281);
nand U19684 (N_19684,N_18733,N_18119);
and U19685 (N_19685,N_18743,N_18674);
and U19686 (N_19686,N_18113,N_18356);
nor U19687 (N_19687,N_18988,N_18722);
nor U19688 (N_19688,N_18714,N_18075);
and U19689 (N_19689,N_18555,N_18070);
nand U19690 (N_19690,N_18523,N_18675);
nor U19691 (N_19691,N_18687,N_18157);
xor U19692 (N_19692,N_18478,N_18270);
and U19693 (N_19693,N_18564,N_18692);
or U19694 (N_19694,N_18508,N_18703);
or U19695 (N_19695,N_18236,N_18313);
and U19696 (N_19696,N_18818,N_18660);
and U19697 (N_19697,N_18221,N_18179);
and U19698 (N_19698,N_18712,N_18561);
nor U19699 (N_19699,N_18147,N_18474);
xor U19700 (N_19700,N_18000,N_18109);
and U19701 (N_19701,N_18858,N_18365);
nand U19702 (N_19702,N_18415,N_18481);
xor U19703 (N_19703,N_18622,N_18929);
xnor U19704 (N_19704,N_18668,N_18027);
nor U19705 (N_19705,N_18071,N_18439);
and U19706 (N_19706,N_18385,N_18897);
or U19707 (N_19707,N_18296,N_18314);
xor U19708 (N_19708,N_18586,N_18219);
or U19709 (N_19709,N_18845,N_18475);
and U19710 (N_19710,N_18607,N_18193);
nor U19711 (N_19711,N_18230,N_18279);
nand U19712 (N_19712,N_18817,N_18187);
and U19713 (N_19713,N_18765,N_18048);
nand U19714 (N_19714,N_18156,N_18024);
nor U19715 (N_19715,N_18089,N_18532);
or U19716 (N_19716,N_18492,N_18850);
nor U19717 (N_19717,N_18823,N_18506);
xnor U19718 (N_19718,N_18603,N_18296);
and U19719 (N_19719,N_18525,N_18082);
nand U19720 (N_19720,N_18401,N_18170);
xor U19721 (N_19721,N_18392,N_18500);
and U19722 (N_19722,N_18753,N_18684);
and U19723 (N_19723,N_18010,N_18170);
and U19724 (N_19724,N_18153,N_18889);
or U19725 (N_19725,N_18299,N_18178);
xnor U19726 (N_19726,N_18083,N_18851);
and U19727 (N_19727,N_18804,N_18992);
and U19728 (N_19728,N_18174,N_18747);
xnor U19729 (N_19729,N_18496,N_18744);
or U19730 (N_19730,N_18413,N_18625);
xor U19731 (N_19731,N_18582,N_18075);
and U19732 (N_19732,N_18225,N_18431);
or U19733 (N_19733,N_18892,N_18876);
xor U19734 (N_19734,N_18662,N_18381);
nand U19735 (N_19735,N_18174,N_18470);
nor U19736 (N_19736,N_18612,N_18188);
xor U19737 (N_19737,N_18243,N_18012);
nand U19738 (N_19738,N_18750,N_18044);
nor U19739 (N_19739,N_18666,N_18100);
or U19740 (N_19740,N_18944,N_18516);
nand U19741 (N_19741,N_18398,N_18625);
and U19742 (N_19742,N_18482,N_18654);
and U19743 (N_19743,N_18420,N_18921);
or U19744 (N_19744,N_18741,N_18961);
nand U19745 (N_19745,N_18407,N_18232);
nor U19746 (N_19746,N_18383,N_18986);
xnor U19747 (N_19747,N_18548,N_18917);
or U19748 (N_19748,N_18278,N_18019);
and U19749 (N_19749,N_18144,N_18806);
nand U19750 (N_19750,N_18388,N_18722);
or U19751 (N_19751,N_18584,N_18771);
or U19752 (N_19752,N_18673,N_18801);
or U19753 (N_19753,N_18394,N_18016);
nor U19754 (N_19754,N_18438,N_18740);
or U19755 (N_19755,N_18669,N_18361);
and U19756 (N_19756,N_18270,N_18810);
xnor U19757 (N_19757,N_18966,N_18830);
nand U19758 (N_19758,N_18583,N_18328);
xnor U19759 (N_19759,N_18811,N_18955);
nor U19760 (N_19760,N_18195,N_18114);
nand U19761 (N_19761,N_18546,N_18884);
nand U19762 (N_19762,N_18631,N_18843);
nand U19763 (N_19763,N_18968,N_18976);
nor U19764 (N_19764,N_18128,N_18844);
and U19765 (N_19765,N_18416,N_18139);
nand U19766 (N_19766,N_18830,N_18296);
nand U19767 (N_19767,N_18041,N_18437);
or U19768 (N_19768,N_18714,N_18578);
or U19769 (N_19769,N_18828,N_18577);
nor U19770 (N_19770,N_18182,N_18113);
and U19771 (N_19771,N_18734,N_18018);
or U19772 (N_19772,N_18846,N_18185);
nor U19773 (N_19773,N_18035,N_18234);
xnor U19774 (N_19774,N_18782,N_18957);
and U19775 (N_19775,N_18923,N_18753);
and U19776 (N_19776,N_18411,N_18825);
and U19777 (N_19777,N_18825,N_18175);
xor U19778 (N_19778,N_18082,N_18776);
and U19779 (N_19779,N_18422,N_18193);
and U19780 (N_19780,N_18421,N_18550);
and U19781 (N_19781,N_18732,N_18464);
xnor U19782 (N_19782,N_18958,N_18706);
nor U19783 (N_19783,N_18059,N_18579);
and U19784 (N_19784,N_18898,N_18506);
xor U19785 (N_19785,N_18685,N_18417);
and U19786 (N_19786,N_18592,N_18114);
and U19787 (N_19787,N_18447,N_18595);
nand U19788 (N_19788,N_18842,N_18898);
or U19789 (N_19789,N_18007,N_18346);
nor U19790 (N_19790,N_18567,N_18335);
xor U19791 (N_19791,N_18954,N_18628);
and U19792 (N_19792,N_18064,N_18565);
and U19793 (N_19793,N_18758,N_18673);
and U19794 (N_19794,N_18510,N_18541);
or U19795 (N_19795,N_18812,N_18877);
xor U19796 (N_19796,N_18548,N_18630);
xnor U19797 (N_19797,N_18412,N_18743);
nor U19798 (N_19798,N_18132,N_18635);
nor U19799 (N_19799,N_18087,N_18331);
and U19800 (N_19800,N_18145,N_18493);
and U19801 (N_19801,N_18766,N_18668);
xor U19802 (N_19802,N_18435,N_18304);
and U19803 (N_19803,N_18359,N_18095);
or U19804 (N_19804,N_18095,N_18144);
and U19805 (N_19805,N_18435,N_18110);
or U19806 (N_19806,N_18060,N_18845);
nor U19807 (N_19807,N_18992,N_18165);
or U19808 (N_19808,N_18206,N_18410);
xor U19809 (N_19809,N_18677,N_18347);
and U19810 (N_19810,N_18286,N_18636);
nand U19811 (N_19811,N_18705,N_18914);
xor U19812 (N_19812,N_18208,N_18445);
or U19813 (N_19813,N_18905,N_18723);
xnor U19814 (N_19814,N_18075,N_18929);
nor U19815 (N_19815,N_18438,N_18875);
or U19816 (N_19816,N_18241,N_18374);
xor U19817 (N_19817,N_18025,N_18056);
nand U19818 (N_19818,N_18565,N_18192);
xnor U19819 (N_19819,N_18585,N_18321);
or U19820 (N_19820,N_18811,N_18143);
and U19821 (N_19821,N_18229,N_18973);
or U19822 (N_19822,N_18033,N_18574);
xnor U19823 (N_19823,N_18039,N_18268);
nand U19824 (N_19824,N_18612,N_18671);
nor U19825 (N_19825,N_18120,N_18596);
nor U19826 (N_19826,N_18802,N_18098);
xor U19827 (N_19827,N_18203,N_18070);
nor U19828 (N_19828,N_18772,N_18961);
and U19829 (N_19829,N_18648,N_18512);
nand U19830 (N_19830,N_18911,N_18288);
nand U19831 (N_19831,N_18181,N_18362);
xnor U19832 (N_19832,N_18128,N_18764);
and U19833 (N_19833,N_18606,N_18896);
and U19834 (N_19834,N_18573,N_18885);
nand U19835 (N_19835,N_18072,N_18036);
xnor U19836 (N_19836,N_18665,N_18946);
nor U19837 (N_19837,N_18372,N_18866);
and U19838 (N_19838,N_18845,N_18565);
xnor U19839 (N_19839,N_18443,N_18978);
nand U19840 (N_19840,N_18381,N_18560);
nor U19841 (N_19841,N_18664,N_18559);
nor U19842 (N_19842,N_18940,N_18885);
xor U19843 (N_19843,N_18061,N_18719);
nor U19844 (N_19844,N_18548,N_18776);
or U19845 (N_19845,N_18356,N_18175);
and U19846 (N_19846,N_18139,N_18093);
or U19847 (N_19847,N_18228,N_18148);
nor U19848 (N_19848,N_18514,N_18727);
xor U19849 (N_19849,N_18047,N_18020);
and U19850 (N_19850,N_18279,N_18451);
and U19851 (N_19851,N_18391,N_18745);
nor U19852 (N_19852,N_18952,N_18448);
or U19853 (N_19853,N_18256,N_18072);
or U19854 (N_19854,N_18089,N_18639);
nor U19855 (N_19855,N_18583,N_18551);
and U19856 (N_19856,N_18681,N_18471);
xor U19857 (N_19857,N_18982,N_18658);
nor U19858 (N_19858,N_18668,N_18725);
nor U19859 (N_19859,N_18080,N_18238);
xor U19860 (N_19860,N_18654,N_18547);
or U19861 (N_19861,N_18633,N_18064);
nor U19862 (N_19862,N_18162,N_18582);
nand U19863 (N_19863,N_18465,N_18867);
or U19864 (N_19864,N_18699,N_18252);
nand U19865 (N_19865,N_18825,N_18494);
and U19866 (N_19866,N_18040,N_18951);
nor U19867 (N_19867,N_18276,N_18185);
and U19868 (N_19868,N_18458,N_18954);
or U19869 (N_19869,N_18103,N_18345);
nor U19870 (N_19870,N_18696,N_18529);
or U19871 (N_19871,N_18684,N_18038);
or U19872 (N_19872,N_18109,N_18091);
nor U19873 (N_19873,N_18335,N_18114);
or U19874 (N_19874,N_18071,N_18450);
nand U19875 (N_19875,N_18919,N_18361);
or U19876 (N_19876,N_18793,N_18084);
xor U19877 (N_19877,N_18757,N_18275);
nand U19878 (N_19878,N_18249,N_18665);
nor U19879 (N_19879,N_18266,N_18243);
nand U19880 (N_19880,N_18598,N_18769);
nand U19881 (N_19881,N_18964,N_18212);
nand U19882 (N_19882,N_18038,N_18460);
or U19883 (N_19883,N_18065,N_18823);
or U19884 (N_19884,N_18772,N_18761);
nor U19885 (N_19885,N_18569,N_18996);
xnor U19886 (N_19886,N_18994,N_18097);
nor U19887 (N_19887,N_18370,N_18693);
and U19888 (N_19888,N_18141,N_18948);
and U19889 (N_19889,N_18641,N_18536);
xor U19890 (N_19890,N_18338,N_18944);
nor U19891 (N_19891,N_18090,N_18753);
nand U19892 (N_19892,N_18531,N_18357);
and U19893 (N_19893,N_18183,N_18672);
and U19894 (N_19894,N_18405,N_18966);
xnor U19895 (N_19895,N_18176,N_18752);
nor U19896 (N_19896,N_18962,N_18841);
nand U19897 (N_19897,N_18096,N_18713);
and U19898 (N_19898,N_18374,N_18297);
nor U19899 (N_19899,N_18102,N_18394);
nand U19900 (N_19900,N_18516,N_18526);
and U19901 (N_19901,N_18324,N_18938);
or U19902 (N_19902,N_18672,N_18574);
nand U19903 (N_19903,N_18939,N_18899);
xor U19904 (N_19904,N_18748,N_18736);
nor U19905 (N_19905,N_18775,N_18298);
or U19906 (N_19906,N_18053,N_18327);
or U19907 (N_19907,N_18472,N_18693);
nand U19908 (N_19908,N_18006,N_18719);
nand U19909 (N_19909,N_18304,N_18891);
xor U19910 (N_19910,N_18769,N_18234);
and U19911 (N_19911,N_18812,N_18429);
and U19912 (N_19912,N_18630,N_18687);
and U19913 (N_19913,N_18056,N_18236);
nor U19914 (N_19914,N_18032,N_18162);
nor U19915 (N_19915,N_18330,N_18012);
nor U19916 (N_19916,N_18594,N_18892);
xnor U19917 (N_19917,N_18907,N_18748);
xor U19918 (N_19918,N_18348,N_18066);
nor U19919 (N_19919,N_18214,N_18940);
nand U19920 (N_19920,N_18248,N_18730);
and U19921 (N_19921,N_18084,N_18776);
and U19922 (N_19922,N_18249,N_18817);
xor U19923 (N_19923,N_18939,N_18086);
and U19924 (N_19924,N_18001,N_18485);
or U19925 (N_19925,N_18249,N_18129);
nor U19926 (N_19926,N_18665,N_18463);
and U19927 (N_19927,N_18837,N_18122);
nand U19928 (N_19928,N_18576,N_18134);
xor U19929 (N_19929,N_18692,N_18483);
xor U19930 (N_19930,N_18637,N_18871);
nor U19931 (N_19931,N_18951,N_18596);
xor U19932 (N_19932,N_18615,N_18320);
or U19933 (N_19933,N_18443,N_18815);
or U19934 (N_19934,N_18686,N_18408);
and U19935 (N_19935,N_18358,N_18465);
nand U19936 (N_19936,N_18623,N_18441);
nand U19937 (N_19937,N_18666,N_18508);
xor U19938 (N_19938,N_18522,N_18043);
and U19939 (N_19939,N_18750,N_18017);
or U19940 (N_19940,N_18740,N_18423);
and U19941 (N_19941,N_18959,N_18605);
or U19942 (N_19942,N_18212,N_18707);
nor U19943 (N_19943,N_18219,N_18391);
nand U19944 (N_19944,N_18863,N_18784);
xnor U19945 (N_19945,N_18727,N_18154);
nand U19946 (N_19946,N_18563,N_18205);
nor U19947 (N_19947,N_18207,N_18917);
and U19948 (N_19948,N_18969,N_18246);
or U19949 (N_19949,N_18244,N_18953);
nor U19950 (N_19950,N_18893,N_18362);
xnor U19951 (N_19951,N_18287,N_18485);
and U19952 (N_19952,N_18562,N_18248);
or U19953 (N_19953,N_18960,N_18174);
or U19954 (N_19954,N_18779,N_18332);
or U19955 (N_19955,N_18705,N_18485);
and U19956 (N_19956,N_18853,N_18682);
or U19957 (N_19957,N_18684,N_18060);
or U19958 (N_19958,N_18966,N_18412);
nand U19959 (N_19959,N_18380,N_18309);
nand U19960 (N_19960,N_18142,N_18528);
or U19961 (N_19961,N_18062,N_18775);
nand U19962 (N_19962,N_18545,N_18581);
nor U19963 (N_19963,N_18937,N_18194);
or U19964 (N_19964,N_18732,N_18374);
and U19965 (N_19965,N_18076,N_18892);
xor U19966 (N_19966,N_18386,N_18664);
xor U19967 (N_19967,N_18722,N_18259);
and U19968 (N_19968,N_18455,N_18971);
and U19969 (N_19969,N_18178,N_18149);
or U19970 (N_19970,N_18431,N_18745);
and U19971 (N_19971,N_18823,N_18682);
nor U19972 (N_19972,N_18112,N_18093);
and U19973 (N_19973,N_18539,N_18686);
xnor U19974 (N_19974,N_18859,N_18290);
and U19975 (N_19975,N_18918,N_18788);
xor U19976 (N_19976,N_18887,N_18807);
and U19977 (N_19977,N_18549,N_18782);
nor U19978 (N_19978,N_18540,N_18058);
nand U19979 (N_19979,N_18282,N_18761);
xor U19980 (N_19980,N_18786,N_18650);
nor U19981 (N_19981,N_18923,N_18641);
nand U19982 (N_19982,N_18921,N_18918);
or U19983 (N_19983,N_18517,N_18879);
and U19984 (N_19984,N_18397,N_18135);
or U19985 (N_19985,N_18110,N_18951);
or U19986 (N_19986,N_18126,N_18389);
and U19987 (N_19987,N_18684,N_18411);
and U19988 (N_19988,N_18538,N_18842);
or U19989 (N_19989,N_18392,N_18598);
nand U19990 (N_19990,N_18270,N_18791);
nor U19991 (N_19991,N_18946,N_18048);
nand U19992 (N_19992,N_18907,N_18299);
or U19993 (N_19993,N_18183,N_18083);
or U19994 (N_19994,N_18013,N_18285);
and U19995 (N_19995,N_18501,N_18132);
nor U19996 (N_19996,N_18295,N_18101);
or U19997 (N_19997,N_18047,N_18517);
xor U19998 (N_19998,N_18663,N_18220);
nor U19999 (N_19999,N_18585,N_18264);
nand UO_0 (O_0,N_19636,N_19915);
nand UO_1 (O_1,N_19369,N_19092);
and UO_2 (O_2,N_19564,N_19960);
nor UO_3 (O_3,N_19345,N_19135);
or UO_4 (O_4,N_19941,N_19339);
nor UO_5 (O_5,N_19824,N_19433);
and UO_6 (O_6,N_19166,N_19570);
or UO_7 (O_7,N_19445,N_19540);
nand UO_8 (O_8,N_19759,N_19288);
nor UO_9 (O_9,N_19844,N_19336);
nor UO_10 (O_10,N_19806,N_19925);
and UO_11 (O_11,N_19178,N_19358);
nor UO_12 (O_12,N_19308,N_19627);
and UO_13 (O_13,N_19195,N_19571);
xor UO_14 (O_14,N_19299,N_19306);
or UO_15 (O_15,N_19828,N_19466);
and UO_16 (O_16,N_19689,N_19513);
or UO_17 (O_17,N_19074,N_19041);
xnor UO_18 (O_18,N_19237,N_19714);
xnor UO_19 (O_19,N_19720,N_19892);
xor UO_20 (O_20,N_19938,N_19108);
xnor UO_21 (O_21,N_19088,N_19334);
xnor UO_22 (O_22,N_19644,N_19352);
nand UO_23 (O_23,N_19103,N_19025);
nor UO_24 (O_24,N_19966,N_19728);
nand UO_25 (O_25,N_19527,N_19648);
nand UO_26 (O_26,N_19120,N_19027);
or UO_27 (O_27,N_19590,N_19046);
nor UO_28 (O_28,N_19335,N_19809);
nor UO_29 (O_29,N_19171,N_19457);
nand UO_30 (O_30,N_19896,N_19365);
xor UO_31 (O_31,N_19266,N_19169);
or UO_32 (O_32,N_19899,N_19616);
nor UO_33 (O_33,N_19837,N_19072);
xnor UO_34 (O_34,N_19536,N_19449);
nand UO_35 (O_35,N_19232,N_19501);
and UO_36 (O_36,N_19823,N_19379);
nand UO_37 (O_37,N_19647,N_19185);
or UO_38 (O_38,N_19414,N_19989);
or UO_39 (O_39,N_19579,N_19164);
nor UO_40 (O_40,N_19881,N_19805);
and UO_41 (O_41,N_19957,N_19482);
xnor UO_42 (O_42,N_19642,N_19833);
nor UO_43 (O_43,N_19131,N_19065);
or UO_44 (O_44,N_19381,N_19081);
or UO_45 (O_45,N_19016,N_19286);
xnor UO_46 (O_46,N_19747,N_19196);
xnor UO_47 (O_47,N_19522,N_19276);
nand UO_48 (O_48,N_19786,N_19404);
nor UO_49 (O_49,N_19511,N_19811);
or UO_50 (O_50,N_19771,N_19702);
or UO_51 (O_51,N_19864,N_19859);
nand UO_52 (O_52,N_19946,N_19223);
xnor UO_53 (O_53,N_19145,N_19662);
or UO_54 (O_54,N_19975,N_19450);
nand UO_55 (O_55,N_19594,N_19520);
and UO_56 (O_56,N_19998,N_19492);
nand UO_57 (O_57,N_19338,N_19248);
nand UO_58 (O_58,N_19877,N_19821);
nor UO_59 (O_59,N_19764,N_19854);
and UO_60 (O_60,N_19641,N_19670);
nand UO_61 (O_61,N_19842,N_19437);
nand UO_62 (O_62,N_19183,N_19763);
nor UO_63 (O_63,N_19271,N_19026);
or UO_64 (O_64,N_19436,N_19556);
and UO_65 (O_65,N_19163,N_19224);
xnor UO_66 (O_66,N_19845,N_19242);
nand UO_67 (O_67,N_19875,N_19420);
or UO_68 (O_68,N_19326,N_19121);
nor UO_69 (O_69,N_19878,N_19887);
nand UO_70 (O_70,N_19235,N_19333);
nand UO_71 (O_71,N_19373,N_19405);
or UO_72 (O_72,N_19356,N_19507);
nor UO_73 (O_73,N_19155,N_19487);
nor UO_74 (O_74,N_19253,N_19661);
xnor UO_75 (O_75,N_19058,N_19261);
nand UO_76 (O_76,N_19586,N_19739);
xor UO_77 (O_77,N_19393,N_19531);
nand UO_78 (O_78,N_19200,N_19734);
xnor UO_79 (O_79,N_19459,N_19607);
and UO_80 (O_80,N_19318,N_19073);
and UO_81 (O_81,N_19790,N_19886);
xnor UO_82 (O_82,N_19969,N_19924);
and UO_83 (O_83,N_19988,N_19015);
or UO_84 (O_84,N_19426,N_19853);
nand UO_85 (O_85,N_19417,N_19995);
or UO_86 (O_86,N_19873,N_19340);
or UO_87 (O_87,N_19172,N_19983);
xor UO_88 (O_88,N_19023,N_19767);
xnor UO_89 (O_89,N_19454,N_19865);
nand UO_90 (O_90,N_19495,N_19708);
or UO_91 (O_91,N_19624,N_19766);
or UO_92 (O_92,N_19706,N_19582);
or UO_93 (O_93,N_19186,N_19246);
and UO_94 (O_94,N_19984,N_19421);
nand UO_95 (O_95,N_19785,N_19528);
nand UO_96 (O_96,N_19751,N_19614);
and UO_97 (O_97,N_19305,N_19187);
xnor UO_98 (O_98,N_19604,N_19555);
nor UO_99 (O_99,N_19496,N_19402);
or UO_100 (O_100,N_19001,N_19355);
nand UO_101 (O_101,N_19990,N_19412);
and UO_102 (O_102,N_19578,N_19640);
nor UO_103 (O_103,N_19125,N_19435);
nand UO_104 (O_104,N_19876,N_19226);
or UO_105 (O_105,N_19156,N_19655);
nand UO_106 (O_106,N_19033,N_19699);
or UO_107 (O_107,N_19961,N_19011);
nor UO_108 (O_108,N_19694,N_19711);
xnor UO_109 (O_109,N_19362,N_19572);
or UO_110 (O_110,N_19043,N_19679);
xor UO_111 (O_111,N_19354,N_19122);
nor UO_112 (O_112,N_19064,N_19498);
or UO_113 (O_113,N_19143,N_19879);
nor UO_114 (O_114,N_19230,N_19419);
or UO_115 (O_115,N_19214,N_19037);
xor UO_116 (O_116,N_19028,N_19439);
and UO_117 (O_117,N_19595,N_19533);
nand UO_118 (O_118,N_19050,N_19815);
xor UO_119 (O_119,N_19676,N_19902);
or UO_120 (O_120,N_19472,N_19465);
and UO_121 (O_121,N_19730,N_19542);
nand UO_122 (O_122,N_19740,N_19069);
nand UO_123 (O_123,N_19722,N_19394);
or UO_124 (O_124,N_19021,N_19204);
nor UO_125 (O_125,N_19280,N_19206);
nand UO_126 (O_126,N_19243,N_19525);
and UO_127 (O_127,N_19664,N_19159);
nor UO_128 (O_128,N_19684,N_19950);
xnor UO_129 (O_129,N_19697,N_19703);
nand UO_130 (O_130,N_19347,N_19577);
nand UO_131 (O_131,N_19973,N_19467);
and UO_132 (O_132,N_19723,N_19245);
nor UO_133 (O_133,N_19396,N_19219);
and UO_134 (O_134,N_19448,N_19851);
nand UO_135 (O_135,N_19403,N_19133);
or UO_136 (O_136,N_19871,N_19275);
xor UO_137 (O_137,N_19959,N_19737);
nor UO_138 (O_138,N_19080,N_19372);
nand UO_139 (O_139,N_19812,N_19067);
and UO_140 (O_140,N_19357,N_19735);
or UO_141 (O_141,N_19677,N_19265);
or UO_142 (O_142,N_19621,N_19907);
and UO_143 (O_143,N_19509,N_19314);
xor UO_144 (O_144,N_19068,N_19905);
nand UO_145 (O_145,N_19963,N_19926);
and UO_146 (O_146,N_19227,N_19388);
xnor UO_147 (O_147,N_19429,N_19160);
nor UO_148 (O_148,N_19093,N_19554);
and UO_149 (O_149,N_19650,N_19778);
and UO_150 (O_150,N_19233,N_19004);
nand UO_151 (O_151,N_19053,N_19954);
nor UO_152 (O_152,N_19300,N_19238);
xor UO_153 (O_153,N_19726,N_19416);
nor UO_154 (O_154,N_19094,N_19502);
and UO_155 (O_155,N_19653,N_19635);
and UO_156 (O_156,N_19168,N_19018);
nand UO_157 (O_157,N_19348,N_19493);
or UO_158 (O_158,N_19087,N_19545);
or UO_159 (O_159,N_19193,N_19399);
or UO_160 (O_160,N_19510,N_19070);
xor UO_161 (O_161,N_19217,N_19803);
or UO_162 (O_162,N_19951,N_19468);
nor UO_163 (O_163,N_19408,N_19297);
nor UO_164 (O_164,N_19424,N_19209);
nor UO_165 (O_165,N_19731,N_19190);
nor UO_166 (O_166,N_19631,N_19138);
nor UO_167 (O_167,N_19535,N_19591);
and UO_168 (O_168,N_19425,N_19293);
nor UO_169 (O_169,N_19458,N_19377);
or UO_170 (O_170,N_19789,N_19952);
nor UO_171 (O_171,N_19287,N_19965);
nand UO_172 (O_172,N_19813,N_19745);
nor UO_173 (O_173,N_19110,N_19964);
nor UO_174 (O_174,N_19724,N_19189);
xnor UO_175 (O_175,N_19061,N_19630);
xor UO_176 (O_176,N_19583,N_19587);
or UO_177 (O_177,N_19547,N_19175);
or UO_178 (O_178,N_19982,N_19974);
nand UO_179 (O_179,N_19484,N_19791);
nor UO_180 (O_180,N_19488,N_19343);
or UO_181 (O_181,N_19981,N_19757);
xnor UO_182 (O_182,N_19788,N_19882);
nor UO_183 (O_183,N_19291,N_19258);
nand UO_184 (O_184,N_19210,N_19158);
or UO_185 (O_185,N_19117,N_19868);
or UO_186 (O_186,N_19561,N_19231);
and UO_187 (O_187,N_19274,N_19104);
nor UO_188 (O_188,N_19282,N_19247);
and UO_189 (O_189,N_19096,N_19637);
or UO_190 (O_190,N_19753,N_19508);
nor UO_191 (O_191,N_19667,N_19850);
and UO_192 (O_192,N_19446,N_19341);
or UO_193 (O_193,N_19380,N_19836);
nand UO_194 (O_194,N_19953,N_19756);
and UO_195 (O_195,N_19503,N_19483);
nand UO_196 (O_196,N_19894,N_19784);
nor UO_197 (O_197,N_19898,N_19830);
nor UO_198 (O_198,N_19395,N_19477);
and UO_199 (O_199,N_19364,N_19869);
or UO_200 (O_200,N_19473,N_19652);
xor UO_201 (O_201,N_19566,N_19212);
nor UO_202 (O_202,N_19781,N_19055);
nor UO_203 (O_203,N_19958,N_19968);
xnor UO_204 (O_204,N_19999,N_19177);
and UO_205 (O_205,N_19367,N_19440);
or UO_206 (O_206,N_19792,N_19769);
xnor UO_207 (O_207,N_19447,N_19602);
or UO_208 (O_208,N_19220,N_19285);
and UO_209 (O_209,N_19962,N_19284);
xor UO_210 (O_210,N_19079,N_19328);
and UO_211 (O_211,N_19124,N_19432);
and UO_212 (O_212,N_19497,N_19040);
xor UO_213 (O_213,N_19514,N_19541);
or UO_214 (O_214,N_19304,N_19315);
xnor UO_215 (O_215,N_19024,N_19903);
nand UO_216 (O_216,N_19770,N_19327);
nor UO_217 (O_217,N_19798,N_19197);
nand UO_218 (O_218,N_19323,N_19491);
nand UO_219 (O_219,N_19213,N_19371);
nand UO_220 (O_220,N_19386,N_19229);
or UO_221 (O_221,N_19576,N_19729);
xor UO_222 (O_222,N_19849,N_19060);
and UO_223 (O_223,N_19669,N_19996);
and UO_224 (O_224,N_19049,N_19029);
xnor UO_225 (O_225,N_19783,N_19366);
nand UO_226 (O_226,N_19234,N_19205);
nand UO_227 (O_227,N_19329,N_19565);
and UO_228 (O_228,N_19428,N_19000);
nand UO_229 (O_229,N_19978,N_19066);
nor UO_230 (O_230,N_19776,N_19153);
nor UO_231 (O_231,N_19310,N_19861);
or UO_232 (O_232,N_19062,N_19599);
nand UO_233 (O_233,N_19617,N_19532);
nor UO_234 (O_234,N_19601,N_19504);
or UO_235 (O_235,N_19967,N_19384);
xor UO_236 (O_236,N_19142,N_19934);
or UO_237 (O_237,N_19410,N_19986);
or UO_238 (O_238,N_19361,N_19109);
nand UO_239 (O_239,N_19516,N_19390);
nand UO_240 (O_240,N_19690,N_19738);
and UO_241 (O_241,N_19283,N_19325);
or UO_242 (O_242,N_19866,N_19980);
nand UO_243 (O_243,N_19939,N_19560);
and UO_244 (O_244,N_19262,N_19620);
or UO_245 (O_245,N_19765,N_19649);
nor UO_246 (O_246,N_19317,N_19972);
nor UO_247 (O_247,N_19800,N_19453);
nand UO_248 (O_248,N_19592,N_19331);
xor UO_249 (O_249,N_19613,N_19758);
or UO_250 (O_250,N_19775,N_19919);
nor UO_251 (O_251,N_19481,N_19411);
or UO_252 (O_252,N_19279,N_19059);
and UO_253 (O_253,N_19134,N_19130);
nor UO_254 (O_254,N_19615,N_19949);
and UO_255 (O_255,N_19378,N_19534);
xor UO_256 (O_256,N_19363,N_19779);
or UO_257 (O_257,N_19102,N_19167);
nor UO_258 (O_258,N_19985,N_19312);
xor UO_259 (O_259,N_19744,N_19626);
xor UO_260 (O_260,N_19793,N_19370);
and UO_261 (O_261,N_19840,N_19693);
xnor UO_262 (O_262,N_19834,N_19044);
nor UO_263 (O_263,N_19207,N_19474);
or UO_264 (O_264,N_19398,N_19415);
or UO_265 (O_265,N_19010,N_19893);
or UO_266 (O_266,N_19918,N_19463);
and UO_267 (O_267,N_19895,N_19180);
xor UO_268 (O_268,N_19943,N_19755);
or UO_269 (O_269,N_19741,N_19500);
or UO_270 (O_270,N_19307,N_19682);
and UO_271 (O_271,N_19872,N_19712);
and UO_272 (O_272,N_19904,N_19606);
or UO_273 (O_273,N_19256,N_19643);
xnor UO_274 (O_274,N_19157,N_19888);
or UO_275 (O_275,N_19321,N_19319);
xor UO_276 (O_276,N_19858,N_19132);
xor UO_277 (O_277,N_19530,N_19856);
xor UO_278 (O_278,N_19006,N_19580);
or UO_279 (O_279,N_19376,N_19475);
and UO_280 (O_280,N_19422,N_19151);
and UO_281 (O_281,N_19956,N_19696);
nand UO_282 (O_282,N_19760,N_19870);
xnor UO_283 (O_283,N_19843,N_19320);
nand UO_284 (O_284,N_19499,N_19401);
xnor UO_285 (O_285,N_19936,N_19825);
and UO_286 (O_286,N_19991,N_19077);
and UO_287 (O_287,N_19434,N_19923);
or UO_288 (O_288,N_19115,N_19353);
nor UO_289 (O_289,N_19588,N_19659);
xor UO_290 (O_290,N_19427,N_19311);
nand UO_291 (O_291,N_19807,N_19589);
nand UO_292 (O_292,N_19019,N_19727);
nand UO_293 (O_293,N_19413,N_19063);
or UO_294 (O_294,N_19848,N_19573);
or UO_295 (O_295,N_19937,N_19057);
nor UO_296 (O_296,N_19176,N_19929);
or UO_297 (O_297,N_19820,N_19660);
xnor UO_298 (O_298,N_19819,N_19761);
nand UO_299 (O_299,N_19239,N_19290);
xor UO_300 (O_300,N_19538,N_19099);
and UO_301 (O_301,N_19713,N_19810);
xnor UO_302 (O_302,N_19240,N_19089);
or UO_303 (O_303,N_19835,N_19469);
nand UO_304 (O_304,N_19486,N_19208);
and UO_305 (O_305,N_19148,N_19773);
nor UO_306 (O_306,N_19633,N_19567);
nor UO_307 (O_307,N_19801,N_19608);
nor UO_308 (O_308,N_19717,N_19584);
and UO_309 (O_309,N_19091,N_19078);
xor UO_310 (O_310,N_19368,N_19452);
xnor UO_311 (O_311,N_19748,N_19444);
or UO_312 (O_312,N_19020,N_19997);
nand UO_313 (O_313,N_19149,N_19005);
xnor UO_314 (O_314,N_19298,N_19251);
or UO_315 (O_315,N_19350,N_19154);
xor UO_316 (O_316,N_19909,N_19846);
nor UO_317 (O_317,N_19052,N_19303);
or UO_318 (O_318,N_19485,N_19032);
or UO_319 (O_319,N_19816,N_19831);
or UO_320 (O_320,N_19139,N_19646);
or UO_321 (O_321,N_19970,N_19736);
nor UO_322 (O_322,N_19927,N_19638);
nor UO_323 (O_323,N_19681,N_19012);
xor UO_324 (O_324,N_19478,N_19847);
nor UO_325 (O_325,N_19056,N_19097);
xor UO_326 (O_326,N_19721,N_19818);
nand UO_327 (O_327,N_19855,N_19596);
nor UO_328 (O_328,N_19263,N_19292);
and UO_329 (O_329,N_19656,N_19826);
and UO_330 (O_330,N_19838,N_19182);
or UO_331 (O_331,N_19658,N_19673);
nand UO_332 (O_332,N_19084,N_19241);
nor UO_333 (O_333,N_19129,N_19344);
xor UO_334 (O_334,N_19928,N_19506);
nor UO_335 (O_335,N_19701,N_19922);
nor UO_336 (O_336,N_19575,N_19316);
and UO_337 (O_337,N_19526,N_19460);
or UO_338 (O_338,N_19675,N_19543);
nand UO_339 (O_339,N_19392,N_19645);
nand UO_340 (O_340,N_19715,N_19600);
and UO_341 (O_341,N_19976,N_19391);
xnor UO_342 (O_342,N_19707,N_19628);
xnor UO_343 (O_343,N_19930,N_19101);
nand UO_344 (O_344,N_19215,N_19552);
xor UO_345 (O_345,N_19302,N_19137);
xnor UO_346 (O_346,N_19948,N_19456);
or UO_347 (O_347,N_19244,N_19451);
or UO_348 (O_348,N_19651,N_19857);
nor UO_349 (O_349,N_19423,N_19891);
or UO_350 (O_350,N_19494,N_19455);
nand UO_351 (O_351,N_19272,N_19462);
xor UO_352 (O_352,N_19400,N_19685);
nor UO_353 (O_353,N_19581,N_19931);
xnor UO_354 (O_354,N_19841,N_19085);
xor UO_355 (O_355,N_19523,N_19802);
and UO_356 (O_356,N_19150,N_19709);
xor UO_357 (O_357,N_19932,N_19038);
and UO_358 (O_358,N_19719,N_19118);
nand UO_359 (O_359,N_19654,N_19048);
xor UO_360 (O_360,N_19022,N_19442);
xor UO_361 (O_361,N_19794,N_19752);
xor UO_362 (O_362,N_19106,N_19553);
nor UO_363 (O_363,N_19671,N_19519);
nand UO_364 (O_364,N_19116,N_19464);
and UO_365 (O_365,N_19035,N_19281);
nand UO_366 (O_366,N_19700,N_19075);
and UO_367 (O_367,N_19249,N_19916);
xor UO_368 (O_368,N_19268,N_19095);
nand UO_369 (O_369,N_19112,N_19550);
nor UO_370 (O_370,N_19598,N_19750);
nand UO_371 (O_371,N_19252,N_19539);
nor UO_372 (O_372,N_19165,N_19746);
or UO_373 (O_373,N_19170,N_19912);
or UO_374 (O_374,N_19942,N_19612);
nor UO_375 (O_375,N_19625,N_19430);
nand UO_376 (O_376,N_19202,N_19585);
or UO_377 (O_377,N_19780,N_19549);
xor UO_378 (O_378,N_19222,N_19762);
and UO_379 (O_379,N_19971,N_19198);
nor UO_380 (O_380,N_19236,N_19774);
and UO_381 (O_381,N_19639,N_19313);
nand UO_382 (O_382,N_19147,N_19407);
nand UO_383 (O_383,N_19688,N_19349);
and UO_384 (O_384,N_19476,N_19610);
xnor UO_385 (O_385,N_19874,N_19623);
nor UO_386 (O_386,N_19322,N_19128);
xnor UO_387 (O_387,N_19885,N_19161);
or UO_388 (O_388,N_19889,N_19505);
or UO_389 (O_389,N_19397,N_19013);
and UO_390 (O_390,N_19277,N_19901);
or UO_391 (O_391,N_19622,N_19977);
xor UO_392 (O_392,N_19039,N_19742);
xor UO_393 (O_393,N_19090,N_19920);
or UO_394 (O_394,N_19832,N_19324);
nor UO_395 (O_395,N_19225,N_19839);
nand UO_396 (O_396,N_19569,N_19441);
or UO_397 (O_397,N_19346,N_19228);
nand UO_398 (O_398,N_19017,N_19192);
nand UO_399 (O_399,N_19668,N_19955);
nor UO_400 (O_400,N_19443,N_19705);
nand UO_401 (O_401,N_19203,N_19890);
nand UO_402 (O_402,N_19933,N_19883);
nor UO_403 (O_403,N_19211,N_19007);
nor UO_404 (O_404,N_19768,N_19559);
xnor UO_405 (O_405,N_19674,N_19083);
or UO_406 (O_406,N_19273,N_19524);
nand UO_407 (O_407,N_19777,N_19993);
and UO_408 (O_408,N_19471,N_19257);
xnor UO_409 (O_409,N_19817,N_19489);
or UO_410 (O_410,N_19908,N_19382);
nor UO_411 (O_411,N_19030,N_19294);
xor UO_412 (O_412,N_19014,N_19808);
xnor UO_413 (O_413,N_19557,N_19518);
nand UO_414 (O_414,N_19611,N_19860);
nor UO_415 (O_415,N_19609,N_19900);
xnor UO_416 (O_416,N_19051,N_19521);
or UO_417 (O_417,N_19672,N_19710);
xnor UO_418 (O_418,N_19698,N_19127);
nand UO_419 (O_419,N_19034,N_19296);
and UO_420 (O_420,N_19692,N_19619);
and UO_421 (O_421,N_19935,N_19944);
nor UO_422 (O_422,N_19255,N_19733);
xor UO_423 (O_423,N_19666,N_19054);
nor UO_424 (O_424,N_19086,N_19605);
nor UO_425 (O_425,N_19512,N_19259);
nand UO_426 (O_426,N_19409,N_19537);
or UO_427 (O_427,N_19544,N_19634);
nor UO_428 (O_428,N_19827,N_19782);
xnor UO_429 (O_429,N_19517,N_19678);
and UO_430 (O_430,N_19479,N_19852);
xor UO_431 (O_431,N_19278,N_19480);
nor UO_432 (O_432,N_19470,N_19260);
nor UO_433 (O_433,N_19359,N_19330);
and UO_434 (O_434,N_19822,N_19686);
and UO_435 (O_435,N_19141,N_19191);
nor UO_436 (O_436,N_19880,N_19114);
and UO_437 (O_437,N_19105,N_19490);
nand UO_438 (O_438,N_19795,N_19267);
and UO_439 (O_439,N_19250,N_19188);
and UO_440 (O_440,N_19657,N_19665);
nand UO_441 (O_441,N_19629,N_19140);
or UO_442 (O_442,N_19289,N_19546);
nor UO_443 (O_443,N_19152,N_19732);
nand UO_444 (O_444,N_19914,N_19515);
or UO_445 (O_445,N_19144,N_19716);
xor UO_446 (O_446,N_19829,N_19337);
xnor UO_447 (O_447,N_19031,N_19562);
nand UO_448 (O_448,N_19917,N_19418);
and UO_449 (O_449,N_19797,N_19375);
nor UO_450 (O_450,N_19563,N_19618);
nand UO_451 (O_451,N_19680,N_19867);
and UO_452 (O_452,N_19173,N_19295);
and UO_453 (O_453,N_19979,N_19431);
nand UO_454 (O_454,N_19725,N_19695);
nand UO_455 (O_455,N_19913,N_19663);
or UO_456 (O_456,N_19179,N_19691);
nor UO_457 (O_457,N_19574,N_19568);
nor UO_458 (O_458,N_19360,N_19111);
and UO_459 (O_459,N_19270,N_19593);
or UO_460 (O_460,N_19749,N_19383);
nor UO_461 (O_461,N_19199,N_19438);
or UO_462 (O_462,N_19184,N_19558);
or UO_463 (O_463,N_19113,N_19548);
nor UO_464 (O_464,N_19863,N_19107);
and UO_465 (O_465,N_19921,N_19126);
and UO_466 (O_466,N_19632,N_19146);
nand UO_467 (O_467,N_19754,N_19987);
xor UO_468 (O_468,N_19772,N_19906);
xnor UO_469 (O_469,N_19897,N_19461);
nand UO_470 (O_470,N_19342,N_19136);
or UO_471 (O_471,N_19045,N_19718);
nand UO_472 (O_472,N_19597,N_19123);
or UO_473 (O_473,N_19814,N_19194);
nor UO_474 (O_474,N_19269,N_19008);
and UO_475 (O_475,N_19076,N_19201);
and UO_476 (O_476,N_19351,N_19221);
and UO_477 (O_477,N_19009,N_19992);
and UO_478 (O_478,N_19603,N_19910);
xor UO_479 (O_479,N_19862,N_19799);
or UO_480 (O_480,N_19254,N_19551);
or UO_481 (O_481,N_19100,N_19218);
xor UO_482 (O_482,N_19385,N_19264);
or UO_483 (O_483,N_19940,N_19332);
and UO_484 (O_484,N_19387,N_19994);
nor UO_485 (O_485,N_19174,N_19743);
xnor UO_486 (O_486,N_19947,N_19301);
nor UO_487 (O_487,N_19529,N_19374);
nand UO_488 (O_488,N_19082,N_19047);
xnor UO_489 (O_489,N_19787,N_19042);
xor UO_490 (O_490,N_19704,N_19406);
nor UO_491 (O_491,N_19687,N_19945);
and UO_492 (O_492,N_19309,N_19003);
nor UO_493 (O_493,N_19911,N_19804);
nand UO_494 (O_494,N_19216,N_19884);
and UO_495 (O_495,N_19683,N_19036);
nor UO_496 (O_496,N_19119,N_19389);
nand UO_497 (O_497,N_19071,N_19098);
nand UO_498 (O_498,N_19162,N_19796);
and UO_499 (O_499,N_19002,N_19181);
nand UO_500 (O_500,N_19719,N_19504);
and UO_501 (O_501,N_19602,N_19032);
and UO_502 (O_502,N_19658,N_19482);
nor UO_503 (O_503,N_19289,N_19993);
nand UO_504 (O_504,N_19948,N_19290);
or UO_505 (O_505,N_19490,N_19145);
nor UO_506 (O_506,N_19083,N_19953);
nor UO_507 (O_507,N_19081,N_19324);
or UO_508 (O_508,N_19518,N_19398);
or UO_509 (O_509,N_19083,N_19031);
nand UO_510 (O_510,N_19556,N_19481);
nand UO_511 (O_511,N_19110,N_19721);
nand UO_512 (O_512,N_19960,N_19281);
or UO_513 (O_513,N_19781,N_19753);
and UO_514 (O_514,N_19836,N_19330);
or UO_515 (O_515,N_19552,N_19287);
nor UO_516 (O_516,N_19639,N_19405);
nand UO_517 (O_517,N_19009,N_19287);
nand UO_518 (O_518,N_19160,N_19616);
and UO_519 (O_519,N_19094,N_19851);
nand UO_520 (O_520,N_19097,N_19010);
nand UO_521 (O_521,N_19674,N_19055);
xor UO_522 (O_522,N_19592,N_19783);
xnor UO_523 (O_523,N_19838,N_19517);
nor UO_524 (O_524,N_19706,N_19595);
xnor UO_525 (O_525,N_19252,N_19541);
nor UO_526 (O_526,N_19163,N_19985);
and UO_527 (O_527,N_19905,N_19240);
nor UO_528 (O_528,N_19962,N_19082);
or UO_529 (O_529,N_19932,N_19487);
or UO_530 (O_530,N_19393,N_19509);
xnor UO_531 (O_531,N_19311,N_19558);
and UO_532 (O_532,N_19687,N_19226);
xnor UO_533 (O_533,N_19091,N_19930);
and UO_534 (O_534,N_19605,N_19309);
and UO_535 (O_535,N_19734,N_19513);
or UO_536 (O_536,N_19452,N_19930);
xnor UO_537 (O_537,N_19269,N_19390);
and UO_538 (O_538,N_19940,N_19340);
nor UO_539 (O_539,N_19435,N_19740);
or UO_540 (O_540,N_19959,N_19876);
and UO_541 (O_541,N_19910,N_19386);
and UO_542 (O_542,N_19682,N_19602);
and UO_543 (O_543,N_19852,N_19567);
nor UO_544 (O_544,N_19455,N_19100);
nand UO_545 (O_545,N_19101,N_19661);
and UO_546 (O_546,N_19250,N_19610);
nand UO_547 (O_547,N_19548,N_19585);
xor UO_548 (O_548,N_19234,N_19064);
or UO_549 (O_549,N_19622,N_19489);
and UO_550 (O_550,N_19663,N_19661);
nand UO_551 (O_551,N_19712,N_19169);
or UO_552 (O_552,N_19984,N_19847);
and UO_553 (O_553,N_19595,N_19509);
nand UO_554 (O_554,N_19995,N_19286);
or UO_555 (O_555,N_19085,N_19649);
nor UO_556 (O_556,N_19602,N_19109);
nand UO_557 (O_557,N_19617,N_19517);
nand UO_558 (O_558,N_19319,N_19704);
or UO_559 (O_559,N_19609,N_19434);
and UO_560 (O_560,N_19837,N_19174);
xnor UO_561 (O_561,N_19320,N_19910);
and UO_562 (O_562,N_19638,N_19177);
and UO_563 (O_563,N_19737,N_19332);
xor UO_564 (O_564,N_19654,N_19832);
nor UO_565 (O_565,N_19209,N_19467);
and UO_566 (O_566,N_19629,N_19356);
or UO_567 (O_567,N_19062,N_19671);
and UO_568 (O_568,N_19209,N_19577);
or UO_569 (O_569,N_19722,N_19420);
xor UO_570 (O_570,N_19836,N_19446);
nor UO_571 (O_571,N_19440,N_19319);
nand UO_572 (O_572,N_19942,N_19304);
or UO_573 (O_573,N_19020,N_19461);
or UO_574 (O_574,N_19467,N_19625);
nor UO_575 (O_575,N_19427,N_19622);
and UO_576 (O_576,N_19580,N_19513);
or UO_577 (O_577,N_19424,N_19914);
and UO_578 (O_578,N_19410,N_19518);
and UO_579 (O_579,N_19492,N_19737);
xnor UO_580 (O_580,N_19782,N_19170);
nand UO_581 (O_581,N_19559,N_19639);
nand UO_582 (O_582,N_19952,N_19222);
or UO_583 (O_583,N_19051,N_19189);
xnor UO_584 (O_584,N_19384,N_19932);
nand UO_585 (O_585,N_19998,N_19559);
xnor UO_586 (O_586,N_19372,N_19834);
or UO_587 (O_587,N_19765,N_19807);
and UO_588 (O_588,N_19116,N_19189);
xnor UO_589 (O_589,N_19899,N_19785);
xor UO_590 (O_590,N_19855,N_19571);
and UO_591 (O_591,N_19679,N_19255);
or UO_592 (O_592,N_19055,N_19899);
nor UO_593 (O_593,N_19848,N_19041);
xnor UO_594 (O_594,N_19062,N_19557);
and UO_595 (O_595,N_19198,N_19317);
and UO_596 (O_596,N_19189,N_19026);
and UO_597 (O_597,N_19678,N_19934);
or UO_598 (O_598,N_19346,N_19107);
xnor UO_599 (O_599,N_19684,N_19696);
and UO_600 (O_600,N_19702,N_19742);
nand UO_601 (O_601,N_19991,N_19491);
and UO_602 (O_602,N_19186,N_19237);
xor UO_603 (O_603,N_19685,N_19604);
xor UO_604 (O_604,N_19058,N_19548);
nor UO_605 (O_605,N_19536,N_19096);
or UO_606 (O_606,N_19883,N_19824);
or UO_607 (O_607,N_19943,N_19561);
or UO_608 (O_608,N_19023,N_19468);
or UO_609 (O_609,N_19310,N_19417);
xor UO_610 (O_610,N_19616,N_19114);
nor UO_611 (O_611,N_19691,N_19675);
nand UO_612 (O_612,N_19810,N_19842);
or UO_613 (O_613,N_19245,N_19460);
and UO_614 (O_614,N_19245,N_19452);
nand UO_615 (O_615,N_19324,N_19139);
or UO_616 (O_616,N_19958,N_19262);
xnor UO_617 (O_617,N_19385,N_19011);
nor UO_618 (O_618,N_19795,N_19469);
and UO_619 (O_619,N_19675,N_19373);
nand UO_620 (O_620,N_19005,N_19018);
xor UO_621 (O_621,N_19480,N_19619);
and UO_622 (O_622,N_19772,N_19968);
nor UO_623 (O_623,N_19088,N_19340);
nor UO_624 (O_624,N_19574,N_19608);
xnor UO_625 (O_625,N_19648,N_19939);
or UO_626 (O_626,N_19109,N_19029);
nand UO_627 (O_627,N_19693,N_19698);
or UO_628 (O_628,N_19720,N_19239);
nor UO_629 (O_629,N_19498,N_19298);
xor UO_630 (O_630,N_19917,N_19956);
nor UO_631 (O_631,N_19511,N_19418);
xor UO_632 (O_632,N_19621,N_19803);
nor UO_633 (O_633,N_19490,N_19628);
nor UO_634 (O_634,N_19977,N_19290);
xor UO_635 (O_635,N_19529,N_19011);
nand UO_636 (O_636,N_19336,N_19809);
or UO_637 (O_637,N_19563,N_19721);
and UO_638 (O_638,N_19349,N_19478);
and UO_639 (O_639,N_19824,N_19902);
or UO_640 (O_640,N_19035,N_19623);
nand UO_641 (O_641,N_19623,N_19917);
and UO_642 (O_642,N_19864,N_19213);
nor UO_643 (O_643,N_19527,N_19928);
nor UO_644 (O_644,N_19474,N_19729);
nor UO_645 (O_645,N_19648,N_19770);
and UO_646 (O_646,N_19250,N_19574);
nand UO_647 (O_647,N_19006,N_19245);
and UO_648 (O_648,N_19930,N_19312);
nor UO_649 (O_649,N_19183,N_19864);
xor UO_650 (O_650,N_19651,N_19679);
xnor UO_651 (O_651,N_19962,N_19835);
and UO_652 (O_652,N_19984,N_19481);
nand UO_653 (O_653,N_19672,N_19731);
nand UO_654 (O_654,N_19215,N_19540);
or UO_655 (O_655,N_19613,N_19936);
xor UO_656 (O_656,N_19509,N_19880);
xor UO_657 (O_657,N_19506,N_19698);
nor UO_658 (O_658,N_19973,N_19735);
and UO_659 (O_659,N_19948,N_19907);
or UO_660 (O_660,N_19731,N_19332);
nor UO_661 (O_661,N_19867,N_19013);
nor UO_662 (O_662,N_19848,N_19917);
nand UO_663 (O_663,N_19897,N_19725);
or UO_664 (O_664,N_19514,N_19530);
or UO_665 (O_665,N_19838,N_19902);
nor UO_666 (O_666,N_19918,N_19236);
nor UO_667 (O_667,N_19017,N_19868);
or UO_668 (O_668,N_19135,N_19780);
and UO_669 (O_669,N_19055,N_19986);
or UO_670 (O_670,N_19464,N_19697);
xor UO_671 (O_671,N_19625,N_19429);
nand UO_672 (O_672,N_19307,N_19755);
xnor UO_673 (O_673,N_19772,N_19710);
and UO_674 (O_674,N_19981,N_19426);
xnor UO_675 (O_675,N_19308,N_19402);
nand UO_676 (O_676,N_19564,N_19128);
nand UO_677 (O_677,N_19161,N_19707);
xnor UO_678 (O_678,N_19601,N_19139);
nor UO_679 (O_679,N_19964,N_19140);
xnor UO_680 (O_680,N_19647,N_19926);
xnor UO_681 (O_681,N_19440,N_19937);
or UO_682 (O_682,N_19515,N_19832);
xor UO_683 (O_683,N_19853,N_19814);
nor UO_684 (O_684,N_19750,N_19027);
or UO_685 (O_685,N_19750,N_19570);
xor UO_686 (O_686,N_19963,N_19837);
nor UO_687 (O_687,N_19688,N_19062);
and UO_688 (O_688,N_19836,N_19682);
xnor UO_689 (O_689,N_19508,N_19916);
nand UO_690 (O_690,N_19018,N_19469);
nand UO_691 (O_691,N_19586,N_19548);
xor UO_692 (O_692,N_19887,N_19809);
nor UO_693 (O_693,N_19461,N_19842);
xnor UO_694 (O_694,N_19175,N_19753);
and UO_695 (O_695,N_19740,N_19425);
or UO_696 (O_696,N_19308,N_19038);
xor UO_697 (O_697,N_19068,N_19347);
nand UO_698 (O_698,N_19827,N_19761);
xnor UO_699 (O_699,N_19779,N_19228);
and UO_700 (O_700,N_19829,N_19862);
and UO_701 (O_701,N_19448,N_19632);
nand UO_702 (O_702,N_19143,N_19043);
and UO_703 (O_703,N_19069,N_19774);
and UO_704 (O_704,N_19435,N_19612);
or UO_705 (O_705,N_19411,N_19256);
nor UO_706 (O_706,N_19147,N_19544);
nor UO_707 (O_707,N_19710,N_19666);
xnor UO_708 (O_708,N_19685,N_19017);
nand UO_709 (O_709,N_19352,N_19168);
nand UO_710 (O_710,N_19168,N_19089);
nor UO_711 (O_711,N_19808,N_19362);
and UO_712 (O_712,N_19795,N_19897);
xnor UO_713 (O_713,N_19681,N_19989);
or UO_714 (O_714,N_19546,N_19433);
nand UO_715 (O_715,N_19058,N_19242);
or UO_716 (O_716,N_19452,N_19663);
xor UO_717 (O_717,N_19172,N_19729);
xnor UO_718 (O_718,N_19196,N_19528);
nor UO_719 (O_719,N_19100,N_19573);
and UO_720 (O_720,N_19722,N_19969);
or UO_721 (O_721,N_19860,N_19300);
or UO_722 (O_722,N_19864,N_19687);
and UO_723 (O_723,N_19547,N_19026);
xnor UO_724 (O_724,N_19148,N_19923);
or UO_725 (O_725,N_19540,N_19656);
or UO_726 (O_726,N_19931,N_19877);
and UO_727 (O_727,N_19053,N_19261);
xor UO_728 (O_728,N_19771,N_19038);
xor UO_729 (O_729,N_19896,N_19318);
and UO_730 (O_730,N_19914,N_19694);
nand UO_731 (O_731,N_19438,N_19550);
xor UO_732 (O_732,N_19821,N_19521);
xnor UO_733 (O_733,N_19275,N_19980);
nand UO_734 (O_734,N_19249,N_19974);
and UO_735 (O_735,N_19551,N_19216);
nand UO_736 (O_736,N_19552,N_19806);
nor UO_737 (O_737,N_19918,N_19888);
xor UO_738 (O_738,N_19865,N_19136);
nand UO_739 (O_739,N_19465,N_19650);
and UO_740 (O_740,N_19744,N_19390);
nand UO_741 (O_741,N_19599,N_19662);
and UO_742 (O_742,N_19325,N_19253);
nor UO_743 (O_743,N_19434,N_19463);
and UO_744 (O_744,N_19938,N_19951);
nand UO_745 (O_745,N_19997,N_19560);
or UO_746 (O_746,N_19416,N_19366);
and UO_747 (O_747,N_19187,N_19283);
nand UO_748 (O_748,N_19428,N_19467);
nor UO_749 (O_749,N_19868,N_19115);
nand UO_750 (O_750,N_19687,N_19192);
nor UO_751 (O_751,N_19759,N_19143);
nand UO_752 (O_752,N_19790,N_19259);
or UO_753 (O_753,N_19770,N_19875);
nand UO_754 (O_754,N_19280,N_19881);
nand UO_755 (O_755,N_19594,N_19366);
xor UO_756 (O_756,N_19209,N_19578);
or UO_757 (O_757,N_19421,N_19988);
or UO_758 (O_758,N_19762,N_19728);
and UO_759 (O_759,N_19906,N_19352);
nor UO_760 (O_760,N_19229,N_19935);
and UO_761 (O_761,N_19077,N_19506);
and UO_762 (O_762,N_19407,N_19367);
or UO_763 (O_763,N_19956,N_19535);
xnor UO_764 (O_764,N_19166,N_19291);
and UO_765 (O_765,N_19199,N_19787);
nand UO_766 (O_766,N_19926,N_19861);
nand UO_767 (O_767,N_19737,N_19504);
nor UO_768 (O_768,N_19669,N_19702);
or UO_769 (O_769,N_19602,N_19776);
or UO_770 (O_770,N_19627,N_19182);
xor UO_771 (O_771,N_19178,N_19136);
nor UO_772 (O_772,N_19360,N_19793);
nor UO_773 (O_773,N_19672,N_19680);
and UO_774 (O_774,N_19236,N_19805);
or UO_775 (O_775,N_19115,N_19364);
nand UO_776 (O_776,N_19151,N_19067);
nand UO_777 (O_777,N_19035,N_19246);
nor UO_778 (O_778,N_19234,N_19309);
nor UO_779 (O_779,N_19038,N_19280);
nor UO_780 (O_780,N_19848,N_19118);
xor UO_781 (O_781,N_19248,N_19935);
nand UO_782 (O_782,N_19760,N_19960);
nand UO_783 (O_783,N_19911,N_19209);
or UO_784 (O_784,N_19993,N_19009);
nand UO_785 (O_785,N_19928,N_19703);
and UO_786 (O_786,N_19877,N_19516);
xnor UO_787 (O_787,N_19620,N_19613);
or UO_788 (O_788,N_19119,N_19285);
and UO_789 (O_789,N_19515,N_19907);
and UO_790 (O_790,N_19905,N_19392);
and UO_791 (O_791,N_19912,N_19839);
nand UO_792 (O_792,N_19434,N_19870);
or UO_793 (O_793,N_19563,N_19434);
xor UO_794 (O_794,N_19215,N_19140);
or UO_795 (O_795,N_19732,N_19194);
or UO_796 (O_796,N_19126,N_19069);
xnor UO_797 (O_797,N_19700,N_19632);
nand UO_798 (O_798,N_19758,N_19724);
or UO_799 (O_799,N_19484,N_19722);
xnor UO_800 (O_800,N_19275,N_19078);
or UO_801 (O_801,N_19481,N_19937);
or UO_802 (O_802,N_19034,N_19253);
and UO_803 (O_803,N_19632,N_19572);
nor UO_804 (O_804,N_19963,N_19583);
and UO_805 (O_805,N_19393,N_19590);
nand UO_806 (O_806,N_19656,N_19017);
xor UO_807 (O_807,N_19637,N_19802);
or UO_808 (O_808,N_19444,N_19532);
or UO_809 (O_809,N_19224,N_19631);
or UO_810 (O_810,N_19406,N_19549);
nor UO_811 (O_811,N_19142,N_19882);
or UO_812 (O_812,N_19153,N_19625);
or UO_813 (O_813,N_19976,N_19718);
xnor UO_814 (O_814,N_19631,N_19241);
nor UO_815 (O_815,N_19732,N_19613);
nand UO_816 (O_816,N_19772,N_19576);
or UO_817 (O_817,N_19782,N_19793);
nand UO_818 (O_818,N_19083,N_19419);
nor UO_819 (O_819,N_19026,N_19482);
or UO_820 (O_820,N_19025,N_19836);
and UO_821 (O_821,N_19241,N_19393);
or UO_822 (O_822,N_19521,N_19910);
xnor UO_823 (O_823,N_19112,N_19070);
xor UO_824 (O_824,N_19650,N_19186);
xor UO_825 (O_825,N_19882,N_19969);
nand UO_826 (O_826,N_19215,N_19590);
nand UO_827 (O_827,N_19647,N_19348);
nand UO_828 (O_828,N_19749,N_19242);
xor UO_829 (O_829,N_19138,N_19452);
or UO_830 (O_830,N_19097,N_19091);
nand UO_831 (O_831,N_19007,N_19240);
or UO_832 (O_832,N_19599,N_19637);
nand UO_833 (O_833,N_19733,N_19522);
nor UO_834 (O_834,N_19899,N_19235);
xnor UO_835 (O_835,N_19121,N_19730);
xor UO_836 (O_836,N_19795,N_19446);
nand UO_837 (O_837,N_19800,N_19991);
or UO_838 (O_838,N_19967,N_19961);
and UO_839 (O_839,N_19698,N_19769);
xnor UO_840 (O_840,N_19700,N_19946);
or UO_841 (O_841,N_19528,N_19418);
or UO_842 (O_842,N_19522,N_19722);
nand UO_843 (O_843,N_19748,N_19837);
xor UO_844 (O_844,N_19463,N_19315);
nor UO_845 (O_845,N_19490,N_19118);
nor UO_846 (O_846,N_19582,N_19796);
xnor UO_847 (O_847,N_19718,N_19346);
and UO_848 (O_848,N_19661,N_19902);
nand UO_849 (O_849,N_19923,N_19309);
and UO_850 (O_850,N_19485,N_19456);
or UO_851 (O_851,N_19205,N_19941);
nand UO_852 (O_852,N_19602,N_19067);
or UO_853 (O_853,N_19262,N_19780);
nand UO_854 (O_854,N_19673,N_19512);
or UO_855 (O_855,N_19241,N_19443);
and UO_856 (O_856,N_19440,N_19014);
and UO_857 (O_857,N_19379,N_19368);
and UO_858 (O_858,N_19008,N_19828);
and UO_859 (O_859,N_19549,N_19123);
and UO_860 (O_860,N_19386,N_19543);
and UO_861 (O_861,N_19318,N_19911);
or UO_862 (O_862,N_19379,N_19473);
nor UO_863 (O_863,N_19297,N_19758);
nand UO_864 (O_864,N_19318,N_19118);
nor UO_865 (O_865,N_19276,N_19160);
nor UO_866 (O_866,N_19588,N_19946);
nand UO_867 (O_867,N_19211,N_19791);
nor UO_868 (O_868,N_19605,N_19274);
nor UO_869 (O_869,N_19243,N_19480);
xnor UO_870 (O_870,N_19695,N_19032);
and UO_871 (O_871,N_19276,N_19915);
xnor UO_872 (O_872,N_19635,N_19698);
and UO_873 (O_873,N_19741,N_19647);
xor UO_874 (O_874,N_19899,N_19102);
xor UO_875 (O_875,N_19812,N_19905);
nor UO_876 (O_876,N_19563,N_19655);
nor UO_877 (O_877,N_19427,N_19610);
nand UO_878 (O_878,N_19438,N_19009);
or UO_879 (O_879,N_19821,N_19680);
nor UO_880 (O_880,N_19894,N_19216);
nand UO_881 (O_881,N_19300,N_19276);
xor UO_882 (O_882,N_19523,N_19909);
and UO_883 (O_883,N_19178,N_19624);
and UO_884 (O_884,N_19092,N_19815);
nor UO_885 (O_885,N_19620,N_19002);
or UO_886 (O_886,N_19934,N_19140);
nor UO_887 (O_887,N_19351,N_19793);
and UO_888 (O_888,N_19586,N_19019);
and UO_889 (O_889,N_19060,N_19435);
and UO_890 (O_890,N_19888,N_19493);
xor UO_891 (O_891,N_19414,N_19190);
or UO_892 (O_892,N_19426,N_19772);
nor UO_893 (O_893,N_19711,N_19987);
xor UO_894 (O_894,N_19505,N_19974);
and UO_895 (O_895,N_19223,N_19879);
or UO_896 (O_896,N_19613,N_19587);
xor UO_897 (O_897,N_19250,N_19013);
and UO_898 (O_898,N_19439,N_19144);
nor UO_899 (O_899,N_19191,N_19573);
nor UO_900 (O_900,N_19041,N_19772);
and UO_901 (O_901,N_19395,N_19692);
xnor UO_902 (O_902,N_19729,N_19355);
xor UO_903 (O_903,N_19976,N_19111);
nand UO_904 (O_904,N_19670,N_19342);
and UO_905 (O_905,N_19746,N_19235);
xor UO_906 (O_906,N_19944,N_19235);
xor UO_907 (O_907,N_19410,N_19359);
and UO_908 (O_908,N_19833,N_19001);
nand UO_909 (O_909,N_19613,N_19244);
or UO_910 (O_910,N_19438,N_19714);
or UO_911 (O_911,N_19673,N_19808);
and UO_912 (O_912,N_19814,N_19520);
nand UO_913 (O_913,N_19234,N_19134);
and UO_914 (O_914,N_19141,N_19442);
or UO_915 (O_915,N_19952,N_19301);
xnor UO_916 (O_916,N_19394,N_19442);
and UO_917 (O_917,N_19399,N_19274);
xnor UO_918 (O_918,N_19082,N_19770);
nor UO_919 (O_919,N_19211,N_19436);
nand UO_920 (O_920,N_19041,N_19818);
and UO_921 (O_921,N_19869,N_19294);
nand UO_922 (O_922,N_19550,N_19624);
nor UO_923 (O_923,N_19428,N_19857);
nor UO_924 (O_924,N_19565,N_19299);
xor UO_925 (O_925,N_19214,N_19234);
nor UO_926 (O_926,N_19503,N_19007);
or UO_927 (O_927,N_19664,N_19626);
and UO_928 (O_928,N_19226,N_19578);
nor UO_929 (O_929,N_19519,N_19535);
nor UO_930 (O_930,N_19954,N_19317);
xnor UO_931 (O_931,N_19477,N_19129);
or UO_932 (O_932,N_19789,N_19044);
nand UO_933 (O_933,N_19134,N_19450);
nand UO_934 (O_934,N_19179,N_19771);
nor UO_935 (O_935,N_19371,N_19272);
and UO_936 (O_936,N_19112,N_19356);
xnor UO_937 (O_937,N_19632,N_19472);
or UO_938 (O_938,N_19188,N_19754);
xor UO_939 (O_939,N_19961,N_19464);
and UO_940 (O_940,N_19063,N_19765);
nand UO_941 (O_941,N_19009,N_19636);
nand UO_942 (O_942,N_19291,N_19158);
and UO_943 (O_943,N_19180,N_19172);
nand UO_944 (O_944,N_19083,N_19347);
and UO_945 (O_945,N_19915,N_19876);
nor UO_946 (O_946,N_19879,N_19944);
and UO_947 (O_947,N_19258,N_19646);
nor UO_948 (O_948,N_19805,N_19409);
or UO_949 (O_949,N_19074,N_19519);
nor UO_950 (O_950,N_19428,N_19815);
nor UO_951 (O_951,N_19788,N_19755);
and UO_952 (O_952,N_19942,N_19650);
and UO_953 (O_953,N_19479,N_19262);
xor UO_954 (O_954,N_19551,N_19435);
nand UO_955 (O_955,N_19653,N_19222);
or UO_956 (O_956,N_19871,N_19890);
and UO_957 (O_957,N_19702,N_19312);
or UO_958 (O_958,N_19736,N_19443);
xnor UO_959 (O_959,N_19540,N_19640);
nor UO_960 (O_960,N_19137,N_19357);
or UO_961 (O_961,N_19438,N_19110);
nand UO_962 (O_962,N_19797,N_19196);
xnor UO_963 (O_963,N_19257,N_19670);
xor UO_964 (O_964,N_19149,N_19045);
nand UO_965 (O_965,N_19365,N_19164);
nand UO_966 (O_966,N_19455,N_19894);
xnor UO_967 (O_967,N_19166,N_19866);
nor UO_968 (O_968,N_19104,N_19129);
and UO_969 (O_969,N_19413,N_19969);
nor UO_970 (O_970,N_19550,N_19891);
nor UO_971 (O_971,N_19597,N_19431);
or UO_972 (O_972,N_19777,N_19441);
and UO_973 (O_973,N_19425,N_19115);
or UO_974 (O_974,N_19398,N_19412);
and UO_975 (O_975,N_19374,N_19604);
nand UO_976 (O_976,N_19973,N_19776);
or UO_977 (O_977,N_19578,N_19072);
nand UO_978 (O_978,N_19483,N_19306);
or UO_979 (O_979,N_19678,N_19397);
nor UO_980 (O_980,N_19514,N_19336);
nand UO_981 (O_981,N_19380,N_19137);
nor UO_982 (O_982,N_19646,N_19228);
nor UO_983 (O_983,N_19584,N_19060);
or UO_984 (O_984,N_19451,N_19794);
or UO_985 (O_985,N_19220,N_19212);
nor UO_986 (O_986,N_19646,N_19384);
nor UO_987 (O_987,N_19591,N_19647);
nand UO_988 (O_988,N_19958,N_19818);
or UO_989 (O_989,N_19136,N_19259);
nand UO_990 (O_990,N_19079,N_19934);
and UO_991 (O_991,N_19293,N_19524);
xor UO_992 (O_992,N_19103,N_19626);
xnor UO_993 (O_993,N_19878,N_19723);
or UO_994 (O_994,N_19099,N_19532);
and UO_995 (O_995,N_19610,N_19049);
nand UO_996 (O_996,N_19182,N_19660);
nand UO_997 (O_997,N_19499,N_19026);
nor UO_998 (O_998,N_19547,N_19318);
and UO_999 (O_999,N_19100,N_19234);
or UO_1000 (O_1000,N_19474,N_19882);
nor UO_1001 (O_1001,N_19752,N_19529);
or UO_1002 (O_1002,N_19921,N_19706);
nand UO_1003 (O_1003,N_19449,N_19117);
or UO_1004 (O_1004,N_19814,N_19063);
or UO_1005 (O_1005,N_19593,N_19981);
and UO_1006 (O_1006,N_19700,N_19648);
nor UO_1007 (O_1007,N_19322,N_19537);
nor UO_1008 (O_1008,N_19579,N_19910);
or UO_1009 (O_1009,N_19730,N_19009);
and UO_1010 (O_1010,N_19245,N_19194);
and UO_1011 (O_1011,N_19426,N_19907);
xnor UO_1012 (O_1012,N_19315,N_19775);
nand UO_1013 (O_1013,N_19689,N_19370);
or UO_1014 (O_1014,N_19784,N_19944);
nor UO_1015 (O_1015,N_19514,N_19840);
nor UO_1016 (O_1016,N_19691,N_19884);
or UO_1017 (O_1017,N_19563,N_19938);
xnor UO_1018 (O_1018,N_19878,N_19017);
or UO_1019 (O_1019,N_19577,N_19959);
nor UO_1020 (O_1020,N_19103,N_19306);
or UO_1021 (O_1021,N_19514,N_19846);
nor UO_1022 (O_1022,N_19523,N_19286);
nor UO_1023 (O_1023,N_19953,N_19305);
and UO_1024 (O_1024,N_19412,N_19324);
or UO_1025 (O_1025,N_19877,N_19820);
xor UO_1026 (O_1026,N_19769,N_19726);
and UO_1027 (O_1027,N_19592,N_19482);
nor UO_1028 (O_1028,N_19280,N_19122);
nor UO_1029 (O_1029,N_19359,N_19312);
xor UO_1030 (O_1030,N_19195,N_19621);
and UO_1031 (O_1031,N_19374,N_19751);
nor UO_1032 (O_1032,N_19004,N_19846);
nor UO_1033 (O_1033,N_19522,N_19695);
xor UO_1034 (O_1034,N_19818,N_19211);
xnor UO_1035 (O_1035,N_19371,N_19010);
or UO_1036 (O_1036,N_19436,N_19845);
nand UO_1037 (O_1037,N_19026,N_19989);
or UO_1038 (O_1038,N_19649,N_19736);
xor UO_1039 (O_1039,N_19885,N_19946);
nor UO_1040 (O_1040,N_19969,N_19043);
xor UO_1041 (O_1041,N_19938,N_19307);
xnor UO_1042 (O_1042,N_19227,N_19536);
xnor UO_1043 (O_1043,N_19624,N_19362);
nand UO_1044 (O_1044,N_19904,N_19637);
nor UO_1045 (O_1045,N_19496,N_19118);
nor UO_1046 (O_1046,N_19021,N_19968);
nand UO_1047 (O_1047,N_19735,N_19444);
nand UO_1048 (O_1048,N_19825,N_19933);
or UO_1049 (O_1049,N_19173,N_19358);
nor UO_1050 (O_1050,N_19633,N_19073);
nand UO_1051 (O_1051,N_19385,N_19309);
and UO_1052 (O_1052,N_19775,N_19721);
or UO_1053 (O_1053,N_19752,N_19810);
nor UO_1054 (O_1054,N_19101,N_19534);
nor UO_1055 (O_1055,N_19534,N_19637);
or UO_1056 (O_1056,N_19005,N_19551);
nand UO_1057 (O_1057,N_19651,N_19131);
xor UO_1058 (O_1058,N_19679,N_19796);
xnor UO_1059 (O_1059,N_19732,N_19292);
nor UO_1060 (O_1060,N_19091,N_19540);
and UO_1061 (O_1061,N_19651,N_19115);
or UO_1062 (O_1062,N_19661,N_19032);
xnor UO_1063 (O_1063,N_19629,N_19840);
and UO_1064 (O_1064,N_19217,N_19171);
or UO_1065 (O_1065,N_19523,N_19881);
or UO_1066 (O_1066,N_19927,N_19995);
nand UO_1067 (O_1067,N_19523,N_19876);
nor UO_1068 (O_1068,N_19620,N_19589);
and UO_1069 (O_1069,N_19208,N_19650);
nor UO_1070 (O_1070,N_19091,N_19883);
nor UO_1071 (O_1071,N_19068,N_19137);
nor UO_1072 (O_1072,N_19589,N_19972);
xor UO_1073 (O_1073,N_19055,N_19101);
nand UO_1074 (O_1074,N_19999,N_19013);
nor UO_1075 (O_1075,N_19989,N_19695);
and UO_1076 (O_1076,N_19709,N_19590);
or UO_1077 (O_1077,N_19671,N_19288);
nand UO_1078 (O_1078,N_19617,N_19691);
or UO_1079 (O_1079,N_19988,N_19335);
nand UO_1080 (O_1080,N_19119,N_19786);
and UO_1081 (O_1081,N_19852,N_19557);
and UO_1082 (O_1082,N_19204,N_19154);
nand UO_1083 (O_1083,N_19402,N_19815);
nand UO_1084 (O_1084,N_19352,N_19489);
or UO_1085 (O_1085,N_19099,N_19718);
xor UO_1086 (O_1086,N_19885,N_19993);
and UO_1087 (O_1087,N_19315,N_19931);
nor UO_1088 (O_1088,N_19810,N_19926);
and UO_1089 (O_1089,N_19609,N_19189);
nor UO_1090 (O_1090,N_19000,N_19078);
xnor UO_1091 (O_1091,N_19688,N_19176);
nand UO_1092 (O_1092,N_19165,N_19293);
nand UO_1093 (O_1093,N_19339,N_19633);
or UO_1094 (O_1094,N_19761,N_19145);
and UO_1095 (O_1095,N_19583,N_19023);
or UO_1096 (O_1096,N_19037,N_19601);
nor UO_1097 (O_1097,N_19493,N_19672);
and UO_1098 (O_1098,N_19031,N_19177);
nand UO_1099 (O_1099,N_19255,N_19482);
nor UO_1100 (O_1100,N_19109,N_19879);
or UO_1101 (O_1101,N_19648,N_19238);
nor UO_1102 (O_1102,N_19354,N_19941);
or UO_1103 (O_1103,N_19850,N_19023);
xnor UO_1104 (O_1104,N_19130,N_19482);
or UO_1105 (O_1105,N_19497,N_19060);
nand UO_1106 (O_1106,N_19537,N_19975);
or UO_1107 (O_1107,N_19278,N_19619);
nand UO_1108 (O_1108,N_19338,N_19573);
and UO_1109 (O_1109,N_19503,N_19346);
or UO_1110 (O_1110,N_19871,N_19731);
or UO_1111 (O_1111,N_19859,N_19158);
or UO_1112 (O_1112,N_19298,N_19412);
nand UO_1113 (O_1113,N_19827,N_19956);
xnor UO_1114 (O_1114,N_19862,N_19246);
nand UO_1115 (O_1115,N_19407,N_19644);
or UO_1116 (O_1116,N_19275,N_19019);
or UO_1117 (O_1117,N_19702,N_19923);
nand UO_1118 (O_1118,N_19913,N_19493);
and UO_1119 (O_1119,N_19221,N_19894);
or UO_1120 (O_1120,N_19021,N_19709);
or UO_1121 (O_1121,N_19607,N_19504);
and UO_1122 (O_1122,N_19410,N_19058);
or UO_1123 (O_1123,N_19153,N_19064);
nand UO_1124 (O_1124,N_19982,N_19386);
xnor UO_1125 (O_1125,N_19967,N_19770);
and UO_1126 (O_1126,N_19382,N_19490);
and UO_1127 (O_1127,N_19418,N_19970);
xnor UO_1128 (O_1128,N_19253,N_19897);
or UO_1129 (O_1129,N_19371,N_19842);
and UO_1130 (O_1130,N_19282,N_19059);
and UO_1131 (O_1131,N_19889,N_19485);
or UO_1132 (O_1132,N_19056,N_19645);
nand UO_1133 (O_1133,N_19370,N_19082);
or UO_1134 (O_1134,N_19646,N_19828);
nor UO_1135 (O_1135,N_19034,N_19887);
and UO_1136 (O_1136,N_19801,N_19284);
or UO_1137 (O_1137,N_19317,N_19845);
nor UO_1138 (O_1138,N_19059,N_19810);
nand UO_1139 (O_1139,N_19396,N_19138);
nand UO_1140 (O_1140,N_19320,N_19179);
and UO_1141 (O_1141,N_19931,N_19939);
and UO_1142 (O_1142,N_19523,N_19128);
nor UO_1143 (O_1143,N_19931,N_19542);
nor UO_1144 (O_1144,N_19113,N_19156);
or UO_1145 (O_1145,N_19037,N_19460);
xor UO_1146 (O_1146,N_19687,N_19745);
nand UO_1147 (O_1147,N_19602,N_19130);
and UO_1148 (O_1148,N_19170,N_19358);
and UO_1149 (O_1149,N_19132,N_19802);
nor UO_1150 (O_1150,N_19110,N_19582);
xor UO_1151 (O_1151,N_19690,N_19344);
and UO_1152 (O_1152,N_19130,N_19274);
nand UO_1153 (O_1153,N_19345,N_19784);
or UO_1154 (O_1154,N_19989,N_19448);
nor UO_1155 (O_1155,N_19953,N_19655);
or UO_1156 (O_1156,N_19427,N_19568);
xor UO_1157 (O_1157,N_19786,N_19647);
nor UO_1158 (O_1158,N_19598,N_19117);
nand UO_1159 (O_1159,N_19577,N_19923);
nand UO_1160 (O_1160,N_19826,N_19629);
nor UO_1161 (O_1161,N_19094,N_19533);
nand UO_1162 (O_1162,N_19916,N_19728);
nor UO_1163 (O_1163,N_19546,N_19921);
nand UO_1164 (O_1164,N_19398,N_19181);
xor UO_1165 (O_1165,N_19349,N_19011);
and UO_1166 (O_1166,N_19710,N_19596);
or UO_1167 (O_1167,N_19531,N_19940);
or UO_1168 (O_1168,N_19848,N_19700);
nand UO_1169 (O_1169,N_19086,N_19527);
nand UO_1170 (O_1170,N_19079,N_19649);
xor UO_1171 (O_1171,N_19919,N_19536);
nor UO_1172 (O_1172,N_19878,N_19644);
xnor UO_1173 (O_1173,N_19928,N_19273);
nand UO_1174 (O_1174,N_19469,N_19403);
nor UO_1175 (O_1175,N_19112,N_19348);
nand UO_1176 (O_1176,N_19555,N_19326);
xor UO_1177 (O_1177,N_19233,N_19282);
and UO_1178 (O_1178,N_19482,N_19881);
nor UO_1179 (O_1179,N_19558,N_19160);
and UO_1180 (O_1180,N_19013,N_19863);
xnor UO_1181 (O_1181,N_19969,N_19626);
or UO_1182 (O_1182,N_19436,N_19191);
nand UO_1183 (O_1183,N_19371,N_19485);
nor UO_1184 (O_1184,N_19848,N_19354);
and UO_1185 (O_1185,N_19997,N_19022);
nor UO_1186 (O_1186,N_19179,N_19956);
xnor UO_1187 (O_1187,N_19300,N_19479);
nor UO_1188 (O_1188,N_19198,N_19936);
or UO_1189 (O_1189,N_19602,N_19458);
nand UO_1190 (O_1190,N_19203,N_19729);
nor UO_1191 (O_1191,N_19630,N_19134);
and UO_1192 (O_1192,N_19408,N_19535);
nand UO_1193 (O_1193,N_19146,N_19702);
nand UO_1194 (O_1194,N_19072,N_19049);
xnor UO_1195 (O_1195,N_19342,N_19250);
nor UO_1196 (O_1196,N_19647,N_19251);
or UO_1197 (O_1197,N_19011,N_19265);
nand UO_1198 (O_1198,N_19865,N_19148);
xnor UO_1199 (O_1199,N_19742,N_19203);
and UO_1200 (O_1200,N_19745,N_19707);
nor UO_1201 (O_1201,N_19628,N_19996);
xor UO_1202 (O_1202,N_19538,N_19015);
xnor UO_1203 (O_1203,N_19538,N_19201);
and UO_1204 (O_1204,N_19757,N_19456);
or UO_1205 (O_1205,N_19144,N_19092);
nand UO_1206 (O_1206,N_19868,N_19056);
nand UO_1207 (O_1207,N_19217,N_19279);
or UO_1208 (O_1208,N_19247,N_19222);
and UO_1209 (O_1209,N_19995,N_19126);
xor UO_1210 (O_1210,N_19549,N_19321);
nand UO_1211 (O_1211,N_19972,N_19379);
xor UO_1212 (O_1212,N_19069,N_19672);
xor UO_1213 (O_1213,N_19253,N_19611);
or UO_1214 (O_1214,N_19172,N_19848);
or UO_1215 (O_1215,N_19209,N_19136);
or UO_1216 (O_1216,N_19659,N_19108);
or UO_1217 (O_1217,N_19434,N_19019);
xor UO_1218 (O_1218,N_19551,N_19209);
and UO_1219 (O_1219,N_19353,N_19644);
xor UO_1220 (O_1220,N_19550,N_19063);
nor UO_1221 (O_1221,N_19779,N_19041);
nor UO_1222 (O_1222,N_19080,N_19170);
nor UO_1223 (O_1223,N_19650,N_19205);
xnor UO_1224 (O_1224,N_19258,N_19939);
and UO_1225 (O_1225,N_19180,N_19797);
nand UO_1226 (O_1226,N_19058,N_19390);
xnor UO_1227 (O_1227,N_19822,N_19212);
nor UO_1228 (O_1228,N_19148,N_19891);
xnor UO_1229 (O_1229,N_19729,N_19718);
and UO_1230 (O_1230,N_19634,N_19874);
nor UO_1231 (O_1231,N_19117,N_19028);
xnor UO_1232 (O_1232,N_19558,N_19993);
or UO_1233 (O_1233,N_19614,N_19528);
or UO_1234 (O_1234,N_19955,N_19249);
xnor UO_1235 (O_1235,N_19427,N_19209);
xor UO_1236 (O_1236,N_19122,N_19253);
xor UO_1237 (O_1237,N_19331,N_19333);
and UO_1238 (O_1238,N_19436,N_19234);
nor UO_1239 (O_1239,N_19017,N_19235);
nand UO_1240 (O_1240,N_19204,N_19662);
and UO_1241 (O_1241,N_19387,N_19024);
or UO_1242 (O_1242,N_19368,N_19489);
nand UO_1243 (O_1243,N_19908,N_19806);
nand UO_1244 (O_1244,N_19069,N_19180);
nand UO_1245 (O_1245,N_19983,N_19494);
xor UO_1246 (O_1246,N_19947,N_19669);
and UO_1247 (O_1247,N_19696,N_19143);
xnor UO_1248 (O_1248,N_19731,N_19867);
nand UO_1249 (O_1249,N_19406,N_19999);
and UO_1250 (O_1250,N_19161,N_19624);
nor UO_1251 (O_1251,N_19060,N_19344);
and UO_1252 (O_1252,N_19655,N_19479);
nor UO_1253 (O_1253,N_19363,N_19189);
and UO_1254 (O_1254,N_19640,N_19260);
xor UO_1255 (O_1255,N_19850,N_19362);
or UO_1256 (O_1256,N_19315,N_19718);
or UO_1257 (O_1257,N_19435,N_19726);
nor UO_1258 (O_1258,N_19043,N_19100);
xor UO_1259 (O_1259,N_19655,N_19456);
nor UO_1260 (O_1260,N_19035,N_19197);
nor UO_1261 (O_1261,N_19527,N_19839);
or UO_1262 (O_1262,N_19250,N_19025);
nor UO_1263 (O_1263,N_19944,N_19227);
or UO_1264 (O_1264,N_19744,N_19335);
nand UO_1265 (O_1265,N_19955,N_19929);
nand UO_1266 (O_1266,N_19937,N_19217);
nor UO_1267 (O_1267,N_19321,N_19510);
nand UO_1268 (O_1268,N_19830,N_19724);
or UO_1269 (O_1269,N_19826,N_19140);
and UO_1270 (O_1270,N_19774,N_19547);
or UO_1271 (O_1271,N_19762,N_19637);
and UO_1272 (O_1272,N_19369,N_19501);
xnor UO_1273 (O_1273,N_19680,N_19429);
nand UO_1274 (O_1274,N_19270,N_19365);
and UO_1275 (O_1275,N_19078,N_19796);
nand UO_1276 (O_1276,N_19498,N_19734);
or UO_1277 (O_1277,N_19707,N_19278);
xor UO_1278 (O_1278,N_19137,N_19696);
or UO_1279 (O_1279,N_19714,N_19372);
xor UO_1280 (O_1280,N_19587,N_19057);
nand UO_1281 (O_1281,N_19325,N_19397);
and UO_1282 (O_1282,N_19623,N_19145);
nand UO_1283 (O_1283,N_19722,N_19268);
and UO_1284 (O_1284,N_19768,N_19955);
xor UO_1285 (O_1285,N_19207,N_19182);
nor UO_1286 (O_1286,N_19701,N_19333);
nand UO_1287 (O_1287,N_19730,N_19857);
nand UO_1288 (O_1288,N_19228,N_19950);
and UO_1289 (O_1289,N_19836,N_19424);
xor UO_1290 (O_1290,N_19028,N_19761);
nand UO_1291 (O_1291,N_19782,N_19707);
or UO_1292 (O_1292,N_19587,N_19908);
and UO_1293 (O_1293,N_19740,N_19679);
or UO_1294 (O_1294,N_19373,N_19892);
or UO_1295 (O_1295,N_19199,N_19814);
and UO_1296 (O_1296,N_19655,N_19873);
or UO_1297 (O_1297,N_19579,N_19022);
and UO_1298 (O_1298,N_19209,N_19203);
or UO_1299 (O_1299,N_19621,N_19558);
nor UO_1300 (O_1300,N_19450,N_19506);
and UO_1301 (O_1301,N_19639,N_19283);
and UO_1302 (O_1302,N_19016,N_19826);
nand UO_1303 (O_1303,N_19540,N_19088);
nand UO_1304 (O_1304,N_19107,N_19975);
nor UO_1305 (O_1305,N_19467,N_19029);
and UO_1306 (O_1306,N_19549,N_19053);
xor UO_1307 (O_1307,N_19978,N_19699);
xor UO_1308 (O_1308,N_19416,N_19308);
and UO_1309 (O_1309,N_19265,N_19859);
and UO_1310 (O_1310,N_19765,N_19075);
nor UO_1311 (O_1311,N_19748,N_19797);
nand UO_1312 (O_1312,N_19373,N_19554);
or UO_1313 (O_1313,N_19698,N_19695);
and UO_1314 (O_1314,N_19548,N_19690);
or UO_1315 (O_1315,N_19326,N_19334);
xor UO_1316 (O_1316,N_19773,N_19291);
xor UO_1317 (O_1317,N_19585,N_19378);
xnor UO_1318 (O_1318,N_19751,N_19027);
nor UO_1319 (O_1319,N_19662,N_19335);
and UO_1320 (O_1320,N_19088,N_19274);
nor UO_1321 (O_1321,N_19491,N_19113);
nand UO_1322 (O_1322,N_19002,N_19119);
nor UO_1323 (O_1323,N_19440,N_19874);
or UO_1324 (O_1324,N_19731,N_19248);
and UO_1325 (O_1325,N_19887,N_19911);
nand UO_1326 (O_1326,N_19405,N_19121);
nand UO_1327 (O_1327,N_19845,N_19367);
nand UO_1328 (O_1328,N_19333,N_19088);
nand UO_1329 (O_1329,N_19354,N_19679);
xor UO_1330 (O_1330,N_19617,N_19536);
nand UO_1331 (O_1331,N_19006,N_19781);
or UO_1332 (O_1332,N_19344,N_19785);
xor UO_1333 (O_1333,N_19918,N_19835);
and UO_1334 (O_1334,N_19675,N_19716);
and UO_1335 (O_1335,N_19511,N_19534);
and UO_1336 (O_1336,N_19170,N_19418);
xnor UO_1337 (O_1337,N_19662,N_19801);
or UO_1338 (O_1338,N_19830,N_19455);
nand UO_1339 (O_1339,N_19274,N_19697);
nor UO_1340 (O_1340,N_19648,N_19411);
nor UO_1341 (O_1341,N_19913,N_19384);
and UO_1342 (O_1342,N_19964,N_19624);
nand UO_1343 (O_1343,N_19521,N_19617);
xnor UO_1344 (O_1344,N_19251,N_19619);
nor UO_1345 (O_1345,N_19394,N_19666);
and UO_1346 (O_1346,N_19169,N_19985);
nor UO_1347 (O_1347,N_19548,N_19475);
xor UO_1348 (O_1348,N_19986,N_19373);
nand UO_1349 (O_1349,N_19813,N_19846);
nor UO_1350 (O_1350,N_19281,N_19047);
nand UO_1351 (O_1351,N_19922,N_19218);
nor UO_1352 (O_1352,N_19323,N_19942);
nand UO_1353 (O_1353,N_19074,N_19923);
and UO_1354 (O_1354,N_19439,N_19075);
nor UO_1355 (O_1355,N_19779,N_19616);
or UO_1356 (O_1356,N_19257,N_19669);
or UO_1357 (O_1357,N_19443,N_19890);
xnor UO_1358 (O_1358,N_19135,N_19836);
nor UO_1359 (O_1359,N_19573,N_19413);
and UO_1360 (O_1360,N_19660,N_19140);
nor UO_1361 (O_1361,N_19000,N_19039);
nand UO_1362 (O_1362,N_19960,N_19334);
nand UO_1363 (O_1363,N_19620,N_19123);
xnor UO_1364 (O_1364,N_19178,N_19829);
nor UO_1365 (O_1365,N_19829,N_19826);
xor UO_1366 (O_1366,N_19603,N_19143);
or UO_1367 (O_1367,N_19456,N_19646);
or UO_1368 (O_1368,N_19363,N_19192);
nand UO_1369 (O_1369,N_19497,N_19587);
or UO_1370 (O_1370,N_19641,N_19470);
nand UO_1371 (O_1371,N_19191,N_19445);
and UO_1372 (O_1372,N_19679,N_19144);
nand UO_1373 (O_1373,N_19250,N_19803);
nor UO_1374 (O_1374,N_19598,N_19451);
nor UO_1375 (O_1375,N_19789,N_19276);
nor UO_1376 (O_1376,N_19707,N_19873);
and UO_1377 (O_1377,N_19997,N_19302);
and UO_1378 (O_1378,N_19601,N_19281);
or UO_1379 (O_1379,N_19672,N_19997);
nand UO_1380 (O_1380,N_19008,N_19706);
and UO_1381 (O_1381,N_19678,N_19387);
or UO_1382 (O_1382,N_19651,N_19141);
nor UO_1383 (O_1383,N_19231,N_19114);
nor UO_1384 (O_1384,N_19299,N_19216);
xor UO_1385 (O_1385,N_19935,N_19449);
or UO_1386 (O_1386,N_19509,N_19719);
and UO_1387 (O_1387,N_19418,N_19033);
nor UO_1388 (O_1388,N_19359,N_19172);
nor UO_1389 (O_1389,N_19127,N_19877);
nand UO_1390 (O_1390,N_19738,N_19762);
and UO_1391 (O_1391,N_19295,N_19716);
nand UO_1392 (O_1392,N_19198,N_19027);
xor UO_1393 (O_1393,N_19285,N_19535);
or UO_1394 (O_1394,N_19636,N_19883);
xor UO_1395 (O_1395,N_19292,N_19583);
nand UO_1396 (O_1396,N_19106,N_19998);
nand UO_1397 (O_1397,N_19603,N_19960);
xor UO_1398 (O_1398,N_19570,N_19798);
or UO_1399 (O_1399,N_19040,N_19130);
or UO_1400 (O_1400,N_19597,N_19330);
nand UO_1401 (O_1401,N_19830,N_19560);
nor UO_1402 (O_1402,N_19597,N_19518);
nor UO_1403 (O_1403,N_19270,N_19545);
nand UO_1404 (O_1404,N_19609,N_19084);
and UO_1405 (O_1405,N_19759,N_19218);
or UO_1406 (O_1406,N_19113,N_19210);
and UO_1407 (O_1407,N_19174,N_19031);
xor UO_1408 (O_1408,N_19112,N_19194);
and UO_1409 (O_1409,N_19102,N_19104);
nand UO_1410 (O_1410,N_19031,N_19855);
nor UO_1411 (O_1411,N_19563,N_19454);
nor UO_1412 (O_1412,N_19458,N_19036);
xor UO_1413 (O_1413,N_19622,N_19403);
or UO_1414 (O_1414,N_19363,N_19184);
and UO_1415 (O_1415,N_19262,N_19481);
or UO_1416 (O_1416,N_19332,N_19153);
nor UO_1417 (O_1417,N_19776,N_19362);
nor UO_1418 (O_1418,N_19285,N_19590);
and UO_1419 (O_1419,N_19904,N_19176);
or UO_1420 (O_1420,N_19877,N_19742);
xnor UO_1421 (O_1421,N_19252,N_19015);
xor UO_1422 (O_1422,N_19630,N_19551);
xnor UO_1423 (O_1423,N_19118,N_19385);
or UO_1424 (O_1424,N_19170,N_19352);
xor UO_1425 (O_1425,N_19963,N_19007);
and UO_1426 (O_1426,N_19745,N_19578);
xor UO_1427 (O_1427,N_19598,N_19222);
or UO_1428 (O_1428,N_19743,N_19550);
xnor UO_1429 (O_1429,N_19798,N_19146);
nand UO_1430 (O_1430,N_19291,N_19735);
or UO_1431 (O_1431,N_19785,N_19036);
and UO_1432 (O_1432,N_19661,N_19435);
and UO_1433 (O_1433,N_19992,N_19541);
and UO_1434 (O_1434,N_19678,N_19706);
or UO_1435 (O_1435,N_19662,N_19068);
and UO_1436 (O_1436,N_19607,N_19805);
or UO_1437 (O_1437,N_19166,N_19091);
xnor UO_1438 (O_1438,N_19911,N_19775);
nor UO_1439 (O_1439,N_19760,N_19181);
nor UO_1440 (O_1440,N_19029,N_19261);
xnor UO_1441 (O_1441,N_19434,N_19965);
nor UO_1442 (O_1442,N_19620,N_19593);
nor UO_1443 (O_1443,N_19331,N_19072);
or UO_1444 (O_1444,N_19811,N_19703);
xnor UO_1445 (O_1445,N_19026,N_19909);
or UO_1446 (O_1446,N_19535,N_19930);
nor UO_1447 (O_1447,N_19198,N_19806);
nand UO_1448 (O_1448,N_19098,N_19529);
xor UO_1449 (O_1449,N_19744,N_19682);
nor UO_1450 (O_1450,N_19408,N_19868);
nand UO_1451 (O_1451,N_19927,N_19793);
nor UO_1452 (O_1452,N_19772,N_19915);
nand UO_1453 (O_1453,N_19614,N_19134);
and UO_1454 (O_1454,N_19729,N_19211);
or UO_1455 (O_1455,N_19358,N_19656);
nand UO_1456 (O_1456,N_19741,N_19425);
nand UO_1457 (O_1457,N_19754,N_19000);
or UO_1458 (O_1458,N_19848,N_19027);
and UO_1459 (O_1459,N_19393,N_19227);
nor UO_1460 (O_1460,N_19337,N_19125);
nor UO_1461 (O_1461,N_19251,N_19826);
nand UO_1462 (O_1462,N_19356,N_19760);
nor UO_1463 (O_1463,N_19076,N_19051);
nand UO_1464 (O_1464,N_19393,N_19938);
and UO_1465 (O_1465,N_19140,N_19152);
xnor UO_1466 (O_1466,N_19066,N_19120);
and UO_1467 (O_1467,N_19126,N_19675);
or UO_1468 (O_1468,N_19694,N_19239);
or UO_1469 (O_1469,N_19421,N_19053);
and UO_1470 (O_1470,N_19163,N_19147);
nor UO_1471 (O_1471,N_19725,N_19153);
nor UO_1472 (O_1472,N_19135,N_19517);
or UO_1473 (O_1473,N_19204,N_19605);
nor UO_1474 (O_1474,N_19682,N_19851);
nand UO_1475 (O_1475,N_19016,N_19252);
nand UO_1476 (O_1476,N_19775,N_19716);
and UO_1477 (O_1477,N_19907,N_19343);
and UO_1478 (O_1478,N_19260,N_19621);
or UO_1479 (O_1479,N_19712,N_19706);
or UO_1480 (O_1480,N_19128,N_19632);
or UO_1481 (O_1481,N_19037,N_19456);
and UO_1482 (O_1482,N_19179,N_19193);
nor UO_1483 (O_1483,N_19772,N_19794);
xor UO_1484 (O_1484,N_19102,N_19251);
or UO_1485 (O_1485,N_19553,N_19731);
nor UO_1486 (O_1486,N_19916,N_19578);
and UO_1487 (O_1487,N_19416,N_19352);
or UO_1488 (O_1488,N_19253,N_19350);
nor UO_1489 (O_1489,N_19299,N_19938);
and UO_1490 (O_1490,N_19439,N_19988);
nor UO_1491 (O_1491,N_19820,N_19383);
xor UO_1492 (O_1492,N_19411,N_19044);
nor UO_1493 (O_1493,N_19824,N_19169);
xor UO_1494 (O_1494,N_19102,N_19157);
xor UO_1495 (O_1495,N_19252,N_19526);
or UO_1496 (O_1496,N_19589,N_19244);
and UO_1497 (O_1497,N_19167,N_19122);
and UO_1498 (O_1498,N_19905,N_19861);
nand UO_1499 (O_1499,N_19417,N_19390);
or UO_1500 (O_1500,N_19395,N_19436);
or UO_1501 (O_1501,N_19961,N_19887);
and UO_1502 (O_1502,N_19650,N_19943);
or UO_1503 (O_1503,N_19512,N_19810);
nand UO_1504 (O_1504,N_19131,N_19378);
nor UO_1505 (O_1505,N_19725,N_19868);
or UO_1506 (O_1506,N_19485,N_19397);
nor UO_1507 (O_1507,N_19891,N_19166);
nor UO_1508 (O_1508,N_19217,N_19748);
xnor UO_1509 (O_1509,N_19597,N_19844);
or UO_1510 (O_1510,N_19148,N_19041);
nand UO_1511 (O_1511,N_19335,N_19952);
or UO_1512 (O_1512,N_19511,N_19552);
nor UO_1513 (O_1513,N_19786,N_19049);
nor UO_1514 (O_1514,N_19808,N_19215);
and UO_1515 (O_1515,N_19821,N_19762);
or UO_1516 (O_1516,N_19989,N_19821);
nor UO_1517 (O_1517,N_19428,N_19045);
nand UO_1518 (O_1518,N_19479,N_19856);
or UO_1519 (O_1519,N_19747,N_19148);
nand UO_1520 (O_1520,N_19887,N_19980);
nand UO_1521 (O_1521,N_19648,N_19487);
xor UO_1522 (O_1522,N_19474,N_19245);
nor UO_1523 (O_1523,N_19836,N_19402);
nand UO_1524 (O_1524,N_19230,N_19599);
and UO_1525 (O_1525,N_19898,N_19459);
xnor UO_1526 (O_1526,N_19263,N_19730);
and UO_1527 (O_1527,N_19398,N_19027);
and UO_1528 (O_1528,N_19698,N_19071);
xor UO_1529 (O_1529,N_19080,N_19252);
nor UO_1530 (O_1530,N_19756,N_19895);
and UO_1531 (O_1531,N_19221,N_19826);
nand UO_1532 (O_1532,N_19404,N_19735);
and UO_1533 (O_1533,N_19446,N_19497);
and UO_1534 (O_1534,N_19438,N_19268);
and UO_1535 (O_1535,N_19399,N_19113);
xor UO_1536 (O_1536,N_19921,N_19832);
nand UO_1537 (O_1537,N_19533,N_19111);
nor UO_1538 (O_1538,N_19126,N_19154);
nor UO_1539 (O_1539,N_19277,N_19724);
xnor UO_1540 (O_1540,N_19081,N_19433);
and UO_1541 (O_1541,N_19498,N_19021);
xor UO_1542 (O_1542,N_19522,N_19176);
xor UO_1543 (O_1543,N_19296,N_19613);
nand UO_1544 (O_1544,N_19271,N_19754);
xnor UO_1545 (O_1545,N_19809,N_19311);
nand UO_1546 (O_1546,N_19718,N_19356);
and UO_1547 (O_1547,N_19031,N_19410);
and UO_1548 (O_1548,N_19809,N_19373);
nor UO_1549 (O_1549,N_19462,N_19323);
or UO_1550 (O_1550,N_19283,N_19036);
and UO_1551 (O_1551,N_19145,N_19357);
xor UO_1552 (O_1552,N_19038,N_19195);
or UO_1553 (O_1553,N_19692,N_19133);
and UO_1554 (O_1554,N_19550,N_19978);
nand UO_1555 (O_1555,N_19127,N_19171);
xnor UO_1556 (O_1556,N_19330,N_19039);
xor UO_1557 (O_1557,N_19748,N_19871);
and UO_1558 (O_1558,N_19354,N_19603);
and UO_1559 (O_1559,N_19890,N_19459);
nand UO_1560 (O_1560,N_19917,N_19536);
xnor UO_1561 (O_1561,N_19215,N_19574);
xor UO_1562 (O_1562,N_19555,N_19573);
xnor UO_1563 (O_1563,N_19568,N_19143);
or UO_1564 (O_1564,N_19042,N_19077);
nor UO_1565 (O_1565,N_19202,N_19318);
and UO_1566 (O_1566,N_19345,N_19602);
and UO_1567 (O_1567,N_19487,N_19016);
xnor UO_1568 (O_1568,N_19034,N_19176);
or UO_1569 (O_1569,N_19423,N_19089);
and UO_1570 (O_1570,N_19817,N_19480);
nor UO_1571 (O_1571,N_19245,N_19280);
nand UO_1572 (O_1572,N_19158,N_19066);
and UO_1573 (O_1573,N_19762,N_19846);
nor UO_1574 (O_1574,N_19910,N_19027);
nor UO_1575 (O_1575,N_19353,N_19335);
nor UO_1576 (O_1576,N_19984,N_19332);
nand UO_1577 (O_1577,N_19711,N_19397);
or UO_1578 (O_1578,N_19066,N_19516);
nor UO_1579 (O_1579,N_19545,N_19299);
nor UO_1580 (O_1580,N_19781,N_19751);
or UO_1581 (O_1581,N_19846,N_19489);
and UO_1582 (O_1582,N_19273,N_19670);
xor UO_1583 (O_1583,N_19151,N_19150);
nor UO_1584 (O_1584,N_19559,N_19845);
nor UO_1585 (O_1585,N_19304,N_19409);
and UO_1586 (O_1586,N_19381,N_19358);
nand UO_1587 (O_1587,N_19550,N_19572);
xor UO_1588 (O_1588,N_19964,N_19567);
xnor UO_1589 (O_1589,N_19746,N_19587);
nor UO_1590 (O_1590,N_19548,N_19534);
xnor UO_1591 (O_1591,N_19806,N_19878);
xnor UO_1592 (O_1592,N_19395,N_19080);
nor UO_1593 (O_1593,N_19212,N_19813);
and UO_1594 (O_1594,N_19917,N_19427);
nor UO_1595 (O_1595,N_19213,N_19765);
or UO_1596 (O_1596,N_19475,N_19794);
xnor UO_1597 (O_1597,N_19443,N_19789);
nand UO_1598 (O_1598,N_19092,N_19254);
or UO_1599 (O_1599,N_19080,N_19494);
xnor UO_1600 (O_1600,N_19052,N_19078);
nor UO_1601 (O_1601,N_19733,N_19570);
nand UO_1602 (O_1602,N_19136,N_19951);
and UO_1603 (O_1603,N_19550,N_19952);
xnor UO_1604 (O_1604,N_19205,N_19360);
xnor UO_1605 (O_1605,N_19315,N_19889);
and UO_1606 (O_1606,N_19704,N_19465);
or UO_1607 (O_1607,N_19687,N_19210);
nor UO_1608 (O_1608,N_19764,N_19239);
nor UO_1609 (O_1609,N_19951,N_19255);
nand UO_1610 (O_1610,N_19097,N_19150);
and UO_1611 (O_1611,N_19032,N_19128);
xnor UO_1612 (O_1612,N_19680,N_19868);
nor UO_1613 (O_1613,N_19455,N_19501);
and UO_1614 (O_1614,N_19412,N_19480);
nor UO_1615 (O_1615,N_19443,N_19416);
nand UO_1616 (O_1616,N_19199,N_19780);
and UO_1617 (O_1617,N_19346,N_19698);
nand UO_1618 (O_1618,N_19737,N_19383);
nor UO_1619 (O_1619,N_19315,N_19930);
nand UO_1620 (O_1620,N_19618,N_19104);
nand UO_1621 (O_1621,N_19309,N_19476);
nor UO_1622 (O_1622,N_19827,N_19997);
xnor UO_1623 (O_1623,N_19199,N_19169);
nand UO_1624 (O_1624,N_19150,N_19446);
xor UO_1625 (O_1625,N_19534,N_19756);
and UO_1626 (O_1626,N_19151,N_19627);
nand UO_1627 (O_1627,N_19027,N_19144);
nand UO_1628 (O_1628,N_19520,N_19730);
xnor UO_1629 (O_1629,N_19326,N_19696);
or UO_1630 (O_1630,N_19984,N_19323);
or UO_1631 (O_1631,N_19807,N_19951);
nor UO_1632 (O_1632,N_19218,N_19974);
nand UO_1633 (O_1633,N_19734,N_19156);
nand UO_1634 (O_1634,N_19171,N_19867);
nand UO_1635 (O_1635,N_19550,N_19843);
nor UO_1636 (O_1636,N_19976,N_19269);
nor UO_1637 (O_1637,N_19421,N_19851);
xnor UO_1638 (O_1638,N_19186,N_19842);
and UO_1639 (O_1639,N_19738,N_19718);
or UO_1640 (O_1640,N_19463,N_19967);
xnor UO_1641 (O_1641,N_19981,N_19716);
and UO_1642 (O_1642,N_19328,N_19034);
nor UO_1643 (O_1643,N_19439,N_19740);
or UO_1644 (O_1644,N_19933,N_19939);
and UO_1645 (O_1645,N_19388,N_19283);
nand UO_1646 (O_1646,N_19238,N_19595);
nand UO_1647 (O_1647,N_19805,N_19078);
and UO_1648 (O_1648,N_19616,N_19228);
nor UO_1649 (O_1649,N_19400,N_19365);
nor UO_1650 (O_1650,N_19613,N_19510);
or UO_1651 (O_1651,N_19469,N_19329);
xor UO_1652 (O_1652,N_19888,N_19552);
and UO_1653 (O_1653,N_19659,N_19563);
nor UO_1654 (O_1654,N_19729,N_19519);
nand UO_1655 (O_1655,N_19621,N_19613);
nand UO_1656 (O_1656,N_19381,N_19956);
nor UO_1657 (O_1657,N_19923,N_19490);
nor UO_1658 (O_1658,N_19413,N_19980);
or UO_1659 (O_1659,N_19558,N_19707);
or UO_1660 (O_1660,N_19840,N_19786);
xnor UO_1661 (O_1661,N_19675,N_19981);
nor UO_1662 (O_1662,N_19639,N_19902);
nor UO_1663 (O_1663,N_19652,N_19557);
xnor UO_1664 (O_1664,N_19641,N_19488);
nor UO_1665 (O_1665,N_19980,N_19457);
or UO_1666 (O_1666,N_19284,N_19814);
and UO_1667 (O_1667,N_19606,N_19767);
or UO_1668 (O_1668,N_19708,N_19559);
nor UO_1669 (O_1669,N_19418,N_19780);
or UO_1670 (O_1670,N_19569,N_19901);
and UO_1671 (O_1671,N_19667,N_19948);
or UO_1672 (O_1672,N_19436,N_19020);
nand UO_1673 (O_1673,N_19607,N_19634);
nand UO_1674 (O_1674,N_19483,N_19055);
nor UO_1675 (O_1675,N_19304,N_19286);
or UO_1676 (O_1676,N_19884,N_19285);
or UO_1677 (O_1677,N_19718,N_19590);
xor UO_1678 (O_1678,N_19604,N_19568);
xnor UO_1679 (O_1679,N_19944,N_19377);
or UO_1680 (O_1680,N_19021,N_19410);
and UO_1681 (O_1681,N_19146,N_19811);
or UO_1682 (O_1682,N_19554,N_19116);
nor UO_1683 (O_1683,N_19045,N_19827);
nand UO_1684 (O_1684,N_19820,N_19973);
nor UO_1685 (O_1685,N_19496,N_19370);
and UO_1686 (O_1686,N_19490,N_19518);
xnor UO_1687 (O_1687,N_19232,N_19653);
nor UO_1688 (O_1688,N_19881,N_19088);
or UO_1689 (O_1689,N_19084,N_19190);
xor UO_1690 (O_1690,N_19172,N_19279);
nor UO_1691 (O_1691,N_19309,N_19642);
nand UO_1692 (O_1692,N_19637,N_19774);
nor UO_1693 (O_1693,N_19785,N_19923);
and UO_1694 (O_1694,N_19116,N_19042);
and UO_1695 (O_1695,N_19620,N_19287);
and UO_1696 (O_1696,N_19264,N_19731);
or UO_1697 (O_1697,N_19933,N_19573);
nand UO_1698 (O_1698,N_19592,N_19143);
xnor UO_1699 (O_1699,N_19588,N_19632);
nand UO_1700 (O_1700,N_19931,N_19075);
nand UO_1701 (O_1701,N_19569,N_19306);
nand UO_1702 (O_1702,N_19538,N_19475);
and UO_1703 (O_1703,N_19138,N_19108);
nor UO_1704 (O_1704,N_19398,N_19455);
nand UO_1705 (O_1705,N_19772,N_19198);
nand UO_1706 (O_1706,N_19782,N_19567);
and UO_1707 (O_1707,N_19948,N_19994);
nor UO_1708 (O_1708,N_19665,N_19431);
and UO_1709 (O_1709,N_19532,N_19981);
nor UO_1710 (O_1710,N_19657,N_19828);
or UO_1711 (O_1711,N_19219,N_19430);
and UO_1712 (O_1712,N_19742,N_19280);
xor UO_1713 (O_1713,N_19318,N_19836);
nand UO_1714 (O_1714,N_19739,N_19765);
nand UO_1715 (O_1715,N_19115,N_19137);
nor UO_1716 (O_1716,N_19899,N_19255);
or UO_1717 (O_1717,N_19365,N_19071);
and UO_1718 (O_1718,N_19314,N_19777);
nand UO_1719 (O_1719,N_19997,N_19195);
and UO_1720 (O_1720,N_19485,N_19308);
xor UO_1721 (O_1721,N_19457,N_19615);
nand UO_1722 (O_1722,N_19435,N_19713);
nor UO_1723 (O_1723,N_19862,N_19450);
xor UO_1724 (O_1724,N_19637,N_19423);
nor UO_1725 (O_1725,N_19692,N_19231);
or UO_1726 (O_1726,N_19565,N_19308);
xor UO_1727 (O_1727,N_19826,N_19736);
and UO_1728 (O_1728,N_19787,N_19461);
nor UO_1729 (O_1729,N_19999,N_19574);
or UO_1730 (O_1730,N_19947,N_19981);
nor UO_1731 (O_1731,N_19063,N_19998);
nor UO_1732 (O_1732,N_19976,N_19498);
xnor UO_1733 (O_1733,N_19739,N_19005);
nor UO_1734 (O_1734,N_19784,N_19968);
xnor UO_1735 (O_1735,N_19564,N_19836);
and UO_1736 (O_1736,N_19167,N_19889);
nand UO_1737 (O_1737,N_19752,N_19287);
xnor UO_1738 (O_1738,N_19132,N_19751);
nor UO_1739 (O_1739,N_19745,N_19330);
nand UO_1740 (O_1740,N_19323,N_19449);
nor UO_1741 (O_1741,N_19628,N_19969);
nor UO_1742 (O_1742,N_19331,N_19393);
nand UO_1743 (O_1743,N_19331,N_19764);
nor UO_1744 (O_1744,N_19768,N_19123);
xor UO_1745 (O_1745,N_19761,N_19663);
xor UO_1746 (O_1746,N_19726,N_19388);
nor UO_1747 (O_1747,N_19750,N_19365);
or UO_1748 (O_1748,N_19419,N_19202);
nand UO_1749 (O_1749,N_19805,N_19593);
and UO_1750 (O_1750,N_19646,N_19574);
xor UO_1751 (O_1751,N_19601,N_19555);
nor UO_1752 (O_1752,N_19863,N_19831);
nand UO_1753 (O_1753,N_19491,N_19896);
and UO_1754 (O_1754,N_19001,N_19675);
and UO_1755 (O_1755,N_19190,N_19443);
nor UO_1756 (O_1756,N_19534,N_19268);
xor UO_1757 (O_1757,N_19202,N_19072);
nor UO_1758 (O_1758,N_19443,N_19233);
xnor UO_1759 (O_1759,N_19717,N_19332);
nor UO_1760 (O_1760,N_19247,N_19516);
or UO_1761 (O_1761,N_19020,N_19600);
xor UO_1762 (O_1762,N_19768,N_19428);
and UO_1763 (O_1763,N_19497,N_19355);
xor UO_1764 (O_1764,N_19575,N_19727);
or UO_1765 (O_1765,N_19038,N_19750);
or UO_1766 (O_1766,N_19732,N_19736);
or UO_1767 (O_1767,N_19194,N_19959);
xor UO_1768 (O_1768,N_19118,N_19884);
nor UO_1769 (O_1769,N_19618,N_19132);
xor UO_1770 (O_1770,N_19006,N_19748);
nor UO_1771 (O_1771,N_19068,N_19611);
or UO_1772 (O_1772,N_19756,N_19129);
xnor UO_1773 (O_1773,N_19986,N_19021);
nand UO_1774 (O_1774,N_19559,N_19873);
or UO_1775 (O_1775,N_19619,N_19894);
nand UO_1776 (O_1776,N_19337,N_19494);
xor UO_1777 (O_1777,N_19343,N_19206);
xnor UO_1778 (O_1778,N_19228,N_19404);
nor UO_1779 (O_1779,N_19326,N_19955);
or UO_1780 (O_1780,N_19081,N_19115);
or UO_1781 (O_1781,N_19239,N_19538);
or UO_1782 (O_1782,N_19566,N_19127);
or UO_1783 (O_1783,N_19545,N_19020);
nor UO_1784 (O_1784,N_19075,N_19658);
and UO_1785 (O_1785,N_19271,N_19767);
and UO_1786 (O_1786,N_19127,N_19901);
xor UO_1787 (O_1787,N_19941,N_19892);
nor UO_1788 (O_1788,N_19324,N_19288);
and UO_1789 (O_1789,N_19237,N_19813);
nor UO_1790 (O_1790,N_19341,N_19584);
nand UO_1791 (O_1791,N_19649,N_19662);
and UO_1792 (O_1792,N_19682,N_19565);
and UO_1793 (O_1793,N_19732,N_19629);
nand UO_1794 (O_1794,N_19696,N_19650);
nand UO_1795 (O_1795,N_19629,N_19452);
or UO_1796 (O_1796,N_19724,N_19283);
or UO_1797 (O_1797,N_19182,N_19671);
and UO_1798 (O_1798,N_19892,N_19522);
or UO_1799 (O_1799,N_19286,N_19831);
xor UO_1800 (O_1800,N_19799,N_19295);
xnor UO_1801 (O_1801,N_19728,N_19438);
and UO_1802 (O_1802,N_19800,N_19393);
or UO_1803 (O_1803,N_19891,N_19979);
xor UO_1804 (O_1804,N_19661,N_19781);
nand UO_1805 (O_1805,N_19489,N_19635);
and UO_1806 (O_1806,N_19031,N_19084);
and UO_1807 (O_1807,N_19342,N_19284);
and UO_1808 (O_1808,N_19368,N_19528);
nand UO_1809 (O_1809,N_19331,N_19239);
nor UO_1810 (O_1810,N_19969,N_19743);
or UO_1811 (O_1811,N_19115,N_19463);
nor UO_1812 (O_1812,N_19138,N_19593);
xor UO_1813 (O_1813,N_19024,N_19863);
or UO_1814 (O_1814,N_19973,N_19111);
nand UO_1815 (O_1815,N_19548,N_19331);
xnor UO_1816 (O_1816,N_19030,N_19790);
nor UO_1817 (O_1817,N_19211,N_19471);
nand UO_1818 (O_1818,N_19186,N_19079);
or UO_1819 (O_1819,N_19817,N_19033);
and UO_1820 (O_1820,N_19701,N_19992);
nand UO_1821 (O_1821,N_19021,N_19192);
or UO_1822 (O_1822,N_19152,N_19100);
nand UO_1823 (O_1823,N_19534,N_19251);
nand UO_1824 (O_1824,N_19750,N_19587);
xor UO_1825 (O_1825,N_19996,N_19774);
nand UO_1826 (O_1826,N_19226,N_19294);
or UO_1827 (O_1827,N_19158,N_19282);
nand UO_1828 (O_1828,N_19156,N_19250);
xnor UO_1829 (O_1829,N_19603,N_19207);
xor UO_1830 (O_1830,N_19453,N_19100);
and UO_1831 (O_1831,N_19071,N_19211);
or UO_1832 (O_1832,N_19776,N_19012);
nor UO_1833 (O_1833,N_19896,N_19393);
xor UO_1834 (O_1834,N_19853,N_19311);
xnor UO_1835 (O_1835,N_19883,N_19587);
or UO_1836 (O_1836,N_19254,N_19324);
nor UO_1837 (O_1837,N_19164,N_19972);
xor UO_1838 (O_1838,N_19339,N_19572);
nor UO_1839 (O_1839,N_19184,N_19909);
nand UO_1840 (O_1840,N_19500,N_19136);
and UO_1841 (O_1841,N_19464,N_19693);
or UO_1842 (O_1842,N_19359,N_19010);
nor UO_1843 (O_1843,N_19683,N_19752);
and UO_1844 (O_1844,N_19781,N_19935);
or UO_1845 (O_1845,N_19360,N_19386);
nor UO_1846 (O_1846,N_19335,N_19068);
and UO_1847 (O_1847,N_19896,N_19969);
nand UO_1848 (O_1848,N_19509,N_19671);
nand UO_1849 (O_1849,N_19230,N_19052);
nand UO_1850 (O_1850,N_19880,N_19050);
xor UO_1851 (O_1851,N_19906,N_19832);
nand UO_1852 (O_1852,N_19240,N_19870);
or UO_1853 (O_1853,N_19817,N_19804);
xor UO_1854 (O_1854,N_19372,N_19008);
nor UO_1855 (O_1855,N_19416,N_19718);
nor UO_1856 (O_1856,N_19969,N_19115);
xor UO_1857 (O_1857,N_19606,N_19224);
nor UO_1858 (O_1858,N_19618,N_19429);
or UO_1859 (O_1859,N_19658,N_19766);
and UO_1860 (O_1860,N_19411,N_19846);
and UO_1861 (O_1861,N_19908,N_19896);
or UO_1862 (O_1862,N_19638,N_19161);
nand UO_1863 (O_1863,N_19906,N_19185);
xor UO_1864 (O_1864,N_19814,N_19537);
or UO_1865 (O_1865,N_19907,N_19427);
nand UO_1866 (O_1866,N_19086,N_19196);
nand UO_1867 (O_1867,N_19603,N_19536);
nor UO_1868 (O_1868,N_19806,N_19151);
nor UO_1869 (O_1869,N_19444,N_19844);
nor UO_1870 (O_1870,N_19182,N_19158);
nand UO_1871 (O_1871,N_19310,N_19848);
xor UO_1872 (O_1872,N_19497,N_19870);
nor UO_1873 (O_1873,N_19780,N_19770);
nand UO_1874 (O_1874,N_19694,N_19463);
xor UO_1875 (O_1875,N_19602,N_19070);
and UO_1876 (O_1876,N_19565,N_19154);
nand UO_1877 (O_1877,N_19575,N_19832);
xnor UO_1878 (O_1878,N_19201,N_19890);
and UO_1879 (O_1879,N_19652,N_19709);
xor UO_1880 (O_1880,N_19212,N_19602);
and UO_1881 (O_1881,N_19629,N_19992);
or UO_1882 (O_1882,N_19045,N_19019);
nor UO_1883 (O_1883,N_19156,N_19823);
or UO_1884 (O_1884,N_19810,N_19962);
nor UO_1885 (O_1885,N_19325,N_19586);
nand UO_1886 (O_1886,N_19626,N_19480);
nor UO_1887 (O_1887,N_19280,N_19795);
nor UO_1888 (O_1888,N_19679,N_19283);
nor UO_1889 (O_1889,N_19981,N_19253);
nand UO_1890 (O_1890,N_19704,N_19307);
or UO_1891 (O_1891,N_19201,N_19862);
xor UO_1892 (O_1892,N_19123,N_19092);
xnor UO_1893 (O_1893,N_19492,N_19816);
xor UO_1894 (O_1894,N_19393,N_19914);
nand UO_1895 (O_1895,N_19141,N_19411);
nand UO_1896 (O_1896,N_19446,N_19941);
nor UO_1897 (O_1897,N_19658,N_19474);
xor UO_1898 (O_1898,N_19140,N_19590);
or UO_1899 (O_1899,N_19450,N_19264);
nand UO_1900 (O_1900,N_19065,N_19330);
nand UO_1901 (O_1901,N_19188,N_19394);
xor UO_1902 (O_1902,N_19420,N_19592);
or UO_1903 (O_1903,N_19357,N_19819);
nor UO_1904 (O_1904,N_19774,N_19279);
nand UO_1905 (O_1905,N_19186,N_19455);
nor UO_1906 (O_1906,N_19518,N_19118);
and UO_1907 (O_1907,N_19714,N_19210);
or UO_1908 (O_1908,N_19793,N_19028);
nor UO_1909 (O_1909,N_19406,N_19137);
and UO_1910 (O_1910,N_19105,N_19836);
or UO_1911 (O_1911,N_19207,N_19477);
and UO_1912 (O_1912,N_19878,N_19747);
or UO_1913 (O_1913,N_19426,N_19999);
and UO_1914 (O_1914,N_19536,N_19301);
xnor UO_1915 (O_1915,N_19297,N_19987);
or UO_1916 (O_1916,N_19622,N_19035);
nor UO_1917 (O_1917,N_19382,N_19539);
or UO_1918 (O_1918,N_19721,N_19556);
nand UO_1919 (O_1919,N_19742,N_19316);
xor UO_1920 (O_1920,N_19564,N_19722);
xnor UO_1921 (O_1921,N_19321,N_19109);
and UO_1922 (O_1922,N_19485,N_19939);
nand UO_1923 (O_1923,N_19679,N_19464);
nand UO_1924 (O_1924,N_19604,N_19387);
or UO_1925 (O_1925,N_19270,N_19030);
nand UO_1926 (O_1926,N_19893,N_19615);
or UO_1927 (O_1927,N_19395,N_19935);
nor UO_1928 (O_1928,N_19663,N_19914);
or UO_1929 (O_1929,N_19288,N_19333);
nand UO_1930 (O_1930,N_19292,N_19623);
xor UO_1931 (O_1931,N_19359,N_19488);
or UO_1932 (O_1932,N_19470,N_19706);
xor UO_1933 (O_1933,N_19714,N_19956);
and UO_1934 (O_1934,N_19873,N_19178);
xnor UO_1935 (O_1935,N_19836,N_19011);
and UO_1936 (O_1936,N_19237,N_19928);
and UO_1937 (O_1937,N_19825,N_19525);
nand UO_1938 (O_1938,N_19236,N_19721);
xor UO_1939 (O_1939,N_19648,N_19133);
and UO_1940 (O_1940,N_19636,N_19914);
nand UO_1941 (O_1941,N_19135,N_19708);
and UO_1942 (O_1942,N_19712,N_19741);
and UO_1943 (O_1943,N_19028,N_19079);
nand UO_1944 (O_1944,N_19386,N_19312);
nand UO_1945 (O_1945,N_19439,N_19705);
nor UO_1946 (O_1946,N_19513,N_19345);
and UO_1947 (O_1947,N_19437,N_19130);
and UO_1948 (O_1948,N_19446,N_19563);
nor UO_1949 (O_1949,N_19721,N_19968);
nand UO_1950 (O_1950,N_19786,N_19629);
nand UO_1951 (O_1951,N_19623,N_19125);
nand UO_1952 (O_1952,N_19350,N_19613);
or UO_1953 (O_1953,N_19270,N_19094);
and UO_1954 (O_1954,N_19604,N_19505);
nand UO_1955 (O_1955,N_19771,N_19709);
and UO_1956 (O_1956,N_19670,N_19952);
or UO_1957 (O_1957,N_19227,N_19444);
or UO_1958 (O_1958,N_19455,N_19730);
or UO_1959 (O_1959,N_19823,N_19548);
or UO_1960 (O_1960,N_19497,N_19248);
nor UO_1961 (O_1961,N_19871,N_19166);
and UO_1962 (O_1962,N_19598,N_19802);
nor UO_1963 (O_1963,N_19319,N_19183);
nand UO_1964 (O_1964,N_19020,N_19773);
nor UO_1965 (O_1965,N_19531,N_19419);
or UO_1966 (O_1966,N_19913,N_19309);
and UO_1967 (O_1967,N_19692,N_19939);
and UO_1968 (O_1968,N_19696,N_19390);
nand UO_1969 (O_1969,N_19259,N_19640);
nand UO_1970 (O_1970,N_19613,N_19177);
and UO_1971 (O_1971,N_19377,N_19420);
nand UO_1972 (O_1972,N_19669,N_19341);
nand UO_1973 (O_1973,N_19419,N_19963);
xor UO_1974 (O_1974,N_19773,N_19494);
and UO_1975 (O_1975,N_19651,N_19243);
xor UO_1976 (O_1976,N_19314,N_19219);
or UO_1977 (O_1977,N_19403,N_19833);
xor UO_1978 (O_1978,N_19772,N_19656);
or UO_1979 (O_1979,N_19082,N_19590);
and UO_1980 (O_1980,N_19616,N_19559);
and UO_1981 (O_1981,N_19279,N_19613);
and UO_1982 (O_1982,N_19758,N_19559);
or UO_1983 (O_1983,N_19136,N_19764);
nand UO_1984 (O_1984,N_19280,N_19261);
and UO_1985 (O_1985,N_19881,N_19087);
nor UO_1986 (O_1986,N_19444,N_19571);
or UO_1987 (O_1987,N_19743,N_19448);
and UO_1988 (O_1988,N_19166,N_19603);
or UO_1989 (O_1989,N_19154,N_19169);
or UO_1990 (O_1990,N_19908,N_19539);
xor UO_1991 (O_1991,N_19468,N_19850);
and UO_1992 (O_1992,N_19053,N_19135);
xor UO_1993 (O_1993,N_19923,N_19565);
or UO_1994 (O_1994,N_19204,N_19082);
or UO_1995 (O_1995,N_19526,N_19861);
nand UO_1996 (O_1996,N_19052,N_19366);
and UO_1997 (O_1997,N_19557,N_19090);
or UO_1998 (O_1998,N_19100,N_19095);
xor UO_1999 (O_1999,N_19923,N_19094);
and UO_2000 (O_2000,N_19607,N_19590);
nand UO_2001 (O_2001,N_19071,N_19717);
xnor UO_2002 (O_2002,N_19905,N_19803);
nor UO_2003 (O_2003,N_19486,N_19411);
xnor UO_2004 (O_2004,N_19817,N_19627);
or UO_2005 (O_2005,N_19091,N_19167);
nand UO_2006 (O_2006,N_19586,N_19942);
xnor UO_2007 (O_2007,N_19263,N_19469);
nand UO_2008 (O_2008,N_19693,N_19085);
or UO_2009 (O_2009,N_19912,N_19023);
and UO_2010 (O_2010,N_19311,N_19405);
and UO_2011 (O_2011,N_19268,N_19926);
and UO_2012 (O_2012,N_19869,N_19912);
or UO_2013 (O_2013,N_19844,N_19599);
or UO_2014 (O_2014,N_19502,N_19324);
or UO_2015 (O_2015,N_19221,N_19017);
and UO_2016 (O_2016,N_19427,N_19933);
nand UO_2017 (O_2017,N_19434,N_19906);
or UO_2018 (O_2018,N_19279,N_19134);
xor UO_2019 (O_2019,N_19727,N_19111);
and UO_2020 (O_2020,N_19872,N_19444);
or UO_2021 (O_2021,N_19378,N_19020);
xnor UO_2022 (O_2022,N_19877,N_19960);
or UO_2023 (O_2023,N_19502,N_19959);
and UO_2024 (O_2024,N_19344,N_19483);
nand UO_2025 (O_2025,N_19155,N_19929);
nand UO_2026 (O_2026,N_19224,N_19673);
nor UO_2027 (O_2027,N_19301,N_19679);
and UO_2028 (O_2028,N_19464,N_19285);
and UO_2029 (O_2029,N_19683,N_19904);
nor UO_2030 (O_2030,N_19675,N_19068);
xor UO_2031 (O_2031,N_19866,N_19787);
xnor UO_2032 (O_2032,N_19058,N_19274);
and UO_2033 (O_2033,N_19199,N_19348);
xnor UO_2034 (O_2034,N_19845,N_19960);
nand UO_2035 (O_2035,N_19331,N_19781);
or UO_2036 (O_2036,N_19537,N_19125);
nor UO_2037 (O_2037,N_19919,N_19896);
nand UO_2038 (O_2038,N_19402,N_19838);
xnor UO_2039 (O_2039,N_19695,N_19885);
or UO_2040 (O_2040,N_19962,N_19765);
or UO_2041 (O_2041,N_19064,N_19014);
xor UO_2042 (O_2042,N_19011,N_19702);
nand UO_2043 (O_2043,N_19586,N_19068);
nor UO_2044 (O_2044,N_19239,N_19853);
nor UO_2045 (O_2045,N_19089,N_19834);
xor UO_2046 (O_2046,N_19316,N_19680);
xnor UO_2047 (O_2047,N_19144,N_19051);
nor UO_2048 (O_2048,N_19237,N_19654);
nor UO_2049 (O_2049,N_19083,N_19172);
xor UO_2050 (O_2050,N_19225,N_19148);
nor UO_2051 (O_2051,N_19444,N_19160);
nor UO_2052 (O_2052,N_19940,N_19643);
and UO_2053 (O_2053,N_19661,N_19587);
or UO_2054 (O_2054,N_19811,N_19584);
and UO_2055 (O_2055,N_19204,N_19974);
and UO_2056 (O_2056,N_19794,N_19441);
nand UO_2057 (O_2057,N_19855,N_19011);
xor UO_2058 (O_2058,N_19583,N_19905);
nor UO_2059 (O_2059,N_19673,N_19411);
or UO_2060 (O_2060,N_19130,N_19258);
or UO_2061 (O_2061,N_19493,N_19719);
and UO_2062 (O_2062,N_19797,N_19409);
xor UO_2063 (O_2063,N_19081,N_19107);
nand UO_2064 (O_2064,N_19053,N_19536);
nand UO_2065 (O_2065,N_19208,N_19518);
nor UO_2066 (O_2066,N_19946,N_19550);
or UO_2067 (O_2067,N_19471,N_19523);
nand UO_2068 (O_2068,N_19852,N_19965);
or UO_2069 (O_2069,N_19103,N_19321);
xnor UO_2070 (O_2070,N_19611,N_19509);
nor UO_2071 (O_2071,N_19240,N_19917);
and UO_2072 (O_2072,N_19387,N_19437);
and UO_2073 (O_2073,N_19795,N_19804);
nor UO_2074 (O_2074,N_19842,N_19800);
or UO_2075 (O_2075,N_19981,N_19215);
nand UO_2076 (O_2076,N_19844,N_19762);
and UO_2077 (O_2077,N_19785,N_19535);
and UO_2078 (O_2078,N_19645,N_19130);
and UO_2079 (O_2079,N_19821,N_19634);
or UO_2080 (O_2080,N_19423,N_19413);
nor UO_2081 (O_2081,N_19608,N_19948);
and UO_2082 (O_2082,N_19184,N_19212);
or UO_2083 (O_2083,N_19233,N_19877);
nand UO_2084 (O_2084,N_19687,N_19419);
nand UO_2085 (O_2085,N_19280,N_19072);
nand UO_2086 (O_2086,N_19663,N_19478);
xnor UO_2087 (O_2087,N_19530,N_19239);
xor UO_2088 (O_2088,N_19310,N_19160);
nand UO_2089 (O_2089,N_19268,N_19316);
nand UO_2090 (O_2090,N_19176,N_19852);
nand UO_2091 (O_2091,N_19241,N_19845);
xnor UO_2092 (O_2092,N_19292,N_19475);
and UO_2093 (O_2093,N_19892,N_19848);
nand UO_2094 (O_2094,N_19386,N_19149);
xor UO_2095 (O_2095,N_19760,N_19631);
xnor UO_2096 (O_2096,N_19482,N_19661);
and UO_2097 (O_2097,N_19178,N_19284);
nand UO_2098 (O_2098,N_19343,N_19554);
and UO_2099 (O_2099,N_19739,N_19974);
and UO_2100 (O_2100,N_19337,N_19161);
and UO_2101 (O_2101,N_19769,N_19570);
nor UO_2102 (O_2102,N_19675,N_19481);
and UO_2103 (O_2103,N_19052,N_19840);
and UO_2104 (O_2104,N_19008,N_19449);
nand UO_2105 (O_2105,N_19474,N_19162);
and UO_2106 (O_2106,N_19452,N_19136);
nand UO_2107 (O_2107,N_19206,N_19269);
xor UO_2108 (O_2108,N_19015,N_19536);
and UO_2109 (O_2109,N_19387,N_19285);
and UO_2110 (O_2110,N_19523,N_19227);
or UO_2111 (O_2111,N_19928,N_19293);
or UO_2112 (O_2112,N_19993,N_19241);
xnor UO_2113 (O_2113,N_19541,N_19240);
and UO_2114 (O_2114,N_19228,N_19472);
or UO_2115 (O_2115,N_19664,N_19613);
and UO_2116 (O_2116,N_19393,N_19978);
nor UO_2117 (O_2117,N_19937,N_19199);
or UO_2118 (O_2118,N_19514,N_19288);
nor UO_2119 (O_2119,N_19036,N_19362);
nor UO_2120 (O_2120,N_19847,N_19405);
nand UO_2121 (O_2121,N_19272,N_19722);
and UO_2122 (O_2122,N_19501,N_19119);
nand UO_2123 (O_2123,N_19693,N_19068);
nand UO_2124 (O_2124,N_19055,N_19171);
and UO_2125 (O_2125,N_19917,N_19103);
nor UO_2126 (O_2126,N_19273,N_19290);
nand UO_2127 (O_2127,N_19254,N_19134);
nand UO_2128 (O_2128,N_19580,N_19839);
nand UO_2129 (O_2129,N_19199,N_19340);
xnor UO_2130 (O_2130,N_19168,N_19090);
nor UO_2131 (O_2131,N_19549,N_19294);
xor UO_2132 (O_2132,N_19428,N_19872);
and UO_2133 (O_2133,N_19211,N_19699);
and UO_2134 (O_2134,N_19078,N_19444);
and UO_2135 (O_2135,N_19920,N_19739);
xor UO_2136 (O_2136,N_19001,N_19696);
nor UO_2137 (O_2137,N_19675,N_19257);
or UO_2138 (O_2138,N_19903,N_19743);
or UO_2139 (O_2139,N_19811,N_19830);
nor UO_2140 (O_2140,N_19285,N_19414);
nand UO_2141 (O_2141,N_19517,N_19029);
and UO_2142 (O_2142,N_19113,N_19903);
or UO_2143 (O_2143,N_19111,N_19240);
nand UO_2144 (O_2144,N_19098,N_19711);
nand UO_2145 (O_2145,N_19459,N_19453);
and UO_2146 (O_2146,N_19873,N_19843);
nor UO_2147 (O_2147,N_19650,N_19881);
xor UO_2148 (O_2148,N_19995,N_19783);
xnor UO_2149 (O_2149,N_19881,N_19202);
and UO_2150 (O_2150,N_19739,N_19969);
nand UO_2151 (O_2151,N_19799,N_19240);
nand UO_2152 (O_2152,N_19779,N_19529);
and UO_2153 (O_2153,N_19408,N_19043);
xnor UO_2154 (O_2154,N_19920,N_19742);
nand UO_2155 (O_2155,N_19013,N_19051);
xor UO_2156 (O_2156,N_19258,N_19772);
xnor UO_2157 (O_2157,N_19059,N_19234);
and UO_2158 (O_2158,N_19938,N_19369);
or UO_2159 (O_2159,N_19741,N_19552);
nor UO_2160 (O_2160,N_19618,N_19321);
xnor UO_2161 (O_2161,N_19951,N_19813);
nor UO_2162 (O_2162,N_19638,N_19431);
or UO_2163 (O_2163,N_19972,N_19330);
and UO_2164 (O_2164,N_19271,N_19705);
xnor UO_2165 (O_2165,N_19473,N_19603);
nor UO_2166 (O_2166,N_19682,N_19541);
and UO_2167 (O_2167,N_19080,N_19776);
nor UO_2168 (O_2168,N_19518,N_19888);
nand UO_2169 (O_2169,N_19662,N_19992);
xnor UO_2170 (O_2170,N_19163,N_19998);
and UO_2171 (O_2171,N_19220,N_19524);
nand UO_2172 (O_2172,N_19259,N_19209);
and UO_2173 (O_2173,N_19436,N_19402);
and UO_2174 (O_2174,N_19450,N_19056);
and UO_2175 (O_2175,N_19818,N_19021);
or UO_2176 (O_2176,N_19182,N_19148);
or UO_2177 (O_2177,N_19337,N_19786);
and UO_2178 (O_2178,N_19763,N_19486);
xor UO_2179 (O_2179,N_19538,N_19619);
nand UO_2180 (O_2180,N_19450,N_19243);
nand UO_2181 (O_2181,N_19364,N_19381);
xor UO_2182 (O_2182,N_19565,N_19989);
xnor UO_2183 (O_2183,N_19691,N_19899);
or UO_2184 (O_2184,N_19764,N_19168);
or UO_2185 (O_2185,N_19919,N_19892);
or UO_2186 (O_2186,N_19274,N_19118);
xnor UO_2187 (O_2187,N_19353,N_19711);
nor UO_2188 (O_2188,N_19073,N_19074);
xnor UO_2189 (O_2189,N_19582,N_19526);
and UO_2190 (O_2190,N_19456,N_19522);
and UO_2191 (O_2191,N_19857,N_19744);
nor UO_2192 (O_2192,N_19162,N_19620);
nor UO_2193 (O_2193,N_19565,N_19226);
nor UO_2194 (O_2194,N_19657,N_19975);
or UO_2195 (O_2195,N_19323,N_19538);
nor UO_2196 (O_2196,N_19997,N_19439);
xnor UO_2197 (O_2197,N_19134,N_19847);
nor UO_2198 (O_2198,N_19442,N_19025);
xnor UO_2199 (O_2199,N_19444,N_19393);
nand UO_2200 (O_2200,N_19960,N_19922);
or UO_2201 (O_2201,N_19926,N_19637);
or UO_2202 (O_2202,N_19999,N_19562);
nor UO_2203 (O_2203,N_19206,N_19737);
nor UO_2204 (O_2204,N_19175,N_19673);
and UO_2205 (O_2205,N_19142,N_19775);
and UO_2206 (O_2206,N_19600,N_19754);
and UO_2207 (O_2207,N_19550,N_19182);
xor UO_2208 (O_2208,N_19871,N_19758);
and UO_2209 (O_2209,N_19792,N_19112);
nor UO_2210 (O_2210,N_19412,N_19693);
nor UO_2211 (O_2211,N_19084,N_19454);
and UO_2212 (O_2212,N_19267,N_19436);
nor UO_2213 (O_2213,N_19818,N_19188);
and UO_2214 (O_2214,N_19521,N_19903);
nand UO_2215 (O_2215,N_19385,N_19745);
nand UO_2216 (O_2216,N_19656,N_19007);
nor UO_2217 (O_2217,N_19421,N_19524);
or UO_2218 (O_2218,N_19534,N_19292);
nor UO_2219 (O_2219,N_19865,N_19438);
xnor UO_2220 (O_2220,N_19112,N_19800);
nand UO_2221 (O_2221,N_19239,N_19865);
or UO_2222 (O_2222,N_19457,N_19904);
nor UO_2223 (O_2223,N_19417,N_19862);
or UO_2224 (O_2224,N_19077,N_19059);
and UO_2225 (O_2225,N_19265,N_19142);
xor UO_2226 (O_2226,N_19723,N_19674);
nand UO_2227 (O_2227,N_19931,N_19121);
and UO_2228 (O_2228,N_19566,N_19392);
or UO_2229 (O_2229,N_19339,N_19593);
nand UO_2230 (O_2230,N_19886,N_19761);
and UO_2231 (O_2231,N_19037,N_19759);
xor UO_2232 (O_2232,N_19938,N_19652);
or UO_2233 (O_2233,N_19958,N_19962);
nor UO_2234 (O_2234,N_19994,N_19602);
or UO_2235 (O_2235,N_19619,N_19636);
xor UO_2236 (O_2236,N_19788,N_19369);
and UO_2237 (O_2237,N_19410,N_19436);
nand UO_2238 (O_2238,N_19202,N_19920);
xnor UO_2239 (O_2239,N_19999,N_19123);
nand UO_2240 (O_2240,N_19721,N_19936);
and UO_2241 (O_2241,N_19386,N_19665);
or UO_2242 (O_2242,N_19791,N_19876);
or UO_2243 (O_2243,N_19020,N_19233);
and UO_2244 (O_2244,N_19948,N_19314);
nand UO_2245 (O_2245,N_19821,N_19226);
nand UO_2246 (O_2246,N_19727,N_19491);
and UO_2247 (O_2247,N_19834,N_19260);
and UO_2248 (O_2248,N_19038,N_19346);
nand UO_2249 (O_2249,N_19738,N_19366);
nor UO_2250 (O_2250,N_19391,N_19001);
nor UO_2251 (O_2251,N_19878,N_19381);
nor UO_2252 (O_2252,N_19614,N_19229);
nand UO_2253 (O_2253,N_19178,N_19707);
nor UO_2254 (O_2254,N_19427,N_19258);
xnor UO_2255 (O_2255,N_19671,N_19218);
or UO_2256 (O_2256,N_19917,N_19345);
and UO_2257 (O_2257,N_19923,N_19688);
xor UO_2258 (O_2258,N_19862,N_19321);
nand UO_2259 (O_2259,N_19024,N_19275);
and UO_2260 (O_2260,N_19351,N_19955);
and UO_2261 (O_2261,N_19324,N_19731);
nand UO_2262 (O_2262,N_19927,N_19496);
nand UO_2263 (O_2263,N_19957,N_19789);
and UO_2264 (O_2264,N_19258,N_19232);
xnor UO_2265 (O_2265,N_19554,N_19013);
and UO_2266 (O_2266,N_19857,N_19053);
and UO_2267 (O_2267,N_19895,N_19448);
nor UO_2268 (O_2268,N_19280,N_19933);
xor UO_2269 (O_2269,N_19640,N_19415);
and UO_2270 (O_2270,N_19548,N_19609);
xnor UO_2271 (O_2271,N_19688,N_19895);
or UO_2272 (O_2272,N_19905,N_19046);
nand UO_2273 (O_2273,N_19699,N_19477);
or UO_2274 (O_2274,N_19530,N_19198);
or UO_2275 (O_2275,N_19553,N_19086);
and UO_2276 (O_2276,N_19978,N_19937);
xnor UO_2277 (O_2277,N_19174,N_19161);
or UO_2278 (O_2278,N_19840,N_19114);
xnor UO_2279 (O_2279,N_19023,N_19571);
xor UO_2280 (O_2280,N_19265,N_19033);
nand UO_2281 (O_2281,N_19006,N_19762);
xnor UO_2282 (O_2282,N_19374,N_19343);
nor UO_2283 (O_2283,N_19685,N_19712);
and UO_2284 (O_2284,N_19806,N_19854);
or UO_2285 (O_2285,N_19023,N_19021);
nand UO_2286 (O_2286,N_19044,N_19250);
xnor UO_2287 (O_2287,N_19344,N_19361);
or UO_2288 (O_2288,N_19455,N_19447);
or UO_2289 (O_2289,N_19504,N_19997);
and UO_2290 (O_2290,N_19894,N_19951);
or UO_2291 (O_2291,N_19767,N_19547);
nor UO_2292 (O_2292,N_19104,N_19669);
and UO_2293 (O_2293,N_19978,N_19889);
nand UO_2294 (O_2294,N_19202,N_19807);
nand UO_2295 (O_2295,N_19311,N_19870);
and UO_2296 (O_2296,N_19415,N_19990);
xor UO_2297 (O_2297,N_19987,N_19645);
nor UO_2298 (O_2298,N_19363,N_19426);
xnor UO_2299 (O_2299,N_19742,N_19250);
and UO_2300 (O_2300,N_19563,N_19060);
nor UO_2301 (O_2301,N_19985,N_19653);
nor UO_2302 (O_2302,N_19083,N_19450);
nand UO_2303 (O_2303,N_19180,N_19973);
or UO_2304 (O_2304,N_19623,N_19514);
nand UO_2305 (O_2305,N_19725,N_19258);
nand UO_2306 (O_2306,N_19271,N_19855);
and UO_2307 (O_2307,N_19982,N_19018);
or UO_2308 (O_2308,N_19660,N_19385);
or UO_2309 (O_2309,N_19482,N_19886);
or UO_2310 (O_2310,N_19399,N_19863);
nand UO_2311 (O_2311,N_19303,N_19074);
nand UO_2312 (O_2312,N_19526,N_19581);
nand UO_2313 (O_2313,N_19219,N_19926);
nand UO_2314 (O_2314,N_19778,N_19658);
nand UO_2315 (O_2315,N_19604,N_19260);
or UO_2316 (O_2316,N_19182,N_19163);
nand UO_2317 (O_2317,N_19029,N_19154);
or UO_2318 (O_2318,N_19786,N_19884);
and UO_2319 (O_2319,N_19510,N_19546);
nand UO_2320 (O_2320,N_19774,N_19982);
or UO_2321 (O_2321,N_19306,N_19559);
nand UO_2322 (O_2322,N_19528,N_19994);
xnor UO_2323 (O_2323,N_19526,N_19771);
nand UO_2324 (O_2324,N_19245,N_19660);
or UO_2325 (O_2325,N_19723,N_19795);
xnor UO_2326 (O_2326,N_19020,N_19173);
nor UO_2327 (O_2327,N_19350,N_19330);
or UO_2328 (O_2328,N_19110,N_19993);
nand UO_2329 (O_2329,N_19311,N_19253);
or UO_2330 (O_2330,N_19112,N_19462);
xor UO_2331 (O_2331,N_19704,N_19039);
and UO_2332 (O_2332,N_19014,N_19277);
nand UO_2333 (O_2333,N_19902,N_19091);
nand UO_2334 (O_2334,N_19034,N_19594);
nor UO_2335 (O_2335,N_19697,N_19204);
or UO_2336 (O_2336,N_19761,N_19799);
and UO_2337 (O_2337,N_19038,N_19986);
nor UO_2338 (O_2338,N_19597,N_19513);
nor UO_2339 (O_2339,N_19133,N_19992);
nand UO_2340 (O_2340,N_19192,N_19533);
and UO_2341 (O_2341,N_19514,N_19626);
or UO_2342 (O_2342,N_19845,N_19846);
xor UO_2343 (O_2343,N_19558,N_19201);
and UO_2344 (O_2344,N_19730,N_19649);
nand UO_2345 (O_2345,N_19696,N_19659);
nand UO_2346 (O_2346,N_19611,N_19524);
xor UO_2347 (O_2347,N_19261,N_19065);
nand UO_2348 (O_2348,N_19297,N_19767);
nand UO_2349 (O_2349,N_19793,N_19232);
nor UO_2350 (O_2350,N_19839,N_19320);
nand UO_2351 (O_2351,N_19158,N_19070);
nand UO_2352 (O_2352,N_19113,N_19878);
nand UO_2353 (O_2353,N_19756,N_19335);
nor UO_2354 (O_2354,N_19814,N_19692);
or UO_2355 (O_2355,N_19851,N_19152);
nor UO_2356 (O_2356,N_19731,N_19025);
nand UO_2357 (O_2357,N_19549,N_19972);
and UO_2358 (O_2358,N_19952,N_19875);
nor UO_2359 (O_2359,N_19322,N_19848);
xor UO_2360 (O_2360,N_19824,N_19848);
or UO_2361 (O_2361,N_19489,N_19679);
and UO_2362 (O_2362,N_19886,N_19349);
or UO_2363 (O_2363,N_19966,N_19607);
and UO_2364 (O_2364,N_19111,N_19378);
nor UO_2365 (O_2365,N_19258,N_19343);
nand UO_2366 (O_2366,N_19039,N_19825);
nor UO_2367 (O_2367,N_19839,N_19216);
and UO_2368 (O_2368,N_19076,N_19430);
and UO_2369 (O_2369,N_19643,N_19434);
nand UO_2370 (O_2370,N_19929,N_19024);
or UO_2371 (O_2371,N_19106,N_19530);
and UO_2372 (O_2372,N_19758,N_19697);
and UO_2373 (O_2373,N_19621,N_19815);
nand UO_2374 (O_2374,N_19889,N_19745);
xnor UO_2375 (O_2375,N_19819,N_19750);
xnor UO_2376 (O_2376,N_19273,N_19178);
nand UO_2377 (O_2377,N_19169,N_19897);
and UO_2378 (O_2378,N_19487,N_19125);
and UO_2379 (O_2379,N_19035,N_19996);
and UO_2380 (O_2380,N_19042,N_19809);
or UO_2381 (O_2381,N_19748,N_19402);
xnor UO_2382 (O_2382,N_19462,N_19689);
or UO_2383 (O_2383,N_19594,N_19189);
nor UO_2384 (O_2384,N_19699,N_19426);
nor UO_2385 (O_2385,N_19387,N_19003);
nor UO_2386 (O_2386,N_19977,N_19203);
nand UO_2387 (O_2387,N_19886,N_19692);
or UO_2388 (O_2388,N_19021,N_19682);
or UO_2389 (O_2389,N_19892,N_19530);
xor UO_2390 (O_2390,N_19243,N_19255);
xnor UO_2391 (O_2391,N_19209,N_19479);
xor UO_2392 (O_2392,N_19407,N_19400);
and UO_2393 (O_2393,N_19599,N_19005);
and UO_2394 (O_2394,N_19525,N_19051);
nand UO_2395 (O_2395,N_19748,N_19072);
xor UO_2396 (O_2396,N_19855,N_19844);
nand UO_2397 (O_2397,N_19511,N_19192);
and UO_2398 (O_2398,N_19119,N_19538);
nand UO_2399 (O_2399,N_19557,N_19949);
nor UO_2400 (O_2400,N_19091,N_19600);
nor UO_2401 (O_2401,N_19694,N_19387);
nand UO_2402 (O_2402,N_19070,N_19200);
nand UO_2403 (O_2403,N_19540,N_19721);
nand UO_2404 (O_2404,N_19460,N_19515);
xnor UO_2405 (O_2405,N_19861,N_19841);
nor UO_2406 (O_2406,N_19089,N_19001);
xor UO_2407 (O_2407,N_19010,N_19880);
nor UO_2408 (O_2408,N_19484,N_19215);
nor UO_2409 (O_2409,N_19260,N_19138);
nand UO_2410 (O_2410,N_19505,N_19397);
or UO_2411 (O_2411,N_19975,N_19082);
nand UO_2412 (O_2412,N_19467,N_19976);
nand UO_2413 (O_2413,N_19528,N_19310);
and UO_2414 (O_2414,N_19759,N_19027);
nor UO_2415 (O_2415,N_19851,N_19543);
and UO_2416 (O_2416,N_19688,N_19656);
nand UO_2417 (O_2417,N_19592,N_19071);
and UO_2418 (O_2418,N_19719,N_19008);
nand UO_2419 (O_2419,N_19002,N_19495);
nand UO_2420 (O_2420,N_19729,N_19451);
xor UO_2421 (O_2421,N_19919,N_19929);
xor UO_2422 (O_2422,N_19715,N_19685);
xor UO_2423 (O_2423,N_19074,N_19295);
and UO_2424 (O_2424,N_19488,N_19838);
and UO_2425 (O_2425,N_19251,N_19325);
and UO_2426 (O_2426,N_19611,N_19799);
nand UO_2427 (O_2427,N_19581,N_19879);
nor UO_2428 (O_2428,N_19215,N_19008);
nand UO_2429 (O_2429,N_19379,N_19022);
nor UO_2430 (O_2430,N_19144,N_19015);
nand UO_2431 (O_2431,N_19956,N_19774);
nor UO_2432 (O_2432,N_19511,N_19254);
nor UO_2433 (O_2433,N_19729,N_19986);
or UO_2434 (O_2434,N_19493,N_19935);
or UO_2435 (O_2435,N_19718,N_19629);
and UO_2436 (O_2436,N_19090,N_19596);
or UO_2437 (O_2437,N_19193,N_19546);
or UO_2438 (O_2438,N_19932,N_19749);
nand UO_2439 (O_2439,N_19424,N_19517);
xnor UO_2440 (O_2440,N_19099,N_19640);
xor UO_2441 (O_2441,N_19177,N_19178);
or UO_2442 (O_2442,N_19884,N_19813);
nand UO_2443 (O_2443,N_19128,N_19189);
nand UO_2444 (O_2444,N_19948,N_19545);
nor UO_2445 (O_2445,N_19338,N_19350);
or UO_2446 (O_2446,N_19008,N_19166);
or UO_2447 (O_2447,N_19197,N_19175);
and UO_2448 (O_2448,N_19850,N_19999);
xor UO_2449 (O_2449,N_19157,N_19379);
nor UO_2450 (O_2450,N_19484,N_19867);
nand UO_2451 (O_2451,N_19933,N_19894);
or UO_2452 (O_2452,N_19909,N_19077);
or UO_2453 (O_2453,N_19420,N_19715);
or UO_2454 (O_2454,N_19296,N_19354);
xnor UO_2455 (O_2455,N_19136,N_19282);
xnor UO_2456 (O_2456,N_19803,N_19024);
nor UO_2457 (O_2457,N_19022,N_19802);
and UO_2458 (O_2458,N_19801,N_19509);
and UO_2459 (O_2459,N_19131,N_19252);
nor UO_2460 (O_2460,N_19284,N_19430);
or UO_2461 (O_2461,N_19686,N_19924);
xor UO_2462 (O_2462,N_19150,N_19718);
nor UO_2463 (O_2463,N_19595,N_19127);
xor UO_2464 (O_2464,N_19185,N_19728);
nor UO_2465 (O_2465,N_19358,N_19366);
or UO_2466 (O_2466,N_19897,N_19586);
xnor UO_2467 (O_2467,N_19110,N_19978);
nor UO_2468 (O_2468,N_19228,N_19331);
xnor UO_2469 (O_2469,N_19604,N_19204);
nand UO_2470 (O_2470,N_19143,N_19664);
xnor UO_2471 (O_2471,N_19506,N_19915);
nand UO_2472 (O_2472,N_19846,N_19567);
and UO_2473 (O_2473,N_19295,N_19498);
or UO_2474 (O_2474,N_19528,N_19165);
or UO_2475 (O_2475,N_19834,N_19014);
or UO_2476 (O_2476,N_19129,N_19994);
nor UO_2477 (O_2477,N_19921,N_19612);
xnor UO_2478 (O_2478,N_19791,N_19276);
nand UO_2479 (O_2479,N_19474,N_19318);
xnor UO_2480 (O_2480,N_19093,N_19039);
or UO_2481 (O_2481,N_19425,N_19032);
and UO_2482 (O_2482,N_19861,N_19451);
or UO_2483 (O_2483,N_19181,N_19298);
nand UO_2484 (O_2484,N_19055,N_19271);
and UO_2485 (O_2485,N_19643,N_19132);
nand UO_2486 (O_2486,N_19835,N_19104);
nand UO_2487 (O_2487,N_19653,N_19179);
nor UO_2488 (O_2488,N_19482,N_19744);
or UO_2489 (O_2489,N_19163,N_19842);
or UO_2490 (O_2490,N_19498,N_19985);
or UO_2491 (O_2491,N_19468,N_19205);
and UO_2492 (O_2492,N_19190,N_19287);
xnor UO_2493 (O_2493,N_19871,N_19601);
nand UO_2494 (O_2494,N_19900,N_19817);
nand UO_2495 (O_2495,N_19341,N_19375);
and UO_2496 (O_2496,N_19029,N_19406);
nand UO_2497 (O_2497,N_19080,N_19808);
and UO_2498 (O_2498,N_19498,N_19962);
or UO_2499 (O_2499,N_19278,N_19501);
endmodule