module basic_5000_50000_5000_100_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nor U0 (N_0,In_4518,In_2589);
and U1 (N_1,In_1462,In_4769);
nor U2 (N_2,In_134,In_1024);
or U3 (N_3,In_1264,In_4446);
nand U4 (N_4,In_2210,In_170);
nor U5 (N_5,In_2239,In_1240);
xor U6 (N_6,In_691,In_4013);
and U7 (N_7,In_3874,In_1442);
or U8 (N_8,In_122,In_1116);
and U9 (N_9,In_1784,In_594);
or U10 (N_10,In_2095,In_4742);
nand U11 (N_11,In_2011,In_264);
xor U12 (N_12,In_496,In_1661);
xnor U13 (N_13,In_1975,In_442);
and U14 (N_14,In_148,In_149);
nand U15 (N_15,In_4749,In_4230);
nor U16 (N_16,In_1514,In_4824);
or U17 (N_17,In_4234,In_3770);
or U18 (N_18,In_4866,In_280);
nand U19 (N_19,In_3401,In_2996);
and U20 (N_20,In_3553,In_3150);
nor U21 (N_21,In_2756,In_958);
xnor U22 (N_22,In_4386,In_3124);
nor U23 (N_23,In_692,In_2271);
or U24 (N_24,In_4081,In_1775);
xnor U25 (N_25,In_210,In_3190);
xor U26 (N_26,In_23,In_4347);
xnor U27 (N_27,In_887,In_1303);
xnor U28 (N_28,In_2433,In_1954);
nor U29 (N_29,In_4397,In_2569);
nand U30 (N_30,In_3162,In_1943);
xnor U31 (N_31,In_4456,In_3308);
nor U32 (N_32,In_2423,In_1557);
xnor U33 (N_33,In_3810,In_1237);
xor U34 (N_34,In_4025,In_3517);
nor U35 (N_35,In_4245,In_3009);
and U36 (N_36,In_855,In_1534);
xor U37 (N_37,In_1750,In_3490);
xor U38 (N_38,In_2751,In_3706);
and U39 (N_39,In_3645,In_3351);
xor U40 (N_40,In_2713,In_2376);
xnor U41 (N_41,In_1829,In_4030);
xor U42 (N_42,In_3236,In_4544);
or U43 (N_43,In_4437,In_3507);
and U44 (N_44,In_1208,In_258);
or U45 (N_45,In_172,In_3172);
or U46 (N_46,In_4335,In_435);
xnor U47 (N_47,In_4843,In_3203);
nand U48 (N_48,In_4402,In_1443);
nor U49 (N_49,In_3878,In_3417);
nand U50 (N_50,In_4344,In_3514);
and U51 (N_51,In_2829,In_4558);
nor U52 (N_52,In_1914,In_758);
nor U53 (N_53,In_2819,In_1586);
and U54 (N_54,In_3361,In_1444);
nand U55 (N_55,In_3885,In_1124);
or U56 (N_56,In_3021,In_3423);
xnor U57 (N_57,In_4032,In_2428);
xnor U58 (N_58,In_3720,In_1753);
nand U59 (N_59,In_4110,In_4348);
nand U60 (N_60,In_2048,In_1603);
xor U61 (N_61,In_1007,In_4736);
or U62 (N_62,In_3750,In_3733);
and U63 (N_63,In_4382,In_1133);
or U64 (N_64,In_3930,In_2692);
nand U65 (N_65,In_4350,In_3126);
and U66 (N_66,In_614,In_4209);
and U67 (N_67,In_198,In_420);
or U68 (N_68,In_493,In_1405);
and U69 (N_69,In_1059,In_3287);
nand U70 (N_70,In_4557,In_1396);
xor U71 (N_71,In_3948,In_2820);
xnor U72 (N_72,In_3356,In_2273);
nor U73 (N_73,In_2491,In_2971);
or U74 (N_74,In_1822,In_4552);
xor U75 (N_75,In_2290,In_2650);
nor U76 (N_76,In_1003,In_2278);
and U77 (N_77,In_1217,In_3574);
nor U78 (N_78,In_1715,In_3786);
nand U79 (N_79,In_3146,In_632);
nand U80 (N_80,In_3915,In_2289);
xor U81 (N_81,In_777,In_555);
xor U82 (N_82,In_4137,In_1823);
and U83 (N_83,In_3484,In_3630);
or U84 (N_84,In_4037,In_2131);
and U85 (N_85,In_3396,In_4265);
and U86 (N_86,In_3034,In_764);
xnor U87 (N_87,In_4249,In_4331);
nor U88 (N_88,In_4683,In_584);
nor U89 (N_89,In_4170,In_797);
nand U90 (N_90,In_3867,In_3041);
and U91 (N_91,In_1229,In_1626);
or U92 (N_92,In_747,In_294);
nand U93 (N_93,In_3188,In_2274);
nor U94 (N_94,In_979,In_59);
and U95 (N_95,In_4050,In_1330);
xnor U96 (N_96,In_4553,In_3555);
nor U97 (N_97,In_1358,In_1723);
xnor U98 (N_98,In_1387,In_1097);
xor U99 (N_99,In_1515,In_3213);
and U100 (N_100,In_4618,In_4722);
nand U101 (N_101,In_377,In_852);
and U102 (N_102,In_3871,In_4120);
nand U103 (N_103,In_2066,In_997);
xnor U104 (N_104,In_1786,In_1493);
nand U105 (N_105,In_61,In_2938);
or U106 (N_106,In_446,In_1367);
nor U107 (N_107,In_1298,In_2633);
xor U108 (N_108,In_4966,In_728);
or U109 (N_109,In_2434,In_3136);
xnor U110 (N_110,In_4235,In_3420);
nand U111 (N_111,In_882,In_663);
and U112 (N_112,In_1041,In_3407);
and U113 (N_113,In_4589,In_1351);
nor U114 (N_114,In_3740,In_2874);
and U115 (N_115,In_638,In_4965);
or U116 (N_116,In_4391,In_3833);
nor U117 (N_117,In_2679,In_4690);
nand U118 (N_118,In_3559,In_2825);
and U119 (N_119,In_1608,In_4969);
nand U120 (N_120,In_3233,In_4284);
xnor U121 (N_121,In_1350,In_3208);
xor U122 (N_122,In_1123,In_2361);
nand U123 (N_123,In_4416,In_3096);
nand U124 (N_124,In_88,In_291);
and U125 (N_125,In_679,In_1166);
or U126 (N_126,In_3971,In_4949);
xnor U127 (N_127,In_2364,In_4474);
xor U128 (N_128,In_1998,In_1917);
or U129 (N_129,In_3301,In_1406);
nor U130 (N_130,In_552,In_4042);
and U131 (N_131,In_4673,In_4621);
nor U132 (N_132,In_3257,In_3191);
and U133 (N_133,In_429,In_1275);
xor U134 (N_134,In_1507,In_4859);
xor U135 (N_135,In_4596,In_4577);
nand U136 (N_136,In_1802,In_26);
xor U137 (N_137,In_383,In_567);
xnor U138 (N_138,In_2074,In_1570);
nor U139 (N_139,In_2069,In_3322);
or U140 (N_140,In_4222,In_4327);
nand U141 (N_141,In_3102,In_1461);
nand U142 (N_142,In_1466,In_1565);
or U143 (N_143,In_2730,In_1252);
nor U144 (N_144,In_3370,In_1294);
or U145 (N_145,In_3105,In_4444);
xor U146 (N_146,In_717,In_3455);
or U147 (N_147,In_635,In_538);
xnor U148 (N_148,In_4164,In_1632);
xor U149 (N_149,In_1291,In_1571);
nor U150 (N_150,In_454,In_4539);
and U151 (N_151,In_2701,In_1747);
and U152 (N_152,In_244,In_844);
nor U153 (N_153,In_4049,In_2107);
nor U154 (N_154,In_3134,In_413);
nor U155 (N_155,In_1642,In_677);
and U156 (N_156,In_2313,In_1238);
or U157 (N_157,In_275,In_1511);
and U158 (N_158,In_1079,In_666);
and U159 (N_159,In_741,In_3580);
and U160 (N_160,In_3563,In_4771);
xor U161 (N_161,In_690,In_2538);
xnor U162 (N_162,In_4306,In_397);
or U163 (N_163,In_4183,In_4920);
and U164 (N_164,In_3234,In_439);
nor U165 (N_165,In_3358,In_1029);
nor U166 (N_166,In_4935,In_1142);
nor U167 (N_167,In_2956,In_1114);
nor U168 (N_168,In_311,In_3639);
nor U169 (N_169,In_4128,In_1796);
or U170 (N_170,In_1213,In_4294);
nor U171 (N_171,In_2417,In_3889);
nor U172 (N_172,In_536,In_3367);
nand U173 (N_173,In_4364,In_2223);
xor U174 (N_174,In_1117,In_1038);
nor U175 (N_175,In_477,In_3073);
and U176 (N_176,In_3952,In_3863);
and U177 (N_177,In_4886,In_3070);
and U178 (N_178,In_4072,In_898);
xor U179 (N_179,In_4520,In_3695);
xnor U180 (N_180,In_4898,In_4658);
nand U181 (N_181,In_3687,In_3088);
or U182 (N_182,In_527,In_4157);
or U183 (N_183,In_3112,In_4940);
nor U184 (N_184,In_742,In_2081);
and U185 (N_185,In_2112,In_1157);
nor U186 (N_186,In_1884,In_1370);
xor U187 (N_187,In_3503,In_2435);
xor U188 (N_188,In_1339,In_4214);
nor U189 (N_189,In_4681,In_4916);
nand U190 (N_190,In_27,In_2916);
nor U191 (N_191,In_3340,In_3918);
nor U192 (N_192,In_3842,In_3520);
nand U193 (N_193,In_1997,In_3155);
and U194 (N_194,In_1471,In_4950);
nor U195 (N_195,In_1563,In_1393);
nand U196 (N_196,In_4146,In_4185);
xor U197 (N_197,In_700,In_3390);
or U198 (N_198,In_2928,In_4560);
nand U199 (N_199,In_4738,In_3543);
and U200 (N_200,In_2685,In_600);
nand U201 (N_201,In_4528,In_873);
nor U202 (N_202,In_287,In_3135);
nor U203 (N_203,In_2248,In_1840);
xnor U204 (N_204,In_3628,In_1309);
xor U205 (N_205,In_4286,In_1055);
nand U206 (N_206,In_1233,In_3201);
and U207 (N_207,In_458,In_2545);
xor U208 (N_208,In_1800,In_3196);
nand U209 (N_209,In_2053,In_3876);
and U210 (N_210,In_2476,In_4430);
nand U211 (N_211,In_1076,In_4776);
or U212 (N_212,In_3068,In_1872);
and U213 (N_213,In_4302,In_4357);
or U214 (N_214,In_4808,In_3209);
nor U215 (N_215,In_1268,In_4063);
or U216 (N_216,In_2805,In_1052);
nor U217 (N_217,In_3526,In_3508);
xor U218 (N_218,In_4586,In_39);
or U219 (N_219,In_1323,In_4166);
and U220 (N_220,In_3785,In_3087);
or U221 (N_221,In_1057,In_4826);
nand U222 (N_222,In_1843,In_987);
xor U223 (N_223,In_2054,In_631);
xor U224 (N_224,In_409,In_2853);
or U225 (N_225,In_908,In_1936);
nand U226 (N_226,In_4133,In_4008);
xnor U227 (N_227,In_2795,In_1799);
or U228 (N_228,In_3716,In_1134);
nor U229 (N_229,In_799,In_4656);
or U230 (N_230,In_593,In_1995);
or U231 (N_231,In_35,In_967);
nor U232 (N_232,In_3540,In_181);
and U233 (N_233,In_1904,In_2903);
or U234 (N_234,In_2905,In_2846);
xor U235 (N_235,In_2587,In_858);
xnor U236 (N_236,In_2940,In_2894);
and U237 (N_237,In_1266,In_3238);
nand U238 (N_238,In_1216,In_1315);
or U239 (N_239,In_206,In_1903);
xor U240 (N_240,In_2534,In_1207);
and U241 (N_241,In_515,In_4454);
xor U242 (N_242,In_1646,In_3374);
nor U243 (N_243,In_2718,In_30);
xnor U244 (N_244,In_2691,In_644);
xor U245 (N_245,In_338,In_4423);
nor U246 (N_246,In_4927,In_4819);
nand U247 (N_247,In_347,In_460);
and U248 (N_248,In_681,In_3935);
xor U249 (N_249,In_3832,In_2533);
xor U250 (N_250,In_1607,In_4129);
nor U251 (N_251,In_1101,In_2407);
nand U252 (N_252,In_2658,In_3524);
nand U253 (N_253,In_924,In_2590);
xor U254 (N_254,In_1824,In_3428);
nand U255 (N_255,In_1736,In_1137);
xnor U256 (N_256,In_1568,In_2686);
or U257 (N_257,In_2158,In_798);
nand U258 (N_258,In_4256,In_619);
nand U259 (N_259,In_3133,In_1011);
nor U260 (N_260,In_1484,In_3035);
or U261 (N_261,In_835,In_621);
nor U262 (N_262,In_748,In_55);
nand U263 (N_263,In_3485,In_467);
nand U264 (N_264,In_4010,In_2960);
nor U265 (N_265,In_1807,In_297);
nor U266 (N_266,In_2327,In_260);
and U267 (N_267,In_4436,In_2465);
or U268 (N_268,In_365,In_994);
and U269 (N_269,In_3166,In_1528);
nor U270 (N_270,In_2839,In_2194);
and U271 (N_271,In_3311,In_4896);
xnor U272 (N_272,In_2547,In_1553);
xnor U273 (N_273,In_3446,In_453);
and U274 (N_274,In_607,In_658);
nor U275 (N_275,In_1707,In_380);
xnor U276 (N_276,In_2866,In_2259);
nor U277 (N_277,In_2108,In_1404);
and U278 (N_278,In_884,In_2989);
nor U279 (N_279,In_2240,In_3788);
nor U280 (N_280,In_2717,In_1815);
xnor U281 (N_281,In_3764,In_3572);
or U282 (N_282,In_4753,In_1619);
nor U283 (N_283,In_1422,In_2539);
and U284 (N_284,In_1714,In_2864);
xnor U285 (N_285,In_3159,In_3506);
nand U286 (N_286,In_976,In_4989);
nor U287 (N_287,In_2260,In_652);
nand U288 (N_288,In_2437,In_2621);
nand U289 (N_289,In_1073,In_1548);
nand U290 (N_290,In_3461,In_808);
and U291 (N_291,In_837,In_2027);
and U292 (N_292,In_3144,In_4404);
xor U293 (N_293,In_434,In_615);
nand U294 (N_294,In_931,In_4317);
nand U295 (N_295,In_4913,In_2325);
or U296 (N_296,In_1105,In_2934);
or U297 (N_297,In_2560,In_4804);
nand U298 (N_298,In_2385,In_426);
or U299 (N_299,In_1956,In_719);
xor U300 (N_300,In_1674,In_4014);
or U301 (N_301,In_2127,In_2766);
or U302 (N_302,In_346,In_216);
nor U303 (N_303,In_647,In_3758);
nand U304 (N_304,In_4221,In_226);
nor U305 (N_305,In_3773,In_1803);
nor U306 (N_306,In_3542,In_2955);
or U307 (N_307,In_3696,In_375);
and U308 (N_308,In_2164,In_281);
nand U309 (N_309,In_403,In_4073);
nor U310 (N_310,In_1968,In_4272);
and U311 (N_311,In_1509,In_1869);
nand U312 (N_312,In_2370,In_4904);
xor U313 (N_313,In_488,In_1670);
nand U314 (N_314,In_1182,In_2077);
and U315 (N_315,In_456,In_613);
nand U316 (N_316,In_2716,In_1795);
nor U317 (N_317,In_1770,In_4239);
xnor U318 (N_318,In_3215,In_2858);
or U319 (N_319,In_1751,In_4017);
xor U320 (N_320,In_2654,In_475);
nand U321 (N_321,In_2205,In_1470);
nand U322 (N_322,In_2337,In_885);
or U323 (N_323,In_3015,In_1749);
or U324 (N_324,In_4887,In_3847);
nor U325 (N_325,In_4938,In_29);
or U326 (N_326,In_1044,In_286);
and U327 (N_327,In_4748,In_94);
nand U328 (N_328,In_4836,In_1641);
nand U329 (N_329,In_1728,In_2332);
nor U330 (N_330,In_4287,In_3307);
xor U331 (N_331,In_2229,In_2034);
or U332 (N_332,In_1478,In_4842);
and U333 (N_333,In_2005,In_2958);
or U334 (N_334,In_1226,In_1644);
nand U335 (N_335,In_3382,In_66);
nor U336 (N_336,In_3327,In_4572);
xnor U337 (N_337,In_1152,In_100);
nor U338 (N_338,In_4136,In_4280);
or U339 (N_339,In_2634,In_3496);
or U340 (N_340,In_1196,In_3268);
and U341 (N_341,In_1527,In_1870);
or U342 (N_342,In_4784,In_4699);
xnor U343 (N_343,In_4298,In_3602);
or U344 (N_344,In_4433,In_1389);
and U345 (N_345,In_1598,In_829);
and U346 (N_346,In_2797,In_560);
nor U347 (N_347,In_2406,In_4864);
or U348 (N_348,In_4297,In_867);
or U349 (N_349,In_96,In_2933);
nor U350 (N_350,In_4768,In_3337);
and U351 (N_351,In_2951,In_492);
xnor U352 (N_352,In_2851,In_2431);
and U353 (N_353,In_3963,In_895);
or U354 (N_354,In_3464,In_3824);
nand U355 (N_355,In_988,In_379);
nand U356 (N_356,In_4107,In_398);
and U357 (N_357,In_2110,In_2963);
nand U358 (N_358,In_361,In_639);
or U359 (N_359,In_1293,In_307);
xnor U360 (N_360,In_788,In_359);
or U361 (N_361,In_2557,In_4964);
xor U362 (N_362,In_2470,In_2604);
nor U363 (N_363,In_2265,In_757);
nand U364 (N_364,In_4777,In_1203);
and U365 (N_365,In_4556,In_1929);
or U366 (N_366,In_3149,In_330);
and U367 (N_367,In_3329,In_1326);
or U368 (N_368,In_597,In_3869);
and U369 (N_369,In_2221,In_3231);
xor U370 (N_370,In_3342,In_3755);
nor U371 (N_371,In_1912,In_938);
nand U372 (N_372,In_2079,In_4999);
nand U373 (N_373,In_610,In_608);
nand U374 (N_374,In_1371,In_3022);
or U375 (N_375,In_4057,In_4570);
nor U376 (N_376,In_2193,In_960);
nor U377 (N_377,In_3681,In_1848);
or U378 (N_378,In_871,In_3056);
xnor U379 (N_379,In_2860,In_1942);
or U380 (N_380,In_3119,In_4853);
nand U381 (N_381,In_2737,In_4499);
or U382 (N_382,In_3586,In_2185);
or U383 (N_383,In_2924,In_1337);
nand U384 (N_384,In_2102,In_2482);
and U385 (N_385,In_1905,In_2136);
xnor U386 (N_386,In_1486,In_498);
and U387 (N_387,In_768,In_4536);
or U388 (N_388,In_2244,In_1899);
xnor U389 (N_389,In_4701,In_2021);
or U390 (N_390,In_3739,In_4532);
and U391 (N_391,In_3798,In_3813);
xnor U392 (N_392,In_1403,In_2809);
xor U393 (N_393,In_2201,In_697);
and U394 (N_394,In_4524,In_1380);
nor U395 (N_395,In_2527,In_1964);
nor U396 (N_396,In_1454,In_1016);
nand U397 (N_397,In_725,In_1179);
nor U398 (N_398,In_3692,In_3592);
and U399 (N_399,In_4840,In_2188);
xor U400 (N_400,In_168,In_2050);
nor U401 (N_401,In_58,In_765);
and U402 (N_402,In_4140,In_2642);
or U403 (N_403,In_2159,In_3550);
or U404 (N_404,In_2782,In_3682);
or U405 (N_405,In_4158,In_1919);
nand U406 (N_406,In_2390,In_1839);
and U407 (N_407,In_4274,In_351);
or U408 (N_408,In_3480,In_4242);
nor U409 (N_409,In_217,In_1666);
or U410 (N_410,In_3416,In_2321);
xnor U411 (N_411,In_4617,In_4193);
nand U412 (N_412,In_2580,In_1577);
nand U413 (N_413,In_1325,In_2520);
xor U414 (N_414,In_2880,In_4269);
or U415 (N_415,In_1139,In_18);
nor U416 (N_416,In_485,In_4376);
or U417 (N_417,In_2807,In_4954);
nand U418 (N_418,In_2485,In_4231);
xor U419 (N_419,In_4075,In_3447);
xor U420 (N_420,In_3046,In_2516);
nand U421 (N_421,In_1622,In_981);
xor U422 (N_422,In_4525,In_1894);
and U423 (N_423,In_2346,In_2635);
xor U424 (N_424,In_4409,In_2123);
and U425 (N_425,In_1920,In_4011);
xnor U426 (N_426,In_3793,In_4545);
nor U427 (N_427,In_1740,In_3491);
nor U428 (N_428,In_2558,In_618);
and U429 (N_429,In_2037,In_2803);
nor U430 (N_430,In_3254,In_3315);
nand U431 (N_431,In_2893,In_2004);
xnor U432 (N_432,In_620,In_3111);
nand U433 (N_433,In_3038,In_611);
xnor U434 (N_434,In_3304,In_4822);
and U435 (N_435,In_3548,In_2007);
or U436 (N_436,In_415,In_1594);
nand U437 (N_437,In_3082,In_3906);
nand U438 (N_438,In_13,In_4559);
nor U439 (N_439,In_4762,In_510);
nand U440 (N_440,In_3128,In_2120);
xor U441 (N_441,In_954,In_4660);
and U442 (N_442,In_4048,In_1763);
nor U443 (N_443,In_4403,In_2811);
xor U444 (N_444,In_3100,In_4761);
nor U445 (N_445,In_3384,In_2502);
or U446 (N_446,In_4004,In_3504);
or U447 (N_447,In_1744,In_2047);
xnor U448 (N_448,In_3411,In_3255);
or U449 (N_449,In_3132,In_660);
xnor U450 (N_450,In_2517,In_1908);
or U451 (N_451,In_2497,In_3151);
nor U452 (N_452,In_2466,In_312);
nor U453 (N_453,In_745,In_1173);
xor U454 (N_454,In_2609,In_4105);
xnor U455 (N_455,In_2626,In_3866);
nand U456 (N_456,In_1399,In_2333);
and U457 (N_457,In_963,In_2020);
nor U458 (N_458,In_3953,In_1967);
xor U459 (N_459,In_3077,In_654);
and U460 (N_460,In_1525,In_3640);
and U461 (N_461,In_4902,In_3698);
or U462 (N_462,In_2241,In_2852);
nand U463 (N_463,In_3988,In_1805);
and U464 (N_464,In_3402,In_3458);
and U465 (N_465,In_270,In_1167);
and U466 (N_466,In_267,In_3229);
or U467 (N_467,In_912,In_2840);
or U468 (N_468,In_322,In_2366);
nor U469 (N_469,In_1364,In_1308);
xnor U470 (N_470,In_4780,In_4585);
and U471 (N_471,In_4321,In_2842);
or U472 (N_472,In_1935,In_471);
nor U473 (N_473,In_2636,In_1524);
or U474 (N_474,In_1397,In_4208);
nor U475 (N_475,In_1755,In_271);
xnor U476 (N_476,In_1765,In_2350);
xor U477 (N_477,In_889,In_2458);
and U478 (N_478,In_452,In_2947);
nand U479 (N_479,In_4101,In_332);
nor U480 (N_480,In_646,In_2688);
or U481 (N_481,In_3909,In_2414);
nor U482 (N_482,In_2978,In_1449);
or U483 (N_483,In_2144,In_3990);
nand U484 (N_484,In_2892,In_1847);
nand U485 (N_485,In_2394,In_2586);
xnor U486 (N_486,In_4582,In_2454);
nand U487 (N_487,In_715,In_1439);
xor U488 (N_488,In_591,In_4797);
nor U489 (N_489,In_3966,In_1789);
xnor U490 (N_490,In_4933,In_2504);
nand U491 (N_491,In_4377,In_4363);
xnor U492 (N_492,In_657,In_1947);
nand U493 (N_493,In_405,In_864);
nor U494 (N_494,In_2577,In_4992);
nor U495 (N_495,In_4649,In_4094);
nand U496 (N_496,In_2206,In_2198);
or U497 (N_497,In_3487,In_2012);
nand U498 (N_498,In_2114,In_540);
xor U499 (N_499,In_2067,In_3352);
nand U500 (N_500,In_2253,In_4429);
and U501 (N_501,In_1153,In_4744);
xnor U502 (N_502,In_4379,N_410);
or U503 (N_503,In_202,In_1895);
or U504 (N_504,In_1810,In_3239);
xor U505 (N_505,In_4349,N_148);
or U506 (N_506,In_3846,In_4305);
and U507 (N_507,In_1926,In_4513);
or U508 (N_508,In_4192,In_1616);
xor U509 (N_509,In_69,In_2392);
or U510 (N_510,N_355,In_2215);
or U511 (N_511,In_196,N_437);
or U512 (N_512,In_2297,In_4512);
or U513 (N_513,In_180,In_1282);
and U514 (N_514,In_4922,In_1726);
and U515 (N_515,In_1916,In_872);
nor U516 (N_516,In_640,N_13);
and U517 (N_517,In_2910,In_724);
or U518 (N_518,In_1668,In_3300);
nor U519 (N_519,In_3470,In_4620);
or U520 (N_520,In_3108,In_2959);
nor U521 (N_521,N_469,In_70);
xnor U522 (N_522,In_1567,In_2001);
or U523 (N_523,In_4441,In_3074);
and U524 (N_524,In_440,In_3576);
nand U525 (N_525,In_2961,In_106);
and U526 (N_526,In_1686,N_365);
nor U527 (N_527,In_1547,In_3912);
xnor U528 (N_528,In_350,In_999);
nand U529 (N_529,In_2478,In_878);
nor U530 (N_530,In_4165,In_125);
xor U531 (N_531,In_2890,In_4277);
nand U532 (N_532,N_307,In_2266);
nor U533 (N_533,In_4588,N_251);
xor U534 (N_534,In_857,In_4601);
nor U535 (N_535,In_284,In_1662);
xor U536 (N_536,In_1250,In_4438);
nand U537 (N_537,In_2125,In_1526);
nor U538 (N_538,In_2070,N_102);
or U539 (N_539,N_50,In_934);
nand U540 (N_540,In_3262,In_3625);
or U541 (N_541,In_2726,In_2536);
and U542 (N_542,In_2412,In_4061);
nor U543 (N_543,In_2424,N_415);
and U544 (N_544,In_2920,N_160);
and U545 (N_545,In_2593,In_807);
or U546 (N_546,In_1901,In_2710);
nand U547 (N_547,In_3968,In_2525);
or U548 (N_548,In_1862,In_3961);
nand U549 (N_549,In_139,In_3752);
nand U550 (N_550,In_3647,In_3158);
nor U551 (N_551,In_34,In_293);
nor U552 (N_552,In_4467,In_1716);
xor U553 (N_553,In_4440,N_127);
or U554 (N_554,In_1255,In_2678);
or U555 (N_555,In_317,N_280);
xor U556 (N_556,N_499,In_1981);
xnor U557 (N_557,In_389,In_3879);
and U558 (N_558,In_4145,In_2699);
xnor U559 (N_559,In_2238,In_4167);
and U560 (N_560,In_4806,In_2543);
or U561 (N_561,In_474,N_352);
and U562 (N_562,In_2884,In_483);
nor U563 (N_563,In_1033,In_784);
nand U564 (N_564,In_4261,In_2147);
nand U565 (N_565,In_1725,In_1771);
and U566 (N_566,N_240,In_3686);
or U567 (N_567,In_4160,N_400);
nand U568 (N_568,In_2663,In_292);
and U569 (N_569,In_2038,In_4932);
nand U570 (N_570,In_436,N_41);
and U571 (N_571,In_303,In_4982);
nand U572 (N_572,In_4636,In_2500);
xnor U573 (N_573,In_1979,In_3697);
nor U574 (N_574,In_3386,In_1312);
nand U575 (N_575,In_20,In_4051);
and U576 (N_576,In_913,In_943);
xor U577 (N_577,In_1887,In_253);
xor U578 (N_578,In_695,In_3214);
nor U579 (N_579,In_1295,In_3872);
nand U580 (N_580,In_537,N_125);
and U581 (N_581,N_392,In_4758);
nand U582 (N_582,In_3445,N_68);
and U583 (N_583,In_2615,In_1656);
or U584 (N_584,In_4442,In_3189);
nand U585 (N_585,N_465,In_4872);
or U586 (N_586,In_2965,In_2213);
and U587 (N_587,In_2156,In_3309);
xnor U588 (N_588,In_4655,N_198);
nor U589 (N_589,In_841,In_3924);
nor U590 (N_590,N_336,In_4607);
nor U591 (N_591,In_2930,In_1578);
nand U592 (N_592,In_1092,N_343);
nand U593 (N_593,In_3328,In_1566);
nand U594 (N_594,In_4219,In_2968);
xor U595 (N_595,In_154,In_3016);
nand U596 (N_596,In_1035,In_3354);
nor U597 (N_597,N_442,In_4168);
xor U598 (N_598,In_511,N_108);
nand U599 (N_599,In_970,In_3293);
nand U600 (N_600,In_177,In_3945);
and U601 (N_601,In_1909,In_246);
nand U602 (N_602,In_4595,In_3537);
nand U603 (N_603,In_4645,In_3762);
and U604 (N_604,N_99,N_470);
nor U605 (N_605,In_2941,In_490);
or U606 (N_606,In_2062,In_4587);
and U607 (N_607,In_3547,In_3061);
or U608 (N_608,In_744,In_2793);
xor U609 (N_609,In_4956,In_4283);
and U610 (N_610,N_463,In_2796);
nand U611 (N_611,In_4876,In_3331);
nand U612 (N_612,In_3228,In_4293);
and U613 (N_613,In_21,In_990);
xnor U614 (N_614,In_316,In_832);
or U615 (N_615,In_3363,In_694);
or U616 (N_616,In_4291,In_1627);
or U617 (N_617,In_4370,In_4514);
xnor U618 (N_618,In_4060,In_1820);
nand U619 (N_619,In_4543,In_9);
nor U620 (N_620,In_2150,In_508);
nand U621 (N_621,N_446,In_750);
nor U622 (N_622,In_781,N_385);
nor U623 (N_623,In_2197,In_2154);
and U624 (N_624,In_3510,In_4934);
or U625 (N_625,In_4019,In_4782);
xnor U626 (N_626,In_2429,In_1300);
and U627 (N_627,In_2816,In_3902);
nand U628 (N_628,In_4654,In_1675);
nor U629 (N_629,In_3024,In_2064);
nand U630 (N_630,In_1317,In_4486);
and U631 (N_631,In_1706,In_1612);
nor U632 (N_632,In_4723,In_756);
nor U633 (N_633,In_4903,In_1858);
nor U634 (N_634,In_3272,In_3059);
nor U635 (N_635,In_4421,In_3326);
nand U636 (N_636,In_718,In_3006);
nor U637 (N_637,N_178,In_2463);
and U638 (N_638,In_2957,In_3156);
nand U639 (N_639,In_242,N_211);
xnor U640 (N_640,In_2867,In_4052);
nor U641 (N_641,In_3596,In_3478);
and U642 (N_642,In_3560,In_68);
or U643 (N_643,In_2997,In_1427);
xnor U644 (N_644,N_200,In_2276);
or U645 (N_645,In_4268,In_1448);
xnor U646 (N_646,In_2711,In_1455);
or U647 (N_647,In_1541,In_2800);
and U648 (N_648,In_4692,In_3699);
nand U649 (N_649,In_3719,In_2786);
or U650 (N_650,In_1270,In_2236);
or U651 (N_651,In_2293,In_2775);
or U652 (N_652,In_4273,In_875);
and U653 (N_653,In_1005,In_507);
or U654 (N_654,In_3724,In_232);
nor U655 (N_655,In_2806,In_3670);
nor U656 (N_656,N_382,N_216);
nand U657 (N_657,In_3393,In_4665);
nor U658 (N_658,In_1520,In_3936);
or U659 (N_659,In_3193,In_4237);
xnor U660 (N_660,In_865,In_2834);
and U661 (N_661,In_1787,In_2045);
xnor U662 (N_662,In_1636,N_349);
and U663 (N_663,In_4251,In_1214);
nand U664 (N_664,In_3037,In_3410);
nor U665 (N_665,In_418,In_144);
nand U666 (N_666,N_215,In_2247);
nand U667 (N_667,In_301,In_3536);
and U668 (N_668,In_3955,In_3649);
xor U669 (N_669,In_3620,In_4646);
or U670 (N_670,In_2977,In_3028);
nor U671 (N_671,In_2148,N_152);
xor U672 (N_672,In_2943,In_4255);
nand U673 (N_673,In_1263,In_308);
xor U674 (N_674,In_3965,In_497);
and U675 (N_675,In_3502,In_3831);
nand U676 (N_676,In_1112,In_4473);
nand U677 (N_677,In_487,In_3283);
or U678 (N_678,In_2324,In_817);
nand U679 (N_679,N_58,In_520);
and U680 (N_680,In_3712,In_229);
nor U681 (N_681,In_3668,In_3383);
nor U682 (N_682,In_4878,In_2984);
xor U683 (N_683,In_1334,In_910);
and U684 (N_684,In_2722,In_2451);
and U685 (N_685,N_11,N_187);
nand U686 (N_686,N_320,In_3197);
nor U687 (N_687,In_4346,In_336);
xnor U688 (N_688,In_1512,In_362);
xor U689 (N_689,In_1834,In_4968);
nor U690 (N_690,In_3372,In_3705);
and U691 (N_691,In_2450,In_2436);
nand U692 (N_692,In_2243,In_2998);
or U693 (N_693,In_522,In_2578);
or U694 (N_694,In_33,In_155);
xor U695 (N_695,N_386,In_4352);
and U696 (N_696,In_2338,N_139);
or U697 (N_697,N_308,In_348);
nand U698 (N_698,In_4450,In_683);
nand U699 (N_699,In_4610,In_4747);
xor U700 (N_700,In_1792,In_4630);
xor U701 (N_701,In_4220,In_1853);
xor U702 (N_702,In_933,In_4162);
or U703 (N_703,N_235,In_716);
and U704 (N_704,In_2315,In_1278);
xnor U705 (N_705,In_3650,In_3679);
or U706 (N_706,In_1871,In_4389);
xor U707 (N_707,In_1835,In_3369);
xnor U708 (N_708,In_4984,N_483);
nand U709 (N_709,In_1985,In_3901);
nand U710 (N_710,In_205,In_4065);
nor U711 (N_711,In_4684,In_1468);
xor U712 (N_712,N_107,In_189);
or U713 (N_713,In_2617,In_539);
and U714 (N_714,In_1410,In_2562);
nand U715 (N_715,In_1910,In_1336);
xor U716 (N_716,In_4388,In_3176);
nand U717 (N_717,In_899,In_3958);
and U718 (N_718,In_3391,In_769);
or U719 (N_719,In_4153,In_3678);
and U720 (N_720,In_1077,In_5);
xor U721 (N_721,In_4150,In_4034);
or U722 (N_722,In_1274,In_2808);
nand U723 (N_723,In_3566,In_2798);
nor U724 (N_724,In_3660,In_1260);
nand U725 (N_725,N_217,N_76);
and U726 (N_726,In_842,N_273);
and U727 (N_727,In_2052,In_1718);
nand U728 (N_728,In_2781,In_2189);
and U729 (N_729,In_17,In_185);
nand U730 (N_730,In_2850,In_4082);
xor U731 (N_731,In_2440,N_298);
nand U732 (N_732,In_2036,N_486);
xor U733 (N_733,In_2091,N_135);
and U734 (N_734,In_3746,In_944);
xnor U735 (N_735,In_2113,In_4213);
or U736 (N_736,In_1121,In_368);
nand U737 (N_737,In_3422,In_3282);
and U738 (N_738,In_2426,N_69);
xnor U739 (N_739,In_1648,In_1536);
and U740 (N_740,In_1398,In_163);
or U741 (N_741,In_2669,In_1054);
nor U742 (N_742,In_689,In_4764);
nor U743 (N_743,In_31,N_12);
xnor U744 (N_744,In_3121,In_2513);
or U745 (N_745,In_328,In_3085);
xnor U746 (N_746,In_4036,In_650);
nor U747 (N_747,In_3927,In_4583);
xnor U748 (N_748,N_19,In_133);
and U749 (N_749,N_250,N_263);
nor U750 (N_750,In_3604,In_161);
xnor U751 (N_751,In_1257,In_2178);
xor U752 (N_752,In_4225,N_15);
xnor U753 (N_753,In_201,In_182);
or U754 (N_754,In_2207,In_255);
or U755 (N_755,In_1192,N_232);
or U756 (N_756,In_1421,N_458);
xor U757 (N_757,In_326,In_1392);
nand U758 (N_758,In_1409,In_2279);
xor U759 (N_759,In_582,In_2326);
or U760 (N_760,In_753,N_218);
and U761 (N_761,In_1933,In_3675);
nor U762 (N_762,In_2420,In_2065);
xnor U763 (N_763,N_321,In_2944);
or U764 (N_764,In_786,In_1602);
and U765 (N_765,In_1297,In_1994);
or U766 (N_766,In_424,N_192);
or U767 (N_767,In_2802,N_480);
nor U768 (N_768,N_72,In_1938);
and U769 (N_769,N_390,In_3303);
nand U770 (N_770,In_3568,In_3023);
and U771 (N_771,In_3081,In_1495);
nor U772 (N_772,In_592,In_3995);
nor U773 (N_773,In_2625,In_1304);
and U774 (N_774,N_103,In_2643);
and U775 (N_775,In_1562,N_360);
or U776 (N_776,N_177,In_1955);
or U777 (N_777,In_1813,In_3919);
or U778 (N_778,In_425,N_478);
nand U779 (N_779,In_4449,N_384);
and U780 (N_780,In_3726,N_453);
and U781 (N_781,In_4592,In_3459);
xor U782 (N_782,In_3765,In_2603);
xor U783 (N_783,In_1425,In_3031);
or U784 (N_784,In_732,In_4817);
nand U785 (N_785,In_325,In_4426);
xnor U786 (N_786,In_2170,In_2368);
or U787 (N_787,In_3760,N_406);
or U788 (N_788,In_4750,In_3093);
nand U789 (N_789,N_471,N_98);
and U790 (N_790,In_2381,In_3453);
and U791 (N_791,In_849,In_4740);
nand U792 (N_792,N_140,In_4281);
or U793 (N_793,N_33,In_586);
or U794 (N_794,In_4087,In_688);
nand U795 (N_795,In_4195,N_132);
and U796 (N_796,In_63,In_1185);
nor U797 (N_797,In_3075,In_324);
nand U798 (N_798,In_1888,In_785);
or U799 (N_799,In_818,In_1098);
nand U800 (N_800,In_2768,In_4367);
and U801 (N_801,In_672,In_3115);
xnor U802 (N_802,In_734,In_1224);
xnor U803 (N_803,In_135,In_4975);
nand U804 (N_804,In_4411,In_2799);
and U805 (N_805,In_1931,In_2877);
and U806 (N_806,In_1288,In_3941);
nand U807 (N_807,In_891,N_242);
and U808 (N_808,In_3665,In_1886);
nor U809 (N_809,In_706,In_1138);
nor U810 (N_810,In_4177,In_2847);
xnor U811 (N_811,In_4093,In_3875);
nor U812 (N_812,In_2563,In_4912);
nor U813 (N_813,In_2275,In_4694);
nor U814 (N_814,In_3769,In_2763);
or U815 (N_815,In_504,In_2876);
nand U816 (N_816,N_179,In_1096);
and U817 (N_817,In_993,In_3767);
xnor U818 (N_818,In_421,In_2343);
nand U819 (N_819,In_1712,In_1230);
or U820 (N_820,In_448,In_3960);
nor U821 (N_821,In_3704,In_2328);
nand U822 (N_822,In_4205,In_4516);
and U823 (N_823,In_4502,In_930);
and U824 (N_824,In_387,In_1533);
nand U825 (N_825,In_4584,In_269);
nor U826 (N_826,In_3232,In_462);
nand U827 (N_827,In_3513,In_530);
and U828 (N_828,In_4970,In_1062);
xnor U829 (N_829,In_2090,In_3782);
nor U830 (N_830,In_791,In_339);
and U831 (N_831,In_564,In_3408);
nand U832 (N_832,N_121,In_2732);
xnor U833 (N_833,In_3226,In_4682);
and U834 (N_834,In_984,In_2181);
xor U835 (N_835,In_3148,In_856);
nand U836 (N_836,N_327,In_1631);
and U837 (N_837,In_3,In_3808);
nand U838 (N_838,In_641,In_1701);
xnor U839 (N_839,N_202,In_521);
nor U840 (N_840,In_1814,In_4977);
nand U841 (N_841,In_2532,In_1280);
or U842 (N_842,In_4508,In_4766);
or U843 (N_843,In_1189,In_213);
nand U844 (N_844,In_4138,In_853);
xnor U845 (N_845,In_265,In_4457);
xnor U846 (N_846,In_3663,N_275);
nand U847 (N_847,In_3711,In_3299);
xor U848 (N_848,In_3207,In_150);
or U849 (N_849,In_3010,In_1063);
or U850 (N_850,In_4691,N_244);
and U851 (N_851,In_2019,In_2033);
xor U852 (N_852,In_408,In_4551);
and U853 (N_853,In_771,In_74);
xor U854 (N_854,In_995,In_1148);
and U855 (N_855,In_3994,In_1830);
or U856 (N_856,In_2791,In_2662);
and U857 (N_857,In_2638,In_1051);
nor U858 (N_858,In_3599,In_1265);
xor U859 (N_859,In_1119,In_1402);
or U860 (N_860,N_4,In_2762);
nand U861 (N_861,In_3653,N_447);
nor U862 (N_862,In_430,In_4275);
nand U863 (N_863,N_78,In_4055);
nand U864 (N_864,In_4196,N_247);
and U865 (N_865,In_1754,In_48);
or U866 (N_866,In_4172,N_52);
nand U867 (N_867,In_4675,In_481);
nand U868 (N_868,In_2100,N_201);
or U869 (N_869,In_4972,In_3018);
or U870 (N_870,In_2813,In_129);
or U871 (N_871,In_4373,In_1070);
nand U872 (N_872,In_3281,In_2522);
or U873 (N_873,In_1496,In_3014);
nor U874 (N_874,N_490,In_636);
xor U875 (N_875,In_2528,In_3253);
or U876 (N_876,In_3672,In_3052);
xnor U877 (N_877,In_2647,In_4307);
nor U878 (N_878,In_1809,In_195);
and U879 (N_879,In_3611,N_42);
xor U880 (N_880,In_1676,In_3092);
and U881 (N_881,In_4711,In_2911);
xor U882 (N_882,In_4616,In_3216);
or U883 (N_883,In_4869,In_4571);
or U884 (N_884,In_2882,In_2929);
and U885 (N_885,In_3881,In_2372);
or U886 (N_886,In_2896,In_385);
or U887 (N_887,In_2230,In_1095);
nor U888 (N_888,In_3147,In_675);
nand U889 (N_889,In_1418,In_2063);
nor U890 (N_890,In_3020,In_4000);
or U891 (N_891,In_840,In_3090);
nand U892 (N_892,In_1990,In_3483);
and U893 (N_893,In_3250,In_395);
nor U894 (N_894,In_4611,In_160);
or U895 (N_895,In_370,In_423);
nand U896 (N_896,In_3648,In_4241);
or U897 (N_897,In_2731,In_4492);
xnor U898 (N_898,In_3336,In_331);
xor U899 (N_899,N_122,In_2550);
and U900 (N_900,In_2237,In_1438);
xnor U901 (N_901,In_3779,In_941);
nor U902 (N_902,In_4127,In_2183);
xor U903 (N_903,In_4546,In_927);
nor U904 (N_904,In_2404,In_76);
nor U905 (N_905,In_923,N_57);
or U906 (N_906,In_3691,In_833);
or U907 (N_907,In_239,In_469);
nor U908 (N_908,In_3748,In_2862);
nor U909 (N_909,In_1618,In_588);
nand U910 (N_910,In_2831,In_2660);
nor U911 (N_911,In_2255,N_319);
and U912 (N_912,In_1854,In_2382);
nand U913 (N_913,In_3515,In_3220);
or U914 (N_914,In_1692,In_4936);
xnor U915 (N_915,N_449,In_2837);
nand U916 (N_916,In_60,In_2991);
and U917 (N_917,In_4248,In_2632);
xnor U918 (N_918,In_4415,In_4126);
xnor U919 (N_919,N_427,In_4194);
xor U920 (N_920,In_3530,In_2263);
nor U921 (N_921,In_4604,N_133);
nand U922 (N_922,In_4715,In_1494);
nand U923 (N_923,In_3501,In_309);
and U924 (N_924,In_4270,In_3934);
nand U925 (N_925,In_2724,In_4865);
xnor U926 (N_926,In_2089,In_543);
nand U927 (N_927,In_1683,In_112);
or U928 (N_928,In_147,In_3305);
nand U929 (N_929,In_4778,In_4785);
and U930 (N_930,In_3364,In_447);
xor U931 (N_931,In_2841,In_2529);
nand U932 (N_932,In_57,In_2833);
or U933 (N_933,N_35,In_4318);
and U934 (N_934,In_333,In_4132);
and U935 (N_935,In_986,In_1806);
or U936 (N_936,In_1161,In_4830);
nor U937 (N_937,In_109,In_1610);
nand U938 (N_938,In_2974,In_3932);
nand U939 (N_939,N_82,In_3612);
xnor U940 (N_940,N_191,In_1306);
nor U941 (N_941,N_197,In_1239);
or U942 (N_942,In_3578,In_3969);
nand U943 (N_943,In_4074,In_2646);
and U944 (N_944,In_4974,In_1499);
xnor U945 (N_945,In_2311,In_1780);
or U946 (N_946,N_322,In_1245);
or U947 (N_947,In_3573,In_4888);
nor U948 (N_948,N_452,In_2481);
xnor U949 (N_949,In_848,In_3145);
and U950 (N_950,In_859,In_831);
and U951 (N_951,In_4889,In_2445);
or U952 (N_952,In_3170,In_4509);
nand U953 (N_953,In_2843,In_936);
xnor U954 (N_954,In_1614,In_1930);
and U955 (N_955,In_2418,In_569);
xnor U956 (N_956,In_1386,In_1345);
nor U957 (N_957,N_450,In_1435);
nand U958 (N_958,In_3320,In_2168);
xnor U959 (N_959,N_411,In_4215);
xor U960 (N_960,In_4818,In_4941);
xor U961 (N_961,In_1053,In_4200);
xnor U962 (N_962,In_544,In_4427);
nand U963 (N_963,In_2245,In_1368);
nor U964 (N_964,In_1655,In_3680);
nor U965 (N_965,In_4729,In_4915);
xnor U966 (N_966,In_1424,In_3512);
or U967 (N_967,In_4385,In_3153);
xor U968 (N_968,In_4568,In_3130);
xor U969 (N_969,In_4279,In_381);
nor U970 (N_970,In_1896,N_93);
and U971 (N_971,In_3891,In_4779);
xnor U972 (N_972,In_2353,In_345);
nor U973 (N_973,In_668,In_3828);
nand U974 (N_974,In_3701,In_2130);
and U975 (N_975,In_2939,In_4662);
or U976 (N_976,In_1590,In_2599);
nand U977 (N_977,In_2142,In_2348);
or U978 (N_978,In_4399,N_224);
xor U979 (N_979,N_315,In_4384);
and U980 (N_980,In_4312,In_164);
or U981 (N_981,In_457,N_402);
nand U982 (N_982,In_2783,N_231);
or U983 (N_983,In_1333,In_343);
or U984 (N_984,In_3983,In_3727);
nand U985 (N_985,In_1171,In_1551);
nand U986 (N_986,In_2339,In_3224);
and U987 (N_987,In_461,In_533);
xnor U988 (N_988,In_3747,In_1774);
or U989 (N_989,In_2671,In_1660);
or U990 (N_990,In_1390,In_1978);
or U991 (N_991,In_1791,In_2483);
or U992 (N_992,N_141,In_1501);
and U993 (N_993,In_4223,In_4731);
xor U994 (N_994,In_1383,In_50);
xnor U995 (N_995,In_110,In_740);
nand U996 (N_996,In_4487,In_3343);
nor U997 (N_997,In_1,In_2854);
nor U998 (N_998,In_4955,In_772);
nor U999 (N_999,In_4342,In_4383);
nand U1000 (N_1000,N_377,In_3778);
xnor U1001 (N_1001,In_2486,In_3042);
nor U1002 (N_1002,In_1673,In_4324);
xnor U1003 (N_1003,In_2787,N_637);
xor U1004 (N_1004,In_4651,In_3030);
nor U1005 (N_1005,N_36,In_2292);
and U1006 (N_1006,In_3120,N_701);
or U1007 (N_1007,In_3661,In_123);
and U1008 (N_1008,In_411,In_215);
nor U1009 (N_1009,In_604,In_1678);
nand U1010 (N_1010,In_1174,In_2966);
nand U1011 (N_1011,In_197,In_156);
nor U1012 (N_1012,In_1825,In_2162);
xnor U1013 (N_1013,In_956,In_2472);
nor U1014 (N_1014,In_642,N_435);
nor U1015 (N_1015,In_2475,N_376);
and U1016 (N_1016,N_354,In_1841);
xnor U1017 (N_1017,N_947,N_451);
or U1018 (N_1018,N_119,In_3438);
nand U1019 (N_1019,N_500,In_3263);
nand U1020 (N_1020,In_2745,In_1988);
or U1021 (N_1021,In_1703,In_1574);
nand U1022 (N_1022,In_3567,N_306);
nor U1023 (N_1023,In_4103,In_1175);
or U1024 (N_1024,In_4677,In_1481);
or U1025 (N_1025,In_2601,In_880);
nand U1026 (N_1026,In_1952,In_581);
nor U1027 (N_1027,In_3066,In_2398);
nor U1028 (N_1028,In_4362,In_4405);
or U1029 (N_1029,In_1115,In_1320);
nand U1030 (N_1030,In_3632,In_124);
nor U1031 (N_1031,In_3289,In_412);
xor U1032 (N_1032,N_927,In_529);
nand U1033 (N_1033,In_3154,In_2388);
nand U1034 (N_1034,In_1107,In_2931);
nand U1035 (N_1035,In_2559,In_4573);
nand U1036 (N_1036,In_1184,In_1071);
xor U1037 (N_1037,In_2597,In_3291);
nor U1038 (N_1038,In_3826,In_2452);
and U1039 (N_1039,In_233,In_1560);
xor U1040 (N_1040,In_625,In_834);
and U1041 (N_1041,In_4466,In_4752);
xnor U1042 (N_1042,N_432,In_7);
xnor U1043 (N_1043,In_4263,In_1544);
xor U1044 (N_1044,N_543,In_3067);
nand U1045 (N_1045,In_1623,In_2973);
and U1046 (N_1046,N_889,N_757);
and U1047 (N_1047,In_2003,In_1635);
and U1048 (N_1048,N_799,In_687);
and U1049 (N_1049,In_4988,In_4918);
or U1050 (N_1050,In_2488,In_10);
xnor U1051 (N_1051,In_3835,In_4228);
nor U1052 (N_1052,N_467,In_2042);
or U1053 (N_1053,In_851,N_174);
or U1054 (N_1054,In_1289,N_531);
and U1055 (N_1055,N_312,In_4031);
xor U1056 (N_1056,In_4445,N_128);
xor U1057 (N_1057,N_43,In_2161);
nor U1058 (N_1058,In_903,In_3987);
nor U1059 (N_1059,In_4996,In_2764);
xor U1060 (N_1060,In_2071,N_567);
and U1061 (N_1061,In_1379,In_3896);
nor U1062 (N_1062,In_2948,In_953);
xor U1063 (N_1063,In_2217,N_112);
nor U1064 (N_1064,In_2868,In_335);
and U1065 (N_1065,In_4852,N_137);
nor U1066 (N_1066,In_438,In_1322);
and U1067 (N_1067,N_115,N_861);
nand U1068 (N_1068,In_1821,In_3997);
nand U1069 (N_1069,In_4098,In_4973);
and U1070 (N_1070,In_509,In_3677);
nand U1071 (N_1071,N_585,N_425);
nor U1072 (N_1072,In_1657,N_464);
xnor U1073 (N_1073,In_1111,In_3495);
nor U1074 (N_1074,In_925,N_755);
nor U1075 (N_1075,In_3353,In_2922);
or U1076 (N_1076,In_783,In_3488);
and U1077 (N_1077,In_2622,In_2299);
or U1078 (N_1078,N_943,In_46);
or U1079 (N_1079,In_1849,In_3703);
xnor U1080 (N_1080,N_763,In_3298);
xor U1081 (N_1081,In_329,In_2487);
xor U1082 (N_1082,In_3904,N_820);
and U1083 (N_1083,In_3317,In_4470);
nand U1084 (N_1084,N_840,In_3169);
nor U1085 (N_1085,In_1474,In_3605);
or U1086 (N_1086,N_980,In_662);
nor U1087 (N_1087,In_4316,In_248);
or U1088 (N_1088,N_195,N_593);
xor U1089 (N_1089,In_2666,In_4603);
and U1090 (N_1090,N_587,In_1677);
xnor U1091 (N_1091,In_4689,In_3802);
or U1092 (N_1092,In_3243,In_2918);
nand U1093 (N_1093,In_4125,In_3644);
nand U1094 (N_1094,N_512,N_316);
or U1095 (N_1095,In_3552,In_602);
xnor U1096 (N_1096,In_4981,N_105);
or U1097 (N_1097,In_1599,In_1530);
xnor U1098 (N_1098,In_3544,In_93);
nor U1099 (N_1099,In_1441,In_2832);
nand U1100 (N_1100,N_241,In_334);
and U1101 (N_1101,N_668,In_4754);
or U1102 (N_1102,In_85,In_4529);
nor U1103 (N_1103,In_107,In_1653);
nor U1104 (N_1104,N_163,In_4631);
and U1105 (N_1105,N_649,In_1369);
nand U1106 (N_1106,In_4624,In_4217);
and U1107 (N_1107,In_3429,In_2129);
xnor U1108 (N_1108,In_2667,In_1876);
xor U1109 (N_1109,In_1010,In_1459);
xor U1110 (N_1110,In_916,N_887);
and U1111 (N_1111,In_3992,N_487);
nand U1112 (N_1112,In_250,In_4963);
xnor U1113 (N_1113,In_273,N_827);
and U1114 (N_1114,In_2257,In_2919);
xor U1115 (N_1115,In_1845,N_375);
or U1116 (N_1116,In_3181,In_4608);
or U1117 (N_1117,In_991,In_612);
nor U1118 (N_1118,N_295,In_1048);
nand U1119 (N_1119,In_3089,In_3083);
or U1120 (N_1120,In_2595,N_955);
nand U1121 (N_1121,N_89,N_313);
xnor U1122 (N_1122,In_4945,In_2231);
or U1123 (N_1123,In_2715,In_3959);
and U1124 (N_1124,In_2008,In_394);
nor U1125 (N_1125,In_4387,In_2403);
nor U1126 (N_1126,In_223,In_2367);
nand U1127 (N_1127,In_3385,In_3771);
nand U1128 (N_1128,In_3123,In_1046);
nand U1129 (N_1129,In_2152,In_1022);
nor U1130 (N_1130,In_3607,In_4829);
nor U1131 (N_1131,In_974,In_2387);
and U1132 (N_1132,In_2583,In_372);
nor U1133 (N_1133,In_262,N_468);
nand U1134 (N_1134,In_4985,N_911);
and U1135 (N_1135,N_888,In_4290);
xor U1136 (N_1136,In_2460,In_3199);
nand U1137 (N_1137,In_4439,In_2661);
xnor U1138 (N_1138,In_3619,In_3129);
nor U1139 (N_1139,In_3683,In_404);
or U1140 (N_1140,N_779,In_4076);
xor U1141 (N_1141,In_2040,In_3815);
nand U1142 (N_1142,In_762,In_3425);
nor U1143 (N_1143,In_1412,N_371);
and U1144 (N_1144,In_2554,In_616);
nand U1145 (N_1145,In_1689,In_4380);
and U1146 (N_1146,In_1878,N_285);
and U1147 (N_1147,In_2714,In_2222);
or U1148 (N_1148,In_2300,N_359);
xor U1149 (N_1149,In_806,In_3736);
xnor U1150 (N_1150,In_3790,In_2296);
or U1151 (N_1151,N_445,In_1490);
nor U1152 (N_1152,In_2119,In_4831);
and U1153 (N_1153,In_3414,In_1940);
nand U1154 (N_1154,In_2043,In_820);
xor U1155 (N_1155,In_561,In_1426);
xnor U1156 (N_1156,In_3643,In_1609);
nand U1157 (N_1157,In_3570,In_4669);
xor U1158 (N_1158,In_4746,In_1355);
or U1159 (N_1159,N_170,In_1811);
nand U1160 (N_1160,In_2702,In_1993);
xor U1161 (N_1161,In_1472,In_146);
nand U1162 (N_1162,In_1595,In_1272);
or U1163 (N_1163,N_809,N_940);
and U1164 (N_1164,In_3800,In_3003);
xnor U1165 (N_1165,In_722,In_2570);
or U1166 (N_1166,In_4726,N_616);
xnor U1167 (N_1167,In_4135,In_1170);
xnor U1168 (N_1168,N_95,In_2640);
or U1169 (N_1169,N_856,In_2909);
and U1170 (N_1170,In_2083,In_1946);
and U1171 (N_1171,In_617,In_563);
or U1172 (N_1172,N_873,N_533);
nand U1173 (N_1173,In_870,In_3606);
and U1174 (N_1174,In_298,In_1889);
and U1175 (N_1175,In_2568,In_87);
nand U1176 (N_1176,N_395,N_822);
or U1177 (N_1177,N_847,N_104);
or U1178 (N_1178,In_2612,In_3359);
xnor U1179 (N_1179,In_812,In_1572);
nor U1180 (N_1180,N_325,In_3858);
and U1181 (N_1181,In_2449,In_495);
nand U1182 (N_1182,In_417,In_4078);
nor U1183 (N_1183,N_248,In_670);
and U1184 (N_1184,In_4629,In_822);
and U1185 (N_1185,In_4755,N_773);
xnor U1186 (N_1186,In_1881,N_941);
nor U1187 (N_1187,In_167,In_4504);
or U1188 (N_1188,In_4605,In_2906);
xor U1189 (N_1189,In_1687,In_4109);
or U1190 (N_1190,In_3768,In_3783);
nand U1191 (N_1191,N_964,N_816);
and U1192 (N_1192,In_3310,In_3171);
nor U1193 (N_1193,In_2789,In_4609);
xor U1194 (N_1194,In_1757,N_430);
and U1195 (N_1195,In_1516,N_419);
or U1196 (N_1196,In_3636,In_3925);
or U1197 (N_1197,In_4171,In_1785);
nor U1198 (N_1198,In_550,In_2748);
nor U1199 (N_1199,In_4895,In_972);
nor U1200 (N_1200,In_823,In_3177);
xor U1201 (N_1201,N_573,In_3376);
or U1202 (N_1202,In_3456,In_2421);
xnor U1203 (N_1203,In_2689,In_587);
nor U1204 (N_1204,In_4453,In_3109);
nand U1205 (N_1205,N_348,In_2844);
nand U1206 (N_1206,In_4247,In_128);
and U1207 (N_1207,N_695,In_1702);
or U1208 (N_1208,In_558,In_2881);
nor U1209 (N_1209,In_518,In_2115);
nand U1210 (N_1210,In_1605,In_1081);
or U1211 (N_1211,In_580,In_557);
or U1212 (N_1212,In_2627,N_874);
nand U1213 (N_1213,In_2921,In_755);
or U1214 (N_1214,In_432,In_1242);
xnor U1215 (N_1215,In_2537,In_296);
or U1216 (N_1216,In_159,N_175);
nor U1217 (N_1217,In_2937,In_3907);
and U1218 (N_1218,In_3637,In_4882);
or U1219 (N_1219,In_801,In_238);
xor U1220 (N_1220,In_1617,In_4410);
or U1221 (N_1221,In_1332,In_302);
xor U1222 (N_1222,In_1457,N_639);
or U1223 (N_1223,In_1709,In_235);
and U1224 (N_1224,In_2725,In_1025);
xnor U1225 (N_1225,In_713,In_1851);
and U1226 (N_1226,N_675,N_56);
or U1227 (N_1227,N_783,In_466);
nor U1228 (N_1228,In_3078,N_586);
nand U1229 (N_1229,In_4046,In_2817);
nor U1230 (N_1230,In_4343,In_199);
xnor U1231 (N_1231,In_4858,In_2600);
xnor U1232 (N_1232,In_4267,In_2072);
or U1233 (N_1233,In_2735,In_1720);
nand U1234 (N_1234,N_672,N_302);
nor U1235 (N_1235,In_1873,In_3230);
or U1236 (N_1236,N_142,In_1432);
xnor U1237 (N_1237,In_2087,N_992);
nand U1238 (N_1238,In_2582,In_4501);
nand U1239 (N_1239,In_2619,N_841);
nor U1240 (N_1240,In_746,In_4458);
nand U1241 (N_1241,In_95,In_3913);
xnor U1242 (N_1242,In_4212,N_190);
and U1243 (N_1243,In_3486,In_4693);
or U1244 (N_1244,In_3057,In_3622);
xor U1245 (N_1245,In_3379,In_3593);
nand U1246 (N_1246,In_4809,In_3843);
or U1247 (N_1247,N_387,In_2812);
nand U1248 (N_1248,In_3734,In_1356);
nand U1249 (N_1249,In_2018,In_1205);
and U1250 (N_1250,N_996,N_618);
nand U1251 (N_1251,N_818,In_664);
and U1252 (N_1252,In_1596,In_2365);
nor U1253 (N_1253,In_4149,In_4351);
or U1254 (N_1254,In_1210,In_1328);
xor U1255 (N_1255,In_545,In_2972);
and U1256 (N_1256,In_4243,In_1731);
or U1257 (N_1257,In_1440,In_3273);
or U1258 (N_1258,In_2810,N_461);
and U1259 (N_1259,In_1400,In_342);
and U1260 (N_1260,In_861,N_689);
xnor U1261 (N_1261,In_2926,In_1018);
nor U1262 (N_1262,In_2530,N_10);
nor U1263 (N_1263,In_2508,N_548);
nand U1264 (N_1264,In_2608,In_1555);
and U1265 (N_1265,In_3993,In_4432);
xor U1266 (N_1266,N_872,In_946);
nand U1267 (N_1267,In_1463,N_860);
nand U1268 (N_1268,N_345,In_1852);
nand U1269 (N_1269,In_254,In_1504);
nor U1270 (N_1270,N_920,N_46);
and U1271 (N_1271,In_1698,N_852);
xnor U1272 (N_1272,In_3294,In_3375);
nand U1273 (N_1273,In_4983,In_3071);
xnor U1274 (N_1274,N_267,In_3460);
xnor U1275 (N_1275,N_394,N_364);
nor U1276 (N_1276,In_400,In_1951);
and U1277 (N_1277,In_4712,In_975);
nand U1278 (N_1278,In_2401,In_1961);
and U1279 (N_1279,In_1433,In_1183);
nand U1280 (N_1280,In_2268,In_1482);
or U1281 (N_1281,In_4480,In_4207);
xnor U1282 (N_1282,In_1882,In_542);
nor U1283 (N_1283,In_431,In_3837);
nand U1284 (N_1284,In_1913,In_1286);
xor U1285 (N_1285,In_3851,In_3914);
nand U1286 (N_1286,In_1783,In_4561);
nor U1287 (N_1287,In_3525,N_971);
or U1288 (N_1288,In_256,In_1262);
and U1289 (N_1289,In_2055,In_1922);
nor U1290 (N_1290,In_4419,In_1695);
nand U1291 (N_1291,N_481,In_3076);
xor U1292 (N_1292,In_65,In_3346);
or U1293 (N_1293,In_4159,In_3219);
nand U1294 (N_1294,In_907,In_1103);
xor U1295 (N_1295,In_4091,N_696);
nor U1296 (N_1296,In_4117,In_12);
nand U1297 (N_1297,N_351,N_994);
nor U1298 (N_1298,In_1385,In_2753);
nand U1299 (N_1299,In_4469,In_1039);
nand U1300 (N_1300,In_3582,In_3839);
or U1301 (N_1301,In_1764,In_3338);
xnor U1302 (N_1302,In_137,In_321);
and U1303 (N_1303,In_4119,In_4563);
and U1304 (N_1304,In_4835,In_1091);
nand U1305 (N_1305,In_499,In_1015);
and U1306 (N_1306,In_2218,N_663);
and U1307 (N_1307,In_2564,In_1630);
nand U1308 (N_1308,In_3922,In_3749);
and U1309 (N_1309,In_4069,In_3476);
nor U1310 (N_1310,In_3449,In_4850);
nand U1311 (N_1311,In_1450,In_2576);
nor U1312 (N_1312,In_3103,In_4006);
nand U1313 (N_1313,N_381,In_171);
xor U1314 (N_1314,In_4039,In_4648);
nand U1315 (N_1315,In_2208,In_4054);
nand U1316 (N_1316,In_4827,In_3097);
nor U1317 (N_1317,N_727,In_1597);
and U1318 (N_1318,In_3916,In_4614);
xnor U1319 (N_1319,N_876,N_230);
nand U1320 (N_1320,N_969,In_3378);
or U1321 (N_1321,In_2226,In_819);
nand U1322 (N_1322,In_1891,In_1911);
nand U1323 (N_1323,In_2347,In_4003);
or U1324 (N_1324,In_1611,N_362);
nand U1325 (N_1325,In_2204,In_1941);
xor U1326 (N_1326,In_2889,N_899);
xnor U1327 (N_1327,In_3054,N_808);
or U1328 (N_1328,In_3985,In_1640);
nand U1329 (N_1329,In_2175,In_1545);
nand U1330 (N_1330,N_652,In_961);
nor U1331 (N_1331,In_1047,In_531);
xor U1332 (N_1332,In_4794,In_4246);
or U1333 (N_1333,In_1788,In_3522);
and U1334 (N_1334,In_4976,In_3178);
nand U1335 (N_1335,N_55,In_4947);
or U1336 (N_1336,In_3855,In_1136);
nand U1337 (N_1337,In_1690,In_98);
or U1338 (N_1338,In_1004,In_3473);
or U1339 (N_1339,In_606,N_725);
xor U1340 (N_1340,In_3218,In_204);
and U1341 (N_1341,N_832,In_4452);
nor U1342 (N_1342,In_4926,In_2655);
and U1343 (N_1343,In_2447,In_4576);
or U1344 (N_1344,In_1349,In_353);
or U1345 (N_1345,In_2495,In_4547);
or U1346 (N_1346,In_4064,In_2886);
xor U1347 (N_1347,In_2301,In_2046);
or U1348 (N_1348,In_468,In_3761);
or U1349 (N_1349,In_4733,In_1581);
and U1350 (N_1350,N_712,N_491);
xnor U1351 (N_1351,In_1067,In_2186);
or U1352 (N_1352,In_838,In_4079);
xor U1353 (N_1353,In_4891,In_1739);
nand U1354 (N_1354,In_2438,In_4108);
nor U1355 (N_1355,In_4635,In_2584);
nand U1356 (N_1356,In_2544,In_3796);
nor U1357 (N_1357,In_1833,In_4931);
or U1358 (N_1358,In_4897,In_2682);
and U1359 (N_1359,N_781,N_117);
and U1360 (N_1360,In_4086,In_3365);
xor U1361 (N_1361,N_156,In_4625);
nand U1362 (N_1362,In_4930,In_998);
nand U1363 (N_1363,N_823,In_378);
nor U1364 (N_1364,In_1040,In_2848);
nand U1365 (N_1365,N_690,In_4686);
or U1366 (N_1366,N_330,In_4674);
nand U1367 (N_1367,In_4676,In_3118);
and U1368 (N_1368,In_4841,In_49);
and U1369 (N_1369,In_2980,In_661);
nor U1370 (N_1370,In_3443,N_628);
nor U1371 (N_1371,N_311,In_1154);
nor U1372 (N_1372,In_2228,N_525);
nor U1373 (N_1373,N_342,In_1244);
or U1374 (N_1374,In_3689,In_2746);
nand U1375 (N_1375,N_598,In_4044);
or U1376 (N_1376,In_1431,In_2165);
xnor U1377 (N_1377,N_811,In_3903);
nor U1378 (N_1378,N_868,In_4541);
xor U1379 (N_1379,In_3058,N_335);
or U1380 (N_1380,In_1613,N_106);
or U1381 (N_1381,In_4900,In_2419);
xor U1382 (N_1382,In_3818,In_1794);
nand U1383 (N_1383,In_162,In_4375);
xor U1384 (N_1384,N_333,In_356);
and U1385 (N_1385,N_94,In_4310);
nand U1386 (N_1386,In_2879,In_4099);
and U1387 (N_1387,In_4018,N_388);
nand U1388 (N_1388,In_4538,In_2822);
and U1389 (N_1389,In_3288,In_1128);
or U1390 (N_1390,In_2891,In_1506);
nand U1391 (N_1391,In_787,N_838);
nand U1392 (N_1392,In_4837,In_4084);
and U1393 (N_1393,In_2838,In_1767);
xor U1394 (N_1394,In_948,In_1158);
or U1395 (N_1395,In_2396,N_765);
and U1396 (N_1396,In_2987,In_3412);
xor U1397 (N_1397,In_1893,N_27);
nor U1398 (N_1398,In_1200,In_3722);
xor U1399 (N_1399,In_4201,In_4191);
and U1400 (N_1400,N_750,N_953);
xnor U1401 (N_1401,In_1639,In_2870);
and U1402 (N_1402,In_3138,In_473);
nand U1403 (N_1403,In_845,In_4807);
nand U1404 (N_1404,In_2873,In_1523);
xor U1405 (N_1405,In_2270,In_1144);
and U1406 (N_1406,In_278,In_4939);
nand U1407 (N_1407,N_64,N_509);
xnor U1408 (N_1408,In_2023,In_709);
nand U1409 (N_1409,In_2932,N_741);
or U1410 (N_1410,In_3266,In_4993);
or U1411 (N_1411,In_3436,In_2954);
and U1412 (N_1412,In_3601,N_631);
and U1413 (N_1413,N_903,N_692);
nand U1414 (N_1414,N_454,In_2988);
or U1415 (N_1415,In_3047,In_3211);
xnor U1416 (N_1416,In_2474,In_2749);
xor U1417 (N_1417,In_4461,In_4491);
and U1418 (N_1418,In_484,In_4015);
or U1419 (N_1419,N_785,N_848);
or U1420 (N_1420,In_2519,In_285);
or U1421 (N_1421,N_891,In_73);
or U1422 (N_1422,N_199,In_78);
or U1423 (N_1423,In_1131,N_96);
and U1424 (N_1424,In_494,In_4258);
and U1425 (N_1425,In_977,In_4637);
and U1426 (N_1426,In_1768,In_2267);
nor U1427 (N_1427,In_2605,In_4035);
nand U1428 (N_1428,In_3053,In_2024);
nand U1429 (N_1429,In_3707,In_3319);
or U1430 (N_1430,In_410,N_337);
or U1431 (N_1431,N_331,In_902);
nor U1432 (N_1432,In_1211,In_2887);
and U1433 (N_1433,N_754,In_2411);
nor U1434 (N_1434,In_1281,In_4047);
and U1435 (N_1435,In_4156,N_624);
nor U1436 (N_1436,In_3450,In_4709);
nand U1437 (N_1437,In_3662,In_1672);
nor U1438 (N_1438,In_4285,In_1973);
and U1439 (N_1439,In_3345,In_80);
or U1440 (N_1440,In_4641,In_3616);
or U1441 (N_1441,N_960,In_4112);
and U1442 (N_1442,N_764,N_721);
or U1443 (N_1443,In_3511,In_3039);
or U1444 (N_1444,In_3251,In_1934);
nor U1445 (N_1445,N_279,N_619);
and U1446 (N_1446,In_2286,In_3735);
and U1447 (N_1447,N_146,In_3362);
and U1448 (N_1448,In_1382,N_79);
and U1449 (N_1449,In_3094,In_693);
and U1450 (N_1450,In_1743,In_4890);
nor U1451 (N_1451,In_2174,In_4679);
or U1452 (N_1452,In_4009,In_673);
and U1453 (N_1453,In_2915,In_4626);
nor U1454 (N_1454,In_4422,In_2084);
nor U1455 (N_1455,In_633,In_3405);
and U1456 (N_1456,In_3277,In_1069);
or U1457 (N_1457,In_1777,In_203);
or U1458 (N_1458,In_3433,In_2122);
nand U1459 (N_1459,In_4353,N_477);
nor U1460 (N_1460,In_3019,In_4737);
nor U1461 (N_1461,N_521,In_1874);
and U1462 (N_1462,In_4113,N_680);
nor U1463 (N_1463,N_849,In_773);
nor U1464 (N_1464,In_4861,N_768);
or U1465 (N_1465,N_633,In_4868);
or U1466 (N_1466,In_4728,In_43);
xor U1467 (N_1467,N_282,In_2294);
nand U1468 (N_1468,N_907,N_869);
xnor U1469 (N_1469,In_283,N_8);
nor U1470 (N_1470,In_4910,In_3198);
xnor U1471 (N_1471,In_3629,N_844);
nor U1472 (N_1472,N_589,In_1106);
or U1473 (N_1473,In_3693,In_4619);
nand U1474 (N_1474,In_25,N_210);
or U1475 (N_1475,N_184,In_2356);
nand U1476 (N_1476,N_677,In_705);
and U1477 (N_1477,In_2652,In_2422);
xnor U1478 (N_1478,In_1537,In_4368);
nor U1479 (N_1479,In_3101,In_1719);
nand U1480 (N_1480,In_1543,In_3323);
nand U1481 (N_1481,In_2801,In_3451);
xnor U1482 (N_1482,In_4238,In_4773);
xnor U1483 (N_1483,In_3194,In_4163);
or U1484 (N_1484,N_711,In_212);
nand U1485 (N_1485,In_3175,In_4417);
nor U1486 (N_1486,In_2814,In_2096);
or U1487 (N_1487,In_1199,N_936);
nand U1488 (N_1488,N_84,In_4633);
xor U1489 (N_1489,N_383,N_414);
xnor U1490 (N_1490,N_147,N_417);
nor U1491 (N_1491,N_503,In_1084);
xor U1492 (N_1492,In_2202,In_3409);
or U1493 (N_1493,In_2399,In_4815);
nor U1494 (N_1494,N_393,In_4851);
and U1495 (N_1495,In_1090,In_2942);
xor U1496 (N_1496,In_1118,In_2835);
xnor U1497 (N_1497,In_4393,In_2907);
and U1498 (N_1498,N_658,In_314);
and U1499 (N_1499,In_4763,In_3984);
nor U1500 (N_1500,In_4998,In_3321);
nand U1501 (N_1501,In_1122,In_1699);
or U1502 (N_1502,In_1721,N_403);
xnor U1503 (N_1503,In_4144,In_4632);
and U1504 (N_1504,In_712,In_2986);
xnor U1505 (N_1505,N_506,In_1163);
or U1506 (N_1506,In_3626,In_1311);
xnor U1507 (N_1507,In_1705,In_2358);
and U1508 (N_1508,N_584,In_3001);
or U1509 (N_1509,In_1150,In_1363);
and U1510 (N_1510,N_1083,N_732);
and U1511 (N_1511,In_221,In_1711);
or U1512 (N_1512,In_2035,In_3937);
nor U1513 (N_1513,In_4459,N_579);
or U1514 (N_1514,N_1243,In_3245);
or U1515 (N_1515,N_747,In_940);
nor U1516 (N_1516,In_1974,In_2531);
xor U1517 (N_1517,N_1012,N_1322);
and U1518 (N_1518,N_669,N_825);
nand U1519 (N_1519,N_1407,N_300);
nor U1520 (N_1520,N_1119,In_4190);
or U1521 (N_1521,In_64,In_1198);
xor U1522 (N_1522,N_1247,In_157);
xnor U1523 (N_1523,N_252,In_919);
or U1524 (N_1524,In_1384,In_2461);
nor U1525 (N_1525,N_706,N_528);
xor U1526 (N_1526,In_4271,In_809);
xnor U1527 (N_1527,In_2618,N_917);
nor U1528 (N_1528,N_831,In_4579);
nor U1529 (N_1529,In_3012,N_1120);
nand U1530 (N_1530,In_3527,In_2039);
xnor U1531 (N_1531,In_574,In_366);
and U1532 (N_1532,In_501,In_2496);
or U1533 (N_1533,In_1588,In_3442);
xnor U1534 (N_1534,N_896,In_1667);
nand U1535 (N_1535,N_991,In_556);
nor U1536 (N_1536,In_4847,In_369);
or U1537 (N_1537,N_1468,In_1970);
nor U1538 (N_1538,In_1125,In_4045);
nor U1539 (N_1539,In_1983,In_4987);
xnor U1540 (N_1540,In_1465,In_2693);
and U1541 (N_1541,N_890,In_2855);
xor U1542 (N_1542,In_1034,In_1729);
or U1543 (N_1543,N_1003,N_1325);
nor U1544 (N_1544,In_4104,In_2792);
nor U1545 (N_1545,In_2836,In_3373);
nand U1546 (N_1546,N_1141,In_2859);
nand U1547 (N_1547,In_2752,N_209);
nand U1548 (N_1548,In_1232,In_4507);
or U1549 (N_1549,In_288,In_252);
nor U1550 (N_1550,In_422,N_426);
nand U1551 (N_1551,In_4023,N_1142);
nor U1552 (N_1552,In_1088,In_1773);
xnor U1553 (N_1553,N_1157,In_52);
or U1554 (N_1554,In_3638,In_3721);
xnor U1555 (N_1555,In_4657,In_119);
and U1556 (N_1556,N_1106,In_4789);
and U1557 (N_1557,In_4703,In_2187);
nor U1558 (N_1558,N_559,N_323);
xnor U1559 (N_1559,In_1366,In_1925);
nand U1560 (N_1560,N_310,N_475);
and U1561 (N_1561,In_3113,N_37);
xor U1562 (N_1562,N_698,In_1953);
nand U1563 (N_1563,N_625,In_1510);
nor U1564 (N_1564,In_3341,In_1099);
xnor U1565 (N_1565,In_1535,N_655);
xor U1566 (N_1566,In_1299,In_3743);
xnor U1567 (N_1567,In_1206,In_3017);
nand U1568 (N_1568,N_1398,In_3587);
xor U1569 (N_1569,N_1246,In_1172);
or U1570 (N_1570,In_45,N_937);
and U1571 (N_1571,In_224,In_4854);
nand U1572 (N_1572,N_667,N_1498);
nand U1573 (N_1573,In_3862,In_4548);
nor U1574 (N_1574,In_1436,In_3588);
or U1575 (N_1575,N_332,In_2287);
xor U1576 (N_1576,In_90,In_2613);
and U1577 (N_1577,N_1211,N_1224);
or U1578 (N_1578,In_4026,In_1021);
or U1579 (N_1579,In_1492,N_1034);
or U1580 (N_1580,In_274,In_549);
nor U1581 (N_1581,N_220,In_1078);
xnor U1582 (N_1582,In_1445,N_1291);
nor U1583 (N_1583,N_1190,In_4187);
nand U1584 (N_1584,In_2211,N_767);
and U1585 (N_1585,N_913,N_274);
and U1586 (N_1586,N_1091,In_1416);
or U1587 (N_1587,In_2030,N_212);
xor U1588 (N_1588,In_1354,In_24);
nand U1589 (N_1589,N_842,In_704);
nor U1590 (N_1590,In_595,N_1273);
or U1591 (N_1591,N_751,N_726);
or U1592 (N_1592,In_4855,In_3962);
nor U1593 (N_1593,In_1939,In_310);
nand U1594 (N_1594,In_433,In_3861);
and U1595 (N_1595,In_699,In_1693);
nor U1596 (N_1596,In_2579,In_971);
and U1597 (N_1597,In_3792,In_2200);
and U1598 (N_1598,N_1495,In_1058);
xor U1599 (N_1599,N_472,In_416);
or U1600 (N_1600,In_4578,In_2704);
xnor U1601 (N_1601,In_1159,N_237);
nor U1602 (N_1602,N_863,In_911);
xnor U1603 (N_1603,In_2707,In_3882);
or U1604 (N_1604,In_3008,In_1734);
nor U1605 (N_1605,N_1450,In_4600);
and U1606 (N_1606,N_870,N_857);
xnor U1607 (N_1607,N_1132,In_2585);
nand U1608 (N_1608,In_2456,In_3463);
and U1609 (N_1609,In_2430,In_3859);
nand U1610 (N_1610,In_4942,In_962);
or U1611 (N_1611,N_1174,In_3533);
nand U1612 (N_1612,N_1428,N_254);
nand U1613 (N_1613,In_3529,In_4790);
or U1614 (N_1614,In_4484,N_281);
or U1615 (N_1615,In_3911,In_2258);
or U1616 (N_1616,In_572,In_344);
or U1617 (N_1617,In_4695,In_4360);
or U1618 (N_1618,N_1114,In_357);
or U1619 (N_1619,N_556,In_2687);
nand U1620 (N_1620,N_958,In_1850);
xnor U1621 (N_1621,In_8,In_3775);
or U1622 (N_1622,In_3477,In_4907);
xnor U1623 (N_1623,In_3314,N_498);
and U1624 (N_1624,In_4355,In_3318);
xnor U1625 (N_1625,In_4443,In_3652);
or U1626 (N_1626,N_1272,N_895);
or U1627 (N_1627,N_1235,In_792);
nor U1628 (N_1628,N_1277,N_932);
or U1629 (N_1629,In_4820,In_4495);
xor U1630 (N_1630,In_1781,In_1832);
and U1631 (N_1631,In_1649,N_775);
nor U1632 (N_1632,N_1275,N_603);
or U1633 (N_1633,In_2824,In_2738);
and U1634 (N_1634,In_2964,In_2309);
xnor U1635 (N_1635,In_1654,N_83);
nand U1636 (N_1636,In_1589,In_4534);
xor U1637 (N_1637,In_4718,In_2765);
xor U1638 (N_1638,N_1290,In_4980);
or U1639 (N_1639,In_2535,In_2818);
or U1640 (N_1640,In_3685,In_4650);
xnor U1641 (N_1641,In_1497,In_1343);
nor U1642 (N_1642,In_2242,In_2695);
xnor U1643 (N_1643,In_4300,In_951);
nor U1644 (N_1644,N_317,N_901);
nor U1645 (N_1645,N_1438,In_3614);
or U1646 (N_1646,In_4756,In_1838);
nand U1647 (N_1647,In_4329,In_2341);
xnor U1648 (N_1648,N_731,In_2203);
nor U1649 (N_1649,In_279,In_102);
xnor U1650 (N_1650,In_678,N_1067);
or U1651 (N_1651,In_1629,In_1338);
nand U1652 (N_1652,N_1315,N_81);
nor U1653 (N_1653,N_114,In_38);
and U1654 (N_1654,In_1060,In_1234);
nor U1655 (N_1655,N_1431,In_763);
and U1656 (N_1656,In_3247,In_1971);
nand U1657 (N_1657,In_3161,N_1011);
nand U1658 (N_1658,In_4877,In_3538);
xor U1659 (N_1659,N_851,N_720);
and U1660 (N_1660,In_4803,In_3347);
xnor U1661 (N_1661,N_292,In_743);
xnor U1662 (N_1662,N_1105,In_4005);
xnor U1663 (N_1663,In_3888,In_2690);
and U1664 (N_1664,In_1186,In_3482);
nand U1665 (N_1665,In_1760,N_1116);
or U1666 (N_1666,In_4424,In_1401);
and U1667 (N_1667,In_4732,N_854);
nor U1668 (N_1668,In_3415,In_4795);
or U1669 (N_1669,In_249,In_4394);
or U1670 (N_1670,In_97,In_795);
nor U1671 (N_1671,In_2029,In_2464);
and U1672 (N_1672,N_289,In_2631);
nor U1673 (N_1673,In_184,N_694);
xor U1674 (N_1674,In_789,N_443);
xnor U1675 (N_1675,N_131,In_4320);
nand U1676 (N_1676,In_1181,In_952);
xnor U1677 (N_1677,In_2302,In_4908);
xnor U1678 (N_1678,N_1193,In_44);
and U1679 (N_1679,In_1628,N_834);
and U1680 (N_1680,N_328,N_1084);
and U1681 (N_1681,In_2484,In_702);
or U1682 (N_1682,N_405,N_1073);
nand U1683 (N_1683,In_1487,In_1549);
and U1684 (N_1684,In_3141,In_1816);
xnor U1685 (N_1685,N_66,In_4948);
and U1686 (N_1686,In_1921,In_1453);
nand U1687 (N_1687,N_1424,In_3534);
or U1688 (N_1688,In_2990,In_4906);
xor U1689 (N_1689,In_2747,N_7);
and U1690 (N_1690,In_4059,N_1478);
xnor U1691 (N_1691,In_645,In_1710);
nor U1692 (N_1692,In_1615,In_2116);
or U1693 (N_1693,In_1251,In_4581);
xor U1694 (N_1694,N_455,In_1945);
and U1695 (N_1695,N_705,N_1433);
xor U1696 (N_1696,N_213,In_3032);
or U1697 (N_1697,In_3168,N_24);
nor U1698 (N_1698,In_4462,In_2760);
or U1699 (N_1699,In_1126,N_859);
nor U1700 (N_1700,In_54,In_996);
nand U1701 (N_1701,In_138,N_1144);
and U1702 (N_1702,In_3812,In_4371);
nor U1703 (N_1703,In_174,In_4772);
nor U1704 (N_1704,N_494,N_798);
nand U1705 (N_1705,In_2298,In_1758);
nor U1706 (N_1706,In_3970,In_151);
xnor U1707 (N_1707,In_3225,In_3799);
nand U1708 (N_1708,In_2979,N_1163);
nand U1709 (N_1709,N_759,In_698);
nand U1710 (N_1710,N_511,N_496);
and U1711 (N_1711,In_1006,N_833);
and U1712 (N_1712,In_4821,In_4254);
nand U1713 (N_1713,In_3271,N_1065);
xnor U1714 (N_1714,In_3192,N_21);
xor U1715 (N_1715,In_2272,N_1154);
nor U1716 (N_1716,In_1140,In_4664);
or U1717 (N_1717,N_1485,In_1241);
nor U1718 (N_1718,In_1331,N_1423);
nand U1719 (N_1719,N_340,In_1842);
nand U1720 (N_1720,N_904,In_92);
nor U1721 (N_1721,In_2471,In_15);
or U1722 (N_1722,N_1343,In_2758);
xor U1723 (N_1723,N_1323,In_2515);
nor U1724 (N_1724,In_3060,In_2374);
nor U1725 (N_1725,In_3569,In_3887);
nor U1726 (N_1726,In_2176,In_188);
or U1727 (N_1727,In_2673,In_2345);
nand U1728 (N_1728,In_4569,In_1865);
xnor U1729 (N_1729,In_627,N_1149);
and U1730 (N_1730,N_552,In_4083);
xor U1731 (N_1731,N_1066,In_4408);
nor U1732 (N_1732,N_196,In_191);
nand U1733 (N_1733,In_4874,In_3584);
or U1734 (N_1734,N_622,In_879);
nand U1735 (N_1735,In_3107,In_2856);
and U1736 (N_1736,N_1487,N_1264);
and U1737 (N_1737,In_502,N_1192);
and U1738 (N_1738,N_1266,N_728);
or U1739 (N_1739,In_3714,In_2773);
or U1740 (N_1740,In_1019,In_1253);
xor U1741 (N_1741,In_1859,In_2212);
nand U1742 (N_1742,N_1439,In_4315);
nor U1743 (N_1743,In_4917,N_707);
and U1744 (N_1744,N_666,In_4951);
xnor U1745 (N_1745,In_2028,N_1446);
xor U1746 (N_1746,In_651,In_4506);
xor U1747 (N_1747,N_922,In_390);
nand U1748 (N_1748,N_800,N_1359);
nor U1749 (N_1749,In_3564,In_711);
xor U1750 (N_1750,In_358,N_1023);
nor U1751 (N_1751,N_1052,In_4262);
nor U1752 (N_1752,In_3204,N_1160);
and U1753 (N_1753,N_1305,In_770);
nand U1754 (N_1754,In_1782,N_931);
and U1755 (N_1755,N_1056,In_2357);
and U1756 (N_1756,N_1176,N_972);
nor U1757 (N_1757,N_708,In_4717);
and U1758 (N_1758,In_4197,In_4455);
nand U1759 (N_1759,In_2614,In_906);
xnor U1760 (N_1760,In_4354,N_1327);
nand U1761 (N_1761,N_1260,N_1121);
xnor U1762 (N_1762,N_318,N_518);
nor U1763 (N_1763,In_77,In_4174);
nor U1764 (N_1764,In_4786,In_1491);
or U1765 (N_1765,In_4883,N_154);
nand U1766 (N_1766,N_1317,N_1090);
and U1767 (N_1767,N_1218,N_256);
nand U1768 (N_1768,In_4414,In_2815);
nand U1769 (N_1769,In_3334,N_1206);
nand U1770 (N_1770,In_730,N_1072);
nand U1771 (N_1771,N_875,N_1469);
or U1772 (N_1772,N_1076,In_2288);
xor U1773 (N_1773,N_378,In_2250);
nor U1774 (N_1774,In_4946,N_353);
nor U1775 (N_1775,N_562,In_1864);
xnor U1776 (N_1776,N_581,In_1087);
nor U1777 (N_1777,In_3549,In_2225);
nor U1778 (N_1778,N_753,In_1521);
xor U1779 (N_1779,N_540,In_1986);
xor U1780 (N_1780,In_4531,In_3339);
or U1781 (N_1781,In_1906,In_176);
nor U1782 (N_1782,N_710,N_682);
and U1783 (N_1783,In_4615,In_2056);
nor U1784 (N_1784,N_1425,In_2551);
or U1785 (N_1785,In_2703,N_269);
or U1786 (N_1786,In_1759,In_2649);
xor U1787 (N_1787,In_3850,N_1415);
xor U1788 (N_1788,In_1357,In_2592);
and U1789 (N_1789,In_2546,In_355);
nand U1790 (N_1790,N_1403,In_105);
xor U1791 (N_1791,In_219,N_214);
nor U1792 (N_1792,N_485,In_2479);
nand U1793 (N_1793,In_91,N_1376);
nor U1794 (N_1794,N_966,N_396);
or U1795 (N_1795,In_2235,N_599);
xor U1796 (N_1796,In_804,N_145);
nand U1797 (N_1797,N_1156,N_905);
and U1798 (N_1798,In_4612,N_1103);
or U1799 (N_1799,In_3516,In_373);
or U1800 (N_1800,In_1818,In_3873);
xor U1801 (N_1801,N_1018,In_2995);
nand U1802 (N_1802,In_1733,In_4198);
nor U1803 (N_1803,N_1029,In_4250);
nor U1804 (N_1804,N_715,In_4447);
nor U1805 (N_1805,N_1347,In_1966);
nand U1806 (N_1806,In_3759,In_3005);
and U1807 (N_1807,In_577,N_459);
and U1808 (N_1808,N_488,N_88);
or U1809 (N_1809,In_3827,N_229);
nor U1810 (N_1810,N_1050,N_433);
nand U1811 (N_1811,In_575,In_4232);
nand U1812 (N_1812,In_3982,N_424);
xor U1813 (N_1813,N_952,In_3666);
nand U1814 (N_1814,In_4555,N_612);
nor U1815 (N_1815,In_4961,N_608);
nor U1816 (N_1816,N_1184,N_1051);
nand U1817 (N_1817,In_3551,In_3099);
and U1818 (N_1818,In_3444,In_111);
or U1819 (N_1819,In_1669,N_770);
xor U1820 (N_1820,In_1352,In_32);
and U1821 (N_1821,In_2648,In_4549);
nand U1822 (N_1822,N_369,In_14);
or U1823 (N_1823,In_926,In_1469);
nor U1824 (N_1824,N_293,In_4565);
or U1825 (N_1825,N_172,In_2303);
and U1826 (N_1826,In_1388,In_1902);
or U1827 (N_1827,In_3324,In_231);
xnor U1828 (N_1828,In_2232,N_804);
nor U1829 (N_1829,In_3127,N_109);
xor U1830 (N_1830,In_3623,In_2155);
nor U1831 (N_1831,N_596,N_324);
nor U1832 (N_1832,N_1016,In_541);
xnor U1833 (N_1833,In_115,In_1271);
xnor U1834 (N_1834,In_89,N_1092);
nor U1835 (N_1835,In_2009,In_4666);
or U1836 (N_1836,N_1000,In_3811);
and U1837 (N_1837,N_979,In_2467);
nor U1838 (N_1838,In_4892,In_4024);
nor U1839 (N_1839,N_1098,In_3801);
xor U1840 (N_1840,In_2823,In_2898);
or U1841 (N_1841,In_3011,In_3844);
and U1842 (N_1842,In_402,In_3857);
xor U1843 (N_1843,In_2723,N_1460);
nand U1844 (N_1844,In_1221,In_3389);
xnor U1845 (N_1845,N_1427,In_2195);
and U1846 (N_1846,N_1296,N_1001);
or U1847 (N_1847,N_1009,In_2917);
and U1848 (N_1848,In_1434,N_1316);
xnor U1849 (N_1849,In_3646,In_3610);
nand U1850 (N_1850,In_4266,N_176);
xnor U1851 (N_1851,N_679,In_225);
and U1852 (N_1852,N_871,N_5);
and U1853 (N_1853,In_1135,In_562);
and U1854 (N_1854,N_264,In_942);
nand U1855 (N_1855,In_2696,In_2994);
nand U1856 (N_1856,In_727,N_1134);
or U1857 (N_1857,In_1542,In_3050);
or U1858 (N_1858,N_1375,In_2323);
or U1859 (N_1859,In_3654,In_2310);
nand U1860 (N_1860,N_722,In_578);
nor U1861 (N_1861,N_776,In_388);
and U1862 (N_1862,In_4967,In_2088);
nor U1863 (N_1863,In_3279,In_3821);
nor U1864 (N_1864,In_396,N_222);
nand U1865 (N_1865,N_92,In_2443);
or U1866 (N_1866,N_1126,In_1156);
and U1867 (N_1867,In_3406,In_4299);
xnor U1868 (N_1868,In_2190,In_4460);
nand U1869 (N_1869,N_180,In_1779);
nand U1870 (N_1870,In_384,N_724);
and U1871 (N_1871,N_942,In_4497);
nor U1872 (N_1872,In_1002,In_2770);
nor U1873 (N_1873,N_723,N_623);
or U1874 (N_1874,N_85,N_519);
and U1875 (N_1875,In_3688,N_373);
or U1876 (N_1876,In_3248,In_4175);
xor U1877 (N_1877,In_4774,In_282);
xor U1878 (N_1878,N_510,In_218);
nor U1879 (N_1879,N_1389,N_223);
or U1880 (N_1880,In_455,In_826);
xor U1881 (N_1881,In_1109,In_830);
and U1882 (N_1882,N_265,N_1219);
nand U1883 (N_1883,In_893,N_482);
and U1884 (N_1884,In_4134,In_779);
or U1885 (N_1885,In_2759,N_54);
and U1886 (N_1886,In_4994,In_4092);
nand U1887 (N_1887,In_3674,In_3836);
nor U1888 (N_1888,N_1047,In_4713);
or U1889 (N_1889,In_4361,In_2044);
nand U1890 (N_1890,In_3531,N_71);
xor U1891 (N_1891,In_4848,In_3657);
nor U1892 (N_1892,N_1022,N_1370);
and U1893 (N_1893,In_649,N_1383);
and U1894 (N_1894,In_3122,In_3979);
nor U1895 (N_1895,In_3671,N_1055);
nand U1896 (N_1896,N_1231,In_1704);
nor U1897 (N_1897,N_673,In_4233);
xor U1898 (N_1898,In_4924,In_1621);
and U1899 (N_1899,N_1213,In_2664);
nand U1900 (N_1900,N_1086,In_1989);
or U1901 (N_1901,In_141,In_1377);
nor U1902 (N_1902,N_1227,In_4613);
xor U1903 (N_1903,In_3942,In_2952);
or U1904 (N_1904,In_3805,N_925);
xor U1905 (N_1905,In_4488,In_3398);
nor U1906 (N_1906,N_1166,N_843);
and U1907 (N_1907,N_1108,N_676);
nor U1908 (N_1908,In_4519,In_3013);
nand U1909 (N_1909,In_2416,In_4131);
nor U1910 (N_1910,N_1364,In_3434);
or U1911 (N_1911,In_3589,N_1430);
and U1912 (N_1912,In_1505,In_2277);
xor U1913 (N_1913,In_3595,In_3676);
xor U1914 (N_1914,In_766,N_30);
nor U1915 (N_1915,N_28,In_1962);
nand U1916 (N_1916,In_2739,In_989);
nand U1917 (N_1917,In_4634,N_801);
or U1918 (N_1918,In_800,In_67);
nand U1919 (N_1919,In_3579,In_2349);
or U1920 (N_1920,In_3738,In_116);
xor U1921 (N_1921,In_3803,In_2697);
or U1922 (N_1922,In_354,N_1220);
or U1923 (N_1923,N_999,In_4688);
xor U1924 (N_1924,In_211,N_23);
xnor U1925 (N_1925,In_4396,N_73);
or U1926 (N_1926,In_3883,In_4139);
nor U1927 (N_1927,In_132,In_4496);
nor U1928 (N_1928,In_3897,N_1278);
nor U1929 (N_1929,In_3950,In_2602);
and U1930 (N_1930,N_1079,In_573);
xnor U1931 (N_1931,In_3841,In_1808);
nor U1932 (N_1932,In_1508,In_548);
and U1933 (N_1933,In_4007,In_2280);
nor U1934 (N_1934,N_219,In_327);
or U1935 (N_1935,In_4997,N_1332);
nor U1936 (N_1936,In_3989,N_627);
nor U1937 (N_1937,In_3174,In_4210);
and U1938 (N_1938,N_44,In_2927);
and U1939 (N_1939,In_2902,N_62);
and U1940 (N_1940,In_3187,In_2058);
or U1941 (N_1941,In_1688,In_3368);
and U1942 (N_1942,In_1222,In_3939);
nand U1943 (N_1943,In_3049,N_397);
nand U1944 (N_1944,In_1996,In_1638);
nand U1945 (N_1945,In_1456,In_3655);
or U1946 (N_1946,In_3285,In_1957);
or U1947 (N_1947,In_2085,In_3820);
nor U1948 (N_1948,N_527,In_1043);
or U1949 (N_1949,In_1276,In_4434);
or U1950 (N_1950,N_738,N_977);
or U1951 (N_1951,N_1130,N_407);
nand U1952 (N_1952,N_1467,In_2117);
or U1953 (N_1953,In_2709,In_3387);
xor U1954 (N_1954,N_1418,In_2391);
nor U1955 (N_1955,In_2336,In_1665);
or U1956 (N_1956,N_1443,N_1301);
or U1957 (N_1957,In_1188,In_304);
or U1958 (N_1958,In_2865,N_1146);
or U1959 (N_1959,N_1417,In_236);
nand U1960 (N_1960,In_876,In_2556);
or U1961 (N_1961,In_2233,In_3523);
nor U1962 (N_1962,In_2073,N_1379);
nor U1963 (N_1963,In_3106,N_1204);
nand U1964 (N_1964,In_1959,In_104);
xnor U1965 (N_1965,In_585,In_3043);
and U1966 (N_1966,In_707,In_2032);
and U1967 (N_1967,In_4801,In_3931);
nand U1968 (N_1968,N_1054,In_796);
nand U1969 (N_1969,N_1031,In_4838);
xor U1970 (N_1970,In_3807,N_1208);
xor U1971 (N_1971,In_1361,In_1681);
or U1972 (N_1972,In_2010,N_1286);
nor U1973 (N_1973,In_2708,In_480);
nor U1974 (N_1974,In_2163,N_1324);
and U1975 (N_1975,N_1395,In_4599);
and U1976 (N_1976,In_1976,In_2249);
or U1977 (N_1977,In_2869,In_583);
nor U1978 (N_1978,In_1301,In_3116);
xnor U1979 (N_1979,N_1447,In_1027);
and U1980 (N_1980,N_1267,N_40);
xnor U1981 (N_1981,In_3260,In_2415);
xnor U1982 (N_1982,In_53,In_4428);
nand U1983 (N_1983,N_576,In_3065);
xor U1984 (N_1984,N_1232,In_3426);
xnor U1985 (N_1985,In_4911,In_4671);
nor U1986 (N_1986,N_225,In_4142);
nand U1987 (N_1987,In_566,In_1735);
or U1988 (N_1988,N_1372,In_2444);
nor U1989 (N_1989,N_1019,In_1327);
xnor U1990 (N_1990,N_713,In_2962);
nor U1991 (N_1991,In_3893,N_1406);
xnor U1992 (N_1992,In_3269,In_4260);
xnor U1993 (N_1993,In_1353,In_2914);
and U1994 (N_1994,In_4328,N_1362);
and U1995 (N_1995,In_914,In_1980);
nand U1996 (N_1996,N_1113,In_1267);
nand U1997 (N_1997,N_1444,In_4598);
and U1998 (N_1998,N_885,In_82);
and U1999 (N_1999,In_4309,In_2827);
and U2000 (N_2000,In_4184,N_1926);
and U2001 (N_2001,N_1666,N_1696);
nor U2002 (N_2002,In_2441,In_4526);
and U2003 (N_2003,N_1996,In_4481);
and U2004 (N_2004,N_1695,N_1230);
nor U2005 (N_2005,N_1843,N_1229);
or U2006 (N_2006,In_3312,In_75);
nand U2007 (N_2007,N_1600,N_664);
nor U2008 (N_2008,N_474,N_648);
nand U2009 (N_2009,In_2082,In_179);
or U2010 (N_2010,N_526,In_1061);
xor U2011 (N_2011,In_1476,N_1862);
or U2012 (N_2012,In_3292,In_2118);
xnor U2013 (N_2013,N_276,N_1550);
nand U2014 (N_2014,In_2641,N_1733);
nand U2015 (N_2015,N_249,In_4178);
xnor U2016 (N_2016,N_688,In_4862);
and U2017 (N_2017,In_601,In_2900);
nand U2018 (N_2018,N_1738,N_536);
and U2019 (N_2019,In_427,In_1652);
nand U2020 (N_2020,In_4028,In_1658);
nand U2021 (N_2021,N_1901,In_2946);
nand U2022 (N_2022,In_1879,N_370);
xnor U2023 (N_2023,In_4668,In_3252);
xnor U2024 (N_2024,In_1072,N_457);
or U2025 (N_2025,N_607,N_1539);
xnor U2026 (N_2026,In_2160,N_1613);
nand U2027 (N_2027,N_1780,N_144);
or U2028 (N_2028,In_3439,N_1556);
nand U2029 (N_2029,N_638,In_4021);
xor U2030 (N_2030,N_1821,N_1580);
nand U2031 (N_2031,In_1346,N_1925);
and U2032 (N_2032,In_3558,N_1123);
nor U2033 (N_2033,N_733,In_1451);
nor U2034 (N_2034,In_2149,N_391);
xnor U2035 (N_2035,In_1285,In_393);
and U2036 (N_2036,In_2637,In_3437);
xor U2037 (N_2037,In_1108,N_1795);
nand U2038 (N_2038,In_4116,N_1205);
nor U2039 (N_2039,In_3973,In_2397);
or U2040 (N_2040,N_1020,In_183);
nand U2041 (N_2041,In_2363,In_3110);
nand U2042 (N_2042,In_4661,In_2575);
xnor U2043 (N_2043,N_1458,In_2744);
and U2044 (N_2044,In_1746,In_802);
nand U2045 (N_2045,N_939,N_129);
nand U2046 (N_2046,N_1697,In_3886);
xor U2047 (N_2047,In_3751,In_419);
and U2048 (N_2048,In_4090,In_3938);
or U2049 (N_2049,N_1619,N_326);
xor U2050 (N_2050,N_1571,In_1190);
and U2051 (N_2051,In_3848,N_444);
and U2052 (N_2052,In_2985,N_1671);
and U2053 (N_2053,N_717,N_1701);
nor U2054 (N_2054,In_854,N_1191);
nor U2055 (N_2055,N_204,In_3246);
and U2056 (N_2056,In_3237,N_1944);
or U2057 (N_2057,In_2706,In_4914);
nand U2058 (N_2058,In_3996,In_1056);
and U2059 (N_2059,N_926,In_3823);
and U2060 (N_2060,In_4644,N_1692);
or U2061 (N_2061,In_243,N_329);
or U2062 (N_2062,In_932,In_4781);
xor U2063 (N_2063,In_2092,In_2772);
and U2064 (N_2064,In_4141,N_1380);
xnor U2065 (N_2065,In_4863,N_448);
and U2066 (N_2066,N_165,In_3723);
nand U2067 (N_2067,N_594,In_4791);
xnor U2068 (N_2068,In_623,In_736);
nand U2069 (N_2069,N_1770,N_1170);
nor U2070 (N_2070,N_1493,In_1187);
nand U2071 (N_2071,N_1030,N_790);
nand U2072 (N_2072,N_626,In_3684);
xor U2073 (N_2073,In_479,In_4218);
nor U2074 (N_2074,In_3316,In_428);
nand U2075 (N_2075,In_4062,N_272);
nand U2076 (N_2076,In_3830,N_1473);
nand U2077 (N_2077,In_2457,N_1905);
xnor U2078 (N_2078,N_1785,N_1577);
nand U2079 (N_2079,In_3242,N_1241);
or U2080 (N_2080,In_3371,N_1339);
or U2081 (N_2081,In_319,In_2312);
xnor U2082 (N_2082,N_150,In_464);
xor U2083 (N_2083,N_1895,N_661);
or U2084 (N_2084,In_860,N_1429);
xnor U2085 (N_2085,In_1129,N_563);
nand U2086 (N_2086,N_588,N_1568);
or U2087 (N_2087,In_4002,N_1508);
nor U2088 (N_2088,N_441,N_1522);
nor U2089 (N_2089,N_700,In_3673);
and U2090 (N_2090,In_3481,In_4359);
and U2091 (N_2091,N_1612,In_843);
and U2092 (N_2092,N_1922,N_436);
xor U2093 (N_2093,In_2246,N_1334);
nor U2094 (N_2094,In_1290,In_4741);
nor U2095 (N_2095,N_810,In_1220);
nor U2096 (N_2096,In_4020,In_2992);
or U2097 (N_2097,N_492,In_3418);
and U2098 (N_2098,N_1829,In_3002);
and U2099 (N_2099,N_1295,N_915);
xor U2100 (N_2100,N_807,In_3202);
nand U2101 (N_2101,In_4482,N_1225);
nor U2102 (N_2102,In_4483,In_517);
nor U2103 (N_2103,N_1356,In_4562);
nand U2104 (N_2104,In_364,In_4724);
and U2105 (N_2105,N_368,In_4602);
nand U2106 (N_2106,N_803,N_837);
nand U2107 (N_2107,In_1564,In_2101);
nor U2108 (N_2108,In_4730,In_2949);
and U2109 (N_2109,N_1769,N_497);
xor U2110 (N_2110,In_4647,In_723);
and U2111 (N_2111,In_4206,N_1969);
nand U2112 (N_2112,In_3594,In_2477);
and U2113 (N_2113,In_4923,N_1963);
xnor U2114 (N_2114,In_2209,N_697);
nor U2115 (N_2115,N_1649,In_1732);
and U2116 (N_2116,In_1467,N_1528);
and U2117 (N_2117,In_1877,In_883);
or U2118 (N_2118,In_1761,In_2330);
nor U2119 (N_2119,In_2192,N_1989);
nor U2120 (N_2120,In_643,In_2359);
nand U2121 (N_2121,In_3335,In_2571);
nand U2122 (N_2122,N_268,N_1946);
nand U2123 (N_2123,N_772,N_1849);
nor U2124 (N_2124,In_3493,N_183);
or U2125 (N_2125,In_3667,N_1841);
nor U2126 (N_2126,In_1228,N_944);
and U2127 (N_2127,N_1392,In_2304);
xnor U2128 (N_2128,In_3165,In_2581);
xnor U2129 (N_2129,N_1835,In_193);
xnor U2130 (N_2130,In_2002,N_914);
nor U2131 (N_2131,N_1,In_4278);
nand U2132 (N_2132,In_2720,In_3498);
and U2133 (N_2133,In_4118,N_389);
and U2134 (N_2134,In_3597,N_1538);
nor U2135 (N_2135,In_1817,In_4471);
nand U2136 (N_2136,N_1760,In_3210);
nand U2137 (N_2137,In_3795,In_1031);
xnor U2138 (N_2138,N_484,In_3163);
and U2139 (N_2139,N_1564,N_439);
or U2140 (N_2140,In_2611,N_1448);
and U2141 (N_2141,In_84,N_1660);
nand U2142 (N_2142,In_866,In_1202);
and U2143 (N_2143,N_1853,In_3431);
nor U2144 (N_2144,In_1420,N_1361);
and U2145 (N_2145,N_1589,In_589);
nor U2146 (N_2146,In_3669,In_4080);
nor U2147 (N_2147,N_1518,In_1513);
or U2148 (N_2148,In_2139,In_4448);
xor U2149 (N_2149,N_1500,N_656);
xor U2150 (N_2150,N_1866,N_61);
nand U2151 (N_2151,In_2656,N_1558);
and U2152 (N_2152,In_3917,In_4407);
nand U2153 (N_2153,N_1186,N_1503);
nand U2154 (N_2154,N_1902,In_579);
xnor U2155 (N_2155,In_1194,In_1861);
or U2156 (N_2156,In_143,N_644);
xor U2157 (N_2157,N_1109,N_1754);
nand U2158 (N_2158,N_1402,In_2453);
xor U2159 (N_2159,N_535,In_3730);
or U2160 (N_2160,In_240,N_1663);
nand U2161 (N_2161,N_123,In_3581);
nor U2162 (N_2162,In_3617,N_1042);
xor U2163 (N_2163,N_670,N_1674);
or U2164 (N_2164,N_1044,In_1283);
nand U2165 (N_2165,In_3380,N_1271);
or U2166 (N_2166,In_2329,In_1160);
xnor U2167 (N_2167,N_1630,In_881);
xor U2168 (N_2168,N_1320,In_3521);
nor U2169 (N_2169,N_910,In_4378);
or U2170 (N_2170,In_4292,N_1879);
nand U2171 (N_2171,In_4323,N_1720);
nor U2172 (N_2172,N_965,N_1777);
xnor U2173 (N_2173,N_1257,N_1555);
nand U2174 (N_2174,In_4077,In_2214);
xor U2175 (N_2175,N_243,In_4628);
or U2176 (N_2176,In_3432,N_1700);
and U2177 (N_2177,In_4464,In_4521);
nor U2178 (N_2178,In_4257,In_2790);
nor U2179 (N_2179,In_4392,In_2179);
nor U2180 (N_2180,N_1151,N_344);
and U2181 (N_2181,In_4659,N_630);
nand U2182 (N_2182,N_166,In_169);
nand U2183 (N_2183,N_1125,In_1488);
nand U2184 (N_2184,N_1188,N_1725);
or U2185 (N_2185,In_2644,In_2318);
or U2186 (N_2186,In_2169,N_539);
and U2187 (N_2187,N_51,N_1153);
nand U2188 (N_2188,In_3794,N_1202);
and U2189 (N_2189,N_812,N_1699);
nor U2190 (N_2190,N_1158,In_4358);
nor U2191 (N_2191,N_1896,In_3217);
xnor U2192 (N_2192,In_622,In_4623);
nand U2193 (N_2193,N_1058,In_3452);
or U2194 (N_2194,In_1344,In_1730);
nand U2195 (N_2195,In_4485,In_305);
xnor U2196 (N_2196,In_1340,In_4873);
xor U2197 (N_2197,N_1851,N_1340);
nand U2198 (N_2198,In_4229,N_1884);
nor U2199 (N_2199,In_1164,In_3717);
nor U2200 (N_2200,In_1414,In_2728);
xnor U2201 (N_2201,N_1985,N_1891);
nor U2202 (N_2202,In_3562,N_1137);
or U2203 (N_2203,In_4542,In_4345);
and U2204 (N_2204,In_245,In_4313);
nor U2205 (N_2205,In_152,N_1390);
nand U2206 (N_2206,In_3182,N_473);
or U2207 (N_2207,In_2124,In_1485);
and U2208 (N_2208,In_2507,In_3350);
nor U2209 (N_2209,N_1413,N_440);
xor U2210 (N_2210,N_835,N_1656);
nand U2211 (N_2211,N_1553,N_1981);
or U2212 (N_2212,N_1887,In_4420);
or U2213 (N_2213,N_334,N_1514);
and U2214 (N_2214,N_830,In_983);
xor U2215 (N_2215,In_2598,In_4580);
xor U2216 (N_2216,N_1999,In_2408);
xnor U2217 (N_2217,In_399,In_1014);
and U2218 (N_2218,N_1653,In_266);
nand U2219 (N_2219,In_3509,N_1986);
or U2220 (N_2220,N_1686,N_546);
nor U2221 (N_2221,In_1992,N_1581);
or U2222 (N_2222,N_253,N_1165);
or U2223 (N_2223,In_2157,N_1739);
nand U2224 (N_2224,N_1823,In_1867);
and U2225 (N_2225,In_3062,In_603);
nor U2226 (N_2226,In_2360,In_1373);
xor U2227 (N_2227,N_1274,In_1620);
or U2228 (N_2228,N_181,In_2308);
and U2229 (N_2229,In_2778,In_3713);
or U2230 (N_2230,In_3590,N_1100);
xnor U2231 (N_2231,N_1570,In_320);
and U2232 (N_2232,In_500,N_1337);
nand U2233 (N_2233,In_1855,In_3244);
xnor U2234 (N_2234,In_4435,In_2133);
nand U2235 (N_2235,In_3598,In_3270);
and U2236 (N_2236,In_3635,In_571);
xor U2237 (N_2237,In_696,In_3399);
xnor U2238 (N_2238,In_2908,In_803);
nor U2239 (N_2239,In_3079,In_1950);
nand U2240 (N_2240,In_4743,In_2080);
or U2241 (N_2241,N_182,N_259);
or U2242 (N_2242,In_1428,In_4944);
nand U2243 (N_2243,In_4533,In_1502);
nand U2244 (N_2244,N_1876,In_3069);
and U2245 (N_2245,N_1677,In_1579);
and U2246 (N_2246,N_45,In_3541);
nand U2247 (N_2247,N_1551,N_1852);
nor U2248 (N_2248,N_1171,N_737);
nor U2249 (N_2249,In_2857,N_207);
nor U2250 (N_2250,N_1796,In_680);
and U2251 (N_2251,In_126,N_1776);
xor U2252 (N_2252,In_1793,N_39);
and U2253 (N_2253,In_3868,In_4844);
nand U2254 (N_2254,N_1248,N_416);
or U2255 (N_2255,In_4330,In_4406);
xor U2256 (N_2256,In_4100,N_1975);
xnor U2257 (N_2257,N_1800,In_2489);
and U2258 (N_2258,N_1346,N_1479);
or U2259 (N_2259,N_523,N_1745);
nand U2260 (N_2260,N_1833,In_4813);
nor U2261 (N_2261,N_1992,N_162);
and U2262 (N_2262,In_1898,In_2442);
and U2263 (N_2263,In_1305,N_1740);
nand U2264 (N_2264,In_11,N_1578);
and U2265 (N_2265,N_1878,N_1382);
or U2266 (N_2266,In_1569,In_4687);
nand U2267 (N_2267,In_1932,N_1936);
or U2268 (N_2268,N_1954,In_1236);
or U2269 (N_2269,In_4567,In_4962);
or U2270 (N_2270,In_4068,N_1270);
nand U2271 (N_2271,N_1249,N_1898);
and U2272 (N_2272,In_2651,In_846);
nand U2273 (N_2273,In_1348,In_3494);
nand U2274 (N_2274,In_684,N_1307);
nand U2275 (N_2275,N_1717,N_1793);
and U2276 (N_2276,In_1151,N_1911);
nand U2277 (N_2277,In_3864,In_1880);
nor U2278 (N_2278,In_1797,In_3880);
nor U2279 (N_2279,In_3556,N_398);
and U2280 (N_2280,N_657,In_554);
nand U2281 (N_2281,N_1948,In_4339);
or U2282 (N_2282,N_1929,In_1037);
nor U2283 (N_2283,N_126,In_178);
xor U2284 (N_2284,In_230,N_1304);
nand U2285 (N_2285,N_1662,N_1712);
nand U2286 (N_2286,In_1696,In_3884);
nand U2287 (N_2287,N_1207,In_2776);
and U2288 (N_2288,In_4893,N_814);
nor U2289 (N_2289,N_1505,In_2923);
or U2290 (N_2290,N_961,N_1909);
nand U2291 (N_2291,In_2145,In_1307);
xnor U2292 (N_2292,N_1920,In_2283);
xnor U2293 (N_2293,N_161,In_4202);
nor U2294 (N_2294,In_4295,N_1088);
xor U2295 (N_2295,In_2784,N_1579);
or U2296 (N_2296,N_1203,N_1180);
and U2297 (N_2297,N_1764,In_2771);
or U2298 (N_2298,In_1201,In_667);
nand U2299 (N_2299,N_1233,N_1694);
nor U2300 (N_2300,In_2402,N_963);
and U2301 (N_2301,In_825,In_2284);
nor U2302 (N_2302,In_1575,In_2712);
nor U2303 (N_2303,N_530,N_1675);
xnor U2304 (N_2304,In_2234,N_1348);
nor U2305 (N_2305,In_3737,N_153);
or U2306 (N_2306,N_1489,In_4720);
nand U2307 (N_2307,N_1057,In_1836);
xor U2308 (N_2308,N_1894,In_1592);
and U2309 (N_2309,In_3306,In_3933);
xor U2310 (N_2310,N_1294,In_2109);
nand U2311 (N_2311,N_1008,In_3774);
nor U2312 (N_2312,N_1609,In_2505);
nand U2313 (N_2313,N_350,In_4787);
and U2314 (N_2314,In_3928,N_1541);
and U2315 (N_2315,In_2754,In_1204);
or U2316 (N_2316,N_660,N_1605);
or U2317 (N_2317,In_2542,N_1434);
nand U2318 (N_2318,In_4953,In_3877);
and U2319 (N_2319,In_2826,In_1742);
xor U2320 (N_2320,In_4053,N_836);
or U2321 (N_2321,In_1685,In_2493);
nor U2322 (N_2322,N_1381,In_2014);
or U2323 (N_2323,In_3615,In_551);
nor U2324 (N_2324,N_1520,In_2872);
and U2325 (N_2325,In_374,N_1504);
and U2326 (N_2326,In_739,N_1214);
and U2327 (N_2327,N_884,N_745);
nor U2328 (N_2328,In_4338,N_260);
or U2329 (N_2329,N_1636,In_3634);
or U2330 (N_2330,In_1375,N_654);
nand U2331 (N_2331,In_629,N_1804);
or U2332 (N_2332,In_2480,N_894);
or U2333 (N_2333,In_3725,In_2314);
or U2334 (N_2334,N_902,In_3448);
and U2335 (N_2335,In_227,N_1838);
and U2336 (N_2336,N_1832,N_246);
nor U2337 (N_2337,In_4412,N_1484);
nor U2338 (N_2338,In_4564,In_1235);
and U2339 (N_2339,In_1643,In_778);
and U2340 (N_2340,In_1013,N_1934);
nor U2341 (N_2341,In_4252,In_969);
and U2342 (N_2342,In_2503,N_1085);
or U2343 (N_2343,In_3033,N_1416);
and U2344 (N_2344,N_1404,N_1143);
xor U2345 (N_2345,N_1928,N_1744);
and U2346 (N_2346,In_4799,N_1194);
nand U2347 (N_2347,In_2677,In_3957);
nand U2348 (N_2348,N_1533,N_1038);
xnor U2349 (N_2349,In_1342,N_18);
or U2350 (N_2350,N_1950,In_437);
or U2351 (N_2351,In_2199,N_1471);
or U2352 (N_2352,N_1352,In_3972);
or U2353 (N_2353,In_2331,In_3349);
nor U2354 (N_2354,In_2097,N_1255);
nand U2355 (N_2355,N_1681,In_980);
nor U2356 (N_2356,N_1507,In_708);
xor U2357 (N_2357,N_1792,In_3838);
or U2358 (N_2358,N_1562,In_1256);
nand U2359 (N_2359,In_760,N_968);
or U2360 (N_2360,In_2981,In_1258);
or U2361 (N_2361,In_4757,N_421);
nand U2362 (N_2362,N_1470,In_3829);
or U2363 (N_2363,In_1738,In_3139);
xnor U2364 (N_2364,N_1093,In_3280);
nand U2365 (N_2365,In_2285,N_1432);
xnor U2366 (N_2366,In_4211,In_4326);
nand U2367 (N_2367,In_2757,N_1167);
and U2368 (N_2368,In_1556,In_3981);
and U2369 (N_2369,In_3200,In_4181);
xor U2370 (N_2370,N_985,In_2016);
xor U2371 (N_2371,N_1480,In_3274);
xor U2372 (N_2372,In_127,N_709);
or U2373 (N_2373,N_572,In_4702);
xor U2374 (N_2374,In_982,In_947);
xnor U2375 (N_2375,In_3427,In_19);
nor U2376 (N_2376,In_3664,In_3895);
nor U2377 (N_2377,N_157,N_1061);
nand U2378 (N_2378,In_4739,In_2895);
nand U2379 (N_2379,N_70,In_2369);
and U2380 (N_2380,N_380,In_3137);
nand U2381 (N_2381,N_1657,In_528);
nand U2382 (N_2382,N_1252,N_729);
xor U2383 (N_2383,N_1743,In_900);
or U2384 (N_2384,N_1068,In_1008);
nand U2385 (N_2385,In_2672,N_1691);
xor U2386 (N_2386,N_1059,N_1655);
xnor U2387 (N_2387,In_2561,In_3185);
or U2388 (N_2388,N_1168,N_1728);
nor U2389 (N_2389,N_1567,N_1546);
xor U2390 (N_2390,In_892,N_1988);
or U2391 (N_2391,N_1787,In_4147);
xnor U2392 (N_2392,N_91,N_288);
nand U2393 (N_2393,In_1023,In_3776);
xnor U2394 (N_2394,In_318,In_272);
and U2395 (N_2395,In_315,N_1452);
and U2396 (N_2396,In_2182,In_685);
or U2397 (N_2397,In_2389,In_4871);
xor U2398 (N_2398,In_3313,In_1068);
xnor U2399 (N_2399,In_209,In_3212);
nor U2400 (N_2400,N_973,N_1400);
or U2401 (N_2401,In_299,In_1284);
xor U2402 (N_2402,In_1120,N_621);
nand U2403 (N_2403,In_1000,In_1500);
or U2404 (N_2404,In_1928,In_3413);
nand U2405 (N_2405,In_3186,N_845);
or U2406 (N_2406,N_1545,In_263);
nor U2407 (N_2407,N_569,N_610);
nor U2408 (N_2408,N_1721,N_1956);
nor U2409 (N_2409,In_4957,In_4642);
nand U2410 (N_2410,N_551,In_523);
nor U2411 (N_2411,In_3806,In_4216);
nand U2412 (N_2412,In_4500,N_1002);
and U2413 (N_2413,N_1287,In_2610);
xor U2414 (N_2414,In_3766,In_337);
nor U2415 (N_2415,N_1462,N_993);
nor U2416 (N_2416,N_1855,In_3142);
or U2417 (N_2417,N_1276,N_778);
nor U2418 (N_2418,N_1906,N_1512);
or U2419 (N_2419,In_4381,In_4719);
xnor U2420 (N_2420,N_1461,N_1369);
or U2421 (N_2421,In_3921,In_503);
xor U2422 (N_2422,In_2455,In_1042);
xor U2423 (N_2423,In_671,In_2567);
xor U2424 (N_2424,In_4919,N_48);
nor U2425 (N_2425,N_297,In_868);
or U2426 (N_2426,In_4901,In_1624);
or U2427 (N_2427,In_145,In_2173);
and U2428 (N_2428,N_1328,In_261);
nand U2429 (N_2429,In_3348,N_493);
or U2430 (N_2430,N_1115,In_4102);
nand U2431 (N_2431,In_596,In_1778);
or U2432 (N_2432,In_2143,N_1299);
nand U2433 (N_2433,In_4236,In_1480);
or U2434 (N_2434,N_1081,N_1138);
or U2435 (N_2435,In_4751,N_1586);
xor U2436 (N_2436,In_4472,In_3809);
nand U2437 (N_2437,N_1775,In_3535);
nand U2438 (N_2438,In_918,In_42);
nand U2439 (N_2439,N_1560,In_4867);
xor U2440 (N_2440,In_2676,N_1915);
xnor U2441 (N_2441,N_1584,In_1218);
xnor U2442 (N_2442,N_1187,N_1060);
or U2443 (N_2443,N_1179,N_1549);
or U2444 (N_2444,In_4334,In_2306);
or U2445 (N_2445,N_1957,In_3295);
xnor U2446 (N_2446,In_4958,N_1917);
or U2447 (N_2447,In_2769,N_824);
or U2448 (N_2448,In_4016,In_2093);
nand U2449 (N_2449,In_2755,In_2553);
and U2450 (N_2450,N_1623,N_924);
and U2451 (N_2451,In_1584,In_2264);
nor U2452 (N_2452,In_4029,In_1316);
xnor U2453 (N_2453,In_1991,N_550);
nor U2454 (N_2454,In_463,In_4314);
xor U2455 (N_2455,N_1614,In_300);
xnor U2456 (N_2456,In_3471,N_412);
nand U2457 (N_2457,N_339,In_686);
xor U2458 (N_2458,N_1637,N_6);
nand U2459 (N_2459,In_2698,N_981);
xnor U2460 (N_2460,N_1408,In_559);
nand U2461 (N_2461,In_3709,N_547);
nand U2462 (N_2462,N_761,N_1940);
xor U2463 (N_2463,N_304,In_2383);
xor U2464 (N_2464,In_2541,N_1961);
nor U2465 (N_2465,In_1324,N_1182);
and U2466 (N_2466,N_1250,N_1396);
and U2467 (N_2467,N_1534,In_3173);
and U2468 (N_2468,In_1659,In_194);
xnor U2469 (N_2469,N_90,N_1112);
or U2470 (N_2470,N_1949,In_917);
xor U2471 (N_2471,N_1913,In_3098);
or U2472 (N_2472,N_580,In_1697);
or U2473 (N_2473,In_4759,N_1040);
nor U2474 (N_2474,In_3929,In_2105);
nand U2475 (N_2475,In_1633,In_922);
nand U2476 (N_2476,In_4040,In_1335);
and U2477 (N_2477,N_789,In_1977);
nand U2478 (N_2478,In_3421,N_1391);
and U2479 (N_2479,N_1634,N_1870);
nor U2480 (N_2480,In_1093,In_1724);
and U2481 (N_2481,N_1135,In_465);
or U2482 (N_2482,N_1082,In_2137);
and U2483 (N_2483,In_815,In_4088);
nand U2484 (N_2484,N_303,N_1590);
xnor U2485 (N_2485,In_2721,In_367);
or U2486 (N_2486,In_3366,In_3791);
or U2487 (N_2487,N_1196,In_767);
and U2488 (N_2488,In_222,In_476);
nor U2489 (N_2489,In_738,In_2378);
nand U2490 (N_2490,N_577,N_864);
nand U2491 (N_2491,N_1711,In_1394);
xor U2492 (N_2492,In_4875,In_445);
or U2493 (N_2493,In_1341,In_634);
or U2494 (N_2494,In_752,In_3898);
or U2495 (N_2495,N_769,In_3609);
xor U2496 (N_2496,N_1665,In_349);
xor U2497 (N_2497,In_1722,N_1868);
xor U2498 (N_2498,In_1745,In_2060);
nand U2499 (N_2499,N_379,In_1531);
xor U2500 (N_2500,N_1932,N_1976);
nand U2501 (N_2501,N_734,N_358);
and U2502 (N_2502,N_935,In_121);
or U2503 (N_2503,In_1741,In_1180);
or U2504 (N_2504,In_774,N_1422);
or U2505 (N_2505,In_2049,N_2148);
or U2506 (N_2506,N_1602,In_3690);
or U2507 (N_2507,N_2042,In_3259);
and U2508 (N_2508,N_1552,N_1872);
xnor U2509 (N_2509,N_271,In_2135);
nor U2510 (N_2510,In_731,N_674);
nor U2511 (N_2511,N_2192,N_1283);
or U2512 (N_2512,In_1273,In_599);
nor U2513 (N_2513,N_892,N_898);
nand U2514 (N_2514,In_2031,In_4986);
xor U2515 (N_2515,N_1736,N_1377);
nor U2516 (N_2516,N_1817,In_1972);
and U2517 (N_2517,N_1474,N_1437);
and U2518 (N_2518,N_681,In_83);
and U2519 (N_2519,In_682,N_1385);
or U2520 (N_2520,N_1850,In_3086);
and U2521 (N_2521,In_2099,N_77);
nand U2522 (N_2522,N_1075,N_2210);
nor U2523 (N_2523,N_2415,In_1132);
and U2524 (N_2524,N_116,In_79);
and U2525 (N_2525,In_3940,In_459);
nand U2526 (N_2526,N_1049,In_1918);
nand U2527 (N_2527,N_159,N_793);
xnor U2528 (N_2528,In_3819,N_2052);
or U2529 (N_2529,In_3777,In_371);
or U2530 (N_2530,N_2454,N_456);
and U2531 (N_2531,N_951,In_3694);
xor U2532 (N_2532,N_1177,In_228);
and U2533 (N_2533,N_1465,N_2170);
xor U2534 (N_2534,In_259,In_2830);
and U2535 (N_2535,In_676,In_1329);
and U2536 (N_2536,N_1531,In_3900);
and U2537 (N_2537,In_4810,N_2110);
xor U2538 (N_2538,In_3258,N_1506);
and U2539 (N_2539,In_3441,N_2005);
and U2540 (N_2540,In_1868,In_2362);
or U2541 (N_2541,In_2140,In_4522);
xnor U2542 (N_2542,N_2402,N_1420);
and U2543 (N_2543,In_2700,N_2290);
nor U2544 (N_2544,In_1812,In_2883);
and U2545 (N_2545,N_1811,N_617);
xor U2546 (N_2546,In_3469,In_1489);
nor U2547 (N_2547,N_2251,In_3710);
nand U2548 (N_2548,In_3275,N_1682);
nand U2549 (N_2549,N_1559,N_2185);
or U2550 (N_2550,In_208,In_340);
nand U2551 (N_2551,N_1735,N_1532);
xnor U2552 (N_2552,In_2492,In_1752);
xnor U2553 (N_2553,N_815,In_570);
nand U2554 (N_2554,In_2821,N_80);
xnor U2555 (N_2555,N_1689,N_1326);
and U2556 (N_2556,In_2078,N_1159);
and U2557 (N_2557,N_2464,In_2681);
nand U2558 (N_2558,In_41,In_2191);
and U2559 (N_2559,In_1310,N_2419);
or U2560 (N_2560,In_726,N_2453);
nor U2561 (N_2561,N_2456,N_2470);
xnor U2562 (N_2562,In_136,N_2315);
or U2563 (N_2563,N_1827,In_3235);
nor U2564 (N_2564,N_865,In_598);
nor U2565 (N_2565,In_2051,N_1426);
nor U2566 (N_2566,N_1527,In_2514);
nor U2567 (N_2567,N_791,N_2428);
and U2568 (N_2568,N_1820,In_1828);
xnor U2569 (N_2569,N_2476,In_1831);
or U2570 (N_2570,N_678,In_4802);
and U2571 (N_2571,In_3817,In_489);
nand U2572 (N_2572,In_4672,In_4716);
nand U2573 (N_2573,N_363,N_1685);
and U2574 (N_2574,In_1650,N_2314);
nand U2575 (N_2575,N_1070,In_4792);
or U2576 (N_2576,N_2141,N_2418);
and U2577 (N_2577,N_2171,In_4431);
nand U2578 (N_2578,N_1289,N_1812);
xor U2579 (N_2579,In_220,N_1742);
xnor U2580 (N_2580,In_2630,N_1669);
or U2581 (N_2581,N_1350,N_900);
xor U2582 (N_2582,In_525,N_1783);
and U2583 (N_2583,N_1013,In_2342);
nand U2584 (N_2584,In_4182,N_744);
or U2585 (N_2585,In_2743,N_1440);
and U2586 (N_2586,In_117,In_3040);
nand U2587 (N_2587,In_36,In_3072);
or U2588 (N_2588,N_529,N_1557);
nand U2589 (N_2589,In_2335,In_3143);
nor U2590 (N_2590,N_988,In_1601);
nor U2591 (N_2591,In_780,In_3577);
xnor U2592 (N_2592,In_3164,In_4554);
nor U2593 (N_2593,In_142,In_3834);
xor U2594 (N_2594,In_2950,In_2912);
and U2595 (N_2595,N_2002,N_1319);
nor U2596 (N_2596,N_1128,N_2274);
nand U2597 (N_2597,N_2443,N_740);
nand U2598 (N_2598,N_582,N_2392);
nor U2599 (N_2599,N_1828,In_1145);
and U2600 (N_2600,In_1423,In_1863);
nor U2601 (N_2601,In_4845,N_2047);
xnor U2602 (N_2602,N_541,N_2487);
or U2603 (N_2603,In_3167,In_1083);
or U2604 (N_2604,In_3991,In_3532);
nor U2605 (N_2605,N_26,N_2126);
xor U2606 (N_2606,N_2468,In_2);
and U2607 (N_2607,N_2012,N_1815);
nor U2608 (N_2608,In_630,N_1336);
xor U2609 (N_2609,N_2118,In_4199);
xor U2610 (N_2610,In_382,N_1673);
nor U2611 (N_2611,N_1903,N_1476);
xnor U2612 (N_2612,N_2383,N_2205);
and U2613 (N_2613,In_22,In_793);
xor U2614 (N_2614,In_3986,N_946);
nand U2615 (N_2615,In_513,N_1646);
nor U2616 (N_2616,N_685,N_923);
nor U2617 (N_2617,N_59,N_2343);
or U2618 (N_2618,N_2271,In_16);
nand U2619 (N_2619,N_1099,In_4498);
nand U2620 (N_2620,In_968,N_262);
nand U2621 (N_2621,N_2050,In_4894);
nand U2622 (N_2622,In_1804,N_2153);
and U2623 (N_2623,N_2112,In_3715);
and U2624 (N_2624,In_175,N_2370);
and U2625 (N_2625,N_2029,N_591);
nor U2626 (N_2626,N_1951,In_1593);
nand U2627 (N_2627,In_939,N_703);
nand U2628 (N_2628,N_2129,N_2480);
and U2629 (N_2629,N_1927,N_1967);
xor U2630 (N_2630,N_1786,N_2082);
nand U2631 (N_2631,N_2200,N_1197);
nor U2632 (N_2632,N_1145,In_4550);
nor U2633 (N_2633,N_1813,N_2373);
xnor U2634 (N_2634,In_2970,In_737);
nand U2635 (N_2635,In_277,N_1414);
nand U2636 (N_2636,In_4319,In_130);
or U2637 (N_2637,N_1931,In_733);
or U2638 (N_2638,In_4811,In_869);
nand U2639 (N_2639,N_1178,N_2224);
nand U2640 (N_2640,In_2512,In_2427);
nor U2641 (N_2641,In_2719,N_2337);
nor U2642 (N_2642,N_2320,In_3325);
or U2643 (N_2643,In_839,N_408);
nor U2644 (N_2644,N_111,In_3600);
xor U2645 (N_2645,N_974,In_3435);
xnor U2646 (N_2646,In_3822,In_2975);
xnor U2647 (N_2647,In_2462,N_954);
xor U2648 (N_2648,In_4527,N_1519);
nor U2649 (N_2649,In_3221,In_890);
xnor U2650 (N_2650,N_671,In_4670);
nand U2651 (N_2651,In_2511,N_2387);
or U2652 (N_2652,N_1150,In_3278);
and U2653 (N_2653,In_3757,N_1136);
or U2654 (N_2654,In_1168,In_1875);
and U2655 (N_2655,N_2382,N_771);
nor U2656 (N_2656,In_1292,In_4510);
nor U2657 (N_2657,In_3585,In_56);
and U2658 (N_2658,In_2138,N_1445);
nor U2659 (N_2659,N_544,In_4204);
nand U2660 (N_2660,N_504,In_828);
and U2661 (N_2661,In_2352,In_2733);
and U2662 (N_2662,N_2179,In_1143);
xor U2663 (N_2663,N_553,In_2498);
or U2664 (N_2664,N_2003,In_449);
nor U2665 (N_2665,N_1310,N_1139);
and U2666 (N_2666,In_703,In_4276);
xnor U2667 (N_2667,In_4839,In_1477);
nand U2668 (N_2668,In_4849,In_3702);
nand U2669 (N_2669,N_2474,N_760);
and U2670 (N_2670,N_1510,In_3700);
nand U2671 (N_2671,N_2360,N_1684);
or U2672 (N_2672,In_2845,In_628);
or U2673 (N_2673,N_75,In_1269);
xnor U2674 (N_2674,In_1012,In_3395);
nor U2675 (N_2675,In_4814,In_2674);
and U2676 (N_2676,N_2368,N_2086);
nor U2677 (N_2677,In_3265,In_905);
xnor U2678 (N_2678,N_632,N_1727);
and U2679 (N_2679,In_1958,N_2070);
nand U2680 (N_2680,N_1036,N_434);
xor U2681 (N_2681,N_1834,N_1164);
xor U2682 (N_2682,N_574,N_291);
nand U2683 (N_2683,N_1282,N_356);
nor U2684 (N_2684,In_4304,In_955);
or U2685 (N_2685,N_1576,In_1965);
nand U2686 (N_2686,In_3613,In_4627);
nor U2687 (N_2687,N_982,N_1842);
nor U2688 (N_2688,N_2049,N_2242);
nand U2689 (N_2689,In_3964,In_4704);
and U2690 (N_2690,In_1554,N_2364);
and U2691 (N_2691,N_1668,N_1537);
xor U2692 (N_2692,N_1464,In_3718);
xor U2693 (N_2693,N_2424,In_4122);
nor U2694 (N_2694,N_2075,In_1009);
or U2695 (N_2695,N_1330,N_1959);
and U2696 (N_2696,In_1576,N_2013);
xor U2697 (N_2697,N_1312,N_2444);
nand U2698 (N_2698,N_2194,N_206);
xor U2699 (N_2699,N_2007,In_1772);
nand U2700 (N_2700,N_1608,N_1877);
nand U2701 (N_2701,N_1536,In_4041);
and U2702 (N_2702,N_1256,In_2572);
xor U2703 (N_2703,In_2540,N_2262);
nor U2704 (N_2704,In_2094,N_489);
nor U2705 (N_2705,N_1111,In_2291);
nor U2706 (N_2706,N_2056,In_811);
or U2707 (N_2707,N_1148,In_3000);
nor U2708 (N_2708,N_1288,In_2167);
and U2709 (N_2709,In_2705,N_431);
nand U2710 (N_2710,N_2134,N_2281);
nand U2711 (N_2711,N_2204,N_1005);
or U2712 (N_2712,N_2258,N_2491);
and U2713 (N_2713,N_2018,N_1937);
nor U2714 (N_2714,In_392,In_4465);
and U2715 (N_2715,In_1446,N_2305);
nor U2716 (N_2716,In_2013,In_1165);
nor U2717 (N_2717,N_1980,N_1710);
nand U2718 (N_2718,N_2132,N_2109);
xnor U2719 (N_2719,In_4366,N_1955);
nand U2720 (N_2720,In_4925,N_1597);
nor U2721 (N_2721,In_2377,N_2240);
and U2722 (N_2722,In_2574,In_3505);
nand U2723 (N_2723,N_950,In_2888);
nor U2724 (N_2724,N_2278,In_3954);
xor U2725 (N_2725,N_1641,N_1859);
nand U2726 (N_2726,N_2460,N_1705);
xor U2727 (N_2727,In_2322,N_505);
nand U2728 (N_2728,In_120,In_2409);
and U2729 (N_2729,N_2199,In_929);
xnor U2730 (N_2730,In_3104,N_2131);
xnor U2731 (N_2731,N_1122,N_1297);
nor U2732 (N_2732,N_1718,In_2219);
xnor U2733 (N_2733,In_4303,N_1610);
xnor U2734 (N_2734,In_3394,N_2025);
or U2735 (N_2735,N_1071,In_3400);
nand U2736 (N_2736,In_3302,In_3114);
and U2737 (N_2737,In_1684,N_1836);
nand U2738 (N_2738,N_1242,N_1063);
xor U2739 (N_2739,In_2683,N_2429);
or U2740 (N_2740,N_2405,In_1798);
or U2741 (N_2741,In_1065,N_1284);
nand U2742 (N_2742,In_3466,N_1535);
nand U2743 (N_2743,In_3608,In_1517);
or U2744 (N_2744,In_1147,N_2340);
xor U2745 (N_2745,In_827,N_916);
xnor U2746 (N_2746,N_2114,N_1102);
nor U2747 (N_2747,N_2485,In_4978);
xnor U2748 (N_2748,N_1611,In_3256);
nand U2749 (N_2749,In_3027,N_1185);
xor U2750 (N_2750,In_4697,N_1569);
or U2751 (N_2751,In_1982,N_2459);
or U2752 (N_2752,N_2441,N_1848);
nand U2753 (N_2753,N_1342,In_4880);
nand U2754 (N_2754,N_2111,N_301);
xor U2755 (N_2755,N_87,N_2053);
nand U2756 (N_2756,N_2285,In_2548);
and U2757 (N_2757,In_1522,In_2828);
nor U2758 (N_2758,N_2223,N_2482);
nor U2759 (N_2759,N_2071,N_774);
or U2760 (N_2760,In_894,In_3545);
xnor U2761 (N_2761,N_2202,In_3627);
nand U2762 (N_2762,N_1517,In_4921);
nand U2763 (N_2763,In_2340,In_3784);
or U2764 (N_2764,N_136,N_2302);
nor U2765 (N_2765,N_1973,N_1490);
xor U2766 (N_2766,In_376,N_221);
nor U2767 (N_2767,N_928,N_1747);
nand U2768 (N_2768,In_4928,N_2297);
nor U2769 (N_2769,In_3355,In_3754);
nand U2770 (N_2770,N_1688,N_1293);
and U2771 (N_2771,N_2073,In_4121);
nand U2772 (N_2772,In_4296,N_1942);
nand U2773 (N_2773,In_1319,In_3951);
and U2774 (N_2774,In_813,N_401);
nor U2775 (N_2775,N_1593,In_1671);
or U2776 (N_2776,In_4705,N_236);
nor U2777 (N_2777,N_338,In_2121);
nor U2778 (N_2778,N_558,N_702);
or U2779 (N_2779,In_935,N_1591);
or U2780 (N_2780,In_4390,In_1969);
or U2781 (N_2781,In_4058,N_2417);
and U2782 (N_2782,N_967,In_1475);
nor U2783 (N_2783,In_2767,In_775);
nor U2784 (N_2784,N_1788,In_1498);
or U2785 (N_2785,In_4111,In_2740);
nand U2786 (N_2786,N_2061,N_2184);
nor U2787 (N_2787,N_2275,N_1982);
nor U2788 (N_2788,In_3264,N_2490);
and U2789 (N_2789,N_2400,N_1048);
and U2790 (N_2790,N_2433,In_2741);
nand U2791 (N_2791,N_2335,N_1488);
and U2792 (N_2792,N_2180,In_782);
and U2793 (N_2793,N_1618,In_3583);
nor U2794 (N_2794,N_2083,In_1604);
or U2795 (N_2795,In_3753,In_360);
xor U2796 (N_2796,In_2252,N_1043);
nand U2797 (N_2797,N_2458,N_1384);
nand U2798 (N_2798,In_2017,In_2616);
nand U2799 (N_2799,N_2181,N_2467);
and U2800 (N_2800,N_1421,N_962);
nor U2801 (N_2801,N_846,N_796);
and U2802 (N_2802,N_1251,In_901);
nand U2803 (N_2803,In_669,In_3240);
nor U2804 (N_2804,N_1809,In_1359);
nand U2805 (N_2805,N_1676,N_1644);
nor U2806 (N_2806,In_62,N_748);
or U2807 (N_2807,In_2993,In_2526);
or U2808 (N_2808,N_561,N_1741);
nor U2809 (N_2809,In_4308,N_1006);
xnor U2810 (N_2810,In_1225,N_2272);
and U2811 (N_2811,In_965,N_797);
nand U2812 (N_2812,N_662,In_1727);
nor U2813 (N_2813,In_749,N_2312);
nand U2814 (N_2814,In_1960,N_205);
or U2815 (N_2815,In_1585,N_2322);
xor U2816 (N_2816,In_1254,N_858);
xnor U2817 (N_2817,N_2218,N_515);
nand U2818 (N_2818,In_3080,In_1915);
and U2819 (N_2819,N_1702,In_1691);
nand U2820 (N_2820,In_4788,In_251);
xor U2821 (N_2821,N_2239,N_2475);
nand U2822 (N_2822,N_1021,N_1321);
nand U2823 (N_2823,N_2156,N_1311);
or U2824 (N_2824,In_131,In_441);
nor U2825 (N_2825,N_1062,In_3025);
nand U2826 (N_2826,In_1866,In_1550);
or U2827 (N_2827,N_2051,In_414);
or U2828 (N_2828,In_2573,In_4971);
or U2829 (N_2829,In_3554,N_2066);
nor U2830 (N_2830,N_2024,In_4400);
nor U2831 (N_2831,N_1583,In_1583);
and U2832 (N_2832,N_284,In_4240);
xnor U2833 (N_2833,In_3728,N_1837);
and U2834 (N_2834,N_2463,In_1857);
nand U2835 (N_2835,N_374,In_2446);
nand U2836 (N_2836,N_788,In_1846);
or U2837 (N_2837,In_3381,In_2549);
xnor U2838 (N_2838,In_2779,N_2398);
and U2839 (N_2839,N_2139,N_2032);
nor U2840 (N_2840,In_1924,N_997);
or U2841 (N_2841,In_6,N_2498);
or U2842 (N_2842,In_4095,In_4707);
nor U2843 (N_2843,In_2171,N_460);
or U2844 (N_2844,N_188,N_636);
or U2845 (N_2845,In_985,In_3756);
or U2846 (N_2846,N_1588,N_613);
or U2847 (N_2847,In_1176,N_975);
nand U2848 (N_2848,In_754,N_1757);
nand U2849 (N_2849,In_2196,In_1032);
nand U2850 (N_2850,In_4885,In_2025);
or U2851 (N_2851,N_1451,In_3744);
or U2852 (N_2852,In_4226,N_2174);
and U2853 (N_2853,N_2284,N_1216);
and U2854 (N_2854,N_1096,N_1672);
or U2855 (N_2855,N_2352,In_4653);
or U2856 (N_2856,In_2785,In_4173);
nand U2857 (N_2857,In_2307,In_3007);
and U2858 (N_2858,In_2395,In_2913);
or U2859 (N_2859,N_2442,In_3518);
xnor U2860 (N_2860,N_557,In_2501);
nor U2861 (N_2861,N_1970,In_4311);
and U2862 (N_2862,N_601,N_1053);
xor U2863 (N_2863,In_0,In_2935);
xor U2864 (N_2864,N_1883,In_4337);
xnor U2865 (N_2865,In_964,N_2206);
nor U2866 (N_2866,In_2684,N_226);
and U2867 (N_2867,In_862,N_1766);
or U2868 (N_2868,N_2306,In_4823);
nor U2869 (N_2869,N_1035,In_821);
nand U2870 (N_2870,In_352,N_2151);
xnor U2871 (N_2871,In_836,N_1511);
and U2872 (N_2872,N_2079,In_313);
xnor U2873 (N_2873,In_2925,In_4597);
and U2874 (N_2874,In_1223,In_2736);
or U2875 (N_2875,In_1944,In_4714);
nand U2876 (N_2876,N_2397,In_4067);
nand U2877 (N_2877,In_4224,N_2027);
xnor U2878 (N_2878,In_2623,In_4022);
nor U2879 (N_2879,In_3926,N_2481);
xor U2880 (N_2880,In_4833,In_257);
xor U2881 (N_2881,In_4812,In_2936);
or U2882 (N_2882,In_659,In_3849);
xor U2883 (N_2883,In_4725,N_659);
nor U2884 (N_2884,In_1075,N_2155);
and U2885 (N_2885,N_2040,In_4640);
nand U2886 (N_2886,N_2336,N_495);
nand U2887 (N_2887,In_2804,N_1554);
and U2888 (N_2888,In_101,In_1558);
nand U2889 (N_2889,In_1651,In_3633);
xor U2890 (N_2890,N_2231,In_478);
nand U2891 (N_2891,In_1197,N_2465);
nand U2892 (N_2892,N_1259,N_168);
nand U2893 (N_2893,N_984,In_2439);
nand U2894 (N_2894,In_897,N_2144);
and U2895 (N_2895,In_2106,N_777);
and U2896 (N_2896,In_81,N_2282);
or U2897 (N_2897,N_1494,N_1026);
or U2898 (N_2898,N_1524,In_1227);
and U2899 (N_2899,In_957,N_1659);
nand U2900 (N_2900,N_1652,N_1028);
and U2901 (N_2901,N_2455,In_4264);
xnor U2902 (N_2902,In_909,N_1638);
nand U2903 (N_2903,In_4288,N_2229);
or U2904 (N_2904,N_2421,N_1654);
nand U2905 (N_2905,In_3091,N_687);
and U2906 (N_2906,In_3241,In_2750);
and U2907 (N_2907,N_2380,N_2201);
and U2908 (N_2908,In_4783,In_2670);
and U2909 (N_2909,N_1472,In_2320);
nand U2910 (N_2910,In_2354,N_2190);
and U2911 (N_2911,N_1007,N_886);
and U2912 (N_2912,N_2308,In_2386);
and U2913 (N_2913,In_2565,N_413);
xnor U2914 (N_2914,In_1937,N_1908);
nand U2915 (N_2915,In_4622,N_1530);
nor U2916 (N_2916,N_2063,In_3565);
xor U2917 (N_2917,N_143,N_1892);
xnor U2918 (N_2918,In_4114,N_290);
and U2919 (N_2919,N_1268,N_1723);
nand U2920 (N_2920,In_401,N_1962);
nor U2921 (N_2921,N_948,N_399);
or U2922 (N_2922,N_2104,N_1355);
nor U2923 (N_2923,In_1900,In_3905);
and U2924 (N_2924,N_921,N_1840);
or U2925 (N_2925,In_959,N_600);
or U2926 (N_2926,In_4798,In_4001);
or U2927 (N_2927,N_261,N_2477);
nor U2928 (N_2928,N_1825,N_2425);
nor U2929 (N_2929,N_1004,N_2168);
and U2930 (N_2930,N_2401,N_1846);
xnor U2931 (N_2931,N_564,N_1737);
xnor U2932 (N_2932,In_553,N_32);
and U2933 (N_2933,In_2380,In_2216);
and U2934 (N_2934,N_2203,In_1407);
nor U2935 (N_2935,In_4857,In_4372);
nor U2936 (N_2936,N_2021,N_1393);
xnor U2937 (N_2937,In_2405,In_3974);
or U2938 (N_2938,N_149,In_2863);
or U2939 (N_2939,N_2145,N_1371);
nand U2940 (N_2940,In_2566,In_790);
and U2941 (N_2941,N_2341,N_850);
nor U2942 (N_2942,In_4169,In_4066);
xor U2943 (N_2943,In_2742,N_1645);
nand U2944 (N_2944,In_1518,N_2296);
and U2945 (N_2945,In_4990,N_1265);
and U2946 (N_2946,In_3157,N_2321);
nor U2947 (N_2947,N_1607,N_1285);
xnor U2948 (N_2948,In_2254,N_1189);
xor U2949 (N_2949,N_1486,N_2198);
xor U2950 (N_2950,In_3131,In_3472);
nand U2951 (N_2951,In_3978,N_2093);
and U2952 (N_2952,N_2259,N_29);
xnor U2953 (N_2953,N_1542,N_786);
nand U2954 (N_2954,In_1287,N_2331);
or U2955 (N_2955,In_1827,In_1503);
and U2956 (N_2956,N_2090,N_164);
and U2957 (N_2957,N_2493,In_1713);
nor U2958 (N_2958,N_1734,In_3561);
or U2959 (N_2959,N_2076,In_2780);
or U2960 (N_2960,N_1761,N_821);
nand U2961 (N_2961,In_3944,In_1243);
or U2962 (N_2962,N_2230,N_641);
nor U2963 (N_2963,N_1353,N_158);
nor U2964 (N_2964,N_2017,In_2141);
nor U2965 (N_2965,N_1226,N_1972);
or U2966 (N_2966,N_258,N_1824);
nand U2967 (N_2967,N_2430,N_2000);
nand U2968 (N_2968,N_1110,In_637);
or U2969 (N_2969,N_2133,In_2904);
nor U2970 (N_2970,N_2318,N_1475);
or U2971 (N_2971,N_169,In_626);
and U2972 (N_2972,In_514,N_2457);
nand U2973 (N_2973,In_4340,In_710);
xor U2974 (N_2974,N_1819,In_2518);
xor U2975 (N_2975,In_190,N_1210);
or U2976 (N_2976,In_3095,N_2396);
xor U2977 (N_2977,N_2222,N_1904);
xnor U2978 (N_2978,N_1616,N_1966);
and U2979 (N_2979,In_1020,In_3227);
or U2980 (N_2980,In_2180,In_3403);
nand U2981 (N_2981,N_2127,N_2207);
nand U2982 (N_2982,In_1682,N_1749);
or U2983 (N_2983,N_1269,N_1667);
xnor U2984 (N_2984,N_1900,In_3036);
and U2985 (N_2985,In_3908,In_1362);
nand U2986 (N_2986,In_2128,N_1411);
xnor U2987 (N_2987,N_283,N_2328);
nor U2988 (N_2988,In_4793,N_1412);
nor U2989 (N_2989,In_4365,N_2123);
and U2990 (N_2990,N_1032,N_1664);
nor U2991 (N_2991,In_3999,In_2000);
and U2992 (N_2992,N_2374,N_1625);
and U2993 (N_2993,N_1117,N_2478);
or U2994 (N_2994,In_1318,In_4909);
nand U2995 (N_2995,N_2057,In_2607);
nor U2996 (N_2996,N_1209,In_3840);
nand U2997 (N_2997,N_1939,N_2089);
nand U2998 (N_2998,In_1546,In_1460);
nand U2999 (N_2999,N_2310,In_3528);
nand U3000 (N_3000,In_2262,In_4413);
nand U3001 (N_3001,N_1753,In_1708);
nor U3002 (N_3002,N_100,N_2416);
or U3003 (N_3003,N_2813,In_761);
xnor U3004 (N_3004,In_4591,N_2764);
nand U3005 (N_3005,N_2573,In_1748);
or U3006 (N_3006,N_2937,N_1814);
nor U3007 (N_3007,In_2885,N_2981);
and U3008 (N_3008,N_2640,N_2072);
nor U3009 (N_3009,N_782,In_3787);
and U3010 (N_3010,N_2232,N_704);
nor U3011 (N_3011,In_3591,N_2754);
or U3012 (N_3012,N_1064,N_2685);
and U3013 (N_3013,N_987,In_3026);
and U3014 (N_3014,N_1436,N_2559);
nor U3015 (N_3015,In_3180,N_1419);
nor U3016 (N_3016,N_2503,N_1899);
and U3017 (N_3017,N_2747,N_2681);
nor U3018 (N_3018,N_1990,N_1298);
or U3019 (N_3019,N_2868,N_2752);
nand U3020 (N_3020,N_2096,N_2953);
and U3021 (N_3021,In_3454,In_2967);
nand U3022 (N_3022,In_4227,In_2006);
or U3023 (N_3023,In_3297,N_309);
and U3024 (N_3024,N_1303,N_2510);
or U3025 (N_3025,In_187,In_1141);
or U3026 (N_3026,N_1606,N_2817);
nand U3027 (N_3027,N_686,N_2875);
nor U3028 (N_3028,N_2346,N_428);
nand U3029 (N_3029,N_34,In_2281);
nand U3030 (N_3030,N_2988,N_2711);
or U3031 (N_3031,N_1598,In_4706);
nand U3032 (N_3032,N_2969,N_2639);
or U3033 (N_3033,N_361,N_647);
nand U3034 (N_3034,N_2803,In_1464);
xnor U3035 (N_3035,N_2515,N_2578);
or U3036 (N_3036,N_2483,In_656);
or U3037 (N_3037,N_2116,In_1559);
nand U3038 (N_3038,In_1209,N_2411);
xnor U3039 (N_3039,N_2246,In_3975);
xnor U3040 (N_3040,In_4096,N_2497);
xnor U3041 (N_3041,N_2786,N_2934);
nor U3042 (N_3042,N_1525,In_4846);
nand U3043 (N_3043,In_4721,N_1341);
and U3044 (N_3044,N_2489,N_739);
or U3045 (N_3045,N_2792,In_3397);
or U3046 (N_3046,N_2805,In_3195);
and U3047 (N_3047,N_1995,N_1253);
or U3048 (N_3048,N_2479,N_1017);
and U3049 (N_3049,N_31,In_3949);
or U3050 (N_3050,In_3223,N_2697);
nand U3051 (N_3051,In_268,N_233);
nor U3052 (N_3052,In_158,N_1865);
nor U3053 (N_3053,In_4515,N_839);
xnor U3054 (N_3054,N_2548,N_2924);
and U3055 (N_3055,In_4490,In_241);
nor U3056 (N_3056,N_609,N_2931);
and U3057 (N_3057,N_1374,In_1737);
xor U3058 (N_3058,N_1544,N_2579);
and U3059 (N_3059,N_2267,In_2469);
nand U3060 (N_3060,N_2004,N_2469);
nand U3061 (N_3061,N_2986,N_1221);
xnor U3062 (N_3062,In_1193,In_1177);
nor U3063 (N_3063,N_2595,In_1248);
nand U3064 (N_3064,In_4180,In_4505);
and U3065 (N_3065,N_1041,N_1627);
xor U3066 (N_3066,N_1463,In_886);
xnor U3067 (N_3067,In_1819,In_4816);
nor U3068 (N_3068,N_2591,N_1523);
nand U3069 (N_3069,N_257,N_2495);
or U3070 (N_3070,In_2675,N_286);
nor U3071 (N_3071,N_2552,In_3430);
nor U3072 (N_3072,N_1789,In_2075);
nor U3073 (N_3073,In_3814,N_1010);
nor U3074 (N_3074,In_1374,N_341);
and U3075 (N_3075,N_2843,N_2266);
nor U3076 (N_3076,In_4943,N_2705);
nand U3077 (N_3077,N_2545,N_897);
nor U3078 (N_3078,N_2678,In_1664);
or U3079 (N_3079,N_2265,In_1376);
xnor U3080 (N_3080,N_2193,N_2991);
nor U3081 (N_3081,N_1351,N_1074);
nor U3082 (N_3082,N_1543,N_2968);
and U3083 (N_3083,N_2794,In_4179);
or U3084 (N_3084,N_2543,N_1261);
nand U3085 (N_3085,N_2703,N_2856);
xnor U3086 (N_3086,N_2757,In_904);
nand U3087 (N_3087,N_1453,N_2734);
and U3088 (N_3088,N_1540,In_1321);
and U3089 (N_3089,N_1803,N_2500);
or U3090 (N_3090,N_2347,N_2877);
or U3091 (N_3091,N_2178,In_3117);
nand U3092 (N_3092,N_2818,N_2238);
nand U3093 (N_3093,N_2149,In_2969);
nand U3094 (N_3094,In_2098,In_1479);
xnor U3095 (N_3095,N_2840,N_2094);
nor U3096 (N_3096,N_2982,N_2546);
or U3097 (N_3097,In_921,In_3404);
xnor U3098 (N_3098,N_2675,N_1799);
xnor U3099 (N_3099,In_4012,N_2219);
nor U3100 (N_3100,In_3943,N_2853);
and U3101 (N_3101,In_4511,In_4106);
or U3102 (N_3102,In_4735,N_1722);
nor U3103 (N_3103,In_1277,N_2121);
xnor U3104 (N_3104,In_1634,N_1496);
nand U3105 (N_3105,In_3205,N_877);
xor U3106 (N_3106,N_2026,N_1387);
nand U3107 (N_3107,N_2157,N_1724);
xor U3108 (N_3108,N_2584,N_2283);
nor U3109 (N_3109,N_2976,N_2790);
nand U3110 (N_3110,N_2288,N_2431);
and U3111 (N_3111,N_934,N_2729);
xnor U3112 (N_3112,N_438,N_2753);
xor U3113 (N_3113,N_2793,N_2227);
nor U3114 (N_3114,In_4770,In_2153);
or U3115 (N_3115,N_1161,N_347);
nor U3116 (N_3116,N_1585,N_2886);
or U3117 (N_3117,N_2531,N_2766);
xnor U3118 (N_3118,In_3772,In_1215);
xnor U3119 (N_3119,In_3804,N_1124);
or U3120 (N_3120,N_1680,N_653);
nand U3121 (N_3121,N_1140,N_1195);
nor U3122 (N_3122,N_2957,N_880);
or U3123 (N_3123,N_1650,In_674);
and U3124 (N_3124,N_2529,N_2164);
nor U3125 (N_3125,In_4937,In_3729);
and U3126 (N_3126,N_2848,N_766);
xnor U3127 (N_3127,N_2329,In_4566);
xor U3128 (N_3128,In_950,N_2623);
nor U3129 (N_3129,N_1409,In_4708);
or U3130 (N_3130,N_1715,In_4401);
or U3131 (N_3131,N_1890,In_4765);
nor U3132 (N_3132,N_2967,In_1261);
or U3133 (N_3133,In_3732,N_2984);
or U3134 (N_3134,N_53,N_2216);
nand U3135 (N_3135,N_1994,In_4960);
xnor U3136 (N_3136,N_642,N_1647);
nand U3137 (N_3137,N_2189,In_166);
nand U3138 (N_3138,N_1762,N_1037);
nand U3139 (N_3139,In_4698,N_2);
or U3140 (N_3140,In_532,N_2146);
nand U3141 (N_3141,N_1670,N_2270);
and U3142 (N_3142,N_2728,N_2620);
xor U3143 (N_3143,N_2117,In_3856);
nand U3144 (N_3144,N_611,N_2019);
or U3145 (N_3145,N_522,In_2261);
or U3146 (N_3146,N_2801,N_2713);
or U3147 (N_3147,N_1314,N_2008);
nor U3148 (N_3148,In_247,N_532);
or U3149 (N_3149,N_1816,N_2438);
nor U3150 (N_3150,N_1784,N_1561);
xor U3151 (N_3151,N_2324,N_2569);
nor U3152 (N_3152,N_2885,N_1095);
nand U3153 (N_3153,N_118,N_2960);
xnor U3154 (N_3154,N_2044,In_1381);
nand U3155 (N_3155,In_1246,N_1349);
nand U3156 (N_3156,In_363,N_239);
xnor U3157 (N_3157,N_1594,In_1984);
xor U3158 (N_3158,N_1797,N_2668);
nor U3159 (N_3159,N_2439,N_2295);
xor U3160 (N_3160,In_3816,In_1625);
nor U3161 (N_3161,In_1001,N_684);
or U3162 (N_3162,N_2850,N_2311);
xor U3163 (N_3163,In_3923,N_2634);
or U3164 (N_3164,In_2976,N_2038);
or U3165 (N_3165,N_2513,N_2892);
nand U3166 (N_3166,N_2137,N_1582);
nor U3167 (N_3167,N_2409,In_3624);
nor U3168 (N_3168,In_2256,N_1778);
or U3169 (N_3169,In_1890,N_2720);
and U3170 (N_3170,N_2159,In_386);
and U3171 (N_3171,N_366,In_1473);
nand U3172 (N_3172,N_1923,N_1097);
nor U3173 (N_3173,In_896,In_1411);
and U3174 (N_3174,In_3064,N_2816);
xor U3175 (N_3175,N_867,N_2700);
nor U3176 (N_3176,N_2248,N_2435);
and U3177 (N_3177,N_2386,N_2619);
nand U3178 (N_3178,In_3651,N_2995);
nand U3179 (N_3179,N_1367,N_2763);
nand U3180 (N_3180,In_3539,In_4341);
nand U3181 (N_3181,In_2076,N_2939);
and U3182 (N_3182,N_1482,N_2600);
or U3183 (N_3183,N_2698,In_406);
xnor U3184 (N_3184,In_140,In_2468);
xnor U3185 (N_3185,In_1372,N_2001);
and U3186 (N_3186,In_3063,N_2601);
nand U3187 (N_3187,In_482,N_1306);
nor U3188 (N_3188,N_2496,N_2158);
and U3189 (N_3189,N_1217,N_2770);
and U3190 (N_3190,N_1651,In_2111);
or U3191 (N_3191,N_2863,In_535);
or U3192 (N_3192,In_928,In_1050);
xnor U3193 (N_3193,In_1378,N_2006);
xor U3194 (N_3194,In_4663,In_1085);
nand U3195 (N_3195,N_1373,N_1280);
nand U3196 (N_3196,In_2373,N_2972);
nand U3197 (N_3197,In_505,N_1394);
nor U3198 (N_3198,N_296,N_2427);
nor U3199 (N_3199,N_683,N_2837);
nand U3200 (N_3200,N_1300,In_1679);
nor U3201 (N_3201,In_4476,N_716);
and U3202 (N_3202,N_2313,N_2388);
or U3203 (N_3203,In_665,N_74);
or U3204 (N_3204,N_2951,In_323);
or U3205 (N_3205,N_650,In_701);
xor U3206 (N_3206,N_2375,N_2944);
and U3207 (N_3207,In_516,N_2881);
or U3208 (N_3208,N_2979,In_4253);
nand U3209 (N_3209,In_519,N_2363);
xnor U3210 (N_3210,In_2184,N_635);
nor U3211 (N_3211,N_780,N_1596);
xnor U3212 (N_3212,N_2606,In_1413);
and U3213 (N_3213,N_2509,In_1769);
nand U3214 (N_3214,N_1791,In_3360);
and U3215 (N_3215,In_2041,In_3894);
nand U3216 (N_3216,In_4395,N_2326);
nor U3217 (N_3217,N_2243,N_2622);
nor U3218 (N_3218,In_3492,N_1924);
nand U3219 (N_3219,In_1897,N_2929);
nand U3220 (N_3220,N_2855,In_2653);
or U3221 (N_3221,N_1212,N_2571);
and U3222 (N_3222,In_2132,N_1822);
and U3223 (N_3223,N_2582,In_1591);
nand U3224 (N_3224,N_2403,In_4979);
nand U3225 (N_3225,N_629,N_2330);
nand U3226 (N_3226,N_2236,N_2554);
or U3227 (N_3227,In_1162,In_653);
and U3228 (N_3228,N_2220,In_2594);
xor U3229 (N_3229,N_2309,N_346);
or U3230 (N_3230,N_238,N_2247);
nor U3231 (N_3231,N_1318,N_1595);
xor U3232 (N_3232,N_1501,N_2099);
or U3233 (N_3233,In_1219,In_3457);
xnor U3234 (N_3234,N_2846,In_978);
and U3235 (N_3235,N_138,In_72);
xnor U3236 (N_3236,N_1910,N_2298);
xor U3237 (N_3237,N_1698,N_2334);
and U3238 (N_3238,N_2390,In_3489);
xnor U3239 (N_3239,In_1539,N_787);
and U3240 (N_3240,N_912,N_2100);
and U3241 (N_3241,In_4593,N_1643);
nand U3242 (N_3242,N_1281,N_2896);
xor U3243 (N_3243,N_1858,N_2921);
nand U3244 (N_3244,N_2605,In_3029);
nor U3245 (N_3245,N_2630,N_2209);
xnor U3246 (N_3246,N_1921,N_2575);
nor U3247 (N_3247,N_1882,N_2484);
nor U3248 (N_3248,N_234,In_4398);
xnor U3249 (N_3249,N_2845,In_1483);
nor U3250 (N_3250,N_1454,N_2750);
nand U3251 (N_3251,In_4056,N_1360);
nor U3252 (N_3252,N_2759,N_2800);
xnor U3253 (N_3253,N_1080,In_4959);
nand U3254 (N_3254,N_287,In_1178);
or U3255 (N_3255,N_2345,N_2521);
xnor U3256 (N_3256,N_1632,In_4188);
nor U3257 (N_3257,N_2799,In_2510);
xnor U3258 (N_3258,In_2983,In_4870);
xor U3259 (N_3259,N_1617,N_2861);
and U3260 (N_3260,In_1826,N_2522);
nor U3261 (N_3261,N_2432,N_2172);
and U3262 (N_3262,N_2974,N_2567);
xnor U3263 (N_3263,In_949,N_1354);
xor U3264 (N_3264,N_2884,In_4535);
nand U3265 (N_3265,N_2665,In_1519);
and U3266 (N_3266,N_466,N_1875);
nand U3267 (N_3267,N_1509,In_4477);
xor U3268 (N_3268,In_605,N_2702);
nor U3269 (N_3269,In_3865,N_1513);
xor U3270 (N_3270,In_824,N_2502);
and U3271 (N_3271,N_2234,N_2609);
nand U3272 (N_3272,In_1279,N_2821);
nand U3273 (N_3273,N_2758,N_1998);
nor U3274 (N_3274,N_1199,N_2617);
nand U3275 (N_3275,N_1592,In_2629);
xor U3276 (N_3276,N_2810,N_2188);
and U3277 (N_3277,N_1566,N_2182);
or U3278 (N_3278,N_1629,N_2844);
nand U3279 (N_3279,N_2723,In_2224);
xor U3280 (N_3280,N_1313,N_2165);
xnor U3281 (N_3281,In_234,N_2046);
nand U3282 (N_3282,N_2880,In_1028);
nor U3283 (N_3283,N_299,N_2412);
xor U3284 (N_3284,N_1565,In_1762);
xor U3285 (N_3285,N_2873,In_2432);
and U3286 (N_3286,N_120,In_3731);
xor U3287 (N_3287,N_2598,N_479);
nand U3288 (N_3288,N_2802,N_736);
and U3289 (N_3289,In_1907,In_1110);
nor U3290 (N_3290,N_1622,In_3357);
nor U3291 (N_3291,N_2244,In_3474);
nand U3292 (N_3292,N_2533,In_888);
or U3293 (N_3293,In_450,In_1700);
nor U3294 (N_3294,N_2699,N_2064);
or U3295 (N_3295,In_114,N_2690);
xor U3296 (N_3296,N_1502,N_2065);
and U3297 (N_3297,N_2852,N_2087);
xor U3298 (N_3298,N_1631,N_1309);
and U3299 (N_3299,N_2532,N_742);
nor U3300 (N_3300,In_1801,In_3656);
nand U3301 (N_3301,N_2916,In_2945);
or U3302 (N_3302,In_2134,N_2900);
and U3303 (N_3303,In_2413,N_2520);
nor U3304 (N_3304,N_2633,N_2876);
xnor U3305 (N_3305,N_2541,N_2214);
xnor U3306 (N_3306,In_2448,N_2451);
nor U3307 (N_3307,N_20,N_2694);
xor U3308 (N_3308,In_3519,N_2492);
xor U3309 (N_3309,N_1378,N_2528);
and U3310 (N_3310,N_1719,In_1247);
nand U3311 (N_3311,N_1952,In_2729);
xnor U3312 (N_3312,In_3296,N_2446);
nor U3313 (N_3313,N_1603,In_470);
xor U3314 (N_3314,N_554,N_2580);
or U3315 (N_3315,N_1731,In_3920);
nor U3316 (N_3316,N_2671,In_2344);
and U3317 (N_3317,N_2908,In_103);
or U3318 (N_3318,N_1492,N_1933);
nor U3319 (N_3319,N_2961,N_2998);
nand U3320 (N_3320,N_227,N_2581);
or U3321 (N_3321,In_4745,In_2490);
xnor U3322 (N_3322,N_1750,N_2627);
nor U3323 (N_3323,N_2536,N_2959);
xor U3324 (N_3324,In_2022,In_4639);
or U3325 (N_3325,N_2695,N_1215);
xor U3326 (N_3326,N_2589,N_2866);
xnor U3327 (N_3327,N_2796,N_228);
nor U3328 (N_3328,N_2196,N_2215);
nand U3329 (N_3329,N_2353,N_1693);
and U3330 (N_3330,In_3860,N_1771);
and U3331 (N_3331,N_2325,In_4590);
or U3332 (N_3332,In_2384,N_2138);
and U3333 (N_3333,N_1874,N_2719);
nand U3334 (N_3334,In_2057,N_2160);
xnor U3335 (N_3335,N_1331,N_746);
nor U3336 (N_3336,In_4468,N_9);
and U3337 (N_3337,N_2461,N_2823);
nor U3338 (N_3338,N_2085,N_2742);
and U3339 (N_3339,N_2925,N_462);
xnor U3340 (N_3340,N_2819,N_2534);
nor U3341 (N_3341,N_524,N_2033);
nand U3342 (N_3342,N_2292,In_2999);
xor U3343 (N_3343,In_3462,In_2425);
or U3344 (N_3344,In_2068,In_1030);
or U3345 (N_3345,In_1089,N_2901);
xnor U3346 (N_3346,In_546,N_2652);
or U3347 (N_3347,In_3557,N_2365);
nor U3348 (N_3348,In_4489,N_167);
nand U3349 (N_3349,N_2323,N_542);
nand U3350 (N_3350,N_1410,N_1516);
xnor U3351 (N_3351,N_2989,N_1107);
nand U3352 (N_3352,N_1223,N_2395);
nor U3353 (N_3353,N_2125,N_1628);
and U3354 (N_3354,N_1435,N_2501);
xor U3355 (N_3355,N_2771,In_3658);
nor U3356 (N_3356,N_2915,In_4189);
or U3357 (N_3357,N_862,N_806);
and U3358 (N_3358,In_1963,N_878);
nor U3359 (N_3359,N_1547,N_2289);
and U3360 (N_3360,N_2659,N_2621);
and U3361 (N_3361,In_4523,N_2186);
nor U3362 (N_3362,N_1015,In_1680);
or U3363 (N_3363,N_2350,N_2043);
or U3364 (N_3364,N_2213,N_817);
nor U3365 (N_3365,N_2379,In_4680);
or U3366 (N_3366,N_1572,In_3642);
and U3367 (N_3367,N_2538,N_1965);
nand U3368 (N_3368,N_520,N_2122);
nand U3369 (N_3369,N_2602,In_1766);
or U3370 (N_3370,N_2406,In_4493);
nand U3371 (N_3371,N_2973,N_1127);
and U3372 (N_3372,In_1082,In_874);
and U3373 (N_3373,N_549,N_2838);
xor U3374 (N_3374,N_2851,N_1234);
nand U3375 (N_3375,N_134,In_4097);
nand U3376 (N_3376,N_2307,N_2993);
xor U3377 (N_3377,N_1703,In_472);
nand U3378 (N_3378,N_1181,In_2334);
nor U3379 (N_3379,N_986,N_2610);
or U3380 (N_3380,N_2834,In_3789);
nor U3381 (N_3381,In_945,N_2811);
nand U3382 (N_3382,In_4115,N_1633);
or U3383 (N_3383,N_2835,N_752);
and U3384 (N_3384,N_2847,In_3852);
nand U3385 (N_3385,In_153,N_2745);
xor U3386 (N_3386,In_2473,N_2965);
xnor U3387 (N_3387,N_2962,N_2080);
nor U3388 (N_3388,N_186,N_508);
and U3389 (N_3389,N_1759,N_2663);
and U3390 (N_3390,N_2526,N_2760);
nand U3391 (N_3391,In_1987,In_2103);
or U3392 (N_3392,In_3967,In_3899);
xnor U3393 (N_3393,N_38,N_1238);
nor U3394 (N_3394,N_2975,N_2037);
nor U3395 (N_3395,In_2509,In_4834);
nor U3396 (N_3396,N_1983,N_2676);
and U3397 (N_3397,N_2828,In_1437);
xor U3398 (N_3398,N_2733,N_945);
nor U3399 (N_3399,N_2173,N_1357);
and U3400 (N_3400,N_2784,N_2410);
nor U3401 (N_3401,N_2587,N_2103);
and U3402 (N_3402,In_4991,In_2657);
nor U3403 (N_3403,In_4517,N_2263);
xnor U3404 (N_3404,N_2562,In_200);
xor U3405 (N_3405,In_568,N_47);
xnor U3406 (N_3406,In_3641,N_2708);
xor U3407 (N_3407,In_2026,N_208);
or U3408 (N_3408,N_2651,N_1808);
nor U3409 (N_3409,N_1779,N_918);
and U3410 (N_3410,N_2943,N_2577);
xor U3411 (N_3411,In_590,N_2692);
or U3412 (N_3412,N_1861,N_2966);
nand U3413 (N_3413,N_938,In_289);
nor U3414 (N_3414,N_1726,N_2888);
or U3415 (N_3415,N_2643,N_949);
xor U3416 (N_3416,N_2177,N_2604);
xnor U3417 (N_3417,N_1869,In_2645);
or U3418 (N_3418,N_2722,N_2369);
nor U3419 (N_3419,N_2618,In_2151);
nor U3420 (N_3420,N_2773,N_1856);
or U3421 (N_3421,N_2102,N_1101);
nor U3422 (N_3422,N_643,N_502);
xnor U3423 (N_3423,N_2436,N_2997);
or U3424 (N_3424,N_1639,In_720);
or U3425 (N_3425,N_1889,In_391);
and U3426 (N_3426,N_2354,N_2636);
or U3427 (N_3427,In_2761,In_4333);
nor U3428 (N_3428,N_0,N_2714);
nand U3429 (N_3429,N_2762,In_443);
and U3430 (N_3430,N_2407,N_735);
and U3431 (N_3431,N_1709,In_40);
nor U3432 (N_3432,In_4332,In_4085);
xor U3433 (N_3433,N_1773,In_2177);
xnor U3434 (N_3434,N_2574,In_2668);
xnor U3435 (N_3435,N_1515,N_2808);
xnor U3436 (N_3436,N_2741,In_2086);
xnor U3437 (N_3437,N_2738,N_2932);
xnor U3438 (N_3438,N_1239,In_1452);
nor U3439 (N_3439,N_422,N_2560);
nand U3440 (N_3440,N_1916,N_2869);
or U3441 (N_3441,N_560,In_4418);
xnor U3442 (N_3442,In_4282,N_2887);
xnor U3443 (N_3443,N_1857,N_2034);
nand U3444 (N_3444,N_2642,N_2135);
and U3445 (N_3445,N_805,In_1948);
or U3446 (N_3446,N_2362,In_1663);
nor U3447 (N_3447,In_3475,N_2250);
nor U3448 (N_3448,N_2787,N_2471);
or U3449 (N_3449,In_3845,N_2933);
nand U3450 (N_3450,In_1049,N_2450);
and U3451 (N_3451,N_1847,In_2901);
or U3452 (N_3452,N_2781,N_1258);
and U3453 (N_3453,N_2987,N_2535);
nor U3454 (N_3454,In_1149,In_2126);
or U3455 (N_3455,In_3546,N_2074);
xnor U3456 (N_3456,N_1363,N_2420);
or U3457 (N_3457,N_2789,N_2682);
nor U3458 (N_3458,N_2393,N_2656);
nor U3459 (N_3459,N_714,N_2009);
and U3460 (N_3460,N_2731,N_795);
nor U3461 (N_3461,N_2473,In_1892);
and U3462 (N_3462,N_908,N_2696);
xor U3463 (N_3463,In_2665,In_1195);
nand U3464 (N_3464,In_1561,N_2954);
or U3465 (N_3465,N_2824,In_937);
or U3466 (N_3466,N_2045,N_2879);
nor U3467 (N_3467,N_2596,N_1624);
nand U3468 (N_3468,In_1856,In_3333);
and U3469 (N_3469,N_2693,N_1599);
or U3470 (N_3470,In_1458,N_1466);
nand U3471 (N_3471,In_814,N_2927);
and U3472 (N_3472,N_1767,In_1860);
and U3473 (N_3473,N_1830,In_491);
xor U3474 (N_3474,N_1844,In_3160);
xnor U3475 (N_3475,In_1146,N_2517);
or U3476 (N_3476,N_651,N_2518);
and U3477 (N_3477,In_108,N_2423);
nand U3478 (N_3478,N_1173,N_2361);
and U3479 (N_3479,In_237,N_2777);
or U3480 (N_3480,N_597,In_4800);
nor U3481 (N_3481,In_1074,N_1798);
nor U3482 (N_3482,N_151,N_2268);
or U3483 (N_3483,N_2594,N_1563);
nand U3484 (N_3484,N_2882,N_2611);
and U3485 (N_3485,N_1529,In_1017);
or U3486 (N_3486,In_1104,N_1497);
nor U3487 (N_3487,N_2870,In_4952);
and U3488 (N_3488,N_1368,N_2333);
nand U3489 (N_3489,N_2098,N_1984);
nor U3490 (N_3490,N_620,N_1228);
and U3491 (N_3491,In_2861,In_2371);
nand U3492 (N_3492,N_2539,N_2893);
nand U3493 (N_3493,In_4155,In_1923);
xnor U3494 (N_3494,In_1094,N_277);
or U3495 (N_3495,In_2953,In_4151);
and U3496 (N_3496,In_2146,In_2727);
nor U3497 (N_3497,N_2820,N_1714);
xnor U3498 (N_3498,N_2561,N_2505);
nor U3499 (N_3499,N_2195,N_2898);
and U3500 (N_3500,N_2414,N_1263);
and U3501 (N_3501,N_294,N_189);
nand U3502 (N_3502,N_3397,N_3265);
and U3503 (N_3503,In_3500,N_3311);
xor U3504 (N_3504,In_1600,N_2780);
or U3505 (N_3505,N_2367,N_2707);
or U3506 (N_3506,N_3071,N_2585);
or U3507 (N_3507,N_1993,N_3127);
nand U3508 (N_3508,N_3055,N_1919);
xnor U3509 (N_3509,N_3386,N_2940);
and U3510 (N_3510,N_1604,N_1222);
nand U3511 (N_3511,In_186,N_3140);
nand U3512 (N_3512,N_2225,N_1236);
nand U3513 (N_3513,N_3017,N_976);
and U3514 (N_3514,N_3136,N_2028);
and U3515 (N_3515,N_3315,N_3253);
nand U3516 (N_3516,N_97,N_3132);
nor U3517 (N_3517,In_2282,N_3349);
xor U3518 (N_3518,N_3451,N_2119);
nand U3519 (N_3519,N_3326,N_3089);
or U3520 (N_3520,In_1130,N_3441);
nor U3521 (N_3521,N_3008,N_2648);
xor U3522 (N_3522,N_3312,N_2524);
and U3523 (N_3523,In_290,N_3323);
and U3524 (N_3524,In_655,N_1456);
and U3525 (N_3525,N_3275,N_1279);
nand U3526 (N_3526,N_2592,In_3780);
or U3527 (N_3527,N_3348,N_2726);
nor U3528 (N_3528,N_3210,N_2525);
nor U3529 (N_3529,N_2936,N_418);
nand U3530 (N_3530,N_3086,N_2359);
xor U3531 (N_3531,N_3338,N_882);
nand U3532 (N_3532,In_4,In_1540);
and U3533 (N_3533,In_3332,N_2276);
xor U3534 (N_3534,N_3081,N_3028);
nor U3535 (N_3535,In_759,In_3183);
nand U3536 (N_3536,N_3058,N_1863);
nand U3537 (N_3537,N_3262,N_2812);
and U3538 (N_3538,In_1408,N_2922);
nor U3539 (N_3539,N_2166,In_2774);
xor U3540 (N_3540,In_1249,N_3103);
and U3541 (N_3541,N_3455,In_2172);
nand U3542 (N_3542,N_1399,In_2220);
nand U3543 (N_3543,N_3432,N_2197);
or U3544 (N_3544,N_3419,N_1620);
nand U3545 (N_3545,In_2494,N_3139);
nand U3546 (N_3546,In_3179,In_2591);
nand U3547 (N_3547,In_2524,N_1679);
nor U3548 (N_3548,In_207,In_4700);
nor U3549 (N_3549,N_3379,In_4734);
and U3550 (N_3550,In_816,N_2629);
and U3551 (N_3551,N_3043,N_3284);
nand U3552 (N_3552,N_60,In_966);
xor U3553 (N_3553,N_634,N_2256);
nand U3554 (N_3554,N_691,In_2788);
xnor U3555 (N_3555,N_1886,In_794);
or U3556 (N_3556,N_3182,In_1776);
and U3557 (N_3557,In_714,N_3310);
or U3558 (N_3558,N_409,N_516);
or U3559 (N_3559,N_2233,N_3307);
nand U3560 (N_3560,N_2730,N_3087);
nor U3561 (N_3561,N_3346,N_2555);
and U3562 (N_3562,N_3,N_2655);
xnor U3563 (N_3563,N_3472,N_1781);
nand U3564 (N_3564,N_2059,In_3708);
nor U3565 (N_3565,N_2593,N_3375);
and U3566 (N_3566,N_2783,N_3293);
or U3567 (N_3567,N_2684,N_3400);
or U3568 (N_3568,N_2664,N_1716);
and U3569 (N_3569,N_2677,N_2599);
nor U3570 (N_3570,N_2661,In_648);
nand U3571 (N_3571,N_1810,N_1358);
nor U3572 (N_3572,N_3014,In_3571);
nand U3573 (N_3573,N_2299,N_2825);
xnor U3574 (N_3574,N_3120,N_3224);
nor U3575 (N_3575,In_4860,N_881);
nor U3576 (N_3576,N_130,N_2277);
xnor U3577 (N_3577,N_1302,N_2120);
nor U3578 (N_3578,N_2644,In_306);
and U3579 (N_3579,N_3299,N_14);
nand U3580 (N_3580,N_3281,N_3289);
nor U3581 (N_3581,N_3487,N_2371);
nand U3582 (N_3582,In_3763,In_1883);
or U3583 (N_3583,N_2011,N_919);
and U3584 (N_3584,N_2366,N_998);
nor U3585 (N_3585,N_3254,N_2241);
nor U3586 (N_3586,N_2437,N_3080);
nor U3587 (N_3587,N_3363,N_3421);
nand U3588 (N_3588,N_2279,N_507);
nor U3589 (N_3589,In_3618,In_2227);
nand U3590 (N_3590,N_3309,In_4479);
or U3591 (N_3591,N_1683,In_1113);
nor U3592 (N_3592,In_4796,N_3385);
nand U3593 (N_3593,In_4186,N_1129);
nand U3594 (N_3594,N_3077,N_2355);
nor U3595 (N_3595,N_3308,N_1978);
nor U3596 (N_3596,In_506,In_2251);
nand U3597 (N_3597,N_3436,N_3423);
xnor U3598 (N_3598,N_1575,N_2426);
xnor U3599 (N_3599,N_2641,N_3484);
and U3600 (N_3600,N_930,In_3825);
and U3601 (N_3601,N_1768,N_3112);
nand U3602 (N_3602,N_2788,In_3125);
nand U3603 (N_3603,In_1191,N_3344);
nor U3604 (N_3604,N_3334,N_2357);
and U3605 (N_3605,N_1918,N_3056);
or U3606 (N_3606,N_1147,In_1999);
or U3607 (N_3607,N_2549,N_3450);
or U3608 (N_3608,N_3366,N_1831);
and U3609 (N_3609,N_893,N_101);
and U3610 (N_3610,N_1752,N_2349);
nor U3611 (N_3611,N_3306,In_4638);
nor U3612 (N_3612,N_2413,N_3033);
xnor U3613 (N_3613,N_245,N_719);
or U3614 (N_3614,In_4537,N_3006);
nand U3615 (N_3615,N_3092,N_989);
xor U3616 (N_3616,N_3414,N_1069);
nor U3617 (N_3617,N_3351,N_2316);
xnor U3618 (N_3618,N_3357,N_3149);
and U3619 (N_3619,N_1169,N_3482);
and U3620 (N_3620,N_1953,N_2092);
nand U3621 (N_3621,N_2739,N_640);
nor U3622 (N_3622,In_1429,N_2105);
nor U3623 (N_3623,N_3395,N_3250);
nand U3624 (N_3624,N_1345,In_4301);
xor U3625 (N_3625,N_3152,N_3465);
and U3626 (N_3626,In_1529,N_2918);
and U3627 (N_3627,In_3980,In_4685);
and U3628 (N_3628,In_2166,N_2023);
nor U3629 (N_3629,N_2748,N_3173);
or U3630 (N_3630,N_2646,N_2769);
nand U3631 (N_3631,N_3096,N_3431);
nand U3632 (N_3632,N_545,N_3453);
xor U3633 (N_3633,N_2576,N_3147);
and U3634 (N_3634,In_4652,N_3012);
or U3635 (N_3635,In_2059,N_3213);
xor U3636 (N_3636,N_3359,In_2400);
nor U3637 (N_3637,In_28,N_3200);
or U3638 (N_3638,N_3413,N_2906);
nand U3639 (N_3639,In_2351,N_1024);
nand U3640 (N_3640,N_2791,In_99);
nand U3641 (N_3641,N_2862,N_605);
nand U3642 (N_3642,N_1104,N_3271);
and U3643 (N_3643,N_3215,N_3019);
and U3644 (N_3644,In_2899,N_2564);
nor U3645 (N_3645,N_3063,N_2717);
or U3646 (N_3646,N_2716,N_2857);
nor U3647 (N_3647,N_3243,N_3042);
nand U3648 (N_3648,In_2628,N_2712);
xnor U3649 (N_3649,N_3354,N_2778);
and U3650 (N_3650,N_2718,N_3418);
xor U3651 (N_3651,N_1871,In_3330);
or U3652 (N_3652,In_3467,N_2565);
xnor U3653 (N_3653,N_2667,N_2280);
xor U3654 (N_3654,N_3216,N_3068);
xor U3655 (N_3655,N_3294,N_194);
or U3656 (N_3656,In_3497,N_3075);
nor U3657 (N_3657,N_2890,In_3854);
nor U3658 (N_3658,N_2832,N_3057);
nor U3659 (N_3659,N_718,N_2628);
or U3660 (N_3660,N_906,N_2176);
xor U3661 (N_3661,N_3187,N_3191);
xnor U3662 (N_3662,N_3239,N_3399);
or U3663 (N_3663,In_735,In_624);
xor U3664 (N_3664,In_1645,In_4540);
nor U3665 (N_3665,N_3364,In_4478);
xnor U3666 (N_3666,N_2399,N_2235);
xor U3667 (N_3667,N_978,N_3342);
xnor U3668 (N_3668,N_2187,N_3264);
and U3669 (N_3669,N_372,N_614);
nand U3670 (N_3670,N_3041,In_4678);
xnor U3671 (N_3671,N_1751,N_1457);
xor U3672 (N_3672,N_3398,N_2985);
or U3673 (N_3673,N_3367,N_3454);
or U3674 (N_3674,N_2106,N_2101);
nor U3675 (N_3675,N_2657,N_2327);
or U3676 (N_3676,N_2449,N_829);
nor U3677 (N_3677,N_1873,N_2378);
and U3678 (N_3678,N_3268,N_2735);
nor U3679 (N_3679,N_3462,N_3322);
nand U3680 (N_3680,N_3031,In_2317);
xor U3681 (N_3681,N_2152,N_2544);
and U3682 (N_3682,N_3218,N_2691);
or U3683 (N_3683,N_1183,In_4123);
xnor U3684 (N_3684,N_3404,N_2721);
nor U3685 (N_3685,N_3094,N_3282);
xnor U3686 (N_3686,N_2704,N_2947);
and U3687 (N_3687,N_1839,N_3480);
xnor U3688 (N_3688,N_2377,N_2867);
nand U3689 (N_3689,In_3742,N_2996);
and U3690 (N_3690,N_2175,In_4574);
xor U3691 (N_3691,N_1201,N_3073);
xnor U3692 (N_3692,N_3405,N_404);
nor U3693 (N_3693,N_2912,N_3230);
or U3694 (N_3694,N_3280,N_3171);
nand U3695 (N_3695,In_444,N_2607);
nand U3696 (N_3696,N_3238,N_3320);
xor U3697 (N_3697,N_1254,N_2950);
or U3698 (N_3698,N_3227,N_2978);
nand U3699 (N_3699,N_1046,N_1455);
xnor U3700 (N_3700,N_2253,N_1888);
xor U3701 (N_3701,N_3297,In_2316);
and U3702 (N_3702,N_3076,N_1087);
xnor U3703 (N_3703,N_3374,N_2130);
or U3704 (N_3704,N_3066,N_1943);
and U3705 (N_3705,N_3412,N_2804);
and U3706 (N_3706,N_2255,N_278);
and U3707 (N_3707,N_2356,N_2035);
or U3708 (N_3708,N_2036,In_3044);
xor U3709 (N_3709,N_2212,N_2920);
nor U3710 (N_3710,N_2452,N_2839);
xor U3711 (N_3711,N_3093,N_2761);
nand U3712 (N_3712,In_3956,N_2540);
xor U3713 (N_3713,N_2689,N_2339);
or U3714 (N_3714,N_3074,N_2797);
and U3715 (N_3715,N_3206,In_4203);
or U3716 (N_3716,N_2874,N_1758);
nand U3717 (N_3717,In_1314,In_2379);
nor U3718 (N_3718,In_1587,N_3483);
and U3719 (N_3719,N_1979,N_3146);
or U3720 (N_3720,N_3095,N_2408);
nand U3721 (N_3721,N_3361,In_1844);
nor U3722 (N_3722,In_2639,N_2154);
or U3723 (N_3723,N_2507,In_3419);
and U3724 (N_3724,In_4089,N_2662);
and U3725 (N_3725,In_3781,N_2645);
xor U3726 (N_3726,In_4038,N_3091);
xnor U3727 (N_3727,In_1127,N_3353);
or U3728 (N_3728,N_3159,N_853);
and U3729 (N_3729,N_2372,N_1958);
or U3730 (N_3730,N_606,N_3272);
nor U3731 (N_3731,N_3179,N_3174);
xor U3732 (N_3732,N_2923,N_3319);
nor U3733 (N_3733,In_192,N_3183);
xor U3734 (N_3734,N_2983,In_4043);
nand U3735 (N_3735,N_3189,In_4929);
xnor U3736 (N_3736,N_3246,N_3137);
nand U3737 (N_3737,N_2191,N_1621);
nand U3738 (N_3738,N_2917,N_1521);
and U3739 (N_3739,In_4124,In_4161);
xor U3740 (N_3740,In_4451,N_2864);
and U3741 (N_3741,N_3048,N_2872);
xnor U3742 (N_3742,N_3013,N_1974);
or U3743 (N_3743,N_3229,N_3290);
nand U3744 (N_3744,N_3065,N_3036);
and U3745 (N_3745,N_2252,N_3027);
or U3746 (N_3746,In_2624,N_3030);
and U3747 (N_3747,N_2563,N_3205);
or U3748 (N_3748,N_956,N_3203);
nor U3749 (N_3749,N_3430,N_3478);
xnor U3750 (N_3750,N_3195,N_2905);
xnor U3751 (N_3751,N_3212,N_3439);
xor U3752 (N_3752,N_1907,N_3356);
and U3753 (N_3753,N_1772,N_3261);
nor U3754 (N_3754,In_1259,N_2779);
nor U3755 (N_3755,In_1064,N_758);
nand U3756 (N_3756,N_595,N_3135);
and U3757 (N_3757,In_3998,In_4425);
nand U3758 (N_3758,N_1707,In_1212);
nand U3759 (N_3759,N_1964,N_583);
xor U3760 (N_3760,N_3304,N_1765);
or U3761 (N_3761,N_1397,In_3048);
nor U3762 (N_3762,N_2384,N_3427);
nor U3763 (N_3763,N_3220,N_2394);
nand U3764 (N_3764,N_555,N_3128);
nor U3765 (N_3765,In_3051,N_3362);
nor U3766 (N_3766,N_3129,N_3105);
or U3767 (N_3767,N_22,In_3465);
xor U3768 (N_3768,In_3499,N_3002);
xor U3769 (N_3769,N_2494,N_1442);
and U3770 (N_3770,N_1818,N_2486);
and U3771 (N_3771,N_2990,N_3394);
nand U3772 (N_3772,In_1582,N_819);
and U3773 (N_3773,N_3347,N_1014);
and U3774 (N_3774,N_3047,N_3188);
xnor U3775 (N_3775,In_3741,N_3154);
nand U3776 (N_3776,N_2649,N_3085);
and U3777 (N_3777,N_1945,N_2068);
xnor U3778 (N_3778,In_2596,N_2654);
and U3779 (N_3779,N_2317,In_1395);
or U3780 (N_3780,N_3251,N_3099);
nand U3781 (N_3781,N_2440,N_2516);
xnor U3782 (N_3782,N_3318,N_3005);
nand U3783 (N_3783,N_1033,In_1538);
and U3784 (N_3784,N_3360,N_3274);
nor U3785 (N_3785,In_3603,In_4828);
and U3786 (N_3786,N_3343,N_2854);
xor U3787 (N_3787,N_3035,N_2514);
and U3788 (N_3788,N_2949,N_1237);
nand U3789 (N_3789,N_3053,In_847);
and U3790 (N_3790,N_2827,N_3381);
nand U3791 (N_3791,In_118,N_3023);
nand U3792 (N_3792,N_3355,N_756);
and U3793 (N_3793,N_1449,N_3167);
nor U3794 (N_3794,N_3464,N_2830);
xnor U3795 (N_3795,N_1730,In_51);
xnor U3796 (N_3796,N_2865,N_3285);
or U3797 (N_3797,In_2410,N_1587);
and U3798 (N_3798,N_3499,N_3222);
xor U3799 (N_3799,N_538,N_2701);
or U3800 (N_3800,N_3350,N_2833);
or U3801 (N_3801,In_2305,N_2556);
xor U3802 (N_3802,N_2254,N_1089);
nor U3803 (N_3803,N_3336,N_3490);
and U3804 (N_3804,N_1483,N_1175);
and U3805 (N_3805,N_3341,N_2660);
xnor U3806 (N_3806,N_2113,N_2894);
nor U3807 (N_3807,N_2650,In_4727);
and U3808 (N_3808,N_2776,In_2982);
and U3809 (N_3809,N_2727,N_3034);
nand U3810 (N_3810,N_2208,N_3166);
xor U3811 (N_3811,N_1947,N_1708);
nand U3812 (N_3812,N_2822,N_3273);
nand U3813 (N_3813,N_3266,N_357);
or U3814 (N_3814,N_63,In_4881);
and U3815 (N_3815,In_609,N_3106);
nor U3816 (N_3816,N_3377,N_155);
or U3817 (N_3817,N_86,N_429);
xor U3818 (N_3818,N_3237,N_124);
and U3819 (N_3819,N_1045,N_2385);
xor U3820 (N_3820,N_2680,In_2606);
nor U3821 (N_3821,In_576,N_3257);
or U3822 (N_3822,N_1678,N_826);
nor U3823 (N_3823,In_2295,N_2775);
and U3824 (N_3824,N_2798,N_3121);
xnor U3825 (N_3825,N_2860,In_3440);
and U3826 (N_3826,N_1687,N_3260);
nand U3827 (N_3827,In_915,N_3471);
and U3828 (N_3828,N_1240,N_3245);
or U3829 (N_3829,N_762,In_1447);
and U3830 (N_3830,N_3169,In_295);
or U3831 (N_3831,N_2257,N_3131);
xor U3832 (N_3832,N_16,N_3233);
nand U3833 (N_3833,N_3329,N_3078);
xor U3834 (N_3834,N_2744,N_1039);
or U3835 (N_3835,N_3124,N_1658);
xor U3836 (N_3836,In_4696,N_3302);
xor U3837 (N_3837,In_165,N_2537);
xor U3838 (N_3838,N_3088,N_3003);
nand U3839 (N_3839,In_3184,N_2999);
nand U3840 (N_3840,N_476,In_2355);
xnor U3841 (N_3841,N_2523,N_2751);
or U3842 (N_3842,N_2935,In_4643);
or U3843 (N_3843,In_1532,In_2061);
xor U3844 (N_3844,In_4710,N_2638);
nor U3845 (N_3845,N_2809,N_2740);
and U3846 (N_3846,N_3082,N_2031);
nor U3847 (N_3847,N_784,N_2091);
nor U3848 (N_3848,N_2971,N_2980);
nand U3849 (N_3849,N_2686,In_276);
or U3850 (N_3850,N_3228,N_3435);
and U3851 (N_3851,In_4244,N_1642);
and U3852 (N_3852,In_1647,N_2653);
and U3853 (N_3853,N_2608,N_2550);
and U3854 (N_3854,In_37,N_2807);
nand U3855 (N_3855,N_3000,N_3138);
nand U3856 (N_3856,N_2055,N_2249);
nor U3857 (N_3857,N_959,In_1100);
or U3858 (N_3858,N_2942,N_2060);
xor U3859 (N_3859,In_721,N_3110);
or U3860 (N_3860,N_3252,N_1635);
or U3861 (N_3861,N_3491,N_2612);
or U3862 (N_3862,N_3434,N_2666);
and U3863 (N_3863,N_2142,In_534);
and U3864 (N_3864,N_3101,In_3055);
nor U3865 (N_3865,N_3051,In_4369);
or U3866 (N_3866,N_3425,N_423);
or U3867 (N_3867,N_2948,N_1386);
or U3868 (N_3868,N_3111,N_3317);
nand U3869 (N_3869,N_2926,In_2794);
nand U3870 (N_3870,In_2555,N_3181);
xor U3871 (N_3871,N_3186,N_2878);
xor U3872 (N_3872,N_665,N_3337);
or U3873 (N_3873,N_1366,N_2746);
xor U3874 (N_3874,N_2755,N_2913);
xor U3875 (N_3875,N_3365,N_3160);
or U3876 (N_3876,N_3217,In_3890);
nand U3877 (N_3877,N_2107,N_2572);
and U3878 (N_3878,N_2928,N_1152);
nand U3879 (N_3879,In_1949,In_3004);
or U3880 (N_3880,N_3161,N_266);
nor U3881 (N_3881,N_1262,N_1690);
and U3882 (N_3882,In_1296,N_2338);
and U3883 (N_3883,In_2694,N_2772);
nor U3884 (N_3884,N_3387,N_3062);
nor U3885 (N_3885,N_3242,N_2930);
xnor U3886 (N_3886,N_2291,N_970);
xor U3887 (N_3887,N_2709,N_1860);
xnor U3888 (N_3888,N_2624,N_693);
nor U3889 (N_3889,In_973,N_2161);
xor U3890 (N_3890,N_3198,N_2859);
xor U3891 (N_3891,N_3175,N_3142);
or U3892 (N_3892,N_171,N_49);
nor U3893 (N_3893,N_3204,N_2795);
nor U3894 (N_3894,In_2588,In_1885);
xor U3895 (N_3895,In_86,In_341);
nand U3896 (N_3896,N_2095,N_2261);
nand U3897 (N_3897,N_3443,N_3372);
and U3898 (N_3898,N_3037,N_3177);
or U3899 (N_3899,N_3018,In_4767);
and U3900 (N_3900,N_2287,N_2169);
xor U3901 (N_3901,N_3100,N_2422);
or U3902 (N_3902,N_2167,N_2785);
and U3903 (N_3903,N_1459,N_2632);
or U3904 (N_3904,N_2015,N_3134);
nand U3905 (N_3905,N_1601,N_3328);
xor U3906 (N_3906,N_2084,N_3192);
nand U3907 (N_3907,N_568,N_2907);
xor U3908 (N_3908,In_3222,N_173);
nor U3909 (N_3909,N_3277,N_1881);
nand U3910 (N_3910,N_2077,In_1365);
and U3911 (N_3911,N_501,N_3352);
nand U3912 (N_3912,N_2162,N_3115);
or U3913 (N_3913,N_604,N_65);
or U3914 (N_3914,N_1880,N_1245);
and U3915 (N_3915,N_3486,N_2530);
nand U3916 (N_3916,N_1078,N_2434);
and U3917 (N_3917,N_3130,N_1960);
and U3918 (N_3918,In_3140,N_1626);
nand U3919 (N_3919,In_4667,In_3910);
nand U3920 (N_3920,N_3049,N_2221);
xor U3921 (N_3921,N_2557,N_3463);
nor U3922 (N_3922,In_920,N_3240);
or U3923 (N_3923,N_3489,In_407);
or U3924 (N_3924,N_3340,N_3158);
nand U3925 (N_3925,In_1717,N_3378);
nor U3926 (N_3926,N_571,N_3321);
nor U3927 (N_3927,N_2889,N_3316);
nor U3928 (N_3928,N_3133,N_3314);
or U3929 (N_3929,N_615,N_3122);
or U3930 (N_3930,In_4070,N_3461);
and U3931 (N_3931,In_4148,N_1704);
and U3932 (N_3932,N_513,In_1756);
and U3933 (N_3933,N_3392,In_3290);
nand U3934 (N_3934,N_3460,N_2765);
and U3935 (N_3935,In_2777,N_2226);
xor U3936 (N_3936,N_802,N_1338);
or U3937 (N_3937,N_2814,N_3108);
or U3938 (N_3938,N_2897,N_1713);
nand U3939 (N_3939,In_4033,N_3278);
nor U3940 (N_3940,N_792,N_2488);
and U3941 (N_3941,N_879,N_3358);
xor U3942 (N_3942,N_3117,N_113);
nand U3943 (N_3943,N_2294,In_2015);
nor U3944 (N_3944,N_2597,N_1131);
nand U3945 (N_3945,N_2938,N_2970);
nor U3946 (N_3946,N_1574,N_3059);
and U3947 (N_3947,In_2523,N_1755);
xnor U3948 (N_3948,N_3157,N_3376);
nor U3949 (N_3949,N_2551,In_2393);
or U3950 (N_3950,In_4336,N_3151);
xor U3951 (N_3951,In_113,N_1329);
and U3952 (N_3952,N_17,N_1661);
xor U3953 (N_3953,N_3444,In_3947);
or U3954 (N_3954,N_1292,N_3313);
nand U3955 (N_3955,N_2030,N_3433);
nand U3956 (N_3956,N_2462,N_2506);
nor U3957 (N_3957,N_1806,N_2992);
or U3958 (N_3958,N_1335,N_2124);
nor U3959 (N_3959,N_3201,In_1837);
or U3960 (N_3960,In_2875,N_2903);
or U3961 (N_3961,N_2389,N_2508);
and U3962 (N_3962,N_3020,N_2715);
nor U3963 (N_3963,N_2183,N_2614);
xnor U3964 (N_3964,In_4475,In_4322);
or U3965 (N_3965,In_776,N_3125);
and U3966 (N_3966,In_1302,N_2732);
and U3967 (N_3967,In_2878,In_2506);
or U3968 (N_3968,N_3396,N_1198);
nand U3969 (N_3969,In_3621,N_1077);
or U3970 (N_3970,N_3370,In_3870);
or U3971 (N_3971,N_3452,In_47);
and U3972 (N_3972,In_4825,N_3473);
and U3973 (N_3973,In_3388,N_3368);
xnor U3974 (N_3974,N_2871,In_1580);
or U3975 (N_3975,N_3114,In_4905);
and U3976 (N_3976,N_2499,N_3170);
or U3977 (N_3977,N_3279,N_3208);
or U3978 (N_3978,N_2376,N_2626);
and U3979 (N_3979,In_2552,N_1763);
or U3980 (N_3980,N_3449,N_1782);
xnor U3981 (N_3981,N_3258,In_3377);
nor U3982 (N_3982,N_3016,N_3305);
xor U3983 (N_3983,N_1807,In_1606);
xor U3984 (N_3984,N_3235,N_3296);
nand U3985 (N_3985,N_3327,In_3206);
nand U3986 (N_3986,N_2956,N_3236);
nand U3987 (N_3987,N_2710,N_3339);
and U3988 (N_3988,N_3098,N_3467);
nand U3989 (N_3989,N_3468,N_3150);
nor U3990 (N_3990,N_2909,N_1941);
nor U3991 (N_3991,In_3853,N_3345);
or U3992 (N_3992,In_3631,N_3331);
xor U3993 (N_3993,N_203,N_3060);
nand U3994 (N_3994,In_3424,N_3244);
nand U3995 (N_3995,N_1893,N_578);
xnor U3996 (N_3996,N_3107,N_2445);
and U3997 (N_3997,N_1615,N_2067);
nand U3998 (N_3998,N_3113,N_2237);
and U3999 (N_3999,N_3070,N_3032);
nand U4000 (N_4000,N_3627,N_3761);
nand U4001 (N_4001,N_305,N_866);
nand U4002 (N_4002,N_3564,N_3919);
nand U4003 (N_4003,In_526,N_3263);
nand U4004 (N_4004,N_2911,N_3283);
or U4005 (N_4005,N_3989,N_3947);
nand U4006 (N_4006,N_3717,N_2831);
nand U4007 (N_4007,N_1333,In_524);
xor U4008 (N_4008,N_2150,N_3816);
or U4009 (N_4009,N_3908,N_3798);
xnor U4010 (N_4010,N_3530,N_3420);
and U4011 (N_4011,In_4530,N_3709);
and U4012 (N_4012,N_3259,In_2680);
or U4013 (N_4013,N_1729,N_3209);
and U4014 (N_4014,N_3555,In_1552);
nor U4015 (N_4015,N_3730,N_3758);
nor U4016 (N_4016,N_3196,N_3595);
nand U4017 (N_4017,N_3779,N_3860);
and U4018 (N_4018,N_3724,N_2039);
nand U4019 (N_4019,N_3689,N_3909);
nand U4020 (N_4020,N_2344,N_1802);
xnor U4021 (N_4021,N_3985,N_3926);
and U4022 (N_4022,N_3211,N_3818);
nor U4023 (N_4023,N_590,N_3675);
or U4024 (N_4024,N_3384,N_933);
or U4025 (N_4025,N_3762,N_3962);
nand U4026 (N_4026,N_855,N_3653);
nor U4027 (N_4027,N_3590,In_4289);
or U4028 (N_4028,N_3097,N_3941);
xor U4029 (N_4029,N_3973,N_2631);
and U4030 (N_4030,N_3025,N_3429);
nand U4031 (N_4031,N_3194,In_1026);
and U4032 (N_4032,N_3990,N_2603);
xnor U4033 (N_4033,N_3069,N_3044);
nor U4034 (N_4034,N_3324,N_3102);
nand U4035 (N_4035,N_3814,N_3647);
xnor U4036 (N_4036,N_3672,N_2081);
xnor U4037 (N_4037,N_3532,N_3734);
nor U4038 (N_4038,N_3807,N_3844);
and U4039 (N_4039,N_2615,N_3738);
and U4040 (N_4040,N_2586,N_3736);
or U4041 (N_4041,N_3492,N_3269);
nor U4042 (N_4042,In_214,N_1308);
nor U4043 (N_4043,N_3702,N_3837);
nor U4044 (N_4044,N_3917,N_3437);
or U4045 (N_4045,N_3967,N_3901);
nand U4046 (N_4046,N_3711,In_4143);
xor U4047 (N_4047,N_3793,N_1027);
or U4048 (N_4048,N_3804,N_3155);
xor U4049 (N_4049,N_3925,N_3872);
nand U4050 (N_4050,In_992,N_3680);
nand U4051 (N_4051,N_3988,N_3972);
or U4052 (N_4052,N_3890,N_3610);
or U4053 (N_4053,N_3603,N_1854);
nor U4054 (N_4054,N_3774,In_1573);
xor U4055 (N_4055,N_2332,N_2304);
xnor U4056 (N_4056,N_3918,In_4071);
nand U4057 (N_4057,N_3813,N_3500);
nor U4058 (N_4058,N_2014,In_3575);
nand U4059 (N_4059,N_699,N_3792);
and U4060 (N_4060,N_2899,N_3679);
nor U4061 (N_4061,N_2570,N_3933);
or U4062 (N_4062,N_3945,N_3475);
nor U4063 (N_4063,N_3232,N_3731);
nor U4064 (N_4064,In_2319,N_3556);
xnor U4065 (N_4065,N_1732,N_3891);
nor U4066 (N_4066,N_3516,In_3946);
or U4067 (N_4067,In_4575,N_3537);
xor U4068 (N_4068,N_3853,N_3791);
nand U4069 (N_4069,N_3518,N_3657);
nand U4070 (N_4070,N_517,N_3409);
or U4071 (N_4071,N_3979,N_3710);
or U4072 (N_4072,N_3604,N_3976);
nand U4073 (N_4073,N_3695,In_2459);
xnor U4074 (N_4074,N_1805,N_3776);
nor U4075 (N_4075,N_2841,N_2994);
nand U4076 (N_4076,N_3373,N_2010);
xnor U4077 (N_4077,N_3930,N_3971);
or U4078 (N_4078,N_3292,In_4152);
nor U4079 (N_4079,N_1867,N_3021);
nor U4080 (N_4080,N_3878,N_3739);
xnor U4081 (N_4081,N_3737,N_3581);
or U4082 (N_4082,N_3503,N_3549);
and U4083 (N_4083,N_565,N_3871);
nand U4084 (N_4084,N_3509,N_3287);
or U4085 (N_4085,N_3223,N_2016);
or U4086 (N_4086,N_3587,N_3846);
nor U4087 (N_4087,N_3732,N_3752);
nand U4088 (N_4088,N_3520,N_3754);
or U4089 (N_4089,N_2706,N_2910);
xnor U4090 (N_4090,N_3303,N_1914);
nor U4091 (N_4091,In_3977,N_3511);
xor U4092 (N_4092,N_3887,N_3893);
and U4093 (N_4093,N_1706,In_1080);
or U4094 (N_4094,N_3219,N_1938);
xnor U4095 (N_4095,N_3716,N_2342);
nor U4096 (N_4096,N_3899,N_1935);
xor U4097 (N_4097,In_810,N_3692);
and U4098 (N_4098,N_3410,N_3607);
nand U4099 (N_4099,N_3045,N_3974);
and U4100 (N_4100,N_3572,N_3867);
nand U4101 (N_4101,N_2858,In_173);
or U4102 (N_4102,N_3984,N_3024);
nand U4103 (N_4103,N_3809,N_3719);
or U4104 (N_4104,N_3857,N_2273);
nor U4105 (N_4105,N_2078,N_3855);
nand U4106 (N_4106,N_3902,N_3596);
nor U4107 (N_4107,In_4879,N_3248);
xnor U4108 (N_4108,N_3965,N_3766);
nand U4109 (N_4109,N_3922,In_2659);
xor U4110 (N_4110,N_1094,N_2658);
xnor U4111 (N_4111,N_3773,N_3288);
xnor U4112 (N_4112,N_1885,N_255);
and U4113 (N_4113,N_3407,N_2568);
and U4114 (N_4114,N_3812,N_3180);
xor U4115 (N_4115,N_3574,In_1927);
nand U4116 (N_4116,N_3640,N_3856);
or U4117 (N_4117,N_3504,N_2673);
xnor U4118 (N_4118,N_3755,In_4884);
nand U4119 (N_4119,N_3440,N_3852);
and U4120 (N_4120,N_3958,N_3832);
xor U4121 (N_4121,N_3767,N_2264);
nand U4122 (N_4122,N_3714,N_602);
or U4123 (N_4123,N_3745,N_3599);
or U4124 (N_4124,In_4805,N_3785);
and U4125 (N_4125,N_3850,N_3998);
and U4126 (N_4126,N_3876,N_3648);
nor U4127 (N_4127,N_1244,N_2260);
nand U4128 (N_4128,N_3369,N_3950);
nand U4129 (N_4129,N_3613,N_3456);
and U4130 (N_4130,N_3506,N_3907);
or U4131 (N_4131,N_3664,In_3468);
nand U4132 (N_4132,N_909,N_3729);
and U4133 (N_4133,N_883,N_3589);
or U4134 (N_4134,N_3858,N_3428);
nor U4135 (N_4135,N_3393,N_646);
nor U4136 (N_4136,N_3527,N_3039);
or U4137 (N_4137,N_3298,In_3479);
nand U4138 (N_4138,N_1388,In_4832);
nor U4139 (N_4139,N_3658,N_3545);
or U4140 (N_4140,N_3141,N_3631);
nand U4141 (N_4141,N_3956,N_645);
nand U4142 (N_4142,N_3911,N_3910);
xor U4143 (N_4143,N_3249,N_3865);
nand U4144 (N_4144,In_3745,N_3707);
nor U4145 (N_4145,N_2647,N_3295);
nor U4146 (N_4146,N_3651,In_805);
or U4147 (N_4147,N_3700,N_3847);
or U4148 (N_4148,N_3474,N_3799);
nor U4149 (N_4149,N_3609,In_3976);
nor U4150 (N_4150,N_3704,N_3932);
or U4151 (N_4151,N_3903,N_2269);
nor U4152 (N_4152,N_3038,N_3827);
nand U4153 (N_4153,N_3863,N_3782);
xor U4154 (N_4154,N_1172,N_2815);
xnor U4155 (N_4155,N_2977,In_2269);
nor U4156 (N_4156,N_3894,N_3952);
nand U4157 (N_4157,N_3753,N_3817);
nand U4158 (N_4158,N_3888,N_3795);
xor U4159 (N_4159,N_3565,N_3948);
nand U4160 (N_4160,N_3960,N_3459);
nand U4161 (N_4161,N_3953,In_4775);
and U4162 (N_4162,N_2466,N_3788);
xor U4163 (N_4163,N_3602,N_3416);
and U4164 (N_4164,N_3961,N_3481);
nand U4165 (N_4165,N_2941,N_3514);
and U4166 (N_4166,N_3643,N_3004);
xnor U4167 (N_4167,N_3403,N_2683);
and U4168 (N_4168,N_3567,N_3551);
nand U4169 (N_4169,In_2871,N_1548);
and U4170 (N_4170,N_3507,N_2128);
xor U4171 (N_4171,N_1748,N_2115);
nand U4172 (N_4172,N_3389,N_3221);
nand U4173 (N_4173,N_3954,N_3601);
nor U4174 (N_4174,In_1231,N_1801);
xnor U4175 (N_4175,N_3015,N_3477);
xnor U4176 (N_4176,In_729,N_2955);
and U4177 (N_4177,N_3199,N_3838);
nor U4178 (N_4178,N_1864,N_3148);
nand U4179 (N_4179,N_3501,N_3805);
and U4180 (N_4180,N_1640,In_1419);
nor U4181 (N_4181,N_3997,N_3978);
or U4182 (N_4182,N_3638,N_1987);
nor U4183 (N_4183,N_3825,N_3022);
nor U4184 (N_4184,N_314,N_3943);
xnor U4185 (N_4185,N_3694,N_3231);
nand U4186 (N_4186,N_3929,N_3566);
nor U4187 (N_4187,N_3733,N_3458);
xor U4188 (N_4188,N_3811,N_2163);
nand U4189 (N_4189,N_3447,N_794);
and U4190 (N_4190,N_3618,N_3781);
xnor U4191 (N_4191,N_3839,N_3176);
or U4192 (N_4192,N_3184,N_3688);
and U4193 (N_4193,N_2637,N_3531);
xnor U4194 (N_4194,N_3701,N_3214);
nor U4195 (N_4195,N_3585,N_1991);
xnor U4196 (N_4196,N_3635,N_2136);
and U4197 (N_4197,In_2897,N_3841);
and U4198 (N_4198,N_2147,N_3915);
or U4199 (N_4199,N_3156,N_3513);
or U4200 (N_4200,N_2020,N_3720);
nand U4201 (N_4201,N_3502,N_2919);
or U4202 (N_4202,N_3936,N_3789);
and U4203 (N_4203,N_3875,N_1826);
xor U4204 (N_4204,N_2097,N_3575);
and U4205 (N_4205,N_3644,N_3756);
nor U4206 (N_4206,N_3959,N_3594);
xnor U4207 (N_4207,N_3234,N_3539);
and U4208 (N_4208,N_3722,N_3084);
xnor U4209 (N_4209,N_270,N_3845);
nand U4210 (N_4210,N_3163,In_850);
xnor U4211 (N_4211,N_3605,In_1169);
nand U4212 (N_4212,N_1756,N_3165);
nor U4213 (N_4213,N_3496,In_4374);
and U4214 (N_4214,N_3806,N_3723);
xor U4215 (N_4215,N_2635,N_3834);
nand U4216 (N_4216,N_3826,N_3744);
nand U4217 (N_4217,N_749,In_4995);
and U4218 (N_4218,N_3286,N_3656);
and U4219 (N_4219,N_3898,N_1491);
and U4220 (N_4220,N_2358,N_1481);
xnor U4221 (N_4221,N_570,N_3333);
xor U4222 (N_4222,N_2566,N_2914);
xor U4223 (N_4223,N_3332,N_1155);
nor U4224 (N_4224,N_3764,N_3446);
nor U4225 (N_4225,N_2670,N_2849);
nand U4226 (N_4226,N_2547,In_3892);
xor U4227 (N_4227,In_4356,N_2527);
nor U4228 (N_4228,N_3645,N_3934);
nand U4229 (N_4229,N_3674,N_3485);
and U4230 (N_4230,N_3064,N_2842);
and U4231 (N_4231,N_193,N_3466);
nand U4232 (N_4232,N_3886,N_3061);
nand U4233 (N_4233,N_3569,N_3712);
and U4234 (N_4234,N_3524,N_3547);
nor U4235 (N_4235,N_3620,N_3445);
xor U4236 (N_4236,In_2620,N_1025);
nor U4237 (N_4237,N_2348,In_4594);
or U4238 (N_4238,N_3083,N_110);
and U4239 (N_4239,N_3276,N_3676);
and U4240 (N_4240,N_3247,N_2768);
nor U4241 (N_4241,N_3900,N_743);
nor U4242 (N_4242,N_3854,N_3560);
nand U4243 (N_4243,N_3523,N_3822);
and U4244 (N_4244,N_3267,N_3476);
or U4245 (N_4245,N_3835,N_3931);
or U4246 (N_4246,In_4130,In_4463);
nor U4247 (N_4247,N_3168,N_3949);
and U4248 (N_4248,N_3868,N_3771);
nor U4249 (N_4249,N_2448,N_3699);
nand U4250 (N_4250,N_3126,N_3185);
nand U4251 (N_4251,N_3760,In_4494);
nor U4252 (N_4252,N_2062,N_3540);
xor U4253 (N_4253,N_3579,N_3696);
nor U4254 (N_4254,N_534,N_3291);
and U4255 (N_4255,N_2725,N_2679);
nand U4256 (N_4256,N_3580,N_3011);
nor U4257 (N_4257,N_3873,N_3649);
xnor U4258 (N_4258,N_3226,N_3914);
xnor U4259 (N_4259,N_1746,N_3780);
or U4260 (N_4260,N_3815,N_3986);
xor U4261 (N_4261,N_3479,In_1347);
and U4262 (N_4262,N_3542,N_3639);
or U4263 (N_4263,N_3144,N_3665);
and U4264 (N_4264,N_3646,In_3249);
nand U4265 (N_4265,N_25,N_3786);
or U4266 (N_4266,N_3667,N_3608);
nand U4267 (N_4267,N_2687,N_828);
xnor U4268 (N_4268,N_3823,N_3964);
nor U4269 (N_4269,N_3488,In_451);
and U4270 (N_4270,N_3515,In_4154);
nor U4271 (N_4271,N_3330,N_3951);
or U4272 (N_4272,N_813,N_3708);
nand U4273 (N_4273,N_3380,N_3874);
xor U4274 (N_4274,N_3654,N_2590);
nand U4275 (N_4275,N_3162,N_3207);
xor U4276 (N_4276,N_3256,N_3685);
nor U4277 (N_4277,In_4325,N_2245);
or U4278 (N_4278,N_3072,N_2404);
and U4279 (N_4279,N_3747,N_3877);
or U4280 (N_4280,N_957,N_3568);
or U4281 (N_4281,N_3632,N_3624);
and U4282 (N_4282,N_2286,N_67);
or U4283 (N_4283,In_2521,N_3442);
nor U4284 (N_4284,N_3391,N_185);
or U4285 (N_4285,In_3261,N_2774);
nand U4286 (N_4286,N_3751,N_3546);
or U4287 (N_4287,N_1162,N_3622);
or U4288 (N_4288,N_3007,N_3705);
and U4289 (N_4289,N_1977,N_3810);
and U4290 (N_4290,N_2447,N_3552);
and U4291 (N_4291,N_3862,N_3510);
xor U4292 (N_4292,N_995,N_3270);
or U4293 (N_4293,N_3659,N_3426);
or U4294 (N_4294,N_2782,N_3906);
and U4295 (N_4295,N_3677,N_2724);
or U4296 (N_4296,In_3267,N_2895);
or U4297 (N_4297,N_3939,N_3937);
nand U4298 (N_4298,N_3470,N_3851);
nand U4299 (N_4299,In_1417,N_3923);
or U4300 (N_4300,N_3079,N_3713);
xnor U4301 (N_4301,N_3662,N_3383);
and U4302 (N_4302,N_3884,N_3678);
or U4303 (N_4303,N_2211,In_547);
xnor U4304 (N_4304,N_3054,In_3084);
and U4305 (N_4305,N_2836,N_3050);
and U4306 (N_4306,N_3775,N_2688);
or U4307 (N_4307,N_2391,N_3684);
or U4308 (N_4308,N_2902,In_3659);
or U4309 (N_4309,In_1313,N_3642);
xnor U4310 (N_4310,N_3497,N_1441);
nor U4311 (N_4311,N_1365,In_3284);
or U4312 (N_4312,N_3831,N_3626);
or U4313 (N_4313,N_2069,N_3869);
or U4314 (N_4314,N_3987,In_1066);
and U4315 (N_4315,N_3424,N_3612);
nand U4316 (N_4316,N_3614,N_3553);
or U4317 (N_4317,N_1997,N_3759);
or U4318 (N_4318,In_3797,N_3994);
and U4319 (N_4319,N_3690,In_1102);
xnor U4320 (N_4320,N_3946,N_3582);
xor U4321 (N_4321,N_3882,N_3550);
and U4322 (N_4322,N_3623,N_3650);
and U4323 (N_4323,N_420,N_2767);
nor U4324 (N_4324,N_3686,N_983);
and U4325 (N_4325,N_3652,N_3969);
nor U4326 (N_4326,N_3944,In_1036);
nand U4327 (N_4327,N_3534,N_3495);
nand U4328 (N_4328,N_3718,N_3996);
nor U4329 (N_4329,N_2511,N_3505);
xnor U4330 (N_4330,N_3406,N_3617);
nor U4331 (N_4331,N_3942,N_3543);
and U4332 (N_4332,N_730,N_3895);
or U4333 (N_4333,In_1415,N_3957);
nor U4334 (N_4334,In_486,N_3864);
nand U4335 (N_4335,N_3691,In_4899);
or U4336 (N_4336,N_2964,N_3803);
xor U4337 (N_4337,In_1430,N_3927);
xor U4338 (N_4338,N_1344,N_3611);
nor U4339 (N_4339,N_3576,N_3797);
nor U4340 (N_4340,N_3508,N_3629);
or U4341 (N_4341,N_3457,N_3558);
xor U4342 (N_4342,N_3577,N_3670);
nor U4343 (N_4343,N_3770,N_3584);
nor U4344 (N_4344,In_2499,N_1401);
or U4345 (N_4345,N_3301,N_2300);
xor U4346 (N_4346,N_2217,N_3571);
nor U4347 (N_4347,N_1477,In_2104);
or U4348 (N_4348,N_2140,N_3778);
and U4349 (N_4349,In_4760,N_3849);
nor U4350 (N_4350,N_3661,N_3469);
nand U4351 (N_4351,N_3666,N_2381);
nor U4352 (N_4352,N_3541,In_1694);
nand U4353 (N_4353,N_3561,N_2319);
nand U4354 (N_4354,N_2946,In_4606);
or U4355 (N_4355,In_1360,N_3993);
and U4356 (N_4356,N_3992,N_3721);
xor U4357 (N_4357,N_3892,N_3557);
or U4358 (N_4358,N_3963,N_2672);
or U4359 (N_4359,N_3559,N_3796);
or U4360 (N_4360,N_3883,N_3742);
nor U4361 (N_4361,In_3152,N_2891);
and U4362 (N_4362,N_3821,N_3920);
nor U4363 (N_4363,N_3802,N_3660);
and U4364 (N_4364,N_3544,N_3833);
nor U4365 (N_4365,N_3225,N_3703);
xor U4366 (N_4366,In_1045,N_3001);
and U4367 (N_4367,N_3525,In_3276);
or U4368 (N_4368,N_3123,N_3528);
nor U4369 (N_4369,N_3619,In_2849);
or U4370 (N_4370,N_2737,N_3202);
xnor U4371 (N_4371,N_2041,N_3683);
or U4372 (N_4372,N_3842,N_3727);
and U4373 (N_4373,N_2542,N_3593);
nor U4374 (N_4374,N_3153,N_3824);
nor U4375 (N_4375,N_2553,N_2303);
xor U4376 (N_4376,N_1133,N_1971);
or U4377 (N_4377,N_3512,N_3570);
or U4378 (N_4378,N_3029,N_3889);
or U4379 (N_4379,N_1499,N_3422);
nor U4380 (N_4380,N_3010,N_3197);
or U4381 (N_4381,N_3750,N_1845);
xnor U4382 (N_4382,N_3840,N_2558);
nand U4383 (N_4383,N_3538,N_3870);
or U4384 (N_4384,N_3765,N_3615);
nor U4385 (N_4385,N_3768,N_3859);
nand U4386 (N_4386,N_1405,N_3980);
and U4387 (N_4387,N_3521,N_566);
or U4388 (N_4388,N_2958,N_3583);
and U4389 (N_4389,N_2806,N_3591);
xor U4390 (N_4390,N_3983,In_751);
and U4391 (N_4391,N_2022,In_512);
xnor U4392 (N_4392,N_3438,N_3630);
or U4393 (N_4393,N_3801,N_3735);
and U4394 (N_4394,N_3009,N_2048);
nor U4395 (N_4395,N_3628,N_3794);
nand U4396 (N_4396,N_3382,N_367);
and U4397 (N_4397,N_3746,N_3255);
xnor U4398 (N_4398,In_4176,N_3586);
nand U4399 (N_4399,N_3693,N_3116);
nor U4400 (N_4400,N_1526,N_3673);
xor U4401 (N_4401,N_2613,N_3119);
nand U4402 (N_4402,N_990,N_2588);
and U4403 (N_4403,N_3143,N_2952);
xnor U4404 (N_4404,N_3067,N_3493);
or U4405 (N_4405,N_3109,N_575);
nor U4406 (N_4406,N_3715,N_3592);
and U4407 (N_4407,N_3916,In_2734);
or U4408 (N_4408,In_1086,In_3286);
nand U4409 (N_4409,N_3668,N_3896);
nand U4410 (N_4410,N_929,N_3190);
nand U4411 (N_4411,N_3681,N_3634);
nor U4412 (N_4412,N_3682,In_1637);
nor U4413 (N_4413,N_3529,N_3828);
nor U4414 (N_4414,N_3178,N_1897);
xor U4415 (N_4415,N_2512,N_2088);
or U4416 (N_4416,N_1794,In_863);
xor U4417 (N_4417,N_3772,In_4027);
nand U4418 (N_4418,N_2963,N_3526);
nand U4419 (N_4419,N_3955,N_3970);
and U4420 (N_4420,N_3697,N_3885);
and U4421 (N_4421,N_3026,N_3905);
xor U4422 (N_4422,N_3928,N_3999);
and U4423 (N_4423,N_3769,N_3118);
and U4424 (N_4424,N_3164,N_3600);
nor U4425 (N_4425,N_3982,N_3390);
nor U4426 (N_4426,N_2756,N_3880);
and U4427 (N_4427,N_3052,N_3881);
or U4428 (N_4428,N_3562,N_3897);
nand U4429 (N_4429,N_1912,N_3663);
xor U4430 (N_4430,N_3641,N_3625);
nor U4431 (N_4431,N_3402,N_3743);
or U4432 (N_4432,N_3921,N_3763);
nand U4433 (N_4433,N_2583,In_3392);
nor U4434 (N_4434,N_3968,In_1790);
nor U4435 (N_4435,N_3517,N_3535);
and U4436 (N_4436,N_2293,N_1573);
or U4437 (N_4437,N_2301,N_2883);
nor U4438 (N_4438,N_3388,N_3783);
and U4439 (N_4439,N_2108,N_3040);
or U4440 (N_4440,N_1790,N_3533);
nor U4441 (N_4441,N_3866,N_3836);
and U4442 (N_4442,N_3335,N_3408);
nand U4443 (N_4443,N_2504,N_3616);
or U4444 (N_4444,In_2375,N_3757);
xor U4445 (N_4445,N_2519,N_3981);
or U4446 (N_4446,In_71,N_3687);
and U4447 (N_4447,N_3966,N_3411);
nor U4448 (N_4448,N_3726,N_3655);
nor U4449 (N_4449,N_3241,In_4259);
nor U4450 (N_4450,N_3401,N_1200);
xor U4451 (N_4451,N_3498,N_3749);
nor U4452 (N_4452,N_3621,N_2736);
and U4453 (N_4453,N_592,N_3935);
nor U4454 (N_4454,N_3588,N_3415);
and U4455 (N_4455,N_3090,N_3819);
xor U4456 (N_4456,N_3904,N_3741);
or U4457 (N_4457,N_3777,In_3045);
and U4458 (N_4458,N_3172,N_2625);
and U4459 (N_4459,N_2829,N_3536);
or U4460 (N_4460,N_1930,In_1155);
or U4461 (N_4461,N_2669,N_3787);
and U4462 (N_4462,In_565,N_2472);
nor U4463 (N_4463,N_3879,N_2749);
nor U4464 (N_4464,In_1391,N_3636);
or U4465 (N_4465,N_3606,In_4856);
nand U4466 (N_4466,N_3548,N_3193);
xnor U4467 (N_4467,N_3940,N_3913);
and U4468 (N_4468,N_3843,N_2743);
nor U4469 (N_4469,N_3725,N_3671);
xor U4470 (N_4470,N_3522,N_3977);
and U4471 (N_4471,N_3820,N_3325);
and U4472 (N_4472,N_537,N_1968);
or U4473 (N_4473,N_2351,N_2826);
and U4474 (N_4474,N_3830,N_2058);
xor U4475 (N_4475,N_3808,N_3417);
nand U4476 (N_4476,N_3706,N_2616);
xor U4477 (N_4477,N_3912,N_3633);
or U4478 (N_4478,N_3995,N_3829);
or U4479 (N_4479,In_3344,N_3800);
xor U4480 (N_4480,N_3597,N_2054);
or U4481 (N_4481,N_3991,N_3104);
xor U4482 (N_4482,N_1774,N_3145);
or U4483 (N_4483,N_3975,N_3924);
or U4484 (N_4484,N_3598,In_4503);
or U4485 (N_4485,N_3790,N_3494);
or U4486 (N_4486,N_3669,N_3300);
nand U4487 (N_4487,N_3371,N_3698);
xnor U4488 (N_4488,N_3748,N_3740);
nand U4489 (N_4489,N_1118,N_3784);
nor U4490 (N_4490,N_3563,N_3573);
nand U4491 (N_4491,N_3578,N_514);
xor U4492 (N_4492,N_2674,N_3938);
nor U4493 (N_4493,N_3861,N_3637);
xor U4494 (N_4494,N_3848,N_2228);
nand U4495 (N_4495,N_3046,N_1648);
and U4496 (N_4496,N_3728,N_2904);
nor U4497 (N_4497,N_3519,N_2945);
and U4498 (N_4498,In_877,N_2143);
and U4499 (N_4499,N_3554,N_3448);
xor U4500 (N_4500,N_4330,N_4245);
nand U4501 (N_4501,N_4347,N_4254);
nand U4502 (N_4502,N_4385,N_4241);
xnor U4503 (N_4503,N_4222,N_4300);
or U4504 (N_4504,N_4010,N_4319);
and U4505 (N_4505,N_4184,N_4444);
or U4506 (N_4506,N_4190,N_4028);
nor U4507 (N_4507,N_4482,N_4080);
nand U4508 (N_4508,N_4020,N_4340);
and U4509 (N_4509,N_4109,N_4499);
nand U4510 (N_4510,N_4147,N_4323);
nand U4511 (N_4511,N_4490,N_4469);
and U4512 (N_4512,N_4393,N_4234);
xnor U4513 (N_4513,N_4011,N_4287);
and U4514 (N_4514,N_4327,N_4349);
xor U4515 (N_4515,N_4361,N_4399);
or U4516 (N_4516,N_4076,N_4232);
and U4517 (N_4517,N_4226,N_4397);
nor U4518 (N_4518,N_4157,N_4029);
and U4519 (N_4519,N_4497,N_4178);
nor U4520 (N_4520,N_4125,N_4244);
nor U4521 (N_4521,N_4373,N_4476);
and U4522 (N_4522,N_4128,N_4446);
xor U4523 (N_4523,N_4483,N_4371);
or U4524 (N_4524,N_4098,N_4177);
and U4525 (N_4525,N_4162,N_4105);
or U4526 (N_4526,N_4243,N_4083);
and U4527 (N_4527,N_4293,N_4013);
nand U4528 (N_4528,N_4003,N_4159);
nand U4529 (N_4529,N_4041,N_4206);
and U4530 (N_4530,N_4317,N_4055);
nor U4531 (N_4531,N_4439,N_4416);
nand U4532 (N_4532,N_4285,N_4430);
or U4533 (N_4533,N_4377,N_4237);
nand U4534 (N_4534,N_4119,N_4056);
nand U4535 (N_4535,N_4018,N_4274);
and U4536 (N_4536,N_4321,N_4295);
nor U4537 (N_4537,N_4388,N_4413);
xnor U4538 (N_4538,N_4152,N_4053);
or U4539 (N_4539,N_4242,N_4464);
and U4540 (N_4540,N_4324,N_4459);
nand U4541 (N_4541,N_4224,N_4441);
nand U4542 (N_4542,N_4197,N_4231);
xor U4543 (N_4543,N_4452,N_4332);
nor U4544 (N_4544,N_4326,N_4333);
nor U4545 (N_4545,N_4185,N_4014);
and U4546 (N_4546,N_4468,N_4493);
xnor U4547 (N_4547,N_4392,N_4496);
nand U4548 (N_4548,N_4478,N_4039);
and U4549 (N_4549,N_4114,N_4175);
nor U4550 (N_4550,N_4168,N_4044);
nor U4551 (N_4551,N_4084,N_4428);
nand U4552 (N_4552,N_4087,N_4461);
nor U4553 (N_4553,N_4425,N_4171);
nor U4554 (N_4554,N_4302,N_4221);
nor U4555 (N_4555,N_4498,N_4134);
or U4556 (N_4556,N_4436,N_4307);
xnor U4557 (N_4557,N_4189,N_4336);
or U4558 (N_4558,N_4289,N_4394);
and U4559 (N_4559,N_4412,N_4365);
nand U4560 (N_4560,N_4213,N_4202);
nand U4561 (N_4561,N_4070,N_4270);
nand U4562 (N_4562,N_4142,N_4216);
nor U4563 (N_4563,N_4002,N_4218);
nand U4564 (N_4564,N_4219,N_4081);
nor U4565 (N_4565,N_4346,N_4443);
nor U4566 (N_4566,N_4036,N_4092);
xor U4567 (N_4567,N_4269,N_4144);
nor U4568 (N_4568,N_4402,N_4238);
nand U4569 (N_4569,N_4296,N_4214);
nand U4570 (N_4570,N_4314,N_4453);
and U4571 (N_4571,N_4024,N_4463);
and U4572 (N_4572,N_4192,N_4131);
and U4573 (N_4573,N_4186,N_4170);
and U4574 (N_4574,N_4487,N_4045);
and U4575 (N_4575,N_4350,N_4484);
xor U4576 (N_4576,N_4048,N_4121);
nor U4577 (N_4577,N_4227,N_4093);
and U4578 (N_4578,N_4460,N_4050);
nand U4579 (N_4579,N_4148,N_4380);
or U4580 (N_4580,N_4072,N_4320);
or U4581 (N_4581,N_4208,N_4467);
or U4582 (N_4582,N_4387,N_4127);
nand U4583 (N_4583,N_4337,N_4278);
nand U4584 (N_4584,N_4331,N_4057);
nand U4585 (N_4585,N_4261,N_4384);
xnor U4586 (N_4586,N_4060,N_4089);
nor U4587 (N_4587,N_4160,N_4239);
nand U4588 (N_4588,N_4389,N_4037);
nand U4589 (N_4589,N_4374,N_4075);
and U4590 (N_4590,N_4137,N_4364);
xnor U4591 (N_4591,N_4117,N_4082);
xor U4592 (N_4592,N_4026,N_4079);
nand U4593 (N_4593,N_4471,N_4410);
xor U4594 (N_4594,N_4448,N_4262);
nor U4595 (N_4595,N_4124,N_4292);
xnor U4596 (N_4596,N_4021,N_4187);
and U4597 (N_4597,N_4429,N_4173);
nor U4598 (N_4598,N_4252,N_4115);
nand U4599 (N_4599,N_4205,N_4183);
and U4600 (N_4600,N_4334,N_4091);
xor U4601 (N_4601,N_4251,N_4067);
nand U4602 (N_4602,N_4138,N_4480);
or U4603 (N_4603,N_4063,N_4282);
or U4604 (N_4604,N_4395,N_4312);
nand U4605 (N_4605,N_4267,N_4322);
nor U4606 (N_4606,N_4376,N_4343);
and U4607 (N_4607,N_4090,N_4209);
xor U4608 (N_4608,N_4465,N_4421);
or U4609 (N_4609,N_4313,N_4027);
nand U4610 (N_4610,N_4466,N_4266);
nor U4611 (N_4611,N_4112,N_4225);
or U4612 (N_4612,N_4012,N_4308);
nand U4613 (N_4613,N_4136,N_4404);
nand U4614 (N_4614,N_4167,N_4215);
and U4615 (N_4615,N_4273,N_4309);
nor U4616 (N_4616,N_4193,N_4042);
nand U4617 (N_4617,N_4470,N_4191);
and U4618 (N_4618,N_4212,N_4294);
nor U4619 (N_4619,N_4288,N_4301);
nor U4620 (N_4620,N_4379,N_4263);
nand U4621 (N_4621,N_4182,N_4210);
nand U4622 (N_4622,N_4275,N_4023);
nand U4623 (N_4623,N_4390,N_4486);
or U4624 (N_4624,N_4315,N_4004);
xor U4625 (N_4625,N_4372,N_4103);
and U4626 (N_4626,N_4061,N_4338);
xnor U4627 (N_4627,N_4325,N_4248);
and U4628 (N_4628,N_4479,N_4422);
and U4629 (N_4629,N_4031,N_4154);
or U4630 (N_4630,N_4298,N_4196);
or U4631 (N_4631,N_4113,N_4492);
nand U4632 (N_4632,N_4120,N_4140);
nor U4633 (N_4633,N_4250,N_4040);
xnor U4634 (N_4634,N_4396,N_4353);
nand U4635 (N_4635,N_4247,N_4179);
or U4636 (N_4636,N_4259,N_4007);
or U4637 (N_4637,N_4101,N_4229);
nor U4638 (N_4638,N_4433,N_4155);
xnor U4639 (N_4639,N_4427,N_4068);
and U4640 (N_4640,N_4495,N_4108);
xor U4641 (N_4641,N_4272,N_4458);
and U4642 (N_4642,N_4032,N_4166);
nor U4643 (N_4643,N_4195,N_4064);
or U4644 (N_4644,N_4279,N_4038);
nor U4645 (N_4645,N_4151,N_4475);
xnor U4646 (N_4646,N_4291,N_4025);
or U4647 (N_4647,N_4073,N_4424);
and U4648 (N_4648,N_4329,N_4046);
nand U4649 (N_4649,N_4417,N_4280);
xnor U4650 (N_4650,N_4382,N_4297);
or U4651 (N_4651,N_4409,N_4260);
nor U4652 (N_4652,N_4097,N_4169);
and U4653 (N_4653,N_4065,N_4200);
nand U4654 (N_4654,N_4230,N_4149);
and U4655 (N_4655,N_4123,N_4201);
xnor U4656 (N_4656,N_4375,N_4378);
and U4657 (N_4657,N_4030,N_4366);
xnor U4658 (N_4658,N_4445,N_4203);
nor U4659 (N_4659,N_4369,N_4405);
xnor U4660 (N_4660,N_4406,N_4129);
nor U4661 (N_4661,N_4284,N_4462);
nand U4662 (N_4662,N_4456,N_4344);
and U4663 (N_4663,N_4001,N_4106);
nand U4664 (N_4664,N_4135,N_4249);
nor U4665 (N_4665,N_4059,N_4016);
nand U4666 (N_4666,N_4408,N_4423);
nand U4667 (N_4667,N_4310,N_4420);
nor U4668 (N_4668,N_4095,N_4188);
xor U4669 (N_4669,N_4088,N_4264);
xnor U4670 (N_4670,N_4485,N_4335);
nand U4671 (N_4671,N_4426,N_4198);
xor U4672 (N_4672,N_4246,N_4086);
nor U4673 (N_4673,N_4419,N_4096);
nand U4674 (N_4674,N_4236,N_4360);
xor U4675 (N_4675,N_4000,N_4450);
nor U4676 (N_4676,N_4281,N_4449);
xor U4677 (N_4677,N_4102,N_4122);
nand U4678 (N_4678,N_4199,N_4223);
and U4679 (N_4679,N_4339,N_4477);
nor U4680 (N_4680,N_4303,N_4432);
or U4681 (N_4681,N_4015,N_4342);
nor U4682 (N_4682,N_4165,N_4110);
nand U4683 (N_4683,N_4401,N_4473);
nor U4684 (N_4684,N_4009,N_4368);
or U4685 (N_4685,N_4489,N_4437);
nor U4686 (N_4686,N_4265,N_4431);
xor U4687 (N_4687,N_4176,N_4415);
nor U4688 (N_4688,N_4043,N_4358);
xor U4689 (N_4689,N_4362,N_4447);
and U4690 (N_4690,N_4434,N_4047);
xnor U4691 (N_4691,N_4204,N_4257);
nand U4692 (N_4692,N_4341,N_4194);
and U4693 (N_4693,N_4414,N_4235);
xnor U4694 (N_4694,N_4407,N_4118);
or U4695 (N_4695,N_4107,N_4286);
nor U4696 (N_4696,N_4006,N_4066);
and U4697 (N_4697,N_4156,N_4158);
nand U4698 (N_4698,N_4318,N_4211);
nand U4699 (N_4699,N_4299,N_4049);
nor U4700 (N_4700,N_4164,N_4116);
nand U4701 (N_4701,N_4348,N_4035);
nor U4702 (N_4702,N_4304,N_4276);
xor U4703 (N_4703,N_4034,N_4005);
nor U4704 (N_4704,N_4491,N_4311);
nand U4705 (N_4705,N_4290,N_4058);
nor U4706 (N_4706,N_4181,N_4078);
nor U4707 (N_4707,N_4100,N_4357);
or U4708 (N_4708,N_4367,N_4451);
and U4709 (N_4709,N_4228,N_4139);
and U4710 (N_4710,N_4455,N_4077);
xnor U4711 (N_4711,N_4418,N_4233);
xor U4712 (N_4712,N_4438,N_4017);
or U4713 (N_4713,N_4398,N_4359);
and U4714 (N_4714,N_4180,N_4391);
xnor U4715 (N_4715,N_4435,N_4411);
xnor U4716 (N_4716,N_4474,N_4132);
nor U4717 (N_4717,N_4381,N_4345);
xnor U4718 (N_4718,N_4283,N_4240);
xor U4719 (N_4719,N_4255,N_4019);
nor U4720 (N_4720,N_4069,N_4104);
and U4721 (N_4721,N_4054,N_4305);
nor U4722 (N_4722,N_4085,N_4494);
xnor U4723 (N_4723,N_4472,N_4442);
xnor U4724 (N_4724,N_4094,N_4133);
xor U4725 (N_4725,N_4363,N_4440);
nand U4726 (N_4726,N_4268,N_4008);
and U4727 (N_4727,N_4271,N_4174);
nand U4728 (N_4728,N_4033,N_4386);
and U4729 (N_4729,N_4454,N_4403);
xnor U4730 (N_4730,N_4488,N_4153);
and U4731 (N_4731,N_4253,N_4126);
xor U4732 (N_4732,N_4099,N_4143);
and U4733 (N_4733,N_4217,N_4258);
nor U4734 (N_4734,N_4356,N_4355);
or U4735 (N_4735,N_4163,N_4150);
xor U4736 (N_4736,N_4352,N_4022);
nand U4737 (N_4737,N_4111,N_4145);
xor U4738 (N_4738,N_4146,N_4161);
or U4739 (N_4739,N_4052,N_4481);
and U4740 (N_4740,N_4400,N_4051);
or U4741 (N_4741,N_4354,N_4074);
nand U4742 (N_4742,N_4062,N_4351);
nand U4743 (N_4743,N_4130,N_4172);
and U4744 (N_4744,N_4457,N_4256);
nor U4745 (N_4745,N_4141,N_4071);
or U4746 (N_4746,N_4383,N_4277);
xor U4747 (N_4747,N_4316,N_4328);
and U4748 (N_4748,N_4207,N_4306);
or U4749 (N_4749,N_4220,N_4370);
nand U4750 (N_4750,N_4045,N_4469);
nor U4751 (N_4751,N_4233,N_4437);
nand U4752 (N_4752,N_4215,N_4150);
xor U4753 (N_4753,N_4492,N_4349);
nand U4754 (N_4754,N_4205,N_4236);
and U4755 (N_4755,N_4324,N_4162);
nand U4756 (N_4756,N_4025,N_4066);
or U4757 (N_4757,N_4414,N_4154);
and U4758 (N_4758,N_4383,N_4389);
or U4759 (N_4759,N_4030,N_4330);
nand U4760 (N_4760,N_4014,N_4328);
nand U4761 (N_4761,N_4179,N_4203);
xor U4762 (N_4762,N_4390,N_4041);
and U4763 (N_4763,N_4460,N_4174);
and U4764 (N_4764,N_4147,N_4356);
nor U4765 (N_4765,N_4159,N_4422);
and U4766 (N_4766,N_4387,N_4369);
nor U4767 (N_4767,N_4139,N_4081);
nand U4768 (N_4768,N_4345,N_4374);
xor U4769 (N_4769,N_4147,N_4212);
or U4770 (N_4770,N_4385,N_4329);
nor U4771 (N_4771,N_4098,N_4340);
or U4772 (N_4772,N_4097,N_4396);
or U4773 (N_4773,N_4311,N_4125);
xor U4774 (N_4774,N_4417,N_4334);
and U4775 (N_4775,N_4180,N_4122);
and U4776 (N_4776,N_4254,N_4482);
or U4777 (N_4777,N_4345,N_4375);
nor U4778 (N_4778,N_4295,N_4181);
or U4779 (N_4779,N_4343,N_4348);
and U4780 (N_4780,N_4065,N_4459);
xor U4781 (N_4781,N_4195,N_4369);
or U4782 (N_4782,N_4085,N_4052);
or U4783 (N_4783,N_4218,N_4376);
and U4784 (N_4784,N_4282,N_4438);
or U4785 (N_4785,N_4151,N_4334);
nor U4786 (N_4786,N_4399,N_4308);
and U4787 (N_4787,N_4104,N_4145);
xnor U4788 (N_4788,N_4074,N_4338);
xnor U4789 (N_4789,N_4294,N_4273);
nand U4790 (N_4790,N_4262,N_4237);
or U4791 (N_4791,N_4357,N_4211);
or U4792 (N_4792,N_4388,N_4120);
nand U4793 (N_4793,N_4173,N_4376);
or U4794 (N_4794,N_4468,N_4184);
and U4795 (N_4795,N_4193,N_4160);
or U4796 (N_4796,N_4157,N_4346);
or U4797 (N_4797,N_4420,N_4439);
nor U4798 (N_4798,N_4365,N_4070);
nor U4799 (N_4799,N_4359,N_4411);
and U4800 (N_4800,N_4267,N_4427);
nand U4801 (N_4801,N_4081,N_4353);
or U4802 (N_4802,N_4269,N_4431);
and U4803 (N_4803,N_4208,N_4249);
nor U4804 (N_4804,N_4247,N_4169);
nand U4805 (N_4805,N_4022,N_4038);
and U4806 (N_4806,N_4162,N_4055);
and U4807 (N_4807,N_4442,N_4428);
and U4808 (N_4808,N_4055,N_4315);
nand U4809 (N_4809,N_4142,N_4350);
or U4810 (N_4810,N_4274,N_4337);
nor U4811 (N_4811,N_4250,N_4201);
and U4812 (N_4812,N_4181,N_4416);
nand U4813 (N_4813,N_4411,N_4419);
xor U4814 (N_4814,N_4005,N_4057);
nand U4815 (N_4815,N_4049,N_4416);
or U4816 (N_4816,N_4482,N_4464);
nand U4817 (N_4817,N_4290,N_4097);
or U4818 (N_4818,N_4050,N_4237);
nand U4819 (N_4819,N_4252,N_4352);
nand U4820 (N_4820,N_4009,N_4422);
nor U4821 (N_4821,N_4494,N_4433);
xor U4822 (N_4822,N_4269,N_4467);
nor U4823 (N_4823,N_4220,N_4262);
or U4824 (N_4824,N_4133,N_4369);
nor U4825 (N_4825,N_4362,N_4317);
and U4826 (N_4826,N_4129,N_4271);
xnor U4827 (N_4827,N_4020,N_4313);
xnor U4828 (N_4828,N_4272,N_4175);
xor U4829 (N_4829,N_4357,N_4118);
xor U4830 (N_4830,N_4059,N_4119);
xor U4831 (N_4831,N_4449,N_4247);
or U4832 (N_4832,N_4261,N_4355);
nand U4833 (N_4833,N_4378,N_4452);
and U4834 (N_4834,N_4394,N_4337);
and U4835 (N_4835,N_4128,N_4105);
xnor U4836 (N_4836,N_4106,N_4493);
xor U4837 (N_4837,N_4144,N_4053);
xor U4838 (N_4838,N_4373,N_4421);
xor U4839 (N_4839,N_4287,N_4393);
xnor U4840 (N_4840,N_4310,N_4410);
xnor U4841 (N_4841,N_4192,N_4364);
or U4842 (N_4842,N_4096,N_4495);
xnor U4843 (N_4843,N_4469,N_4394);
nand U4844 (N_4844,N_4464,N_4077);
xor U4845 (N_4845,N_4063,N_4209);
nor U4846 (N_4846,N_4231,N_4085);
xor U4847 (N_4847,N_4443,N_4436);
xor U4848 (N_4848,N_4393,N_4316);
xor U4849 (N_4849,N_4092,N_4473);
nand U4850 (N_4850,N_4242,N_4467);
and U4851 (N_4851,N_4025,N_4118);
xor U4852 (N_4852,N_4367,N_4200);
nor U4853 (N_4853,N_4056,N_4210);
nor U4854 (N_4854,N_4287,N_4309);
xor U4855 (N_4855,N_4043,N_4171);
nor U4856 (N_4856,N_4427,N_4467);
and U4857 (N_4857,N_4160,N_4104);
or U4858 (N_4858,N_4491,N_4315);
nor U4859 (N_4859,N_4267,N_4067);
nand U4860 (N_4860,N_4327,N_4205);
nand U4861 (N_4861,N_4374,N_4104);
nand U4862 (N_4862,N_4322,N_4435);
or U4863 (N_4863,N_4420,N_4370);
nand U4864 (N_4864,N_4154,N_4085);
xor U4865 (N_4865,N_4123,N_4035);
nor U4866 (N_4866,N_4401,N_4316);
nand U4867 (N_4867,N_4373,N_4089);
nor U4868 (N_4868,N_4227,N_4218);
nand U4869 (N_4869,N_4052,N_4109);
nor U4870 (N_4870,N_4320,N_4311);
and U4871 (N_4871,N_4078,N_4075);
or U4872 (N_4872,N_4261,N_4241);
nor U4873 (N_4873,N_4087,N_4256);
xor U4874 (N_4874,N_4140,N_4364);
nor U4875 (N_4875,N_4160,N_4363);
xor U4876 (N_4876,N_4016,N_4418);
nand U4877 (N_4877,N_4206,N_4222);
and U4878 (N_4878,N_4356,N_4296);
or U4879 (N_4879,N_4292,N_4060);
nor U4880 (N_4880,N_4224,N_4397);
xor U4881 (N_4881,N_4399,N_4046);
or U4882 (N_4882,N_4051,N_4093);
xnor U4883 (N_4883,N_4386,N_4451);
or U4884 (N_4884,N_4404,N_4098);
or U4885 (N_4885,N_4084,N_4057);
or U4886 (N_4886,N_4175,N_4209);
and U4887 (N_4887,N_4001,N_4078);
nor U4888 (N_4888,N_4375,N_4275);
xor U4889 (N_4889,N_4406,N_4254);
nand U4890 (N_4890,N_4146,N_4426);
or U4891 (N_4891,N_4118,N_4348);
nand U4892 (N_4892,N_4197,N_4164);
xnor U4893 (N_4893,N_4027,N_4291);
xnor U4894 (N_4894,N_4277,N_4347);
xnor U4895 (N_4895,N_4063,N_4383);
or U4896 (N_4896,N_4139,N_4297);
xor U4897 (N_4897,N_4187,N_4302);
and U4898 (N_4898,N_4480,N_4061);
and U4899 (N_4899,N_4148,N_4136);
nor U4900 (N_4900,N_4260,N_4105);
xnor U4901 (N_4901,N_4174,N_4154);
xor U4902 (N_4902,N_4344,N_4389);
nor U4903 (N_4903,N_4242,N_4076);
nor U4904 (N_4904,N_4404,N_4033);
nor U4905 (N_4905,N_4021,N_4207);
and U4906 (N_4906,N_4184,N_4043);
and U4907 (N_4907,N_4237,N_4151);
xor U4908 (N_4908,N_4349,N_4470);
and U4909 (N_4909,N_4032,N_4315);
nand U4910 (N_4910,N_4000,N_4345);
xnor U4911 (N_4911,N_4231,N_4348);
and U4912 (N_4912,N_4382,N_4437);
or U4913 (N_4913,N_4274,N_4040);
and U4914 (N_4914,N_4114,N_4445);
and U4915 (N_4915,N_4194,N_4347);
xnor U4916 (N_4916,N_4258,N_4413);
or U4917 (N_4917,N_4305,N_4214);
xor U4918 (N_4918,N_4428,N_4490);
xor U4919 (N_4919,N_4372,N_4345);
nand U4920 (N_4920,N_4409,N_4011);
nand U4921 (N_4921,N_4220,N_4243);
or U4922 (N_4922,N_4075,N_4393);
nand U4923 (N_4923,N_4075,N_4034);
xnor U4924 (N_4924,N_4065,N_4326);
nand U4925 (N_4925,N_4218,N_4239);
nand U4926 (N_4926,N_4085,N_4144);
xor U4927 (N_4927,N_4048,N_4236);
nand U4928 (N_4928,N_4012,N_4051);
nand U4929 (N_4929,N_4330,N_4242);
and U4930 (N_4930,N_4085,N_4053);
and U4931 (N_4931,N_4381,N_4421);
or U4932 (N_4932,N_4076,N_4387);
and U4933 (N_4933,N_4311,N_4052);
nor U4934 (N_4934,N_4176,N_4152);
xor U4935 (N_4935,N_4418,N_4268);
nor U4936 (N_4936,N_4118,N_4193);
or U4937 (N_4937,N_4256,N_4084);
xor U4938 (N_4938,N_4428,N_4110);
nand U4939 (N_4939,N_4459,N_4298);
nor U4940 (N_4940,N_4303,N_4461);
nor U4941 (N_4941,N_4388,N_4130);
nand U4942 (N_4942,N_4356,N_4403);
xnor U4943 (N_4943,N_4129,N_4260);
nand U4944 (N_4944,N_4156,N_4248);
or U4945 (N_4945,N_4279,N_4043);
nor U4946 (N_4946,N_4475,N_4166);
and U4947 (N_4947,N_4359,N_4309);
xnor U4948 (N_4948,N_4151,N_4176);
and U4949 (N_4949,N_4344,N_4361);
or U4950 (N_4950,N_4287,N_4017);
nor U4951 (N_4951,N_4128,N_4492);
and U4952 (N_4952,N_4379,N_4479);
nand U4953 (N_4953,N_4197,N_4441);
nor U4954 (N_4954,N_4420,N_4270);
nand U4955 (N_4955,N_4126,N_4127);
nor U4956 (N_4956,N_4147,N_4182);
and U4957 (N_4957,N_4389,N_4378);
xor U4958 (N_4958,N_4112,N_4431);
nand U4959 (N_4959,N_4122,N_4377);
xnor U4960 (N_4960,N_4194,N_4460);
or U4961 (N_4961,N_4084,N_4126);
xnor U4962 (N_4962,N_4003,N_4371);
nand U4963 (N_4963,N_4292,N_4382);
nor U4964 (N_4964,N_4081,N_4039);
and U4965 (N_4965,N_4293,N_4058);
nor U4966 (N_4966,N_4077,N_4230);
nor U4967 (N_4967,N_4302,N_4132);
and U4968 (N_4968,N_4333,N_4028);
xor U4969 (N_4969,N_4077,N_4437);
and U4970 (N_4970,N_4468,N_4481);
xnor U4971 (N_4971,N_4297,N_4414);
and U4972 (N_4972,N_4352,N_4174);
nor U4973 (N_4973,N_4302,N_4254);
nand U4974 (N_4974,N_4158,N_4342);
xnor U4975 (N_4975,N_4447,N_4121);
nor U4976 (N_4976,N_4008,N_4045);
or U4977 (N_4977,N_4115,N_4060);
xnor U4978 (N_4978,N_4389,N_4380);
nand U4979 (N_4979,N_4117,N_4088);
nand U4980 (N_4980,N_4497,N_4430);
or U4981 (N_4981,N_4065,N_4313);
or U4982 (N_4982,N_4428,N_4300);
nand U4983 (N_4983,N_4067,N_4380);
or U4984 (N_4984,N_4387,N_4061);
nand U4985 (N_4985,N_4334,N_4317);
and U4986 (N_4986,N_4320,N_4109);
xnor U4987 (N_4987,N_4148,N_4468);
or U4988 (N_4988,N_4253,N_4208);
and U4989 (N_4989,N_4254,N_4183);
nor U4990 (N_4990,N_4259,N_4065);
or U4991 (N_4991,N_4341,N_4337);
and U4992 (N_4992,N_4060,N_4086);
nand U4993 (N_4993,N_4252,N_4060);
xnor U4994 (N_4994,N_4459,N_4343);
nor U4995 (N_4995,N_4446,N_4011);
nand U4996 (N_4996,N_4098,N_4333);
nand U4997 (N_4997,N_4136,N_4217);
or U4998 (N_4998,N_4323,N_4347);
nor U4999 (N_4999,N_4116,N_4216);
or U5000 (N_5000,N_4629,N_4720);
nand U5001 (N_5001,N_4699,N_4694);
or U5002 (N_5002,N_4973,N_4938);
nor U5003 (N_5003,N_4724,N_4965);
nor U5004 (N_5004,N_4529,N_4588);
nor U5005 (N_5005,N_4651,N_4516);
and U5006 (N_5006,N_4502,N_4533);
and U5007 (N_5007,N_4759,N_4542);
nor U5008 (N_5008,N_4803,N_4886);
or U5009 (N_5009,N_4646,N_4754);
and U5010 (N_5010,N_4524,N_4895);
or U5011 (N_5011,N_4961,N_4619);
nand U5012 (N_5012,N_4781,N_4547);
nand U5013 (N_5013,N_4732,N_4689);
nand U5014 (N_5014,N_4986,N_4608);
xor U5015 (N_5015,N_4728,N_4537);
or U5016 (N_5016,N_4826,N_4650);
nand U5017 (N_5017,N_4740,N_4985);
or U5018 (N_5018,N_4791,N_4702);
nand U5019 (N_5019,N_4868,N_4814);
nand U5020 (N_5020,N_4628,N_4823);
nor U5021 (N_5021,N_4565,N_4851);
or U5022 (N_5022,N_4648,N_4804);
and U5023 (N_5023,N_4585,N_4596);
nand U5024 (N_5024,N_4854,N_4794);
nor U5025 (N_5025,N_4857,N_4856);
nor U5026 (N_5026,N_4654,N_4936);
nand U5027 (N_5027,N_4848,N_4891);
nand U5028 (N_5028,N_4786,N_4534);
nand U5029 (N_5029,N_4815,N_4785);
nand U5030 (N_5030,N_4704,N_4896);
nor U5031 (N_5031,N_4575,N_4977);
nor U5032 (N_5032,N_4697,N_4945);
nor U5033 (N_5033,N_4976,N_4601);
xnor U5034 (N_5034,N_4538,N_4679);
nand U5035 (N_5035,N_4739,N_4706);
nand U5036 (N_5036,N_4636,N_4507);
and U5037 (N_5037,N_4951,N_4899);
or U5038 (N_5038,N_4933,N_4782);
and U5039 (N_5039,N_4989,N_4784);
or U5040 (N_5040,N_4701,N_4847);
xnor U5041 (N_5041,N_4626,N_4586);
and U5042 (N_5042,N_4764,N_4672);
or U5043 (N_5043,N_4966,N_4902);
nand U5044 (N_5044,N_4621,N_4705);
xor U5045 (N_5045,N_4684,N_4605);
nor U5046 (N_5046,N_4535,N_4816);
nor U5047 (N_5047,N_4944,N_4540);
nor U5048 (N_5048,N_4971,N_4526);
and U5049 (N_5049,N_4780,N_4836);
xor U5050 (N_5050,N_4578,N_4914);
and U5051 (N_5051,N_4934,N_4674);
nor U5052 (N_5052,N_4683,N_4927);
nor U5053 (N_5053,N_4928,N_4910);
xor U5054 (N_5054,N_4911,N_4801);
nand U5055 (N_5055,N_4503,N_4835);
nor U5056 (N_5056,N_4760,N_4504);
xnor U5057 (N_5057,N_4962,N_4845);
nand U5058 (N_5058,N_4758,N_4591);
nand U5059 (N_5059,N_4680,N_4984);
or U5060 (N_5060,N_4752,N_4594);
or U5061 (N_5061,N_4630,N_4888);
or U5062 (N_5062,N_4867,N_4866);
nor U5063 (N_5063,N_4963,N_4772);
or U5064 (N_5064,N_4611,N_4862);
or U5065 (N_5065,N_4665,N_4900);
and U5066 (N_5066,N_4842,N_4713);
or U5067 (N_5067,N_4964,N_4508);
and U5068 (N_5068,N_4572,N_4799);
nand U5069 (N_5069,N_4841,N_4743);
xor U5070 (N_5070,N_4860,N_4746);
nor U5071 (N_5071,N_4511,N_4510);
nand U5072 (N_5072,N_4873,N_4916);
nor U5073 (N_5073,N_4885,N_4741);
xnor U5074 (N_5074,N_4663,N_4771);
xor U5075 (N_5075,N_4956,N_4880);
and U5076 (N_5076,N_4818,N_4970);
nor U5077 (N_5077,N_4929,N_4921);
or U5078 (N_5078,N_4620,N_4649);
or U5079 (N_5079,N_4906,N_4988);
or U5080 (N_5080,N_4573,N_4755);
or U5081 (N_5081,N_4882,N_4756);
nor U5082 (N_5082,N_4864,N_4632);
nor U5083 (N_5083,N_4641,N_4872);
xor U5084 (N_5084,N_4924,N_4523);
nor U5085 (N_5085,N_4981,N_4750);
nand U5086 (N_5086,N_4948,N_4825);
xnor U5087 (N_5087,N_4564,N_4673);
nor U5088 (N_5088,N_4676,N_4528);
xnor U5089 (N_5089,N_4567,N_4513);
nand U5090 (N_5090,N_4656,N_4747);
and U5091 (N_5091,N_4990,N_4576);
nand U5092 (N_5092,N_4797,N_4718);
xor U5093 (N_5093,N_4558,N_4789);
xor U5094 (N_5094,N_4995,N_4822);
nor U5095 (N_5095,N_4942,N_4839);
xor U5096 (N_5096,N_4837,N_4686);
nor U5097 (N_5097,N_4774,N_4670);
or U5098 (N_5098,N_4505,N_4552);
and U5099 (N_5099,N_4668,N_4725);
or U5100 (N_5100,N_4590,N_4999);
and U5101 (N_5101,N_4580,N_4691);
nand U5102 (N_5102,N_4553,N_4824);
nand U5103 (N_5103,N_4644,N_4883);
and U5104 (N_5104,N_4708,N_4931);
xnor U5105 (N_5105,N_4768,N_4647);
xor U5106 (N_5106,N_4993,N_4833);
nor U5107 (N_5107,N_4954,N_4871);
xor U5108 (N_5108,N_4521,N_4881);
nor U5109 (N_5109,N_4737,N_4821);
nand U5110 (N_5110,N_4714,N_4863);
xnor U5111 (N_5111,N_4742,N_4918);
nand U5112 (N_5112,N_4778,N_4582);
nand U5113 (N_5113,N_4829,N_4522);
nor U5114 (N_5114,N_4678,N_4861);
and U5115 (N_5115,N_4587,N_4852);
xnor U5116 (N_5116,N_4531,N_4884);
xor U5117 (N_5117,N_4597,N_4696);
xnor U5118 (N_5118,N_4710,N_4827);
and U5119 (N_5119,N_4796,N_4666);
and U5120 (N_5120,N_4579,N_4667);
nor U5121 (N_5121,N_4645,N_4727);
and U5122 (N_5122,N_4959,N_4753);
xnor U5123 (N_5123,N_4834,N_4612);
xor U5124 (N_5124,N_4787,N_4769);
nand U5125 (N_5125,N_4849,N_4717);
xor U5126 (N_5126,N_4569,N_4606);
xor U5127 (N_5127,N_4947,N_4655);
nor U5128 (N_5128,N_4744,N_4726);
nor U5129 (N_5129,N_4729,N_4887);
or U5130 (N_5130,N_4767,N_4811);
and U5131 (N_5131,N_4719,N_4721);
nor U5132 (N_5132,N_4926,N_4898);
nor U5133 (N_5133,N_4935,N_4905);
and U5134 (N_5134,N_4643,N_4736);
or U5135 (N_5135,N_4978,N_4994);
nand U5136 (N_5136,N_4876,N_4917);
nor U5137 (N_5137,N_4637,N_4979);
nand U5138 (N_5138,N_4991,N_4879);
nor U5139 (N_5139,N_4525,N_4583);
nand U5140 (N_5140,N_4904,N_4890);
nor U5141 (N_5141,N_4806,N_4574);
xnor U5142 (N_5142,N_4541,N_4707);
nor U5143 (N_5143,N_4539,N_4869);
and U5144 (N_5144,N_4844,N_4997);
and U5145 (N_5145,N_4603,N_4878);
nor U5146 (N_5146,N_4716,N_4775);
xnor U5147 (N_5147,N_4681,N_4763);
or U5148 (N_5148,N_4703,N_4974);
nand U5149 (N_5149,N_4692,N_4949);
nor U5150 (N_5150,N_4544,N_4698);
nand U5151 (N_5151,N_4709,N_4773);
or U5152 (N_5152,N_4820,N_4635);
xor U5153 (N_5153,N_4599,N_4802);
nor U5154 (N_5154,N_4500,N_4874);
nand U5155 (N_5155,N_4515,N_4577);
nor U5156 (N_5156,N_4658,N_4996);
nor U5157 (N_5157,N_4512,N_4613);
nor U5158 (N_5158,N_4711,N_4687);
nor U5159 (N_5159,N_4623,N_4568);
and U5160 (N_5160,N_4618,N_4519);
or U5161 (N_5161,N_4514,N_4897);
and U5162 (N_5162,N_4749,N_4671);
xor U5163 (N_5163,N_4602,N_4915);
and U5164 (N_5164,N_4757,N_4909);
nand U5165 (N_5165,N_4738,N_4893);
nand U5166 (N_5166,N_4952,N_4660);
xor U5167 (N_5167,N_4627,N_4817);
or U5168 (N_5168,N_4664,N_4566);
nor U5169 (N_5169,N_4501,N_4960);
xnor U5170 (N_5170,N_4735,N_4634);
xnor U5171 (N_5171,N_4604,N_4748);
xnor U5172 (N_5172,N_4751,N_4913);
or U5173 (N_5173,N_4761,N_4930);
xnor U5174 (N_5174,N_4563,N_4831);
nand U5175 (N_5175,N_4555,N_4581);
or U5176 (N_5176,N_4551,N_4809);
nor U5177 (N_5177,N_4722,N_4682);
nor U5178 (N_5178,N_4607,N_4685);
nor U5179 (N_5179,N_4932,N_4617);
nor U5180 (N_5180,N_4830,N_4571);
and U5181 (N_5181,N_4908,N_4765);
xnor U5182 (N_5182,N_4777,N_4652);
xnor U5183 (N_5183,N_4638,N_4907);
nor U5184 (N_5184,N_4950,N_4939);
xnor U5185 (N_5185,N_4762,N_4943);
or U5186 (N_5186,N_4832,N_4788);
xor U5187 (N_5187,N_4559,N_4598);
and U5188 (N_5188,N_4920,N_4792);
xnor U5189 (N_5189,N_4624,N_4813);
nand U5190 (N_5190,N_4520,N_4779);
and U5191 (N_5191,N_4838,N_4631);
or U5192 (N_5192,N_4807,N_4955);
nand U5193 (N_5193,N_4610,N_4870);
nand U5194 (N_5194,N_4790,N_4912);
xor U5195 (N_5195,N_4600,N_4662);
nand U5196 (N_5196,N_4730,N_4892);
xnor U5197 (N_5197,N_4690,N_4987);
and U5198 (N_5198,N_4975,N_4509);
or U5199 (N_5199,N_4642,N_4615);
and U5200 (N_5200,N_4998,N_4875);
xnor U5201 (N_5201,N_4903,N_4640);
nor U5202 (N_5202,N_4653,N_4633);
nor U5203 (N_5203,N_4967,N_4592);
and U5204 (N_5204,N_4850,N_4693);
and U5205 (N_5205,N_4946,N_4570);
nand U5206 (N_5206,N_4625,N_4715);
nor U5207 (N_5207,N_4554,N_4941);
nor U5208 (N_5208,N_4622,N_4734);
or U5209 (N_5209,N_4609,N_4828);
and U5210 (N_5210,N_4543,N_4783);
xor U5211 (N_5211,N_4506,N_4853);
or U5212 (N_5212,N_4661,N_4695);
xor U5213 (N_5213,N_4840,N_4901);
and U5214 (N_5214,N_4530,N_4675);
nor U5215 (N_5215,N_4770,N_4595);
xor U5216 (N_5216,N_4982,N_4969);
nand U5217 (N_5217,N_4557,N_4798);
nand U5218 (N_5218,N_4843,N_4894);
and U5219 (N_5219,N_4808,N_4614);
or U5220 (N_5220,N_4657,N_4937);
xnor U5221 (N_5221,N_4527,N_4688);
nor U5222 (N_5222,N_4919,N_4733);
xnor U5223 (N_5223,N_4923,N_4865);
or U5224 (N_5224,N_4855,N_4712);
and U5225 (N_5225,N_4561,N_4972);
nor U5226 (N_5226,N_4980,N_4925);
xor U5227 (N_5227,N_4846,N_4745);
or U5228 (N_5228,N_4819,N_4793);
nand U5229 (N_5229,N_4677,N_4957);
and U5230 (N_5230,N_4669,N_4731);
or U5231 (N_5231,N_4639,N_4795);
nand U5232 (N_5232,N_4536,N_4548);
and U5233 (N_5233,N_4560,N_4958);
or U5234 (N_5234,N_4518,N_4858);
or U5235 (N_5235,N_4723,N_4940);
nand U5236 (N_5236,N_4659,N_4616);
and U5237 (N_5237,N_4545,N_4922);
or U5238 (N_5238,N_4766,N_4983);
or U5239 (N_5239,N_4992,N_4546);
and U5240 (N_5240,N_4968,N_4700);
or U5241 (N_5241,N_4805,N_4549);
nand U5242 (N_5242,N_4810,N_4800);
and U5243 (N_5243,N_4550,N_4593);
nand U5244 (N_5244,N_4889,N_4812);
xnor U5245 (N_5245,N_4517,N_4776);
nand U5246 (N_5246,N_4859,N_4584);
nor U5247 (N_5247,N_4556,N_4877);
nor U5248 (N_5248,N_4953,N_4532);
and U5249 (N_5249,N_4589,N_4562);
and U5250 (N_5250,N_4574,N_4614);
xor U5251 (N_5251,N_4977,N_4656);
nor U5252 (N_5252,N_4548,N_4521);
xnor U5253 (N_5253,N_4727,N_4757);
xor U5254 (N_5254,N_4614,N_4536);
or U5255 (N_5255,N_4699,N_4727);
and U5256 (N_5256,N_4528,N_4985);
nor U5257 (N_5257,N_4793,N_4966);
xnor U5258 (N_5258,N_4522,N_4667);
or U5259 (N_5259,N_4581,N_4708);
xnor U5260 (N_5260,N_4628,N_4843);
nor U5261 (N_5261,N_4558,N_4668);
or U5262 (N_5262,N_4763,N_4780);
xor U5263 (N_5263,N_4794,N_4732);
nand U5264 (N_5264,N_4670,N_4917);
nand U5265 (N_5265,N_4508,N_4547);
xor U5266 (N_5266,N_4697,N_4639);
nor U5267 (N_5267,N_4925,N_4881);
or U5268 (N_5268,N_4708,N_4960);
xnor U5269 (N_5269,N_4599,N_4905);
xor U5270 (N_5270,N_4878,N_4969);
and U5271 (N_5271,N_4847,N_4704);
or U5272 (N_5272,N_4726,N_4863);
or U5273 (N_5273,N_4833,N_4510);
and U5274 (N_5274,N_4896,N_4557);
and U5275 (N_5275,N_4930,N_4569);
xor U5276 (N_5276,N_4930,N_4921);
and U5277 (N_5277,N_4753,N_4666);
nor U5278 (N_5278,N_4569,N_4658);
nand U5279 (N_5279,N_4941,N_4871);
and U5280 (N_5280,N_4555,N_4502);
nand U5281 (N_5281,N_4674,N_4900);
and U5282 (N_5282,N_4847,N_4771);
or U5283 (N_5283,N_4713,N_4851);
or U5284 (N_5284,N_4698,N_4889);
nor U5285 (N_5285,N_4632,N_4612);
or U5286 (N_5286,N_4502,N_4952);
xnor U5287 (N_5287,N_4749,N_4646);
nand U5288 (N_5288,N_4755,N_4694);
or U5289 (N_5289,N_4955,N_4783);
xnor U5290 (N_5290,N_4753,N_4912);
nand U5291 (N_5291,N_4939,N_4879);
and U5292 (N_5292,N_4931,N_4786);
xor U5293 (N_5293,N_4834,N_4804);
or U5294 (N_5294,N_4627,N_4820);
nand U5295 (N_5295,N_4681,N_4740);
or U5296 (N_5296,N_4673,N_4883);
nor U5297 (N_5297,N_4817,N_4801);
xnor U5298 (N_5298,N_4693,N_4662);
and U5299 (N_5299,N_4830,N_4593);
nand U5300 (N_5300,N_4962,N_4794);
and U5301 (N_5301,N_4844,N_4836);
nand U5302 (N_5302,N_4965,N_4761);
or U5303 (N_5303,N_4778,N_4596);
or U5304 (N_5304,N_4958,N_4765);
and U5305 (N_5305,N_4671,N_4943);
xor U5306 (N_5306,N_4599,N_4745);
or U5307 (N_5307,N_4761,N_4959);
nor U5308 (N_5308,N_4726,N_4971);
xnor U5309 (N_5309,N_4791,N_4652);
nor U5310 (N_5310,N_4975,N_4815);
nand U5311 (N_5311,N_4639,N_4631);
or U5312 (N_5312,N_4570,N_4581);
xnor U5313 (N_5313,N_4872,N_4913);
xnor U5314 (N_5314,N_4634,N_4860);
or U5315 (N_5315,N_4516,N_4830);
or U5316 (N_5316,N_4647,N_4729);
or U5317 (N_5317,N_4980,N_4736);
and U5318 (N_5318,N_4963,N_4572);
xnor U5319 (N_5319,N_4519,N_4879);
xnor U5320 (N_5320,N_4789,N_4538);
nand U5321 (N_5321,N_4706,N_4897);
or U5322 (N_5322,N_4692,N_4573);
xor U5323 (N_5323,N_4789,N_4817);
nand U5324 (N_5324,N_4922,N_4550);
nor U5325 (N_5325,N_4623,N_4917);
and U5326 (N_5326,N_4511,N_4521);
and U5327 (N_5327,N_4676,N_4727);
or U5328 (N_5328,N_4847,N_4515);
nor U5329 (N_5329,N_4777,N_4956);
and U5330 (N_5330,N_4690,N_4899);
and U5331 (N_5331,N_4535,N_4580);
nand U5332 (N_5332,N_4958,N_4651);
xnor U5333 (N_5333,N_4702,N_4800);
xnor U5334 (N_5334,N_4775,N_4907);
or U5335 (N_5335,N_4875,N_4828);
nand U5336 (N_5336,N_4761,N_4697);
nand U5337 (N_5337,N_4881,N_4598);
nand U5338 (N_5338,N_4659,N_4504);
nand U5339 (N_5339,N_4754,N_4703);
xor U5340 (N_5340,N_4650,N_4855);
nand U5341 (N_5341,N_4908,N_4675);
xnor U5342 (N_5342,N_4779,N_4500);
nor U5343 (N_5343,N_4708,N_4672);
nand U5344 (N_5344,N_4743,N_4662);
nor U5345 (N_5345,N_4530,N_4897);
nand U5346 (N_5346,N_4748,N_4545);
xnor U5347 (N_5347,N_4580,N_4614);
nor U5348 (N_5348,N_4991,N_4876);
xor U5349 (N_5349,N_4759,N_4529);
or U5350 (N_5350,N_4962,N_4592);
nand U5351 (N_5351,N_4971,N_4710);
xor U5352 (N_5352,N_4658,N_4547);
xnor U5353 (N_5353,N_4992,N_4694);
and U5354 (N_5354,N_4678,N_4896);
and U5355 (N_5355,N_4951,N_4666);
and U5356 (N_5356,N_4639,N_4574);
xor U5357 (N_5357,N_4913,N_4868);
and U5358 (N_5358,N_4963,N_4849);
nor U5359 (N_5359,N_4549,N_4709);
nor U5360 (N_5360,N_4860,N_4919);
and U5361 (N_5361,N_4930,N_4841);
xnor U5362 (N_5362,N_4598,N_4948);
xor U5363 (N_5363,N_4739,N_4836);
nor U5364 (N_5364,N_4650,N_4807);
and U5365 (N_5365,N_4558,N_4597);
nand U5366 (N_5366,N_4592,N_4831);
xnor U5367 (N_5367,N_4502,N_4594);
or U5368 (N_5368,N_4502,N_4916);
nand U5369 (N_5369,N_4589,N_4735);
nand U5370 (N_5370,N_4891,N_4715);
nand U5371 (N_5371,N_4652,N_4772);
or U5372 (N_5372,N_4530,N_4814);
xor U5373 (N_5373,N_4888,N_4872);
nand U5374 (N_5374,N_4649,N_4500);
xor U5375 (N_5375,N_4662,N_4818);
and U5376 (N_5376,N_4532,N_4720);
nor U5377 (N_5377,N_4946,N_4824);
or U5378 (N_5378,N_4848,N_4972);
and U5379 (N_5379,N_4672,N_4733);
nor U5380 (N_5380,N_4708,N_4527);
nor U5381 (N_5381,N_4863,N_4607);
nor U5382 (N_5382,N_4930,N_4822);
nor U5383 (N_5383,N_4846,N_4597);
nand U5384 (N_5384,N_4748,N_4953);
xnor U5385 (N_5385,N_4862,N_4753);
nor U5386 (N_5386,N_4587,N_4575);
nor U5387 (N_5387,N_4988,N_4911);
nand U5388 (N_5388,N_4709,N_4944);
and U5389 (N_5389,N_4977,N_4713);
xnor U5390 (N_5390,N_4961,N_4892);
and U5391 (N_5391,N_4826,N_4636);
xnor U5392 (N_5392,N_4831,N_4716);
and U5393 (N_5393,N_4834,N_4859);
nand U5394 (N_5394,N_4827,N_4851);
xor U5395 (N_5395,N_4753,N_4722);
nand U5396 (N_5396,N_4979,N_4951);
or U5397 (N_5397,N_4792,N_4933);
nand U5398 (N_5398,N_4979,N_4889);
xnor U5399 (N_5399,N_4751,N_4632);
nand U5400 (N_5400,N_4921,N_4559);
xnor U5401 (N_5401,N_4577,N_4619);
nand U5402 (N_5402,N_4960,N_4872);
nor U5403 (N_5403,N_4640,N_4585);
and U5404 (N_5404,N_4975,N_4608);
xor U5405 (N_5405,N_4742,N_4505);
and U5406 (N_5406,N_4572,N_4918);
nor U5407 (N_5407,N_4532,N_4524);
xnor U5408 (N_5408,N_4842,N_4666);
xor U5409 (N_5409,N_4723,N_4823);
nor U5410 (N_5410,N_4785,N_4581);
or U5411 (N_5411,N_4847,N_4673);
nand U5412 (N_5412,N_4872,N_4795);
and U5413 (N_5413,N_4876,N_4838);
nand U5414 (N_5414,N_4948,N_4673);
xor U5415 (N_5415,N_4500,N_4567);
xnor U5416 (N_5416,N_4620,N_4621);
nor U5417 (N_5417,N_4746,N_4790);
or U5418 (N_5418,N_4569,N_4889);
xor U5419 (N_5419,N_4553,N_4604);
nand U5420 (N_5420,N_4574,N_4604);
xor U5421 (N_5421,N_4686,N_4515);
xor U5422 (N_5422,N_4835,N_4966);
xnor U5423 (N_5423,N_4591,N_4616);
nand U5424 (N_5424,N_4832,N_4995);
nand U5425 (N_5425,N_4747,N_4547);
nor U5426 (N_5426,N_4969,N_4970);
nand U5427 (N_5427,N_4908,N_4971);
nor U5428 (N_5428,N_4550,N_4542);
xor U5429 (N_5429,N_4727,N_4723);
xnor U5430 (N_5430,N_4755,N_4874);
and U5431 (N_5431,N_4701,N_4673);
nor U5432 (N_5432,N_4948,N_4506);
or U5433 (N_5433,N_4662,N_4726);
nor U5434 (N_5434,N_4973,N_4871);
nand U5435 (N_5435,N_4761,N_4876);
or U5436 (N_5436,N_4548,N_4838);
or U5437 (N_5437,N_4765,N_4526);
or U5438 (N_5438,N_4694,N_4804);
nand U5439 (N_5439,N_4671,N_4640);
and U5440 (N_5440,N_4671,N_4699);
xor U5441 (N_5441,N_4988,N_4855);
and U5442 (N_5442,N_4839,N_4524);
nand U5443 (N_5443,N_4505,N_4667);
or U5444 (N_5444,N_4600,N_4905);
nand U5445 (N_5445,N_4793,N_4547);
and U5446 (N_5446,N_4922,N_4733);
nand U5447 (N_5447,N_4777,N_4564);
nor U5448 (N_5448,N_4800,N_4972);
nand U5449 (N_5449,N_4746,N_4617);
xnor U5450 (N_5450,N_4568,N_4866);
and U5451 (N_5451,N_4626,N_4984);
xor U5452 (N_5452,N_4760,N_4512);
nand U5453 (N_5453,N_4886,N_4890);
and U5454 (N_5454,N_4854,N_4718);
or U5455 (N_5455,N_4703,N_4911);
nor U5456 (N_5456,N_4778,N_4846);
or U5457 (N_5457,N_4974,N_4536);
nor U5458 (N_5458,N_4556,N_4964);
and U5459 (N_5459,N_4959,N_4970);
nand U5460 (N_5460,N_4688,N_4644);
xnor U5461 (N_5461,N_4947,N_4943);
nor U5462 (N_5462,N_4674,N_4730);
xnor U5463 (N_5463,N_4541,N_4706);
and U5464 (N_5464,N_4793,N_4799);
nor U5465 (N_5465,N_4684,N_4584);
or U5466 (N_5466,N_4840,N_4926);
nand U5467 (N_5467,N_4919,N_4952);
xnor U5468 (N_5468,N_4933,N_4612);
and U5469 (N_5469,N_4758,N_4908);
xnor U5470 (N_5470,N_4549,N_4978);
or U5471 (N_5471,N_4810,N_4709);
and U5472 (N_5472,N_4516,N_4837);
nand U5473 (N_5473,N_4824,N_4530);
and U5474 (N_5474,N_4587,N_4948);
nor U5475 (N_5475,N_4547,N_4995);
nor U5476 (N_5476,N_4963,N_4886);
nand U5477 (N_5477,N_4629,N_4636);
or U5478 (N_5478,N_4846,N_4915);
nand U5479 (N_5479,N_4532,N_4619);
or U5480 (N_5480,N_4959,N_4966);
nand U5481 (N_5481,N_4793,N_4721);
xnor U5482 (N_5482,N_4614,N_4934);
or U5483 (N_5483,N_4565,N_4788);
and U5484 (N_5484,N_4799,N_4970);
nor U5485 (N_5485,N_4839,N_4918);
nor U5486 (N_5486,N_4615,N_4744);
and U5487 (N_5487,N_4638,N_4984);
and U5488 (N_5488,N_4732,N_4682);
nand U5489 (N_5489,N_4733,N_4765);
nor U5490 (N_5490,N_4733,N_4564);
and U5491 (N_5491,N_4527,N_4932);
xor U5492 (N_5492,N_4819,N_4936);
and U5493 (N_5493,N_4822,N_4721);
and U5494 (N_5494,N_4848,N_4727);
or U5495 (N_5495,N_4803,N_4661);
or U5496 (N_5496,N_4941,N_4862);
and U5497 (N_5497,N_4592,N_4544);
xor U5498 (N_5498,N_4624,N_4798);
nor U5499 (N_5499,N_4724,N_4994);
or U5500 (N_5500,N_5055,N_5074);
nor U5501 (N_5501,N_5144,N_5091);
or U5502 (N_5502,N_5194,N_5051);
xnor U5503 (N_5503,N_5056,N_5233);
xor U5504 (N_5504,N_5421,N_5426);
or U5505 (N_5505,N_5489,N_5449);
xnor U5506 (N_5506,N_5198,N_5414);
and U5507 (N_5507,N_5161,N_5188);
nand U5508 (N_5508,N_5431,N_5040);
xnor U5509 (N_5509,N_5248,N_5106);
or U5510 (N_5510,N_5471,N_5433);
and U5511 (N_5511,N_5183,N_5011);
or U5512 (N_5512,N_5270,N_5023);
nor U5513 (N_5513,N_5484,N_5424);
nor U5514 (N_5514,N_5235,N_5175);
or U5515 (N_5515,N_5015,N_5010);
nor U5516 (N_5516,N_5383,N_5117);
nand U5517 (N_5517,N_5336,N_5070);
xor U5518 (N_5518,N_5276,N_5076);
xnor U5519 (N_5519,N_5408,N_5264);
or U5520 (N_5520,N_5192,N_5310);
xor U5521 (N_5521,N_5151,N_5013);
nor U5522 (N_5522,N_5080,N_5267);
nor U5523 (N_5523,N_5031,N_5227);
nand U5524 (N_5524,N_5283,N_5485);
and U5525 (N_5525,N_5320,N_5045);
and U5526 (N_5526,N_5016,N_5126);
or U5527 (N_5527,N_5348,N_5444);
nand U5528 (N_5528,N_5001,N_5277);
and U5529 (N_5529,N_5492,N_5361);
xor U5530 (N_5530,N_5138,N_5116);
xor U5531 (N_5531,N_5105,N_5285);
nand U5532 (N_5532,N_5354,N_5075);
and U5533 (N_5533,N_5462,N_5493);
and U5534 (N_5534,N_5178,N_5236);
nor U5535 (N_5535,N_5366,N_5041);
nor U5536 (N_5536,N_5316,N_5048);
nand U5537 (N_5537,N_5347,N_5002);
xor U5538 (N_5538,N_5231,N_5109);
or U5539 (N_5539,N_5226,N_5305);
nand U5540 (N_5540,N_5423,N_5456);
nand U5541 (N_5541,N_5306,N_5465);
xor U5542 (N_5542,N_5382,N_5396);
and U5543 (N_5543,N_5266,N_5262);
nand U5544 (N_5544,N_5490,N_5079);
and U5545 (N_5545,N_5049,N_5165);
nand U5546 (N_5546,N_5077,N_5129);
xor U5547 (N_5547,N_5084,N_5344);
or U5548 (N_5548,N_5272,N_5085);
or U5549 (N_5549,N_5249,N_5498);
or U5550 (N_5550,N_5038,N_5281);
or U5551 (N_5551,N_5030,N_5054);
xnor U5552 (N_5552,N_5438,N_5258);
xor U5553 (N_5553,N_5179,N_5416);
nand U5554 (N_5554,N_5278,N_5368);
xnor U5555 (N_5555,N_5323,N_5430);
nand U5556 (N_5556,N_5228,N_5429);
nand U5557 (N_5557,N_5389,N_5250);
nor U5558 (N_5558,N_5241,N_5229);
nand U5559 (N_5559,N_5434,N_5384);
xor U5560 (N_5560,N_5393,N_5359);
and U5561 (N_5561,N_5378,N_5474);
nor U5562 (N_5562,N_5140,N_5318);
nor U5563 (N_5563,N_5113,N_5173);
nand U5564 (N_5564,N_5162,N_5202);
nor U5565 (N_5565,N_5349,N_5370);
or U5566 (N_5566,N_5166,N_5042);
nor U5567 (N_5567,N_5339,N_5033);
xnor U5568 (N_5568,N_5428,N_5328);
nor U5569 (N_5569,N_5148,N_5478);
nand U5570 (N_5570,N_5333,N_5146);
xnor U5571 (N_5571,N_5253,N_5448);
nand U5572 (N_5572,N_5286,N_5170);
nor U5573 (N_5573,N_5189,N_5362);
nand U5574 (N_5574,N_5331,N_5123);
xnor U5575 (N_5575,N_5122,N_5037);
xor U5576 (N_5576,N_5487,N_5163);
nand U5577 (N_5577,N_5211,N_5247);
nand U5578 (N_5578,N_5068,N_5413);
nor U5579 (N_5579,N_5254,N_5441);
xor U5580 (N_5580,N_5006,N_5093);
and U5581 (N_5581,N_5386,N_5172);
nand U5582 (N_5582,N_5089,N_5311);
nor U5583 (N_5583,N_5353,N_5000);
and U5584 (N_5584,N_5225,N_5324);
nand U5585 (N_5585,N_5398,N_5210);
nand U5586 (N_5586,N_5299,N_5381);
and U5587 (N_5587,N_5181,N_5304);
and U5588 (N_5588,N_5083,N_5418);
nor U5589 (N_5589,N_5152,N_5346);
nor U5590 (N_5590,N_5268,N_5209);
or U5591 (N_5591,N_5097,N_5313);
nor U5592 (N_5592,N_5150,N_5303);
nand U5593 (N_5593,N_5447,N_5193);
xnor U5594 (N_5594,N_5375,N_5103);
nand U5595 (N_5595,N_5222,N_5427);
or U5596 (N_5596,N_5307,N_5059);
nor U5597 (N_5597,N_5100,N_5364);
xor U5598 (N_5598,N_5288,N_5240);
or U5599 (N_5599,N_5452,N_5115);
nor U5600 (N_5600,N_5176,N_5203);
nor U5601 (N_5601,N_5201,N_5153);
or U5602 (N_5602,N_5439,N_5317);
nor U5603 (N_5603,N_5101,N_5403);
or U5604 (N_5604,N_5341,N_5459);
xnor U5605 (N_5605,N_5132,N_5380);
nand U5606 (N_5606,N_5340,N_5125);
and U5607 (N_5607,N_5371,N_5357);
and U5608 (N_5608,N_5294,N_5481);
xnor U5609 (N_5609,N_5350,N_5321);
nor U5610 (N_5610,N_5453,N_5415);
or U5611 (N_5611,N_5302,N_5450);
xor U5612 (N_5612,N_5252,N_5464);
xnor U5613 (N_5613,N_5468,N_5399);
nor U5614 (N_5614,N_5355,N_5190);
nor U5615 (N_5615,N_5219,N_5182);
nand U5616 (N_5616,N_5088,N_5213);
and U5617 (N_5617,N_5218,N_5168);
or U5618 (N_5618,N_5147,N_5477);
and U5619 (N_5619,N_5437,N_5275);
or U5620 (N_5620,N_5470,N_5377);
and U5621 (N_5621,N_5026,N_5058);
nor U5622 (N_5622,N_5238,N_5110);
nand U5623 (N_5623,N_5047,N_5345);
nor U5624 (N_5624,N_5257,N_5032);
or U5625 (N_5625,N_5186,N_5496);
or U5626 (N_5626,N_5269,N_5039);
and U5627 (N_5627,N_5358,N_5284);
xor U5628 (N_5628,N_5099,N_5149);
nor U5629 (N_5629,N_5400,N_5034);
nor U5630 (N_5630,N_5312,N_5356);
and U5631 (N_5631,N_5325,N_5142);
and U5632 (N_5632,N_5021,N_5208);
and U5633 (N_5633,N_5488,N_5187);
and U5634 (N_5634,N_5363,N_5245);
xnor U5635 (N_5635,N_5206,N_5003);
nor U5636 (N_5636,N_5061,N_5141);
xnor U5637 (N_5637,N_5197,N_5046);
and U5638 (N_5638,N_5273,N_5029);
nand U5639 (N_5639,N_5184,N_5315);
xnor U5640 (N_5640,N_5133,N_5025);
and U5641 (N_5641,N_5171,N_5145);
xnor U5642 (N_5642,N_5155,N_5096);
nor U5643 (N_5643,N_5078,N_5329);
nand U5644 (N_5644,N_5024,N_5274);
xnor U5645 (N_5645,N_5330,N_5118);
nand U5646 (N_5646,N_5215,N_5425);
nor U5647 (N_5647,N_5296,N_5053);
and U5648 (N_5648,N_5018,N_5308);
and U5649 (N_5649,N_5369,N_5407);
nor U5650 (N_5650,N_5212,N_5230);
nor U5651 (N_5651,N_5458,N_5028);
xor U5652 (N_5652,N_5052,N_5290);
xor U5653 (N_5653,N_5164,N_5107);
nor U5654 (N_5654,N_5137,N_5195);
nand U5655 (N_5655,N_5461,N_5090);
and U5656 (N_5656,N_5397,N_5300);
nand U5657 (N_5657,N_5191,N_5160);
xor U5658 (N_5658,N_5388,N_5221);
xnor U5659 (N_5659,N_5136,N_5483);
or U5660 (N_5660,N_5005,N_5027);
nand U5661 (N_5661,N_5014,N_5261);
nand U5662 (N_5662,N_5334,N_5092);
nor U5663 (N_5663,N_5204,N_5255);
or U5664 (N_5664,N_5094,N_5174);
xor U5665 (N_5665,N_5319,N_5224);
xnor U5666 (N_5666,N_5259,N_5177);
or U5667 (N_5667,N_5409,N_5495);
nor U5668 (N_5668,N_5385,N_5360);
nand U5669 (N_5669,N_5337,N_5063);
and U5670 (N_5670,N_5108,N_5419);
xor U5671 (N_5671,N_5469,N_5480);
and U5672 (N_5672,N_5019,N_5012);
nand U5673 (N_5673,N_5373,N_5376);
xnor U5674 (N_5674,N_5223,N_5067);
nand U5675 (N_5675,N_5292,N_5072);
nor U5676 (N_5676,N_5217,N_5020);
xor U5677 (N_5677,N_5124,N_5243);
nand U5678 (N_5678,N_5422,N_5232);
or U5679 (N_5679,N_5128,N_5069);
xnor U5680 (N_5680,N_5499,N_5234);
or U5681 (N_5681,N_5466,N_5494);
or U5682 (N_5682,N_5404,N_5401);
and U5683 (N_5683,N_5180,N_5446);
xor U5684 (N_5684,N_5265,N_5295);
and U5685 (N_5685,N_5279,N_5017);
or U5686 (N_5686,N_5159,N_5411);
nand U5687 (N_5687,N_5064,N_5081);
or U5688 (N_5688,N_5256,N_5332);
or U5689 (N_5689,N_5237,N_5342);
nand U5690 (N_5690,N_5395,N_5417);
nor U5691 (N_5691,N_5475,N_5473);
nand U5692 (N_5692,N_5086,N_5087);
and U5693 (N_5693,N_5293,N_5390);
xor U5694 (N_5694,N_5050,N_5406);
and U5695 (N_5695,N_5322,N_5073);
nand U5696 (N_5696,N_5135,N_5467);
or U5697 (N_5697,N_5007,N_5239);
nor U5698 (N_5698,N_5440,N_5082);
nand U5699 (N_5699,N_5130,N_5271);
xor U5700 (N_5700,N_5291,N_5289);
xnor U5701 (N_5701,N_5491,N_5102);
nor U5702 (N_5702,N_5120,N_5062);
nand U5703 (N_5703,N_5112,N_5482);
and U5704 (N_5704,N_5309,N_5199);
nand U5705 (N_5705,N_5216,N_5095);
xor U5706 (N_5706,N_5451,N_5119);
nand U5707 (N_5707,N_5287,N_5314);
or U5708 (N_5708,N_5391,N_5443);
nor U5709 (N_5709,N_5022,N_5139);
or U5710 (N_5710,N_5326,N_5200);
xor U5711 (N_5711,N_5435,N_5167);
nor U5712 (N_5712,N_5134,N_5098);
and U5713 (N_5713,N_5121,N_5442);
xnor U5714 (N_5714,N_5214,N_5169);
nor U5715 (N_5715,N_5457,N_5158);
nand U5716 (N_5716,N_5060,N_5402);
nor U5717 (N_5717,N_5104,N_5035);
nand U5718 (N_5718,N_5154,N_5405);
or U5719 (N_5719,N_5043,N_5352);
nand U5720 (N_5720,N_5242,N_5066);
nor U5721 (N_5721,N_5367,N_5486);
nand U5722 (N_5722,N_5479,N_5036);
or U5723 (N_5723,N_5420,N_5301);
xor U5724 (N_5724,N_5205,N_5460);
and U5725 (N_5725,N_5327,N_5143);
or U5726 (N_5726,N_5131,N_5185);
xnor U5727 (N_5727,N_5338,N_5057);
nor U5728 (N_5728,N_5387,N_5298);
xnor U5729 (N_5729,N_5263,N_5282);
nand U5730 (N_5730,N_5412,N_5220);
nand U5731 (N_5731,N_5351,N_5476);
xnor U5732 (N_5732,N_5207,N_5374);
and U5733 (N_5733,N_5009,N_5157);
nand U5734 (N_5734,N_5280,N_5071);
and U5735 (N_5735,N_5432,N_5365);
or U5736 (N_5736,N_5251,N_5472);
nand U5737 (N_5737,N_5410,N_5196);
nand U5738 (N_5738,N_5044,N_5392);
nor U5739 (N_5739,N_5244,N_5114);
nor U5740 (N_5740,N_5065,N_5111);
and U5741 (N_5741,N_5463,N_5127);
and U5742 (N_5742,N_5455,N_5004);
or U5743 (N_5743,N_5156,N_5497);
or U5744 (N_5744,N_5436,N_5335);
or U5745 (N_5745,N_5297,N_5379);
xor U5746 (N_5746,N_5445,N_5372);
xnor U5747 (N_5747,N_5394,N_5008);
xor U5748 (N_5748,N_5260,N_5343);
and U5749 (N_5749,N_5246,N_5454);
or U5750 (N_5750,N_5201,N_5316);
nand U5751 (N_5751,N_5324,N_5311);
nand U5752 (N_5752,N_5140,N_5172);
xnor U5753 (N_5753,N_5482,N_5236);
nand U5754 (N_5754,N_5290,N_5493);
and U5755 (N_5755,N_5143,N_5084);
nor U5756 (N_5756,N_5216,N_5134);
xnor U5757 (N_5757,N_5249,N_5028);
nand U5758 (N_5758,N_5126,N_5358);
nor U5759 (N_5759,N_5181,N_5427);
or U5760 (N_5760,N_5224,N_5046);
nor U5761 (N_5761,N_5466,N_5145);
nor U5762 (N_5762,N_5355,N_5082);
or U5763 (N_5763,N_5487,N_5457);
nor U5764 (N_5764,N_5167,N_5077);
xor U5765 (N_5765,N_5069,N_5429);
or U5766 (N_5766,N_5327,N_5039);
xnor U5767 (N_5767,N_5157,N_5418);
or U5768 (N_5768,N_5444,N_5371);
xor U5769 (N_5769,N_5240,N_5334);
nand U5770 (N_5770,N_5008,N_5437);
nor U5771 (N_5771,N_5064,N_5321);
and U5772 (N_5772,N_5295,N_5469);
xnor U5773 (N_5773,N_5438,N_5376);
or U5774 (N_5774,N_5416,N_5189);
nand U5775 (N_5775,N_5421,N_5084);
or U5776 (N_5776,N_5295,N_5115);
or U5777 (N_5777,N_5443,N_5143);
nor U5778 (N_5778,N_5005,N_5372);
and U5779 (N_5779,N_5404,N_5120);
and U5780 (N_5780,N_5129,N_5243);
and U5781 (N_5781,N_5031,N_5470);
and U5782 (N_5782,N_5163,N_5129);
nand U5783 (N_5783,N_5407,N_5445);
nand U5784 (N_5784,N_5417,N_5131);
xnor U5785 (N_5785,N_5491,N_5277);
nand U5786 (N_5786,N_5037,N_5227);
and U5787 (N_5787,N_5008,N_5270);
nor U5788 (N_5788,N_5050,N_5188);
and U5789 (N_5789,N_5498,N_5264);
nand U5790 (N_5790,N_5122,N_5326);
nor U5791 (N_5791,N_5445,N_5282);
nor U5792 (N_5792,N_5245,N_5491);
xor U5793 (N_5793,N_5156,N_5313);
or U5794 (N_5794,N_5195,N_5304);
or U5795 (N_5795,N_5358,N_5231);
and U5796 (N_5796,N_5291,N_5097);
nor U5797 (N_5797,N_5428,N_5185);
or U5798 (N_5798,N_5269,N_5232);
nand U5799 (N_5799,N_5409,N_5312);
or U5800 (N_5800,N_5156,N_5422);
or U5801 (N_5801,N_5405,N_5267);
nor U5802 (N_5802,N_5057,N_5329);
or U5803 (N_5803,N_5027,N_5224);
nand U5804 (N_5804,N_5173,N_5213);
nor U5805 (N_5805,N_5186,N_5007);
nor U5806 (N_5806,N_5115,N_5098);
xor U5807 (N_5807,N_5312,N_5463);
nor U5808 (N_5808,N_5204,N_5449);
or U5809 (N_5809,N_5400,N_5372);
nand U5810 (N_5810,N_5472,N_5232);
and U5811 (N_5811,N_5281,N_5042);
nor U5812 (N_5812,N_5325,N_5241);
nand U5813 (N_5813,N_5104,N_5033);
nor U5814 (N_5814,N_5474,N_5278);
nand U5815 (N_5815,N_5392,N_5452);
nand U5816 (N_5816,N_5082,N_5199);
nor U5817 (N_5817,N_5273,N_5456);
and U5818 (N_5818,N_5171,N_5364);
or U5819 (N_5819,N_5363,N_5304);
xnor U5820 (N_5820,N_5344,N_5267);
xor U5821 (N_5821,N_5383,N_5002);
or U5822 (N_5822,N_5032,N_5049);
nor U5823 (N_5823,N_5318,N_5252);
nand U5824 (N_5824,N_5261,N_5338);
or U5825 (N_5825,N_5061,N_5131);
nand U5826 (N_5826,N_5046,N_5460);
xnor U5827 (N_5827,N_5088,N_5425);
nor U5828 (N_5828,N_5312,N_5109);
or U5829 (N_5829,N_5249,N_5155);
nand U5830 (N_5830,N_5155,N_5390);
or U5831 (N_5831,N_5306,N_5100);
xnor U5832 (N_5832,N_5003,N_5189);
nand U5833 (N_5833,N_5451,N_5092);
xor U5834 (N_5834,N_5144,N_5205);
nor U5835 (N_5835,N_5244,N_5493);
nand U5836 (N_5836,N_5201,N_5183);
nor U5837 (N_5837,N_5291,N_5416);
xnor U5838 (N_5838,N_5460,N_5424);
xor U5839 (N_5839,N_5289,N_5316);
nor U5840 (N_5840,N_5032,N_5489);
or U5841 (N_5841,N_5259,N_5266);
or U5842 (N_5842,N_5290,N_5489);
xor U5843 (N_5843,N_5316,N_5278);
or U5844 (N_5844,N_5043,N_5084);
nor U5845 (N_5845,N_5134,N_5132);
nor U5846 (N_5846,N_5228,N_5261);
or U5847 (N_5847,N_5378,N_5389);
nor U5848 (N_5848,N_5019,N_5240);
nand U5849 (N_5849,N_5277,N_5187);
and U5850 (N_5850,N_5366,N_5280);
xnor U5851 (N_5851,N_5036,N_5174);
nand U5852 (N_5852,N_5293,N_5110);
nor U5853 (N_5853,N_5190,N_5421);
and U5854 (N_5854,N_5076,N_5181);
or U5855 (N_5855,N_5328,N_5020);
and U5856 (N_5856,N_5268,N_5437);
nor U5857 (N_5857,N_5061,N_5377);
or U5858 (N_5858,N_5439,N_5321);
xor U5859 (N_5859,N_5314,N_5422);
or U5860 (N_5860,N_5131,N_5178);
xnor U5861 (N_5861,N_5170,N_5356);
nor U5862 (N_5862,N_5326,N_5195);
nor U5863 (N_5863,N_5394,N_5037);
or U5864 (N_5864,N_5156,N_5110);
nor U5865 (N_5865,N_5167,N_5371);
nor U5866 (N_5866,N_5252,N_5168);
nor U5867 (N_5867,N_5132,N_5302);
nand U5868 (N_5868,N_5244,N_5451);
nor U5869 (N_5869,N_5018,N_5251);
nor U5870 (N_5870,N_5315,N_5107);
nor U5871 (N_5871,N_5488,N_5349);
and U5872 (N_5872,N_5205,N_5268);
nor U5873 (N_5873,N_5411,N_5221);
or U5874 (N_5874,N_5383,N_5031);
or U5875 (N_5875,N_5430,N_5169);
nand U5876 (N_5876,N_5364,N_5224);
xnor U5877 (N_5877,N_5266,N_5149);
xnor U5878 (N_5878,N_5444,N_5164);
nor U5879 (N_5879,N_5007,N_5317);
nand U5880 (N_5880,N_5011,N_5072);
nand U5881 (N_5881,N_5354,N_5299);
nand U5882 (N_5882,N_5150,N_5475);
nor U5883 (N_5883,N_5192,N_5431);
or U5884 (N_5884,N_5008,N_5390);
and U5885 (N_5885,N_5194,N_5311);
nor U5886 (N_5886,N_5087,N_5471);
xnor U5887 (N_5887,N_5107,N_5329);
nand U5888 (N_5888,N_5063,N_5296);
nand U5889 (N_5889,N_5172,N_5119);
xor U5890 (N_5890,N_5141,N_5292);
or U5891 (N_5891,N_5114,N_5313);
and U5892 (N_5892,N_5312,N_5457);
and U5893 (N_5893,N_5139,N_5006);
xnor U5894 (N_5894,N_5474,N_5360);
xor U5895 (N_5895,N_5284,N_5215);
xor U5896 (N_5896,N_5371,N_5008);
and U5897 (N_5897,N_5263,N_5487);
nand U5898 (N_5898,N_5009,N_5220);
or U5899 (N_5899,N_5355,N_5147);
nor U5900 (N_5900,N_5486,N_5066);
nor U5901 (N_5901,N_5486,N_5495);
nand U5902 (N_5902,N_5350,N_5220);
nand U5903 (N_5903,N_5089,N_5366);
xnor U5904 (N_5904,N_5321,N_5409);
or U5905 (N_5905,N_5181,N_5338);
nand U5906 (N_5906,N_5120,N_5224);
nor U5907 (N_5907,N_5445,N_5035);
nor U5908 (N_5908,N_5010,N_5191);
and U5909 (N_5909,N_5451,N_5114);
nor U5910 (N_5910,N_5475,N_5068);
xnor U5911 (N_5911,N_5432,N_5051);
or U5912 (N_5912,N_5079,N_5351);
and U5913 (N_5913,N_5241,N_5201);
xor U5914 (N_5914,N_5002,N_5016);
nand U5915 (N_5915,N_5340,N_5332);
nand U5916 (N_5916,N_5499,N_5109);
and U5917 (N_5917,N_5463,N_5332);
or U5918 (N_5918,N_5028,N_5048);
or U5919 (N_5919,N_5335,N_5149);
nand U5920 (N_5920,N_5042,N_5306);
nand U5921 (N_5921,N_5324,N_5198);
nand U5922 (N_5922,N_5047,N_5260);
xnor U5923 (N_5923,N_5035,N_5298);
xnor U5924 (N_5924,N_5415,N_5089);
nor U5925 (N_5925,N_5499,N_5140);
nor U5926 (N_5926,N_5096,N_5332);
xor U5927 (N_5927,N_5037,N_5138);
nand U5928 (N_5928,N_5285,N_5352);
xnor U5929 (N_5929,N_5237,N_5223);
xnor U5930 (N_5930,N_5327,N_5384);
xor U5931 (N_5931,N_5269,N_5305);
nand U5932 (N_5932,N_5269,N_5249);
nand U5933 (N_5933,N_5017,N_5473);
or U5934 (N_5934,N_5057,N_5050);
xnor U5935 (N_5935,N_5107,N_5308);
nor U5936 (N_5936,N_5010,N_5360);
xnor U5937 (N_5937,N_5294,N_5250);
nand U5938 (N_5938,N_5053,N_5218);
xor U5939 (N_5939,N_5023,N_5353);
nand U5940 (N_5940,N_5473,N_5366);
and U5941 (N_5941,N_5413,N_5484);
nand U5942 (N_5942,N_5137,N_5014);
or U5943 (N_5943,N_5346,N_5430);
and U5944 (N_5944,N_5486,N_5373);
or U5945 (N_5945,N_5402,N_5098);
nand U5946 (N_5946,N_5009,N_5113);
xor U5947 (N_5947,N_5189,N_5223);
or U5948 (N_5948,N_5331,N_5294);
or U5949 (N_5949,N_5142,N_5056);
nor U5950 (N_5950,N_5337,N_5096);
xnor U5951 (N_5951,N_5238,N_5098);
or U5952 (N_5952,N_5282,N_5391);
xnor U5953 (N_5953,N_5082,N_5015);
nand U5954 (N_5954,N_5291,N_5022);
nor U5955 (N_5955,N_5255,N_5212);
and U5956 (N_5956,N_5318,N_5254);
nor U5957 (N_5957,N_5204,N_5132);
xnor U5958 (N_5958,N_5445,N_5274);
xor U5959 (N_5959,N_5396,N_5016);
or U5960 (N_5960,N_5096,N_5072);
xnor U5961 (N_5961,N_5433,N_5395);
nand U5962 (N_5962,N_5418,N_5276);
nor U5963 (N_5963,N_5427,N_5157);
or U5964 (N_5964,N_5247,N_5106);
or U5965 (N_5965,N_5297,N_5316);
xor U5966 (N_5966,N_5467,N_5397);
nand U5967 (N_5967,N_5176,N_5035);
nor U5968 (N_5968,N_5327,N_5044);
nor U5969 (N_5969,N_5114,N_5398);
and U5970 (N_5970,N_5417,N_5036);
xor U5971 (N_5971,N_5367,N_5251);
and U5972 (N_5972,N_5351,N_5245);
xnor U5973 (N_5973,N_5248,N_5351);
and U5974 (N_5974,N_5163,N_5085);
nand U5975 (N_5975,N_5431,N_5463);
nor U5976 (N_5976,N_5049,N_5133);
nand U5977 (N_5977,N_5304,N_5353);
and U5978 (N_5978,N_5110,N_5353);
nand U5979 (N_5979,N_5229,N_5414);
nand U5980 (N_5980,N_5115,N_5469);
or U5981 (N_5981,N_5416,N_5135);
xnor U5982 (N_5982,N_5046,N_5492);
nor U5983 (N_5983,N_5252,N_5222);
xnor U5984 (N_5984,N_5291,N_5253);
xnor U5985 (N_5985,N_5354,N_5076);
nand U5986 (N_5986,N_5218,N_5365);
xor U5987 (N_5987,N_5214,N_5241);
and U5988 (N_5988,N_5040,N_5098);
nor U5989 (N_5989,N_5292,N_5353);
nor U5990 (N_5990,N_5278,N_5246);
nand U5991 (N_5991,N_5008,N_5237);
xor U5992 (N_5992,N_5199,N_5266);
or U5993 (N_5993,N_5340,N_5345);
nand U5994 (N_5994,N_5471,N_5292);
xnor U5995 (N_5995,N_5392,N_5071);
or U5996 (N_5996,N_5261,N_5040);
nor U5997 (N_5997,N_5273,N_5376);
nand U5998 (N_5998,N_5085,N_5244);
nor U5999 (N_5999,N_5088,N_5420);
xor U6000 (N_6000,N_5850,N_5639);
and U6001 (N_6001,N_5827,N_5592);
or U6002 (N_6002,N_5959,N_5787);
nand U6003 (N_6003,N_5544,N_5699);
nand U6004 (N_6004,N_5947,N_5507);
nor U6005 (N_6005,N_5951,N_5804);
xnor U6006 (N_6006,N_5504,N_5894);
xnor U6007 (N_6007,N_5984,N_5574);
nand U6008 (N_6008,N_5734,N_5861);
nand U6009 (N_6009,N_5884,N_5832);
nand U6010 (N_6010,N_5610,N_5879);
nand U6011 (N_6011,N_5669,N_5591);
and U6012 (N_6012,N_5649,N_5874);
nand U6013 (N_6013,N_5571,N_5617);
and U6014 (N_6014,N_5908,N_5904);
or U6015 (N_6015,N_5612,N_5725);
nor U6016 (N_6016,N_5722,N_5663);
and U6017 (N_6017,N_5922,N_5944);
xor U6018 (N_6018,N_5829,N_5748);
or U6019 (N_6019,N_5731,N_5958);
or U6020 (N_6020,N_5541,N_5596);
and U6021 (N_6021,N_5935,N_5856);
and U6022 (N_6022,N_5750,N_5940);
or U6023 (N_6023,N_5522,N_5964);
nor U6024 (N_6024,N_5939,N_5893);
nand U6025 (N_6025,N_5989,N_5517);
nor U6026 (N_6026,N_5578,N_5733);
or U6027 (N_6027,N_5720,N_5611);
and U6028 (N_6028,N_5500,N_5636);
nor U6029 (N_6029,N_5868,N_5713);
nor U6030 (N_6030,N_5744,N_5718);
or U6031 (N_6031,N_5691,N_5943);
xor U6032 (N_6032,N_5569,N_5672);
xnor U6033 (N_6033,N_5647,N_5878);
and U6034 (N_6034,N_5509,N_5533);
xor U6035 (N_6035,N_5564,N_5668);
xor U6036 (N_6036,N_5621,N_5890);
or U6037 (N_6037,N_5687,N_5988);
xnor U6038 (N_6038,N_5705,N_5983);
nor U6039 (N_6039,N_5948,N_5973);
or U6040 (N_6040,N_5747,N_5682);
nand U6041 (N_6041,N_5588,N_5993);
nand U6042 (N_6042,N_5764,N_5797);
or U6043 (N_6043,N_5825,N_5506);
xnor U6044 (N_6044,N_5971,N_5917);
and U6045 (N_6045,N_5809,N_5537);
or U6046 (N_6046,N_5659,N_5585);
or U6047 (N_6047,N_5981,N_5801);
or U6048 (N_6048,N_5550,N_5587);
and U6049 (N_6049,N_5715,N_5763);
or U6050 (N_6050,N_5817,N_5549);
nor U6051 (N_6051,N_5936,N_5781);
and U6052 (N_6052,N_5824,N_5690);
nand U6053 (N_6053,N_5976,N_5812);
or U6054 (N_6054,N_5880,N_5969);
or U6055 (N_6055,N_5642,N_5651);
xor U6056 (N_6056,N_5540,N_5627);
and U6057 (N_6057,N_5816,N_5580);
nor U6058 (N_6058,N_5654,N_5698);
nand U6059 (N_6059,N_5711,N_5980);
xnor U6060 (N_6060,N_5521,N_5576);
and U6061 (N_6061,N_5778,N_5568);
and U6062 (N_6062,N_5901,N_5761);
nor U6063 (N_6063,N_5883,N_5814);
xor U6064 (N_6064,N_5967,N_5745);
nor U6065 (N_6065,N_5683,N_5789);
nor U6066 (N_6066,N_5534,N_5903);
nor U6067 (N_6067,N_5799,N_5674);
nand U6068 (N_6068,N_5990,N_5717);
nor U6069 (N_6069,N_5754,N_5561);
or U6070 (N_6070,N_5756,N_5932);
and U6071 (N_6071,N_5772,N_5759);
xnor U6072 (N_6072,N_5707,N_5567);
nand U6073 (N_6073,N_5842,N_5891);
or U6074 (N_6074,N_5701,N_5526);
xnor U6075 (N_6075,N_5595,N_5520);
and U6076 (N_6076,N_5834,N_5599);
or U6077 (N_6077,N_5539,N_5865);
nand U6078 (N_6078,N_5706,N_5782);
nand U6079 (N_6079,N_5860,N_5593);
nor U6080 (N_6080,N_5635,N_5511);
and U6081 (N_6081,N_5590,N_5552);
xnor U6082 (N_6082,N_5608,N_5977);
and U6083 (N_6083,N_5524,N_5972);
nand U6084 (N_6084,N_5907,N_5862);
and U6085 (N_6085,N_5873,N_5529);
or U6086 (N_6086,N_5937,N_5985);
or U6087 (N_6087,N_5996,N_5695);
nor U6088 (N_6088,N_5543,N_5645);
or U6089 (N_6089,N_5565,N_5700);
or U6090 (N_6090,N_5791,N_5783);
nand U6091 (N_6091,N_5805,N_5963);
nand U6092 (N_6092,N_5557,N_5650);
and U6093 (N_6093,N_5968,N_5726);
and U6094 (N_6094,N_5955,N_5995);
xor U6095 (N_6095,N_5910,N_5729);
nor U6096 (N_6096,N_5548,N_5965);
and U6097 (N_6097,N_5508,N_5531);
xnor U6098 (N_6098,N_5808,N_5954);
nor U6099 (N_6099,N_5577,N_5501);
nand U6100 (N_6100,N_5830,N_5502);
nand U6101 (N_6101,N_5685,N_5952);
xnor U6102 (N_6102,N_5620,N_5589);
xor U6103 (N_6103,N_5758,N_5515);
nand U6104 (N_6104,N_5542,N_5623);
nor U6105 (N_6105,N_5709,N_5871);
and U6106 (N_6106,N_5898,N_5696);
and U6107 (N_6107,N_5933,N_5606);
or U6108 (N_6108,N_5582,N_5742);
nand U6109 (N_6109,N_5949,N_5819);
and U6110 (N_6110,N_5689,N_5870);
nand U6111 (N_6111,N_5982,N_5902);
or U6112 (N_6112,N_5770,N_5974);
and U6113 (N_6113,N_5840,N_5633);
xnor U6114 (N_6114,N_5785,N_5628);
xnor U6115 (N_6115,N_5660,N_5924);
nor U6116 (N_6116,N_5609,N_5930);
or U6117 (N_6117,N_5762,N_5641);
or U6118 (N_6118,N_5530,N_5553);
or U6119 (N_6119,N_5743,N_5766);
and U6120 (N_6120,N_5941,N_5777);
and U6121 (N_6121,N_5913,N_5931);
and U6122 (N_6122,N_5950,N_5652);
nor U6123 (N_6123,N_5875,N_5869);
nor U6124 (N_6124,N_5723,N_5822);
nor U6125 (N_6125,N_5516,N_5684);
and U6126 (N_6126,N_5677,N_5887);
nand U6127 (N_6127,N_5831,N_5638);
nand U6128 (N_6128,N_5960,N_5518);
xor U6129 (N_6129,N_5992,N_5844);
nor U6130 (N_6130,N_5602,N_5845);
xor U6131 (N_6131,N_5876,N_5979);
xnor U6132 (N_6132,N_5795,N_5556);
nand U6133 (N_6133,N_5843,N_5688);
and U6134 (N_6134,N_5790,N_5545);
and U6135 (N_6135,N_5818,N_5661);
nor U6136 (N_6136,N_5572,N_5538);
xnor U6137 (N_6137,N_5528,N_5821);
xnor U6138 (N_6138,N_5676,N_5667);
xor U6139 (N_6139,N_5704,N_5839);
nor U6140 (N_6140,N_5841,N_5735);
xnor U6141 (N_6141,N_5694,N_5736);
nand U6142 (N_6142,N_5788,N_5523);
or U6143 (N_6143,N_5853,N_5820);
xnor U6144 (N_6144,N_5888,N_5916);
nor U6145 (N_6145,N_5811,N_5712);
or U6146 (N_6146,N_5721,N_5503);
nand U6147 (N_6147,N_5987,N_5673);
xor U6148 (N_6148,N_5746,N_5566);
and U6149 (N_6149,N_5961,N_5899);
or U6150 (N_6150,N_5732,N_5519);
or U6151 (N_6151,N_5915,N_5847);
nand U6152 (N_6152,N_5803,N_5665);
and U6153 (N_6153,N_5598,N_5863);
or U6154 (N_6154,N_5532,N_5896);
nand U6155 (N_6155,N_5838,N_5881);
nor U6156 (N_6156,N_5769,N_5823);
nor U6157 (N_6157,N_5505,N_5584);
and U6158 (N_6158,N_5885,N_5826);
or U6159 (N_6159,N_5757,N_5653);
or U6160 (N_6160,N_5909,N_5921);
or U6161 (N_6161,N_5798,N_5536);
or U6162 (N_6162,N_5905,N_5513);
nand U6163 (N_6163,N_5586,N_5562);
or U6164 (N_6164,N_5807,N_5767);
xnor U6165 (N_6165,N_5784,N_5854);
nand U6166 (N_6166,N_5877,N_5618);
nand U6167 (N_6167,N_5702,N_5752);
or U6168 (N_6168,N_5708,N_5716);
nand U6169 (N_6169,N_5792,N_5664);
nand U6170 (N_6170,N_5622,N_5895);
or U6171 (N_6171,N_5925,N_5575);
xnor U6172 (N_6172,N_5670,N_5573);
and U6173 (N_6173,N_5928,N_5710);
nor U6174 (N_6174,N_5857,N_5558);
and U6175 (N_6175,N_5859,N_5919);
nand U6176 (N_6176,N_5741,N_5942);
or U6177 (N_6177,N_5662,N_5833);
xnor U6178 (N_6178,N_5666,N_5866);
xnor U6179 (N_6179,N_5998,N_5900);
nand U6180 (N_6180,N_5625,N_5999);
nor U6181 (N_6181,N_5938,N_5837);
or U6182 (N_6182,N_5771,N_5889);
nand U6183 (N_6183,N_5906,N_5728);
xnor U6184 (N_6184,N_5815,N_5793);
xor U6185 (N_6185,N_5886,N_5648);
nor U6186 (N_6186,N_5546,N_5923);
nor U6187 (N_6187,N_5946,N_5624);
nor U6188 (N_6188,N_5813,N_5510);
xor U6189 (N_6189,N_5864,N_5927);
xor U6190 (N_6190,N_5594,N_5634);
nand U6191 (N_6191,N_5929,N_5724);
or U6192 (N_6192,N_5920,N_5926);
and U6193 (N_6193,N_5957,N_5962);
nor U6194 (N_6194,N_5644,N_5714);
nand U6195 (N_6195,N_5774,N_5892);
xor U6196 (N_6196,N_5911,N_5626);
and U6197 (N_6197,N_5678,N_5600);
or U6198 (N_6198,N_5855,N_5934);
nand U6199 (N_6199,N_5914,N_5882);
and U6200 (N_6200,N_5760,N_5835);
or U6201 (N_6201,N_5681,N_5535);
and U6202 (N_6202,N_5802,N_5755);
nor U6203 (N_6203,N_5851,N_5806);
xnor U6204 (N_6204,N_5604,N_5867);
nand U6205 (N_6205,N_5719,N_5849);
xor U6206 (N_6206,N_5675,N_5780);
and U6207 (N_6207,N_5740,N_5945);
nor U6208 (N_6208,N_5570,N_5697);
nor U6209 (N_6209,N_5629,N_5679);
and U6210 (N_6210,N_5828,N_5703);
nand U6211 (N_6211,N_5994,N_5616);
and U6212 (N_6212,N_5991,N_5607);
or U6213 (N_6213,N_5753,N_5615);
xnor U6214 (N_6214,N_5800,N_5727);
nor U6215 (N_6215,N_5581,N_5794);
nor U6216 (N_6216,N_5912,N_5512);
xnor U6217 (N_6217,N_5601,N_5640);
xor U6218 (N_6218,N_5656,N_5978);
xor U6219 (N_6219,N_5514,N_5597);
or U6220 (N_6220,N_5751,N_5657);
xnor U6221 (N_6221,N_5605,N_5637);
nor U6222 (N_6222,N_5614,N_5872);
or U6223 (N_6223,N_5554,N_5779);
or U6224 (N_6224,N_5786,N_5773);
nor U6225 (N_6225,N_5560,N_5768);
or U6226 (N_6226,N_5559,N_5986);
and U6227 (N_6227,N_5613,N_5630);
nor U6228 (N_6228,N_5631,N_5632);
and U6229 (N_6229,N_5970,N_5555);
nand U6230 (N_6230,N_5776,N_5848);
and U6231 (N_6231,N_5646,N_5680);
and U6232 (N_6232,N_5643,N_5527);
xnor U6233 (N_6233,N_5765,N_5563);
nor U6234 (N_6234,N_5775,N_5749);
or U6235 (N_6235,N_5852,N_5836);
and U6236 (N_6236,N_5547,N_5693);
and U6237 (N_6237,N_5810,N_5738);
xnor U6238 (N_6238,N_5975,N_5655);
nand U6239 (N_6239,N_5692,N_5966);
xor U6240 (N_6240,N_5603,N_5583);
nor U6241 (N_6241,N_5525,N_5858);
or U6242 (N_6242,N_5897,N_5730);
xor U6243 (N_6243,N_5739,N_5796);
nand U6244 (N_6244,N_5551,N_5956);
or U6245 (N_6245,N_5997,N_5686);
xnor U6246 (N_6246,N_5918,N_5671);
and U6247 (N_6247,N_5658,N_5579);
nand U6248 (N_6248,N_5737,N_5846);
and U6249 (N_6249,N_5953,N_5619);
nand U6250 (N_6250,N_5770,N_5562);
xor U6251 (N_6251,N_5650,N_5627);
and U6252 (N_6252,N_5762,N_5883);
or U6253 (N_6253,N_5679,N_5577);
or U6254 (N_6254,N_5778,N_5684);
xnor U6255 (N_6255,N_5878,N_5869);
xor U6256 (N_6256,N_5750,N_5529);
and U6257 (N_6257,N_5536,N_5525);
nor U6258 (N_6258,N_5788,N_5679);
nand U6259 (N_6259,N_5743,N_5846);
xnor U6260 (N_6260,N_5664,N_5502);
nor U6261 (N_6261,N_5961,N_5682);
and U6262 (N_6262,N_5947,N_5798);
xnor U6263 (N_6263,N_5570,N_5556);
and U6264 (N_6264,N_5834,N_5884);
xor U6265 (N_6265,N_5728,N_5921);
or U6266 (N_6266,N_5994,N_5790);
nor U6267 (N_6267,N_5884,N_5623);
nand U6268 (N_6268,N_5849,N_5505);
nor U6269 (N_6269,N_5800,N_5677);
or U6270 (N_6270,N_5966,N_5784);
or U6271 (N_6271,N_5777,N_5975);
or U6272 (N_6272,N_5770,N_5943);
and U6273 (N_6273,N_5854,N_5848);
nand U6274 (N_6274,N_5603,N_5892);
and U6275 (N_6275,N_5620,N_5570);
xor U6276 (N_6276,N_5917,N_5625);
and U6277 (N_6277,N_5690,N_5708);
or U6278 (N_6278,N_5732,N_5644);
nor U6279 (N_6279,N_5727,N_5768);
or U6280 (N_6280,N_5909,N_5502);
nand U6281 (N_6281,N_5621,N_5998);
nor U6282 (N_6282,N_5994,N_5626);
nand U6283 (N_6283,N_5648,N_5851);
xor U6284 (N_6284,N_5881,N_5633);
or U6285 (N_6285,N_5946,N_5824);
and U6286 (N_6286,N_5685,N_5986);
or U6287 (N_6287,N_5538,N_5685);
and U6288 (N_6288,N_5668,N_5875);
or U6289 (N_6289,N_5721,N_5769);
and U6290 (N_6290,N_5935,N_5783);
nand U6291 (N_6291,N_5668,N_5634);
xor U6292 (N_6292,N_5699,N_5978);
nand U6293 (N_6293,N_5870,N_5807);
and U6294 (N_6294,N_5837,N_5694);
and U6295 (N_6295,N_5507,N_5547);
xnor U6296 (N_6296,N_5507,N_5962);
nor U6297 (N_6297,N_5737,N_5569);
or U6298 (N_6298,N_5992,N_5796);
xnor U6299 (N_6299,N_5696,N_5837);
nor U6300 (N_6300,N_5880,N_5550);
or U6301 (N_6301,N_5741,N_5534);
nand U6302 (N_6302,N_5737,N_5829);
nor U6303 (N_6303,N_5879,N_5676);
and U6304 (N_6304,N_5967,N_5609);
nand U6305 (N_6305,N_5634,N_5951);
nor U6306 (N_6306,N_5857,N_5691);
nor U6307 (N_6307,N_5648,N_5803);
nand U6308 (N_6308,N_5843,N_5743);
and U6309 (N_6309,N_5690,N_5933);
or U6310 (N_6310,N_5920,N_5682);
xnor U6311 (N_6311,N_5502,N_5776);
or U6312 (N_6312,N_5918,N_5921);
or U6313 (N_6313,N_5818,N_5524);
xnor U6314 (N_6314,N_5521,N_5681);
nand U6315 (N_6315,N_5724,N_5906);
xnor U6316 (N_6316,N_5743,N_5998);
nand U6317 (N_6317,N_5778,N_5618);
and U6318 (N_6318,N_5549,N_5508);
or U6319 (N_6319,N_5977,N_5759);
nand U6320 (N_6320,N_5620,N_5778);
and U6321 (N_6321,N_5968,N_5509);
and U6322 (N_6322,N_5798,N_5985);
nand U6323 (N_6323,N_5619,N_5838);
xor U6324 (N_6324,N_5689,N_5970);
nand U6325 (N_6325,N_5935,N_5967);
or U6326 (N_6326,N_5977,N_5903);
xor U6327 (N_6327,N_5655,N_5960);
xnor U6328 (N_6328,N_5863,N_5557);
xor U6329 (N_6329,N_5806,N_5839);
nand U6330 (N_6330,N_5834,N_5752);
nor U6331 (N_6331,N_5870,N_5894);
and U6332 (N_6332,N_5839,N_5567);
nor U6333 (N_6333,N_5740,N_5536);
nor U6334 (N_6334,N_5957,N_5810);
xor U6335 (N_6335,N_5788,N_5872);
or U6336 (N_6336,N_5830,N_5626);
nand U6337 (N_6337,N_5812,N_5840);
or U6338 (N_6338,N_5809,N_5691);
xor U6339 (N_6339,N_5907,N_5790);
nand U6340 (N_6340,N_5652,N_5655);
nand U6341 (N_6341,N_5871,N_5950);
or U6342 (N_6342,N_5868,N_5973);
and U6343 (N_6343,N_5908,N_5660);
xor U6344 (N_6344,N_5728,N_5749);
xor U6345 (N_6345,N_5991,N_5772);
xnor U6346 (N_6346,N_5666,N_5827);
nand U6347 (N_6347,N_5832,N_5661);
or U6348 (N_6348,N_5623,N_5782);
xnor U6349 (N_6349,N_5740,N_5733);
nor U6350 (N_6350,N_5684,N_5548);
nand U6351 (N_6351,N_5675,N_5600);
nor U6352 (N_6352,N_5733,N_5848);
nor U6353 (N_6353,N_5708,N_5551);
nor U6354 (N_6354,N_5883,N_5968);
nor U6355 (N_6355,N_5763,N_5922);
or U6356 (N_6356,N_5969,N_5604);
xnor U6357 (N_6357,N_5670,N_5599);
nor U6358 (N_6358,N_5519,N_5675);
nand U6359 (N_6359,N_5841,N_5818);
xnor U6360 (N_6360,N_5992,N_5766);
nor U6361 (N_6361,N_5752,N_5563);
xnor U6362 (N_6362,N_5993,N_5861);
nand U6363 (N_6363,N_5569,N_5812);
or U6364 (N_6364,N_5692,N_5893);
and U6365 (N_6365,N_5822,N_5761);
and U6366 (N_6366,N_5721,N_5919);
and U6367 (N_6367,N_5844,N_5717);
and U6368 (N_6368,N_5835,N_5629);
xnor U6369 (N_6369,N_5922,N_5655);
or U6370 (N_6370,N_5597,N_5558);
xor U6371 (N_6371,N_5621,N_5827);
xnor U6372 (N_6372,N_5522,N_5999);
and U6373 (N_6373,N_5844,N_5943);
nand U6374 (N_6374,N_5903,N_5649);
or U6375 (N_6375,N_5679,N_5797);
nand U6376 (N_6376,N_5854,N_5834);
nand U6377 (N_6377,N_5661,N_5532);
xor U6378 (N_6378,N_5517,N_5801);
and U6379 (N_6379,N_5524,N_5739);
nand U6380 (N_6380,N_5761,N_5680);
xor U6381 (N_6381,N_5648,N_5790);
xnor U6382 (N_6382,N_5643,N_5558);
xor U6383 (N_6383,N_5735,N_5625);
and U6384 (N_6384,N_5677,N_5955);
or U6385 (N_6385,N_5683,N_5711);
nor U6386 (N_6386,N_5660,N_5584);
or U6387 (N_6387,N_5675,N_5659);
or U6388 (N_6388,N_5585,N_5582);
and U6389 (N_6389,N_5627,N_5720);
xnor U6390 (N_6390,N_5672,N_5564);
xnor U6391 (N_6391,N_5786,N_5966);
and U6392 (N_6392,N_5618,N_5770);
xor U6393 (N_6393,N_5839,N_5727);
xor U6394 (N_6394,N_5762,N_5754);
xnor U6395 (N_6395,N_5853,N_5511);
xnor U6396 (N_6396,N_5526,N_5544);
nor U6397 (N_6397,N_5616,N_5979);
or U6398 (N_6398,N_5711,N_5599);
nand U6399 (N_6399,N_5966,N_5590);
nand U6400 (N_6400,N_5842,N_5942);
nor U6401 (N_6401,N_5742,N_5723);
nor U6402 (N_6402,N_5553,N_5801);
nand U6403 (N_6403,N_5564,N_5624);
nor U6404 (N_6404,N_5898,N_5508);
xnor U6405 (N_6405,N_5630,N_5566);
or U6406 (N_6406,N_5858,N_5885);
or U6407 (N_6407,N_5607,N_5984);
nor U6408 (N_6408,N_5919,N_5825);
and U6409 (N_6409,N_5743,N_5751);
nand U6410 (N_6410,N_5948,N_5992);
xnor U6411 (N_6411,N_5763,N_5797);
and U6412 (N_6412,N_5573,N_5874);
nand U6413 (N_6413,N_5538,N_5910);
xnor U6414 (N_6414,N_5955,N_5530);
nor U6415 (N_6415,N_5785,N_5599);
nand U6416 (N_6416,N_5841,N_5529);
and U6417 (N_6417,N_5996,N_5968);
xnor U6418 (N_6418,N_5775,N_5510);
nand U6419 (N_6419,N_5917,N_5718);
nor U6420 (N_6420,N_5876,N_5766);
nand U6421 (N_6421,N_5882,N_5604);
nand U6422 (N_6422,N_5571,N_5796);
nand U6423 (N_6423,N_5863,N_5780);
nor U6424 (N_6424,N_5933,N_5769);
nor U6425 (N_6425,N_5522,N_5666);
or U6426 (N_6426,N_5580,N_5704);
nor U6427 (N_6427,N_5743,N_5950);
nand U6428 (N_6428,N_5754,N_5694);
xnor U6429 (N_6429,N_5810,N_5813);
or U6430 (N_6430,N_5578,N_5972);
xnor U6431 (N_6431,N_5606,N_5694);
nor U6432 (N_6432,N_5733,N_5889);
nand U6433 (N_6433,N_5859,N_5914);
or U6434 (N_6434,N_5602,N_5803);
or U6435 (N_6435,N_5760,N_5944);
xnor U6436 (N_6436,N_5589,N_5571);
or U6437 (N_6437,N_5743,N_5918);
and U6438 (N_6438,N_5938,N_5895);
nand U6439 (N_6439,N_5890,N_5884);
or U6440 (N_6440,N_5599,N_5733);
nor U6441 (N_6441,N_5804,N_5772);
and U6442 (N_6442,N_5614,N_5652);
or U6443 (N_6443,N_5754,N_5861);
and U6444 (N_6444,N_5979,N_5973);
xnor U6445 (N_6445,N_5609,N_5811);
xnor U6446 (N_6446,N_5794,N_5729);
nor U6447 (N_6447,N_5973,N_5537);
xnor U6448 (N_6448,N_5523,N_5787);
xor U6449 (N_6449,N_5581,N_5547);
nor U6450 (N_6450,N_5915,N_5898);
or U6451 (N_6451,N_5726,N_5579);
xor U6452 (N_6452,N_5868,N_5675);
nand U6453 (N_6453,N_5725,N_5893);
xnor U6454 (N_6454,N_5621,N_5944);
or U6455 (N_6455,N_5746,N_5888);
and U6456 (N_6456,N_5893,N_5608);
nand U6457 (N_6457,N_5872,N_5932);
and U6458 (N_6458,N_5644,N_5592);
xnor U6459 (N_6459,N_5755,N_5918);
nor U6460 (N_6460,N_5540,N_5694);
nor U6461 (N_6461,N_5948,N_5909);
or U6462 (N_6462,N_5921,N_5739);
and U6463 (N_6463,N_5984,N_5962);
nor U6464 (N_6464,N_5579,N_5623);
xor U6465 (N_6465,N_5716,N_5916);
nand U6466 (N_6466,N_5960,N_5749);
nor U6467 (N_6467,N_5716,N_5680);
nand U6468 (N_6468,N_5727,N_5741);
or U6469 (N_6469,N_5943,N_5775);
and U6470 (N_6470,N_5828,N_5697);
xor U6471 (N_6471,N_5556,N_5750);
and U6472 (N_6472,N_5575,N_5540);
nor U6473 (N_6473,N_5863,N_5660);
nor U6474 (N_6474,N_5858,N_5920);
or U6475 (N_6475,N_5617,N_5858);
xor U6476 (N_6476,N_5836,N_5688);
nor U6477 (N_6477,N_5728,N_5934);
or U6478 (N_6478,N_5732,N_5810);
and U6479 (N_6479,N_5550,N_5599);
and U6480 (N_6480,N_5535,N_5962);
nand U6481 (N_6481,N_5678,N_5700);
nor U6482 (N_6482,N_5865,N_5673);
and U6483 (N_6483,N_5506,N_5723);
xnor U6484 (N_6484,N_5622,N_5923);
nand U6485 (N_6485,N_5882,N_5921);
nand U6486 (N_6486,N_5946,N_5577);
nand U6487 (N_6487,N_5918,N_5782);
nor U6488 (N_6488,N_5678,N_5653);
nor U6489 (N_6489,N_5697,N_5959);
or U6490 (N_6490,N_5589,N_5515);
xnor U6491 (N_6491,N_5557,N_5746);
and U6492 (N_6492,N_5663,N_5675);
nor U6493 (N_6493,N_5799,N_5856);
nor U6494 (N_6494,N_5784,N_5672);
nor U6495 (N_6495,N_5938,N_5781);
nand U6496 (N_6496,N_5785,N_5679);
nand U6497 (N_6497,N_5900,N_5911);
or U6498 (N_6498,N_5649,N_5652);
or U6499 (N_6499,N_5676,N_5553);
nand U6500 (N_6500,N_6075,N_6334);
or U6501 (N_6501,N_6320,N_6023);
nor U6502 (N_6502,N_6025,N_6410);
nand U6503 (N_6503,N_6148,N_6159);
nand U6504 (N_6504,N_6365,N_6049);
and U6505 (N_6505,N_6323,N_6019);
and U6506 (N_6506,N_6324,N_6057);
and U6507 (N_6507,N_6110,N_6138);
nand U6508 (N_6508,N_6402,N_6013);
nor U6509 (N_6509,N_6037,N_6146);
nor U6510 (N_6510,N_6234,N_6186);
and U6511 (N_6511,N_6317,N_6038);
nand U6512 (N_6512,N_6034,N_6300);
or U6513 (N_6513,N_6281,N_6102);
and U6514 (N_6514,N_6386,N_6253);
and U6515 (N_6515,N_6134,N_6087);
nor U6516 (N_6516,N_6380,N_6100);
nor U6517 (N_6517,N_6198,N_6329);
or U6518 (N_6518,N_6116,N_6047);
xor U6519 (N_6519,N_6214,N_6274);
or U6520 (N_6520,N_6178,N_6242);
nand U6521 (N_6521,N_6245,N_6330);
or U6522 (N_6522,N_6020,N_6003);
xnor U6523 (N_6523,N_6017,N_6346);
or U6524 (N_6524,N_6237,N_6293);
nor U6525 (N_6525,N_6239,N_6267);
nor U6526 (N_6526,N_6255,N_6392);
nand U6527 (N_6527,N_6130,N_6268);
or U6528 (N_6528,N_6090,N_6092);
and U6529 (N_6529,N_6283,N_6459);
nor U6530 (N_6530,N_6168,N_6128);
and U6531 (N_6531,N_6262,N_6304);
xnor U6532 (N_6532,N_6289,N_6141);
nor U6533 (N_6533,N_6097,N_6415);
or U6534 (N_6534,N_6144,N_6012);
and U6535 (N_6535,N_6095,N_6467);
nor U6536 (N_6536,N_6139,N_6411);
and U6537 (N_6537,N_6355,N_6246);
nor U6538 (N_6538,N_6041,N_6021);
nand U6539 (N_6539,N_6477,N_6424);
xnor U6540 (N_6540,N_6111,N_6084);
xnor U6541 (N_6541,N_6230,N_6481);
nand U6542 (N_6542,N_6256,N_6363);
nand U6543 (N_6543,N_6301,N_6290);
and U6544 (N_6544,N_6121,N_6350);
nor U6545 (N_6545,N_6269,N_6180);
nand U6546 (N_6546,N_6263,N_6188);
and U6547 (N_6547,N_6107,N_6094);
xor U6548 (N_6548,N_6124,N_6444);
or U6549 (N_6549,N_6399,N_6279);
nor U6550 (N_6550,N_6493,N_6018);
and U6551 (N_6551,N_6101,N_6002);
or U6552 (N_6552,N_6387,N_6270);
xnor U6553 (N_6553,N_6160,N_6089);
nand U6554 (N_6554,N_6378,N_6383);
or U6555 (N_6555,N_6154,N_6202);
and U6556 (N_6556,N_6035,N_6074);
and U6557 (N_6557,N_6462,N_6054);
xor U6558 (N_6558,N_6059,N_6026);
and U6559 (N_6559,N_6409,N_6352);
or U6560 (N_6560,N_6498,N_6241);
nor U6561 (N_6561,N_6321,N_6260);
or U6562 (N_6562,N_6105,N_6266);
or U6563 (N_6563,N_6446,N_6431);
or U6564 (N_6564,N_6413,N_6199);
and U6565 (N_6565,N_6428,N_6476);
or U6566 (N_6566,N_6337,N_6227);
nor U6567 (N_6567,N_6332,N_6435);
nand U6568 (N_6568,N_6236,N_6053);
and U6569 (N_6569,N_6073,N_6419);
and U6570 (N_6570,N_6479,N_6308);
nand U6571 (N_6571,N_6447,N_6361);
nor U6572 (N_6572,N_6457,N_6078);
nor U6573 (N_6573,N_6229,N_6081);
or U6574 (N_6574,N_6135,N_6485);
xor U6575 (N_6575,N_6287,N_6357);
and U6576 (N_6576,N_6055,N_6120);
nand U6577 (N_6577,N_6076,N_6150);
or U6578 (N_6578,N_6052,N_6328);
nand U6579 (N_6579,N_6096,N_6473);
nor U6580 (N_6580,N_6179,N_6125);
and U6581 (N_6581,N_6187,N_6488);
or U6582 (N_6582,N_6405,N_6182);
or U6583 (N_6583,N_6398,N_6296);
or U6584 (N_6584,N_6219,N_6295);
or U6585 (N_6585,N_6109,N_6458);
nand U6586 (N_6586,N_6379,N_6369);
or U6587 (N_6587,N_6496,N_6151);
xnor U6588 (N_6588,N_6343,N_6085);
or U6589 (N_6589,N_6408,N_6396);
nor U6590 (N_6590,N_6194,N_6181);
nand U6591 (N_6591,N_6440,N_6292);
xor U6592 (N_6592,N_6068,N_6011);
nor U6593 (N_6593,N_6086,N_6401);
nor U6594 (N_6594,N_6032,N_6454);
xor U6595 (N_6595,N_6338,N_6185);
xnor U6596 (N_6596,N_6136,N_6311);
nor U6597 (N_6597,N_6484,N_6172);
xnor U6598 (N_6598,N_6000,N_6327);
and U6599 (N_6599,N_6114,N_6316);
xor U6600 (N_6600,N_6165,N_6288);
nor U6601 (N_6601,N_6122,N_6231);
nor U6602 (N_6602,N_6249,N_6204);
and U6603 (N_6603,N_6232,N_6046);
nor U6604 (N_6604,N_6455,N_6252);
nand U6605 (N_6605,N_6433,N_6403);
nor U6606 (N_6606,N_6247,N_6036);
xor U6607 (N_6607,N_6235,N_6077);
nand U6608 (N_6608,N_6226,N_6258);
nor U6609 (N_6609,N_6039,N_6208);
nor U6610 (N_6610,N_6091,N_6307);
nand U6611 (N_6611,N_6390,N_6388);
xor U6612 (N_6612,N_6098,N_6248);
nor U6613 (N_6613,N_6257,N_6360);
nand U6614 (N_6614,N_6063,N_6129);
or U6615 (N_6615,N_6315,N_6184);
or U6616 (N_6616,N_6341,N_6471);
and U6617 (N_6617,N_6282,N_6452);
nand U6618 (N_6618,N_6067,N_6340);
nor U6619 (N_6619,N_6143,N_6448);
and U6620 (N_6620,N_6351,N_6066);
xor U6621 (N_6621,N_6407,N_6381);
and U6622 (N_6622,N_6491,N_6264);
nand U6623 (N_6623,N_6275,N_6142);
or U6624 (N_6624,N_6394,N_6395);
nor U6625 (N_6625,N_6309,N_6382);
nor U6626 (N_6626,N_6276,N_6492);
nor U6627 (N_6627,N_6193,N_6028);
nand U6628 (N_6628,N_6104,N_6016);
or U6629 (N_6629,N_6430,N_6303);
nor U6630 (N_6630,N_6359,N_6490);
nor U6631 (N_6631,N_6072,N_6201);
nor U6632 (N_6632,N_6277,N_6022);
and U6633 (N_6633,N_6031,N_6313);
or U6634 (N_6634,N_6156,N_6212);
and U6635 (N_6635,N_6374,N_6335);
xnor U6636 (N_6636,N_6007,N_6456);
xor U6637 (N_6637,N_6216,N_6206);
nand U6638 (N_6638,N_6213,N_6432);
nand U6639 (N_6639,N_6305,N_6064);
or U6640 (N_6640,N_6118,N_6483);
nand U6641 (N_6641,N_6099,N_6243);
nor U6642 (N_6642,N_6065,N_6450);
nor U6643 (N_6643,N_6207,N_6210);
nand U6644 (N_6644,N_6157,N_6298);
nor U6645 (N_6645,N_6469,N_6008);
xor U6646 (N_6646,N_6489,N_6342);
nand U6647 (N_6647,N_6058,N_6362);
and U6648 (N_6648,N_6487,N_6333);
nand U6649 (N_6649,N_6171,N_6190);
nor U6650 (N_6650,N_6325,N_6368);
or U6651 (N_6651,N_6238,N_6437);
xor U6652 (N_6652,N_6434,N_6117);
or U6653 (N_6653,N_6347,N_6113);
and U6654 (N_6654,N_6108,N_6438);
nand U6655 (N_6655,N_6261,N_6391);
or U6656 (N_6656,N_6149,N_6417);
nor U6657 (N_6657,N_6331,N_6163);
or U6658 (N_6658,N_6414,N_6429);
nor U6659 (N_6659,N_6056,N_6441);
nor U6660 (N_6660,N_6140,N_6285);
xnor U6661 (N_6661,N_6251,N_6051);
nand U6662 (N_6662,N_6166,N_6233);
and U6663 (N_6663,N_6494,N_6044);
nand U6664 (N_6664,N_6222,N_6162);
nor U6665 (N_6665,N_6197,N_6451);
nand U6666 (N_6666,N_6196,N_6299);
and U6667 (N_6667,N_6254,N_6426);
or U6668 (N_6668,N_6131,N_6286);
xor U6669 (N_6669,N_6468,N_6083);
and U6670 (N_6670,N_6291,N_6348);
nor U6671 (N_6671,N_6112,N_6319);
nor U6672 (N_6672,N_6412,N_6209);
or U6673 (N_6673,N_6497,N_6133);
or U6674 (N_6674,N_6137,N_6442);
and U6675 (N_6675,N_6228,N_6119);
xnor U6676 (N_6676,N_6082,N_6284);
nor U6677 (N_6677,N_6106,N_6445);
nor U6678 (N_6678,N_6192,N_6421);
nand U6679 (N_6679,N_6215,N_6371);
nor U6680 (N_6680,N_6322,N_6191);
and U6681 (N_6681,N_6372,N_6080);
xor U6682 (N_6682,N_6155,N_6294);
or U6683 (N_6683,N_6079,N_6048);
and U6684 (N_6684,N_6225,N_6427);
nand U6685 (N_6685,N_6326,N_6480);
nor U6686 (N_6686,N_6203,N_6306);
and U6687 (N_6687,N_6061,N_6014);
and U6688 (N_6688,N_6376,N_6093);
nor U6689 (N_6689,N_6377,N_6170);
and U6690 (N_6690,N_6029,N_6443);
and U6691 (N_6691,N_6393,N_6297);
and U6692 (N_6692,N_6069,N_6189);
nand U6693 (N_6693,N_6482,N_6474);
xor U6694 (N_6694,N_6418,N_6318);
nand U6695 (N_6695,N_6259,N_6265);
and U6696 (N_6696,N_6453,N_6070);
nor U6697 (N_6697,N_6218,N_6183);
xor U6698 (N_6698,N_6177,N_6273);
nand U6699 (N_6699,N_6406,N_6010);
nor U6700 (N_6700,N_6103,N_6499);
nand U6701 (N_6701,N_6280,N_6153);
nor U6702 (N_6702,N_6466,N_6123);
nor U6703 (N_6703,N_6486,N_6420);
nand U6704 (N_6704,N_6167,N_6158);
xnor U6705 (N_6705,N_6161,N_6354);
nand U6706 (N_6706,N_6176,N_6436);
nor U6707 (N_6707,N_6464,N_6416);
nand U6708 (N_6708,N_6404,N_6302);
nor U6709 (N_6709,N_6200,N_6224);
xor U6710 (N_6710,N_6221,N_6071);
or U6711 (N_6711,N_6004,N_6353);
xor U6712 (N_6712,N_6175,N_6005);
or U6713 (N_6713,N_6145,N_6358);
or U6714 (N_6714,N_6126,N_6024);
or U6715 (N_6715,N_6423,N_6195);
or U6716 (N_6716,N_6062,N_6240);
and U6717 (N_6717,N_6147,N_6475);
xnor U6718 (N_6718,N_6088,N_6278);
nor U6719 (N_6719,N_6336,N_6042);
nand U6720 (N_6720,N_6356,N_6132);
nor U6721 (N_6721,N_6060,N_6439);
xor U6722 (N_6722,N_6271,N_6465);
nor U6723 (N_6723,N_6152,N_6272);
or U6724 (N_6724,N_6470,N_6173);
and U6725 (N_6725,N_6223,N_6015);
and U6726 (N_6726,N_6389,N_6367);
nand U6727 (N_6727,N_6366,N_6030);
xor U6728 (N_6728,N_6478,N_6040);
or U6729 (N_6729,N_6463,N_6495);
and U6730 (N_6730,N_6460,N_6375);
nand U6731 (N_6731,N_6314,N_6205);
and U6732 (N_6732,N_6312,N_6449);
or U6733 (N_6733,N_6220,N_6244);
or U6734 (N_6734,N_6250,N_6349);
or U6735 (N_6735,N_6127,N_6400);
xnor U6736 (N_6736,N_6310,N_6164);
or U6737 (N_6737,N_6009,N_6425);
or U6738 (N_6738,N_6027,N_6422);
xor U6739 (N_6739,N_6345,N_6373);
xnor U6740 (N_6740,N_6174,N_6472);
or U6741 (N_6741,N_6115,N_6370);
xnor U6742 (N_6742,N_6006,N_6033);
and U6743 (N_6743,N_6397,N_6385);
or U6744 (N_6744,N_6217,N_6461);
xor U6745 (N_6745,N_6364,N_6050);
or U6746 (N_6746,N_6344,N_6339);
nor U6747 (N_6747,N_6211,N_6169);
nand U6748 (N_6748,N_6045,N_6384);
or U6749 (N_6749,N_6001,N_6043);
or U6750 (N_6750,N_6256,N_6221);
nand U6751 (N_6751,N_6134,N_6440);
or U6752 (N_6752,N_6453,N_6164);
xor U6753 (N_6753,N_6421,N_6405);
and U6754 (N_6754,N_6398,N_6487);
and U6755 (N_6755,N_6024,N_6337);
or U6756 (N_6756,N_6220,N_6490);
xor U6757 (N_6757,N_6409,N_6261);
nand U6758 (N_6758,N_6409,N_6375);
xnor U6759 (N_6759,N_6418,N_6227);
or U6760 (N_6760,N_6419,N_6266);
nand U6761 (N_6761,N_6340,N_6225);
or U6762 (N_6762,N_6087,N_6364);
or U6763 (N_6763,N_6472,N_6175);
nand U6764 (N_6764,N_6419,N_6175);
xor U6765 (N_6765,N_6495,N_6163);
and U6766 (N_6766,N_6274,N_6195);
or U6767 (N_6767,N_6275,N_6071);
nor U6768 (N_6768,N_6351,N_6147);
xnor U6769 (N_6769,N_6008,N_6483);
or U6770 (N_6770,N_6082,N_6048);
or U6771 (N_6771,N_6372,N_6467);
or U6772 (N_6772,N_6051,N_6078);
nand U6773 (N_6773,N_6243,N_6052);
or U6774 (N_6774,N_6283,N_6091);
nor U6775 (N_6775,N_6276,N_6287);
or U6776 (N_6776,N_6046,N_6280);
xnor U6777 (N_6777,N_6275,N_6045);
and U6778 (N_6778,N_6312,N_6254);
and U6779 (N_6779,N_6341,N_6081);
and U6780 (N_6780,N_6362,N_6475);
or U6781 (N_6781,N_6266,N_6333);
nor U6782 (N_6782,N_6419,N_6262);
or U6783 (N_6783,N_6275,N_6031);
xor U6784 (N_6784,N_6137,N_6146);
or U6785 (N_6785,N_6474,N_6376);
nand U6786 (N_6786,N_6469,N_6350);
nand U6787 (N_6787,N_6012,N_6463);
nand U6788 (N_6788,N_6227,N_6301);
xor U6789 (N_6789,N_6221,N_6135);
and U6790 (N_6790,N_6378,N_6231);
nand U6791 (N_6791,N_6473,N_6245);
nor U6792 (N_6792,N_6221,N_6038);
or U6793 (N_6793,N_6118,N_6141);
and U6794 (N_6794,N_6380,N_6335);
nand U6795 (N_6795,N_6086,N_6274);
nand U6796 (N_6796,N_6309,N_6159);
nand U6797 (N_6797,N_6283,N_6269);
or U6798 (N_6798,N_6368,N_6235);
nand U6799 (N_6799,N_6182,N_6491);
xor U6800 (N_6800,N_6342,N_6427);
xor U6801 (N_6801,N_6002,N_6490);
nand U6802 (N_6802,N_6136,N_6063);
xnor U6803 (N_6803,N_6240,N_6415);
and U6804 (N_6804,N_6433,N_6475);
nor U6805 (N_6805,N_6473,N_6272);
or U6806 (N_6806,N_6369,N_6302);
nand U6807 (N_6807,N_6433,N_6261);
or U6808 (N_6808,N_6316,N_6068);
or U6809 (N_6809,N_6354,N_6251);
xor U6810 (N_6810,N_6312,N_6137);
xor U6811 (N_6811,N_6134,N_6366);
nand U6812 (N_6812,N_6085,N_6336);
or U6813 (N_6813,N_6444,N_6197);
nand U6814 (N_6814,N_6426,N_6078);
nor U6815 (N_6815,N_6033,N_6476);
nor U6816 (N_6816,N_6143,N_6303);
xnor U6817 (N_6817,N_6171,N_6179);
nor U6818 (N_6818,N_6353,N_6455);
nand U6819 (N_6819,N_6288,N_6230);
or U6820 (N_6820,N_6244,N_6054);
nor U6821 (N_6821,N_6258,N_6311);
xor U6822 (N_6822,N_6030,N_6063);
nor U6823 (N_6823,N_6290,N_6231);
xnor U6824 (N_6824,N_6116,N_6262);
xnor U6825 (N_6825,N_6221,N_6183);
nor U6826 (N_6826,N_6429,N_6296);
nor U6827 (N_6827,N_6402,N_6168);
and U6828 (N_6828,N_6122,N_6053);
or U6829 (N_6829,N_6405,N_6456);
xor U6830 (N_6830,N_6094,N_6221);
or U6831 (N_6831,N_6136,N_6046);
and U6832 (N_6832,N_6065,N_6114);
xnor U6833 (N_6833,N_6473,N_6427);
and U6834 (N_6834,N_6358,N_6002);
and U6835 (N_6835,N_6040,N_6441);
nand U6836 (N_6836,N_6161,N_6139);
nor U6837 (N_6837,N_6213,N_6061);
xor U6838 (N_6838,N_6158,N_6182);
nor U6839 (N_6839,N_6154,N_6153);
nor U6840 (N_6840,N_6150,N_6115);
and U6841 (N_6841,N_6280,N_6056);
and U6842 (N_6842,N_6002,N_6169);
nor U6843 (N_6843,N_6497,N_6417);
and U6844 (N_6844,N_6034,N_6479);
and U6845 (N_6845,N_6032,N_6357);
nor U6846 (N_6846,N_6201,N_6191);
xor U6847 (N_6847,N_6087,N_6155);
nor U6848 (N_6848,N_6073,N_6026);
or U6849 (N_6849,N_6043,N_6276);
and U6850 (N_6850,N_6456,N_6286);
and U6851 (N_6851,N_6065,N_6448);
nor U6852 (N_6852,N_6218,N_6474);
and U6853 (N_6853,N_6396,N_6028);
or U6854 (N_6854,N_6027,N_6222);
xor U6855 (N_6855,N_6334,N_6357);
nor U6856 (N_6856,N_6392,N_6113);
and U6857 (N_6857,N_6094,N_6364);
and U6858 (N_6858,N_6299,N_6230);
or U6859 (N_6859,N_6189,N_6270);
or U6860 (N_6860,N_6418,N_6488);
nand U6861 (N_6861,N_6155,N_6467);
nor U6862 (N_6862,N_6490,N_6328);
and U6863 (N_6863,N_6374,N_6059);
and U6864 (N_6864,N_6403,N_6048);
nand U6865 (N_6865,N_6128,N_6177);
and U6866 (N_6866,N_6394,N_6427);
and U6867 (N_6867,N_6072,N_6309);
or U6868 (N_6868,N_6345,N_6485);
nor U6869 (N_6869,N_6448,N_6260);
nand U6870 (N_6870,N_6068,N_6024);
nor U6871 (N_6871,N_6459,N_6114);
and U6872 (N_6872,N_6136,N_6320);
xnor U6873 (N_6873,N_6154,N_6253);
xor U6874 (N_6874,N_6252,N_6243);
xnor U6875 (N_6875,N_6023,N_6460);
nor U6876 (N_6876,N_6152,N_6090);
or U6877 (N_6877,N_6079,N_6244);
and U6878 (N_6878,N_6056,N_6368);
nand U6879 (N_6879,N_6299,N_6273);
nand U6880 (N_6880,N_6360,N_6202);
nor U6881 (N_6881,N_6012,N_6374);
or U6882 (N_6882,N_6142,N_6083);
xnor U6883 (N_6883,N_6401,N_6468);
nand U6884 (N_6884,N_6198,N_6078);
nand U6885 (N_6885,N_6381,N_6099);
xnor U6886 (N_6886,N_6458,N_6041);
or U6887 (N_6887,N_6234,N_6068);
or U6888 (N_6888,N_6285,N_6329);
or U6889 (N_6889,N_6056,N_6453);
nand U6890 (N_6890,N_6049,N_6027);
and U6891 (N_6891,N_6285,N_6179);
xnor U6892 (N_6892,N_6442,N_6210);
and U6893 (N_6893,N_6002,N_6469);
xor U6894 (N_6894,N_6409,N_6017);
or U6895 (N_6895,N_6352,N_6432);
nor U6896 (N_6896,N_6000,N_6207);
and U6897 (N_6897,N_6057,N_6136);
and U6898 (N_6898,N_6013,N_6480);
nor U6899 (N_6899,N_6127,N_6013);
nand U6900 (N_6900,N_6129,N_6323);
and U6901 (N_6901,N_6353,N_6473);
or U6902 (N_6902,N_6322,N_6100);
nor U6903 (N_6903,N_6165,N_6324);
nor U6904 (N_6904,N_6310,N_6320);
nand U6905 (N_6905,N_6321,N_6188);
nor U6906 (N_6906,N_6405,N_6124);
nand U6907 (N_6907,N_6051,N_6267);
and U6908 (N_6908,N_6083,N_6146);
nor U6909 (N_6909,N_6217,N_6005);
nand U6910 (N_6910,N_6337,N_6177);
nand U6911 (N_6911,N_6097,N_6128);
and U6912 (N_6912,N_6408,N_6317);
xor U6913 (N_6913,N_6211,N_6010);
nand U6914 (N_6914,N_6158,N_6016);
nand U6915 (N_6915,N_6044,N_6485);
or U6916 (N_6916,N_6201,N_6044);
xnor U6917 (N_6917,N_6314,N_6256);
or U6918 (N_6918,N_6248,N_6383);
nand U6919 (N_6919,N_6058,N_6118);
nor U6920 (N_6920,N_6121,N_6282);
and U6921 (N_6921,N_6338,N_6102);
and U6922 (N_6922,N_6086,N_6110);
xor U6923 (N_6923,N_6108,N_6006);
and U6924 (N_6924,N_6463,N_6434);
nand U6925 (N_6925,N_6303,N_6272);
or U6926 (N_6926,N_6236,N_6452);
xor U6927 (N_6927,N_6327,N_6072);
nor U6928 (N_6928,N_6042,N_6221);
and U6929 (N_6929,N_6353,N_6304);
nor U6930 (N_6930,N_6438,N_6061);
and U6931 (N_6931,N_6223,N_6491);
xor U6932 (N_6932,N_6050,N_6491);
nand U6933 (N_6933,N_6277,N_6299);
and U6934 (N_6934,N_6301,N_6427);
and U6935 (N_6935,N_6487,N_6422);
or U6936 (N_6936,N_6205,N_6085);
or U6937 (N_6937,N_6074,N_6454);
and U6938 (N_6938,N_6153,N_6201);
and U6939 (N_6939,N_6225,N_6434);
xnor U6940 (N_6940,N_6195,N_6251);
nor U6941 (N_6941,N_6087,N_6182);
xnor U6942 (N_6942,N_6309,N_6476);
or U6943 (N_6943,N_6472,N_6364);
and U6944 (N_6944,N_6337,N_6396);
and U6945 (N_6945,N_6228,N_6250);
and U6946 (N_6946,N_6473,N_6230);
nor U6947 (N_6947,N_6056,N_6434);
xor U6948 (N_6948,N_6097,N_6051);
and U6949 (N_6949,N_6002,N_6015);
xnor U6950 (N_6950,N_6253,N_6461);
nand U6951 (N_6951,N_6347,N_6010);
and U6952 (N_6952,N_6205,N_6323);
nand U6953 (N_6953,N_6235,N_6000);
xor U6954 (N_6954,N_6208,N_6168);
xor U6955 (N_6955,N_6133,N_6457);
or U6956 (N_6956,N_6186,N_6327);
nand U6957 (N_6957,N_6078,N_6202);
xnor U6958 (N_6958,N_6397,N_6104);
and U6959 (N_6959,N_6143,N_6325);
xor U6960 (N_6960,N_6042,N_6444);
and U6961 (N_6961,N_6467,N_6054);
nor U6962 (N_6962,N_6486,N_6256);
and U6963 (N_6963,N_6162,N_6108);
xnor U6964 (N_6964,N_6128,N_6457);
or U6965 (N_6965,N_6404,N_6101);
or U6966 (N_6966,N_6247,N_6257);
or U6967 (N_6967,N_6181,N_6044);
xor U6968 (N_6968,N_6433,N_6305);
nand U6969 (N_6969,N_6039,N_6322);
xor U6970 (N_6970,N_6438,N_6115);
and U6971 (N_6971,N_6497,N_6486);
nand U6972 (N_6972,N_6218,N_6041);
and U6973 (N_6973,N_6267,N_6432);
or U6974 (N_6974,N_6347,N_6392);
xor U6975 (N_6975,N_6098,N_6009);
xnor U6976 (N_6976,N_6387,N_6346);
nand U6977 (N_6977,N_6315,N_6447);
or U6978 (N_6978,N_6415,N_6254);
nor U6979 (N_6979,N_6007,N_6258);
nand U6980 (N_6980,N_6389,N_6181);
nor U6981 (N_6981,N_6395,N_6063);
nor U6982 (N_6982,N_6444,N_6061);
or U6983 (N_6983,N_6021,N_6044);
nor U6984 (N_6984,N_6459,N_6105);
xor U6985 (N_6985,N_6067,N_6483);
nand U6986 (N_6986,N_6408,N_6363);
nor U6987 (N_6987,N_6088,N_6327);
nand U6988 (N_6988,N_6096,N_6252);
xor U6989 (N_6989,N_6031,N_6213);
or U6990 (N_6990,N_6176,N_6292);
nand U6991 (N_6991,N_6415,N_6185);
nand U6992 (N_6992,N_6333,N_6238);
nand U6993 (N_6993,N_6039,N_6210);
nor U6994 (N_6994,N_6260,N_6024);
xnor U6995 (N_6995,N_6304,N_6326);
nand U6996 (N_6996,N_6479,N_6117);
and U6997 (N_6997,N_6276,N_6243);
xnor U6998 (N_6998,N_6346,N_6301);
xor U6999 (N_6999,N_6235,N_6447);
xor U7000 (N_7000,N_6513,N_6820);
xnor U7001 (N_7001,N_6719,N_6612);
nand U7002 (N_7002,N_6787,N_6843);
xor U7003 (N_7003,N_6879,N_6611);
or U7004 (N_7004,N_6914,N_6949);
xor U7005 (N_7005,N_6774,N_6892);
nand U7006 (N_7006,N_6502,N_6673);
nand U7007 (N_7007,N_6662,N_6872);
nor U7008 (N_7008,N_6970,N_6882);
nand U7009 (N_7009,N_6973,N_6635);
nor U7010 (N_7010,N_6830,N_6508);
and U7011 (N_7011,N_6689,N_6595);
or U7012 (N_7012,N_6541,N_6964);
xor U7013 (N_7013,N_6526,N_6702);
or U7014 (N_7014,N_6760,N_6993);
nand U7015 (N_7015,N_6940,N_6838);
or U7016 (N_7016,N_6590,N_6659);
and U7017 (N_7017,N_6714,N_6919);
or U7018 (N_7018,N_6986,N_6530);
nand U7019 (N_7019,N_6568,N_6740);
xor U7020 (N_7020,N_6581,N_6965);
nand U7021 (N_7021,N_6672,N_6693);
and U7022 (N_7022,N_6766,N_6971);
xor U7023 (N_7023,N_6622,N_6755);
or U7024 (N_7024,N_6745,N_6792);
nor U7025 (N_7025,N_6731,N_6790);
nor U7026 (N_7026,N_6870,N_6738);
nand U7027 (N_7027,N_6916,N_6982);
nor U7028 (N_7028,N_6674,N_6527);
or U7029 (N_7029,N_6725,N_6899);
and U7030 (N_7030,N_6898,N_6942);
and U7031 (N_7031,N_6620,N_6761);
xor U7032 (N_7032,N_6763,N_6996);
nand U7033 (N_7033,N_6871,N_6796);
nor U7034 (N_7034,N_6715,N_6900);
and U7035 (N_7035,N_6684,N_6580);
and U7036 (N_7036,N_6555,N_6851);
and U7037 (N_7037,N_6592,N_6698);
and U7038 (N_7038,N_6607,N_6987);
nor U7039 (N_7039,N_6700,N_6545);
nand U7040 (N_7040,N_6500,N_6921);
nor U7041 (N_7041,N_6972,N_6748);
or U7042 (N_7042,N_6791,N_6969);
and U7043 (N_7043,N_6514,N_6544);
nor U7044 (N_7044,N_6877,N_6891);
nor U7045 (N_7045,N_6887,N_6976);
nor U7046 (N_7046,N_6565,N_6924);
nand U7047 (N_7047,N_6678,N_6805);
and U7048 (N_7048,N_6634,N_6742);
and U7049 (N_7049,N_6506,N_6998);
or U7050 (N_7050,N_6605,N_6951);
and U7051 (N_7051,N_6632,N_6923);
nand U7052 (N_7052,N_6886,N_6618);
nand U7053 (N_7053,N_6586,N_6551);
xor U7054 (N_7054,N_6546,N_6999);
or U7055 (N_7055,N_6572,N_6703);
nor U7056 (N_7056,N_6813,N_6517);
xnor U7057 (N_7057,N_6915,N_6571);
nand U7058 (N_7058,N_6859,N_6690);
nand U7059 (N_7059,N_6995,N_6627);
xor U7060 (N_7060,N_6944,N_6683);
nor U7061 (N_7061,N_6802,N_6840);
nand U7062 (N_7062,N_6962,N_6873);
and U7063 (N_7063,N_6656,N_6515);
nor U7064 (N_7064,N_6668,N_6988);
or U7065 (N_7065,N_6729,N_6904);
nor U7066 (N_7066,N_6633,N_6650);
or U7067 (N_7067,N_6855,N_6799);
or U7068 (N_7068,N_6960,N_6599);
nand U7069 (N_7069,N_6510,N_6936);
xnor U7070 (N_7070,N_6905,N_6516);
nand U7071 (N_7071,N_6903,N_6628);
or U7072 (N_7072,N_6528,N_6707);
xor U7073 (N_7073,N_6817,N_6560);
or U7074 (N_7074,N_6614,N_6952);
nor U7075 (N_7075,N_6676,N_6681);
and U7076 (N_7076,N_6959,N_6889);
and U7077 (N_7077,N_6688,N_6549);
nor U7078 (N_7078,N_6902,N_6857);
xnor U7079 (N_7079,N_6569,N_6721);
or U7080 (N_7080,N_6888,N_6630);
and U7081 (N_7081,N_6573,N_6542);
xor U7082 (N_7082,N_6806,N_6613);
nor U7083 (N_7083,N_6833,N_6687);
nand U7084 (N_7084,N_6600,N_6558);
xnor U7085 (N_7085,N_6928,N_6778);
nor U7086 (N_7086,N_6822,N_6686);
xor U7087 (N_7087,N_6780,N_6847);
nor U7088 (N_7088,N_6594,N_6744);
and U7089 (N_7089,N_6804,N_6538);
nor U7090 (N_7090,N_6846,N_6750);
nor U7091 (N_7091,N_6785,N_6974);
nand U7092 (N_7092,N_6699,N_6677);
and U7093 (N_7093,N_6570,N_6694);
xor U7094 (N_7094,N_6732,N_6543);
nand U7095 (N_7095,N_6669,N_6927);
nand U7096 (N_7096,N_6654,N_6926);
or U7097 (N_7097,N_6625,N_6598);
or U7098 (N_7098,N_6741,N_6578);
or U7099 (N_7099,N_6685,N_6657);
nor U7100 (N_7100,N_6810,N_6910);
nor U7101 (N_7101,N_6624,N_6647);
or U7102 (N_7102,N_6884,N_6705);
and U7103 (N_7103,N_6579,N_6680);
or U7104 (N_7104,N_6563,N_6756);
nand U7105 (N_7105,N_6653,N_6880);
or U7106 (N_7106,N_6733,N_6616);
nor U7107 (N_7107,N_6621,N_6757);
xor U7108 (N_7108,N_6772,N_6786);
or U7109 (N_7109,N_6861,N_6821);
nand U7110 (N_7110,N_6896,N_6701);
xor U7111 (N_7111,N_6961,N_6588);
nand U7112 (N_7112,N_6779,N_6597);
nand U7113 (N_7113,N_6713,N_6539);
nand U7114 (N_7114,N_6979,N_6907);
or U7115 (N_7115,N_6853,N_6519);
nand U7116 (N_7116,N_6845,N_6561);
xnor U7117 (N_7117,N_6909,N_6920);
and U7118 (N_7118,N_6946,N_6564);
or U7119 (N_7119,N_6764,N_6858);
nor U7120 (N_7120,N_6868,N_6795);
nand U7121 (N_7121,N_6617,N_6576);
nor U7122 (N_7122,N_6874,N_6990);
nand U7123 (N_7123,N_6797,N_6950);
nand U7124 (N_7124,N_6531,N_6644);
xor U7125 (N_7125,N_6582,N_6826);
nor U7126 (N_7126,N_6807,N_6692);
nand U7127 (N_7127,N_6878,N_6525);
or U7128 (N_7128,N_6665,N_6704);
xor U7129 (N_7129,N_6623,N_6587);
xor U7130 (N_7130,N_6913,N_6609);
nor U7131 (N_7131,N_6777,N_6606);
and U7132 (N_7132,N_6963,N_6636);
xnor U7133 (N_7133,N_6512,N_6574);
xnor U7134 (N_7134,N_6863,N_6717);
xor U7135 (N_7135,N_6844,N_6997);
or U7136 (N_7136,N_6893,N_6504);
and U7137 (N_7137,N_6610,N_6945);
xnor U7138 (N_7138,N_6752,N_6897);
or U7139 (N_7139,N_6697,N_6934);
and U7140 (N_7140,N_6724,N_6890);
xor U7141 (N_7141,N_6985,N_6929);
xnor U7142 (N_7142,N_6815,N_6941);
xor U7143 (N_7143,N_6743,N_6726);
or U7144 (N_7144,N_6661,N_6984);
xor U7145 (N_7145,N_6825,N_6955);
nor U7146 (N_7146,N_6768,N_6708);
nand U7147 (N_7147,N_6849,N_6521);
and U7148 (N_7148,N_6585,N_6666);
or U7149 (N_7149,N_6601,N_6832);
nor U7150 (N_7150,N_6770,N_6501);
and U7151 (N_7151,N_6781,N_6842);
nor U7152 (N_7152,N_6789,N_6735);
xor U7153 (N_7153,N_6591,N_6869);
or U7154 (N_7154,N_6948,N_6975);
xor U7155 (N_7155,N_6589,N_6819);
nand U7156 (N_7156,N_6619,N_6818);
nor U7157 (N_7157,N_6922,N_6667);
xnor U7158 (N_7158,N_6522,N_6981);
xor U7159 (N_7159,N_6556,N_6682);
and U7160 (N_7160,N_6524,N_6720);
nor U7161 (N_7161,N_6566,N_6584);
or U7162 (N_7162,N_6912,N_6631);
nor U7163 (N_7163,N_6583,N_6559);
nand U7164 (N_7164,N_6552,N_6860);
xnor U7165 (N_7165,N_6954,N_6968);
nor U7166 (N_7166,N_6529,N_6992);
nor U7167 (N_7167,N_6728,N_6824);
nor U7168 (N_7168,N_6794,N_6862);
or U7169 (N_7169,N_6876,N_6722);
nand U7170 (N_7170,N_6933,N_6577);
xnor U7171 (N_7171,N_6638,N_6856);
nor U7172 (N_7172,N_6557,N_6671);
or U7173 (N_7173,N_6894,N_6604);
xnor U7174 (N_7174,N_6727,N_6739);
and U7175 (N_7175,N_6901,N_6935);
xor U7176 (N_7176,N_6536,N_6937);
and U7177 (N_7177,N_6540,N_6753);
or U7178 (N_7178,N_6788,N_6643);
or U7179 (N_7179,N_6664,N_6850);
or U7180 (N_7180,N_6749,N_6637);
or U7181 (N_7181,N_6608,N_6931);
or U7182 (N_7182,N_6831,N_6652);
nand U7183 (N_7183,N_6696,N_6983);
xnor U7184 (N_7184,N_6706,N_6930);
nor U7185 (N_7185,N_6641,N_6509);
or U7186 (N_7186,N_6864,N_6837);
nor U7187 (N_7187,N_6759,N_6827);
xor U7188 (N_7188,N_6645,N_6505);
or U7189 (N_7189,N_6518,N_6814);
xor U7190 (N_7190,N_6523,N_6852);
nand U7191 (N_7191,N_6917,N_6783);
or U7192 (N_7192,N_6736,N_6782);
nor U7193 (N_7193,N_6553,N_6660);
nand U7194 (N_7194,N_6989,N_6670);
nor U7195 (N_7195,N_6865,N_6503);
nand U7196 (N_7196,N_6593,N_6642);
or U7197 (N_7197,N_6746,N_6829);
nor U7198 (N_7198,N_6567,N_6991);
nand U7199 (N_7199,N_6554,N_6562);
or U7200 (N_7200,N_6771,N_6550);
nor U7201 (N_7201,N_6776,N_6867);
nor U7202 (N_7202,N_6754,N_6906);
or U7203 (N_7203,N_6547,N_6751);
xnor U7204 (N_7204,N_6640,N_6953);
nand U7205 (N_7205,N_6798,N_6811);
and U7206 (N_7206,N_6812,N_6875);
xor U7207 (N_7207,N_6532,N_6691);
nand U7208 (N_7208,N_6658,N_6977);
or U7209 (N_7209,N_6793,N_6932);
or U7210 (N_7210,N_6994,N_6695);
nor U7211 (N_7211,N_6648,N_6758);
nor U7212 (N_7212,N_6535,N_6773);
nor U7213 (N_7213,N_6967,N_6957);
xor U7214 (N_7214,N_6679,N_6651);
nor U7215 (N_7215,N_6978,N_6767);
nor U7216 (N_7216,N_6784,N_6711);
nor U7217 (N_7217,N_6956,N_6841);
and U7218 (N_7218,N_6834,N_6762);
nand U7219 (N_7219,N_6747,N_6908);
nor U7220 (N_7220,N_6866,N_6675);
and U7221 (N_7221,N_6626,N_6801);
nor U7222 (N_7222,N_6943,N_6548);
xnor U7223 (N_7223,N_6663,N_6615);
and U7224 (N_7224,N_6734,N_6854);
and U7225 (N_7225,N_6712,N_6958);
nand U7226 (N_7226,N_6533,N_6839);
nand U7227 (N_7227,N_6716,N_6918);
nand U7228 (N_7228,N_6723,N_6808);
or U7229 (N_7229,N_6596,N_6718);
nor U7230 (N_7230,N_6649,N_6629);
or U7231 (N_7231,N_6534,N_6639);
nand U7232 (N_7232,N_6881,N_6730);
or U7233 (N_7233,N_6769,N_6511);
and U7234 (N_7234,N_6520,N_6537);
and U7235 (N_7235,N_6848,N_6947);
or U7236 (N_7236,N_6828,N_6646);
or U7237 (N_7237,N_6885,N_6765);
xor U7238 (N_7238,N_6911,N_6816);
xor U7239 (N_7239,N_6980,N_6823);
nand U7240 (N_7240,N_6883,N_6655);
and U7241 (N_7241,N_6803,N_6895);
xnor U7242 (N_7242,N_6775,N_6737);
xor U7243 (N_7243,N_6575,N_6603);
or U7244 (N_7244,N_6800,N_6925);
and U7245 (N_7245,N_6835,N_6710);
xor U7246 (N_7246,N_6709,N_6809);
nand U7247 (N_7247,N_6939,N_6966);
nor U7248 (N_7248,N_6602,N_6836);
xnor U7249 (N_7249,N_6507,N_6938);
nand U7250 (N_7250,N_6783,N_6736);
or U7251 (N_7251,N_6836,N_6812);
and U7252 (N_7252,N_6692,N_6645);
and U7253 (N_7253,N_6764,N_6873);
nand U7254 (N_7254,N_6599,N_6601);
or U7255 (N_7255,N_6679,N_6839);
nor U7256 (N_7256,N_6619,N_6712);
or U7257 (N_7257,N_6643,N_6747);
and U7258 (N_7258,N_6660,N_6893);
nor U7259 (N_7259,N_6789,N_6581);
and U7260 (N_7260,N_6538,N_6594);
nand U7261 (N_7261,N_6832,N_6776);
or U7262 (N_7262,N_6927,N_6828);
and U7263 (N_7263,N_6642,N_6635);
nor U7264 (N_7264,N_6564,N_6621);
and U7265 (N_7265,N_6884,N_6902);
and U7266 (N_7266,N_6965,N_6925);
and U7267 (N_7267,N_6984,N_6637);
nor U7268 (N_7268,N_6673,N_6996);
and U7269 (N_7269,N_6933,N_6516);
and U7270 (N_7270,N_6552,N_6974);
and U7271 (N_7271,N_6577,N_6834);
nand U7272 (N_7272,N_6931,N_6969);
and U7273 (N_7273,N_6711,N_6528);
or U7274 (N_7274,N_6587,N_6983);
and U7275 (N_7275,N_6527,N_6769);
and U7276 (N_7276,N_6863,N_6971);
nand U7277 (N_7277,N_6690,N_6540);
xor U7278 (N_7278,N_6925,N_6517);
or U7279 (N_7279,N_6743,N_6759);
nand U7280 (N_7280,N_6885,N_6985);
nor U7281 (N_7281,N_6793,N_6787);
and U7282 (N_7282,N_6772,N_6727);
and U7283 (N_7283,N_6599,N_6565);
nor U7284 (N_7284,N_6974,N_6766);
nor U7285 (N_7285,N_6564,N_6899);
xnor U7286 (N_7286,N_6903,N_6955);
nand U7287 (N_7287,N_6528,N_6739);
nor U7288 (N_7288,N_6953,N_6860);
xnor U7289 (N_7289,N_6778,N_6500);
nand U7290 (N_7290,N_6630,N_6692);
xnor U7291 (N_7291,N_6957,N_6698);
and U7292 (N_7292,N_6909,N_6972);
xor U7293 (N_7293,N_6829,N_6687);
nand U7294 (N_7294,N_6537,N_6803);
nor U7295 (N_7295,N_6762,N_6982);
xnor U7296 (N_7296,N_6557,N_6956);
nand U7297 (N_7297,N_6812,N_6621);
nor U7298 (N_7298,N_6738,N_6998);
nand U7299 (N_7299,N_6963,N_6597);
nor U7300 (N_7300,N_6716,N_6736);
nand U7301 (N_7301,N_6983,N_6876);
xor U7302 (N_7302,N_6992,N_6964);
or U7303 (N_7303,N_6865,N_6730);
and U7304 (N_7304,N_6872,N_6625);
and U7305 (N_7305,N_6740,N_6553);
and U7306 (N_7306,N_6693,N_6871);
xnor U7307 (N_7307,N_6948,N_6658);
or U7308 (N_7308,N_6919,N_6672);
xor U7309 (N_7309,N_6600,N_6752);
nand U7310 (N_7310,N_6893,N_6538);
or U7311 (N_7311,N_6794,N_6843);
or U7312 (N_7312,N_6691,N_6915);
or U7313 (N_7313,N_6703,N_6900);
xnor U7314 (N_7314,N_6852,N_6793);
nor U7315 (N_7315,N_6658,N_6553);
xor U7316 (N_7316,N_6717,N_6834);
or U7317 (N_7317,N_6704,N_6643);
nand U7318 (N_7318,N_6716,N_6919);
and U7319 (N_7319,N_6714,N_6911);
xor U7320 (N_7320,N_6654,N_6586);
nor U7321 (N_7321,N_6596,N_6890);
or U7322 (N_7322,N_6761,N_6771);
nor U7323 (N_7323,N_6607,N_6846);
nand U7324 (N_7324,N_6649,N_6811);
nor U7325 (N_7325,N_6918,N_6665);
or U7326 (N_7326,N_6759,N_6852);
nor U7327 (N_7327,N_6705,N_6640);
nand U7328 (N_7328,N_6951,N_6628);
nor U7329 (N_7329,N_6951,N_6697);
or U7330 (N_7330,N_6899,N_6829);
and U7331 (N_7331,N_6875,N_6729);
nor U7332 (N_7332,N_6515,N_6752);
or U7333 (N_7333,N_6743,N_6506);
xnor U7334 (N_7334,N_6549,N_6738);
nor U7335 (N_7335,N_6695,N_6720);
nor U7336 (N_7336,N_6572,N_6791);
and U7337 (N_7337,N_6667,N_6513);
and U7338 (N_7338,N_6547,N_6597);
xor U7339 (N_7339,N_6518,N_6812);
nor U7340 (N_7340,N_6870,N_6666);
and U7341 (N_7341,N_6696,N_6646);
and U7342 (N_7342,N_6831,N_6645);
and U7343 (N_7343,N_6500,N_6750);
nand U7344 (N_7344,N_6776,N_6904);
nor U7345 (N_7345,N_6768,N_6643);
and U7346 (N_7346,N_6898,N_6570);
or U7347 (N_7347,N_6613,N_6989);
or U7348 (N_7348,N_6708,N_6980);
and U7349 (N_7349,N_6620,N_6898);
xnor U7350 (N_7350,N_6545,N_6868);
nor U7351 (N_7351,N_6608,N_6930);
nand U7352 (N_7352,N_6681,N_6621);
xor U7353 (N_7353,N_6801,N_6871);
or U7354 (N_7354,N_6947,N_6863);
and U7355 (N_7355,N_6743,N_6546);
or U7356 (N_7356,N_6913,N_6560);
and U7357 (N_7357,N_6949,N_6811);
or U7358 (N_7358,N_6950,N_6968);
nor U7359 (N_7359,N_6710,N_6754);
nor U7360 (N_7360,N_6636,N_6984);
nor U7361 (N_7361,N_6721,N_6785);
xnor U7362 (N_7362,N_6929,N_6715);
nor U7363 (N_7363,N_6534,N_6945);
nor U7364 (N_7364,N_6592,N_6580);
xnor U7365 (N_7365,N_6913,N_6627);
nor U7366 (N_7366,N_6659,N_6796);
xnor U7367 (N_7367,N_6511,N_6593);
nand U7368 (N_7368,N_6877,N_6923);
or U7369 (N_7369,N_6817,N_6859);
xor U7370 (N_7370,N_6528,N_6596);
and U7371 (N_7371,N_6655,N_6998);
nand U7372 (N_7372,N_6997,N_6741);
nor U7373 (N_7373,N_6776,N_6579);
xor U7374 (N_7374,N_6975,N_6784);
nand U7375 (N_7375,N_6882,N_6702);
and U7376 (N_7376,N_6941,N_6501);
nand U7377 (N_7377,N_6753,N_6758);
xor U7378 (N_7378,N_6773,N_6981);
nor U7379 (N_7379,N_6602,N_6604);
and U7380 (N_7380,N_6871,N_6725);
nand U7381 (N_7381,N_6896,N_6931);
nor U7382 (N_7382,N_6758,N_6894);
nand U7383 (N_7383,N_6586,N_6946);
nand U7384 (N_7384,N_6745,N_6854);
nor U7385 (N_7385,N_6639,N_6624);
or U7386 (N_7386,N_6838,N_6714);
xor U7387 (N_7387,N_6602,N_6876);
nand U7388 (N_7388,N_6833,N_6726);
or U7389 (N_7389,N_6927,N_6978);
nor U7390 (N_7390,N_6975,N_6942);
nand U7391 (N_7391,N_6872,N_6692);
and U7392 (N_7392,N_6583,N_6808);
xor U7393 (N_7393,N_6512,N_6682);
nor U7394 (N_7394,N_6782,N_6901);
xor U7395 (N_7395,N_6761,N_6728);
and U7396 (N_7396,N_6595,N_6876);
or U7397 (N_7397,N_6570,N_6774);
xnor U7398 (N_7398,N_6983,N_6875);
and U7399 (N_7399,N_6858,N_6694);
nand U7400 (N_7400,N_6536,N_6523);
and U7401 (N_7401,N_6968,N_6669);
or U7402 (N_7402,N_6788,N_6769);
nor U7403 (N_7403,N_6857,N_6878);
or U7404 (N_7404,N_6961,N_6823);
nand U7405 (N_7405,N_6818,N_6947);
xnor U7406 (N_7406,N_6523,N_6799);
or U7407 (N_7407,N_6508,N_6735);
or U7408 (N_7408,N_6759,N_6697);
nor U7409 (N_7409,N_6565,N_6678);
nand U7410 (N_7410,N_6645,N_6512);
and U7411 (N_7411,N_6784,N_6587);
xnor U7412 (N_7412,N_6814,N_6516);
xnor U7413 (N_7413,N_6556,N_6767);
xnor U7414 (N_7414,N_6896,N_6679);
nor U7415 (N_7415,N_6544,N_6758);
nor U7416 (N_7416,N_6971,N_6788);
nand U7417 (N_7417,N_6910,N_6596);
nor U7418 (N_7418,N_6726,N_6916);
and U7419 (N_7419,N_6870,N_6900);
and U7420 (N_7420,N_6915,N_6679);
and U7421 (N_7421,N_6643,N_6703);
nand U7422 (N_7422,N_6502,N_6945);
or U7423 (N_7423,N_6593,N_6757);
nor U7424 (N_7424,N_6946,N_6682);
xnor U7425 (N_7425,N_6531,N_6879);
and U7426 (N_7426,N_6598,N_6943);
or U7427 (N_7427,N_6665,N_6700);
nor U7428 (N_7428,N_6625,N_6949);
nor U7429 (N_7429,N_6580,N_6890);
nand U7430 (N_7430,N_6543,N_6748);
xnor U7431 (N_7431,N_6799,N_6775);
or U7432 (N_7432,N_6561,N_6546);
nand U7433 (N_7433,N_6853,N_6515);
nor U7434 (N_7434,N_6823,N_6830);
nor U7435 (N_7435,N_6686,N_6606);
xor U7436 (N_7436,N_6538,N_6828);
nor U7437 (N_7437,N_6873,N_6907);
nor U7438 (N_7438,N_6565,N_6723);
and U7439 (N_7439,N_6631,N_6765);
nand U7440 (N_7440,N_6670,N_6774);
and U7441 (N_7441,N_6617,N_6667);
and U7442 (N_7442,N_6653,N_6588);
or U7443 (N_7443,N_6932,N_6539);
or U7444 (N_7444,N_6521,N_6899);
xor U7445 (N_7445,N_6931,N_6929);
xor U7446 (N_7446,N_6876,N_6899);
or U7447 (N_7447,N_6617,N_6915);
and U7448 (N_7448,N_6528,N_6791);
or U7449 (N_7449,N_6939,N_6974);
and U7450 (N_7450,N_6695,N_6778);
nor U7451 (N_7451,N_6747,N_6509);
and U7452 (N_7452,N_6517,N_6673);
and U7453 (N_7453,N_6662,N_6610);
and U7454 (N_7454,N_6918,N_6732);
and U7455 (N_7455,N_6533,N_6876);
or U7456 (N_7456,N_6895,N_6663);
xnor U7457 (N_7457,N_6753,N_6842);
or U7458 (N_7458,N_6669,N_6529);
nor U7459 (N_7459,N_6553,N_6543);
xor U7460 (N_7460,N_6851,N_6547);
xnor U7461 (N_7461,N_6857,N_6836);
nand U7462 (N_7462,N_6586,N_6645);
xnor U7463 (N_7463,N_6666,N_6861);
xor U7464 (N_7464,N_6505,N_6884);
and U7465 (N_7465,N_6507,N_6762);
and U7466 (N_7466,N_6604,N_6699);
xnor U7467 (N_7467,N_6500,N_6515);
and U7468 (N_7468,N_6821,N_6780);
and U7469 (N_7469,N_6537,N_6516);
xnor U7470 (N_7470,N_6546,N_6979);
and U7471 (N_7471,N_6977,N_6936);
nor U7472 (N_7472,N_6809,N_6972);
and U7473 (N_7473,N_6797,N_6862);
nand U7474 (N_7474,N_6623,N_6681);
nand U7475 (N_7475,N_6893,N_6790);
nand U7476 (N_7476,N_6826,N_6991);
nand U7477 (N_7477,N_6609,N_6900);
xor U7478 (N_7478,N_6942,N_6882);
or U7479 (N_7479,N_6520,N_6893);
nor U7480 (N_7480,N_6742,N_6733);
nor U7481 (N_7481,N_6904,N_6689);
and U7482 (N_7482,N_6507,N_6505);
and U7483 (N_7483,N_6750,N_6964);
nand U7484 (N_7484,N_6979,N_6924);
nor U7485 (N_7485,N_6697,N_6975);
and U7486 (N_7486,N_6650,N_6923);
nand U7487 (N_7487,N_6600,N_6795);
or U7488 (N_7488,N_6783,N_6954);
or U7489 (N_7489,N_6881,N_6617);
and U7490 (N_7490,N_6624,N_6599);
nor U7491 (N_7491,N_6575,N_6777);
xnor U7492 (N_7492,N_6534,N_6953);
nand U7493 (N_7493,N_6748,N_6772);
or U7494 (N_7494,N_6925,N_6904);
xor U7495 (N_7495,N_6749,N_6868);
nor U7496 (N_7496,N_6687,N_6794);
xnor U7497 (N_7497,N_6802,N_6937);
nor U7498 (N_7498,N_6844,N_6603);
and U7499 (N_7499,N_6657,N_6746);
nand U7500 (N_7500,N_7089,N_7469);
nor U7501 (N_7501,N_7360,N_7167);
nor U7502 (N_7502,N_7064,N_7411);
xor U7503 (N_7503,N_7148,N_7434);
nand U7504 (N_7504,N_7039,N_7102);
and U7505 (N_7505,N_7430,N_7462);
or U7506 (N_7506,N_7497,N_7441);
nor U7507 (N_7507,N_7380,N_7228);
nor U7508 (N_7508,N_7284,N_7223);
xor U7509 (N_7509,N_7108,N_7169);
nor U7510 (N_7510,N_7128,N_7371);
nor U7511 (N_7511,N_7447,N_7330);
or U7512 (N_7512,N_7409,N_7000);
nor U7513 (N_7513,N_7395,N_7298);
and U7514 (N_7514,N_7345,N_7154);
and U7515 (N_7515,N_7304,N_7106);
nand U7516 (N_7516,N_7214,N_7467);
or U7517 (N_7517,N_7481,N_7254);
and U7518 (N_7518,N_7276,N_7138);
nand U7519 (N_7519,N_7165,N_7094);
xnor U7520 (N_7520,N_7315,N_7428);
nand U7521 (N_7521,N_7087,N_7268);
nor U7522 (N_7522,N_7008,N_7237);
and U7523 (N_7523,N_7445,N_7029);
nand U7524 (N_7524,N_7376,N_7009);
xnor U7525 (N_7525,N_7056,N_7435);
nor U7526 (N_7526,N_7136,N_7016);
and U7527 (N_7527,N_7240,N_7294);
nand U7528 (N_7528,N_7369,N_7152);
and U7529 (N_7529,N_7377,N_7090);
xnor U7530 (N_7530,N_7220,N_7389);
or U7531 (N_7531,N_7006,N_7425);
and U7532 (N_7532,N_7110,N_7471);
or U7533 (N_7533,N_7137,N_7224);
or U7534 (N_7534,N_7019,N_7446);
and U7535 (N_7535,N_7143,N_7341);
nor U7536 (N_7536,N_7199,N_7200);
nand U7537 (N_7537,N_7300,N_7118);
nand U7538 (N_7538,N_7069,N_7005);
nor U7539 (N_7539,N_7272,N_7114);
and U7540 (N_7540,N_7092,N_7473);
or U7541 (N_7541,N_7034,N_7286);
nand U7542 (N_7542,N_7235,N_7242);
xnor U7543 (N_7543,N_7403,N_7212);
nor U7544 (N_7544,N_7363,N_7429);
nand U7545 (N_7545,N_7465,N_7076);
and U7546 (N_7546,N_7097,N_7335);
and U7547 (N_7547,N_7193,N_7252);
nor U7548 (N_7548,N_7227,N_7017);
xor U7549 (N_7549,N_7303,N_7078);
and U7550 (N_7550,N_7324,N_7147);
xor U7551 (N_7551,N_7067,N_7474);
or U7552 (N_7552,N_7221,N_7157);
nand U7553 (N_7553,N_7264,N_7073);
xor U7554 (N_7554,N_7156,N_7354);
or U7555 (N_7555,N_7129,N_7436);
nor U7556 (N_7556,N_7144,N_7450);
xnor U7557 (N_7557,N_7386,N_7260);
or U7558 (N_7558,N_7295,N_7424);
nand U7559 (N_7559,N_7011,N_7236);
or U7560 (N_7560,N_7291,N_7209);
and U7561 (N_7561,N_7247,N_7490);
xor U7562 (N_7562,N_7385,N_7026);
or U7563 (N_7563,N_7265,N_7329);
nand U7564 (N_7564,N_7099,N_7004);
nor U7565 (N_7565,N_7479,N_7478);
and U7566 (N_7566,N_7406,N_7070);
nand U7567 (N_7567,N_7115,N_7437);
nand U7568 (N_7568,N_7244,N_7058);
nor U7569 (N_7569,N_7343,N_7210);
xnor U7570 (N_7570,N_7483,N_7328);
or U7571 (N_7571,N_7122,N_7396);
nand U7572 (N_7572,N_7045,N_7266);
or U7573 (N_7573,N_7100,N_7133);
xor U7574 (N_7574,N_7458,N_7077);
or U7575 (N_7575,N_7140,N_7101);
or U7576 (N_7576,N_7312,N_7392);
nand U7577 (N_7577,N_7250,N_7241);
and U7578 (N_7578,N_7179,N_7239);
xnor U7579 (N_7579,N_7040,N_7095);
and U7580 (N_7580,N_7263,N_7256);
nor U7581 (N_7581,N_7205,N_7440);
nor U7582 (N_7582,N_7270,N_7031);
and U7583 (N_7583,N_7439,N_7074);
xnor U7584 (N_7584,N_7121,N_7225);
and U7585 (N_7585,N_7498,N_7043);
nand U7586 (N_7586,N_7387,N_7365);
nor U7587 (N_7587,N_7417,N_7030);
or U7588 (N_7588,N_7466,N_7086);
xor U7589 (N_7589,N_7468,N_7146);
and U7590 (N_7590,N_7285,N_7062);
or U7591 (N_7591,N_7103,N_7248);
and U7592 (N_7592,N_7307,N_7278);
nor U7593 (N_7593,N_7277,N_7112);
or U7594 (N_7594,N_7361,N_7057);
nand U7595 (N_7595,N_7060,N_7433);
nand U7596 (N_7596,N_7289,N_7340);
nand U7597 (N_7597,N_7238,N_7160);
nor U7598 (N_7598,N_7038,N_7318);
and U7599 (N_7599,N_7491,N_7052);
or U7600 (N_7600,N_7423,N_7370);
nand U7601 (N_7601,N_7414,N_7400);
or U7602 (N_7602,N_7135,N_7302);
xor U7603 (N_7603,N_7326,N_7053);
or U7604 (N_7604,N_7310,N_7487);
nor U7605 (N_7605,N_7448,N_7041);
or U7606 (N_7606,N_7342,N_7384);
nand U7607 (N_7607,N_7454,N_7035);
xor U7608 (N_7608,N_7290,N_7150);
nor U7609 (N_7609,N_7233,N_7444);
nand U7610 (N_7610,N_7207,N_7461);
xor U7611 (N_7611,N_7174,N_7182);
nor U7612 (N_7612,N_7470,N_7332);
or U7613 (N_7613,N_7388,N_7269);
or U7614 (N_7614,N_7050,N_7066);
and U7615 (N_7615,N_7338,N_7164);
xnor U7616 (N_7616,N_7292,N_7463);
and U7617 (N_7617,N_7134,N_7175);
nand U7618 (N_7618,N_7022,N_7047);
xnor U7619 (N_7619,N_7357,N_7416);
and U7620 (N_7620,N_7378,N_7049);
and U7621 (N_7621,N_7251,N_7211);
xnor U7622 (N_7622,N_7486,N_7001);
xnor U7623 (N_7623,N_7367,N_7145);
and U7624 (N_7624,N_7373,N_7464);
or U7625 (N_7625,N_7494,N_7130);
or U7626 (N_7626,N_7158,N_7142);
nor U7627 (N_7627,N_7368,N_7098);
and U7628 (N_7628,N_7096,N_7333);
or U7629 (N_7629,N_7163,N_7245);
nor U7630 (N_7630,N_7405,N_7168);
or U7631 (N_7631,N_7495,N_7201);
xnor U7632 (N_7632,N_7311,N_7359);
nor U7633 (N_7633,N_7230,N_7177);
xnor U7634 (N_7634,N_7317,N_7181);
nand U7635 (N_7635,N_7024,N_7422);
xnor U7636 (N_7636,N_7484,N_7021);
nand U7637 (N_7637,N_7351,N_7217);
nand U7638 (N_7638,N_7390,N_7093);
nor U7639 (N_7639,N_7383,N_7374);
or U7640 (N_7640,N_7197,N_7296);
or U7641 (N_7641,N_7187,N_7229);
or U7642 (N_7642,N_7299,N_7253);
nand U7643 (N_7643,N_7489,N_7432);
and U7644 (N_7644,N_7394,N_7012);
and U7645 (N_7645,N_7132,N_7356);
and U7646 (N_7646,N_7202,N_7282);
xor U7647 (N_7647,N_7499,N_7274);
xor U7648 (N_7648,N_7306,N_7170);
nor U7649 (N_7649,N_7316,N_7349);
xnor U7650 (N_7650,N_7155,N_7375);
nand U7651 (N_7651,N_7048,N_7183);
and U7652 (N_7652,N_7313,N_7051);
or U7653 (N_7653,N_7257,N_7319);
or U7654 (N_7654,N_7192,N_7496);
xnor U7655 (N_7655,N_7127,N_7267);
nor U7656 (N_7656,N_7126,N_7309);
or U7657 (N_7657,N_7305,N_7082);
nand U7658 (N_7658,N_7459,N_7018);
or U7659 (N_7659,N_7149,N_7032);
xor U7660 (N_7660,N_7243,N_7085);
and U7661 (N_7661,N_7382,N_7194);
and U7662 (N_7662,N_7427,N_7492);
or U7663 (N_7663,N_7191,N_7204);
xnor U7664 (N_7664,N_7344,N_7184);
xnor U7665 (N_7665,N_7336,N_7071);
nor U7666 (N_7666,N_7015,N_7141);
or U7667 (N_7667,N_7273,N_7081);
xnor U7668 (N_7668,N_7219,N_7449);
and U7669 (N_7669,N_7123,N_7055);
xor U7670 (N_7670,N_7297,N_7189);
nor U7671 (N_7671,N_7153,N_7443);
nor U7672 (N_7672,N_7218,N_7171);
xor U7673 (N_7673,N_7275,N_7412);
nor U7674 (N_7674,N_7493,N_7418);
xor U7675 (N_7675,N_7401,N_7063);
nor U7676 (N_7676,N_7046,N_7027);
or U7677 (N_7677,N_7279,N_7117);
nor U7678 (N_7678,N_7013,N_7216);
and U7679 (N_7679,N_7065,N_7258);
or U7680 (N_7680,N_7460,N_7116);
or U7681 (N_7681,N_7420,N_7195);
nor U7682 (N_7682,N_7322,N_7482);
xor U7683 (N_7683,N_7325,N_7350);
and U7684 (N_7684,N_7358,N_7255);
xnor U7685 (N_7685,N_7393,N_7188);
xnor U7686 (N_7686,N_7334,N_7271);
nand U7687 (N_7687,N_7339,N_7259);
xnor U7688 (N_7688,N_7472,N_7222);
nand U7689 (N_7689,N_7407,N_7215);
and U7690 (N_7690,N_7119,N_7083);
or U7691 (N_7691,N_7213,N_7176);
xnor U7692 (N_7692,N_7002,N_7190);
xor U7693 (N_7693,N_7079,N_7072);
or U7694 (N_7694,N_7404,N_7075);
and U7695 (N_7695,N_7007,N_7226);
and U7696 (N_7696,N_7353,N_7261);
xor U7697 (N_7697,N_7262,N_7415);
nor U7698 (N_7698,N_7111,N_7480);
xnor U7699 (N_7699,N_7366,N_7421);
nor U7700 (N_7700,N_7485,N_7025);
or U7701 (N_7701,N_7280,N_7180);
or U7702 (N_7702,N_7419,N_7287);
xnor U7703 (N_7703,N_7020,N_7475);
and U7704 (N_7704,N_7331,N_7288);
and U7705 (N_7705,N_7346,N_7036);
or U7706 (N_7706,N_7159,N_7453);
xor U7707 (N_7707,N_7372,N_7249);
or U7708 (N_7708,N_7379,N_7455);
nor U7709 (N_7709,N_7438,N_7203);
nor U7710 (N_7710,N_7452,N_7246);
or U7711 (N_7711,N_7413,N_7301);
nand U7712 (N_7712,N_7185,N_7186);
xor U7713 (N_7713,N_7234,N_7125);
nor U7714 (N_7714,N_7113,N_7162);
nor U7715 (N_7715,N_7131,N_7451);
nor U7716 (N_7716,N_7431,N_7139);
or U7717 (N_7717,N_7281,N_7391);
and U7718 (N_7718,N_7044,N_7003);
or U7719 (N_7719,N_7084,N_7308);
and U7720 (N_7720,N_7042,N_7231);
and U7721 (N_7721,N_7397,N_7178);
nor U7722 (N_7722,N_7232,N_7091);
nand U7723 (N_7723,N_7323,N_7033);
and U7724 (N_7724,N_7327,N_7061);
nor U7725 (N_7725,N_7105,N_7120);
and U7726 (N_7726,N_7107,N_7151);
and U7727 (N_7727,N_7293,N_7104);
or U7728 (N_7728,N_7321,N_7457);
or U7729 (N_7729,N_7442,N_7399);
xnor U7730 (N_7730,N_7198,N_7109);
and U7731 (N_7731,N_7054,N_7172);
nand U7732 (N_7732,N_7037,N_7068);
or U7733 (N_7733,N_7166,N_7362);
xor U7734 (N_7734,N_7059,N_7088);
xor U7735 (N_7735,N_7476,N_7283);
or U7736 (N_7736,N_7426,N_7456);
nand U7737 (N_7737,N_7398,N_7381);
nor U7738 (N_7738,N_7408,N_7364);
nand U7739 (N_7739,N_7410,N_7347);
or U7740 (N_7740,N_7348,N_7320);
nand U7741 (N_7741,N_7173,N_7028);
nand U7742 (N_7742,N_7337,N_7196);
nand U7743 (N_7743,N_7080,N_7023);
or U7744 (N_7744,N_7161,N_7014);
or U7745 (N_7745,N_7488,N_7208);
nor U7746 (N_7746,N_7352,N_7206);
nand U7747 (N_7747,N_7477,N_7010);
and U7748 (N_7748,N_7124,N_7402);
nor U7749 (N_7749,N_7355,N_7314);
and U7750 (N_7750,N_7313,N_7123);
nor U7751 (N_7751,N_7054,N_7312);
nand U7752 (N_7752,N_7180,N_7101);
nor U7753 (N_7753,N_7050,N_7422);
nand U7754 (N_7754,N_7276,N_7018);
nand U7755 (N_7755,N_7048,N_7401);
nand U7756 (N_7756,N_7371,N_7192);
or U7757 (N_7757,N_7209,N_7355);
nand U7758 (N_7758,N_7287,N_7386);
and U7759 (N_7759,N_7150,N_7206);
or U7760 (N_7760,N_7167,N_7277);
and U7761 (N_7761,N_7266,N_7154);
and U7762 (N_7762,N_7308,N_7349);
or U7763 (N_7763,N_7280,N_7227);
nor U7764 (N_7764,N_7435,N_7130);
xnor U7765 (N_7765,N_7463,N_7065);
and U7766 (N_7766,N_7454,N_7481);
nand U7767 (N_7767,N_7314,N_7171);
or U7768 (N_7768,N_7166,N_7286);
or U7769 (N_7769,N_7078,N_7342);
and U7770 (N_7770,N_7071,N_7108);
and U7771 (N_7771,N_7161,N_7081);
nand U7772 (N_7772,N_7081,N_7477);
or U7773 (N_7773,N_7048,N_7376);
nand U7774 (N_7774,N_7394,N_7115);
and U7775 (N_7775,N_7045,N_7193);
xor U7776 (N_7776,N_7032,N_7235);
or U7777 (N_7777,N_7058,N_7313);
nor U7778 (N_7778,N_7012,N_7058);
nor U7779 (N_7779,N_7390,N_7101);
and U7780 (N_7780,N_7413,N_7177);
nand U7781 (N_7781,N_7136,N_7496);
or U7782 (N_7782,N_7067,N_7195);
xnor U7783 (N_7783,N_7454,N_7163);
nand U7784 (N_7784,N_7484,N_7152);
xnor U7785 (N_7785,N_7316,N_7134);
and U7786 (N_7786,N_7306,N_7224);
nand U7787 (N_7787,N_7197,N_7243);
xor U7788 (N_7788,N_7331,N_7083);
nor U7789 (N_7789,N_7315,N_7084);
nand U7790 (N_7790,N_7281,N_7324);
xnor U7791 (N_7791,N_7015,N_7098);
nand U7792 (N_7792,N_7014,N_7312);
nor U7793 (N_7793,N_7385,N_7014);
xnor U7794 (N_7794,N_7314,N_7245);
nand U7795 (N_7795,N_7279,N_7461);
xor U7796 (N_7796,N_7049,N_7301);
xnor U7797 (N_7797,N_7071,N_7074);
nand U7798 (N_7798,N_7285,N_7159);
xnor U7799 (N_7799,N_7241,N_7472);
and U7800 (N_7800,N_7370,N_7391);
and U7801 (N_7801,N_7480,N_7180);
nor U7802 (N_7802,N_7038,N_7450);
nand U7803 (N_7803,N_7286,N_7450);
nand U7804 (N_7804,N_7416,N_7131);
and U7805 (N_7805,N_7232,N_7051);
and U7806 (N_7806,N_7229,N_7399);
and U7807 (N_7807,N_7452,N_7134);
xor U7808 (N_7808,N_7141,N_7061);
xor U7809 (N_7809,N_7176,N_7497);
xor U7810 (N_7810,N_7257,N_7284);
xor U7811 (N_7811,N_7364,N_7167);
nand U7812 (N_7812,N_7272,N_7121);
nand U7813 (N_7813,N_7225,N_7024);
and U7814 (N_7814,N_7381,N_7223);
nor U7815 (N_7815,N_7378,N_7407);
or U7816 (N_7816,N_7364,N_7292);
or U7817 (N_7817,N_7329,N_7045);
xnor U7818 (N_7818,N_7164,N_7284);
nor U7819 (N_7819,N_7050,N_7210);
nor U7820 (N_7820,N_7175,N_7348);
nor U7821 (N_7821,N_7496,N_7299);
nand U7822 (N_7822,N_7122,N_7325);
nor U7823 (N_7823,N_7109,N_7027);
nor U7824 (N_7824,N_7006,N_7223);
xor U7825 (N_7825,N_7073,N_7128);
or U7826 (N_7826,N_7241,N_7402);
and U7827 (N_7827,N_7400,N_7425);
xor U7828 (N_7828,N_7397,N_7057);
xnor U7829 (N_7829,N_7093,N_7195);
or U7830 (N_7830,N_7036,N_7187);
or U7831 (N_7831,N_7448,N_7355);
xnor U7832 (N_7832,N_7226,N_7199);
or U7833 (N_7833,N_7271,N_7034);
xnor U7834 (N_7834,N_7303,N_7329);
nor U7835 (N_7835,N_7215,N_7064);
and U7836 (N_7836,N_7438,N_7409);
nand U7837 (N_7837,N_7117,N_7071);
and U7838 (N_7838,N_7262,N_7104);
nor U7839 (N_7839,N_7455,N_7236);
and U7840 (N_7840,N_7311,N_7334);
xor U7841 (N_7841,N_7161,N_7494);
xor U7842 (N_7842,N_7326,N_7320);
xor U7843 (N_7843,N_7131,N_7125);
xnor U7844 (N_7844,N_7394,N_7481);
xnor U7845 (N_7845,N_7499,N_7401);
nor U7846 (N_7846,N_7012,N_7049);
and U7847 (N_7847,N_7158,N_7427);
xor U7848 (N_7848,N_7011,N_7097);
xnor U7849 (N_7849,N_7482,N_7126);
or U7850 (N_7850,N_7287,N_7075);
and U7851 (N_7851,N_7079,N_7322);
and U7852 (N_7852,N_7355,N_7433);
xor U7853 (N_7853,N_7374,N_7126);
nand U7854 (N_7854,N_7228,N_7343);
nand U7855 (N_7855,N_7127,N_7453);
nor U7856 (N_7856,N_7142,N_7439);
nor U7857 (N_7857,N_7339,N_7432);
or U7858 (N_7858,N_7274,N_7057);
and U7859 (N_7859,N_7114,N_7278);
xnor U7860 (N_7860,N_7105,N_7438);
xnor U7861 (N_7861,N_7241,N_7158);
xnor U7862 (N_7862,N_7492,N_7403);
or U7863 (N_7863,N_7430,N_7270);
or U7864 (N_7864,N_7302,N_7232);
and U7865 (N_7865,N_7039,N_7262);
nand U7866 (N_7866,N_7278,N_7101);
nand U7867 (N_7867,N_7007,N_7330);
or U7868 (N_7868,N_7435,N_7395);
xnor U7869 (N_7869,N_7399,N_7489);
nor U7870 (N_7870,N_7033,N_7417);
xor U7871 (N_7871,N_7311,N_7375);
nor U7872 (N_7872,N_7095,N_7224);
or U7873 (N_7873,N_7329,N_7238);
xor U7874 (N_7874,N_7282,N_7101);
xnor U7875 (N_7875,N_7299,N_7135);
xnor U7876 (N_7876,N_7264,N_7109);
or U7877 (N_7877,N_7040,N_7104);
nand U7878 (N_7878,N_7286,N_7147);
nor U7879 (N_7879,N_7355,N_7310);
and U7880 (N_7880,N_7130,N_7017);
and U7881 (N_7881,N_7245,N_7379);
xnor U7882 (N_7882,N_7059,N_7261);
nor U7883 (N_7883,N_7045,N_7134);
nor U7884 (N_7884,N_7393,N_7125);
nand U7885 (N_7885,N_7288,N_7157);
nor U7886 (N_7886,N_7202,N_7228);
or U7887 (N_7887,N_7414,N_7450);
nand U7888 (N_7888,N_7383,N_7088);
and U7889 (N_7889,N_7005,N_7343);
xnor U7890 (N_7890,N_7022,N_7317);
nand U7891 (N_7891,N_7497,N_7460);
nor U7892 (N_7892,N_7395,N_7224);
xor U7893 (N_7893,N_7091,N_7115);
nand U7894 (N_7894,N_7010,N_7183);
nor U7895 (N_7895,N_7490,N_7423);
xnor U7896 (N_7896,N_7495,N_7305);
or U7897 (N_7897,N_7319,N_7177);
nor U7898 (N_7898,N_7087,N_7431);
or U7899 (N_7899,N_7054,N_7438);
or U7900 (N_7900,N_7261,N_7043);
nand U7901 (N_7901,N_7189,N_7338);
nand U7902 (N_7902,N_7077,N_7158);
or U7903 (N_7903,N_7296,N_7104);
nor U7904 (N_7904,N_7215,N_7435);
nand U7905 (N_7905,N_7391,N_7173);
or U7906 (N_7906,N_7365,N_7062);
and U7907 (N_7907,N_7173,N_7217);
nand U7908 (N_7908,N_7361,N_7152);
nand U7909 (N_7909,N_7248,N_7480);
nor U7910 (N_7910,N_7148,N_7136);
xor U7911 (N_7911,N_7294,N_7070);
nand U7912 (N_7912,N_7318,N_7217);
or U7913 (N_7913,N_7172,N_7408);
or U7914 (N_7914,N_7241,N_7373);
xor U7915 (N_7915,N_7468,N_7056);
or U7916 (N_7916,N_7377,N_7155);
and U7917 (N_7917,N_7245,N_7169);
xnor U7918 (N_7918,N_7146,N_7194);
and U7919 (N_7919,N_7450,N_7056);
and U7920 (N_7920,N_7261,N_7368);
or U7921 (N_7921,N_7356,N_7212);
or U7922 (N_7922,N_7145,N_7120);
or U7923 (N_7923,N_7443,N_7053);
xor U7924 (N_7924,N_7311,N_7332);
and U7925 (N_7925,N_7153,N_7460);
xnor U7926 (N_7926,N_7296,N_7200);
xnor U7927 (N_7927,N_7149,N_7478);
and U7928 (N_7928,N_7047,N_7474);
and U7929 (N_7929,N_7106,N_7253);
or U7930 (N_7930,N_7347,N_7110);
xor U7931 (N_7931,N_7330,N_7193);
xnor U7932 (N_7932,N_7196,N_7134);
xor U7933 (N_7933,N_7331,N_7482);
and U7934 (N_7934,N_7228,N_7072);
and U7935 (N_7935,N_7153,N_7314);
xor U7936 (N_7936,N_7223,N_7073);
or U7937 (N_7937,N_7364,N_7154);
and U7938 (N_7938,N_7372,N_7102);
and U7939 (N_7939,N_7284,N_7018);
nor U7940 (N_7940,N_7285,N_7466);
nand U7941 (N_7941,N_7189,N_7346);
nand U7942 (N_7942,N_7012,N_7402);
and U7943 (N_7943,N_7154,N_7361);
xnor U7944 (N_7944,N_7484,N_7225);
nand U7945 (N_7945,N_7392,N_7395);
or U7946 (N_7946,N_7287,N_7341);
or U7947 (N_7947,N_7254,N_7285);
nand U7948 (N_7948,N_7264,N_7091);
xor U7949 (N_7949,N_7381,N_7121);
and U7950 (N_7950,N_7373,N_7466);
nor U7951 (N_7951,N_7462,N_7491);
xor U7952 (N_7952,N_7498,N_7294);
xor U7953 (N_7953,N_7055,N_7198);
or U7954 (N_7954,N_7214,N_7087);
xnor U7955 (N_7955,N_7104,N_7498);
or U7956 (N_7956,N_7004,N_7201);
nor U7957 (N_7957,N_7015,N_7131);
nor U7958 (N_7958,N_7479,N_7418);
xor U7959 (N_7959,N_7155,N_7225);
and U7960 (N_7960,N_7330,N_7368);
xnor U7961 (N_7961,N_7236,N_7299);
nand U7962 (N_7962,N_7222,N_7129);
xnor U7963 (N_7963,N_7201,N_7341);
or U7964 (N_7964,N_7338,N_7314);
nand U7965 (N_7965,N_7162,N_7443);
xor U7966 (N_7966,N_7064,N_7294);
nor U7967 (N_7967,N_7369,N_7007);
or U7968 (N_7968,N_7155,N_7455);
and U7969 (N_7969,N_7304,N_7289);
nand U7970 (N_7970,N_7098,N_7046);
nand U7971 (N_7971,N_7279,N_7302);
or U7972 (N_7972,N_7103,N_7453);
nor U7973 (N_7973,N_7497,N_7120);
nand U7974 (N_7974,N_7209,N_7041);
nand U7975 (N_7975,N_7128,N_7228);
xor U7976 (N_7976,N_7391,N_7440);
or U7977 (N_7977,N_7211,N_7488);
nor U7978 (N_7978,N_7186,N_7028);
and U7979 (N_7979,N_7167,N_7321);
or U7980 (N_7980,N_7062,N_7303);
xor U7981 (N_7981,N_7079,N_7066);
or U7982 (N_7982,N_7049,N_7443);
xnor U7983 (N_7983,N_7046,N_7167);
and U7984 (N_7984,N_7363,N_7200);
xor U7985 (N_7985,N_7086,N_7236);
nand U7986 (N_7986,N_7070,N_7344);
or U7987 (N_7987,N_7045,N_7263);
nand U7988 (N_7988,N_7471,N_7100);
and U7989 (N_7989,N_7250,N_7133);
and U7990 (N_7990,N_7370,N_7246);
nor U7991 (N_7991,N_7234,N_7367);
and U7992 (N_7992,N_7322,N_7344);
and U7993 (N_7993,N_7347,N_7134);
and U7994 (N_7994,N_7367,N_7236);
xnor U7995 (N_7995,N_7189,N_7171);
nor U7996 (N_7996,N_7115,N_7036);
nand U7997 (N_7997,N_7319,N_7424);
nand U7998 (N_7998,N_7107,N_7396);
xor U7999 (N_7999,N_7439,N_7292);
or U8000 (N_8000,N_7903,N_7747);
or U8001 (N_8001,N_7649,N_7929);
nand U8002 (N_8002,N_7917,N_7622);
and U8003 (N_8003,N_7686,N_7807);
nand U8004 (N_8004,N_7783,N_7715);
nand U8005 (N_8005,N_7605,N_7897);
and U8006 (N_8006,N_7533,N_7771);
nand U8007 (N_8007,N_7583,N_7642);
or U8008 (N_8008,N_7581,N_7837);
xor U8009 (N_8009,N_7600,N_7976);
or U8010 (N_8010,N_7597,N_7697);
and U8011 (N_8011,N_7626,N_7617);
and U8012 (N_8012,N_7639,N_7623);
nand U8013 (N_8013,N_7789,N_7908);
xor U8014 (N_8014,N_7750,N_7734);
nor U8015 (N_8015,N_7966,N_7518);
and U8016 (N_8016,N_7914,N_7778);
or U8017 (N_8017,N_7863,N_7776);
xnor U8018 (N_8018,N_7873,N_7958);
nor U8019 (N_8019,N_7509,N_7521);
nand U8020 (N_8020,N_7843,N_7792);
and U8021 (N_8021,N_7551,N_7636);
nand U8022 (N_8022,N_7894,N_7749);
or U8023 (N_8023,N_7969,N_7695);
and U8024 (N_8024,N_7785,N_7865);
nand U8025 (N_8025,N_7670,N_7585);
xnor U8026 (N_8026,N_7540,N_7943);
or U8027 (N_8027,N_7510,N_7650);
nor U8028 (N_8028,N_7885,N_7919);
nand U8029 (N_8029,N_7543,N_7504);
and U8030 (N_8030,N_7683,N_7514);
nand U8031 (N_8031,N_7840,N_7982);
nor U8032 (N_8032,N_7796,N_7502);
xnor U8033 (N_8033,N_7564,N_7962);
nand U8034 (N_8034,N_7631,N_7781);
nor U8035 (N_8035,N_7531,N_7950);
or U8036 (N_8036,N_7580,N_7916);
or U8037 (N_8037,N_7800,N_7710);
and U8038 (N_8038,N_7856,N_7822);
nand U8039 (N_8039,N_7530,N_7983);
nor U8040 (N_8040,N_7755,N_7714);
xnor U8041 (N_8041,N_7938,N_7845);
xnor U8042 (N_8042,N_7604,N_7759);
and U8043 (N_8043,N_7944,N_7911);
or U8044 (N_8044,N_7980,N_7861);
nand U8045 (N_8045,N_7555,N_7978);
or U8046 (N_8046,N_7891,N_7561);
xor U8047 (N_8047,N_7782,N_7507);
or U8048 (N_8048,N_7816,N_7556);
and U8049 (N_8049,N_7529,N_7732);
and U8050 (N_8050,N_7820,N_7939);
and U8051 (N_8051,N_7888,N_7562);
or U8052 (N_8052,N_7606,N_7825);
nor U8053 (N_8053,N_7501,N_7754);
and U8054 (N_8054,N_7515,N_7904);
or U8055 (N_8055,N_7691,N_7779);
xor U8056 (N_8056,N_7967,N_7788);
or U8057 (N_8057,N_7989,N_7599);
nor U8058 (N_8058,N_7954,N_7591);
xnor U8059 (N_8059,N_7932,N_7602);
or U8060 (N_8060,N_7769,N_7548);
nor U8061 (N_8061,N_7620,N_7719);
nor U8062 (N_8062,N_7557,N_7974);
and U8063 (N_8063,N_7860,N_7651);
or U8064 (N_8064,N_7610,N_7787);
xnor U8065 (N_8065,N_7965,N_7831);
or U8066 (N_8066,N_7640,N_7508);
nand U8067 (N_8067,N_7726,N_7669);
nor U8068 (N_8068,N_7731,N_7842);
or U8069 (N_8069,N_7678,N_7665);
and U8070 (N_8070,N_7575,N_7853);
xor U8071 (N_8071,N_7641,N_7573);
nand U8072 (N_8072,N_7828,N_7574);
or U8073 (N_8073,N_7560,N_7524);
xnor U8074 (N_8074,N_7659,N_7536);
and U8075 (N_8075,N_7798,N_7517);
or U8076 (N_8076,N_7957,N_7857);
xor U8077 (N_8077,N_7777,N_7871);
and U8078 (N_8078,N_7823,N_7542);
and U8079 (N_8079,N_7698,N_7702);
xor U8080 (N_8080,N_7892,N_7993);
nor U8081 (N_8081,N_7968,N_7513);
nor U8082 (N_8082,N_7544,N_7748);
xor U8083 (N_8083,N_7721,N_7538);
and U8084 (N_8084,N_7537,N_7752);
and U8085 (N_8085,N_7723,N_7793);
xnor U8086 (N_8086,N_7987,N_7883);
nor U8087 (N_8087,N_7770,N_7925);
or U8088 (N_8088,N_7913,N_7701);
nand U8089 (N_8089,N_7708,N_7619);
or U8090 (N_8090,N_7689,N_7578);
nand U8091 (N_8091,N_7625,N_7566);
xor U8092 (N_8092,N_7762,N_7907);
nand U8093 (N_8093,N_7528,N_7775);
or U8094 (N_8094,N_7884,N_7616);
nand U8095 (N_8095,N_7572,N_7571);
or U8096 (N_8096,N_7512,N_7826);
and U8097 (N_8097,N_7746,N_7926);
nor U8098 (N_8098,N_7935,N_7952);
nand U8099 (N_8099,N_7921,N_7733);
nor U8100 (N_8100,N_7841,N_7608);
and U8101 (N_8101,N_7881,N_7844);
nand U8102 (N_8102,N_7963,N_7811);
or U8103 (N_8103,N_7964,N_7658);
nor U8104 (N_8104,N_7614,N_7643);
nand U8105 (N_8105,N_7764,N_7946);
xor U8106 (N_8106,N_7931,N_7886);
and U8107 (N_8107,N_7985,N_7900);
and U8108 (N_8108,N_7596,N_7687);
xnor U8109 (N_8109,N_7955,N_7933);
nand U8110 (N_8110,N_7744,N_7997);
xnor U8111 (N_8111,N_7549,N_7677);
or U8112 (N_8112,N_7868,N_7986);
nand U8113 (N_8113,N_7738,N_7766);
or U8114 (N_8114,N_7835,N_7864);
nor U8115 (N_8115,N_7672,N_7657);
and U8116 (N_8116,N_7582,N_7662);
nand U8117 (N_8117,N_7654,N_7869);
and U8118 (N_8118,N_7674,N_7615);
and U8119 (N_8119,N_7712,N_7682);
xor U8120 (N_8120,N_7526,N_7799);
nand U8121 (N_8121,N_7628,N_7730);
nand U8122 (N_8122,N_7772,N_7603);
nand U8123 (N_8123,N_7924,N_7696);
or U8124 (N_8124,N_7713,N_7645);
and U8125 (N_8125,N_7711,N_7994);
xnor U8126 (N_8126,N_7898,N_7758);
nand U8127 (N_8127,N_7589,N_7804);
and U8128 (N_8128,N_7768,N_7613);
nand U8129 (N_8129,N_7829,N_7813);
nor U8130 (N_8130,N_7960,N_7739);
nand U8131 (N_8131,N_7821,N_7928);
or U8132 (N_8132,N_7652,N_7920);
nand U8133 (N_8133,N_7506,N_7527);
nand U8134 (N_8134,N_7927,N_7761);
or U8135 (N_8135,N_7996,N_7814);
and U8136 (N_8136,N_7790,N_7902);
or U8137 (N_8137,N_7848,N_7534);
and U8138 (N_8138,N_7847,N_7663);
nand U8139 (N_8139,N_7972,N_7661);
xnor U8140 (N_8140,N_7786,N_7523);
nand U8141 (N_8141,N_7593,N_7791);
and U8142 (N_8142,N_7618,N_7638);
xor U8143 (N_8143,N_7552,N_7675);
xnor U8144 (N_8144,N_7751,N_7520);
xor U8145 (N_8145,N_7546,N_7878);
or U8146 (N_8146,N_7977,N_7569);
nand U8147 (N_8147,N_7539,N_7707);
and U8148 (N_8148,N_7889,N_7765);
or U8149 (N_8149,N_7653,N_7817);
xnor U8150 (N_8150,N_7554,N_7901);
nand U8151 (N_8151,N_7601,N_7999);
xnor U8152 (N_8152,N_7718,N_7949);
nand U8153 (N_8153,N_7780,N_7809);
xnor U8154 (N_8154,N_7936,N_7852);
xor U8155 (N_8155,N_7541,N_7699);
or U8156 (N_8156,N_7704,N_7722);
xor U8157 (N_8157,N_7700,N_7671);
nor U8158 (N_8158,N_7995,N_7934);
nor U8159 (N_8159,N_7953,N_7680);
and U8160 (N_8160,N_7627,N_7849);
and U8161 (N_8161,N_7558,N_7930);
xor U8162 (N_8162,N_7630,N_7991);
nor U8163 (N_8163,N_7612,N_7893);
nand U8164 (N_8164,N_7611,N_7525);
nand U8165 (N_8165,N_7945,N_7984);
nor U8166 (N_8166,N_7729,N_7644);
or U8167 (N_8167,N_7879,N_7942);
xnor U8168 (N_8168,N_7815,N_7915);
xor U8169 (N_8169,N_7547,N_7896);
or U8170 (N_8170,N_7988,N_7668);
nand U8171 (N_8171,N_7875,N_7516);
and U8172 (N_8172,N_7660,N_7688);
or U8173 (N_8173,N_7545,N_7767);
and U8174 (N_8174,N_7895,N_7819);
or U8175 (N_8175,N_7839,N_7757);
xnor U8176 (N_8176,N_7940,N_7784);
or U8177 (N_8177,N_7947,N_7808);
nor U8178 (N_8178,N_7805,N_7629);
or U8179 (N_8179,N_7676,N_7632);
xor U8180 (N_8180,N_7836,N_7576);
or U8181 (N_8181,N_7801,N_7690);
nand U8182 (N_8182,N_7740,N_7961);
nor U8183 (N_8183,N_7812,N_7609);
or U8184 (N_8184,N_7909,N_7664);
xor U8185 (N_8185,N_7838,N_7797);
nor U8186 (N_8186,N_7855,N_7563);
nand U8187 (N_8187,N_7773,N_7876);
nor U8188 (N_8188,N_7553,N_7727);
xnor U8189 (N_8189,N_7567,N_7854);
or U8190 (N_8190,N_7763,N_7590);
nor U8191 (N_8191,N_7866,N_7979);
or U8192 (N_8192,N_7586,N_7753);
nand U8193 (N_8193,N_7906,N_7693);
or U8194 (N_8194,N_7834,N_7874);
and U8195 (N_8195,N_7720,N_7795);
nor U8196 (N_8196,N_7832,N_7736);
and U8197 (N_8197,N_7511,N_7912);
nand U8198 (N_8198,N_7890,N_7685);
nand U8199 (N_8199,N_7519,N_7568);
and U8200 (N_8200,N_7635,N_7634);
nand U8201 (N_8201,N_7637,N_7716);
nor U8202 (N_8202,N_7703,N_7910);
or U8203 (N_8203,N_7532,N_7948);
and U8204 (N_8204,N_7565,N_7802);
nand U8205 (N_8205,N_7503,N_7922);
nand U8206 (N_8206,N_7877,N_7656);
and U8207 (N_8207,N_7973,N_7717);
xor U8208 (N_8208,N_7998,N_7918);
nand U8209 (N_8209,N_7742,N_7887);
nand U8210 (N_8210,N_7743,N_7810);
nor U8211 (N_8211,N_7937,N_7830);
nor U8212 (N_8212,N_7846,N_7741);
and U8213 (N_8213,N_7706,N_7880);
or U8214 (N_8214,N_7647,N_7550);
or U8215 (N_8215,N_7760,N_7794);
and U8216 (N_8216,N_7607,N_7679);
nand U8217 (N_8217,N_7858,N_7595);
nand U8218 (N_8218,N_7981,N_7774);
nor U8219 (N_8219,N_7756,N_7971);
nand U8220 (N_8220,N_7941,N_7850);
xor U8221 (N_8221,N_7522,N_7870);
xnor U8222 (N_8222,N_7818,N_7990);
nand U8223 (N_8223,N_7633,N_7588);
and U8224 (N_8224,N_7673,N_7737);
and U8225 (N_8225,N_7724,N_7694);
xnor U8226 (N_8226,N_7592,N_7970);
and U8227 (N_8227,N_7905,N_7505);
nand U8228 (N_8228,N_7882,N_7725);
nand U8229 (N_8229,N_7584,N_7624);
nand U8230 (N_8230,N_7598,N_7621);
nor U8231 (N_8231,N_7867,N_7728);
xor U8232 (N_8232,N_7587,N_7500);
and U8233 (N_8233,N_7667,N_7579);
or U8234 (N_8234,N_7594,N_7570);
nand U8235 (N_8235,N_7681,N_7735);
nand U8236 (N_8236,N_7806,N_7824);
or U8237 (N_8237,N_7577,N_7851);
nand U8238 (N_8238,N_7646,N_7803);
and U8239 (N_8239,N_7535,N_7648);
and U8240 (N_8240,N_7692,N_7992);
or U8241 (N_8241,N_7862,N_7709);
nor U8242 (N_8242,N_7899,N_7872);
nand U8243 (N_8243,N_7975,N_7923);
nand U8244 (N_8244,N_7655,N_7684);
or U8245 (N_8245,N_7745,N_7833);
nand U8246 (N_8246,N_7959,N_7859);
and U8247 (N_8247,N_7956,N_7705);
nand U8248 (N_8248,N_7951,N_7666);
xnor U8249 (N_8249,N_7827,N_7559);
nor U8250 (N_8250,N_7590,N_7649);
nand U8251 (N_8251,N_7575,N_7531);
nor U8252 (N_8252,N_7805,N_7580);
or U8253 (N_8253,N_7553,N_7775);
nor U8254 (N_8254,N_7640,N_7922);
nor U8255 (N_8255,N_7596,N_7932);
nand U8256 (N_8256,N_7709,N_7943);
or U8257 (N_8257,N_7760,N_7868);
nand U8258 (N_8258,N_7500,N_7957);
nor U8259 (N_8259,N_7763,N_7753);
xnor U8260 (N_8260,N_7503,N_7798);
nand U8261 (N_8261,N_7735,N_7918);
nand U8262 (N_8262,N_7570,N_7575);
nand U8263 (N_8263,N_7943,N_7666);
xnor U8264 (N_8264,N_7558,N_7698);
and U8265 (N_8265,N_7984,N_7795);
nand U8266 (N_8266,N_7767,N_7779);
xnor U8267 (N_8267,N_7752,N_7992);
and U8268 (N_8268,N_7619,N_7767);
xnor U8269 (N_8269,N_7592,N_7855);
xnor U8270 (N_8270,N_7916,N_7899);
nor U8271 (N_8271,N_7700,N_7746);
or U8272 (N_8272,N_7504,N_7621);
and U8273 (N_8273,N_7612,N_7596);
or U8274 (N_8274,N_7833,N_7876);
nand U8275 (N_8275,N_7575,N_7982);
nand U8276 (N_8276,N_7916,N_7605);
xnor U8277 (N_8277,N_7775,N_7523);
and U8278 (N_8278,N_7641,N_7620);
or U8279 (N_8279,N_7781,N_7699);
nand U8280 (N_8280,N_7835,N_7605);
or U8281 (N_8281,N_7829,N_7816);
nand U8282 (N_8282,N_7544,N_7873);
or U8283 (N_8283,N_7717,N_7508);
nor U8284 (N_8284,N_7690,N_7735);
nor U8285 (N_8285,N_7939,N_7690);
and U8286 (N_8286,N_7773,N_7886);
or U8287 (N_8287,N_7804,N_7952);
nor U8288 (N_8288,N_7919,N_7837);
and U8289 (N_8289,N_7977,N_7792);
nand U8290 (N_8290,N_7701,N_7884);
nor U8291 (N_8291,N_7877,N_7544);
nand U8292 (N_8292,N_7978,N_7795);
or U8293 (N_8293,N_7999,N_7958);
and U8294 (N_8294,N_7587,N_7941);
nor U8295 (N_8295,N_7552,N_7659);
or U8296 (N_8296,N_7961,N_7544);
nor U8297 (N_8297,N_7689,N_7691);
nand U8298 (N_8298,N_7963,N_7668);
xnor U8299 (N_8299,N_7802,N_7858);
or U8300 (N_8300,N_7969,N_7642);
nand U8301 (N_8301,N_7627,N_7572);
or U8302 (N_8302,N_7743,N_7554);
and U8303 (N_8303,N_7926,N_7713);
and U8304 (N_8304,N_7757,N_7516);
nor U8305 (N_8305,N_7760,N_7890);
or U8306 (N_8306,N_7997,N_7516);
and U8307 (N_8307,N_7986,N_7588);
and U8308 (N_8308,N_7953,N_7821);
nor U8309 (N_8309,N_7969,N_7593);
nor U8310 (N_8310,N_7522,N_7726);
xor U8311 (N_8311,N_7785,N_7981);
or U8312 (N_8312,N_7763,N_7871);
or U8313 (N_8313,N_7926,N_7982);
xnor U8314 (N_8314,N_7582,N_7768);
nor U8315 (N_8315,N_7969,N_7551);
or U8316 (N_8316,N_7599,N_7813);
and U8317 (N_8317,N_7648,N_7730);
nor U8318 (N_8318,N_7884,N_7925);
xor U8319 (N_8319,N_7794,N_7564);
xor U8320 (N_8320,N_7995,N_7970);
and U8321 (N_8321,N_7687,N_7947);
nor U8322 (N_8322,N_7649,N_7864);
or U8323 (N_8323,N_7580,N_7654);
nor U8324 (N_8324,N_7827,N_7605);
or U8325 (N_8325,N_7888,N_7702);
and U8326 (N_8326,N_7609,N_7732);
xor U8327 (N_8327,N_7770,N_7951);
and U8328 (N_8328,N_7793,N_7736);
nand U8329 (N_8329,N_7991,N_7613);
xnor U8330 (N_8330,N_7741,N_7874);
and U8331 (N_8331,N_7608,N_7552);
xnor U8332 (N_8332,N_7726,N_7803);
xnor U8333 (N_8333,N_7513,N_7827);
or U8334 (N_8334,N_7933,N_7712);
nand U8335 (N_8335,N_7771,N_7583);
or U8336 (N_8336,N_7891,N_7555);
and U8337 (N_8337,N_7937,N_7844);
or U8338 (N_8338,N_7981,N_7980);
or U8339 (N_8339,N_7644,N_7918);
xnor U8340 (N_8340,N_7971,N_7514);
nor U8341 (N_8341,N_7995,N_7762);
nor U8342 (N_8342,N_7842,N_7717);
nor U8343 (N_8343,N_7725,N_7946);
or U8344 (N_8344,N_7825,N_7687);
or U8345 (N_8345,N_7806,N_7816);
nor U8346 (N_8346,N_7929,N_7940);
nand U8347 (N_8347,N_7902,N_7862);
or U8348 (N_8348,N_7748,N_7547);
nand U8349 (N_8349,N_7986,N_7540);
nand U8350 (N_8350,N_7725,N_7919);
and U8351 (N_8351,N_7972,N_7630);
nor U8352 (N_8352,N_7624,N_7758);
nand U8353 (N_8353,N_7759,N_7601);
xor U8354 (N_8354,N_7620,N_7709);
xnor U8355 (N_8355,N_7744,N_7814);
or U8356 (N_8356,N_7657,N_7956);
or U8357 (N_8357,N_7659,N_7948);
xor U8358 (N_8358,N_7601,N_7917);
xor U8359 (N_8359,N_7842,N_7682);
and U8360 (N_8360,N_7588,N_7561);
nor U8361 (N_8361,N_7740,N_7577);
and U8362 (N_8362,N_7679,N_7672);
nor U8363 (N_8363,N_7641,N_7955);
nand U8364 (N_8364,N_7555,N_7778);
and U8365 (N_8365,N_7704,N_7937);
nand U8366 (N_8366,N_7721,N_7964);
xor U8367 (N_8367,N_7941,N_7803);
and U8368 (N_8368,N_7717,N_7583);
xor U8369 (N_8369,N_7866,N_7579);
nand U8370 (N_8370,N_7769,N_7651);
xnor U8371 (N_8371,N_7773,N_7849);
xor U8372 (N_8372,N_7819,N_7967);
or U8373 (N_8373,N_7948,N_7516);
or U8374 (N_8374,N_7818,N_7525);
and U8375 (N_8375,N_7581,N_7529);
nand U8376 (N_8376,N_7530,N_7696);
xnor U8377 (N_8377,N_7730,N_7783);
nor U8378 (N_8378,N_7622,N_7810);
nor U8379 (N_8379,N_7519,N_7993);
and U8380 (N_8380,N_7553,N_7806);
xnor U8381 (N_8381,N_7685,N_7633);
or U8382 (N_8382,N_7869,N_7902);
and U8383 (N_8383,N_7581,N_7667);
nand U8384 (N_8384,N_7903,N_7674);
xnor U8385 (N_8385,N_7652,N_7723);
xor U8386 (N_8386,N_7642,N_7903);
nand U8387 (N_8387,N_7914,N_7753);
or U8388 (N_8388,N_7683,N_7792);
or U8389 (N_8389,N_7632,N_7928);
nor U8390 (N_8390,N_7987,N_7538);
nor U8391 (N_8391,N_7771,N_7609);
xor U8392 (N_8392,N_7603,N_7758);
or U8393 (N_8393,N_7600,N_7655);
xor U8394 (N_8394,N_7712,N_7975);
and U8395 (N_8395,N_7582,N_7775);
nand U8396 (N_8396,N_7736,N_7798);
xnor U8397 (N_8397,N_7995,N_7518);
nand U8398 (N_8398,N_7629,N_7641);
nand U8399 (N_8399,N_7696,N_7618);
or U8400 (N_8400,N_7960,N_7916);
nor U8401 (N_8401,N_7982,N_7723);
and U8402 (N_8402,N_7873,N_7845);
nor U8403 (N_8403,N_7630,N_7617);
or U8404 (N_8404,N_7715,N_7659);
and U8405 (N_8405,N_7564,N_7776);
xnor U8406 (N_8406,N_7726,N_7545);
xor U8407 (N_8407,N_7737,N_7874);
or U8408 (N_8408,N_7664,N_7740);
nand U8409 (N_8409,N_7942,N_7697);
and U8410 (N_8410,N_7752,N_7751);
xnor U8411 (N_8411,N_7731,N_7571);
and U8412 (N_8412,N_7570,N_7833);
or U8413 (N_8413,N_7562,N_7506);
or U8414 (N_8414,N_7673,N_7935);
or U8415 (N_8415,N_7632,N_7748);
nand U8416 (N_8416,N_7734,N_7837);
and U8417 (N_8417,N_7972,N_7743);
or U8418 (N_8418,N_7664,N_7991);
nand U8419 (N_8419,N_7804,N_7976);
nand U8420 (N_8420,N_7741,N_7982);
or U8421 (N_8421,N_7515,N_7829);
and U8422 (N_8422,N_7608,N_7970);
or U8423 (N_8423,N_7765,N_7756);
nand U8424 (N_8424,N_7595,N_7896);
xor U8425 (N_8425,N_7612,N_7538);
and U8426 (N_8426,N_7596,N_7582);
and U8427 (N_8427,N_7785,N_7527);
or U8428 (N_8428,N_7693,N_7701);
nor U8429 (N_8429,N_7862,N_7771);
xor U8430 (N_8430,N_7615,N_7662);
nor U8431 (N_8431,N_7529,N_7749);
or U8432 (N_8432,N_7744,N_7854);
nor U8433 (N_8433,N_7738,N_7767);
and U8434 (N_8434,N_7631,N_7884);
nand U8435 (N_8435,N_7936,N_7536);
nand U8436 (N_8436,N_7824,N_7937);
nor U8437 (N_8437,N_7901,N_7970);
nand U8438 (N_8438,N_7576,N_7795);
or U8439 (N_8439,N_7763,N_7904);
or U8440 (N_8440,N_7694,N_7903);
xnor U8441 (N_8441,N_7859,N_7693);
nor U8442 (N_8442,N_7539,N_7835);
xnor U8443 (N_8443,N_7667,N_7836);
and U8444 (N_8444,N_7817,N_7646);
and U8445 (N_8445,N_7925,N_7779);
nand U8446 (N_8446,N_7883,N_7844);
and U8447 (N_8447,N_7745,N_7552);
nor U8448 (N_8448,N_7649,N_7751);
nand U8449 (N_8449,N_7771,N_7693);
or U8450 (N_8450,N_7560,N_7507);
or U8451 (N_8451,N_7601,N_7960);
nand U8452 (N_8452,N_7926,N_7590);
or U8453 (N_8453,N_7942,N_7887);
nand U8454 (N_8454,N_7680,N_7558);
and U8455 (N_8455,N_7771,N_7540);
or U8456 (N_8456,N_7827,N_7803);
xor U8457 (N_8457,N_7675,N_7744);
and U8458 (N_8458,N_7742,N_7697);
or U8459 (N_8459,N_7770,N_7668);
or U8460 (N_8460,N_7632,N_7890);
and U8461 (N_8461,N_7947,N_7571);
nor U8462 (N_8462,N_7749,N_7786);
and U8463 (N_8463,N_7543,N_7567);
nand U8464 (N_8464,N_7957,N_7998);
and U8465 (N_8465,N_7588,N_7760);
nor U8466 (N_8466,N_7628,N_7784);
and U8467 (N_8467,N_7986,N_7700);
nand U8468 (N_8468,N_7566,N_7721);
nor U8469 (N_8469,N_7554,N_7933);
xor U8470 (N_8470,N_7884,N_7526);
xnor U8471 (N_8471,N_7827,N_7968);
and U8472 (N_8472,N_7507,N_7953);
or U8473 (N_8473,N_7861,N_7641);
xor U8474 (N_8474,N_7950,N_7842);
nand U8475 (N_8475,N_7847,N_7566);
nor U8476 (N_8476,N_7916,N_7561);
or U8477 (N_8477,N_7830,N_7727);
nor U8478 (N_8478,N_7582,N_7844);
nand U8479 (N_8479,N_7515,N_7633);
nand U8480 (N_8480,N_7749,N_7952);
xor U8481 (N_8481,N_7749,N_7930);
nand U8482 (N_8482,N_7735,N_7669);
xor U8483 (N_8483,N_7684,N_7567);
xnor U8484 (N_8484,N_7776,N_7986);
or U8485 (N_8485,N_7710,N_7759);
xnor U8486 (N_8486,N_7562,N_7655);
xor U8487 (N_8487,N_7545,N_7647);
xnor U8488 (N_8488,N_7887,N_7897);
and U8489 (N_8489,N_7786,N_7545);
and U8490 (N_8490,N_7594,N_7996);
nor U8491 (N_8491,N_7806,N_7924);
nor U8492 (N_8492,N_7996,N_7599);
and U8493 (N_8493,N_7512,N_7948);
nor U8494 (N_8494,N_7573,N_7508);
and U8495 (N_8495,N_7595,N_7810);
and U8496 (N_8496,N_7934,N_7817);
nor U8497 (N_8497,N_7936,N_7786);
xor U8498 (N_8498,N_7792,N_7705);
nor U8499 (N_8499,N_7699,N_7979);
or U8500 (N_8500,N_8048,N_8389);
and U8501 (N_8501,N_8449,N_8386);
nor U8502 (N_8502,N_8353,N_8152);
nand U8503 (N_8503,N_8246,N_8422);
and U8504 (N_8504,N_8354,N_8089);
nor U8505 (N_8505,N_8226,N_8129);
and U8506 (N_8506,N_8049,N_8034);
xor U8507 (N_8507,N_8312,N_8085);
and U8508 (N_8508,N_8088,N_8341);
xor U8509 (N_8509,N_8496,N_8280);
nor U8510 (N_8510,N_8397,N_8402);
xor U8511 (N_8511,N_8008,N_8004);
and U8512 (N_8512,N_8398,N_8027);
or U8513 (N_8513,N_8487,N_8388);
xnor U8514 (N_8514,N_8207,N_8335);
xnor U8515 (N_8515,N_8407,N_8482);
nand U8516 (N_8516,N_8208,N_8116);
or U8517 (N_8517,N_8118,N_8411);
xor U8518 (N_8518,N_8431,N_8159);
nand U8519 (N_8519,N_8454,N_8416);
nand U8520 (N_8520,N_8275,N_8426);
and U8521 (N_8521,N_8236,N_8241);
nand U8522 (N_8522,N_8419,N_8443);
nand U8523 (N_8523,N_8425,N_8459);
nor U8524 (N_8524,N_8465,N_8289);
or U8525 (N_8525,N_8286,N_8003);
nand U8526 (N_8526,N_8175,N_8051);
xnor U8527 (N_8527,N_8259,N_8043);
nor U8528 (N_8528,N_8359,N_8342);
xor U8529 (N_8529,N_8221,N_8038);
xnor U8530 (N_8530,N_8072,N_8379);
nor U8531 (N_8531,N_8460,N_8127);
or U8532 (N_8532,N_8110,N_8257);
nand U8533 (N_8533,N_8172,N_8084);
nand U8534 (N_8534,N_8391,N_8151);
nor U8535 (N_8535,N_8028,N_8093);
nor U8536 (N_8536,N_8390,N_8392);
nor U8537 (N_8537,N_8115,N_8166);
and U8538 (N_8538,N_8000,N_8169);
and U8539 (N_8539,N_8213,N_8047);
xnor U8540 (N_8540,N_8483,N_8440);
nor U8541 (N_8541,N_8070,N_8373);
or U8542 (N_8542,N_8247,N_8130);
or U8543 (N_8543,N_8446,N_8382);
nand U8544 (N_8544,N_8202,N_8396);
and U8545 (N_8545,N_8380,N_8098);
or U8546 (N_8546,N_8090,N_8451);
and U8547 (N_8547,N_8385,N_8320);
and U8548 (N_8548,N_8481,N_8078);
or U8549 (N_8549,N_8077,N_8435);
nand U8550 (N_8550,N_8405,N_8186);
xor U8551 (N_8551,N_8351,N_8020);
or U8552 (N_8552,N_8306,N_8105);
nor U8553 (N_8553,N_8216,N_8310);
xnor U8554 (N_8554,N_8432,N_8137);
or U8555 (N_8555,N_8498,N_8173);
and U8556 (N_8556,N_8233,N_8288);
xnor U8557 (N_8557,N_8472,N_8430);
nand U8558 (N_8558,N_8346,N_8434);
nor U8559 (N_8559,N_8318,N_8324);
xor U8560 (N_8560,N_8201,N_8160);
nor U8561 (N_8561,N_8150,N_8271);
and U8562 (N_8562,N_8058,N_8319);
and U8563 (N_8563,N_8339,N_8067);
and U8564 (N_8564,N_8330,N_8184);
or U8565 (N_8565,N_8229,N_8326);
nor U8566 (N_8566,N_8249,N_8138);
xor U8567 (N_8567,N_8122,N_8064);
nor U8568 (N_8568,N_8193,N_8300);
xnor U8569 (N_8569,N_8337,N_8283);
xnor U8570 (N_8570,N_8479,N_8444);
xor U8571 (N_8571,N_8071,N_8418);
xor U8572 (N_8572,N_8204,N_8083);
nor U8573 (N_8573,N_8304,N_8139);
nand U8574 (N_8574,N_8448,N_8189);
nor U8575 (N_8575,N_8102,N_8096);
xnor U8576 (N_8576,N_8023,N_8142);
xor U8577 (N_8577,N_8367,N_8113);
nand U8578 (N_8578,N_8101,N_8143);
and U8579 (N_8579,N_8366,N_8250);
nor U8580 (N_8580,N_8106,N_8258);
nor U8581 (N_8581,N_8290,N_8269);
or U8582 (N_8582,N_8183,N_8327);
xor U8583 (N_8583,N_8458,N_8270);
nand U8584 (N_8584,N_8281,N_8291);
or U8585 (N_8585,N_8156,N_8042);
and U8586 (N_8586,N_8178,N_8420);
xor U8587 (N_8587,N_8220,N_8225);
nor U8588 (N_8588,N_8117,N_8181);
or U8589 (N_8589,N_8428,N_8447);
xnor U8590 (N_8590,N_8006,N_8120);
or U8591 (N_8591,N_8413,N_8403);
and U8592 (N_8592,N_8494,N_8365);
nor U8593 (N_8593,N_8211,N_8153);
xnor U8594 (N_8594,N_8490,N_8414);
and U8595 (N_8595,N_8338,N_8358);
and U8596 (N_8596,N_8171,N_8329);
or U8597 (N_8597,N_8344,N_8296);
nand U8598 (N_8598,N_8148,N_8356);
or U8599 (N_8599,N_8182,N_8266);
nand U8600 (N_8600,N_8328,N_8360);
xnor U8601 (N_8601,N_8141,N_8161);
or U8602 (N_8602,N_8384,N_8316);
nand U8603 (N_8603,N_8194,N_8378);
nor U8604 (N_8604,N_8303,N_8033);
xor U8605 (N_8605,N_8251,N_8230);
xor U8606 (N_8606,N_8239,N_8214);
xor U8607 (N_8607,N_8493,N_8484);
nand U8608 (N_8608,N_8375,N_8215);
nor U8609 (N_8609,N_8469,N_8167);
nor U8610 (N_8610,N_8073,N_8144);
nand U8611 (N_8611,N_8024,N_8199);
xnor U8612 (N_8612,N_8170,N_8321);
xor U8613 (N_8613,N_8491,N_8188);
and U8614 (N_8614,N_8069,N_8471);
xor U8615 (N_8615,N_8054,N_8134);
or U8616 (N_8616,N_8046,N_8087);
nand U8617 (N_8617,N_8442,N_8001);
or U8618 (N_8618,N_8252,N_8376);
nand U8619 (N_8619,N_8061,N_8383);
or U8620 (N_8620,N_8499,N_8017);
or U8621 (N_8621,N_8176,N_8313);
or U8622 (N_8622,N_8273,N_8347);
xnor U8623 (N_8623,N_8010,N_8438);
or U8624 (N_8624,N_8298,N_8021);
xor U8625 (N_8625,N_8417,N_8475);
xnor U8626 (N_8626,N_8415,N_8371);
nor U8627 (N_8627,N_8470,N_8157);
xnor U8628 (N_8628,N_8031,N_8197);
nor U8629 (N_8629,N_8045,N_8466);
xnor U8630 (N_8630,N_8268,N_8095);
nor U8631 (N_8631,N_8334,N_8336);
xor U8632 (N_8632,N_8149,N_8164);
nor U8633 (N_8633,N_8489,N_8456);
and U8634 (N_8634,N_8076,N_8155);
and U8635 (N_8635,N_8002,N_8133);
nand U8636 (N_8636,N_8112,N_8315);
nand U8637 (N_8637,N_8492,N_8476);
xnor U8638 (N_8638,N_8497,N_8185);
nand U8639 (N_8639,N_8399,N_8349);
or U8640 (N_8640,N_8158,N_8311);
or U8641 (N_8641,N_8372,N_8192);
nor U8642 (N_8642,N_8111,N_8488);
or U8643 (N_8643,N_8212,N_8473);
nand U8644 (N_8644,N_8114,N_8410);
nor U8645 (N_8645,N_8195,N_8040);
and U8646 (N_8646,N_8007,N_8361);
and U8647 (N_8647,N_8009,N_8092);
nor U8648 (N_8648,N_8323,N_8474);
nor U8649 (N_8649,N_8041,N_8053);
or U8650 (N_8650,N_8065,N_8278);
nor U8651 (N_8651,N_8455,N_8218);
nand U8652 (N_8652,N_8277,N_8074);
and U8653 (N_8653,N_8132,N_8025);
nand U8654 (N_8654,N_8191,N_8299);
nand U8655 (N_8655,N_8343,N_8265);
or U8656 (N_8656,N_8394,N_8154);
xor U8657 (N_8657,N_8279,N_8421);
nand U8658 (N_8658,N_8307,N_8174);
and U8659 (N_8659,N_8301,N_8068);
nand U8660 (N_8660,N_8357,N_8210);
or U8661 (N_8661,N_8467,N_8352);
and U8662 (N_8662,N_8284,N_8203);
xor U8663 (N_8663,N_8036,N_8267);
and U8664 (N_8664,N_8406,N_8099);
xnor U8665 (N_8665,N_8468,N_8231);
and U8666 (N_8666,N_8457,N_8295);
xnor U8667 (N_8667,N_8039,N_8103);
or U8668 (N_8668,N_8285,N_8245);
and U8669 (N_8669,N_8136,N_8276);
nand U8670 (N_8670,N_8350,N_8264);
nand U8671 (N_8671,N_8005,N_8395);
nand U8672 (N_8672,N_8332,N_8260);
and U8673 (N_8673,N_8056,N_8445);
and U8674 (N_8674,N_8362,N_8486);
nand U8675 (N_8675,N_8016,N_8128);
nand U8676 (N_8676,N_8363,N_8125);
nand U8677 (N_8677,N_8165,N_8228);
or U8678 (N_8678,N_8223,N_8082);
xnor U8679 (N_8679,N_8035,N_8075);
xnor U8680 (N_8680,N_8248,N_8044);
nor U8681 (N_8681,N_8408,N_8393);
nor U8682 (N_8682,N_8333,N_8062);
or U8683 (N_8683,N_8119,N_8109);
xnor U8684 (N_8684,N_8253,N_8294);
and U8685 (N_8685,N_8305,N_8091);
nor U8686 (N_8686,N_8209,N_8377);
xor U8687 (N_8687,N_8108,N_8495);
xnor U8688 (N_8688,N_8453,N_8463);
xor U8689 (N_8689,N_8345,N_8217);
or U8690 (N_8690,N_8196,N_8135);
nand U8691 (N_8691,N_8079,N_8029);
or U8692 (N_8692,N_8477,N_8055);
nor U8693 (N_8693,N_8274,N_8317);
nand U8694 (N_8694,N_8013,N_8019);
nor U8695 (N_8695,N_8187,N_8050);
xnor U8696 (N_8696,N_8374,N_8439);
nand U8697 (N_8697,N_8032,N_8409);
and U8698 (N_8698,N_8063,N_8145);
and U8699 (N_8699,N_8429,N_8424);
and U8700 (N_8700,N_8401,N_8018);
or U8701 (N_8701,N_8126,N_8404);
or U8702 (N_8702,N_8146,N_8011);
or U8703 (N_8703,N_8370,N_8427);
xor U8704 (N_8704,N_8180,N_8355);
xor U8705 (N_8705,N_8292,N_8433);
nor U8706 (N_8706,N_8309,N_8066);
xnor U8707 (N_8707,N_8256,N_8314);
xor U8708 (N_8708,N_8014,N_8400);
and U8709 (N_8709,N_8081,N_8302);
and U8710 (N_8710,N_8255,N_8121);
xor U8711 (N_8711,N_8205,N_8412);
and U8712 (N_8712,N_8262,N_8124);
xnor U8713 (N_8713,N_8094,N_8147);
or U8714 (N_8714,N_8308,N_8131);
nor U8715 (N_8715,N_8190,N_8198);
or U8716 (N_8716,N_8026,N_8261);
or U8717 (N_8717,N_8348,N_8107);
and U8718 (N_8718,N_8387,N_8086);
and U8719 (N_8719,N_8297,N_8104);
nand U8720 (N_8720,N_8224,N_8200);
nand U8721 (N_8721,N_8238,N_8485);
nand U8722 (N_8722,N_8462,N_8162);
and U8723 (N_8723,N_8480,N_8461);
nor U8724 (N_8724,N_8037,N_8287);
nand U8725 (N_8725,N_8022,N_8464);
and U8726 (N_8726,N_8234,N_8293);
nand U8727 (N_8727,N_8254,N_8015);
nor U8728 (N_8728,N_8282,N_8235);
xor U8729 (N_8729,N_8206,N_8059);
xnor U8730 (N_8730,N_8097,N_8478);
or U8731 (N_8731,N_8060,N_8237);
nor U8732 (N_8732,N_8242,N_8423);
xnor U8733 (N_8733,N_8140,N_8177);
nor U8734 (N_8734,N_8368,N_8437);
and U8735 (N_8735,N_8325,N_8179);
xnor U8736 (N_8736,N_8222,N_8244);
xor U8737 (N_8737,N_8452,N_8052);
nand U8738 (N_8738,N_8100,N_8163);
xor U8739 (N_8739,N_8369,N_8168);
nand U8740 (N_8740,N_8080,N_8450);
xnor U8741 (N_8741,N_8436,N_8331);
or U8742 (N_8742,N_8030,N_8272);
nand U8743 (N_8743,N_8263,N_8340);
nand U8744 (N_8744,N_8322,N_8012);
nand U8745 (N_8745,N_8232,N_8057);
or U8746 (N_8746,N_8227,N_8240);
nand U8747 (N_8747,N_8381,N_8219);
or U8748 (N_8748,N_8364,N_8123);
nor U8749 (N_8749,N_8243,N_8441);
or U8750 (N_8750,N_8296,N_8077);
nand U8751 (N_8751,N_8064,N_8489);
or U8752 (N_8752,N_8402,N_8312);
nor U8753 (N_8753,N_8000,N_8024);
xor U8754 (N_8754,N_8367,N_8478);
or U8755 (N_8755,N_8480,N_8089);
xnor U8756 (N_8756,N_8069,N_8473);
nor U8757 (N_8757,N_8410,N_8238);
and U8758 (N_8758,N_8079,N_8485);
xor U8759 (N_8759,N_8063,N_8111);
and U8760 (N_8760,N_8045,N_8088);
and U8761 (N_8761,N_8276,N_8342);
and U8762 (N_8762,N_8137,N_8128);
or U8763 (N_8763,N_8230,N_8133);
or U8764 (N_8764,N_8101,N_8394);
nor U8765 (N_8765,N_8499,N_8189);
nand U8766 (N_8766,N_8482,N_8365);
or U8767 (N_8767,N_8171,N_8266);
nand U8768 (N_8768,N_8267,N_8488);
or U8769 (N_8769,N_8298,N_8059);
xor U8770 (N_8770,N_8410,N_8443);
xor U8771 (N_8771,N_8379,N_8094);
nor U8772 (N_8772,N_8111,N_8359);
nand U8773 (N_8773,N_8208,N_8344);
nand U8774 (N_8774,N_8108,N_8282);
or U8775 (N_8775,N_8227,N_8061);
nor U8776 (N_8776,N_8208,N_8052);
nand U8777 (N_8777,N_8392,N_8288);
nor U8778 (N_8778,N_8285,N_8132);
and U8779 (N_8779,N_8228,N_8367);
or U8780 (N_8780,N_8138,N_8300);
nor U8781 (N_8781,N_8115,N_8331);
xor U8782 (N_8782,N_8079,N_8420);
or U8783 (N_8783,N_8356,N_8073);
nor U8784 (N_8784,N_8232,N_8074);
and U8785 (N_8785,N_8130,N_8210);
nor U8786 (N_8786,N_8335,N_8465);
or U8787 (N_8787,N_8494,N_8216);
nor U8788 (N_8788,N_8275,N_8451);
nand U8789 (N_8789,N_8417,N_8186);
or U8790 (N_8790,N_8195,N_8416);
xor U8791 (N_8791,N_8019,N_8353);
nor U8792 (N_8792,N_8441,N_8453);
nor U8793 (N_8793,N_8163,N_8187);
nand U8794 (N_8794,N_8153,N_8464);
and U8795 (N_8795,N_8346,N_8348);
nor U8796 (N_8796,N_8000,N_8479);
nand U8797 (N_8797,N_8359,N_8117);
or U8798 (N_8798,N_8379,N_8131);
xor U8799 (N_8799,N_8177,N_8042);
nand U8800 (N_8800,N_8176,N_8264);
nand U8801 (N_8801,N_8365,N_8206);
nor U8802 (N_8802,N_8248,N_8128);
or U8803 (N_8803,N_8113,N_8305);
nor U8804 (N_8804,N_8425,N_8298);
and U8805 (N_8805,N_8335,N_8048);
nand U8806 (N_8806,N_8182,N_8367);
nand U8807 (N_8807,N_8059,N_8427);
nor U8808 (N_8808,N_8070,N_8065);
or U8809 (N_8809,N_8481,N_8205);
nor U8810 (N_8810,N_8078,N_8144);
nor U8811 (N_8811,N_8172,N_8026);
nand U8812 (N_8812,N_8342,N_8466);
and U8813 (N_8813,N_8072,N_8358);
and U8814 (N_8814,N_8379,N_8431);
nor U8815 (N_8815,N_8346,N_8444);
and U8816 (N_8816,N_8065,N_8129);
nand U8817 (N_8817,N_8320,N_8116);
xnor U8818 (N_8818,N_8145,N_8262);
or U8819 (N_8819,N_8018,N_8213);
or U8820 (N_8820,N_8492,N_8483);
nand U8821 (N_8821,N_8369,N_8062);
or U8822 (N_8822,N_8370,N_8342);
or U8823 (N_8823,N_8474,N_8387);
or U8824 (N_8824,N_8304,N_8189);
nor U8825 (N_8825,N_8044,N_8107);
nand U8826 (N_8826,N_8426,N_8064);
xor U8827 (N_8827,N_8476,N_8302);
or U8828 (N_8828,N_8227,N_8347);
or U8829 (N_8829,N_8321,N_8184);
xnor U8830 (N_8830,N_8026,N_8478);
and U8831 (N_8831,N_8367,N_8063);
nand U8832 (N_8832,N_8099,N_8428);
xor U8833 (N_8833,N_8009,N_8447);
and U8834 (N_8834,N_8055,N_8483);
or U8835 (N_8835,N_8136,N_8449);
nor U8836 (N_8836,N_8372,N_8096);
nand U8837 (N_8837,N_8180,N_8261);
xnor U8838 (N_8838,N_8288,N_8413);
nand U8839 (N_8839,N_8134,N_8156);
xor U8840 (N_8840,N_8378,N_8331);
nor U8841 (N_8841,N_8469,N_8339);
or U8842 (N_8842,N_8101,N_8161);
and U8843 (N_8843,N_8212,N_8475);
xnor U8844 (N_8844,N_8001,N_8030);
xor U8845 (N_8845,N_8048,N_8180);
xor U8846 (N_8846,N_8414,N_8282);
nand U8847 (N_8847,N_8139,N_8275);
or U8848 (N_8848,N_8011,N_8033);
nor U8849 (N_8849,N_8472,N_8041);
or U8850 (N_8850,N_8311,N_8204);
xor U8851 (N_8851,N_8050,N_8002);
nor U8852 (N_8852,N_8262,N_8032);
and U8853 (N_8853,N_8315,N_8182);
or U8854 (N_8854,N_8073,N_8440);
or U8855 (N_8855,N_8062,N_8430);
and U8856 (N_8856,N_8002,N_8413);
or U8857 (N_8857,N_8072,N_8261);
nor U8858 (N_8858,N_8303,N_8055);
and U8859 (N_8859,N_8488,N_8197);
xnor U8860 (N_8860,N_8416,N_8363);
nand U8861 (N_8861,N_8453,N_8246);
nand U8862 (N_8862,N_8022,N_8450);
nor U8863 (N_8863,N_8394,N_8239);
nand U8864 (N_8864,N_8025,N_8137);
nor U8865 (N_8865,N_8089,N_8466);
nand U8866 (N_8866,N_8328,N_8303);
xor U8867 (N_8867,N_8125,N_8194);
nor U8868 (N_8868,N_8095,N_8367);
and U8869 (N_8869,N_8391,N_8023);
xnor U8870 (N_8870,N_8017,N_8431);
or U8871 (N_8871,N_8247,N_8216);
or U8872 (N_8872,N_8486,N_8431);
nor U8873 (N_8873,N_8350,N_8303);
nand U8874 (N_8874,N_8224,N_8033);
nand U8875 (N_8875,N_8427,N_8317);
and U8876 (N_8876,N_8242,N_8324);
and U8877 (N_8877,N_8100,N_8212);
or U8878 (N_8878,N_8140,N_8244);
nand U8879 (N_8879,N_8481,N_8076);
or U8880 (N_8880,N_8025,N_8475);
xnor U8881 (N_8881,N_8167,N_8121);
or U8882 (N_8882,N_8144,N_8306);
xnor U8883 (N_8883,N_8467,N_8368);
nor U8884 (N_8884,N_8303,N_8480);
xnor U8885 (N_8885,N_8174,N_8232);
nand U8886 (N_8886,N_8495,N_8107);
xnor U8887 (N_8887,N_8253,N_8068);
nor U8888 (N_8888,N_8339,N_8014);
or U8889 (N_8889,N_8433,N_8204);
nor U8890 (N_8890,N_8086,N_8379);
or U8891 (N_8891,N_8178,N_8045);
nand U8892 (N_8892,N_8399,N_8385);
nor U8893 (N_8893,N_8439,N_8271);
nand U8894 (N_8894,N_8401,N_8293);
or U8895 (N_8895,N_8179,N_8053);
or U8896 (N_8896,N_8265,N_8162);
xnor U8897 (N_8897,N_8488,N_8057);
nand U8898 (N_8898,N_8328,N_8411);
xor U8899 (N_8899,N_8474,N_8245);
nand U8900 (N_8900,N_8092,N_8135);
xnor U8901 (N_8901,N_8241,N_8069);
nor U8902 (N_8902,N_8135,N_8189);
or U8903 (N_8903,N_8451,N_8260);
nand U8904 (N_8904,N_8199,N_8209);
xnor U8905 (N_8905,N_8438,N_8298);
or U8906 (N_8906,N_8001,N_8325);
xor U8907 (N_8907,N_8133,N_8366);
and U8908 (N_8908,N_8097,N_8222);
nor U8909 (N_8909,N_8465,N_8405);
and U8910 (N_8910,N_8402,N_8334);
nor U8911 (N_8911,N_8146,N_8323);
and U8912 (N_8912,N_8370,N_8275);
nand U8913 (N_8913,N_8340,N_8146);
and U8914 (N_8914,N_8340,N_8431);
nand U8915 (N_8915,N_8314,N_8254);
and U8916 (N_8916,N_8300,N_8436);
nor U8917 (N_8917,N_8405,N_8309);
xnor U8918 (N_8918,N_8059,N_8333);
nor U8919 (N_8919,N_8394,N_8017);
and U8920 (N_8920,N_8037,N_8014);
nor U8921 (N_8921,N_8166,N_8146);
or U8922 (N_8922,N_8266,N_8141);
nor U8923 (N_8923,N_8242,N_8202);
and U8924 (N_8924,N_8411,N_8060);
or U8925 (N_8925,N_8063,N_8169);
and U8926 (N_8926,N_8344,N_8348);
and U8927 (N_8927,N_8412,N_8467);
nand U8928 (N_8928,N_8196,N_8349);
or U8929 (N_8929,N_8164,N_8301);
nand U8930 (N_8930,N_8202,N_8162);
or U8931 (N_8931,N_8439,N_8137);
nand U8932 (N_8932,N_8283,N_8288);
nor U8933 (N_8933,N_8015,N_8491);
nand U8934 (N_8934,N_8442,N_8338);
or U8935 (N_8935,N_8313,N_8478);
and U8936 (N_8936,N_8034,N_8349);
nor U8937 (N_8937,N_8030,N_8239);
or U8938 (N_8938,N_8476,N_8093);
nand U8939 (N_8939,N_8036,N_8020);
xor U8940 (N_8940,N_8233,N_8392);
nor U8941 (N_8941,N_8144,N_8131);
xnor U8942 (N_8942,N_8002,N_8108);
nor U8943 (N_8943,N_8326,N_8081);
xor U8944 (N_8944,N_8127,N_8105);
or U8945 (N_8945,N_8230,N_8073);
nor U8946 (N_8946,N_8174,N_8435);
nor U8947 (N_8947,N_8228,N_8010);
or U8948 (N_8948,N_8476,N_8382);
xnor U8949 (N_8949,N_8138,N_8471);
or U8950 (N_8950,N_8418,N_8368);
or U8951 (N_8951,N_8057,N_8318);
nand U8952 (N_8952,N_8226,N_8014);
or U8953 (N_8953,N_8368,N_8133);
xor U8954 (N_8954,N_8259,N_8422);
and U8955 (N_8955,N_8385,N_8137);
or U8956 (N_8956,N_8203,N_8155);
nor U8957 (N_8957,N_8271,N_8112);
nor U8958 (N_8958,N_8353,N_8369);
or U8959 (N_8959,N_8177,N_8394);
nor U8960 (N_8960,N_8194,N_8401);
xor U8961 (N_8961,N_8130,N_8399);
nand U8962 (N_8962,N_8277,N_8423);
nand U8963 (N_8963,N_8017,N_8190);
nor U8964 (N_8964,N_8157,N_8015);
and U8965 (N_8965,N_8406,N_8449);
or U8966 (N_8966,N_8137,N_8323);
xor U8967 (N_8967,N_8396,N_8220);
and U8968 (N_8968,N_8341,N_8371);
and U8969 (N_8969,N_8217,N_8254);
nand U8970 (N_8970,N_8191,N_8232);
and U8971 (N_8971,N_8121,N_8086);
nor U8972 (N_8972,N_8318,N_8308);
and U8973 (N_8973,N_8471,N_8290);
xor U8974 (N_8974,N_8432,N_8039);
xor U8975 (N_8975,N_8411,N_8061);
or U8976 (N_8976,N_8125,N_8460);
and U8977 (N_8977,N_8464,N_8236);
or U8978 (N_8978,N_8185,N_8180);
xor U8979 (N_8979,N_8342,N_8255);
nor U8980 (N_8980,N_8126,N_8253);
xnor U8981 (N_8981,N_8095,N_8048);
and U8982 (N_8982,N_8364,N_8098);
or U8983 (N_8983,N_8102,N_8375);
nand U8984 (N_8984,N_8042,N_8237);
xor U8985 (N_8985,N_8297,N_8429);
xor U8986 (N_8986,N_8309,N_8198);
and U8987 (N_8987,N_8120,N_8362);
xnor U8988 (N_8988,N_8388,N_8299);
nor U8989 (N_8989,N_8257,N_8240);
and U8990 (N_8990,N_8407,N_8287);
nor U8991 (N_8991,N_8086,N_8188);
xnor U8992 (N_8992,N_8212,N_8370);
and U8993 (N_8993,N_8249,N_8345);
xor U8994 (N_8994,N_8341,N_8089);
or U8995 (N_8995,N_8134,N_8378);
and U8996 (N_8996,N_8043,N_8263);
xnor U8997 (N_8997,N_8429,N_8323);
and U8998 (N_8998,N_8349,N_8047);
or U8999 (N_8999,N_8347,N_8358);
or U9000 (N_9000,N_8979,N_8618);
nand U9001 (N_9001,N_8691,N_8938);
nor U9002 (N_9002,N_8789,N_8993);
nor U9003 (N_9003,N_8505,N_8779);
and U9004 (N_9004,N_8630,N_8797);
nor U9005 (N_9005,N_8626,N_8513);
and U9006 (N_9006,N_8893,N_8917);
and U9007 (N_9007,N_8560,N_8610);
and U9008 (N_9008,N_8621,N_8906);
nor U9009 (N_9009,N_8943,N_8780);
or U9010 (N_9010,N_8972,N_8937);
nor U9011 (N_9011,N_8619,N_8720);
xnor U9012 (N_9012,N_8654,N_8996);
xnor U9013 (N_9013,N_8612,N_8567);
or U9014 (N_9014,N_8553,N_8737);
nand U9015 (N_9015,N_8948,N_8601);
nor U9016 (N_9016,N_8705,N_8859);
or U9017 (N_9017,N_8604,N_8650);
nor U9018 (N_9018,N_8633,N_8933);
or U9019 (N_9019,N_8734,N_8540);
nand U9020 (N_9020,N_8754,N_8947);
or U9021 (N_9021,N_8594,N_8827);
nand U9022 (N_9022,N_8868,N_8985);
nor U9023 (N_9023,N_8945,N_8728);
nand U9024 (N_9024,N_8932,N_8561);
and U9025 (N_9025,N_8642,N_8687);
or U9026 (N_9026,N_8834,N_8558);
and U9027 (N_9027,N_8711,N_8964);
xor U9028 (N_9028,N_8719,N_8651);
xnor U9029 (N_9029,N_8989,N_8586);
and U9030 (N_9030,N_8925,N_8915);
xor U9031 (N_9031,N_8931,N_8628);
xnor U9032 (N_9032,N_8702,N_8710);
and U9033 (N_9033,N_8544,N_8795);
and U9034 (N_9034,N_8950,N_8721);
or U9035 (N_9035,N_8579,N_8872);
xor U9036 (N_9036,N_8584,N_8799);
or U9037 (N_9037,N_8707,N_8590);
or U9038 (N_9038,N_8631,N_8848);
or U9039 (N_9039,N_8507,N_8758);
or U9040 (N_9040,N_8747,N_8693);
xnor U9041 (N_9041,N_8546,N_8967);
xor U9042 (N_9042,N_8879,N_8767);
nor U9043 (N_9043,N_8823,N_8955);
nand U9044 (N_9044,N_8919,N_8547);
xnor U9045 (N_9045,N_8537,N_8713);
xor U9046 (N_9046,N_8817,N_8966);
xnor U9047 (N_9047,N_8785,N_8965);
nor U9048 (N_9048,N_8697,N_8974);
xor U9049 (N_9049,N_8674,N_8733);
and U9050 (N_9050,N_8929,N_8946);
or U9051 (N_9051,N_8995,N_8752);
or U9052 (N_9052,N_8842,N_8942);
and U9053 (N_9053,N_8577,N_8895);
xnor U9054 (N_9054,N_8746,N_8531);
nand U9055 (N_9055,N_8908,N_8769);
nand U9056 (N_9056,N_8690,N_8638);
nor U9057 (N_9057,N_8539,N_8564);
and U9058 (N_9058,N_8784,N_8506);
nand U9059 (N_9059,N_8944,N_8936);
nor U9060 (N_9060,N_8732,N_8835);
nor U9061 (N_9061,N_8562,N_8639);
nand U9062 (N_9062,N_8583,N_8788);
nor U9063 (N_9063,N_8951,N_8910);
or U9064 (N_9064,N_8682,N_8962);
xor U9065 (N_9065,N_8881,N_8837);
or U9066 (N_9066,N_8865,N_8658);
nand U9067 (N_9067,N_8709,N_8692);
and U9068 (N_9068,N_8724,N_8749);
and U9069 (N_9069,N_8646,N_8649);
nor U9070 (N_9070,N_8609,N_8627);
and U9071 (N_9071,N_8880,N_8864);
nand U9072 (N_9072,N_8502,N_8600);
and U9073 (N_9073,N_8636,N_8524);
nor U9074 (N_9074,N_8635,N_8884);
nand U9075 (N_9075,N_8998,N_8886);
or U9076 (N_9076,N_8503,N_8681);
nand U9077 (N_9077,N_8653,N_8568);
and U9078 (N_9078,N_8751,N_8529);
or U9079 (N_9079,N_8829,N_8555);
or U9080 (N_9080,N_8963,N_8850);
nor U9081 (N_9081,N_8602,N_8914);
and U9082 (N_9082,N_8822,N_8866);
nor U9083 (N_9083,N_8666,N_8888);
nor U9084 (N_9084,N_8997,N_8510);
nand U9085 (N_9085,N_8640,N_8695);
nand U9086 (N_9086,N_8934,N_8545);
nor U9087 (N_9087,N_8718,N_8870);
xor U9088 (N_9088,N_8987,N_8836);
nor U9089 (N_9089,N_8740,N_8973);
xor U9090 (N_9090,N_8607,N_8615);
xor U9091 (N_9091,N_8620,N_8844);
nand U9092 (N_9092,N_8890,N_8912);
nand U9093 (N_9093,N_8854,N_8731);
nor U9094 (N_9094,N_8899,N_8730);
or U9095 (N_9095,N_8833,N_8891);
or U9096 (N_9096,N_8556,N_8768);
xor U9097 (N_9097,N_8552,N_8701);
xor U9098 (N_9098,N_8875,N_8782);
and U9099 (N_9099,N_8971,N_8764);
xnor U9100 (N_9100,N_8957,N_8675);
or U9101 (N_9101,N_8725,N_8763);
or U9102 (N_9102,N_8592,N_8885);
nand U9103 (N_9103,N_8559,N_8887);
and U9104 (N_9104,N_8841,N_8664);
nor U9105 (N_9105,N_8909,N_8988);
or U9106 (N_9106,N_8533,N_8500);
or U9107 (N_9107,N_8663,N_8598);
nand U9108 (N_9108,N_8597,N_8519);
nand U9109 (N_9109,N_8786,N_8976);
and U9110 (N_9110,N_8516,N_8977);
xor U9111 (N_9111,N_8678,N_8569);
xor U9112 (N_9112,N_8566,N_8548);
nor U9113 (N_9113,N_8831,N_8698);
or U9114 (N_9114,N_8905,N_8657);
nor U9115 (N_9115,N_8755,N_8587);
or U9116 (N_9116,N_8637,N_8862);
or U9117 (N_9117,N_8750,N_8696);
or U9118 (N_9118,N_8742,N_8603);
and U9119 (N_9119,N_8729,N_8515);
nand U9120 (N_9120,N_8816,N_8745);
xor U9121 (N_9121,N_8846,N_8794);
nand U9122 (N_9122,N_8813,N_8765);
xnor U9123 (N_9123,N_8787,N_8916);
nand U9124 (N_9124,N_8853,N_8595);
and U9125 (N_9125,N_8680,N_8772);
nand U9126 (N_9126,N_8699,N_8645);
nand U9127 (N_9127,N_8832,N_8800);
or U9128 (N_9128,N_8775,N_8588);
or U9129 (N_9129,N_8700,N_8857);
and U9130 (N_9130,N_8542,N_8551);
nand U9131 (N_9131,N_8806,N_8792);
and U9132 (N_9132,N_8736,N_8528);
nand U9133 (N_9133,N_8670,N_8926);
or U9134 (N_9134,N_8928,N_8903);
xor U9135 (N_9135,N_8541,N_8994);
xnor U9136 (N_9136,N_8571,N_8756);
or U9137 (N_9137,N_8543,N_8669);
or U9138 (N_9138,N_8830,N_8953);
xor U9139 (N_9139,N_8982,N_8520);
xnor U9140 (N_9140,N_8530,N_8992);
and U9141 (N_9141,N_8793,N_8554);
nor U9142 (N_9142,N_8574,N_8770);
or U9143 (N_9143,N_8525,N_8518);
or U9144 (N_9144,N_8739,N_8694);
xnor U9145 (N_9145,N_8757,N_8999);
xor U9146 (N_9146,N_8802,N_8907);
nor U9147 (N_9147,N_8759,N_8796);
and U9148 (N_9148,N_8761,N_8815);
or U9149 (N_9149,N_8743,N_8896);
nor U9150 (N_9150,N_8689,N_8686);
nor U9151 (N_9151,N_8660,N_8589);
and U9152 (N_9152,N_8673,N_8980);
nor U9153 (N_9153,N_8894,N_8825);
nand U9154 (N_9154,N_8573,N_8712);
nand U9155 (N_9155,N_8941,N_8869);
nand U9156 (N_9156,N_8593,N_8956);
and U9157 (N_9157,N_8504,N_8801);
and U9158 (N_9158,N_8617,N_8634);
or U9159 (N_9159,N_8521,N_8726);
or U9160 (N_9160,N_8762,N_8824);
xor U9161 (N_9161,N_8582,N_8852);
nor U9162 (N_9162,N_8684,N_8613);
nor U9163 (N_9163,N_8662,N_8969);
or U9164 (N_9164,N_8904,N_8549);
nor U9165 (N_9165,N_8706,N_8580);
xor U9166 (N_9166,N_8748,N_8652);
nor U9167 (N_9167,N_8523,N_8898);
xor U9168 (N_9168,N_8930,N_8803);
and U9169 (N_9169,N_8576,N_8808);
nand U9170 (N_9170,N_8984,N_8727);
xor U9171 (N_9171,N_8717,N_8809);
xor U9172 (N_9172,N_8897,N_8672);
and U9173 (N_9173,N_8778,N_8508);
nor U9174 (N_9174,N_8883,N_8991);
xnor U9175 (N_9175,N_8596,N_8623);
xor U9176 (N_9176,N_8585,N_8819);
or U9177 (N_9177,N_8921,N_8981);
nor U9178 (N_9178,N_8867,N_8661);
nor U9179 (N_9179,N_8954,N_8920);
nand U9180 (N_9180,N_8616,N_8856);
nand U9181 (N_9181,N_8847,N_8622);
nand U9182 (N_9182,N_8591,N_8771);
nor U9183 (N_9183,N_8723,N_8791);
xor U9184 (N_9184,N_8683,N_8961);
xnor U9185 (N_9185,N_8704,N_8629);
xor U9186 (N_9186,N_8714,N_8667);
and U9187 (N_9187,N_8860,N_8676);
or U9188 (N_9188,N_8889,N_8668);
xor U9189 (N_9189,N_8911,N_8685);
or U9190 (N_9190,N_8798,N_8570);
xnor U9191 (N_9191,N_8970,N_8708);
nand U9192 (N_9192,N_8876,N_8818);
and U9193 (N_9193,N_8838,N_8949);
and U9194 (N_9194,N_8608,N_8647);
xor U9195 (N_9195,N_8952,N_8820);
nor U9196 (N_9196,N_8783,N_8509);
or U9197 (N_9197,N_8812,N_8923);
nor U9198 (N_9198,N_8959,N_8536);
xor U9199 (N_9199,N_8858,N_8563);
nor U9200 (N_9200,N_8511,N_8871);
and U9201 (N_9201,N_8849,N_8804);
nor U9202 (N_9202,N_8679,N_8873);
or U9203 (N_9203,N_8656,N_8924);
xnor U9204 (N_9204,N_8703,N_8828);
or U9205 (N_9205,N_8927,N_8735);
nor U9206 (N_9206,N_8611,N_8773);
xor U9207 (N_9207,N_8760,N_8581);
xnor U9208 (N_9208,N_8643,N_8922);
and U9209 (N_9209,N_8538,N_8671);
xor U9210 (N_9210,N_8918,N_8781);
or U9211 (N_9211,N_8978,N_8665);
nand U9212 (N_9212,N_8632,N_8527);
nand U9213 (N_9213,N_8940,N_8776);
nand U9214 (N_9214,N_8526,N_8753);
nand U9215 (N_9215,N_8535,N_8655);
nand U9216 (N_9216,N_8902,N_8990);
nor U9217 (N_9217,N_8572,N_8624);
and U9218 (N_9218,N_8805,N_8741);
nand U9219 (N_9219,N_8715,N_8861);
and U9220 (N_9220,N_8968,N_8913);
nand U9221 (N_9221,N_8550,N_8565);
xor U9222 (N_9222,N_8557,N_8790);
or U9223 (N_9223,N_8863,N_8855);
xnor U9224 (N_9224,N_8648,N_8578);
nand U9225 (N_9225,N_8532,N_8935);
and U9226 (N_9226,N_8814,N_8975);
and U9227 (N_9227,N_8892,N_8983);
or U9228 (N_9228,N_8878,N_8625);
nor U9229 (N_9229,N_8738,N_8874);
and U9230 (N_9230,N_8659,N_8722);
nor U9231 (N_9231,N_8939,N_8774);
and U9232 (N_9232,N_8826,N_8614);
nand U9233 (N_9233,N_8534,N_8512);
xor U9234 (N_9234,N_8840,N_8821);
or U9235 (N_9235,N_8744,N_8517);
and U9236 (N_9236,N_8606,N_8811);
or U9237 (N_9237,N_8688,N_8716);
or U9238 (N_9238,N_8900,N_8501);
nand U9239 (N_9239,N_8644,N_8986);
or U9240 (N_9240,N_8958,N_8851);
nor U9241 (N_9241,N_8575,N_8960);
nand U9242 (N_9242,N_8777,N_8522);
xnor U9243 (N_9243,N_8514,N_8599);
and U9244 (N_9244,N_8677,N_8845);
xor U9245 (N_9245,N_8605,N_8641);
and U9246 (N_9246,N_8877,N_8843);
or U9247 (N_9247,N_8766,N_8839);
xnor U9248 (N_9248,N_8810,N_8807);
nand U9249 (N_9249,N_8882,N_8901);
nor U9250 (N_9250,N_8899,N_8836);
nor U9251 (N_9251,N_8639,N_8772);
nor U9252 (N_9252,N_8900,N_8506);
and U9253 (N_9253,N_8802,N_8864);
nor U9254 (N_9254,N_8978,N_8961);
nor U9255 (N_9255,N_8685,N_8651);
xnor U9256 (N_9256,N_8907,N_8603);
nor U9257 (N_9257,N_8642,N_8806);
nand U9258 (N_9258,N_8806,N_8945);
nor U9259 (N_9259,N_8749,N_8739);
and U9260 (N_9260,N_8844,N_8783);
nor U9261 (N_9261,N_8524,N_8812);
or U9262 (N_9262,N_8794,N_8929);
xor U9263 (N_9263,N_8956,N_8853);
and U9264 (N_9264,N_8736,N_8828);
nor U9265 (N_9265,N_8539,N_8804);
or U9266 (N_9266,N_8830,N_8756);
or U9267 (N_9267,N_8623,N_8775);
nand U9268 (N_9268,N_8857,N_8619);
or U9269 (N_9269,N_8881,N_8517);
nand U9270 (N_9270,N_8921,N_8522);
xor U9271 (N_9271,N_8990,N_8528);
and U9272 (N_9272,N_8959,N_8523);
nand U9273 (N_9273,N_8714,N_8887);
and U9274 (N_9274,N_8739,N_8773);
and U9275 (N_9275,N_8563,N_8860);
or U9276 (N_9276,N_8988,N_8626);
or U9277 (N_9277,N_8585,N_8756);
or U9278 (N_9278,N_8662,N_8874);
or U9279 (N_9279,N_8522,N_8697);
and U9280 (N_9280,N_8599,N_8585);
xnor U9281 (N_9281,N_8984,N_8948);
xor U9282 (N_9282,N_8698,N_8669);
nand U9283 (N_9283,N_8745,N_8774);
xnor U9284 (N_9284,N_8640,N_8737);
nor U9285 (N_9285,N_8975,N_8619);
and U9286 (N_9286,N_8519,N_8765);
or U9287 (N_9287,N_8802,N_8647);
xor U9288 (N_9288,N_8659,N_8605);
nand U9289 (N_9289,N_8829,N_8729);
or U9290 (N_9290,N_8562,N_8894);
or U9291 (N_9291,N_8734,N_8633);
nor U9292 (N_9292,N_8931,N_8739);
xor U9293 (N_9293,N_8502,N_8991);
xor U9294 (N_9294,N_8983,N_8920);
nor U9295 (N_9295,N_8618,N_8559);
or U9296 (N_9296,N_8666,N_8957);
nand U9297 (N_9297,N_8718,N_8690);
nor U9298 (N_9298,N_8704,N_8951);
or U9299 (N_9299,N_8545,N_8822);
nand U9300 (N_9300,N_8792,N_8689);
nor U9301 (N_9301,N_8525,N_8938);
or U9302 (N_9302,N_8583,N_8779);
nor U9303 (N_9303,N_8931,N_8595);
or U9304 (N_9304,N_8700,N_8611);
or U9305 (N_9305,N_8519,N_8748);
nand U9306 (N_9306,N_8752,N_8585);
nor U9307 (N_9307,N_8992,N_8741);
nor U9308 (N_9308,N_8703,N_8777);
nor U9309 (N_9309,N_8531,N_8888);
nor U9310 (N_9310,N_8805,N_8614);
and U9311 (N_9311,N_8881,N_8595);
and U9312 (N_9312,N_8722,N_8595);
or U9313 (N_9313,N_8541,N_8727);
nand U9314 (N_9314,N_8616,N_8683);
and U9315 (N_9315,N_8894,N_8773);
nor U9316 (N_9316,N_8983,N_8658);
xor U9317 (N_9317,N_8828,N_8755);
nor U9318 (N_9318,N_8741,N_8731);
or U9319 (N_9319,N_8694,N_8582);
and U9320 (N_9320,N_8880,N_8602);
nand U9321 (N_9321,N_8703,N_8532);
or U9322 (N_9322,N_8720,N_8998);
xor U9323 (N_9323,N_8660,N_8509);
and U9324 (N_9324,N_8771,N_8979);
and U9325 (N_9325,N_8768,N_8585);
nand U9326 (N_9326,N_8644,N_8808);
and U9327 (N_9327,N_8576,N_8706);
and U9328 (N_9328,N_8707,N_8643);
or U9329 (N_9329,N_8883,N_8738);
nor U9330 (N_9330,N_8560,N_8834);
and U9331 (N_9331,N_8994,N_8625);
xnor U9332 (N_9332,N_8719,N_8539);
xor U9333 (N_9333,N_8643,N_8630);
nand U9334 (N_9334,N_8981,N_8579);
nand U9335 (N_9335,N_8997,N_8595);
nor U9336 (N_9336,N_8502,N_8862);
nor U9337 (N_9337,N_8944,N_8609);
and U9338 (N_9338,N_8672,N_8668);
or U9339 (N_9339,N_8550,N_8611);
and U9340 (N_9340,N_8542,N_8537);
nor U9341 (N_9341,N_8655,N_8751);
nand U9342 (N_9342,N_8894,N_8611);
nor U9343 (N_9343,N_8934,N_8568);
nor U9344 (N_9344,N_8509,N_8620);
xnor U9345 (N_9345,N_8698,N_8940);
or U9346 (N_9346,N_8946,N_8942);
nand U9347 (N_9347,N_8617,N_8936);
nor U9348 (N_9348,N_8720,N_8891);
nand U9349 (N_9349,N_8917,N_8981);
nand U9350 (N_9350,N_8918,N_8675);
nand U9351 (N_9351,N_8587,N_8786);
xor U9352 (N_9352,N_8818,N_8632);
nor U9353 (N_9353,N_8829,N_8591);
nand U9354 (N_9354,N_8620,N_8624);
or U9355 (N_9355,N_8612,N_8578);
nor U9356 (N_9356,N_8805,N_8567);
nand U9357 (N_9357,N_8839,N_8980);
xnor U9358 (N_9358,N_8828,N_8617);
nand U9359 (N_9359,N_8873,N_8525);
nand U9360 (N_9360,N_8804,N_8651);
and U9361 (N_9361,N_8799,N_8562);
xnor U9362 (N_9362,N_8623,N_8835);
and U9363 (N_9363,N_8615,N_8912);
or U9364 (N_9364,N_8510,N_8618);
nor U9365 (N_9365,N_8571,N_8737);
nand U9366 (N_9366,N_8771,N_8860);
nand U9367 (N_9367,N_8759,N_8637);
nor U9368 (N_9368,N_8675,N_8554);
xor U9369 (N_9369,N_8611,N_8644);
xnor U9370 (N_9370,N_8766,N_8825);
xnor U9371 (N_9371,N_8801,N_8765);
nor U9372 (N_9372,N_8559,N_8693);
and U9373 (N_9373,N_8677,N_8501);
or U9374 (N_9374,N_8618,N_8647);
nor U9375 (N_9375,N_8657,N_8788);
xnor U9376 (N_9376,N_8541,N_8625);
nand U9377 (N_9377,N_8986,N_8544);
or U9378 (N_9378,N_8567,N_8774);
or U9379 (N_9379,N_8989,N_8961);
nor U9380 (N_9380,N_8984,N_8577);
and U9381 (N_9381,N_8664,N_8986);
nand U9382 (N_9382,N_8588,N_8759);
nand U9383 (N_9383,N_8558,N_8827);
or U9384 (N_9384,N_8963,N_8954);
nand U9385 (N_9385,N_8967,N_8614);
nand U9386 (N_9386,N_8763,N_8851);
or U9387 (N_9387,N_8765,N_8983);
xnor U9388 (N_9388,N_8838,N_8674);
nor U9389 (N_9389,N_8861,N_8630);
nand U9390 (N_9390,N_8570,N_8679);
and U9391 (N_9391,N_8998,N_8870);
or U9392 (N_9392,N_8857,N_8660);
and U9393 (N_9393,N_8759,N_8612);
nor U9394 (N_9394,N_8619,N_8634);
or U9395 (N_9395,N_8569,N_8592);
or U9396 (N_9396,N_8914,N_8791);
nand U9397 (N_9397,N_8921,N_8863);
nand U9398 (N_9398,N_8604,N_8871);
nor U9399 (N_9399,N_8618,N_8861);
nand U9400 (N_9400,N_8729,N_8939);
and U9401 (N_9401,N_8514,N_8922);
nand U9402 (N_9402,N_8800,N_8817);
or U9403 (N_9403,N_8947,N_8833);
nand U9404 (N_9404,N_8749,N_8906);
nand U9405 (N_9405,N_8909,N_8981);
or U9406 (N_9406,N_8569,N_8652);
nor U9407 (N_9407,N_8551,N_8568);
or U9408 (N_9408,N_8902,N_8805);
and U9409 (N_9409,N_8754,N_8530);
nand U9410 (N_9410,N_8526,N_8765);
nand U9411 (N_9411,N_8803,N_8907);
nor U9412 (N_9412,N_8561,N_8747);
or U9413 (N_9413,N_8517,N_8555);
and U9414 (N_9414,N_8511,N_8506);
and U9415 (N_9415,N_8586,N_8914);
nor U9416 (N_9416,N_8878,N_8978);
or U9417 (N_9417,N_8633,N_8982);
xor U9418 (N_9418,N_8699,N_8721);
and U9419 (N_9419,N_8643,N_8808);
and U9420 (N_9420,N_8544,N_8827);
nand U9421 (N_9421,N_8512,N_8599);
nand U9422 (N_9422,N_8730,N_8989);
nand U9423 (N_9423,N_8547,N_8502);
nor U9424 (N_9424,N_8754,N_8833);
nand U9425 (N_9425,N_8609,N_8527);
or U9426 (N_9426,N_8532,N_8921);
nor U9427 (N_9427,N_8509,N_8823);
nor U9428 (N_9428,N_8750,N_8957);
and U9429 (N_9429,N_8532,N_8818);
and U9430 (N_9430,N_8528,N_8788);
and U9431 (N_9431,N_8559,N_8578);
xor U9432 (N_9432,N_8622,N_8961);
nor U9433 (N_9433,N_8643,N_8581);
xor U9434 (N_9434,N_8609,N_8869);
nor U9435 (N_9435,N_8941,N_8584);
xnor U9436 (N_9436,N_8545,N_8726);
or U9437 (N_9437,N_8659,N_8607);
and U9438 (N_9438,N_8729,N_8517);
nand U9439 (N_9439,N_8972,N_8570);
nor U9440 (N_9440,N_8795,N_8810);
nand U9441 (N_9441,N_8885,N_8930);
nor U9442 (N_9442,N_8887,N_8730);
xor U9443 (N_9443,N_8515,N_8651);
nand U9444 (N_9444,N_8881,N_8831);
or U9445 (N_9445,N_8508,N_8503);
or U9446 (N_9446,N_8606,N_8549);
nand U9447 (N_9447,N_8949,N_8847);
nor U9448 (N_9448,N_8515,N_8745);
or U9449 (N_9449,N_8785,N_8763);
xor U9450 (N_9450,N_8677,N_8858);
nor U9451 (N_9451,N_8658,N_8568);
or U9452 (N_9452,N_8925,N_8983);
xor U9453 (N_9453,N_8845,N_8827);
nand U9454 (N_9454,N_8990,N_8769);
nand U9455 (N_9455,N_8831,N_8708);
and U9456 (N_9456,N_8998,N_8608);
nand U9457 (N_9457,N_8953,N_8937);
or U9458 (N_9458,N_8878,N_8809);
nand U9459 (N_9459,N_8821,N_8950);
and U9460 (N_9460,N_8764,N_8818);
nand U9461 (N_9461,N_8955,N_8908);
and U9462 (N_9462,N_8640,N_8956);
xor U9463 (N_9463,N_8543,N_8946);
and U9464 (N_9464,N_8804,N_8597);
and U9465 (N_9465,N_8631,N_8591);
nand U9466 (N_9466,N_8705,N_8820);
and U9467 (N_9467,N_8686,N_8672);
or U9468 (N_9468,N_8693,N_8507);
and U9469 (N_9469,N_8886,N_8962);
xnor U9470 (N_9470,N_8650,N_8536);
and U9471 (N_9471,N_8672,N_8780);
xor U9472 (N_9472,N_8550,N_8624);
and U9473 (N_9473,N_8627,N_8711);
or U9474 (N_9474,N_8512,N_8545);
or U9475 (N_9475,N_8782,N_8570);
and U9476 (N_9476,N_8866,N_8921);
or U9477 (N_9477,N_8700,N_8647);
nand U9478 (N_9478,N_8842,N_8926);
xor U9479 (N_9479,N_8773,N_8837);
xnor U9480 (N_9480,N_8653,N_8657);
or U9481 (N_9481,N_8757,N_8647);
xnor U9482 (N_9482,N_8757,N_8916);
or U9483 (N_9483,N_8568,N_8855);
nand U9484 (N_9484,N_8747,N_8978);
or U9485 (N_9485,N_8589,N_8532);
xnor U9486 (N_9486,N_8599,N_8546);
and U9487 (N_9487,N_8774,N_8500);
xor U9488 (N_9488,N_8584,N_8748);
nand U9489 (N_9489,N_8844,N_8974);
nor U9490 (N_9490,N_8709,N_8801);
xnor U9491 (N_9491,N_8655,N_8681);
nor U9492 (N_9492,N_8722,N_8966);
xnor U9493 (N_9493,N_8779,N_8703);
xnor U9494 (N_9494,N_8503,N_8586);
xnor U9495 (N_9495,N_8639,N_8729);
nor U9496 (N_9496,N_8576,N_8872);
and U9497 (N_9497,N_8821,N_8744);
xnor U9498 (N_9498,N_8694,N_8526);
and U9499 (N_9499,N_8821,N_8920);
and U9500 (N_9500,N_9381,N_9456);
and U9501 (N_9501,N_9289,N_9180);
and U9502 (N_9502,N_9075,N_9020);
nand U9503 (N_9503,N_9401,N_9414);
and U9504 (N_9504,N_9417,N_9394);
or U9505 (N_9505,N_9123,N_9205);
or U9506 (N_9506,N_9151,N_9344);
xor U9507 (N_9507,N_9101,N_9340);
and U9508 (N_9508,N_9014,N_9279);
xnor U9509 (N_9509,N_9326,N_9231);
nand U9510 (N_9510,N_9089,N_9094);
or U9511 (N_9511,N_9405,N_9469);
and U9512 (N_9512,N_9422,N_9461);
and U9513 (N_9513,N_9479,N_9114);
or U9514 (N_9514,N_9388,N_9441);
nor U9515 (N_9515,N_9130,N_9272);
xnor U9516 (N_9516,N_9271,N_9309);
nand U9517 (N_9517,N_9131,N_9187);
xnor U9518 (N_9518,N_9413,N_9190);
nand U9519 (N_9519,N_9323,N_9008);
nor U9520 (N_9520,N_9029,N_9030);
or U9521 (N_9521,N_9162,N_9066);
or U9522 (N_9522,N_9305,N_9111);
or U9523 (N_9523,N_9328,N_9297);
xor U9524 (N_9524,N_9005,N_9332);
nor U9525 (N_9525,N_9063,N_9474);
and U9526 (N_9526,N_9443,N_9356);
xor U9527 (N_9527,N_9428,N_9113);
or U9528 (N_9528,N_9085,N_9433);
and U9529 (N_9529,N_9412,N_9498);
nand U9530 (N_9530,N_9380,N_9056);
xnor U9531 (N_9531,N_9216,N_9172);
and U9532 (N_9532,N_9354,N_9124);
nand U9533 (N_9533,N_9165,N_9472);
or U9534 (N_9534,N_9319,N_9200);
and U9535 (N_9535,N_9310,N_9296);
and U9536 (N_9536,N_9438,N_9211);
nor U9537 (N_9537,N_9107,N_9415);
or U9538 (N_9538,N_9228,N_9459);
nand U9539 (N_9539,N_9320,N_9284);
xor U9540 (N_9540,N_9084,N_9269);
or U9541 (N_9541,N_9496,N_9062);
nand U9542 (N_9542,N_9206,N_9440);
xor U9543 (N_9543,N_9432,N_9213);
and U9544 (N_9544,N_9159,N_9396);
xor U9545 (N_9545,N_9455,N_9343);
nand U9546 (N_9546,N_9088,N_9349);
or U9547 (N_9547,N_9091,N_9482);
xnor U9548 (N_9548,N_9135,N_9152);
and U9549 (N_9549,N_9032,N_9120);
or U9550 (N_9550,N_9076,N_9402);
nor U9551 (N_9551,N_9458,N_9290);
and U9552 (N_9552,N_9308,N_9072);
and U9553 (N_9553,N_9341,N_9292);
nor U9554 (N_9554,N_9490,N_9257);
and U9555 (N_9555,N_9092,N_9436);
xnor U9556 (N_9556,N_9125,N_9225);
or U9557 (N_9557,N_9423,N_9036);
xnor U9558 (N_9558,N_9361,N_9002);
xnor U9559 (N_9559,N_9276,N_9170);
nor U9560 (N_9560,N_9024,N_9480);
nand U9561 (N_9561,N_9406,N_9463);
or U9562 (N_9562,N_9383,N_9424);
nor U9563 (N_9563,N_9258,N_9015);
or U9564 (N_9564,N_9444,N_9301);
and U9565 (N_9565,N_9363,N_9001);
and U9566 (N_9566,N_9453,N_9194);
and U9567 (N_9567,N_9153,N_9095);
and U9568 (N_9568,N_9337,N_9163);
nand U9569 (N_9569,N_9389,N_9046);
nand U9570 (N_9570,N_9334,N_9379);
nand U9571 (N_9571,N_9287,N_9099);
nand U9572 (N_9572,N_9179,N_9331);
nor U9573 (N_9573,N_9100,N_9385);
nor U9574 (N_9574,N_9188,N_9298);
xnor U9575 (N_9575,N_9398,N_9322);
xnor U9576 (N_9576,N_9336,N_9057);
and U9577 (N_9577,N_9265,N_9311);
and U9578 (N_9578,N_9294,N_9350);
nor U9579 (N_9579,N_9446,N_9223);
nand U9580 (N_9580,N_9460,N_9467);
nor U9581 (N_9581,N_9329,N_9489);
nand U9582 (N_9582,N_9366,N_9359);
nand U9583 (N_9583,N_9185,N_9318);
nand U9584 (N_9584,N_9355,N_9249);
xor U9585 (N_9585,N_9374,N_9477);
xnor U9586 (N_9586,N_9220,N_9207);
and U9587 (N_9587,N_9410,N_9486);
and U9588 (N_9588,N_9182,N_9462);
nor U9589 (N_9589,N_9164,N_9173);
xor U9590 (N_9590,N_9019,N_9260);
and U9591 (N_9591,N_9420,N_9251);
and U9592 (N_9592,N_9430,N_9321);
xor U9593 (N_9593,N_9468,N_9484);
nand U9594 (N_9594,N_9222,N_9497);
or U9595 (N_9595,N_9244,N_9335);
xnor U9596 (N_9596,N_9006,N_9115);
nor U9597 (N_9597,N_9055,N_9028);
and U9598 (N_9598,N_9473,N_9390);
nor U9599 (N_9599,N_9080,N_9395);
xnor U9600 (N_9600,N_9313,N_9058);
and U9601 (N_9601,N_9189,N_9407);
or U9602 (N_9602,N_9312,N_9226);
or U9603 (N_9603,N_9397,N_9068);
or U9604 (N_9604,N_9348,N_9262);
and U9605 (N_9605,N_9302,N_9465);
nor U9606 (N_9606,N_9176,N_9218);
nand U9607 (N_9607,N_9049,N_9025);
and U9608 (N_9608,N_9481,N_9122);
nor U9609 (N_9609,N_9300,N_9248);
nor U9610 (N_9610,N_9096,N_9007);
nand U9611 (N_9611,N_9060,N_9450);
nand U9612 (N_9612,N_9045,N_9384);
nor U9613 (N_9613,N_9017,N_9471);
nand U9614 (N_9614,N_9035,N_9147);
and U9615 (N_9615,N_9202,N_9138);
nand U9616 (N_9616,N_9104,N_9171);
nand U9617 (N_9617,N_9016,N_9454);
or U9618 (N_9618,N_9050,N_9105);
xor U9619 (N_9619,N_9476,N_9373);
and U9620 (N_9620,N_9169,N_9464);
xor U9621 (N_9621,N_9090,N_9181);
xor U9622 (N_9622,N_9252,N_9408);
or U9623 (N_9623,N_9375,N_9266);
nand U9624 (N_9624,N_9042,N_9175);
or U9625 (N_9625,N_9421,N_9203);
or U9626 (N_9626,N_9136,N_9208);
xor U9627 (N_9627,N_9209,N_9283);
and U9628 (N_9628,N_9419,N_9010);
and U9629 (N_9629,N_9259,N_9437);
or U9630 (N_9630,N_9439,N_9198);
nor U9631 (N_9631,N_9186,N_9011);
nor U9632 (N_9632,N_9143,N_9134);
or U9633 (N_9633,N_9132,N_9081);
xnor U9634 (N_9634,N_9447,N_9493);
nor U9635 (N_9635,N_9478,N_9048);
or U9636 (N_9636,N_9177,N_9280);
or U9637 (N_9637,N_9038,N_9235);
or U9638 (N_9638,N_9061,N_9485);
and U9639 (N_9639,N_9285,N_9103);
or U9640 (N_9640,N_9369,N_9118);
nor U9641 (N_9641,N_9195,N_9034);
and U9642 (N_9642,N_9346,N_9362);
xor U9643 (N_9643,N_9204,N_9238);
or U9644 (N_9644,N_9256,N_9387);
nor U9645 (N_9645,N_9315,N_9426);
nor U9646 (N_9646,N_9360,N_9261);
xnor U9647 (N_9647,N_9393,N_9012);
nand U9648 (N_9648,N_9357,N_9270);
nand U9649 (N_9649,N_9009,N_9133);
nor U9650 (N_9650,N_9316,N_9110);
and U9651 (N_9651,N_9021,N_9377);
and U9652 (N_9652,N_9221,N_9031);
and U9653 (N_9653,N_9126,N_9342);
nand U9654 (N_9654,N_9214,N_9442);
nor U9655 (N_9655,N_9303,N_9037);
and U9656 (N_9656,N_9364,N_9119);
xor U9657 (N_9657,N_9102,N_9215);
or U9658 (N_9658,N_9137,N_9347);
and U9659 (N_9659,N_9083,N_9059);
nor U9660 (N_9660,N_9196,N_9033);
and U9661 (N_9661,N_9053,N_9487);
nor U9662 (N_9662,N_9026,N_9404);
nor U9663 (N_9663,N_9418,N_9027);
nand U9664 (N_9664,N_9212,N_9082);
nand U9665 (N_9665,N_9155,N_9064);
nor U9666 (N_9666,N_9365,N_9087);
and U9667 (N_9667,N_9466,N_9086);
nand U9668 (N_9668,N_9191,N_9229);
xor U9669 (N_9669,N_9116,N_9304);
and U9670 (N_9670,N_9254,N_9041);
or U9671 (N_9671,N_9077,N_9161);
nor U9672 (N_9672,N_9098,N_9451);
xnor U9673 (N_9673,N_9241,N_9475);
and U9674 (N_9674,N_9386,N_9178);
nor U9675 (N_9675,N_9399,N_9149);
or U9676 (N_9676,N_9314,N_9047);
or U9677 (N_9677,N_9234,N_9367);
nor U9678 (N_9678,N_9370,N_9154);
nor U9679 (N_9679,N_9106,N_9307);
or U9680 (N_9680,N_9192,N_9470);
nor U9681 (N_9681,N_9457,N_9264);
or U9682 (N_9682,N_9071,N_9250);
nor U9683 (N_9683,N_9267,N_9378);
nand U9684 (N_9684,N_9184,N_9112);
xor U9685 (N_9685,N_9376,N_9141);
xor U9686 (N_9686,N_9158,N_9070);
nor U9687 (N_9687,N_9148,N_9452);
nor U9688 (N_9688,N_9140,N_9293);
nand U9689 (N_9689,N_9109,N_9353);
xnor U9690 (N_9690,N_9074,N_9183);
nand U9691 (N_9691,N_9324,N_9278);
xnor U9692 (N_9692,N_9274,N_9492);
nand U9693 (N_9693,N_9330,N_9067);
nand U9694 (N_9694,N_9345,N_9372);
or U9695 (N_9695,N_9145,N_9239);
nand U9696 (N_9696,N_9224,N_9051);
or U9697 (N_9697,N_9160,N_9210);
xnor U9698 (N_9698,N_9243,N_9142);
and U9699 (N_9699,N_9128,N_9144);
or U9700 (N_9700,N_9127,N_9448);
nand U9701 (N_9701,N_9351,N_9167);
and U9702 (N_9702,N_9429,N_9277);
xor U9703 (N_9703,N_9227,N_9263);
nand U9704 (N_9704,N_9018,N_9382);
nand U9705 (N_9705,N_9317,N_9201);
or U9706 (N_9706,N_9236,N_9065);
and U9707 (N_9707,N_9282,N_9295);
nor U9708 (N_9708,N_9168,N_9232);
and U9709 (N_9709,N_9499,N_9233);
or U9710 (N_9710,N_9425,N_9445);
nand U9711 (N_9711,N_9253,N_9416);
nor U9712 (N_9712,N_9157,N_9409);
or U9713 (N_9713,N_9255,N_9327);
nand U9714 (N_9714,N_9146,N_9245);
nor U9715 (N_9715,N_9400,N_9097);
or U9716 (N_9716,N_9054,N_9039);
and U9717 (N_9717,N_9022,N_9219);
and U9718 (N_9718,N_9197,N_9411);
xnor U9719 (N_9719,N_9495,N_9281);
and U9720 (N_9720,N_9242,N_9273);
and U9721 (N_9721,N_9494,N_9358);
nand U9722 (N_9722,N_9434,N_9325);
and U9723 (N_9723,N_9000,N_9431);
and U9724 (N_9724,N_9139,N_9093);
or U9725 (N_9725,N_9275,N_9427);
nor U9726 (N_9726,N_9043,N_9117);
and U9727 (N_9727,N_9291,N_9352);
xnor U9728 (N_9728,N_9023,N_9286);
nand U9729 (N_9729,N_9392,N_9217);
or U9730 (N_9730,N_9013,N_9052);
nand U9731 (N_9731,N_9240,N_9488);
nor U9732 (N_9732,N_9069,N_9150);
and U9733 (N_9733,N_9199,N_9333);
nor U9734 (N_9734,N_9193,N_9491);
xor U9735 (N_9735,N_9166,N_9247);
nand U9736 (N_9736,N_9368,N_9079);
nand U9737 (N_9737,N_9403,N_9371);
nor U9738 (N_9738,N_9044,N_9268);
or U9739 (N_9739,N_9156,N_9078);
or U9740 (N_9740,N_9230,N_9338);
nor U9741 (N_9741,N_9174,N_9435);
and U9742 (N_9742,N_9003,N_9121);
and U9743 (N_9743,N_9391,N_9483);
xor U9744 (N_9744,N_9246,N_9299);
nand U9745 (N_9745,N_9306,N_9288);
and U9746 (N_9746,N_9129,N_9449);
and U9747 (N_9747,N_9040,N_9339);
nand U9748 (N_9748,N_9073,N_9108);
nand U9749 (N_9749,N_9237,N_9004);
nand U9750 (N_9750,N_9369,N_9386);
nor U9751 (N_9751,N_9161,N_9085);
nand U9752 (N_9752,N_9370,N_9276);
nor U9753 (N_9753,N_9230,N_9134);
nand U9754 (N_9754,N_9192,N_9246);
or U9755 (N_9755,N_9463,N_9346);
and U9756 (N_9756,N_9427,N_9370);
xnor U9757 (N_9757,N_9290,N_9376);
xor U9758 (N_9758,N_9329,N_9403);
xnor U9759 (N_9759,N_9142,N_9378);
or U9760 (N_9760,N_9023,N_9106);
nand U9761 (N_9761,N_9097,N_9180);
nand U9762 (N_9762,N_9359,N_9251);
and U9763 (N_9763,N_9011,N_9328);
xnor U9764 (N_9764,N_9463,N_9282);
nor U9765 (N_9765,N_9288,N_9477);
nor U9766 (N_9766,N_9297,N_9350);
and U9767 (N_9767,N_9177,N_9381);
xnor U9768 (N_9768,N_9164,N_9263);
xor U9769 (N_9769,N_9021,N_9405);
nor U9770 (N_9770,N_9456,N_9284);
nor U9771 (N_9771,N_9141,N_9163);
xnor U9772 (N_9772,N_9392,N_9445);
nand U9773 (N_9773,N_9062,N_9032);
and U9774 (N_9774,N_9247,N_9281);
nand U9775 (N_9775,N_9072,N_9330);
nor U9776 (N_9776,N_9421,N_9336);
nor U9777 (N_9777,N_9047,N_9457);
or U9778 (N_9778,N_9490,N_9477);
and U9779 (N_9779,N_9460,N_9342);
and U9780 (N_9780,N_9181,N_9081);
xor U9781 (N_9781,N_9087,N_9498);
nor U9782 (N_9782,N_9450,N_9336);
nand U9783 (N_9783,N_9275,N_9280);
or U9784 (N_9784,N_9099,N_9342);
and U9785 (N_9785,N_9491,N_9090);
xor U9786 (N_9786,N_9180,N_9383);
xor U9787 (N_9787,N_9293,N_9021);
and U9788 (N_9788,N_9128,N_9206);
xor U9789 (N_9789,N_9054,N_9416);
xor U9790 (N_9790,N_9124,N_9075);
or U9791 (N_9791,N_9446,N_9181);
or U9792 (N_9792,N_9095,N_9076);
xnor U9793 (N_9793,N_9223,N_9375);
nand U9794 (N_9794,N_9316,N_9049);
nor U9795 (N_9795,N_9443,N_9285);
and U9796 (N_9796,N_9377,N_9014);
nand U9797 (N_9797,N_9385,N_9053);
and U9798 (N_9798,N_9358,N_9482);
nand U9799 (N_9799,N_9136,N_9259);
xor U9800 (N_9800,N_9076,N_9018);
and U9801 (N_9801,N_9368,N_9062);
and U9802 (N_9802,N_9223,N_9246);
xor U9803 (N_9803,N_9274,N_9182);
and U9804 (N_9804,N_9356,N_9084);
or U9805 (N_9805,N_9101,N_9433);
nand U9806 (N_9806,N_9115,N_9360);
nor U9807 (N_9807,N_9098,N_9400);
or U9808 (N_9808,N_9415,N_9455);
xnor U9809 (N_9809,N_9488,N_9228);
and U9810 (N_9810,N_9238,N_9358);
nor U9811 (N_9811,N_9066,N_9253);
or U9812 (N_9812,N_9139,N_9165);
and U9813 (N_9813,N_9447,N_9496);
nand U9814 (N_9814,N_9009,N_9293);
xnor U9815 (N_9815,N_9462,N_9160);
xor U9816 (N_9816,N_9443,N_9101);
nand U9817 (N_9817,N_9380,N_9412);
and U9818 (N_9818,N_9306,N_9378);
xor U9819 (N_9819,N_9158,N_9498);
and U9820 (N_9820,N_9330,N_9488);
and U9821 (N_9821,N_9087,N_9350);
nand U9822 (N_9822,N_9325,N_9066);
xor U9823 (N_9823,N_9143,N_9233);
xor U9824 (N_9824,N_9027,N_9001);
or U9825 (N_9825,N_9006,N_9323);
xnor U9826 (N_9826,N_9435,N_9115);
nand U9827 (N_9827,N_9178,N_9129);
nand U9828 (N_9828,N_9031,N_9278);
xnor U9829 (N_9829,N_9485,N_9318);
or U9830 (N_9830,N_9233,N_9251);
nor U9831 (N_9831,N_9370,N_9067);
and U9832 (N_9832,N_9135,N_9389);
and U9833 (N_9833,N_9036,N_9337);
and U9834 (N_9834,N_9217,N_9123);
xnor U9835 (N_9835,N_9131,N_9210);
and U9836 (N_9836,N_9253,N_9118);
nor U9837 (N_9837,N_9362,N_9116);
or U9838 (N_9838,N_9324,N_9251);
nor U9839 (N_9839,N_9225,N_9039);
xor U9840 (N_9840,N_9054,N_9266);
nand U9841 (N_9841,N_9222,N_9408);
nor U9842 (N_9842,N_9299,N_9261);
nand U9843 (N_9843,N_9057,N_9122);
xor U9844 (N_9844,N_9426,N_9048);
xnor U9845 (N_9845,N_9354,N_9271);
or U9846 (N_9846,N_9398,N_9138);
nor U9847 (N_9847,N_9162,N_9438);
or U9848 (N_9848,N_9444,N_9365);
or U9849 (N_9849,N_9176,N_9120);
or U9850 (N_9850,N_9268,N_9133);
and U9851 (N_9851,N_9026,N_9343);
and U9852 (N_9852,N_9364,N_9329);
and U9853 (N_9853,N_9337,N_9013);
or U9854 (N_9854,N_9119,N_9291);
and U9855 (N_9855,N_9088,N_9237);
and U9856 (N_9856,N_9057,N_9267);
xor U9857 (N_9857,N_9222,N_9042);
nand U9858 (N_9858,N_9402,N_9399);
or U9859 (N_9859,N_9013,N_9100);
and U9860 (N_9860,N_9408,N_9396);
xnor U9861 (N_9861,N_9054,N_9315);
nor U9862 (N_9862,N_9121,N_9153);
and U9863 (N_9863,N_9153,N_9455);
nand U9864 (N_9864,N_9135,N_9435);
or U9865 (N_9865,N_9035,N_9480);
or U9866 (N_9866,N_9151,N_9122);
nand U9867 (N_9867,N_9424,N_9161);
nor U9868 (N_9868,N_9197,N_9452);
and U9869 (N_9869,N_9103,N_9008);
xnor U9870 (N_9870,N_9225,N_9218);
nor U9871 (N_9871,N_9403,N_9464);
nor U9872 (N_9872,N_9308,N_9393);
nor U9873 (N_9873,N_9007,N_9232);
xor U9874 (N_9874,N_9458,N_9017);
nand U9875 (N_9875,N_9446,N_9028);
nand U9876 (N_9876,N_9492,N_9093);
nor U9877 (N_9877,N_9423,N_9357);
and U9878 (N_9878,N_9391,N_9298);
and U9879 (N_9879,N_9473,N_9009);
and U9880 (N_9880,N_9293,N_9160);
nand U9881 (N_9881,N_9493,N_9075);
nand U9882 (N_9882,N_9030,N_9283);
nand U9883 (N_9883,N_9254,N_9138);
xnor U9884 (N_9884,N_9089,N_9348);
xnor U9885 (N_9885,N_9445,N_9298);
nor U9886 (N_9886,N_9478,N_9234);
nand U9887 (N_9887,N_9024,N_9295);
nand U9888 (N_9888,N_9191,N_9257);
nor U9889 (N_9889,N_9062,N_9302);
and U9890 (N_9890,N_9467,N_9005);
or U9891 (N_9891,N_9311,N_9163);
and U9892 (N_9892,N_9174,N_9176);
nor U9893 (N_9893,N_9349,N_9482);
nand U9894 (N_9894,N_9409,N_9499);
xnor U9895 (N_9895,N_9110,N_9056);
or U9896 (N_9896,N_9101,N_9193);
xor U9897 (N_9897,N_9088,N_9047);
xor U9898 (N_9898,N_9385,N_9058);
nor U9899 (N_9899,N_9337,N_9325);
nand U9900 (N_9900,N_9269,N_9453);
nand U9901 (N_9901,N_9494,N_9043);
nor U9902 (N_9902,N_9033,N_9148);
nand U9903 (N_9903,N_9016,N_9088);
xor U9904 (N_9904,N_9112,N_9307);
or U9905 (N_9905,N_9064,N_9121);
or U9906 (N_9906,N_9058,N_9125);
nor U9907 (N_9907,N_9015,N_9035);
and U9908 (N_9908,N_9180,N_9471);
nor U9909 (N_9909,N_9189,N_9183);
xor U9910 (N_9910,N_9346,N_9073);
and U9911 (N_9911,N_9457,N_9210);
and U9912 (N_9912,N_9400,N_9015);
nand U9913 (N_9913,N_9296,N_9092);
nand U9914 (N_9914,N_9132,N_9000);
or U9915 (N_9915,N_9361,N_9229);
nand U9916 (N_9916,N_9389,N_9304);
nand U9917 (N_9917,N_9130,N_9126);
xnor U9918 (N_9918,N_9168,N_9162);
nand U9919 (N_9919,N_9424,N_9362);
nand U9920 (N_9920,N_9069,N_9049);
and U9921 (N_9921,N_9053,N_9223);
or U9922 (N_9922,N_9121,N_9080);
xor U9923 (N_9923,N_9167,N_9010);
or U9924 (N_9924,N_9464,N_9295);
xnor U9925 (N_9925,N_9474,N_9447);
or U9926 (N_9926,N_9046,N_9297);
nand U9927 (N_9927,N_9302,N_9311);
or U9928 (N_9928,N_9251,N_9088);
xnor U9929 (N_9929,N_9040,N_9319);
xor U9930 (N_9930,N_9401,N_9333);
and U9931 (N_9931,N_9065,N_9282);
and U9932 (N_9932,N_9337,N_9250);
and U9933 (N_9933,N_9375,N_9384);
and U9934 (N_9934,N_9273,N_9122);
or U9935 (N_9935,N_9280,N_9325);
and U9936 (N_9936,N_9399,N_9322);
nor U9937 (N_9937,N_9243,N_9365);
or U9938 (N_9938,N_9299,N_9148);
or U9939 (N_9939,N_9155,N_9012);
xor U9940 (N_9940,N_9264,N_9108);
and U9941 (N_9941,N_9305,N_9255);
nand U9942 (N_9942,N_9059,N_9423);
and U9943 (N_9943,N_9205,N_9105);
nand U9944 (N_9944,N_9426,N_9436);
and U9945 (N_9945,N_9062,N_9470);
nor U9946 (N_9946,N_9439,N_9074);
or U9947 (N_9947,N_9246,N_9023);
nand U9948 (N_9948,N_9349,N_9041);
nand U9949 (N_9949,N_9241,N_9013);
nor U9950 (N_9950,N_9108,N_9472);
xor U9951 (N_9951,N_9441,N_9466);
nor U9952 (N_9952,N_9065,N_9170);
nor U9953 (N_9953,N_9213,N_9026);
nand U9954 (N_9954,N_9053,N_9311);
nand U9955 (N_9955,N_9275,N_9375);
or U9956 (N_9956,N_9416,N_9240);
or U9957 (N_9957,N_9388,N_9396);
and U9958 (N_9958,N_9025,N_9147);
xor U9959 (N_9959,N_9417,N_9174);
xor U9960 (N_9960,N_9323,N_9415);
and U9961 (N_9961,N_9400,N_9195);
nor U9962 (N_9962,N_9028,N_9189);
nand U9963 (N_9963,N_9215,N_9024);
and U9964 (N_9964,N_9448,N_9383);
nor U9965 (N_9965,N_9432,N_9405);
nor U9966 (N_9966,N_9421,N_9365);
nand U9967 (N_9967,N_9307,N_9473);
nand U9968 (N_9968,N_9465,N_9228);
nand U9969 (N_9969,N_9014,N_9287);
nor U9970 (N_9970,N_9198,N_9328);
and U9971 (N_9971,N_9425,N_9378);
nand U9972 (N_9972,N_9349,N_9043);
xor U9973 (N_9973,N_9108,N_9290);
xor U9974 (N_9974,N_9025,N_9162);
nand U9975 (N_9975,N_9039,N_9232);
and U9976 (N_9976,N_9068,N_9000);
xnor U9977 (N_9977,N_9083,N_9016);
nand U9978 (N_9978,N_9156,N_9258);
nor U9979 (N_9979,N_9498,N_9062);
and U9980 (N_9980,N_9433,N_9200);
nor U9981 (N_9981,N_9277,N_9445);
nand U9982 (N_9982,N_9194,N_9458);
nand U9983 (N_9983,N_9104,N_9351);
or U9984 (N_9984,N_9421,N_9348);
and U9985 (N_9985,N_9218,N_9215);
nor U9986 (N_9986,N_9120,N_9303);
or U9987 (N_9987,N_9082,N_9402);
or U9988 (N_9988,N_9340,N_9129);
xnor U9989 (N_9989,N_9147,N_9451);
or U9990 (N_9990,N_9491,N_9280);
xor U9991 (N_9991,N_9107,N_9484);
and U9992 (N_9992,N_9190,N_9298);
nand U9993 (N_9993,N_9163,N_9449);
and U9994 (N_9994,N_9060,N_9186);
nor U9995 (N_9995,N_9211,N_9270);
nand U9996 (N_9996,N_9294,N_9278);
and U9997 (N_9997,N_9197,N_9162);
nand U9998 (N_9998,N_9153,N_9241);
and U9999 (N_9999,N_9200,N_9291);
nand U10000 (N_10000,N_9753,N_9621);
nand U10001 (N_10001,N_9817,N_9906);
nand U10002 (N_10002,N_9530,N_9628);
or U10003 (N_10003,N_9934,N_9733);
xnor U10004 (N_10004,N_9611,N_9637);
and U10005 (N_10005,N_9552,N_9822);
and U10006 (N_10006,N_9506,N_9879);
nor U10007 (N_10007,N_9760,N_9531);
nor U10008 (N_10008,N_9781,N_9728);
xor U10009 (N_10009,N_9620,N_9612);
and U10010 (N_10010,N_9588,N_9654);
nor U10011 (N_10011,N_9955,N_9695);
xor U10012 (N_10012,N_9761,N_9785);
and U10013 (N_10013,N_9547,N_9975);
nand U10014 (N_10014,N_9502,N_9820);
nor U10015 (N_10015,N_9591,N_9756);
nor U10016 (N_10016,N_9882,N_9897);
nor U10017 (N_10017,N_9856,N_9965);
and U10018 (N_10018,N_9925,N_9952);
nor U10019 (N_10019,N_9851,N_9682);
nand U10020 (N_10020,N_9824,N_9624);
nor U10021 (N_10021,N_9902,N_9796);
nor U10022 (N_10022,N_9821,N_9566);
nor U10023 (N_10023,N_9572,N_9544);
nor U10024 (N_10024,N_9729,N_9545);
nand U10025 (N_10025,N_9635,N_9935);
nand U10026 (N_10026,N_9770,N_9992);
or U10027 (N_10027,N_9896,N_9751);
nor U10028 (N_10028,N_9859,N_9833);
nor U10029 (N_10029,N_9720,N_9806);
nor U10030 (N_10030,N_9782,N_9762);
xnor U10031 (N_10031,N_9765,N_9528);
nand U10032 (N_10032,N_9581,N_9798);
xor U10033 (N_10033,N_9533,N_9589);
nor U10034 (N_10034,N_9959,N_9986);
nand U10035 (N_10035,N_9954,N_9501);
nand U10036 (N_10036,N_9972,N_9605);
nor U10037 (N_10037,N_9854,N_9692);
nand U10038 (N_10038,N_9800,N_9953);
xnor U10039 (N_10039,N_9691,N_9799);
nor U10040 (N_10040,N_9909,N_9746);
or U10041 (N_10041,N_9601,N_9869);
nor U10042 (N_10042,N_9863,N_9521);
and U10043 (N_10043,N_9561,N_9562);
nand U10044 (N_10044,N_9776,N_9685);
or U10045 (N_10045,N_9910,N_9650);
nor U10046 (N_10046,N_9716,N_9939);
nor U10047 (N_10047,N_9744,N_9858);
nand U10048 (N_10048,N_9919,N_9597);
nand U10049 (N_10049,N_9632,N_9887);
and U10050 (N_10050,N_9513,N_9641);
xor U10051 (N_10051,N_9922,N_9725);
nand U10052 (N_10052,N_9866,N_9842);
nand U10053 (N_10053,N_9884,N_9907);
and U10054 (N_10054,N_9646,N_9715);
nand U10055 (N_10055,N_9895,N_9898);
and U10056 (N_10056,N_9633,N_9793);
nor U10057 (N_10057,N_9541,N_9996);
or U10058 (N_10058,N_9764,N_9981);
nand U10059 (N_10059,N_9525,N_9985);
nor U10060 (N_10060,N_9915,N_9890);
xor U10061 (N_10061,N_9701,N_9623);
nor U10062 (N_10062,N_9938,N_9787);
nor U10063 (N_10063,N_9629,N_9943);
or U10064 (N_10064,N_9510,N_9571);
nand U10065 (N_10065,N_9698,N_9536);
and U10066 (N_10066,N_9944,N_9679);
or U10067 (N_10067,N_9757,N_9994);
nor U10068 (N_10068,N_9941,N_9747);
nor U10069 (N_10069,N_9845,N_9967);
xnor U10070 (N_10070,N_9860,N_9738);
and U10071 (N_10071,N_9559,N_9514);
nand U10072 (N_10072,N_9576,N_9529);
nand U10073 (N_10073,N_9853,N_9710);
nor U10074 (N_10074,N_9989,N_9619);
nand U10075 (N_10075,N_9532,N_9644);
and U10076 (N_10076,N_9964,N_9655);
nor U10077 (N_10077,N_9553,N_9917);
xor U10078 (N_10078,N_9665,N_9862);
or U10079 (N_10079,N_9668,N_9814);
xor U10080 (N_10080,N_9946,N_9554);
nor U10081 (N_10081,N_9880,N_9690);
nor U10082 (N_10082,N_9750,N_9921);
or U10083 (N_10083,N_9936,N_9693);
or U10084 (N_10084,N_9997,N_9899);
nand U10085 (N_10085,N_9719,N_9737);
nand U10086 (N_10086,N_9920,N_9871);
and U10087 (N_10087,N_9557,N_9609);
and U10088 (N_10088,N_9984,N_9976);
nor U10089 (N_10089,N_9789,N_9539);
xnor U10090 (N_10090,N_9763,N_9639);
xor U10091 (N_10091,N_9999,N_9930);
and U10092 (N_10092,N_9675,N_9974);
nor U10093 (N_10093,N_9878,N_9648);
or U10094 (N_10094,N_9963,N_9610);
xnor U10095 (N_10095,N_9512,N_9773);
or U10096 (N_10096,N_9828,N_9689);
nand U10097 (N_10097,N_9647,N_9962);
xor U10098 (N_10098,N_9673,N_9657);
nand U10099 (N_10099,N_9709,N_9927);
nor U10100 (N_10100,N_9543,N_9783);
xnor U10101 (N_10101,N_9593,N_9861);
nor U10102 (N_10102,N_9596,N_9929);
and U10103 (N_10103,N_9741,N_9734);
and U10104 (N_10104,N_9604,N_9815);
xnor U10105 (N_10105,N_9855,N_9590);
xnor U10106 (N_10106,N_9721,N_9669);
and U10107 (N_10107,N_9867,N_9706);
nor U10108 (N_10108,N_9908,N_9956);
xnor U10109 (N_10109,N_9810,N_9507);
xor U10110 (N_10110,N_9844,N_9827);
and U10111 (N_10111,N_9697,N_9876);
xor U10112 (N_10112,N_9874,N_9835);
or U10113 (N_10113,N_9829,N_9670);
or U10114 (N_10114,N_9755,N_9931);
and U10115 (N_10115,N_9819,N_9684);
or U10116 (N_10116,N_9535,N_9918);
and U10117 (N_10117,N_9872,N_9847);
nand U10118 (N_10118,N_9680,N_9534);
nand U10119 (N_10119,N_9852,N_9991);
nand U10120 (N_10120,N_9615,N_9813);
nor U10121 (N_10121,N_9519,N_9585);
xnor U10122 (N_10122,N_9708,N_9803);
and U10123 (N_10123,N_9801,N_9993);
and U10124 (N_10124,N_9926,N_9900);
xnor U10125 (N_10125,N_9575,N_9983);
nor U10126 (N_10126,N_9517,N_9881);
and U10127 (N_10127,N_9988,N_9700);
nor U10128 (N_10128,N_9546,N_9980);
xnor U10129 (N_10129,N_9795,N_9904);
nand U10130 (N_10130,N_9949,N_9666);
nor U10131 (N_10131,N_9883,N_9940);
xnor U10132 (N_10132,N_9932,N_9743);
and U10133 (N_10133,N_9555,N_9652);
and U10134 (N_10134,N_9618,N_9914);
nor U10135 (N_10135,N_9504,N_9772);
xor U10136 (N_10136,N_9752,N_9839);
xor U10137 (N_10137,N_9837,N_9966);
and U10138 (N_10138,N_9631,N_9831);
nor U10139 (N_10139,N_9663,N_9834);
or U10140 (N_10140,N_9602,N_9617);
or U10141 (N_10141,N_9982,N_9740);
nor U10142 (N_10142,N_9667,N_9758);
nand U10143 (N_10143,N_9569,N_9841);
nor U10144 (N_10144,N_9523,N_9794);
nor U10145 (N_10145,N_9791,N_9865);
nand U10146 (N_10146,N_9778,N_9973);
nand U10147 (N_10147,N_9613,N_9823);
nor U10148 (N_10148,N_9767,N_9705);
nand U10149 (N_10149,N_9968,N_9707);
nor U10150 (N_10150,N_9516,N_9634);
nand U10151 (N_10151,N_9995,N_9661);
and U10152 (N_10152,N_9550,N_9509);
nor U10153 (N_10153,N_9676,N_9774);
nor U10154 (N_10154,N_9888,N_9998);
nor U10155 (N_10155,N_9873,N_9727);
xnor U10156 (N_10156,N_9825,N_9574);
xor U10157 (N_10157,N_9889,N_9687);
xnor U10158 (N_10158,N_9775,N_9712);
nor U10159 (N_10159,N_9784,N_9768);
nor U10160 (N_10160,N_9771,N_9846);
and U10161 (N_10161,N_9748,N_9978);
nor U10162 (N_10162,N_9586,N_9704);
and U10163 (N_10163,N_9522,N_9526);
or U10164 (N_10164,N_9903,N_9560);
or U10165 (N_10165,N_9500,N_9731);
nor U10166 (N_10166,N_9924,N_9797);
nand U10167 (N_10167,N_9662,N_9653);
xor U10168 (N_10168,N_9868,N_9524);
and U10169 (N_10169,N_9542,N_9945);
xnor U10170 (N_10170,N_9625,N_9606);
nor U10171 (N_10171,N_9699,N_9659);
nand U10172 (N_10172,N_9818,N_9503);
nand U10173 (N_10173,N_9816,N_9608);
nor U10174 (N_10174,N_9812,N_9717);
xnor U10175 (N_10175,N_9711,N_9960);
nor U10176 (N_10176,N_9811,N_9722);
nand U10177 (N_10177,N_9714,N_9891);
nand U10178 (N_10178,N_9508,N_9563);
nand U10179 (N_10179,N_9970,N_9892);
nor U10180 (N_10180,N_9702,N_9779);
nor U10181 (N_10181,N_9805,N_9570);
nand U10182 (N_10182,N_9732,N_9875);
nor U10183 (N_10183,N_9558,N_9913);
xnor U10184 (N_10184,N_9979,N_9723);
or U10185 (N_10185,N_9848,N_9780);
or U10186 (N_10186,N_9951,N_9527);
nand U10187 (N_10187,N_9577,N_9958);
nor U10188 (N_10188,N_9877,N_9515);
nor U10189 (N_10189,N_9683,N_9933);
nor U10190 (N_10190,N_9832,N_9660);
nor U10191 (N_10191,N_9580,N_9990);
nor U10192 (N_10192,N_9518,N_9724);
and U10193 (N_10193,N_9573,N_9649);
xnor U10194 (N_10194,N_9870,N_9627);
and U10195 (N_10195,N_9950,N_9584);
nor U10196 (N_10196,N_9901,N_9948);
xnor U10197 (N_10197,N_9583,N_9694);
nand U10198 (N_10198,N_9885,N_9664);
or U10199 (N_10199,N_9749,N_9893);
nand U10200 (N_10200,N_9671,N_9674);
nand U10201 (N_10201,N_9540,N_9894);
nand U10202 (N_10202,N_9592,N_9638);
and U10203 (N_10203,N_9537,N_9836);
or U10204 (N_10204,N_9607,N_9640);
nand U10205 (N_10205,N_9759,N_9777);
nand U10206 (N_10206,N_9857,N_9804);
nand U10207 (N_10207,N_9905,N_9726);
or U10208 (N_10208,N_9603,N_9622);
nor U10209 (N_10209,N_9686,N_9840);
or U10210 (N_10210,N_9942,N_9645);
xor U10211 (N_10211,N_9961,N_9579);
nand U10212 (N_10212,N_9769,N_9568);
nand U10213 (N_10213,N_9672,N_9742);
or U10214 (N_10214,N_9643,N_9786);
xnor U10215 (N_10215,N_9551,N_9971);
nor U10216 (N_10216,N_9808,N_9718);
xnor U10217 (N_10217,N_9843,N_9957);
xor U10218 (N_10218,N_9754,N_9850);
and U10219 (N_10219,N_9788,N_9730);
xnor U10220 (N_10220,N_9616,N_9916);
or U10221 (N_10221,N_9923,N_9745);
nand U10222 (N_10222,N_9594,N_9658);
and U10223 (N_10223,N_9582,N_9587);
and U10224 (N_10224,N_9651,N_9630);
and U10225 (N_10225,N_9677,N_9567);
nand U10226 (N_10226,N_9807,N_9688);
xor U10227 (N_10227,N_9520,N_9826);
xor U10228 (N_10228,N_9678,N_9987);
xnor U10229 (N_10229,N_9505,N_9626);
nand U10230 (N_10230,N_9928,N_9830);
nor U10231 (N_10231,N_9766,N_9809);
xnor U10232 (N_10232,N_9538,N_9802);
xor U10233 (N_10233,N_9614,N_9578);
or U10234 (N_10234,N_9790,N_9656);
and U10235 (N_10235,N_9595,N_9556);
nand U10236 (N_10236,N_9977,N_9735);
xor U10237 (N_10237,N_9739,N_9947);
or U10238 (N_10238,N_9681,N_9838);
nand U10239 (N_10239,N_9911,N_9636);
xnor U10240 (N_10240,N_9565,N_9713);
nand U10241 (N_10241,N_9511,N_9864);
xor U10242 (N_10242,N_9696,N_9564);
or U10243 (N_10243,N_9792,N_9548);
nor U10244 (N_10244,N_9600,N_9912);
or U10245 (N_10245,N_9703,N_9969);
nor U10246 (N_10246,N_9849,N_9937);
nor U10247 (N_10247,N_9642,N_9736);
nor U10248 (N_10248,N_9599,N_9549);
xnor U10249 (N_10249,N_9598,N_9886);
or U10250 (N_10250,N_9660,N_9871);
or U10251 (N_10251,N_9588,N_9536);
nand U10252 (N_10252,N_9888,N_9767);
or U10253 (N_10253,N_9772,N_9537);
or U10254 (N_10254,N_9710,N_9634);
nor U10255 (N_10255,N_9603,N_9642);
nand U10256 (N_10256,N_9663,N_9653);
nor U10257 (N_10257,N_9573,N_9950);
nand U10258 (N_10258,N_9553,N_9974);
or U10259 (N_10259,N_9958,N_9645);
nand U10260 (N_10260,N_9851,N_9768);
or U10261 (N_10261,N_9623,N_9847);
and U10262 (N_10262,N_9572,N_9995);
nand U10263 (N_10263,N_9637,N_9604);
and U10264 (N_10264,N_9644,N_9927);
xnor U10265 (N_10265,N_9507,N_9990);
or U10266 (N_10266,N_9543,N_9789);
nor U10267 (N_10267,N_9602,N_9872);
nor U10268 (N_10268,N_9721,N_9748);
or U10269 (N_10269,N_9894,N_9810);
and U10270 (N_10270,N_9812,N_9897);
xor U10271 (N_10271,N_9671,N_9611);
nor U10272 (N_10272,N_9834,N_9990);
and U10273 (N_10273,N_9707,N_9651);
nor U10274 (N_10274,N_9866,N_9847);
xor U10275 (N_10275,N_9729,N_9781);
nor U10276 (N_10276,N_9676,N_9707);
xor U10277 (N_10277,N_9707,N_9680);
and U10278 (N_10278,N_9726,N_9729);
xnor U10279 (N_10279,N_9593,N_9840);
nor U10280 (N_10280,N_9693,N_9659);
or U10281 (N_10281,N_9593,N_9542);
nor U10282 (N_10282,N_9922,N_9597);
nor U10283 (N_10283,N_9996,N_9932);
nor U10284 (N_10284,N_9786,N_9801);
nand U10285 (N_10285,N_9823,N_9808);
and U10286 (N_10286,N_9991,N_9723);
or U10287 (N_10287,N_9583,N_9979);
or U10288 (N_10288,N_9660,N_9910);
nand U10289 (N_10289,N_9772,N_9888);
nand U10290 (N_10290,N_9875,N_9815);
nand U10291 (N_10291,N_9776,N_9603);
and U10292 (N_10292,N_9764,N_9677);
xor U10293 (N_10293,N_9878,N_9851);
xnor U10294 (N_10294,N_9526,N_9842);
nor U10295 (N_10295,N_9771,N_9704);
and U10296 (N_10296,N_9621,N_9647);
and U10297 (N_10297,N_9807,N_9516);
or U10298 (N_10298,N_9804,N_9768);
nand U10299 (N_10299,N_9665,N_9732);
nor U10300 (N_10300,N_9698,N_9859);
xnor U10301 (N_10301,N_9892,N_9933);
nor U10302 (N_10302,N_9756,N_9809);
nor U10303 (N_10303,N_9685,N_9502);
and U10304 (N_10304,N_9803,N_9580);
nor U10305 (N_10305,N_9721,N_9996);
nand U10306 (N_10306,N_9756,N_9929);
xnor U10307 (N_10307,N_9937,N_9579);
xor U10308 (N_10308,N_9571,N_9921);
or U10309 (N_10309,N_9597,N_9615);
xnor U10310 (N_10310,N_9565,N_9901);
nand U10311 (N_10311,N_9929,N_9748);
and U10312 (N_10312,N_9817,N_9919);
or U10313 (N_10313,N_9633,N_9574);
nor U10314 (N_10314,N_9726,N_9841);
nor U10315 (N_10315,N_9778,N_9823);
or U10316 (N_10316,N_9745,N_9570);
xor U10317 (N_10317,N_9553,N_9717);
xor U10318 (N_10318,N_9903,N_9639);
nor U10319 (N_10319,N_9888,N_9937);
and U10320 (N_10320,N_9533,N_9812);
or U10321 (N_10321,N_9873,N_9591);
xnor U10322 (N_10322,N_9975,N_9817);
or U10323 (N_10323,N_9836,N_9701);
or U10324 (N_10324,N_9566,N_9859);
or U10325 (N_10325,N_9970,N_9812);
or U10326 (N_10326,N_9898,N_9994);
or U10327 (N_10327,N_9844,N_9919);
xor U10328 (N_10328,N_9792,N_9889);
nor U10329 (N_10329,N_9742,N_9707);
or U10330 (N_10330,N_9529,N_9904);
or U10331 (N_10331,N_9784,N_9611);
and U10332 (N_10332,N_9989,N_9645);
nand U10333 (N_10333,N_9569,N_9915);
and U10334 (N_10334,N_9659,N_9771);
and U10335 (N_10335,N_9714,N_9566);
or U10336 (N_10336,N_9519,N_9671);
and U10337 (N_10337,N_9615,N_9900);
or U10338 (N_10338,N_9514,N_9733);
xor U10339 (N_10339,N_9706,N_9638);
and U10340 (N_10340,N_9664,N_9526);
nor U10341 (N_10341,N_9884,N_9506);
and U10342 (N_10342,N_9912,N_9764);
or U10343 (N_10343,N_9769,N_9660);
xor U10344 (N_10344,N_9533,N_9628);
nand U10345 (N_10345,N_9667,N_9815);
and U10346 (N_10346,N_9549,N_9694);
xnor U10347 (N_10347,N_9747,N_9723);
xnor U10348 (N_10348,N_9567,N_9904);
nand U10349 (N_10349,N_9923,N_9894);
and U10350 (N_10350,N_9792,N_9883);
and U10351 (N_10351,N_9898,N_9518);
or U10352 (N_10352,N_9941,N_9564);
and U10353 (N_10353,N_9564,N_9924);
nand U10354 (N_10354,N_9714,N_9536);
and U10355 (N_10355,N_9618,N_9981);
xor U10356 (N_10356,N_9993,N_9538);
and U10357 (N_10357,N_9511,N_9640);
and U10358 (N_10358,N_9568,N_9797);
nand U10359 (N_10359,N_9578,N_9510);
nor U10360 (N_10360,N_9789,N_9607);
and U10361 (N_10361,N_9509,N_9858);
nand U10362 (N_10362,N_9696,N_9582);
nor U10363 (N_10363,N_9502,N_9736);
and U10364 (N_10364,N_9842,N_9691);
xor U10365 (N_10365,N_9827,N_9536);
and U10366 (N_10366,N_9599,N_9627);
and U10367 (N_10367,N_9647,N_9567);
xor U10368 (N_10368,N_9520,N_9796);
xnor U10369 (N_10369,N_9704,N_9805);
or U10370 (N_10370,N_9984,N_9725);
or U10371 (N_10371,N_9504,N_9594);
nor U10372 (N_10372,N_9995,N_9742);
nor U10373 (N_10373,N_9617,N_9955);
and U10374 (N_10374,N_9792,N_9858);
nor U10375 (N_10375,N_9810,N_9502);
nor U10376 (N_10376,N_9581,N_9999);
nand U10377 (N_10377,N_9890,N_9840);
or U10378 (N_10378,N_9588,N_9530);
xor U10379 (N_10379,N_9630,N_9655);
xor U10380 (N_10380,N_9894,N_9723);
nand U10381 (N_10381,N_9762,N_9972);
or U10382 (N_10382,N_9622,N_9816);
and U10383 (N_10383,N_9660,N_9836);
nand U10384 (N_10384,N_9954,N_9955);
xnor U10385 (N_10385,N_9802,N_9940);
or U10386 (N_10386,N_9587,N_9931);
or U10387 (N_10387,N_9617,N_9577);
nand U10388 (N_10388,N_9882,N_9843);
nand U10389 (N_10389,N_9603,N_9778);
nand U10390 (N_10390,N_9979,N_9549);
and U10391 (N_10391,N_9793,N_9852);
nand U10392 (N_10392,N_9670,N_9812);
xor U10393 (N_10393,N_9803,N_9605);
and U10394 (N_10394,N_9500,N_9563);
nor U10395 (N_10395,N_9917,N_9506);
xor U10396 (N_10396,N_9843,N_9628);
nor U10397 (N_10397,N_9724,N_9680);
xnor U10398 (N_10398,N_9838,N_9505);
xor U10399 (N_10399,N_9589,N_9831);
nand U10400 (N_10400,N_9581,N_9730);
or U10401 (N_10401,N_9829,N_9996);
or U10402 (N_10402,N_9631,N_9510);
nand U10403 (N_10403,N_9935,N_9554);
xnor U10404 (N_10404,N_9757,N_9649);
or U10405 (N_10405,N_9543,N_9622);
and U10406 (N_10406,N_9610,N_9611);
and U10407 (N_10407,N_9644,N_9718);
xor U10408 (N_10408,N_9917,N_9759);
nand U10409 (N_10409,N_9593,N_9762);
or U10410 (N_10410,N_9851,N_9509);
nand U10411 (N_10411,N_9852,N_9726);
nand U10412 (N_10412,N_9527,N_9931);
nor U10413 (N_10413,N_9967,N_9807);
nor U10414 (N_10414,N_9968,N_9637);
nor U10415 (N_10415,N_9504,N_9668);
and U10416 (N_10416,N_9774,N_9930);
and U10417 (N_10417,N_9533,N_9782);
nor U10418 (N_10418,N_9636,N_9986);
nand U10419 (N_10419,N_9956,N_9827);
or U10420 (N_10420,N_9997,N_9514);
and U10421 (N_10421,N_9646,N_9836);
or U10422 (N_10422,N_9759,N_9738);
nor U10423 (N_10423,N_9987,N_9791);
and U10424 (N_10424,N_9725,N_9776);
nand U10425 (N_10425,N_9541,N_9683);
nor U10426 (N_10426,N_9670,N_9533);
and U10427 (N_10427,N_9818,N_9555);
nor U10428 (N_10428,N_9813,N_9649);
xnor U10429 (N_10429,N_9770,N_9547);
or U10430 (N_10430,N_9749,N_9713);
xnor U10431 (N_10431,N_9791,N_9906);
nor U10432 (N_10432,N_9721,N_9838);
or U10433 (N_10433,N_9877,N_9783);
and U10434 (N_10434,N_9908,N_9933);
nand U10435 (N_10435,N_9580,N_9512);
nand U10436 (N_10436,N_9642,N_9918);
and U10437 (N_10437,N_9988,N_9841);
or U10438 (N_10438,N_9947,N_9684);
or U10439 (N_10439,N_9740,N_9811);
nor U10440 (N_10440,N_9930,N_9994);
and U10441 (N_10441,N_9725,N_9505);
nor U10442 (N_10442,N_9937,N_9936);
nand U10443 (N_10443,N_9854,N_9513);
nor U10444 (N_10444,N_9653,N_9973);
and U10445 (N_10445,N_9506,N_9599);
xnor U10446 (N_10446,N_9935,N_9807);
nor U10447 (N_10447,N_9878,N_9748);
nand U10448 (N_10448,N_9733,N_9545);
nand U10449 (N_10449,N_9740,N_9664);
nand U10450 (N_10450,N_9693,N_9760);
xnor U10451 (N_10451,N_9807,N_9661);
xnor U10452 (N_10452,N_9581,N_9941);
nor U10453 (N_10453,N_9760,N_9858);
and U10454 (N_10454,N_9571,N_9845);
xor U10455 (N_10455,N_9989,N_9597);
xor U10456 (N_10456,N_9949,N_9706);
xnor U10457 (N_10457,N_9794,N_9566);
nand U10458 (N_10458,N_9728,N_9909);
xnor U10459 (N_10459,N_9702,N_9546);
nand U10460 (N_10460,N_9873,N_9560);
and U10461 (N_10461,N_9669,N_9946);
nand U10462 (N_10462,N_9760,N_9712);
nand U10463 (N_10463,N_9814,N_9892);
xor U10464 (N_10464,N_9615,N_9592);
or U10465 (N_10465,N_9995,N_9741);
nor U10466 (N_10466,N_9955,N_9997);
or U10467 (N_10467,N_9712,N_9797);
nand U10468 (N_10468,N_9862,N_9956);
nand U10469 (N_10469,N_9534,N_9508);
xnor U10470 (N_10470,N_9731,N_9895);
or U10471 (N_10471,N_9866,N_9604);
nand U10472 (N_10472,N_9793,N_9526);
and U10473 (N_10473,N_9907,N_9999);
and U10474 (N_10474,N_9700,N_9961);
xnor U10475 (N_10475,N_9816,N_9512);
xnor U10476 (N_10476,N_9847,N_9833);
xor U10477 (N_10477,N_9878,N_9573);
and U10478 (N_10478,N_9629,N_9710);
xor U10479 (N_10479,N_9578,N_9819);
nor U10480 (N_10480,N_9781,N_9542);
nand U10481 (N_10481,N_9806,N_9867);
xnor U10482 (N_10482,N_9634,N_9753);
or U10483 (N_10483,N_9807,N_9868);
or U10484 (N_10484,N_9542,N_9983);
nor U10485 (N_10485,N_9524,N_9659);
nor U10486 (N_10486,N_9698,N_9520);
xnor U10487 (N_10487,N_9956,N_9838);
or U10488 (N_10488,N_9723,N_9546);
and U10489 (N_10489,N_9514,N_9820);
or U10490 (N_10490,N_9616,N_9728);
nor U10491 (N_10491,N_9891,N_9779);
nand U10492 (N_10492,N_9942,N_9973);
nor U10493 (N_10493,N_9676,N_9954);
xor U10494 (N_10494,N_9976,N_9626);
or U10495 (N_10495,N_9855,N_9691);
or U10496 (N_10496,N_9558,N_9600);
nor U10497 (N_10497,N_9740,N_9866);
or U10498 (N_10498,N_9934,N_9838);
nor U10499 (N_10499,N_9602,N_9893);
xor U10500 (N_10500,N_10124,N_10052);
and U10501 (N_10501,N_10484,N_10156);
nand U10502 (N_10502,N_10424,N_10045);
nand U10503 (N_10503,N_10090,N_10064);
or U10504 (N_10504,N_10425,N_10269);
nand U10505 (N_10505,N_10204,N_10494);
nand U10506 (N_10506,N_10070,N_10341);
and U10507 (N_10507,N_10397,N_10063);
nand U10508 (N_10508,N_10366,N_10214);
and U10509 (N_10509,N_10266,N_10228);
and U10510 (N_10510,N_10237,N_10039);
nor U10511 (N_10511,N_10056,N_10413);
xor U10512 (N_10512,N_10312,N_10187);
xnor U10513 (N_10513,N_10234,N_10114);
nand U10514 (N_10514,N_10270,N_10203);
or U10515 (N_10515,N_10351,N_10272);
nor U10516 (N_10516,N_10206,N_10191);
xnor U10517 (N_10517,N_10025,N_10365);
nor U10518 (N_10518,N_10033,N_10073);
nor U10519 (N_10519,N_10222,N_10327);
xnor U10520 (N_10520,N_10078,N_10288);
nand U10521 (N_10521,N_10490,N_10043);
nor U10522 (N_10522,N_10473,N_10445);
xnor U10523 (N_10523,N_10480,N_10182);
nor U10524 (N_10524,N_10251,N_10162);
xnor U10525 (N_10525,N_10136,N_10155);
and U10526 (N_10526,N_10326,N_10008);
and U10527 (N_10527,N_10210,N_10364);
or U10528 (N_10528,N_10497,N_10194);
nand U10529 (N_10529,N_10159,N_10409);
xor U10530 (N_10530,N_10379,N_10456);
nor U10531 (N_10531,N_10154,N_10051);
nor U10532 (N_10532,N_10392,N_10329);
nor U10533 (N_10533,N_10355,N_10450);
and U10534 (N_10534,N_10447,N_10461);
and U10535 (N_10535,N_10097,N_10346);
nor U10536 (N_10536,N_10429,N_10278);
nor U10537 (N_10537,N_10440,N_10075);
and U10538 (N_10538,N_10492,N_10230);
nand U10539 (N_10539,N_10127,N_10290);
or U10540 (N_10540,N_10112,N_10174);
or U10541 (N_10541,N_10350,N_10000);
nand U10542 (N_10542,N_10475,N_10274);
nor U10543 (N_10543,N_10465,N_10010);
and U10544 (N_10544,N_10486,N_10438);
xnor U10545 (N_10545,N_10152,N_10171);
xnor U10546 (N_10546,N_10232,N_10306);
or U10547 (N_10547,N_10246,N_10106);
nor U10548 (N_10548,N_10004,N_10360);
and U10549 (N_10549,N_10087,N_10400);
xnor U10550 (N_10550,N_10128,N_10249);
nor U10551 (N_10551,N_10307,N_10011);
and U10552 (N_10552,N_10368,N_10195);
or U10553 (N_10553,N_10394,N_10250);
nor U10554 (N_10554,N_10021,N_10105);
nand U10555 (N_10555,N_10479,N_10079);
or U10556 (N_10556,N_10081,N_10017);
nand U10557 (N_10557,N_10121,N_10319);
xor U10558 (N_10558,N_10100,N_10036);
nand U10559 (N_10559,N_10188,N_10263);
nor U10560 (N_10560,N_10374,N_10476);
nor U10561 (N_10561,N_10295,N_10068);
nor U10562 (N_10562,N_10356,N_10323);
or U10563 (N_10563,N_10134,N_10453);
and U10564 (N_10564,N_10072,N_10089);
xnor U10565 (N_10565,N_10333,N_10047);
or U10566 (N_10566,N_10287,N_10189);
nor U10567 (N_10567,N_10102,N_10432);
and U10568 (N_10568,N_10111,N_10357);
nor U10569 (N_10569,N_10371,N_10145);
nor U10570 (N_10570,N_10197,N_10150);
xor U10571 (N_10571,N_10183,N_10303);
xnor U10572 (N_10572,N_10018,N_10255);
and U10573 (N_10573,N_10361,N_10498);
nand U10574 (N_10574,N_10173,N_10190);
nand U10575 (N_10575,N_10338,N_10388);
nand U10576 (N_10576,N_10221,N_10029);
xor U10577 (N_10577,N_10141,N_10259);
nor U10578 (N_10578,N_10207,N_10393);
nand U10579 (N_10579,N_10403,N_10436);
nor U10580 (N_10580,N_10344,N_10448);
or U10581 (N_10581,N_10140,N_10095);
xor U10582 (N_10582,N_10225,N_10254);
nor U10583 (N_10583,N_10318,N_10378);
and U10584 (N_10584,N_10220,N_10466);
nand U10585 (N_10585,N_10468,N_10455);
and U10586 (N_10586,N_10314,N_10199);
nand U10587 (N_10587,N_10442,N_10014);
xor U10588 (N_10588,N_10340,N_10116);
or U10589 (N_10589,N_10229,N_10399);
or U10590 (N_10590,N_10441,N_10275);
xor U10591 (N_10591,N_10477,N_10370);
nor U10592 (N_10592,N_10024,N_10418);
and U10593 (N_10593,N_10027,N_10235);
xor U10594 (N_10594,N_10264,N_10049);
nand U10595 (N_10595,N_10324,N_10420);
nand U10596 (N_10596,N_10335,N_10139);
nand U10597 (N_10597,N_10493,N_10164);
or U10598 (N_10598,N_10451,N_10163);
xnor U10599 (N_10599,N_10175,N_10491);
or U10600 (N_10600,N_10135,N_10439);
or U10601 (N_10601,N_10218,N_10099);
xor U10602 (N_10602,N_10454,N_10130);
or U10603 (N_10603,N_10240,N_10487);
nor U10604 (N_10604,N_10489,N_10458);
and U10605 (N_10605,N_10305,N_10169);
nand U10606 (N_10606,N_10311,N_10209);
and U10607 (N_10607,N_10343,N_10321);
and U10608 (N_10608,N_10383,N_10345);
nand U10609 (N_10609,N_10098,N_10302);
nor U10610 (N_10610,N_10241,N_10469);
nand U10611 (N_10611,N_10339,N_10108);
or U10612 (N_10612,N_10067,N_10396);
xor U10613 (N_10613,N_10336,N_10196);
and U10614 (N_10614,N_10459,N_10062);
xnor U10615 (N_10615,N_10386,N_10488);
or U10616 (N_10616,N_10283,N_10299);
and U10617 (N_10617,N_10030,N_10382);
and U10618 (N_10618,N_10224,N_10349);
or U10619 (N_10619,N_10271,N_10300);
or U10620 (N_10620,N_10212,N_10103);
nor U10621 (N_10621,N_10082,N_10119);
and U10622 (N_10622,N_10227,N_10367);
nor U10623 (N_10623,N_10353,N_10244);
nand U10624 (N_10624,N_10320,N_10423);
or U10625 (N_10625,N_10474,N_10422);
or U10626 (N_10626,N_10092,N_10058);
nor U10627 (N_10627,N_10467,N_10178);
or U10628 (N_10628,N_10007,N_10342);
and U10629 (N_10629,N_10015,N_10471);
nand U10630 (N_10630,N_10460,N_10464);
nor U10631 (N_10631,N_10462,N_10020);
xnor U10632 (N_10632,N_10296,N_10416);
nand U10633 (N_10633,N_10291,N_10219);
nor U10634 (N_10634,N_10284,N_10470);
or U10635 (N_10635,N_10138,N_10006);
nor U10636 (N_10636,N_10358,N_10482);
nand U10637 (N_10637,N_10449,N_10446);
or U10638 (N_10638,N_10405,N_10410);
or U10639 (N_10639,N_10042,N_10258);
xnor U10640 (N_10640,N_10304,N_10301);
nor U10641 (N_10641,N_10028,N_10261);
or U10642 (N_10642,N_10481,N_10016);
xor U10643 (N_10643,N_10093,N_10050);
xor U10644 (N_10644,N_10292,N_10389);
or U10645 (N_10645,N_10213,N_10337);
or U10646 (N_10646,N_10120,N_10208);
xor U10647 (N_10647,N_10402,N_10243);
nand U10648 (N_10648,N_10122,N_10427);
and U10649 (N_10649,N_10217,N_10252);
or U10650 (N_10650,N_10023,N_10401);
xor U10651 (N_10651,N_10236,N_10363);
and U10652 (N_10652,N_10348,N_10347);
xnor U10653 (N_10653,N_10430,N_10012);
nand U10654 (N_10654,N_10282,N_10273);
nor U10655 (N_10655,N_10309,N_10168);
or U10656 (N_10656,N_10009,N_10077);
and U10657 (N_10657,N_10066,N_10317);
nand U10658 (N_10658,N_10391,N_10123);
nor U10659 (N_10659,N_10279,N_10071);
or U10660 (N_10660,N_10125,N_10180);
nor U10661 (N_10661,N_10257,N_10026);
xnor U10662 (N_10662,N_10463,N_10385);
xor U10663 (N_10663,N_10238,N_10242);
xnor U10664 (N_10664,N_10046,N_10001);
nand U10665 (N_10665,N_10256,N_10352);
nor U10666 (N_10666,N_10297,N_10215);
xnor U10667 (N_10667,N_10267,N_10472);
nand U10668 (N_10668,N_10193,N_10177);
nor U10669 (N_10669,N_10104,N_10115);
nand U10670 (N_10670,N_10133,N_10496);
and U10671 (N_10671,N_10426,N_10041);
nand U10672 (N_10672,N_10005,N_10076);
and U10673 (N_10673,N_10437,N_10315);
nor U10674 (N_10674,N_10457,N_10354);
and U10675 (N_10675,N_10406,N_10216);
nand U10676 (N_10676,N_10268,N_10404);
and U10677 (N_10677,N_10185,N_10146);
nand U10678 (N_10678,N_10143,N_10048);
nand U10679 (N_10679,N_10057,N_10372);
or U10680 (N_10680,N_10415,N_10031);
nor U10681 (N_10681,N_10265,N_10144);
xor U10682 (N_10682,N_10132,N_10359);
nand U10683 (N_10683,N_10091,N_10147);
nand U10684 (N_10684,N_10433,N_10094);
nor U10685 (N_10685,N_10142,N_10316);
or U10686 (N_10686,N_10172,N_10153);
nand U10687 (N_10687,N_10157,N_10044);
xor U10688 (N_10688,N_10186,N_10381);
or U10689 (N_10689,N_10126,N_10131);
nand U10690 (N_10690,N_10285,N_10298);
xnor U10691 (N_10691,N_10444,N_10205);
xnor U10692 (N_10692,N_10239,N_10330);
and U10693 (N_10693,N_10084,N_10003);
xnor U10694 (N_10694,N_10331,N_10165);
or U10695 (N_10695,N_10248,N_10109);
and U10696 (N_10696,N_10040,N_10149);
and U10697 (N_10697,N_10101,N_10167);
nand U10698 (N_10698,N_10431,N_10308);
and U10699 (N_10699,N_10034,N_10198);
nand U10700 (N_10700,N_10060,N_10384);
or U10701 (N_10701,N_10158,N_10074);
nor U10702 (N_10702,N_10377,N_10485);
and U10703 (N_10703,N_10211,N_10019);
or U10704 (N_10704,N_10038,N_10176);
and U10705 (N_10705,N_10032,N_10233);
and U10706 (N_10706,N_10061,N_10037);
and U10707 (N_10707,N_10247,N_10055);
xnor U10708 (N_10708,N_10398,N_10054);
nor U10709 (N_10709,N_10478,N_10151);
nand U10710 (N_10710,N_10110,N_10226);
nand U10711 (N_10711,N_10161,N_10086);
or U10712 (N_10712,N_10260,N_10408);
or U10713 (N_10713,N_10277,N_10387);
xor U10714 (N_10714,N_10452,N_10421);
nor U10715 (N_10715,N_10313,N_10499);
nor U10716 (N_10716,N_10322,N_10419);
nand U10717 (N_10717,N_10411,N_10376);
xnor U10718 (N_10718,N_10231,N_10148);
nor U10719 (N_10719,N_10117,N_10276);
xnor U10720 (N_10720,N_10129,N_10435);
xnor U10721 (N_10721,N_10407,N_10080);
nor U10722 (N_10722,N_10380,N_10083);
or U10723 (N_10723,N_10373,N_10443);
and U10724 (N_10724,N_10310,N_10395);
nor U10725 (N_10725,N_10262,N_10088);
xnor U10726 (N_10726,N_10059,N_10085);
and U10727 (N_10727,N_10184,N_10483);
or U10728 (N_10728,N_10166,N_10202);
or U10729 (N_10729,N_10428,N_10495);
and U10730 (N_10730,N_10200,N_10096);
nor U10731 (N_10731,N_10118,N_10412);
or U10732 (N_10732,N_10417,N_10281);
nor U10733 (N_10733,N_10053,N_10294);
nand U10734 (N_10734,N_10362,N_10179);
or U10735 (N_10735,N_10434,N_10002);
nand U10736 (N_10736,N_10334,N_10181);
nand U10737 (N_10737,N_10035,N_10223);
xnor U10738 (N_10738,N_10328,N_10065);
xnor U10739 (N_10739,N_10332,N_10013);
or U10740 (N_10740,N_10022,N_10069);
and U10741 (N_10741,N_10293,N_10192);
and U10742 (N_10742,N_10375,N_10280);
and U10743 (N_10743,N_10201,N_10289);
or U10744 (N_10744,N_10253,N_10369);
xor U10745 (N_10745,N_10137,N_10414);
nand U10746 (N_10746,N_10113,N_10286);
nand U10747 (N_10747,N_10325,N_10160);
xnor U10748 (N_10748,N_10390,N_10245);
and U10749 (N_10749,N_10170,N_10107);
xnor U10750 (N_10750,N_10242,N_10266);
nor U10751 (N_10751,N_10003,N_10329);
xnor U10752 (N_10752,N_10051,N_10174);
nand U10753 (N_10753,N_10051,N_10396);
nand U10754 (N_10754,N_10047,N_10403);
nand U10755 (N_10755,N_10082,N_10368);
and U10756 (N_10756,N_10305,N_10042);
and U10757 (N_10757,N_10130,N_10062);
nor U10758 (N_10758,N_10425,N_10453);
or U10759 (N_10759,N_10316,N_10215);
and U10760 (N_10760,N_10433,N_10303);
xnor U10761 (N_10761,N_10157,N_10244);
or U10762 (N_10762,N_10202,N_10147);
nand U10763 (N_10763,N_10415,N_10417);
or U10764 (N_10764,N_10091,N_10483);
xor U10765 (N_10765,N_10449,N_10254);
xnor U10766 (N_10766,N_10310,N_10088);
or U10767 (N_10767,N_10334,N_10027);
xor U10768 (N_10768,N_10037,N_10462);
xnor U10769 (N_10769,N_10296,N_10010);
nand U10770 (N_10770,N_10132,N_10377);
or U10771 (N_10771,N_10191,N_10379);
xnor U10772 (N_10772,N_10302,N_10430);
nand U10773 (N_10773,N_10186,N_10008);
or U10774 (N_10774,N_10388,N_10458);
xor U10775 (N_10775,N_10070,N_10348);
and U10776 (N_10776,N_10122,N_10177);
nand U10777 (N_10777,N_10293,N_10142);
and U10778 (N_10778,N_10227,N_10313);
and U10779 (N_10779,N_10048,N_10331);
and U10780 (N_10780,N_10089,N_10405);
xnor U10781 (N_10781,N_10302,N_10014);
nand U10782 (N_10782,N_10164,N_10258);
nand U10783 (N_10783,N_10306,N_10065);
or U10784 (N_10784,N_10056,N_10357);
nand U10785 (N_10785,N_10492,N_10392);
or U10786 (N_10786,N_10331,N_10181);
nand U10787 (N_10787,N_10114,N_10360);
nor U10788 (N_10788,N_10148,N_10059);
nand U10789 (N_10789,N_10210,N_10321);
and U10790 (N_10790,N_10228,N_10157);
or U10791 (N_10791,N_10462,N_10372);
and U10792 (N_10792,N_10249,N_10452);
xor U10793 (N_10793,N_10218,N_10224);
xor U10794 (N_10794,N_10376,N_10378);
nand U10795 (N_10795,N_10312,N_10461);
nor U10796 (N_10796,N_10355,N_10280);
xnor U10797 (N_10797,N_10340,N_10211);
xnor U10798 (N_10798,N_10228,N_10192);
or U10799 (N_10799,N_10197,N_10371);
and U10800 (N_10800,N_10210,N_10347);
or U10801 (N_10801,N_10281,N_10095);
nand U10802 (N_10802,N_10052,N_10159);
nor U10803 (N_10803,N_10369,N_10038);
nor U10804 (N_10804,N_10112,N_10416);
xor U10805 (N_10805,N_10330,N_10315);
and U10806 (N_10806,N_10058,N_10114);
nand U10807 (N_10807,N_10164,N_10252);
nor U10808 (N_10808,N_10126,N_10385);
or U10809 (N_10809,N_10159,N_10492);
and U10810 (N_10810,N_10398,N_10492);
xor U10811 (N_10811,N_10273,N_10122);
or U10812 (N_10812,N_10133,N_10403);
nand U10813 (N_10813,N_10114,N_10244);
nor U10814 (N_10814,N_10180,N_10114);
or U10815 (N_10815,N_10448,N_10159);
xnor U10816 (N_10816,N_10106,N_10242);
or U10817 (N_10817,N_10158,N_10327);
xnor U10818 (N_10818,N_10099,N_10260);
nand U10819 (N_10819,N_10329,N_10391);
or U10820 (N_10820,N_10463,N_10411);
xnor U10821 (N_10821,N_10109,N_10392);
and U10822 (N_10822,N_10154,N_10024);
nor U10823 (N_10823,N_10037,N_10333);
or U10824 (N_10824,N_10051,N_10435);
nand U10825 (N_10825,N_10260,N_10391);
nor U10826 (N_10826,N_10111,N_10085);
or U10827 (N_10827,N_10486,N_10068);
xor U10828 (N_10828,N_10101,N_10219);
and U10829 (N_10829,N_10461,N_10008);
and U10830 (N_10830,N_10488,N_10114);
or U10831 (N_10831,N_10364,N_10341);
nand U10832 (N_10832,N_10300,N_10214);
nand U10833 (N_10833,N_10447,N_10006);
xnor U10834 (N_10834,N_10459,N_10466);
nand U10835 (N_10835,N_10499,N_10030);
and U10836 (N_10836,N_10462,N_10403);
nand U10837 (N_10837,N_10215,N_10303);
xnor U10838 (N_10838,N_10402,N_10248);
xor U10839 (N_10839,N_10307,N_10236);
nand U10840 (N_10840,N_10161,N_10241);
xnor U10841 (N_10841,N_10263,N_10459);
and U10842 (N_10842,N_10185,N_10175);
and U10843 (N_10843,N_10457,N_10224);
xor U10844 (N_10844,N_10041,N_10497);
xnor U10845 (N_10845,N_10384,N_10125);
nor U10846 (N_10846,N_10336,N_10115);
xnor U10847 (N_10847,N_10352,N_10306);
or U10848 (N_10848,N_10006,N_10408);
or U10849 (N_10849,N_10361,N_10268);
nor U10850 (N_10850,N_10441,N_10470);
or U10851 (N_10851,N_10035,N_10084);
nor U10852 (N_10852,N_10363,N_10060);
nand U10853 (N_10853,N_10040,N_10236);
and U10854 (N_10854,N_10099,N_10216);
or U10855 (N_10855,N_10292,N_10062);
nand U10856 (N_10856,N_10256,N_10051);
nor U10857 (N_10857,N_10344,N_10481);
and U10858 (N_10858,N_10015,N_10027);
and U10859 (N_10859,N_10318,N_10163);
nand U10860 (N_10860,N_10016,N_10208);
nor U10861 (N_10861,N_10146,N_10426);
xnor U10862 (N_10862,N_10080,N_10276);
and U10863 (N_10863,N_10229,N_10081);
nand U10864 (N_10864,N_10456,N_10237);
nand U10865 (N_10865,N_10028,N_10451);
xor U10866 (N_10866,N_10168,N_10076);
nand U10867 (N_10867,N_10139,N_10004);
nand U10868 (N_10868,N_10409,N_10078);
or U10869 (N_10869,N_10230,N_10244);
xor U10870 (N_10870,N_10150,N_10286);
xor U10871 (N_10871,N_10009,N_10239);
or U10872 (N_10872,N_10036,N_10436);
xnor U10873 (N_10873,N_10497,N_10478);
and U10874 (N_10874,N_10030,N_10059);
nor U10875 (N_10875,N_10220,N_10182);
xnor U10876 (N_10876,N_10363,N_10201);
nand U10877 (N_10877,N_10491,N_10127);
and U10878 (N_10878,N_10077,N_10225);
nor U10879 (N_10879,N_10151,N_10119);
and U10880 (N_10880,N_10425,N_10159);
nand U10881 (N_10881,N_10296,N_10152);
or U10882 (N_10882,N_10064,N_10442);
xor U10883 (N_10883,N_10312,N_10108);
and U10884 (N_10884,N_10349,N_10468);
nand U10885 (N_10885,N_10086,N_10182);
and U10886 (N_10886,N_10187,N_10258);
nand U10887 (N_10887,N_10466,N_10245);
or U10888 (N_10888,N_10423,N_10178);
nand U10889 (N_10889,N_10015,N_10331);
nand U10890 (N_10890,N_10012,N_10450);
and U10891 (N_10891,N_10339,N_10020);
nand U10892 (N_10892,N_10371,N_10455);
or U10893 (N_10893,N_10189,N_10255);
xnor U10894 (N_10894,N_10134,N_10350);
and U10895 (N_10895,N_10237,N_10403);
xnor U10896 (N_10896,N_10432,N_10215);
nor U10897 (N_10897,N_10130,N_10174);
xnor U10898 (N_10898,N_10482,N_10198);
and U10899 (N_10899,N_10404,N_10060);
xor U10900 (N_10900,N_10326,N_10027);
or U10901 (N_10901,N_10341,N_10164);
xnor U10902 (N_10902,N_10065,N_10485);
and U10903 (N_10903,N_10291,N_10210);
or U10904 (N_10904,N_10164,N_10181);
and U10905 (N_10905,N_10056,N_10289);
nand U10906 (N_10906,N_10284,N_10296);
xor U10907 (N_10907,N_10268,N_10121);
nand U10908 (N_10908,N_10046,N_10493);
and U10909 (N_10909,N_10204,N_10449);
nand U10910 (N_10910,N_10257,N_10158);
xnor U10911 (N_10911,N_10110,N_10314);
nand U10912 (N_10912,N_10297,N_10423);
xnor U10913 (N_10913,N_10333,N_10249);
nor U10914 (N_10914,N_10162,N_10007);
xnor U10915 (N_10915,N_10289,N_10386);
nand U10916 (N_10916,N_10355,N_10164);
xnor U10917 (N_10917,N_10035,N_10243);
xnor U10918 (N_10918,N_10313,N_10058);
or U10919 (N_10919,N_10143,N_10061);
or U10920 (N_10920,N_10151,N_10321);
xnor U10921 (N_10921,N_10059,N_10152);
nand U10922 (N_10922,N_10284,N_10293);
nor U10923 (N_10923,N_10259,N_10393);
or U10924 (N_10924,N_10340,N_10139);
nand U10925 (N_10925,N_10134,N_10364);
nand U10926 (N_10926,N_10081,N_10398);
or U10927 (N_10927,N_10014,N_10311);
nand U10928 (N_10928,N_10128,N_10063);
or U10929 (N_10929,N_10074,N_10421);
nor U10930 (N_10930,N_10148,N_10154);
xor U10931 (N_10931,N_10093,N_10081);
or U10932 (N_10932,N_10071,N_10000);
xnor U10933 (N_10933,N_10167,N_10383);
xor U10934 (N_10934,N_10292,N_10230);
xor U10935 (N_10935,N_10154,N_10249);
nand U10936 (N_10936,N_10052,N_10267);
or U10937 (N_10937,N_10150,N_10217);
and U10938 (N_10938,N_10087,N_10425);
or U10939 (N_10939,N_10484,N_10193);
nand U10940 (N_10940,N_10296,N_10125);
xor U10941 (N_10941,N_10148,N_10220);
nand U10942 (N_10942,N_10062,N_10226);
or U10943 (N_10943,N_10331,N_10019);
and U10944 (N_10944,N_10341,N_10382);
nand U10945 (N_10945,N_10228,N_10410);
xor U10946 (N_10946,N_10000,N_10222);
nor U10947 (N_10947,N_10128,N_10357);
xor U10948 (N_10948,N_10295,N_10167);
nor U10949 (N_10949,N_10279,N_10148);
xor U10950 (N_10950,N_10153,N_10102);
xor U10951 (N_10951,N_10012,N_10401);
xor U10952 (N_10952,N_10496,N_10011);
and U10953 (N_10953,N_10396,N_10461);
nor U10954 (N_10954,N_10371,N_10378);
or U10955 (N_10955,N_10454,N_10435);
nor U10956 (N_10956,N_10040,N_10112);
xor U10957 (N_10957,N_10167,N_10156);
or U10958 (N_10958,N_10203,N_10227);
nor U10959 (N_10959,N_10487,N_10275);
nand U10960 (N_10960,N_10353,N_10417);
nand U10961 (N_10961,N_10438,N_10249);
nor U10962 (N_10962,N_10351,N_10167);
or U10963 (N_10963,N_10131,N_10113);
nand U10964 (N_10964,N_10345,N_10159);
xor U10965 (N_10965,N_10258,N_10143);
xnor U10966 (N_10966,N_10043,N_10337);
or U10967 (N_10967,N_10138,N_10247);
xnor U10968 (N_10968,N_10272,N_10038);
xnor U10969 (N_10969,N_10234,N_10257);
and U10970 (N_10970,N_10434,N_10166);
and U10971 (N_10971,N_10423,N_10395);
nor U10972 (N_10972,N_10108,N_10179);
or U10973 (N_10973,N_10169,N_10337);
nor U10974 (N_10974,N_10400,N_10479);
and U10975 (N_10975,N_10067,N_10252);
and U10976 (N_10976,N_10486,N_10192);
and U10977 (N_10977,N_10231,N_10103);
nand U10978 (N_10978,N_10198,N_10249);
nand U10979 (N_10979,N_10458,N_10252);
and U10980 (N_10980,N_10466,N_10171);
xor U10981 (N_10981,N_10294,N_10264);
or U10982 (N_10982,N_10320,N_10380);
and U10983 (N_10983,N_10033,N_10184);
or U10984 (N_10984,N_10124,N_10092);
nor U10985 (N_10985,N_10433,N_10279);
or U10986 (N_10986,N_10366,N_10217);
nand U10987 (N_10987,N_10358,N_10363);
and U10988 (N_10988,N_10369,N_10068);
and U10989 (N_10989,N_10212,N_10418);
nand U10990 (N_10990,N_10116,N_10143);
nand U10991 (N_10991,N_10334,N_10242);
nand U10992 (N_10992,N_10129,N_10023);
and U10993 (N_10993,N_10182,N_10332);
or U10994 (N_10994,N_10330,N_10234);
and U10995 (N_10995,N_10048,N_10098);
nand U10996 (N_10996,N_10116,N_10002);
nand U10997 (N_10997,N_10003,N_10220);
or U10998 (N_10998,N_10469,N_10111);
nand U10999 (N_10999,N_10063,N_10214);
nor U11000 (N_11000,N_10859,N_10727);
nor U11001 (N_11001,N_10886,N_10583);
nand U11002 (N_11002,N_10789,N_10599);
and U11003 (N_11003,N_10629,N_10742);
nand U11004 (N_11004,N_10720,N_10885);
xnor U11005 (N_11005,N_10970,N_10768);
nand U11006 (N_11006,N_10525,N_10581);
xnor U11007 (N_11007,N_10516,N_10878);
nand U11008 (N_11008,N_10526,N_10632);
nor U11009 (N_11009,N_10941,N_10823);
and U11010 (N_11010,N_10557,N_10853);
or U11011 (N_11011,N_10820,N_10567);
xor U11012 (N_11012,N_10999,N_10961);
xnor U11013 (N_11013,N_10685,N_10834);
and U11014 (N_11014,N_10739,N_10741);
nor U11015 (N_11015,N_10986,N_10717);
and U11016 (N_11016,N_10817,N_10712);
nor U11017 (N_11017,N_10625,N_10651);
nand U11018 (N_11018,N_10579,N_10566);
xor U11019 (N_11019,N_10863,N_10860);
xor U11020 (N_11020,N_10657,N_10641);
and U11021 (N_11021,N_10618,N_10934);
xnor U11022 (N_11022,N_10563,N_10888);
or U11023 (N_11023,N_10938,N_10591);
xor U11024 (N_11024,N_10541,N_10907);
or U11025 (N_11025,N_10679,N_10848);
nand U11026 (N_11026,N_10946,N_10622);
or U11027 (N_11027,N_10723,N_10792);
nor U11028 (N_11028,N_10812,N_10835);
nand U11029 (N_11029,N_10913,N_10626);
or U11030 (N_11030,N_10613,N_10537);
xor U11031 (N_11031,N_10511,N_10695);
nand U11032 (N_11032,N_10915,N_10957);
nor U11033 (N_11033,N_10936,N_10677);
xnor U11034 (N_11034,N_10620,N_10642);
xnor U11035 (N_11035,N_10771,N_10652);
and U11036 (N_11036,N_10507,N_10821);
xnor U11037 (N_11037,N_10929,N_10730);
and U11038 (N_11038,N_10933,N_10655);
nand U11039 (N_11039,N_10521,N_10518);
nor U11040 (N_11040,N_10875,N_10752);
nor U11041 (N_11041,N_10676,N_10952);
and U11042 (N_11042,N_10932,N_10906);
nand U11043 (N_11043,N_10611,N_10945);
and U11044 (N_11044,N_10761,N_10992);
nand U11045 (N_11045,N_10773,N_10724);
or U11046 (N_11046,N_10635,N_10740);
xnor U11047 (N_11047,N_10964,N_10816);
nand U11048 (N_11048,N_10889,N_10683);
or U11049 (N_11049,N_10791,N_10598);
nand U11050 (N_11050,N_10953,N_10813);
nor U11051 (N_11051,N_10686,N_10593);
xor U11052 (N_11052,N_10989,N_10726);
and U11053 (N_11053,N_10700,N_10621);
xnor U11054 (N_11054,N_10770,N_10993);
nand U11055 (N_11055,N_10732,N_10956);
nor U11056 (N_11056,N_10671,N_10841);
nor U11057 (N_11057,N_10803,N_10614);
or U11058 (N_11058,N_10856,N_10669);
nand U11059 (N_11059,N_10766,N_10610);
or U11060 (N_11060,N_10763,N_10509);
or U11061 (N_11061,N_10811,N_10561);
or U11062 (N_11062,N_10777,N_10751);
nor U11063 (N_11063,N_10833,N_10728);
nand U11064 (N_11064,N_10678,N_10680);
xnor U11065 (N_11065,N_10667,N_10535);
nand U11066 (N_11066,N_10824,N_10909);
or U11067 (N_11067,N_10706,N_10568);
xor U11068 (N_11068,N_10882,N_10782);
nor U11069 (N_11069,N_10804,N_10505);
nor U11070 (N_11070,N_10601,N_10881);
nand U11071 (N_11071,N_10715,N_10951);
or U11072 (N_11072,N_10991,N_10666);
nor U11073 (N_11073,N_10832,N_10691);
xnor U11074 (N_11074,N_10865,N_10852);
nor U11075 (N_11075,N_10830,N_10974);
and U11076 (N_11076,N_10924,N_10573);
xnor U11077 (N_11077,N_10744,N_10617);
nor U11078 (N_11078,N_10809,N_10928);
nor U11079 (N_11079,N_10556,N_10844);
nand U11080 (N_11080,N_10714,N_10687);
xor U11081 (N_11081,N_10866,N_10628);
and U11082 (N_11082,N_10903,N_10653);
or U11083 (N_11083,N_10604,N_10754);
nand U11084 (N_11084,N_10719,N_10877);
xor U11085 (N_11085,N_10746,N_10796);
nor U11086 (N_11086,N_10810,N_10858);
xnor U11087 (N_11087,N_10774,N_10520);
xor U11088 (N_11088,N_10587,N_10552);
xnor U11089 (N_11089,N_10849,N_10840);
nand U11090 (N_11090,N_10538,N_10627);
xor U11091 (N_11091,N_10555,N_10985);
or U11092 (N_11092,N_10867,N_10958);
nor U11093 (N_11093,N_10862,N_10519);
and U11094 (N_11094,N_10914,N_10721);
nand U11095 (N_11095,N_10775,N_10837);
or U11096 (N_11096,N_10994,N_10697);
nor U11097 (N_11097,N_10549,N_10708);
or U11098 (N_11098,N_10805,N_10959);
xor U11099 (N_11099,N_10762,N_10864);
or U11100 (N_11100,N_10883,N_10948);
nand U11101 (N_11101,N_10544,N_10845);
or U11102 (N_11102,N_10800,N_10524);
or U11103 (N_11103,N_10902,N_10701);
nand U11104 (N_11104,N_10968,N_10797);
nand U11105 (N_11105,N_10749,N_10815);
and U11106 (N_11106,N_10979,N_10600);
xor U11107 (N_11107,N_10536,N_10590);
nor U11108 (N_11108,N_10976,N_10553);
nor U11109 (N_11109,N_10869,N_10916);
xnor U11110 (N_11110,N_10884,N_10887);
nand U11111 (N_11111,N_10910,N_10850);
or U11112 (N_11112,N_10854,N_10503);
xor U11113 (N_11113,N_10682,N_10533);
or U11114 (N_11114,N_10838,N_10890);
nand U11115 (N_11115,N_10582,N_10955);
nor U11116 (N_11116,N_10760,N_10650);
xor U11117 (N_11117,N_10758,N_10793);
xor U11118 (N_11118,N_10624,N_10692);
nand U11119 (N_11119,N_10784,N_10722);
nand U11120 (N_11120,N_10818,N_10870);
nand U11121 (N_11121,N_10972,N_10702);
xor U11122 (N_11122,N_10602,N_10935);
nor U11123 (N_11123,N_10922,N_10785);
and U11124 (N_11124,N_10729,N_10780);
and U11125 (N_11125,N_10980,N_10672);
nor U11126 (N_11126,N_10759,N_10580);
xor U11127 (N_11127,N_10969,N_10569);
or U11128 (N_11128,N_10608,N_10900);
or U11129 (N_11129,N_10512,N_10745);
nand U11130 (N_11130,N_10735,N_10925);
nand U11131 (N_11131,N_10988,N_10637);
or U11132 (N_11132,N_10716,N_10543);
or U11133 (N_11133,N_10967,N_10983);
nor U11134 (N_11134,N_10638,N_10799);
nand U11135 (N_11135,N_10943,N_10839);
or U11136 (N_11136,N_10788,N_10908);
or U11137 (N_11137,N_10843,N_10879);
nor U11138 (N_11138,N_10753,N_10595);
xor U11139 (N_11139,N_10738,N_10631);
xnor U11140 (N_11140,N_10851,N_10901);
nand U11141 (N_11141,N_10531,N_10779);
nor U11142 (N_11142,N_10790,N_10649);
nor U11143 (N_11143,N_10787,N_10855);
or U11144 (N_11144,N_10829,N_10904);
and U11145 (N_11145,N_10675,N_10645);
nor U11146 (N_11146,N_10950,N_10828);
nand U11147 (N_11147,N_10940,N_10656);
xor U11148 (N_11148,N_10584,N_10550);
xnor U11149 (N_11149,N_10660,N_10609);
nand U11150 (N_11150,N_10530,N_10806);
and U11151 (N_11151,N_10560,N_10684);
nand U11152 (N_11152,N_10765,N_10963);
nor U11153 (N_11153,N_10892,N_10654);
and U11154 (N_11154,N_10794,N_10918);
nor U11155 (N_11155,N_10673,N_10564);
and U11156 (N_11156,N_10515,N_10688);
and U11157 (N_11157,N_10558,N_10554);
nor U11158 (N_11158,N_10623,N_10588);
xnor U11159 (N_11159,N_10990,N_10736);
nor U11160 (N_11160,N_10501,N_10597);
nor U11161 (N_11161,N_10966,N_10594);
nor U11162 (N_11162,N_10747,N_10571);
nand U11163 (N_11163,N_10891,N_10978);
and U11164 (N_11164,N_10548,N_10731);
xor U11165 (N_11165,N_10822,N_10644);
and U11166 (N_11166,N_10984,N_10529);
or U11167 (N_11167,N_10802,N_10846);
nor U11168 (N_11168,N_10647,N_10895);
or U11169 (N_11169,N_10872,N_10508);
xor U11170 (N_11170,N_10939,N_10757);
nor U11171 (N_11171,N_10664,N_10577);
or U11172 (N_11172,N_10504,N_10574);
or U11173 (N_11173,N_10670,N_10917);
xnor U11174 (N_11174,N_10603,N_10897);
nor U11175 (N_11175,N_10658,N_10827);
nand U11176 (N_11176,N_10527,N_10572);
nand U11177 (N_11177,N_10661,N_10781);
and U11178 (N_11178,N_10857,N_10965);
nand U11179 (N_11179,N_10921,N_10905);
xor U11180 (N_11180,N_10693,N_10842);
xor U11181 (N_11181,N_10931,N_10586);
nor U11182 (N_11182,N_10646,N_10710);
or U11183 (N_11183,N_10876,N_10570);
xor U11184 (N_11184,N_10836,N_10500);
and U11185 (N_11185,N_10926,N_10944);
or U11186 (N_11186,N_10880,N_10659);
nor U11187 (N_11187,N_10748,N_10562);
or U11188 (N_11188,N_10899,N_10709);
xor U11189 (N_11189,N_10596,N_10927);
xor U11190 (N_11190,N_10547,N_10546);
xnor U11191 (N_11191,N_10923,N_10634);
nand U11192 (N_11192,N_10750,N_10559);
nand U11193 (N_11193,N_10973,N_10534);
nand U11194 (N_11194,N_10703,N_10874);
nor U11195 (N_11195,N_10681,N_10894);
or U11196 (N_11196,N_10513,N_10756);
xnor U11197 (N_11197,N_10819,N_10737);
and U11198 (N_11198,N_10718,N_10607);
and U11199 (N_11199,N_10630,N_10847);
xor U11200 (N_11200,N_10826,N_10585);
nand U11201 (N_11201,N_10539,N_10725);
nand U11202 (N_11202,N_10919,N_10517);
nor U11203 (N_11203,N_10592,N_10542);
nor U11204 (N_11204,N_10801,N_10942);
or U11205 (N_11205,N_10772,N_10764);
nor U11206 (N_11206,N_10674,N_10639);
and U11207 (N_11207,N_10615,N_10616);
nand U11208 (N_11208,N_10522,N_10606);
nor U11209 (N_11209,N_10743,N_10532);
and U11210 (N_11210,N_10997,N_10551);
nand U11211 (N_11211,N_10937,N_10733);
or U11212 (N_11212,N_10893,N_10663);
or U11213 (N_11213,N_10589,N_10640);
nor U11214 (N_11214,N_10636,N_10778);
nor U11215 (N_11215,N_10998,N_10540);
nand U11216 (N_11216,N_10662,N_10696);
xor U11217 (N_11217,N_10578,N_10633);
xnor U11218 (N_11218,N_10545,N_10514);
or U11219 (N_11219,N_10506,N_10996);
and U11220 (N_11220,N_10612,N_10808);
xor U11221 (N_11221,N_10911,N_10705);
nor U11222 (N_11222,N_10912,N_10699);
nand U11223 (N_11223,N_10698,N_10798);
xnor U11224 (N_11224,N_10896,N_10930);
xnor U11225 (N_11225,N_10975,N_10977);
xor U11226 (N_11226,N_10575,N_10898);
xor U11227 (N_11227,N_10769,N_10643);
nand U11228 (N_11228,N_10868,N_10807);
xor U11229 (N_11229,N_10668,N_10981);
or U11230 (N_11230,N_10648,N_10954);
or U11231 (N_11231,N_10995,N_10665);
xnor U11232 (N_11232,N_10949,N_10755);
nand U11233 (N_11233,N_10690,N_10711);
nor U11234 (N_11234,N_10814,N_10694);
nand U11235 (N_11235,N_10689,N_10920);
or U11236 (N_11236,N_10962,N_10783);
and U11237 (N_11237,N_10795,N_10734);
nand U11238 (N_11238,N_10502,N_10619);
and U11239 (N_11239,N_10528,N_10565);
nand U11240 (N_11240,N_10971,N_10767);
nor U11241 (N_11241,N_10947,N_10871);
or U11242 (N_11242,N_10704,N_10982);
and U11243 (N_11243,N_10861,N_10825);
nor U11244 (N_11244,N_10510,N_10776);
xnor U11245 (N_11245,N_10523,N_10960);
nor U11246 (N_11246,N_10786,N_10987);
nand U11247 (N_11247,N_10576,N_10831);
nor U11248 (N_11248,N_10605,N_10707);
nand U11249 (N_11249,N_10713,N_10873);
nand U11250 (N_11250,N_10727,N_10996);
or U11251 (N_11251,N_10551,N_10879);
or U11252 (N_11252,N_10664,N_10970);
nand U11253 (N_11253,N_10796,N_10975);
or U11254 (N_11254,N_10559,N_10599);
or U11255 (N_11255,N_10746,N_10843);
or U11256 (N_11256,N_10521,N_10736);
nor U11257 (N_11257,N_10852,N_10519);
nand U11258 (N_11258,N_10578,N_10561);
nor U11259 (N_11259,N_10968,N_10553);
xnor U11260 (N_11260,N_10567,N_10578);
or U11261 (N_11261,N_10864,N_10691);
xor U11262 (N_11262,N_10840,N_10853);
xnor U11263 (N_11263,N_10728,N_10786);
or U11264 (N_11264,N_10525,N_10895);
nand U11265 (N_11265,N_10504,N_10866);
or U11266 (N_11266,N_10691,N_10942);
nand U11267 (N_11267,N_10853,N_10878);
nor U11268 (N_11268,N_10943,N_10824);
nor U11269 (N_11269,N_10767,N_10867);
xor U11270 (N_11270,N_10645,N_10862);
or U11271 (N_11271,N_10687,N_10668);
nor U11272 (N_11272,N_10654,N_10544);
nor U11273 (N_11273,N_10679,N_10509);
xnor U11274 (N_11274,N_10694,N_10791);
nand U11275 (N_11275,N_10567,N_10958);
nand U11276 (N_11276,N_10588,N_10919);
nor U11277 (N_11277,N_10748,N_10812);
nand U11278 (N_11278,N_10700,N_10503);
or U11279 (N_11279,N_10585,N_10755);
nand U11280 (N_11280,N_10542,N_10745);
nand U11281 (N_11281,N_10605,N_10817);
xor U11282 (N_11282,N_10687,N_10629);
or U11283 (N_11283,N_10632,N_10976);
xnor U11284 (N_11284,N_10805,N_10602);
nand U11285 (N_11285,N_10578,N_10846);
nor U11286 (N_11286,N_10659,N_10815);
nor U11287 (N_11287,N_10851,N_10942);
nand U11288 (N_11288,N_10514,N_10965);
nor U11289 (N_11289,N_10527,N_10736);
and U11290 (N_11290,N_10537,N_10574);
and U11291 (N_11291,N_10752,N_10982);
xnor U11292 (N_11292,N_10850,N_10894);
nand U11293 (N_11293,N_10911,N_10843);
nor U11294 (N_11294,N_10842,N_10665);
nor U11295 (N_11295,N_10765,N_10545);
nor U11296 (N_11296,N_10602,N_10897);
or U11297 (N_11297,N_10647,N_10502);
or U11298 (N_11298,N_10737,N_10860);
and U11299 (N_11299,N_10519,N_10812);
and U11300 (N_11300,N_10979,N_10989);
xor U11301 (N_11301,N_10641,N_10905);
xnor U11302 (N_11302,N_10818,N_10824);
or U11303 (N_11303,N_10776,N_10813);
nor U11304 (N_11304,N_10597,N_10650);
nand U11305 (N_11305,N_10600,N_10574);
nor U11306 (N_11306,N_10802,N_10906);
and U11307 (N_11307,N_10844,N_10623);
or U11308 (N_11308,N_10863,N_10961);
nor U11309 (N_11309,N_10964,N_10573);
nor U11310 (N_11310,N_10885,N_10737);
nand U11311 (N_11311,N_10589,N_10901);
xor U11312 (N_11312,N_10843,N_10898);
nand U11313 (N_11313,N_10776,N_10522);
and U11314 (N_11314,N_10665,N_10529);
xnor U11315 (N_11315,N_10735,N_10945);
nand U11316 (N_11316,N_10938,N_10832);
and U11317 (N_11317,N_10535,N_10909);
nand U11318 (N_11318,N_10687,N_10765);
xnor U11319 (N_11319,N_10737,N_10911);
xnor U11320 (N_11320,N_10849,N_10691);
nor U11321 (N_11321,N_10922,N_10604);
nor U11322 (N_11322,N_10796,N_10897);
and U11323 (N_11323,N_10776,N_10805);
and U11324 (N_11324,N_10612,N_10778);
or U11325 (N_11325,N_10558,N_10833);
or U11326 (N_11326,N_10923,N_10700);
and U11327 (N_11327,N_10793,N_10558);
and U11328 (N_11328,N_10792,N_10515);
or U11329 (N_11329,N_10513,N_10749);
nor U11330 (N_11330,N_10953,N_10973);
xnor U11331 (N_11331,N_10599,N_10617);
xnor U11332 (N_11332,N_10741,N_10565);
or U11333 (N_11333,N_10808,N_10831);
and U11334 (N_11334,N_10825,N_10853);
nor U11335 (N_11335,N_10666,N_10906);
nand U11336 (N_11336,N_10597,N_10941);
and U11337 (N_11337,N_10999,N_10830);
nand U11338 (N_11338,N_10656,N_10729);
or U11339 (N_11339,N_10899,N_10849);
and U11340 (N_11340,N_10678,N_10877);
nand U11341 (N_11341,N_10942,N_10760);
xnor U11342 (N_11342,N_10898,N_10788);
nor U11343 (N_11343,N_10594,N_10860);
or U11344 (N_11344,N_10902,N_10749);
or U11345 (N_11345,N_10501,N_10708);
nand U11346 (N_11346,N_10906,N_10992);
nor U11347 (N_11347,N_10567,N_10991);
and U11348 (N_11348,N_10783,N_10760);
or U11349 (N_11349,N_10525,N_10942);
and U11350 (N_11350,N_10716,N_10695);
nor U11351 (N_11351,N_10931,N_10918);
nand U11352 (N_11352,N_10956,N_10634);
and U11353 (N_11353,N_10649,N_10515);
or U11354 (N_11354,N_10700,N_10924);
or U11355 (N_11355,N_10540,N_10765);
nand U11356 (N_11356,N_10560,N_10612);
nor U11357 (N_11357,N_10720,N_10568);
nor U11358 (N_11358,N_10628,N_10699);
or U11359 (N_11359,N_10817,N_10944);
and U11360 (N_11360,N_10797,N_10810);
nand U11361 (N_11361,N_10593,N_10925);
and U11362 (N_11362,N_10502,N_10819);
nor U11363 (N_11363,N_10692,N_10598);
nand U11364 (N_11364,N_10998,N_10914);
xnor U11365 (N_11365,N_10913,N_10603);
nor U11366 (N_11366,N_10506,N_10514);
xnor U11367 (N_11367,N_10874,N_10999);
nand U11368 (N_11368,N_10645,N_10590);
nand U11369 (N_11369,N_10906,N_10955);
nand U11370 (N_11370,N_10563,N_10879);
or U11371 (N_11371,N_10715,N_10583);
xnor U11372 (N_11372,N_10630,N_10898);
nor U11373 (N_11373,N_10618,N_10609);
nand U11374 (N_11374,N_10562,N_10507);
xnor U11375 (N_11375,N_10794,N_10705);
nand U11376 (N_11376,N_10649,N_10929);
nand U11377 (N_11377,N_10771,N_10665);
nand U11378 (N_11378,N_10882,N_10772);
nand U11379 (N_11379,N_10935,N_10731);
xnor U11380 (N_11380,N_10687,N_10759);
nor U11381 (N_11381,N_10887,N_10637);
xor U11382 (N_11382,N_10614,N_10663);
or U11383 (N_11383,N_10970,N_10959);
nand U11384 (N_11384,N_10728,N_10967);
or U11385 (N_11385,N_10617,N_10830);
nand U11386 (N_11386,N_10866,N_10777);
and U11387 (N_11387,N_10687,N_10949);
or U11388 (N_11388,N_10847,N_10722);
nor U11389 (N_11389,N_10525,N_10566);
nand U11390 (N_11390,N_10967,N_10984);
xor U11391 (N_11391,N_10970,N_10872);
xor U11392 (N_11392,N_10604,N_10835);
nand U11393 (N_11393,N_10687,N_10931);
xnor U11394 (N_11394,N_10535,N_10776);
and U11395 (N_11395,N_10572,N_10797);
or U11396 (N_11396,N_10502,N_10750);
nor U11397 (N_11397,N_10740,N_10587);
nand U11398 (N_11398,N_10973,N_10826);
nor U11399 (N_11399,N_10665,N_10605);
xnor U11400 (N_11400,N_10685,N_10698);
nand U11401 (N_11401,N_10688,N_10593);
and U11402 (N_11402,N_10698,N_10650);
and U11403 (N_11403,N_10931,N_10741);
xor U11404 (N_11404,N_10617,N_10856);
xnor U11405 (N_11405,N_10673,N_10952);
nand U11406 (N_11406,N_10925,N_10622);
or U11407 (N_11407,N_10738,N_10805);
or U11408 (N_11408,N_10816,N_10743);
nor U11409 (N_11409,N_10500,N_10652);
or U11410 (N_11410,N_10513,N_10529);
xor U11411 (N_11411,N_10971,N_10639);
nand U11412 (N_11412,N_10915,N_10929);
and U11413 (N_11413,N_10758,N_10552);
nand U11414 (N_11414,N_10541,N_10636);
xor U11415 (N_11415,N_10908,N_10533);
nand U11416 (N_11416,N_10587,N_10545);
xor U11417 (N_11417,N_10813,N_10578);
and U11418 (N_11418,N_10609,N_10548);
xor U11419 (N_11419,N_10876,N_10927);
nor U11420 (N_11420,N_10709,N_10941);
and U11421 (N_11421,N_10718,N_10778);
nor U11422 (N_11422,N_10968,N_10990);
nor U11423 (N_11423,N_10977,N_10632);
xor U11424 (N_11424,N_10751,N_10663);
nand U11425 (N_11425,N_10648,N_10606);
xor U11426 (N_11426,N_10857,N_10709);
nor U11427 (N_11427,N_10692,N_10664);
and U11428 (N_11428,N_10799,N_10981);
nor U11429 (N_11429,N_10922,N_10577);
xnor U11430 (N_11430,N_10708,N_10770);
xor U11431 (N_11431,N_10817,N_10622);
nand U11432 (N_11432,N_10578,N_10611);
and U11433 (N_11433,N_10637,N_10502);
nand U11434 (N_11434,N_10862,N_10858);
and U11435 (N_11435,N_10662,N_10704);
or U11436 (N_11436,N_10672,N_10502);
nor U11437 (N_11437,N_10950,N_10813);
nand U11438 (N_11438,N_10886,N_10628);
and U11439 (N_11439,N_10511,N_10516);
nand U11440 (N_11440,N_10715,N_10909);
nor U11441 (N_11441,N_10986,N_10984);
and U11442 (N_11442,N_10561,N_10537);
nor U11443 (N_11443,N_10624,N_10885);
and U11444 (N_11444,N_10659,N_10687);
nor U11445 (N_11445,N_10906,N_10829);
nor U11446 (N_11446,N_10748,N_10784);
or U11447 (N_11447,N_10743,N_10710);
or U11448 (N_11448,N_10693,N_10983);
or U11449 (N_11449,N_10535,N_10669);
and U11450 (N_11450,N_10797,N_10683);
nor U11451 (N_11451,N_10713,N_10770);
nor U11452 (N_11452,N_10820,N_10898);
nand U11453 (N_11453,N_10597,N_10569);
or U11454 (N_11454,N_10909,N_10955);
nand U11455 (N_11455,N_10688,N_10931);
xor U11456 (N_11456,N_10974,N_10534);
xor U11457 (N_11457,N_10970,N_10910);
or U11458 (N_11458,N_10734,N_10988);
or U11459 (N_11459,N_10750,N_10894);
xnor U11460 (N_11460,N_10885,N_10900);
and U11461 (N_11461,N_10723,N_10507);
nor U11462 (N_11462,N_10849,N_10857);
or U11463 (N_11463,N_10986,N_10711);
nor U11464 (N_11464,N_10869,N_10709);
and U11465 (N_11465,N_10593,N_10561);
nand U11466 (N_11466,N_10591,N_10614);
nor U11467 (N_11467,N_10905,N_10882);
xnor U11468 (N_11468,N_10733,N_10758);
and U11469 (N_11469,N_10646,N_10791);
xor U11470 (N_11470,N_10573,N_10594);
or U11471 (N_11471,N_10793,N_10547);
xnor U11472 (N_11472,N_10947,N_10966);
nor U11473 (N_11473,N_10771,N_10737);
nor U11474 (N_11474,N_10895,N_10966);
xnor U11475 (N_11475,N_10886,N_10954);
xor U11476 (N_11476,N_10649,N_10708);
xor U11477 (N_11477,N_10587,N_10556);
nand U11478 (N_11478,N_10828,N_10966);
nand U11479 (N_11479,N_10993,N_10974);
nand U11480 (N_11480,N_10730,N_10633);
or U11481 (N_11481,N_10701,N_10749);
xor U11482 (N_11482,N_10859,N_10946);
xor U11483 (N_11483,N_10506,N_10999);
nor U11484 (N_11484,N_10911,N_10661);
nand U11485 (N_11485,N_10779,N_10624);
or U11486 (N_11486,N_10554,N_10592);
nor U11487 (N_11487,N_10799,N_10752);
or U11488 (N_11488,N_10628,N_10981);
nand U11489 (N_11489,N_10680,N_10730);
nand U11490 (N_11490,N_10647,N_10937);
nand U11491 (N_11491,N_10908,N_10894);
and U11492 (N_11492,N_10565,N_10516);
or U11493 (N_11493,N_10505,N_10925);
or U11494 (N_11494,N_10872,N_10648);
and U11495 (N_11495,N_10640,N_10534);
nand U11496 (N_11496,N_10710,N_10632);
nand U11497 (N_11497,N_10756,N_10561);
nor U11498 (N_11498,N_10659,N_10613);
nor U11499 (N_11499,N_10613,N_10739);
and U11500 (N_11500,N_11100,N_11327);
nand U11501 (N_11501,N_11298,N_11037);
xnor U11502 (N_11502,N_11186,N_11326);
xor U11503 (N_11503,N_11272,N_11023);
or U11504 (N_11504,N_11480,N_11178);
and U11505 (N_11505,N_11073,N_11123);
xor U11506 (N_11506,N_11174,N_11161);
and U11507 (N_11507,N_11315,N_11034);
or U11508 (N_11508,N_11493,N_11072);
nor U11509 (N_11509,N_11187,N_11429);
and U11510 (N_11510,N_11191,N_11454);
xnor U11511 (N_11511,N_11013,N_11038);
nor U11512 (N_11512,N_11200,N_11455);
nand U11513 (N_11513,N_11258,N_11403);
nor U11514 (N_11514,N_11088,N_11299);
nor U11515 (N_11515,N_11470,N_11251);
nand U11516 (N_11516,N_11410,N_11134);
nor U11517 (N_11517,N_11222,N_11496);
or U11518 (N_11518,N_11135,N_11069);
nor U11519 (N_11519,N_11061,N_11042);
nor U11520 (N_11520,N_11341,N_11428);
nor U11521 (N_11521,N_11059,N_11414);
nand U11522 (N_11522,N_11442,N_11147);
nand U11523 (N_11523,N_11494,N_11351);
and U11524 (N_11524,N_11364,N_11209);
nor U11525 (N_11525,N_11450,N_11342);
nor U11526 (N_11526,N_11130,N_11372);
nor U11527 (N_11527,N_11004,N_11089);
and U11528 (N_11528,N_11462,N_11374);
xnor U11529 (N_11529,N_11291,N_11482);
xor U11530 (N_11530,N_11030,N_11121);
or U11531 (N_11531,N_11395,N_11055);
nand U11532 (N_11532,N_11111,N_11153);
nand U11533 (N_11533,N_11360,N_11173);
nor U11534 (N_11534,N_11391,N_11213);
nand U11535 (N_11535,N_11460,N_11126);
nand U11536 (N_11536,N_11467,N_11129);
and U11537 (N_11537,N_11400,N_11456);
xor U11538 (N_11538,N_11443,N_11384);
and U11539 (N_11539,N_11057,N_11273);
nand U11540 (N_11540,N_11184,N_11216);
xnor U11541 (N_11541,N_11011,N_11353);
nand U11542 (N_11542,N_11307,N_11006);
and U11543 (N_11543,N_11346,N_11485);
and U11544 (N_11544,N_11194,N_11473);
nor U11545 (N_11545,N_11104,N_11045);
nor U11546 (N_11546,N_11425,N_11189);
and U11547 (N_11547,N_11260,N_11090);
or U11548 (N_11548,N_11483,N_11359);
xnor U11549 (N_11549,N_11431,N_11438);
or U11550 (N_11550,N_11257,N_11167);
xnor U11551 (N_11551,N_11052,N_11349);
and U11552 (N_11552,N_11312,N_11097);
xor U11553 (N_11553,N_11065,N_11110);
xor U11554 (N_11554,N_11196,N_11382);
nand U11555 (N_11555,N_11318,N_11303);
nand U11556 (N_11556,N_11305,N_11152);
and U11557 (N_11557,N_11197,N_11226);
nor U11558 (N_11558,N_11084,N_11387);
nand U11559 (N_11559,N_11475,N_11201);
nor U11560 (N_11560,N_11118,N_11219);
and U11561 (N_11561,N_11249,N_11019);
and U11562 (N_11562,N_11117,N_11220);
nand U11563 (N_11563,N_11381,N_11247);
or U11564 (N_11564,N_11175,N_11279);
xor U11565 (N_11565,N_11350,N_11422);
and U11566 (N_11566,N_11096,N_11000);
nand U11567 (N_11567,N_11266,N_11445);
and U11568 (N_11568,N_11099,N_11120);
and U11569 (N_11569,N_11434,N_11008);
nand U11570 (N_11570,N_11385,N_11457);
xor U11571 (N_11571,N_11239,N_11234);
xor U11572 (N_11572,N_11176,N_11396);
nor U11573 (N_11573,N_11012,N_11102);
nor U11574 (N_11574,N_11285,N_11363);
nand U11575 (N_11575,N_11250,N_11155);
and U11576 (N_11576,N_11078,N_11029);
and U11577 (N_11577,N_11166,N_11062);
xor U11578 (N_11578,N_11205,N_11053);
and U11579 (N_11579,N_11344,N_11369);
or U11580 (N_11580,N_11394,N_11339);
xnor U11581 (N_11581,N_11109,N_11486);
and U11582 (N_11582,N_11469,N_11106);
or U11583 (N_11583,N_11417,N_11143);
nor U11584 (N_11584,N_11499,N_11420);
xnor U11585 (N_11585,N_11287,N_11108);
xor U11586 (N_11586,N_11406,N_11018);
or U11587 (N_11587,N_11498,N_11066);
and U11588 (N_11588,N_11058,N_11028);
nand U11589 (N_11589,N_11484,N_11095);
nand U11590 (N_11590,N_11290,N_11325);
nand U11591 (N_11591,N_11481,N_11142);
nor U11592 (N_11592,N_11271,N_11337);
nand U11593 (N_11593,N_11440,N_11254);
or U11594 (N_11594,N_11221,N_11087);
and U11595 (N_11595,N_11208,N_11025);
xor U11596 (N_11596,N_11014,N_11301);
nand U11597 (N_11597,N_11217,N_11433);
nand U11598 (N_11598,N_11043,N_11446);
xnor U11599 (N_11599,N_11242,N_11017);
and U11600 (N_11600,N_11373,N_11465);
and U11601 (N_11601,N_11003,N_11094);
and U11602 (N_11602,N_11083,N_11060);
nor U11603 (N_11603,N_11032,N_11265);
nor U11604 (N_11604,N_11302,N_11453);
or U11605 (N_11605,N_11383,N_11471);
xor U11606 (N_11606,N_11340,N_11461);
nor U11607 (N_11607,N_11228,N_11050);
xnor U11608 (N_11608,N_11159,N_11252);
or U11609 (N_11609,N_11048,N_11160);
nor U11610 (N_11610,N_11421,N_11439);
or U11611 (N_11611,N_11296,N_11281);
and U11612 (N_11612,N_11039,N_11474);
nor U11613 (N_11613,N_11122,N_11136);
xnor U11614 (N_11614,N_11101,N_11026);
or U11615 (N_11615,N_11079,N_11235);
nand U11616 (N_11616,N_11098,N_11068);
nand U11617 (N_11617,N_11230,N_11033);
or U11618 (N_11618,N_11144,N_11211);
nor U11619 (N_11619,N_11386,N_11016);
nand U11620 (N_11620,N_11127,N_11168);
nand U11621 (N_11621,N_11323,N_11366);
xor U11622 (N_11622,N_11086,N_11437);
nand U11623 (N_11623,N_11031,N_11092);
xor U11624 (N_11624,N_11022,N_11172);
xor U11625 (N_11625,N_11085,N_11362);
and U11626 (N_11626,N_11367,N_11289);
nor U11627 (N_11627,N_11378,N_11427);
nand U11628 (N_11628,N_11401,N_11277);
nor U11629 (N_11629,N_11040,N_11371);
nand U11630 (N_11630,N_11046,N_11049);
nand U11631 (N_11631,N_11077,N_11492);
nor U11632 (N_11632,N_11407,N_11165);
xnor U11633 (N_11633,N_11182,N_11148);
nand U11634 (N_11634,N_11080,N_11444);
nor U11635 (N_11635,N_11105,N_11185);
nor U11636 (N_11636,N_11304,N_11063);
nand U11637 (N_11637,N_11036,N_11274);
nand U11638 (N_11638,N_11044,N_11286);
or U11639 (N_11639,N_11259,N_11365);
nand U11640 (N_11640,N_11157,N_11335);
xnor U11641 (N_11641,N_11308,N_11024);
nand U11642 (N_11642,N_11293,N_11392);
xnor U11643 (N_11643,N_11424,N_11261);
nand U11644 (N_11644,N_11449,N_11466);
and U11645 (N_11645,N_11270,N_11103);
and U11646 (N_11646,N_11495,N_11150);
nor U11647 (N_11647,N_11267,N_11477);
xor U11648 (N_11648,N_11310,N_11452);
xnor U11649 (N_11649,N_11206,N_11463);
nand U11650 (N_11650,N_11361,N_11133);
or U11651 (N_11651,N_11107,N_11294);
and U11652 (N_11652,N_11375,N_11070);
and U11653 (N_11653,N_11231,N_11114);
or U11654 (N_11654,N_11131,N_11227);
or U11655 (N_11655,N_11115,N_11202);
or U11656 (N_11656,N_11447,N_11021);
or U11657 (N_11657,N_11332,N_11156);
xnor U11658 (N_11658,N_11472,N_11334);
and U11659 (N_11659,N_11262,N_11284);
nand U11660 (N_11660,N_11190,N_11064);
or U11661 (N_11661,N_11275,N_11370);
or U11662 (N_11662,N_11204,N_11183);
xor U11663 (N_11663,N_11140,N_11354);
nor U11664 (N_11664,N_11311,N_11215);
or U11665 (N_11665,N_11380,N_11358);
nand U11666 (N_11666,N_11280,N_11181);
nor U11667 (N_11667,N_11238,N_11398);
nor U11668 (N_11668,N_11237,N_11321);
nor U11669 (N_11669,N_11336,N_11347);
and U11670 (N_11670,N_11419,N_11164);
nor U11671 (N_11671,N_11233,N_11243);
and U11672 (N_11672,N_11119,N_11459);
or U11673 (N_11673,N_11199,N_11405);
xnor U11674 (N_11674,N_11112,N_11268);
nand U11675 (N_11675,N_11348,N_11313);
xnor U11676 (N_11676,N_11377,N_11151);
or U11677 (N_11677,N_11316,N_11263);
or U11678 (N_11678,N_11116,N_11320);
nand U11679 (N_11679,N_11488,N_11487);
and U11680 (N_11680,N_11343,N_11352);
nor U11681 (N_11681,N_11020,N_11416);
nor U11682 (N_11682,N_11476,N_11379);
or U11683 (N_11683,N_11203,N_11253);
nand U11684 (N_11684,N_11244,N_11389);
nor U11685 (N_11685,N_11413,N_11137);
and U11686 (N_11686,N_11212,N_11232);
nor U11687 (N_11687,N_11225,N_11399);
and U11688 (N_11688,N_11338,N_11163);
nor U11689 (N_11689,N_11015,N_11468);
nor U11690 (N_11690,N_11322,N_11317);
or U11691 (N_11691,N_11328,N_11207);
nor U11692 (N_11692,N_11248,N_11179);
nand U11693 (N_11693,N_11397,N_11193);
nor U11694 (N_11694,N_11314,N_11376);
nand U11695 (N_11695,N_11412,N_11093);
nor U11696 (N_11696,N_11005,N_11458);
nor U11697 (N_11697,N_11241,N_11451);
xor U11698 (N_11698,N_11162,N_11229);
xor U11699 (N_11699,N_11051,N_11356);
nor U11700 (N_11700,N_11324,N_11132);
and U11701 (N_11701,N_11388,N_11245);
and U11702 (N_11702,N_11169,N_11441);
nor U11703 (N_11703,N_11368,N_11464);
xor U11704 (N_11704,N_11306,N_11214);
nor U11705 (N_11705,N_11223,N_11448);
and U11706 (N_11706,N_11218,N_11393);
nor U11707 (N_11707,N_11075,N_11423);
or U11708 (N_11708,N_11195,N_11479);
or U11709 (N_11709,N_11188,N_11141);
and U11710 (N_11710,N_11418,N_11282);
and U11711 (N_11711,N_11224,N_11124);
xor U11712 (N_11712,N_11139,N_11319);
xnor U11713 (N_11713,N_11297,N_11177);
nand U11714 (N_11714,N_11404,N_11435);
xnor U11715 (N_11715,N_11430,N_11180);
or U11716 (N_11716,N_11113,N_11255);
and U11717 (N_11717,N_11170,N_11478);
or U11718 (N_11718,N_11128,N_11278);
nor U11719 (N_11719,N_11149,N_11256);
nor U11720 (N_11720,N_11076,N_11357);
nand U11721 (N_11721,N_11411,N_11490);
or U11722 (N_11722,N_11091,N_11295);
and U11723 (N_11723,N_11035,N_11292);
nor U11724 (N_11724,N_11402,N_11192);
or U11725 (N_11725,N_11138,N_11283);
or U11726 (N_11726,N_11210,N_11047);
or U11727 (N_11727,N_11491,N_11288);
nor U11728 (N_11728,N_11027,N_11390);
nor U11729 (N_11729,N_11355,N_11007);
and U11730 (N_11730,N_11002,N_11125);
nor U11731 (N_11731,N_11236,N_11146);
nor U11732 (N_11732,N_11154,N_11300);
xnor U11733 (N_11733,N_11409,N_11331);
xnor U11734 (N_11734,N_11269,N_11067);
and U11735 (N_11735,N_11436,N_11309);
or U11736 (N_11736,N_11009,N_11082);
nor U11737 (N_11737,N_11246,N_11198);
xnor U11738 (N_11738,N_11001,N_11408);
nor U11739 (N_11739,N_11010,N_11240);
or U11740 (N_11740,N_11329,N_11330);
and U11741 (N_11741,N_11145,N_11171);
xnor U11742 (N_11742,N_11497,N_11158);
nor U11743 (N_11743,N_11426,N_11056);
nand U11744 (N_11744,N_11074,N_11264);
xnor U11745 (N_11745,N_11276,N_11415);
nor U11746 (N_11746,N_11489,N_11071);
or U11747 (N_11747,N_11041,N_11333);
xnor U11748 (N_11748,N_11081,N_11432);
nor U11749 (N_11749,N_11054,N_11345);
and U11750 (N_11750,N_11087,N_11440);
nor U11751 (N_11751,N_11128,N_11255);
and U11752 (N_11752,N_11467,N_11122);
xor U11753 (N_11753,N_11120,N_11224);
or U11754 (N_11754,N_11037,N_11195);
nor U11755 (N_11755,N_11385,N_11375);
nand U11756 (N_11756,N_11357,N_11336);
or U11757 (N_11757,N_11428,N_11386);
and U11758 (N_11758,N_11417,N_11482);
nand U11759 (N_11759,N_11022,N_11281);
nand U11760 (N_11760,N_11125,N_11280);
nor U11761 (N_11761,N_11454,N_11220);
xnor U11762 (N_11762,N_11208,N_11372);
or U11763 (N_11763,N_11319,N_11493);
nand U11764 (N_11764,N_11459,N_11160);
xor U11765 (N_11765,N_11082,N_11184);
and U11766 (N_11766,N_11490,N_11172);
or U11767 (N_11767,N_11264,N_11212);
and U11768 (N_11768,N_11352,N_11390);
xnor U11769 (N_11769,N_11069,N_11472);
or U11770 (N_11770,N_11205,N_11352);
and U11771 (N_11771,N_11233,N_11407);
xnor U11772 (N_11772,N_11493,N_11321);
xor U11773 (N_11773,N_11024,N_11051);
nor U11774 (N_11774,N_11404,N_11137);
xor U11775 (N_11775,N_11024,N_11036);
nand U11776 (N_11776,N_11165,N_11042);
nor U11777 (N_11777,N_11459,N_11162);
nand U11778 (N_11778,N_11036,N_11414);
xnor U11779 (N_11779,N_11103,N_11280);
xor U11780 (N_11780,N_11334,N_11018);
nand U11781 (N_11781,N_11223,N_11459);
nand U11782 (N_11782,N_11403,N_11439);
and U11783 (N_11783,N_11226,N_11466);
nor U11784 (N_11784,N_11251,N_11119);
xnor U11785 (N_11785,N_11420,N_11152);
and U11786 (N_11786,N_11083,N_11202);
or U11787 (N_11787,N_11140,N_11083);
or U11788 (N_11788,N_11351,N_11123);
nor U11789 (N_11789,N_11490,N_11008);
or U11790 (N_11790,N_11175,N_11318);
or U11791 (N_11791,N_11486,N_11498);
nand U11792 (N_11792,N_11308,N_11491);
xor U11793 (N_11793,N_11176,N_11261);
xor U11794 (N_11794,N_11298,N_11049);
xnor U11795 (N_11795,N_11168,N_11276);
or U11796 (N_11796,N_11385,N_11127);
xor U11797 (N_11797,N_11387,N_11293);
nor U11798 (N_11798,N_11324,N_11007);
or U11799 (N_11799,N_11245,N_11116);
and U11800 (N_11800,N_11344,N_11108);
nor U11801 (N_11801,N_11367,N_11228);
nand U11802 (N_11802,N_11295,N_11444);
nor U11803 (N_11803,N_11129,N_11174);
and U11804 (N_11804,N_11232,N_11006);
nor U11805 (N_11805,N_11083,N_11495);
xor U11806 (N_11806,N_11081,N_11377);
nor U11807 (N_11807,N_11286,N_11111);
nor U11808 (N_11808,N_11199,N_11330);
or U11809 (N_11809,N_11480,N_11471);
xnor U11810 (N_11810,N_11426,N_11408);
or U11811 (N_11811,N_11343,N_11406);
nand U11812 (N_11812,N_11468,N_11201);
nand U11813 (N_11813,N_11394,N_11157);
and U11814 (N_11814,N_11188,N_11473);
nand U11815 (N_11815,N_11445,N_11273);
or U11816 (N_11816,N_11437,N_11388);
xor U11817 (N_11817,N_11254,N_11449);
xnor U11818 (N_11818,N_11090,N_11353);
xnor U11819 (N_11819,N_11232,N_11311);
and U11820 (N_11820,N_11131,N_11026);
or U11821 (N_11821,N_11073,N_11192);
nor U11822 (N_11822,N_11466,N_11392);
or U11823 (N_11823,N_11102,N_11482);
xnor U11824 (N_11824,N_11491,N_11138);
xnor U11825 (N_11825,N_11103,N_11169);
nand U11826 (N_11826,N_11252,N_11375);
xor U11827 (N_11827,N_11192,N_11324);
nor U11828 (N_11828,N_11309,N_11129);
nand U11829 (N_11829,N_11110,N_11166);
nor U11830 (N_11830,N_11058,N_11422);
xnor U11831 (N_11831,N_11249,N_11391);
and U11832 (N_11832,N_11341,N_11187);
nor U11833 (N_11833,N_11336,N_11242);
xor U11834 (N_11834,N_11395,N_11243);
xnor U11835 (N_11835,N_11046,N_11172);
nand U11836 (N_11836,N_11130,N_11417);
or U11837 (N_11837,N_11064,N_11336);
or U11838 (N_11838,N_11476,N_11074);
and U11839 (N_11839,N_11315,N_11218);
nand U11840 (N_11840,N_11373,N_11164);
xnor U11841 (N_11841,N_11288,N_11225);
xor U11842 (N_11842,N_11376,N_11308);
and U11843 (N_11843,N_11300,N_11436);
xor U11844 (N_11844,N_11247,N_11143);
and U11845 (N_11845,N_11019,N_11476);
and U11846 (N_11846,N_11372,N_11222);
nand U11847 (N_11847,N_11366,N_11371);
and U11848 (N_11848,N_11243,N_11299);
nand U11849 (N_11849,N_11248,N_11121);
nand U11850 (N_11850,N_11021,N_11300);
or U11851 (N_11851,N_11172,N_11269);
and U11852 (N_11852,N_11428,N_11323);
and U11853 (N_11853,N_11189,N_11201);
xnor U11854 (N_11854,N_11396,N_11000);
nor U11855 (N_11855,N_11303,N_11454);
nor U11856 (N_11856,N_11381,N_11493);
and U11857 (N_11857,N_11433,N_11466);
and U11858 (N_11858,N_11027,N_11325);
or U11859 (N_11859,N_11160,N_11431);
and U11860 (N_11860,N_11157,N_11476);
nor U11861 (N_11861,N_11096,N_11220);
xnor U11862 (N_11862,N_11338,N_11000);
nor U11863 (N_11863,N_11496,N_11056);
nor U11864 (N_11864,N_11161,N_11394);
xor U11865 (N_11865,N_11245,N_11073);
or U11866 (N_11866,N_11466,N_11241);
or U11867 (N_11867,N_11369,N_11460);
xor U11868 (N_11868,N_11066,N_11470);
xnor U11869 (N_11869,N_11184,N_11113);
nor U11870 (N_11870,N_11086,N_11495);
nor U11871 (N_11871,N_11282,N_11351);
nand U11872 (N_11872,N_11013,N_11101);
nor U11873 (N_11873,N_11209,N_11354);
and U11874 (N_11874,N_11127,N_11158);
xnor U11875 (N_11875,N_11199,N_11417);
or U11876 (N_11876,N_11099,N_11127);
and U11877 (N_11877,N_11033,N_11156);
and U11878 (N_11878,N_11475,N_11345);
or U11879 (N_11879,N_11379,N_11435);
and U11880 (N_11880,N_11037,N_11104);
and U11881 (N_11881,N_11229,N_11282);
xnor U11882 (N_11882,N_11315,N_11401);
nand U11883 (N_11883,N_11374,N_11079);
nor U11884 (N_11884,N_11032,N_11217);
nand U11885 (N_11885,N_11261,N_11488);
xor U11886 (N_11886,N_11226,N_11209);
and U11887 (N_11887,N_11283,N_11056);
nor U11888 (N_11888,N_11194,N_11479);
or U11889 (N_11889,N_11358,N_11438);
or U11890 (N_11890,N_11316,N_11340);
and U11891 (N_11891,N_11351,N_11024);
nand U11892 (N_11892,N_11485,N_11408);
and U11893 (N_11893,N_11050,N_11022);
xnor U11894 (N_11894,N_11260,N_11170);
xor U11895 (N_11895,N_11224,N_11270);
and U11896 (N_11896,N_11386,N_11028);
nor U11897 (N_11897,N_11498,N_11264);
nand U11898 (N_11898,N_11161,N_11156);
or U11899 (N_11899,N_11394,N_11101);
xor U11900 (N_11900,N_11422,N_11382);
and U11901 (N_11901,N_11016,N_11148);
nor U11902 (N_11902,N_11330,N_11389);
and U11903 (N_11903,N_11233,N_11391);
xor U11904 (N_11904,N_11149,N_11215);
nor U11905 (N_11905,N_11307,N_11222);
nand U11906 (N_11906,N_11035,N_11200);
or U11907 (N_11907,N_11483,N_11267);
nand U11908 (N_11908,N_11127,N_11175);
or U11909 (N_11909,N_11017,N_11143);
nand U11910 (N_11910,N_11093,N_11221);
nor U11911 (N_11911,N_11323,N_11248);
or U11912 (N_11912,N_11129,N_11240);
or U11913 (N_11913,N_11347,N_11243);
nand U11914 (N_11914,N_11384,N_11194);
xnor U11915 (N_11915,N_11093,N_11084);
xor U11916 (N_11916,N_11188,N_11205);
nand U11917 (N_11917,N_11165,N_11174);
nor U11918 (N_11918,N_11024,N_11030);
or U11919 (N_11919,N_11394,N_11090);
nand U11920 (N_11920,N_11164,N_11472);
or U11921 (N_11921,N_11322,N_11206);
xor U11922 (N_11922,N_11334,N_11010);
and U11923 (N_11923,N_11384,N_11489);
nor U11924 (N_11924,N_11316,N_11264);
and U11925 (N_11925,N_11356,N_11288);
xnor U11926 (N_11926,N_11091,N_11133);
and U11927 (N_11927,N_11075,N_11381);
xnor U11928 (N_11928,N_11315,N_11006);
nand U11929 (N_11929,N_11267,N_11207);
or U11930 (N_11930,N_11148,N_11224);
or U11931 (N_11931,N_11064,N_11417);
nand U11932 (N_11932,N_11252,N_11115);
nand U11933 (N_11933,N_11119,N_11301);
nor U11934 (N_11934,N_11245,N_11211);
nand U11935 (N_11935,N_11103,N_11484);
or U11936 (N_11936,N_11053,N_11405);
nor U11937 (N_11937,N_11394,N_11184);
xnor U11938 (N_11938,N_11494,N_11270);
nor U11939 (N_11939,N_11470,N_11369);
and U11940 (N_11940,N_11478,N_11090);
and U11941 (N_11941,N_11469,N_11349);
and U11942 (N_11942,N_11228,N_11064);
nor U11943 (N_11943,N_11471,N_11496);
or U11944 (N_11944,N_11363,N_11104);
or U11945 (N_11945,N_11097,N_11063);
or U11946 (N_11946,N_11337,N_11037);
nor U11947 (N_11947,N_11008,N_11020);
and U11948 (N_11948,N_11328,N_11348);
or U11949 (N_11949,N_11106,N_11141);
and U11950 (N_11950,N_11399,N_11086);
or U11951 (N_11951,N_11265,N_11069);
and U11952 (N_11952,N_11013,N_11458);
nand U11953 (N_11953,N_11197,N_11440);
nor U11954 (N_11954,N_11015,N_11285);
xnor U11955 (N_11955,N_11260,N_11318);
and U11956 (N_11956,N_11083,N_11258);
xor U11957 (N_11957,N_11115,N_11286);
nand U11958 (N_11958,N_11402,N_11285);
nor U11959 (N_11959,N_11418,N_11123);
nor U11960 (N_11960,N_11394,N_11289);
nor U11961 (N_11961,N_11046,N_11103);
or U11962 (N_11962,N_11303,N_11296);
xnor U11963 (N_11963,N_11136,N_11495);
xnor U11964 (N_11964,N_11474,N_11025);
or U11965 (N_11965,N_11268,N_11395);
and U11966 (N_11966,N_11207,N_11403);
xor U11967 (N_11967,N_11264,N_11275);
nand U11968 (N_11968,N_11310,N_11444);
nor U11969 (N_11969,N_11447,N_11251);
nor U11970 (N_11970,N_11142,N_11036);
or U11971 (N_11971,N_11456,N_11442);
nor U11972 (N_11972,N_11370,N_11152);
nand U11973 (N_11973,N_11459,N_11024);
or U11974 (N_11974,N_11467,N_11110);
nand U11975 (N_11975,N_11471,N_11189);
nand U11976 (N_11976,N_11451,N_11252);
and U11977 (N_11977,N_11021,N_11368);
or U11978 (N_11978,N_11447,N_11422);
xor U11979 (N_11979,N_11106,N_11350);
xor U11980 (N_11980,N_11193,N_11211);
and U11981 (N_11981,N_11454,N_11424);
xnor U11982 (N_11982,N_11132,N_11069);
xnor U11983 (N_11983,N_11060,N_11329);
nor U11984 (N_11984,N_11473,N_11353);
nor U11985 (N_11985,N_11256,N_11205);
nand U11986 (N_11986,N_11165,N_11482);
or U11987 (N_11987,N_11244,N_11077);
nand U11988 (N_11988,N_11485,N_11370);
or U11989 (N_11989,N_11178,N_11207);
nor U11990 (N_11990,N_11146,N_11391);
or U11991 (N_11991,N_11224,N_11344);
xnor U11992 (N_11992,N_11203,N_11226);
or U11993 (N_11993,N_11432,N_11487);
nand U11994 (N_11994,N_11144,N_11434);
and U11995 (N_11995,N_11305,N_11318);
and U11996 (N_11996,N_11468,N_11321);
and U11997 (N_11997,N_11271,N_11276);
nor U11998 (N_11998,N_11323,N_11108);
or U11999 (N_11999,N_11118,N_11424);
nand U12000 (N_12000,N_11989,N_11860);
xnor U12001 (N_12001,N_11620,N_11711);
xnor U12002 (N_12002,N_11914,N_11726);
nand U12003 (N_12003,N_11763,N_11773);
nor U12004 (N_12004,N_11863,N_11800);
xor U12005 (N_12005,N_11881,N_11651);
or U12006 (N_12006,N_11782,N_11909);
nand U12007 (N_12007,N_11589,N_11984);
xnor U12008 (N_12008,N_11585,N_11619);
nor U12009 (N_12009,N_11802,N_11890);
nand U12010 (N_12010,N_11736,N_11981);
or U12011 (N_12011,N_11835,N_11727);
xor U12012 (N_12012,N_11621,N_11673);
nor U12013 (N_12013,N_11513,N_11794);
and U12014 (N_12014,N_11930,N_11861);
nor U12015 (N_12015,N_11707,N_11745);
nand U12016 (N_12016,N_11821,N_11533);
or U12017 (N_12017,N_11531,N_11778);
or U12018 (N_12018,N_11864,N_11983);
and U12019 (N_12019,N_11614,N_11574);
nand U12020 (N_12020,N_11561,N_11929);
or U12021 (N_12021,N_11940,N_11946);
nand U12022 (N_12022,N_11600,N_11719);
nand U12023 (N_12023,N_11739,N_11941);
and U12024 (N_12024,N_11575,N_11742);
nand U12025 (N_12025,N_11937,N_11862);
and U12026 (N_12026,N_11820,N_11622);
nor U12027 (N_12027,N_11826,N_11729);
nor U12028 (N_12028,N_11750,N_11968);
nor U12029 (N_12029,N_11834,N_11885);
or U12030 (N_12030,N_11550,N_11667);
xor U12031 (N_12031,N_11509,N_11807);
xnor U12032 (N_12032,N_11560,N_11936);
nand U12033 (N_12033,N_11738,N_11891);
nor U12034 (N_12034,N_11698,N_11646);
xor U12035 (N_12035,N_11846,N_11843);
nor U12036 (N_12036,N_11524,N_11920);
and U12037 (N_12037,N_11594,N_11757);
xnor U12038 (N_12038,N_11756,N_11808);
xor U12039 (N_12039,N_11894,N_11605);
nand U12040 (N_12040,N_11770,N_11876);
and U12041 (N_12041,N_11643,N_11565);
and U12042 (N_12042,N_11631,N_11693);
nand U12043 (N_12043,N_11922,N_11657);
and U12044 (N_12044,N_11805,N_11896);
or U12045 (N_12045,N_11710,N_11969);
nand U12046 (N_12046,N_11705,N_11677);
nand U12047 (N_12047,N_11943,N_11776);
nor U12048 (N_12048,N_11674,N_11767);
or U12049 (N_12049,N_11523,N_11957);
nor U12050 (N_12050,N_11558,N_11685);
or U12051 (N_12051,N_11919,N_11918);
xor U12052 (N_12052,N_11700,N_11966);
xor U12053 (N_12053,N_11534,N_11901);
or U12054 (N_12054,N_11851,N_11748);
nor U12055 (N_12055,N_11633,N_11869);
or U12056 (N_12056,N_11666,N_11987);
xnor U12057 (N_12057,N_11539,N_11988);
or U12058 (N_12058,N_11716,N_11598);
or U12059 (N_12059,N_11582,N_11768);
and U12060 (N_12060,N_11978,N_11601);
xor U12061 (N_12061,N_11553,N_11661);
nand U12062 (N_12062,N_11500,N_11559);
and U12063 (N_12063,N_11771,N_11516);
nand U12064 (N_12064,N_11734,N_11731);
and U12065 (N_12065,N_11687,N_11549);
xnor U12066 (N_12066,N_11766,N_11648);
nor U12067 (N_12067,N_11892,N_11917);
or U12068 (N_12068,N_11706,N_11905);
nor U12069 (N_12069,N_11916,N_11961);
nand U12070 (N_12070,N_11889,N_11508);
or U12071 (N_12071,N_11799,N_11662);
nor U12072 (N_12072,N_11725,N_11535);
or U12073 (N_12073,N_11686,N_11743);
nor U12074 (N_12074,N_11712,N_11762);
and U12075 (N_12075,N_11714,N_11609);
nand U12076 (N_12076,N_11564,N_11668);
nor U12077 (N_12077,N_11530,N_11840);
or U12078 (N_12078,N_11853,N_11828);
nor U12079 (N_12079,N_11596,N_11975);
nand U12080 (N_12080,N_11733,N_11570);
xor U12081 (N_12081,N_11624,N_11723);
nand U12082 (N_12082,N_11997,N_11584);
or U12083 (N_12083,N_11954,N_11977);
and U12084 (N_12084,N_11528,N_11907);
or U12085 (N_12085,N_11649,N_11640);
nor U12086 (N_12086,N_11688,N_11991);
nand U12087 (N_12087,N_11947,N_11897);
and U12088 (N_12088,N_11856,N_11709);
nor U12089 (N_12089,N_11903,N_11854);
nor U12090 (N_12090,N_11658,N_11525);
nor U12091 (N_12091,N_11985,N_11795);
nand U12092 (N_12092,N_11563,N_11730);
or U12093 (N_12093,N_11963,N_11680);
or U12094 (N_12094,N_11557,N_11728);
xnor U12095 (N_12095,N_11844,N_11838);
and U12096 (N_12096,N_11964,N_11702);
nor U12097 (N_12097,N_11599,N_11942);
and U12098 (N_12098,N_11664,N_11960);
and U12099 (N_12099,N_11696,N_11514);
and U12100 (N_12100,N_11502,N_11653);
nor U12101 (N_12101,N_11537,N_11852);
nor U12102 (N_12102,N_11694,N_11724);
nor U12103 (N_12103,N_11676,N_11758);
and U12104 (N_12104,N_11990,N_11986);
xnor U12105 (N_12105,N_11591,N_11813);
nand U12106 (N_12106,N_11720,N_11546);
or U12107 (N_12107,N_11971,N_11924);
and U12108 (N_12108,N_11635,N_11842);
and U12109 (N_12109,N_11634,N_11832);
nand U12110 (N_12110,N_11573,N_11612);
xnor U12111 (N_12111,N_11697,N_11928);
nand U12112 (N_12112,N_11519,N_11944);
nand U12113 (N_12113,N_11979,N_11779);
xnor U12114 (N_12114,N_11911,N_11865);
xor U12115 (N_12115,N_11543,N_11934);
nand U12116 (N_12116,N_11814,N_11717);
and U12117 (N_12117,N_11858,N_11749);
nand U12118 (N_12118,N_11790,N_11593);
or U12119 (N_12119,N_11850,N_11886);
and U12120 (N_12120,N_11684,N_11517);
xor U12121 (N_12121,N_11913,N_11735);
xor U12122 (N_12122,N_11998,N_11789);
or U12123 (N_12123,N_11970,N_11777);
nand U12124 (N_12124,N_11615,N_11660);
and U12125 (N_12125,N_11769,N_11610);
nand U12126 (N_12126,N_11837,N_11568);
or U12127 (N_12127,N_11713,N_11587);
and U12128 (N_12128,N_11857,N_11926);
nand U12129 (N_12129,N_11877,N_11921);
and U12130 (N_12130,N_11650,N_11812);
nor U12131 (N_12131,N_11787,N_11751);
xor U12132 (N_12132,N_11831,N_11786);
nand U12133 (N_12133,N_11670,N_11722);
nor U12134 (N_12134,N_11611,N_11547);
or U12135 (N_12135,N_11671,N_11900);
nor U12136 (N_12136,N_11718,N_11949);
and U12137 (N_12137,N_11950,N_11849);
and U12138 (N_12138,N_11999,N_11656);
and U12139 (N_12139,N_11761,N_11642);
and U12140 (N_12140,N_11695,N_11822);
nand U12141 (N_12141,N_11506,N_11578);
xor U12142 (N_12142,N_11566,N_11915);
and U12143 (N_12143,N_11772,N_11527);
nor U12144 (N_12144,N_11597,N_11616);
or U12145 (N_12145,N_11792,N_11791);
nor U12146 (N_12146,N_11625,N_11839);
nor U12147 (N_12147,N_11545,N_11816);
and U12148 (N_12148,N_11781,N_11654);
and U12149 (N_12149,N_11875,N_11953);
nand U12150 (N_12150,N_11632,N_11945);
nand U12151 (N_12151,N_11902,N_11793);
and U12152 (N_12152,N_11630,N_11753);
or U12153 (N_12153,N_11590,N_11692);
and U12154 (N_12154,N_11562,N_11636);
nor U12155 (N_12155,N_11827,N_11627);
xor U12156 (N_12156,N_11938,N_11811);
xnor U12157 (N_12157,N_11737,N_11689);
xnor U12158 (N_12158,N_11883,N_11880);
nor U12159 (N_12159,N_11867,N_11878);
nor U12160 (N_12160,N_11577,N_11606);
or U12161 (N_12161,N_11638,N_11955);
nor U12162 (N_12162,N_11899,N_11752);
xnor U12163 (N_12163,N_11721,N_11607);
and U12164 (N_12164,N_11933,N_11645);
nand U12165 (N_12165,N_11588,N_11829);
nor U12166 (N_12166,N_11796,N_11980);
or U12167 (N_12167,N_11542,N_11603);
nor U12168 (N_12168,N_11608,N_11912);
nand U12169 (N_12169,N_11927,N_11744);
and U12170 (N_12170,N_11996,N_11520);
nand U12171 (N_12171,N_11617,N_11595);
nand U12172 (N_12172,N_11974,N_11626);
nor U12173 (N_12173,N_11956,N_11823);
xor U12174 (N_12174,N_11583,N_11701);
nor U12175 (N_12175,N_11893,N_11592);
or U12176 (N_12176,N_11873,N_11629);
nor U12177 (N_12177,N_11879,N_11830);
xnor U12178 (N_12178,N_11683,N_11925);
and U12179 (N_12179,N_11521,N_11868);
and U12180 (N_12180,N_11848,N_11665);
xor U12181 (N_12181,N_11904,N_11503);
nor U12182 (N_12182,N_11958,N_11908);
or U12183 (N_12183,N_11678,N_11526);
nand U12184 (N_12184,N_11871,N_11623);
or U12185 (N_12185,N_11774,N_11544);
and U12186 (N_12186,N_11866,N_11884);
or U12187 (N_12187,N_11679,N_11572);
and U12188 (N_12188,N_11571,N_11505);
and U12189 (N_12189,N_11939,N_11872);
or U12190 (N_12190,N_11847,N_11501);
nor U12191 (N_12191,N_11579,N_11555);
nand U12192 (N_12192,N_11511,N_11510);
xor U12193 (N_12193,N_11699,N_11982);
or U12194 (N_12194,N_11952,N_11759);
and U12195 (N_12195,N_11888,N_11906);
nor U12196 (N_12196,N_11554,N_11551);
nand U12197 (N_12197,N_11825,N_11576);
xor U12198 (N_12198,N_11746,N_11740);
and U12199 (N_12199,N_11604,N_11931);
nor U12200 (N_12200,N_11715,N_11586);
xnor U12201 (N_12201,N_11552,N_11882);
or U12202 (N_12202,N_11910,N_11529);
or U12203 (N_12203,N_11798,N_11581);
nand U12204 (N_12204,N_11959,N_11644);
and U12205 (N_12205,N_11515,N_11817);
nor U12206 (N_12206,N_11784,N_11760);
xor U12207 (N_12207,N_11628,N_11874);
and U12208 (N_12208,N_11898,N_11732);
xor U12209 (N_12209,N_11538,N_11806);
nor U12210 (N_12210,N_11613,N_11652);
or U12211 (N_12211,N_11659,N_11704);
nor U12212 (N_12212,N_11703,N_11993);
xnor U12213 (N_12213,N_11672,N_11754);
xnor U12214 (N_12214,N_11948,N_11540);
nor U12215 (N_12215,N_11818,N_11895);
xnor U12216 (N_12216,N_11747,N_11994);
nor U12217 (N_12217,N_11788,N_11755);
and U12218 (N_12218,N_11841,N_11691);
xnor U12219 (N_12219,N_11962,N_11618);
nor U12220 (N_12220,N_11532,N_11965);
nand U12221 (N_12221,N_11815,N_11972);
nor U12222 (N_12222,N_11923,N_11803);
and U12223 (N_12223,N_11932,N_11836);
xnor U12224 (N_12224,N_11580,N_11859);
or U12225 (N_12225,N_11541,N_11602);
or U12226 (N_12226,N_11569,N_11976);
nand U12227 (N_12227,N_11522,N_11507);
xnor U12228 (N_12228,N_11512,N_11870);
nand U12229 (N_12229,N_11785,N_11775);
xor U12230 (N_12230,N_11663,N_11567);
xor U12231 (N_12231,N_11855,N_11973);
nand U12232 (N_12232,N_11675,N_11556);
xnor U12233 (N_12233,N_11819,N_11809);
nand U12234 (N_12234,N_11887,N_11797);
and U12235 (N_12235,N_11833,N_11783);
xnor U12236 (N_12236,N_11639,N_11504);
nor U12237 (N_12237,N_11804,N_11669);
or U12238 (N_12238,N_11708,N_11741);
xnor U12239 (N_12239,N_11951,N_11995);
or U12240 (N_12240,N_11655,N_11810);
nor U12241 (N_12241,N_11824,N_11967);
and U12242 (N_12242,N_11682,N_11641);
nand U12243 (N_12243,N_11536,N_11780);
and U12244 (N_12244,N_11845,N_11801);
nor U12245 (N_12245,N_11548,N_11637);
xor U12246 (N_12246,N_11647,N_11681);
and U12247 (N_12247,N_11935,N_11690);
and U12248 (N_12248,N_11518,N_11764);
nand U12249 (N_12249,N_11992,N_11765);
nand U12250 (N_12250,N_11667,N_11929);
nand U12251 (N_12251,N_11839,N_11744);
nand U12252 (N_12252,N_11838,N_11706);
or U12253 (N_12253,N_11979,N_11792);
or U12254 (N_12254,N_11868,N_11790);
nor U12255 (N_12255,N_11801,N_11799);
nand U12256 (N_12256,N_11613,N_11804);
and U12257 (N_12257,N_11611,N_11865);
or U12258 (N_12258,N_11887,N_11555);
and U12259 (N_12259,N_11998,N_11723);
or U12260 (N_12260,N_11712,N_11788);
nor U12261 (N_12261,N_11816,N_11731);
nand U12262 (N_12262,N_11682,N_11739);
xnor U12263 (N_12263,N_11814,N_11596);
xnor U12264 (N_12264,N_11639,N_11796);
and U12265 (N_12265,N_11973,N_11653);
xor U12266 (N_12266,N_11805,N_11930);
nor U12267 (N_12267,N_11745,N_11886);
xnor U12268 (N_12268,N_11711,N_11633);
and U12269 (N_12269,N_11922,N_11958);
xnor U12270 (N_12270,N_11518,N_11674);
nor U12271 (N_12271,N_11844,N_11796);
nand U12272 (N_12272,N_11654,N_11885);
or U12273 (N_12273,N_11730,N_11523);
and U12274 (N_12274,N_11627,N_11721);
nor U12275 (N_12275,N_11915,N_11582);
and U12276 (N_12276,N_11957,N_11735);
and U12277 (N_12277,N_11838,N_11590);
nand U12278 (N_12278,N_11688,N_11968);
nor U12279 (N_12279,N_11988,N_11925);
or U12280 (N_12280,N_11738,N_11776);
and U12281 (N_12281,N_11712,N_11533);
or U12282 (N_12282,N_11742,N_11648);
xnor U12283 (N_12283,N_11920,N_11742);
nand U12284 (N_12284,N_11671,N_11521);
nor U12285 (N_12285,N_11695,N_11780);
or U12286 (N_12286,N_11968,N_11878);
and U12287 (N_12287,N_11956,N_11913);
xnor U12288 (N_12288,N_11670,N_11781);
nand U12289 (N_12289,N_11923,N_11842);
xnor U12290 (N_12290,N_11908,N_11737);
nor U12291 (N_12291,N_11911,N_11658);
nor U12292 (N_12292,N_11734,N_11501);
xnor U12293 (N_12293,N_11836,N_11951);
or U12294 (N_12294,N_11638,N_11848);
nor U12295 (N_12295,N_11961,N_11571);
nand U12296 (N_12296,N_11885,N_11665);
or U12297 (N_12297,N_11904,N_11579);
and U12298 (N_12298,N_11954,N_11590);
and U12299 (N_12299,N_11896,N_11635);
nand U12300 (N_12300,N_11515,N_11932);
nand U12301 (N_12301,N_11650,N_11760);
xnor U12302 (N_12302,N_11590,N_11979);
or U12303 (N_12303,N_11985,N_11922);
nand U12304 (N_12304,N_11967,N_11764);
xor U12305 (N_12305,N_11770,N_11525);
nand U12306 (N_12306,N_11908,N_11876);
and U12307 (N_12307,N_11997,N_11626);
xor U12308 (N_12308,N_11650,N_11520);
nor U12309 (N_12309,N_11931,N_11986);
xor U12310 (N_12310,N_11732,N_11866);
and U12311 (N_12311,N_11623,N_11939);
and U12312 (N_12312,N_11530,N_11656);
nand U12313 (N_12313,N_11842,N_11718);
or U12314 (N_12314,N_11792,N_11952);
nor U12315 (N_12315,N_11651,N_11747);
and U12316 (N_12316,N_11714,N_11728);
xor U12317 (N_12317,N_11612,N_11725);
nor U12318 (N_12318,N_11580,N_11667);
xnor U12319 (N_12319,N_11741,N_11879);
and U12320 (N_12320,N_11755,N_11664);
xor U12321 (N_12321,N_11509,N_11973);
or U12322 (N_12322,N_11739,N_11517);
xor U12323 (N_12323,N_11844,N_11732);
xor U12324 (N_12324,N_11797,N_11631);
or U12325 (N_12325,N_11793,N_11907);
nor U12326 (N_12326,N_11536,N_11579);
or U12327 (N_12327,N_11682,N_11882);
nand U12328 (N_12328,N_11755,N_11581);
and U12329 (N_12329,N_11774,N_11504);
and U12330 (N_12330,N_11739,N_11735);
and U12331 (N_12331,N_11756,N_11574);
xnor U12332 (N_12332,N_11679,N_11881);
xor U12333 (N_12333,N_11642,N_11771);
nand U12334 (N_12334,N_11862,N_11836);
nor U12335 (N_12335,N_11970,N_11807);
or U12336 (N_12336,N_11536,N_11524);
xor U12337 (N_12337,N_11791,N_11739);
nand U12338 (N_12338,N_11868,N_11640);
nand U12339 (N_12339,N_11550,N_11801);
or U12340 (N_12340,N_11607,N_11743);
or U12341 (N_12341,N_11699,N_11690);
or U12342 (N_12342,N_11769,N_11685);
xnor U12343 (N_12343,N_11566,N_11980);
nand U12344 (N_12344,N_11731,N_11526);
nor U12345 (N_12345,N_11824,N_11809);
xor U12346 (N_12346,N_11862,N_11869);
or U12347 (N_12347,N_11552,N_11902);
nor U12348 (N_12348,N_11623,N_11776);
nand U12349 (N_12349,N_11973,N_11684);
or U12350 (N_12350,N_11864,N_11715);
and U12351 (N_12351,N_11855,N_11844);
or U12352 (N_12352,N_11815,N_11581);
xnor U12353 (N_12353,N_11902,N_11576);
nor U12354 (N_12354,N_11647,N_11650);
and U12355 (N_12355,N_11702,N_11897);
or U12356 (N_12356,N_11818,N_11874);
nor U12357 (N_12357,N_11559,N_11711);
xnor U12358 (N_12358,N_11799,N_11640);
nand U12359 (N_12359,N_11898,N_11503);
and U12360 (N_12360,N_11539,N_11618);
and U12361 (N_12361,N_11534,N_11800);
nand U12362 (N_12362,N_11646,N_11967);
or U12363 (N_12363,N_11989,N_11579);
or U12364 (N_12364,N_11875,N_11937);
xnor U12365 (N_12365,N_11713,N_11763);
xor U12366 (N_12366,N_11661,N_11887);
or U12367 (N_12367,N_11530,N_11581);
and U12368 (N_12368,N_11899,N_11565);
xor U12369 (N_12369,N_11723,N_11697);
nor U12370 (N_12370,N_11738,N_11558);
or U12371 (N_12371,N_11542,N_11776);
xnor U12372 (N_12372,N_11753,N_11813);
nor U12373 (N_12373,N_11568,N_11599);
xor U12374 (N_12374,N_11765,N_11604);
nor U12375 (N_12375,N_11893,N_11944);
nor U12376 (N_12376,N_11556,N_11704);
and U12377 (N_12377,N_11790,N_11715);
nand U12378 (N_12378,N_11751,N_11867);
or U12379 (N_12379,N_11524,N_11657);
nand U12380 (N_12380,N_11645,N_11717);
and U12381 (N_12381,N_11950,N_11834);
or U12382 (N_12382,N_11835,N_11710);
and U12383 (N_12383,N_11995,N_11846);
nor U12384 (N_12384,N_11732,N_11500);
or U12385 (N_12385,N_11947,N_11555);
nor U12386 (N_12386,N_11554,N_11892);
xor U12387 (N_12387,N_11829,N_11560);
nand U12388 (N_12388,N_11941,N_11729);
or U12389 (N_12389,N_11904,N_11943);
and U12390 (N_12390,N_11523,N_11623);
or U12391 (N_12391,N_11528,N_11504);
nand U12392 (N_12392,N_11537,N_11638);
xnor U12393 (N_12393,N_11693,N_11718);
or U12394 (N_12394,N_11506,N_11889);
and U12395 (N_12395,N_11887,N_11705);
and U12396 (N_12396,N_11807,N_11784);
or U12397 (N_12397,N_11823,N_11515);
and U12398 (N_12398,N_11692,N_11852);
nand U12399 (N_12399,N_11739,N_11704);
or U12400 (N_12400,N_11983,N_11894);
nand U12401 (N_12401,N_11562,N_11976);
xnor U12402 (N_12402,N_11692,N_11837);
and U12403 (N_12403,N_11547,N_11509);
xor U12404 (N_12404,N_11889,N_11964);
xor U12405 (N_12405,N_11860,N_11995);
nand U12406 (N_12406,N_11575,N_11978);
or U12407 (N_12407,N_11522,N_11985);
nor U12408 (N_12408,N_11754,N_11612);
xor U12409 (N_12409,N_11765,N_11735);
or U12410 (N_12410,N_11609,N_11840);
and U12411 (N_12411,N_11880,N_11948);
xnor U12412 (N_12412,N_11974,N_11899);
xor U12413 (N_12413,N_11683,N_11671);
and U12414 (N_12414,N_11717,N_11983);
nor U12415 (N_12415,N_11577,N_11634);
and U12416 (N_12416,N_11631,N_11993);
xnor U12417 (N_12417,N_11586,N_11610);
nor U12418 (N_12418,N_11931,N_11997);
nand U12419 (N_12419,N_11950,N_11915);
or U12420 (N_12420,N_11795,N_11846);
nor U12421 (N_12421,N_11825,N_11922);
or U12422 (N_12422,N_11581,N_11924);
nor U12423 (N_12423,N_11658,N_11514);
nor U12424 (N_12424,N_11565,N_11993);
xor U12425 (N_12425,N_11670,N_11944);
nor U12426 (N_12426,N_11673,N_11786);
nand U12427 (N_12427,N_11928,N_11507);
nand U12428 (N_12428,N_11731,N_11994);
or U12429 (N_12429,N_11514,N_11944);
nor U12430 (N_12430,N_11615,N_11897);
nand U12431 (N_12431,N_11879,N_11864);
and U12432 (N_12432,N_11882,N_11693);
nand U12433 (N_12433,N_11972,N_11951);
and U12434 (N_12434,N_11617,N_11821);
nor U12435 (N_12435,N_11606,N_11924);
and U12436 (N_12436,N_11757,N_11741);
and U12437 (N_12437,N_11794,N_11512);
nand U12438 (N_12438,N_11919,N_11668);
and U12439 (N_12439,N_11897,N_11801);
xor U12440 (N_12440,N_11700,N_11979);
and U12441 (N_12441,N_11534,N_11867);
nor U12442 (N_12442,N_11723,N_11555);
or U12443 (N_12443,N_11547,N_11816);
xnor U12444 (N_12444,N_11690,N_11829);
and U12445 (N_12445,N_11909,N_11525);
nor U12446 (N_12446,N_11607,N_11805);
or U12447 (N_12447,N_11877,N_11616);
or U12448 (N_12448,N_11622,N_11680);
or U12449 (N_12449,N_11741,N_11816);
nor U12450 (N_12450,N_11575,N_11991);
xnor U12451 (N_12451,N_11523,N_11630);
or U12452 (N_12452,N_11898,N_11782);
nand U12453 (N_12453,N_11890,N_11627);
nor U12454 (N_12454,N_11656,N_11675);
nor U12455 (N_12455,N_11876,N_11786);
xnor U12456 (N_12456,N_11567,N_11986);
xnor U12457 (N_12457,N_11652,N_11564);
nor U12458 (N_12458,N_11979,N_11546);
nor U12459 (N_12459,N_11640,N_11674);
and U12460 (N_12460,N_11529,N_11647);
nor U12461 (N_12461,N_11545,N_11795);
or U12462 (N_12462,N_11802,N_11858);
xor U12463 (N_12463,N_11837,N_11705);
or U12464 (N_12464,N_11693,N_11641);
and U12465 (N_12465,N_11525,N_11782);
nand U12466 (N_12466,N_11728,N_11976);
nand U12467 (N_12467,N_11511,N_11667);
xnor U12468 (N_12468,N_11683,N_11612);
nand U12469 (N_12469,N_11923,N_11925);
nand U12470 (N_12470,N_11986,N_11810);
nand U12471 (N_12471,N_11884,N_11612);
xor U12472 (N_12472,N_11686,N_11673);
nand U12473 (N_12473,N_11987,N_11870);
xor U12474 (N_12474,N_11738,N_11762);
nand U12475 (N_12475,N_11834,N_11675);
nor U12476 (N_12476,N_11534,N_11974);
nand U12477 (N_12477,N_11835,N_11804);
and U12478 (N_12478,N_11852,N_11523);
nand U12479 (N_12479,N_11537,N_11936);
nand U12480 (N_12480,N_11899,N_11538);
nand U12481 (N_12481,N_11661,N_11554);
and U12482 (N_12482,N_11770,N_11898);
and U12483 (N_12483,N_11664,N_11534);
xor U12484 (N_12484,N_11529,N_11636);
nor U12485 (N_12485,N_11593,N_11994);
xor U12486 (N_12486,N_11836,N_11777);
or U12487 (N_12487,N_11757,N_11937);
and U12488 (N_12488,N_11614,N_11570);
and U12489 (N_12489,N_11970,N_11530);
xnor U12490 (N_12490,N_11938,N_11813);
nand U12491 (N_12491,N_11652,N_11969);
xor U12492 (N_12492,N_11592,N_11542);
nand U12493 (N_12493,N_11881,N_11998);
and U12494 (N_12494,N_11713,N_11507);
and U12495 (N_12495,N_11627,N_11589);
xor U12496 (N_12496,N_11610,N_11619);
nor U12497 (N_12497,N_11667,N_11890);
nand U12498 (N_12498,N_11819,N_11628);
xnor U12499 (N_12499,N_11894,N_11765);
or U12500 (N_12500,N_12270,N_12493);
nor U12501 (N_12501,N_12437,N_12370);
or U12502 (N_12502,N_12241,N_12231);
xnor U12503 (N_12503,N_12349,N_12117);
nand U12504 (N_12504,N_12175,N_12113);
and U12505 (N_12505,N_12305,N_12386);
xnor U12506 (N_12506,N_12411,N_12445);
xnor U12507 (N_12507,N_12329,N_12194);
or U12508 (N_12508,N_12348,N_12212);
nor U12509 (N_12509,N_12120,N_12234);
nand U12510 (N_12510,N_12224,N_12243);
or U12511 (N_12511,N_12337,N_12235);
nor U12512 (N_12512,N_12354,N_12443);
nor U12513 (N_12513,N_12080,N_12280);
nor U12514 (N_12514,N_12090,N_12127);
xor U12515 (N_12515,N_12003,N_12303);
nand U12516 (N_12516,N_12133,N_12424);
or U12517 (N_12517,N_12099,N_12442);
nor U12518 (N_12518,N_12053,N_12483);
and U12519 (N_12519,N_12195,N_12159);
and U12520 (N_12520,N_12131,N_12473);
and U12521 (N_12521,N_12388,N_12332);
xnor U12522 (N_12522,N_12236,N_12446);
xor U12523 (N_12523,N_12309,N_12086);
and U12524 (N_12524,N_12485,N_12032);
or U12525 (N_12525,N_12230,N_12060);
nor U12526 (N_12526,N_12497,N_12326);
nor U12527 (N_12527,N_12094,N_12266);
nor U12528 (N_12528,N_12284,N_12366);
nand U12529 (N_12529,N_12110,N_12167);
xnor U12530 (N_12530,N_12142,N_12017);
and U12531 (N_12531,N_12097,N_12440);
and U12532 (N_12532,N_12342,N_12359);
nor U12533 (N_12533,N_12433,N_12256);
nor U12534 (N_12534,N_12286,N_12168);
nor U12535 (N_12535,N_12338,N_12277);
or U12536 (N_12536,N_12290,N_12129);
and U12537 (N_12537,N_12197,N_12271);
or U12538 (N_12538,N_12054,N_12148);
and U12539 (N_12539,N_12403,N_12237);
nand U12540 (N_12540,N_12317,N_12265);
nand U12541 (N_12541,N_12066,N_12061);
nor U12542 (N_12542,N_12334,N_12164);
nor U12543 (N_12543,N_12124,N_12415);
xor U12544 (N_12544,N_12019,N_12021);
and U12545 (N_12545,N_12052,N_12214);
nor U12546 (N_12546,N_12367,N_12145);
or U12547 (N_12547,N_12034,N_12268);
xor U12548 (N_12548,N_12383,N_12050);
nor U12549 (N_12549,N_12183,N_12478);
and U12550 (N_12550,N_12315,N_12176);
nor U12551 (N_12551,N_12161,N_12213);
nand U12552 (N_12552,N_12389,N_12081);
or U12553 (N_12553,N_12378,N_12249);
xor U12554 (N_12554,N_12227,N_12414);
and U12555 (N_12555,N_12360,N_12391);
and U12556 (N_12556,N_12393,N_12458);
xnor U12557 (N_12557,N_12084,N_12384);
nor U12558 (N_12558,N_12375,N_12122);
and U12559 (N_12559,N_12104,N_12217);
or U12560 (N_12560,N_12198,N_12158);
nand U12561 (N_12561,N_12327,N_12455);
nand U12562 (N_12562,N_12079,N_12258);
nor U12563 (N_12563,N_12312,N_12347);
xnor U12564 (N_12564,N_12273,N_12428);
or U12565 (N_12565,N_12007,N_12188);
nand U12566 (N_12566,N_12035,N_12068);
xor U12567 (N_12567,N_12141,N_12123);
and U12568 (N_12568,N_12373,N_12336);
or U12569 (N_12569,N_12390,N_12065);
and U12570 (N_12570,N_12335,N_12288);
xor U12571 (N_12571,N_12192,N_12490);
and U12572 (N_12572,N_12203,N_12207);
xnor U12573 (N_12573,N_12024,N_12229);
nand U12574 (N_12574,N_12029,N_12102);
or U12575 (N_12575,N_12208,N_12301);
xnor U12576 (N_12576,N_12018,N_12308);
nand U12577 (N_12577,N_12444,N_12289);
and U12578 (N_12578,N_12431,N_12240);
or U12579 (N_12579,N_12162,N_12394);
nor U12580 (N_12580,N_12355,N_12330);
nor U12581 (N_12581,N_12452,N_12044);
and U12582 (N_12582,N_12457,N_12484);
and U12583 (N_12583,N_12014,N_12477);
or U12584 (N_12584,N_12170,N_12196);
and U12585 (N_12585,N_12321,N_12278);
and U12586 (N_12586,N_12404,N_12260);
nand U12587 (N_12587,N_12298,N_12331);
and U12588 (N_12588,N_12441,N_12163);
and U12589 (N_12589,N_12041,N_12223);
and U12590 (N_12590,N_12460,N_12180);
and U12591 (N_12591,N_12151,N_12185);
nand U12592 (N_12592,N_12296,N_12328);
and U12593 (N_12593,N_12062,N_12089);
and U12594 (N_12594,N_12105,N_12263);
and U12595 (N_12595,N_12177,N_12209);
xor U12596 (N_12596,N_12250,N_12135);
xor U12597 (N_12597,N_12439,N_12339);
xnor U12598 (N_12598,N_12106,N_12480);
nand U12599 (N_12599,N_12323,N_12146);
xor U12600 (N_12600,N_12039,N_12137);
and U12601 (N_12601,N_12115,N_12472);
nor U12602 (N_12602,N_12109,N_12076);
nor U12603 (N_12603,N_12487,N_12307);
nor U12604 (N_12604,N_12495,N_12351);
and U12605 (N_12605,N_12365,N_12184);
xnor U12606 (N_12606,N_12417,N_12125);
and U12607 (N_12607,N_12160,N_12190);
nor U12608 (N_12608,N_12087,N_12130);
nand U12609 (N_12609,N_12095,N_12465);
nor U12610 (N_12610,N_12252,N_12325);
nor U12611 (N_12611,N_12239,N_12363);
or U12612 (N_12612,N_12179,N_12282);
nor U12613 (N_12613,N_12055,N_12222);
nor U12614 (N_12614,N_12456,N_12299);
xor U12615 (N_12615,N_12311,N_12369);
or U12616 (N_12616,N_12413,N_12264);
or U12617 (N_12617,N_12259,N_12011);
xor U12618 (N_12618,N_12418,N_12462);
or U12619 (N_12619,N_12476,N_12000);
and U12620 (N_12620,N_12381,N_12344);
nor U12621 (N_12621,N_12049,N_12242);
nor U12622 (N_12622,N_12324,N_12147);
or U12623 (N_12623,N_12279,N_12205);
nor U12624 (N_12624,N_12453,N_12416);
or U12625 (N_12625,N_12356,N_12255);
xor U12626 (N_12626,N_12199,N_12316);
xor U12627 (N_12627,N_12063,N_12475);
and U12628 (N_12628,N_12406,N_12215);
or U12629 (N_12629,N_12319,N_12101);
or U12630 (N_12630,N_12267,N_12353);
and U12631 (N_12631,N_12362,N_12025);
or U12632 (N_12632,N_12096,N_12173);
and U12633 (N_12633,N_12494,N_12488);
xnor U12634 (N_12634,N_12139,N_12376);
nor U12635 (N_12635,N_12272,N_12281);
nor U12636 (N_12636,N_12067,N_12352);
nor U12637 (N_12637,N_12009,N_12333);
xor U12638 (N_12638,N_12200,N_12165);
nand U12639 (N_12639,N_12379,N_12189);
or U12640 (N_12640,N_12112,N_12100);
nor U12641 (N_12641,N_12470,N_12037);
or U12642 (N_12642,N_12471,N_12346);
and U12643 (N_12643,N_12128,N_12374);
nand U12644 (N_12644,N_12191,N_12233);
xnor U12645 (N_12645,N_12064,N_12447);
nor U12646 (N_12646,N_12499,N_12006);
nor U12647 (N_12647,N_12297,N_12496);
xnor U12648 (N_12648,N_12253,N_12091);
nor U12649 (N_12649,N_12116,N_12345);
nand U12650 (N_12650,N_12341,N_12204);
and U12651 (N_12651,N_12078,N_12144);
and U12652 (N_12652,N_12201,N_12459);
or U12653 (N_12653,N_12225,N_12082);
xor U12654 (N_12654,N_12031,N_12482);
and U12655 (N_12655,N_12318,N_12069);
nor U12656 (N_12656,N_12038,N_12294);
or U12657 (N_12657,N_12045,N_12040);
nor U12658 (N_12658,N_12121,N_12461);
nor U12659 (N_12659,N_12057,N_12464);
and U12660 (N_12660,N_12292,N_12397);
and U12661 (N_12661,N_12005,N_12155);
nand U12662 (N_12662,N_12036,N_12254);
or U12663 (N_12663,N_12410,N_12219);
and U12664 (N_12664,N_12436,N_12398);
xor U12665 (N_12665,N_12412,N_12186);
or U12666 (N_12666,N_12275,N_12310);
nor U12667 (N_12667,N_12300,N_12467);
or U12668 (N_12668,N_12246,N_12020);
nand U12669 (N_12669,N_12430,N_12111);
xnor U12670 (N_12670,N_12427,N_12257);
and U12671 (N_12671,N_12153,N_12401);
and U12672 (N_12672,N_12276,N_12274);
and U12673 (N_12673,N_12372,N_12429);
nor U12674 (N_12674,N_12469,N_12202);
and U12675 (N_12675,N_12407,N_12293);
xor U12676 (N_12676,N_12498,N_12387);
or U12677 (N_12677,N_12134,N_12371);
xnor U12678 (N_12678,N_12451,N_12466);
or U12679 (N_12679,N_12103,N_12450);
nand U12680 (N_12680,N_12232,N_12088);
nor U12681 (N_12681,N_12075,N_12420);
xnor U12682 (N_12682,N_12262,N_12304);
nand U12683 (N_12683,N_12357,N_12491);
xor U12684 (N_12684,N_12419,N_12479);
or U12685 (N_12685,N_12350,N_12178);
xnor U12686 (N_12686,N_12313,N_12056);
nand U12687 (N_12687,N_12030,N_12216);
xor U12688 (N_12688,N_12166,N_12405);
nand U12689 (N_12689,N_12238,N_12211);
and U12690 (N_12690,N_12048,N_12320);
xor U12691 (N_12691,N_12098,N_12013);
nand U12692 (N_12692,N_12107,N_12042);
nor U12693 (N_12693,N_12193,N_12154);
and U12694 (N_12694,N_12187,N_12138);
nand U12695 (N_12695,N_12181,N_12156);
nand U12696 (N_12696,N_12409,N_12454);
or U12697 (N_12697,N_12395,N_12059);
and U12698 (N_12698,N_12364,N_12382);
nand U12699 (N_12699,N_12283,N_12400);
nand U12700 (N_12700,N_12302,N_12343);
xor U12701 (N_12701,N_12248,N_12314);
or U12702 (N_12702,N_12072,N_12152);
or U12703 (N_12703,N_12463,N_12285);
nor U12704 (N_12704,N_12399,N_12426);
nand U12705 (N_12705,N_12468,N_12244);
xnor U12706 (N_12706,N_12171,N_12033);
and U12707 (N_12707,N_12093,N_12221);
and U12708 (N_12708,N_12486,N_12015);
nand U12709 (N_12709,N_12027,N_12001);
nand U12710 (N_12710,N_12247,N_12008);
xor U12711 (N_12711,N_12118,N_12026);
nand U12712 (N_12712,N_12322,N_12425);
nor U12713 (N_12713,N_12172,N_12492);
or U12714 (N_12714,N_12421,N_12182);
or U12715 (N_12715,N_12140,N_12157);
nor U12716 (N_12716,N_12004,N_12119);
xnor U12717 (N_12717,N_12210,N_12083);
nor U12718 (N_12718,N_12228,N_12028);
xnor U12719 (N_12719,N_12402,N_12022);
xor U12720 (N_12720,N_12114,N_12070);
nand U12721 (N_12721,N_12012,N_12010);
nor U12722 (N_12722,N_12051,N_12408);
xor U12723 (N_12723,N_12474,N_12432);
and U12724 (N_12724,N_12377,N_12269);
and U12725 (N_12725,N_12218,N_12380);
xor U12726 (N_12726,N_12291,N_12449);
xor U12727 (N_12727,N_12058,N_12132);
xor U12728 (N_12728,N_12143,N_12092);
nor U12729 (N_12729,N_12149,N_12169);
nand U12730 (N_12730,N_12047,N_12226);
or U12731 (N_12731,N_12043,N_12023);
xnor U12732 (N_12732,N_12002,N_12392);
nor U12733 (N_12733,N_12074,N_12287);
nor U12734 (N_12734,N_12108,N_12448);
or U12735 (N_12735,N_12245,N_12016);
xor U12736 (N_12736,N_12126,N_12396);
or U12737 (N_12737,N_12368,N_12435);
and U12738 (N_12738,N_12434,N_12261);
xnor U12739 (N_12739,N_12046,N_12295);
and U12740 (N_12740,N_12220,N_12085);
xnor U12741 (N_12741,N_12306,N_12385);
xor U12742 (N_12742,N_12340,N_12358);
nor U12743 (N_12743,N_12071,N_12174);
nor U12744 (N_12744,N_12438,N_12251);
xor U12745 (N_12745,N_12206,N_12489);
or U12746 (N_12746,N_12423,N_12422);
xnor U12747 (N_12747,N_12150,N_12136);
or U12748 (N_12748,N_12481,N_12361);
xor U12749 (N_12749,N_12073,N_12077);
nand U12750 (N_12750,N_12494,N_12019);
xor U12751 (N_12751,N_12174,N_12011);
nand U12752 (N_12752,N_12103,N_12341);
or U12753 (N_12753,N_12271,N_12215);
nand U12754 (N_12754,N_12046,N_12058);
nand U12755 (N_12755,N_12288,N_12392);
nor U12756 (N_12756,N_12499,N_12097);
and U12757 (N_12757,N_12197,N_12391);
or U12758 (N_12758,N_12494,N_12253);
and U12759 (N_12759,N_12123,N_12488);
nor U12760 (N_12760,N_12462,N_12295);
nor U12761 (N_12761,N_12035,N_12078);
nor U12762 (N_12762,N_12439,N_12191);
nand U12763 (N_12763,N_12226,N_12421);
nor U12764 (N_12764,N_12005,N_12022);
xnor U12765 (N_12765,N_12155,N_12080);
xor U12766 (N_12766,N_12254,N_12394);
or U12767 (N_12767,N_12041,N_12376);
or U12768 (N_12768,N_12141,N_12133);
xor U12769 (N_12769,N_12001,N_12489);
nand U12770 (N_12770,N_12471,N_12198);
nor U12771 (N_12771,N_12081,N_12295);
xor U12772 (N_12772,N_12241,N_12084);
nand U12773 (N_12773,N_12306,N_12394);
nor U12774 (N_12774,N_12209,N_12479);
or U12775 (N_12775,N_12474,N_12472);
nand U12776 (N_12776,N_12275,N_12195);
nand U12777 (N_12777,N_12138,N_12148);
or U12778 (N_12778,N_12284,N_12138);
and U12779 (N_12779,N_12438,N_12155);
xnor U12780 (N_12780,N_12263,N_12070);
and U12781 (N_12781,N_12442,N_12429);
and U12782 (N_12782,N_12104,N_12261);
or U12783 (N_12783,N_12263,N_12124);
or U12784 (N_12784,N_12326,N_12092);
xor U12785 (N_12785,N_12439,N_12120);
xor U12786 (N_12786,N_12199,N_12165);
xnor U12787 (N_12787,N_12184,N_12140);
nor U12788 (N_12788,N_12153,N_12138);
nand U12789 (N_12789,N_12299,N_12225);
or U12790 (N_12790,N_12307,N_12186);
and U12791 (N_12791,N_12321,N_12094);
xnor U12792 (N_12792,N_12339,N_12397);
xnor U12793 (N_12793,N_12274,N_12483);
or U12794 (N_12794,N_12441,N_12056);
and U12795 (N_12795,N_12492,N_12229);
and U12796 (N_12796,N_12017,N_12387);
and U12797 (N_12797,N_12157,N_12309);
nor U12798 (N_12798,N_12281,N_12237);
or U12799 (N_12799,N_12067,N_12097);
or U12800 (N_12800,N_12230,N_12161);
nor U12801 (N_12801,N_12462,N_12439);
and U12802 (N_12802,N_12068,N_12444);
nand U12803 (N_12803,N_12012,N_12195);
nand U12804 (N_12804,N_12040,N_12255);
nand U12805 (N_12805,N_12464,N_12117);
or U12806 (N_12806,N_12389,N_12058);
or U12807 (N_12807,N_12334,N_12007);
nor U12808 (N_12808,N_12364,N_12294);
or U12809 (N_12809,N_12237,N_12179);
xnor U12810 (N_12810,N_12396,N_12171);
nand U12811 (N_12811,N_12167,N_12337);
xnor U12812 (N_12812,N_12270,N_12453);
xor U12813 (N_12813,N_12157,N_12243);
nor U12814 (N_12814,N_12211,N_12493);
nor U12815 (N_12815,N_12324,N_12442);
xor U12816 (N_12816,N_12490,N_12066);
or U12817 (N_12817,N_12395,N_12093);
nand U12818 (N_12818,N_12183,N_12179);
or U12819 (N_12819,N_12375,N_12015);
nand U12820 (N_12820,N_12366,N_12264);
nand U12821 (N_12821,N_12088,N_12165);
xor U12822 (N_12822,N_12375,N_12335);
or U12823 (N_12823,N_12234,N_12276);
or U12824 (N_12824,N_12051,N_12192);
or U12825 (N_12825,N_12385,N_12487);
or U12826 (N_12826,N_12449,N_12212);
xor U12827 (N_12827,N_12304,N_12288);
and U12828 (N_12828,N_12216,N_12051);
xnor U12829 (N_12829,N_12086,N_12379);
nor U12830 (N_12830,N_12133,N_12209);
nand U12831 (N_12831,N_12201,N_12211);
and U12832 (N_12832,N_12308,N_12316);
nor U12833 (N_12833,N_12392,N_12049);
xnor U12834 (N_12834,N_12283,N_12342);
or U12835 (N_12835,N_12002,N_12042);
xor U12836 (N_12836,N_12068,N_12454);
nand U12837 (N_12837,N_12302,N_12471);
nor U12838 (N_12838,N_12283,N_12493);
nor U12839 (N_12839,N_12155,N_12398);
and U12840 (N_12840,N_12465,N_12230);
and U12841 (N_12841,N_12220,N_12160);
and U12842 (N_12842,N_12208,N_12487);
nand U12843 (N_12843,N_12279,N_12118);
nand U12844 (N_12844,N_12040,N_12046);
xnor U12845 (N_12845,N_12305,N_12216);
or U12846 (N_12846,N_12231,N_12149);
xnor U12847 (N_12847,N_12003,N_12434);
and U12848 (N_12848,N_12170,N_12290);
and U12849 (N_12849,N_12147,N_12014);
nand U12850 (N_12850,N_12316,N_12485);
and U12851 (N_12851,N_12387,N_12022);
nor U12852 (N_12852,N_12057,N_12142);
nand U12853 (N_12853,N_12428,N_12418);
or U12854 (N_12854,N_12249,N_12360);
or U12855 (N_12855,N_12103,N_12160);
nor U12856 (N_12856,N_12441,N_12101);
and U12857 (N_12857,N_12422,N_12146);
and U12858 (N_12858,N_12080,N_12466);
xnor U12859 (N_12859,N_12176,N_12393);
nor U12860 (N_12860,N_12261,N_12150);
and U12861 (N_12861,N_12014,N_12372);
xnor U12862 (N_12862,N_12175,N_12352);
nand U12863 (N_12863,N_12431,N_12495);
xnor U12864 (N_12864,N_12210,N_12284);
and U12865 (N_12865,N_12247,N_12244);
nor U12866 (N_12866,N_12481,N_12262);
nor U12867 (N_12867,N_12059,N_12213);
nor U12868 (N_12868,N_12434,N_12086);
and U12869 (N_12869,N_12183,N_12019);
or U12870 (N_12870,N_12326,N_12455);
nand U12871 (N_12871,N_12380,N_12272);
or U12872 (N_12872,N_12073,N_12193);
or U12873 (N_12873,N_12117,N_12488);
nand U12874 (N_12874,N_12337,N_12350);
and U12875 (N_12875,N_12224,N_12343);
or U12876 (N_12876,N_12494,N_12037);
nand U12877 (N_12877,N_12469,N_12435);
or U12878 (N_12878,N_12112,N_12235);
nor U12879 (N_12879,N_12426,N_12015);
nor U12880 (N_12880,N_12457,N_12480);
and U12881 (N_12881,N_12043,N_12429);
xnor U12882 (N_12882,N_12252,N_12333);
and U12883 (N_12883,N_12281,N_12251);
and U12884 (N_12884,N_12334,N_12450);
xnor U12885 (N_12885,N_12287,N_12127);
and U12886 (N_12886,N_12177,N_12380);
nand U12887 (N_12887,N_12461,N_12080);
or U12888 (N_12888,N_12344,N_12477);
xnor U12889 (N_12889,N_12062,N_12347);
nor U12890 (N_12890,N_12009,N_12164);
or U12891 (N_12891,N_12376,N_12356);
or U12892 (N_12892,N_12279,N_12490);
nor U12893 (N_12893,N_12103,N_12305);
and U12894 (N_12894,N_12413,N_12062);
nand U12895 (N_12895,N_12220,N_12427);
xor U12896 (N_12896,N_12090,N_12184);
or U12897 (N_12897,N_12266,N_12119);
and U12898 (N_12898,N_12324,N_12388);
or U12899 (N_12899,N_12467,N_12374);
or U12900 (N_12900,N_12316,N_12208);
nand U12901 (N_12901,N_12208,N_12453);
nand U12902 (N_12902,N_12114,N_12044);
nand U12903 (N_12903,N_12467,N_12488);
nand U12904 (N_12904,N_12428,N_12332);
xor U12905 (N_12905,N_12249,N_12398);
or U12906 (N_12906,N_12022,N_12278);
or U12907 (N_12907,N_12105,N_12236);
or U12908 (N_12908,N_12452,N_12050);
or U12909 (N_12909,N_12401,N_12085);
or U12910 (N_12910,N_12440,N_12132);
nor U12911 (N_12911,N_12143,N_12389);
nor U12912 (N_12912,N_12430,N_12395);
or U12913 (N_12913,N_12413,N_12022);
nor U12914 (N_12914,N_12478,N_12373);
nand U12915 (N_12915,N_12029,N_12387);
and U12916 (N_12916,N_12219,N_12283);
and U12917 (N_12917,N_12407,N_12476);
nand U12918 (N_12918,N_12376,N_12233);
xor U12919 (N_12919,N_12153,N_12434);
and U12920 (N_12920,N_12289,N_12443);
xnor U12921 (N_12921,N_12357,N_12343);
or U12922 (N_12922,N_12169,N_12400);
and U12923 (N_12923,N_12346,N_12105);
or U12924 (N_12924,N_12442,N_12217);
xnor U12925 (N_12925,N_12443,N_12305);
nand U12926 (N_12926,N_12208,N_12266);
xnor U12927 (N_12927,N_12051,N_12188);
xor U12928 (N_12928,N_12385,N_12266);
xnor U12929 (N_12929,N_12300,N_12098);
and U12930 (N_12930,N_12395,N_12472);
and U12931 (N_12931,N_12053,N_12253);
or U12932 (N_12932,N_12325,N_12200);
nor U12933 (N_12933,N_12427,N_12223);
xor U12934 (N_12934,N_12415,N_12336);
and U12935 (N_12935,N_12284,N_12047);
and U12936 (N_12936,N_12332,N_12392);
nor U12937 (N_12937,N_12258,N_12401);
nor U12938 (N_12938,N_12093,N_12003);
nor U12939 (N_12939,N_12149,N_12102);
nor U12940 (N_12940,N_12289,N_12439);
nand U12941 (N_12941,N_12442,N_12204);
nor U12942 (N_12942,N_12071,N_12388);
nor U12943 (N_12943,N_12285,N_12383);
nor U12944 (N_12944,N_12360,N_12317);
and U12945 (N_12945,N_12070,N_12201);
nor U12946 (N_12946,N_12096,N_12428);
nand U12947 (N_12947,N_12062,N_12003);
or U12948 (N_12948,N_12137,N_12177);
nor U12949 (N_12949,N_12494,N_12495);
xor U12950 (N_12950,N_12297,N_12232);
nor U12951 (N_12951,N_12028,N_12054);
nor U12952 (N_12952,N_12479,N_12194);
and U12953 (N_12953,N_12178,N_12154);
nand U12954 (N_12954,N_12020,N_12374);
xnor U12955 (N_12955,N_12202,N_12371);
xnor U12956 (N_12956,N_12247,N_12070);
xnor U12957 (N_12957,N_12155,N_12012);
nor U12958 (N_12958,N_12166,N_12284);
or U12959 (N_12959,N_12444,N_12265);
nand U12960 (N_12960,N_12094,N_12050);
and U12961 (N_12961,N_12303,N_12234);
nor U12962 (N_12962,N_12128,N_12081);
or U12963 (N_12963,N_12023,N_12385);
nand U12964 (N_12964,N_12213,N_12347);
nor U12965 (N_12965,N_12493,N_12409);
xnor U12966 (N_12966,N_12072,N_12231);
xor U12967 (N_12967,N_12356,N_12318);
xnor U12968 (N_12968,N_12369,N_12253);
nand U12969 (N_12969,N_12227,N_12123);
or U12970 (N_12970,N_12425,N_12309);
nand U12971 (N_12971,N_12041,N_12372);
nor U12972 (N_12972,N_12047,N_12399);
xor U12973 (N_12973,N_12402,N_12031);
nand U12974 (N_12974,N_12210,N_12368);
or U12975 (N_12975,N_12317,N_12071);
or U12976 (N_12976,N_12430,N_12398);
and U12977 (N_12977,N_12152,N_12160);
or U12978 (N_12978,N_12305,N_12170);
nand U12979 (N_12979,N_12439,N_12310);
nor U12980 (N_12980,N_12079,N_12040);
xor U12981 (N_12981,N_12328,N_12356);
nor U12982 (N_12982,N_12376,N_12479);
and U12983 (N_12983,N_12163,N_12013);
nand U12984 (N_12984,N_12382,N_12075);
nor U12985 (N_12985,N_12398,N_12484);
nor U12986 (N_12986,N_12465,N_12166);
nand U12987 (N_12987,N_12087,N_12417);
nand U12988 (N_12988,N_12313,N_12405);
nor U12989 (N_12989,N_12493,N_12216);
and U12990 (N_12990,N_12216,N_12274);
or U12991 (N_12991,N_12064,N_12430);
xnor U12992 (N_12992,N_12333,N_12355);
nand U12993 (N_12993,N_12246,N_12346);
nor U12994 (N_12994,N_12467,N_12446);
nor U12995 (N_12995,N_12097,N_12386);
xnor U12996 (N_12996,N_12046,N_12024);
nor U12997 (N_12997,N_12183,N_12370);
nor U12998 (N_12998,N_12357,N_12042);
xnor U12999 (N_12999,N_12085,N_12112);
nand U13000 (N_13000,N_12970,N_12616);
xor U13001 (N_13001,N_12750,N_12764);
xnor U13002 (N_13002,N_12996,N_12737);
xor U13003 (N_13003,N_12515,N_12520);
xor U13004 (N_13004,N_12783,N_12661);
or U13005 (N_13005,N_12571,N_12686);
nand U13006 (N_13006,N_12842,N_12554);
nor U13007 (N_13007,N_12645,N_12572);
or U13008 (N_13008,N_12672,N_12622);
nor U13009 (N_13009,N_12684,N_12723);
xor U13010 (N_13010,N_12959,N_12594);
or U13011 (N_13011,N_12745,N_12674);
xnor U13012 (N_13012,N_12906,N_12696);
or U13013 (N_13013,N_12564,N_12715);
or U13014 (N_13014,N_12628,N_12759);
nand U13015 (N_13015,N_12608,N_12943);
and U13016 (N_13016,N_12631,N_12518);
xnor U13017 (N_13017,N_12688,N_12530);
and U13018 (N_13018,N_12802,N_12738);
nor U13019 (N_13019,N_12597,N_12523);
nor U13020 (N_13020,N_12853,N_12944);
or U13021 (N_13021,N_12805,N_12614);
and U13022 (N_13022,N_12820,N_12592);
xnor U13023 (N_13023,N_12671,N_12990);
and U13024 (N_13024,N_12877,N_12505);
xnor U13025 (N_13025,N_12639,N_12563);
and U13026 (N_13026,N_12956,N_12690);
or U13027 (N_13027,N_12543,N_12620);
nor U13028 (N_13028,N_12646,N_12985);
and U13029 (N_13029,N_12630,N_12559);
nor U13030 (N_13030,N_12579,N_12586);
and U13031 (N_13031,N_12643,N_12799);
nand U13032 (N_13032,N_12937,N_12514);
and U13033 (N_13033,N_12891,N_12606);
nand U13034 (N_13034,N_12811,N_12555);
nor U13035 (N_13035,N_12871,N_12786);
nand U13036 (N_13036,N_12742,N_12668);
nor U13037 (N_13037,N_12950,N_12755);
nor U13038 (N_13038,N_12829,N_12741);
or U13039 (N_13039,N_12790,N_12733);
and U13040 (N_13040,N_12940,N_12503);
nand U13041 (N_13041,N_12669,N_12912);
or U13042 (N_13042,N_12699,N_12854);
nor U13043 (N_13043,N_12731,N_12659);
or U13044 (N_13044,N_12525,N_12581);
nand U13045 (N_13045,N_12859,N_12792);
xnor U13046 (N_13046,N_12968,N_12734);
nor U13047 (N_13047,N_12513,N_12654);
xnor U13048 (N_13048,N_12774,N_12747);
nor U13049 (N_13049,N_12640,N_12595);
nand U13050 (N_13050,N_12857,N_12584);
nor U13051 (N_13051,N_12587,N_12813);
nand U13052 (N_13052,N_12931,N_12568);
nand U13053 (N_13053,N_12965,N_12839);
nand U13054 (N_13054,N_12617,N_12508);
or U13055 (N_13055,N_12962,N_12512);
and U13056 (N_13056,N_12975,N_12627);
or U13057 (N_13057,N_12702,N_12652);
nand U13058 (N_13058,N_12547,N_12718);
nand U13059 (N_13059,N_12504,N_12717);
nor U13060 (N_13060,N_12952,N_12576);
and U13061 (N_13061,N_12551,N_12847);
xnor U13062 (N_13062,N_12872,N_12934);
xnor U13063 (N_13063,N_12585,N_12607);
xor U13064 (N_13064,N_12549,N_12719);
xnor U13065 (N_13065,N_12830,N_12921);
nand U13066 (N_13066,N_12787,N_12818);
nor U13067 (N_13067,N_12634,N_12981);
nor U13068 (N_13068,N_12812,N_12574);
and U13069 (N_13069,N_12889,N_12960);
and U13070 (N_13070,N_12920,N_12822);
or U13071 (N_13071,N_12983,N_12649);
nand U13072 (N_13072,N_12929,N_12936);
xor U13073 (N_13073,N_12991,N_12545);
and U13074 (N_13074,N_12516,N_12544);
nor U13075 (N_13075,N_12570,N_12957);
nand U13076 (N_13076,N_12838,N_12771);
and U13077 (N_13077,N_12900,N_12775);
and U13078 (N_13078,N_12843,N_12782);
nor U13079 (N_13079,N_12966,N_12511);
nor U13080 (N_13080,N_12765,N_12914);
xor U13081 (N_13081,N_12548,N_12507);
nor U13082 (N_13082,N_12724,N_12501);
xor U13083 (N_13083,N_12806,N_12602);
nor U13084 (N_13084,N_12666,N_12899);
and U13085 (N_13085,N_12730,N_12770);
or U13086 (N_13086,N_12561,N_12777);
xor U13087 (N_13087,N_12817,N_12815);
or U13088 (N_13088,N_12835,N_12919);
and U13089 (N_13089,N_12685,N_12837);
or U13090 (N_13090,N_12867,N_12667);
and U13091 (N_13091,N_12946,N_12658);
nor U13092 (N_13092,N_12863,N_12677);
or U13093 (N_13093,N_12788,N_12762);
or U13094 (N_13094,N_12687,N_12908);
nand U13095 (N_13095,N_12612,N_12884);
nand U13096 (N_13096,N_12673,N_12540);
nor U13097 (N_13097,N_12632,N_12746);
or U13098 (N_13098,N_12998,N_12917);
or U13099 (N_13099,N_12691,N_12605);
nor U13100 (N_13100,N_12532,N_12633);
nor U13101 (N_13101,N_12763,N_12648);
and U13102 (N_13102,N_12980,N_12735);
and U13103 (N_13103,N_12729,N_12878);
or U13104 (N_13104,N_12744,N_12825);
or U13105 (N_13105,N_12541,N_12767);
nand U13106 (N_13106,N_12714,N_12573);
xnor U13107 (N_13107,N_12697,N_12938);
or U13108 (N_13108,N_12828,N_12973);
or U13109 (N_13109,N_12798,N_12720);
xnor U13110 (N_13110,N_12675,N_12641);
or U13111 (N_13111,N_12901,N_12947);
nand U13112 (N_13112,N_12880,N_12888);
nor U13113 (N_13113,N_12550,N_12784);
and U13114 (N_13114,N_12862,N_12961);
and U13115 (N_13115,N_12848,N_12749);
nand U13116 (N_13116,N_12604,N_12701);
xnor U13117 (N_13117,N_12580,N_12683);
xor U13118 (N_13118,N_12909,N_12955);
or U13119 (N_13119,N_12995,N_12809);
and U13120 (N_13120,N_12689,N_12926);
xnor U13121 (N_13121,N_12752,N_12986);
nand U13122 (N_13122,N_12542,N_12974);
nand U13123 (N_13123,N_12716,N_12932);
and U13124 (N_13124,N_12754,N_12897);
and U13125 (N_13125,N_12886,N_12949);
nand U13126 (N_13126,N_12819,N_12567);
and U13127 (N_13127,N_12560,N_12904);
or U13128 (N_13128,N_12760,N_12610);
and U13129 (N_13129,N_12660,N_12893);
or U13130 (N_13130,N_12533,N_12976);
nor U13131 (N_13131,N_12922,N_12722);
nor U13132 (N_13132,N_12903,N_12521);
xnor U13133 (N_13133,N_12902,N_12836);
or U13134 (N_13134,N_12693,N_12662);
nand U13135 (N_13135,N_12933,N_12870);
nor U13136 (N_13136,N_12681,N_12858);
and U13137 (N_13137,N_12528,N_12558);
nand U13138 (N_13138,N_12779,N_12682);
xor U13139 (N_13139,N_12539,N_12565);
nor U13140 (N_13140,N_12789,N_12500);
and U13141 (N_13141,N_12624,N_12849);
and U13142 (N_13142,N_12844,N_12566);
nor U13143 (N_13143,N_12776,N_12856);
and U13144 (N_13144,N_12865,N_12885);
and U13145 (N_13145,N_12845,N_12653);
or U13146 (N_13146,N_12527,N_12892);
nand U13147 (N_13147,N_12999,N_12502);
nand U13148 (N_13148,N_12625,N_12941);
or U13149 (N_13149,N_12993,N_12954);
and U13150 (N_13150,N_12656,N_12948);
nand U13151 (N_13151,N_12827,N_12953);
nor U13152 (N_13152,N_12876,N_12930);
and U13153 (N_13153,N_12894,N_12619);
nand U13154 (N_13154,N_12562,N_12583);
or U13155 (N_13155,N_12650,N_12589);
and U13156 (N_13156,N_12978,N_12538);
nor U13157 (N_13157,N_12757,N_12772);
nand U13158 (N_13158,N_12773,N_12593);
xor U13159 (N_13159,N_12510,N_12846);
or U13160 (N_13160,N_12740,N_12860);
or U13161 (N_13161,N_12637,N_12728);
xor U13162 (N_13162,N_12801,N_12778);
and U13163 (N_13163,N_12705,N_12826);
and U13164 (N_13164,N_12866,N_12569);
nand U13165 (N_13165,N_12800,N_12869);
xnor U13166 (N_13166,N_12536,N_12824);
xnor U13167 (N_13167,N_12879,N_12793);
or U13168 (N_13168,N_12972,N_12881);
and U13169 (N_13169,N_12713,N_12781);
nand U13170 (N_13170,N_12522,N_12939);
xor U13171 (N_13171,N_12651,N_12599);
and U13172 (N_13172,N_12678,N_12517);
or U13173 (N_13173,N_12794,N_12935);
nor U13174 (N_13174,N_12761,N_12623);
xnor U13175 (N_13175,N_12924,N_12618);
nor U13176 (N_13176,N_12708,N_12964);
and U13177 (N_13177,N_12552,N_12994);
nand U13178 (N_13178,N_12911,N_12875);
nand U13179 (N_13179,N_12663,N_12832);
nand U13180 (N_13180,N_12590,N_12615);
or U13181 (N_13181,N_12557,N_12913);
and U13182 (N_13182,N_12706,N_12537);
nor U13183 (N_13183,N_12841,N_12647);
or U13184 (N_13184,N_12664,N_12732);
or U13185 (N_13185,N_12700,N_12577);
and U13186 (N_13186,N_12905,N_12785);
xor U13187 (N_13187,N_12709,N_12600);
nor U13188 (N_13188,N_12916,N_12780);
nor U13189 (N_13189,N_12636,N_12629);
nor U13190 (N_13190,N_12851,N_12670);
xor U13191 (N_13191,N_12804,N_12655);
xnor U13192 (N_13192,N_12534,N_12831);
or U13193 (N_13193,N_12766,N_12603);
nand U13194 (N_13194,N_12553,N_12868);
xor U13195 (N_13195,N_12910,N_12598);
xor U13196 (N_13196,N_12694,N_12751);
xnor U13197 (N_13197,N_12963,N_12601);
xor U13198 (N_13198,N_12613,N_12987);
nand U13199 (N_13199,N_12808,N_12873);
or U13200 (N_13200,N_12967,N_12797);
and U13201 (N_13201,N_12834,N_12582);
and U13202 (N_13202,N_12882,N_12642);
or U13203 (N_13203,N_12861,N_12918);
or U13204 (N_13204,N_12840,N_12971);
nor U13205 (N_13205,N_12529,N_12852);
nor U13206 (N_13206,N_12988,N_12942);
nor U13207 (N_13207,N_12923,N_12864);
nand U13208 (N_13208,N_12644,N_12524);
xor U13209 (N_13209,N_12748,N_12578);
and U13210 (N_13210,N_12997,N_12707);
nor U13211 (N_13211,N_12575,N_12739);
or U13212 (N_13212,N_12925,N_12814);
nor U13213 (N_13213,N_12611,N_12726);
xor U13214 (N_13214,N_12890,N_12526);
nand U13215 (N_13215,N_12769,N_12833);
nor U13216 (N_13216,N_12756,N_12768);
and U13217 (N_13217,N_12704,N_12895);
or U13218 (N_13218,N_12535,N_12509);
xnor U13219 (N_13219,N_12743,N_12977);
or U13220 (N_13220,N_12855,N_12657);
and U13221 (N_13221,N_12823,N_12591);
xnor U13222 (N_13222,N_12887,N_12519);
and U13223 (N_13223,N_12638,N_12821);
or U13224 (N_13224,N_12989,N_12758);
and U13225 (N_13225,N_12795,N_12807);
nor U13226 (N_13226,N_12915,N_12703);
and U13227 (N_13227,N_12609,N_12736);
nand U13228 (N_13228,N_12898,N_12979);
xor U13229 (N_13229,N_12710,N_12679);
nor U13230 (N_13230,N_12588,N_12816);
or U13231 (N_13231,N_12928,N_12907);
and U13232 (N_13232,N_12711,N_12665);
nor U13233 (N_13233,N_12596,N_12621);
nor U13234 (N_13234,N_12531,N_12721);
nor U13235 (N_13235,N_12883,N_12626);
and U13236 (N_13236,N_12992,N_12680);
or U13237 (N_13237,N_12753,N_12969);
or U13238 (N_13238,N_12698,N_12927);
nor U13239 (N_13239,N_12676,N_12556);
nand U13240 (N_13240,N_12945,N_12712);
nor U13241 (N_13241,N_12896,N_12850);
or U13242 (N_13242,N_12506,N_12874);
nor U13243 (N_13243,N_12692,N_12810);
nor U13244 (N_13244,N_12951,N_12984);
xor U13245 (N_13245,N_12695,N_12546);
nand U13246 (N_13246,N_12725,N_12791);
and U13247 (N_13247,N_12958,N_12803);
nand U13248 (N_13248,N_12982,N_12635);
and U13249 (N_13249,N_12796,N_12727);
xnor U13250 (N_13250,N_12730,N_12867);
nand U13251 (N_13251,N_12503,N_12973);
and U13252 (N_13252,N_12515,N_12985);
nand U13253 (N_13253,N_12792,N_12519);
and U13254 (N_13254,N_12643,N_12889);
xor U13255 (N_13255,N_12735,N_12717);
and U13256 (N_13256,N_12624,N_12677);
xor U13257 (N_13257,N_12540,N_12812);
and U13258 (N_13258,N_12586,N_12707);
nand U13259 (N_13259,N_12718,N_12517);
xnor U13260 (N_13260,N_12713,N_12864);
xnor U13261 (N_13261,N_12643,N_12577);
and U13262 (N_13262,N_12745,N_12805);
or U13263 (N_13263,N_12656,N_12772);
and U13264 (N_13264,N_12569,N_12912);
xor U13265 (N_13265,N_12524,N_12841);
xor U13266 (N_13266,N_12581,N_12981);
nor U13267 (N_13267,N_12709,N_12960);
or U13268 (N_13268,N_12897,N_12624);
xnor U13269 (N_13269,N_12913,N_12686);
nand U13270 (N_13270,N_12795,N_12566);
nor U13271 (N_13271,N_12579,N_12913);
or U13272 (N_13272,N_12606,N_12686);
nand U13273 (N_13273,N_12522,N_12862);
and U13274 (N_13274,N_12962,N_12753);
nor U13275 (N_13275,N_12634,N_12970);
nor U13276 (N_13276,N_12635,N_12548);
xnor U13277 (N_13277,N_12992,N_12845);
and U13278 (N_13278,N_12572,N_12735);
xnor U13279 (N_13279,N_12506,N_12695);
xnor U13280 (N_13280,N_12986,N_12690);
nor U13281 (N_13281,N_12526,N_12628);
or U13282 (N_13282,N_12546,N_12560);
xnor U13283 (N_13283,N_12931,N_12870);
and U13284 (N_13284,N_12807,N_12910);
xnor U13285 (N_13285,N_12993,N_12791);
nor U13286 (N_13286,N_12711,N_12911);
nor U13287 (N_13287,N_12594,N_12645);
and U13288 (N_13288,N_12961,N_12619);
xnor U13289 (N_13289,N_12727,N_12580);
nand U13290 (N_13290,N_12579,N_12710);
nand U13291 (N_13291,N_12727,N_12681);
nor U13292 (N_13292,N_12737,N_12975);
and U13293 (N_13293,N_12576,N_12795);
and U13294 (N_13294,N_12877,N_12570);
nor U13295 (N_13295,N_12576,N_12510);
nor U13296 (N_13296,N_12844,N_12710);
nor U13297 (N_13297,N_12690,N_12657);
or U13298 (N_13298,N_12951,N_12658);
nand U13299 (N_13299,N_12626,N_12786);
nand U13300 (N_13300,N_12685,N_12813);
nor U13301 (N_13301,N_12516,N_12807);
or U13302 (N_13302,N_12958,N_12544);
xor U13303 (N_13303,N_12633,N_12719);
nand U13304 (N_13304,N_12798,N_12997);
or U13305 (N_13305,N_12710,N_12727);
and U13306 (N_13306,N_12665,N_12503);
nor U13307 (N_13307,N_12838,N_12834);
nand U13308 (N_13308,N_12637,N_12833);
or U13309 (N_13309,N_12847,N_12790);
and U13310 (N_13310,N_12627,N_12599);
or U13311 (N_13311,N_12732,N_12546);
nand U13312 (N_13312,N_12827,N_12869);
and U13313 (N_13313,N_12594,N_12766);
xor U13314 (N_13314,N_12718,N_12515);
and U13315 (N_13315,N_12850,N_12529);
nand U13316 (N_13316,N_12835,N_12809);
and U13317 (N_13317,N_12575,N_12729);
and U13318 (N_13318,N_12779,N_12573);
and U13319 (N_13319,N_12712,N_12951);
and U13320 (N_13320,N_12985,N_12956);
and U13321 (N_13321,N_12508,N_12739);
and U13322 (N_13322,N_12567,N_12595);
nor U13323 (N_13323,N_12695,N_12934);
and U13324 (N_13324,N_12931,N_12728);
xor U13325 (N_13325,N_12867,N_12626);
nor U13326 (N_13326,N_12809,N_12846);
nand U13327 (N_13327,N_12987,N_12810);
and U13328 (N_13328,N_12794,N_12641);
xnor U13329 (N_13329,N_12884,N_12583);
or U13330 (N_13330,N_12774,N_12617);
nor U13331 (N_13331,N_12584,N_12571);
nor U13332 (N_13332,N_12633,N_12991);
nor U13333 (N_13333,N_12964,N_12617);
nand U13334 (N_13334,N_12876,N_12754);
xor U13335 (N_13335,N_12966,N_12946);
xor U13336 (N_13336,N_12693,N_12579);
nand U13337 (N_13337,N_12668,N_12565);
nand U13338 (N_13338,N_12604,N_12732);
or U13339 (N_13339,N_12681,N_12609);
nor U13340 (N_13340,N_12579,N_12949);
nor U13341 (N_13341,N_12967,N_12779);
nand U13342 (N_13342,N_12844,N_12508);
or U13343 (N_13343,N_12739,N_12548);
nand U13344 (N_13344,N_12588,N_12804);
or U13345 (N_13345,N_12585,N_12708);
and U13346 (N_13346,N_12914,N_12814);
and U13347 (N_13347,N_12794,N_12924);
nor U13348 (N_13348,N_12560,N_12828);
nor U13349 (N_13349,N_12803,N_12928);
xor U13350 (N_13350,N_12522,N_12904);
and U13351 (N_13351,N_12815,N_12744);
xnor U13352 (N_13352,N_12860,N_12849);
and U13353 (N_13353,N_12685,N_12993);
xor U13354 (N_13354,N_12786,N_12998);
nand U13355 (N_13355,N_12538,N_12952);
nor U13356 (N_13356,N_12994,N_12638);
xnor U13357 (N_13357,N_12653,N_12838);
and U13358 (N_13358,N_12803,N_12584);
and U13359 (N_13359,N_12830,N_12849);
xor U13360 (N_13360,N_12558,N_12666);
or U13361 (N_13361,N_12971,N_12818);
nand U13362 (N_13362,N_12881,N_12663);
xor U13363 (N_13363,N_12939,N_12783);
or U13364 (N_13364,N_12954,N_12902);
nor U13365 (N_13365,N_12918,N_12679);
or U13366 (N_13366,N_12968,N_12993);
or U13367 (N_13367,N_12541,N_12868);
nor U13368 (N_13368,N_12907,N_12534);
nand U13369 (N_13369,N_12988,N_12998);
xor U13370 (N_13370,N_12552,N_12963);
and U13371 (N_13371,N_12625,N_12635);
xor U13372 (N_13372,N_12590,N_12761);
xor U13373 (N_13373,N_12648,N_12732);
xor U13374 (N_13374,N_12876,N_12674);
nand U13375 (N_13375,N_12776,N_12658);
or U13376 (N_13376,N_12671,N_12649);
or U13377 (N_13377,N_12909,N_12934);
xnor U13378 (N_13378,N_12873,N_12778);
nand U13379 (N_13379,N_12538,N_12923);
or U13380 (N_13380,N_12847,N_12716);
and U13381 (N_13381,N_12817,N_12942);
nor U13382 (N_13382,N_12807,N_12652);
nand U13383 (N_13383,N_12688,N_12592);
and U13384 (N_13384,N_12514,N_12627);
nor U13385 (N_13385,N_12942,N_12669);
xor U13386 (N_13386,N_12552,N_12520);
xor U13387 (N_13387,N_12768,N_12769);
nor U13388 (N_13388,N_12718,N_12548);
nor U13389 (N_13389,N_12780,N_12867);
or U13390 (N_13390,N_12522,N_12658);
or U13391 (N_13391,N_12675,N_12533);
or U13392 (N_13392,N_12963,N_12844);
xor U13393 (N_13393,N_12698,N_12755);
and U13394 (N_13394,N_12873,N_12980);
nand U13395 (N_13395,N_12661,N_12751);
xnor U13396 (N_13396,N_12850,N_12861);
or U13397 (N_13397,N_12625,N_12533);
nor U13398 (N_13398,N_12815,N_12516);
or U13399 (N_13399,N_12535,N_12906);
and U13400 (N_13400,N_12980,N_12564);
nand U13401 (N_13401,N_12681,N_12995);
nor U13402 (N_13402,N_12971,N_12552);
and U13403 (N_13403,N_12860,N_12994);
and U13404 (N_13404,N_12646,N_12588);
and U13405 (N_13405,N_12608,N_12628);
nand U13406 (N_13406,N_12861,N_12982);
nor U13407 (N_13407,N_12884,N_12803);
nand U13408 (N_13408,N_12918,N_12505);
nor U13409 (N_13409,N_12607,N_12933);
and U13410 (N_13410,N_12521,N_12614);
and U13411 (N_13411,N_12747,N_12687);
nand U13412 (N_13412,N_12646,N_12848);
nor U13413 (N_13413,N_12921,N_12687);
and U13414 (N_13414,N_12678,N_12973);
or U13415 (N_13415,N_12954,N_12930);
or U13416 (N_13416,N_12828,N_12822);
nor U13417 (N_13417,N_12875,N_12500);
and U13418 (N_13418,N_12926,N_12768);
and U13419 (N_13419,N_12822,N_12981);
nand U13420 (N_13420,N_12935,N_12977);
nor U13421 (N_13421,N_12792,N_12709);
or U13422 (N_13422,N_12782,N_12716);
nor U13423 (N_13423,N_12707,N_12980);
xor U13424 (N_13424,N_12886,N_12726);
and U13425 (N_13425,N_12769,N_12842);
nor U13426 (N_13426,N_12785,N_12814);
nand U13427 (N_13427,N_12578,N_12686);
xnor U13428 (N_13428,N_12582,N_12659);
nor U13429 (N_13429,N_12664,N_12645);
nand U13430 (N_13430,N_12735,N_12931);
nand U13431 (N_13431,N_12964,N_12848);
and U13432 (N_13432,N_12947,N_12817);
xnor U13433 (N_13433,N_12706,N_12822);
nand U13434 (N_13434,N_12631,N_12705);
nand U13435 (N_13435,N_12985,N_12692);
nor U13436 (N_13436,N_12720,N_12597);
xor U13437 (N_13437,N_12769,N_12903);
nand U13438 (N_13438,N_12692,N_12767);
nor U13439 (N_13439,N_12562,N_12729);
nand U13440 (N_13440,N_12867,N_12546);
xnor U13441 (N_13441,N_12980,N_12721);
and U13442 (N_13442,N_12920,N_12710);
or U13443 (N_13443,N_12898,N_12813);
nand U13444 (N_13444,N_12596,N_12889);
and U13445 (N_13445,N_12728,N_12826);
xnor U13446 (N_13446,N_12618,N_12761);
nor U13447 (N_13447,N_12852,N_12896);
nand U13448 (N_13448,N_12635,N_12919);
xor U13449 (N_13449,N_12515,N_12646);
and U13450 (N_13450,N_12573,N_12570);
nand U13451 (N_13451,N_12916,N_12614);
and U13452 (N_13452,N_12610,N_12587);
xor U13453 (N_13453,N_12728,N_12571);
xor U13454 (N_13454,N_12917,N_12738);
xnor U13455 (N_13455,N_12980,N_12541);
or U13456 (N_13456,N_12947,N_12962);
nand U13457 (N_13457,N_12515,N_12777);
xnor U13458 (N_13458,N_12986,N_12853);
or U13459 (N_13459,N_12901,N_12990);
xnor U13460 (N_13460,N_12783,N_12882);
or U13461 (N_13461,N_12591,N_12830);
or U13462 (N_13462,N_12825,N_12815);
nand U13463 (N_13463,N_12601,N_12678);
xnor U13464 (N_13464,N_12996,N_12765);
nand U13465 (N_13465,N_12600,N_12505);
nand U13466 (N_13466,N_12712,N_12598);
xnor U13467 (N_13467,N_12517,N_12631);
nand U13468 (N_13468,N_12765,N_12745);
or U13469 (N_13469,N_12771,N_12736);
nand U13470 (N_13470,N_12837,N_12768);
xnor U13471 (N_13471,N_12541,N_12752);
nand U13472 (N_13472,N_12503,N_12620);
nor U13473 (N_13473,N_12802,N_12807);
and U13474 (N_13474,N_12821,N_12793);
nor U13475 (N_13475,N_12945,N_12606);
nand U13476 (N_13476,N_12521,N_12766);
nor U13477 (N_13477,N_12711,N_12747);
and U13478 (N_13478,N_12992,N_12868);
xnor U13479 (N_13479,N_12841,N_12876);
nand U13480 (N_13480,N_12949,N_12742);
or U13481 (N_13481,N_12748,N_12841);
xnor U13482 (N_13482,N_12513,N_12794);
nor U13483 (N_13483,N_12908,N_12904);
nand U13484 (N_13484,N_12503,N_12790);
nor U13485 (N_13485,N_12706,N_12873);
and U13486 (N_13486,N_12512,N_12532);
and U13487 (N_13487,N_12636,N_12974);
nand U13488 (N_13488,N_12625,N_12568);
or U13489 (N_13489,N_12912,N_12800);
and U13490 (N_13490,N_12821,N_12661);
or U13491 (N_13491,N_12674,N_12508);
or U13492 (N_13492,N_12780,N_12640);
nand U13493 (N_13493,N_12952,N_12551);
nor U13494 (N_13494,N_12612,N_12713);
xnor U13495 (N_13495,N_12553,N_12679);
nand U13496 (N_13496,N_12665,N_12622);
nand U13497 (N_13497,N_12541,N_12608);
or U13498 (N_13498,N_12803,N_12523);
or U13499 (N_13499,N_12725,N_12970);
xnor U13500 (N_13500,N_13204,N_13172);
nand U13501 (N_13501,N_13176,N_13296);
nor U13502 (N_13502,N_13441,N_13257);
nor U13503 (N_13503,N_13207,N_13114);
nor U13504 (N_13504,N_13115,N_13261);
nand U13505 (N_13505,N_13471,N_13369);
nor U13506 (N_13506,N_13111,N_13373);
and U13507 (N_13507,N_13436,N_13142);
xnor U13508 (N_13508,N_13028,N_13490);
nor U13509 (N_13509,N_13327,N_13360);
nor U13510 (N_13510,N_13250,N_13254);
nor U13511 (N_13511,N_13174,N_13316);
nand U13512 (N_13512,N_13492,N_13305);
and U13513 (N_13513,N_13046,N_13245);
xor U13514 (N_13514,N_13155,N_13399);
nor U13515 (N_13515,N_13255,N_13160);
xnor U13516 (N_13516,N_13145,N_13484);
xor U13517 (N_13517,N_13408,N_13166);
and U13518 (N_13518,N_13061,N_13454);
nand U13519 (N_13519,N_13129,N_13152);
nor U13520 (N_13520,N_13124,N_13417);
nor U13521 (N_13521,N_13081,N_13188);
or U13522 (N_13522,N_13354,N_13268);
xnor U13523 (N_13523,N_13322,N_13153);
and U13524 (N_13524,N_13428,N_13424);
or U13525 (N_13525,N_13384,N_13324);
nand U13526 (N_13526,N_13054,N_13089);
or U13527 (N_13527,N_13029,N_13213);
or U13528 (N_13528,N_13448,N_13333);
nor U13529 (N_13529,N_13258,N_13264);
xor U13530 (N_13530,N_13236,N_13049);
nand U13531 (N_13531,N_13367,N_13022);
nor U13532 (N_13532,N_13112,N_13456);
xnor U13533 (N_13533,N_13133,N_13475);
and U13534 (N_13534,N_13420,N_13064);
or U13535 (N_13535,N_13003,N_13170);
xnor U13536 (N_13536,N_13226,N_13286);
nor U13537 (N_13537,N_13234,N_13351);
and U13538 (N_13538,N_13498,N_13135);
and U13539 (N_13539,N_13389,N_13069);
and U13540 (N_13540,N_13410,N_13362);
xor U13541 (N_13541,N_13052,N_13229);
or U13542 (N_13542,N_13209,N_13335);
nor U13543 (N_13543,N_13210,N_13319);
and U13544 (N_13544,N_13165,N_13019);
nand U13545 (N_13545,N_13038,N_13192);
nor U13546 (N_13546,N_13223,N_13221);
and U13547 (N_13547,N_13307,N_13232);
nor U13548 (N_13548,N_13442,N_13096);
nand U13549 (N_13549,N_13489,N_13432);
or U13550 (N_13550,N_13073,N_13281);
xor U13551 (N_13551,N_13020,N_13464);
xnor U13552 (N_13552,N_13200,N_13119);
or U13553 (N_13553,N_13072,N_13405);
and U13554 (N_13554,N_13297,N_13010);
xor U13555 (N_13555,N_13211,N_13051);
xnor U13556 (N_13556,N_13128,N_13311);
xnor U13557 (N_13557,N_13121,N_13280);
and U13558 (N_13558,N_13308,N_13198);
and U13559 (N_13559,N_13274,N_13392);
or U13560 (N_13560,N_13108,N_13048);
nand U13561 (N_13561,N_13186,N_13034);
or U13562 (N_13562,N_13247,N_13080);
xnor U13563 (N_13563,N_13467,N_13380);
nor U13564 (N_13564,N_13491,N_13164);
and U13565 (N_13565,N_13196,N_13058);
nand U13566 (N_13566,N_13151,N_13159);
and U13567 (N_13567,N_13377,N_13091);
and U13568 (N_13568,N_13187,N_13149);
or U13569 (N_13569,N_13027,N_13162);
or U13570 (N_13570,N_13088,N_13090);
nand U13571 (N_13571,N_13497,N_13481);
xor U13572 (N_13572,N_13147,N_13256);
xor U13573 (N_13573,N_13318,N_13270);
nand U13574 (N_13574,N_13216,N_13055);
nand U13575 (N_13575,N_13295,N_13449);
and U13576 (N_13576,N_13169,N_13321);
or U13577 (N_13577,N_13004,N_13132);
nor U13578 (N_13578,N_13284,N_13314);
nand U13579 (N_13579,N_13079,N_13473);
or U13580 (N_13580,N_13341,N_13141);
or U13581 (N_13581,N_13348,N_13244);
nor U13582 (N_13582,N_13439,N_13383);
nor U13583 (N_13583,N_13451,N_13292);
or U13584 (N_13584,N_13134,N_13483);
or U13585 (N_13585,N_13304,N_13366);
nand U13586 (N_13586,N_13293,N_13440);
and U13587 (N_13587,N_13433,N_13037);
xnor U13588 (N_13588,N_13184,N_13370);
and U13589 (N_13589,N_13240,N_13237);
nor U13590 (N_13590,N_13302,N_13482);
or U13591 (N_13591,N_13418,N_13126);
nor U13592 (N_13592,N_13282,N_13182);
nand U13593 (N_13593,N_13263,N_13045);
or U13594 (N_13594,N_13138,N_13246);
and U13595 (N_13595,N_13390,N_13063);
nor U13596 (N_13596,N_13279,N_13336);
or U13597 (N_13597,N_13422,N_13397);
and U13598 (N_13598,N_13178,N_13154);
nor U13599 (N_13599,N_13403,N_13218);
nor U13600 (N_13600,N_13249,N_13444);
and U13601 (N_13601,N_13356,N_13374);
or U13602 (N_13602,N_13487,N_13201);
and U13603 (N_13603,N_13331,N_13271);
xor U13604 (N_13604,N_13447,N_13056);
and U13605 (N_13605,N_13393,N_13183);
or U13606 (N_13606,N_13098,N_13289);
nor U13607 (N_13607,N_13161,N_13287);
nor U13608 (N_13608,N_13299,N_13053);
nand U13609 (N_13609,N_13071,N_13050);
xnor U13610 (N_13610,N_13269,N_13346);
nor U13611 (N_13611,N_13076,N_13459);
or U13612 (N_13612,N_13339,N_13202);
or U13613 (N_13613,N_13332,N_13125);
nand U13614 (N_13614,N_13337,N_13425);
and U13615 (N_13615,N_13021,N_13101);
nor U13616 (N_13616,N_13298,N_13349);
nor U13617 (N_13617,N_13315,N_13175);
and U13618 (N_13618,N_13233,N_13372);
nor U13619 (N_13619,N_13180,N_13388);
nand U13620 (N_13620,N_13328,N_13347);
xor U13621 (N_13621,N_13100,N_13041);
or U13622 (N_13622,N_13394,N_13320);
xnor U13623 (N_13623,N_13214,N_13260);
nor U13624 (N_13624,N_13361,N_13031);
nand U13625 (N_13625,N_13463,N_13083);
nor U13626 (N_13626,N_13171,N_13468);
and U13627 (N_13627,N_13371,N_13057);
or U13628 (N_13628,N_13220,N_13032);
and U13629 (N_13629,N_13102,N_13205);
xnor U13630 (N_13630,N_13310,N_13103);
and U13631 (N_13631,N_13382,N_13044);
or U13632 (N_13632,N_13375,N_13030);
nor U13633 (N_13633,N_13143,N_13059);
xor U13634 (N_13634,N_13478,N_13043);
nor U13635 (N_13635,N_13185,N_13406);
and U13636 (N_13636,N_13093,N_13163);
xor U13637 (N_13637,N_13342,N_13496);
nor U13638 (N_13638,N_13285,N_13006);
nand U13639 (N_13639,N_13402,N_13303);
nand U13640 (N_13640,N_13493,N_13469);
xnor U13641 (N_13641,N_13248,N_13173);
nor U13642 (N_13642,N_13313,N_13087);
xnor U13643 (N_13643,N_13065,N_13013);
nand U13644 (N_13644,N_13238,N_13066);
xnor U13645 (N_13645,N_13191,N_13082);
nor U13646 (N_13646,N_13097,N_13479);
xor U13647 (N_13647,N_13294,N_13446);
nand U13648 (N_13648,N_13167,N_13413);
or U13649 (N_13649,N_13401,N_13212);
nor U13650 (N_13650,N_13025,N_13387);
nand U13651 (N_13651,N_13116,N_13113);
or U13652 (N_13652,N_13002,N_13156);
xnor U13653 (N_13653,N_13437,N_13122);
nand U13654 (N_13654,N_13074,N_13386);
and U13655 (N_13655,N_13352,N_13376);
nor U13656 (N_13656,N_13477,N_13009);
nor U13657 (N_13657,N_13344,N_13430);
nor U13658 (N_13658,N_13105,N_13365);
nand U13659 (N_13659,N_13068,N_13455);
nand U13660 (N_13660,N_13457,N_13197);
or U13661 (N_13661,N_13450,N_13262);
xor U13662 (N_13662,N_13494,N_13230);
nand U13663 (N_13663,N_13136,N_13011);
nor U13664 (N_13664,N_13018,N_13014);
nor U13665 (N_13665,N_13290,N_13033);
xnor U13666 (N_13666,N_13343,N_13499);
nor U13667 (N_13667,N_13358,N_13094);
xnor U13668 (N_13668,N_13368,N_13194);
xnor U13669 (N_13669,N_13330,N_13485);
or U13670 (N_13670,N_13231,N_13435);
nor U13671 (N_13671,N_13085,N_13144);
nor U13672 (N_13672,N_13400,N_13458);
xnor U13673 (N_13673,N_13381,N_13012);
nand U13674 (N_13674,N_13008,N_13326);
or U13675 (N_13675,N_13016,N_13005);
nand U13676 (N_13676,N_13222,N_13275);
nand U13677 (N_13677,N_13495,N_13219);
nor U13678 (N_13678,N_13363,N_13426);
xor U13679 (N_13679,N_13217,N_13084);
nand U13680 (N_13680,N_13118,N_13146);
and U13681 (N_13681,N_13139,N_13107);
or U13682 (N_13682,N_13411,N_13193);
nor U13683 (N_13683,N_13273,N_13325);
xnor U13684 (N_13684,N_13415,N_13309);
nand U13685 (N_13685,N_13224,N_13095);
nand U13686 (N_13686,N_13120,N_13150);
or U13687 (N_13687,N_13385,N_13266);
nor U13688 (N_13688,N_13465,N_13364);
xor U13689 (N_13689,N_13106,N_13259);
or U13690 (N_13690,N_13137,N_13203);
nor U13691 (N_13691,N_13357,N_13235);
and U13692 (N_13692,N_13416,N_13078);
nand U13693 (N_13693,N_13039,N_13228);
and U13694 (N_13694,N_13278,N_13474);
and U13695 (N_13695,N_13452,N_13404);
or U13696 (N_13696,N_13409,N_13272);
nand U13697 (N_13697,N_13131,N_13427);
or U13698 (N_13698,N_13355,N_13023);
nand U13699 (N_13699,N_13189,N_13225);
nor U13700 (N_13700,N_13239,N_13243);
and U13701 (N_13701,N_13334,N_13140);
and U13702 (N_13702,N_13195,N_13015);
and U13703 (N_13703,N_13288,N_13329);
xnor U13704 (N_13704,N_13379,N_13359);
nand U13705 (N_13705,N_13423,N_13431);
xor U13706 (N_13706,N_13208,N_13291);
nor U13707 (N_13707,N_13391,N_13077);
nand U13708 (N_13708,N_13466,N_13267);
and U13709 (N_13709,N_13434,N_13040);
or U13710 (N_13710,N_13242,N_13398);
and U13711 (N_13711,N_13317,N_13215);
nor U13712 (N_13712,N_13007,N_13099);
or U13713 (N_13713,N_13443,N_13000);
nor U13714 (N_13714,N_13148,N_13488);
or U13715 (N_13715,N_13476,N_13110);
nand U13716 (N_13716,N_13179,N_13241);
and U13717 (N_13717,N_13092,N_13345);
nand U13718 (N_13718,N_13453,N_13036);
nor U13719 (N_13719,N_13353,N_13395);
and U13720 (N_13720,N_13421,N_13300);
nor U13721 (N_13721,N_13301,N_13312);
or U13722 (N_13722,N_13277,N_13461);
and U13723 (N_13723,N_13414,N_13190);
nor U13724 (N_13724,N_13206,N_13472);
nor U13725 (N_13725,N_13306,N_13062);
and U13726 (N_13726,N_13130,N_13024);
xor U13727 (N_13727,N_13378,N_13486);
or U13728 (N_13728,N_13462,N_13075);
and U13729 (N_13729,N_13104,N_13123);
nand U13730 (N_13730,N_13412,N_13199);
and U13731 (N_13731,N_13067,N_13042);
and U13732 (N_13732,N_13177,N_13060);
xor U13733 (N_13733,N_13445,N_13253);
nand U13734 (N_13734,N_13283,N_13252);
xnor U13735 (N_13735,N_13396,N_13350);
and U13736 (N_13736,N_13438,N_13117);
or U13737 (N_13737,N_13470,N_13001);
nor U13738 (N_13738,N_13340,N_13168);
xnor U13739 (N_13739,N_13047,N_13429);
nand U13740 (N_13740,N_13017,N_13109);
or U13741 (N_13741,N_13070,N_13338);
xor U13742 (N_13742,N_13086,N_13158);
and U13743 (N_13743,N_13227,N_13407);
and U13744 (N_13744,N_13460,N_13265);
or U13745 (N_13745,N_13157,N_13127);
nor U13746 (N_13746,N_13323,N_13251);
and U13747 (N_13747,N_13035,N_13419);
nor U13748 (N_13748,N_13026,N_13181);
nor U13749 (N_13749,N_13480,N_13276);
nand U13750 (N_13750,N_13114,N_13058);
or U13751 (N_13751,N_13073,N_13317);
xnor U13752 (N_13752,N_13226,N_13479);
or U13753 (N_13753,N_13182,N_13358);
nor U13754 (N_13754,N_13223,N_13070);
nand U13755 (N_13755,N_13195,N_13176);
or U13756 (N_13756,N_13204,N_13358);
and U13757 (N_13757,N_13249,N_13352);
xnor U13758 (N_13758,N_13353,N_13169);
and U13759 (N_13759,N_13282,N_13368);
and U13760 (N_13760,N_13213,N_13042);
xnor U13761 (N_13761,N_13025,N_13177);
xnor U13762 (N_13762,N_13427,N_13241);
or U13763 (N_13763,N_13270,N_13336);
and U13764 (N_13764,N_13176,N_13179);
nand U13765 (N_13765,N_13498,N_13247);
and U13766 (N_13766,N_13150,N_13235);
or U13767 (N_13767,N_13147,N_13346);
xor U13768 (N_13768,N_13438,N_13132);
nor U13769 (N_13769,N_13450,N_13018);
nor U13770 (N_13770,N_13324,N_13369);
and U13771 (N_13771,N_13088,N_13165);
and U13772 (N_13772,N_13306,N_13273);
and U13773 (N_13773,N_13363,N_13104);
and U13774 (N_13774,N_13012,N_13004);
or U13775 (N_13775,N_13396,N_13082);
or U13776 (N_13776,N_13108,N_13470);
and U13777 (N_13777,N_13260,N_13204);
or U13778 (N_13778,N_13089,N_13164);
or U13779 (N_13779,N_13067,N_13158);
and U13780 (N_13780,N_13413,N_13386);
or U13781 (N_13781,N_13356,N_13025);
and U13782 (N_13782,N_13239,N_13420);
xor U13783 (N_13783,N_13447,N_13237);
nor U13784 (N_13784,N_13425,N_13346);
xor U13785 (N_13785,N_13254,N_13204);
nor U13786 (N_13786,N_13038,N_13263);
nand U13787 (N_13787,N_13258,N_13219);
or U13788 (N_13788,N_13190,N_13272);
and U13789 (N_13789,N_13249,N_13309);
or U13790 (N_13790,N_13234,N_13428);
nor U13791 (N_13791,N_13097,N_13083);
or U13792 (N_13792,N_13076,N_13336);
or U13793 (N_13793,N_13205,N_13448);
or U13794 (N_13794,N_13321,N_13055);
and U13795 (N_13795,N_13333,N_13377);
nand U13796 (N_13796,N_13494,N_13027);
nand U13797 (N_13797,N_13398,N_13147);
xnor U13798 (N_13798,N_13166,N_13427);
xor U13799 (N_13799,N_13012,N_13145);
nor U13800 (N_13800,N_13185,N_13262);
and U13801 (N_13801,N_13224,N_13090);
nand U13802 (N_13802,N_13413,N_13455);
nor U13803 (N_13803,N_13336,N_13265);
or U13804 (N_13804,N_13332,N_13133);
nor U13805 (N_13805,N_13017,N_13072);
or U13806 (N_13806,N_13036,N_13439);
and U13807 (N_13807,N_13444,N_13201);
xnor U13808 (N_13808,N_13068,N_13222);
and U13809 (N_13809,N_13238,N_13019);
or U13810 (N_13810,N_13486,N_13437);
xor U13811 (N_13811,N_13483,N_13175);
or U13812 (N_13812,N_13368,N_13134);
nand U13813 (N_13813,N_13222,N_13442);
and U13814 (N_13814,N_13386,N_13382);
and U13815 (N_13815,N_13210,N_13093);
nand U13816 (N_13816,N_13256,N_13095);
or U13817 (N_13817,N_13234,N_13005);
or U13818 (N_13818,N_13353,N_13272);
or U13819 (N_13819,N_13276,N_13454);
nor U13820 (N_13820,N_13130,N_13117);
nand U13821 (N_13821,N_13143,N_13314);
or U13822 (N_13822,N_13206,N_13123);
and U13823 (N_13823,N_13490,N_13103);
or U13824 (N_13824,N_13320,N_13400);
or U13825 (N_13825,N_13130,N_13009);
nand U13826 (N_13826,N_13230,N_13048);
xor U13827 (N_13827,N_13035,N_13179);
xnor U13828 (N_13828,N_13102,N_13349);
and U13829 (N_13829,N_13020,N_13300);
and U13830 (N_13830,N_13101,N_13240);
nand U13831 (N_13831,N_13364,N_13090);
nand U13832 (N_13832,N_13145,N_13283);
nand U13833 (N_13833,N_13344,N_13153);
nor U13834 (N_13834,N_13204,N_13100);
or U13835 (N_13835,N_13332,N_13271);
nand U13836 (N_13836,N_13102,N_13061);
nor U13837 (N_13837,N_13187,N_13494);
xor U13838 (N_13838,N_13307,N_13107);
nor U13839 (N_13839,N_13109,N_13297);
nor U13840 (N_13840,N_13004,N_13219);
xor U13841 (N_13841,N_13264,N_13014);
nor U13842 (N_13842,N_13270,N_13314);
nand U13843 (N_13843,N_13178,N_13236);
xnor U13844 (N_13844,N_13228,N_13056);
or U13845 (N_13845,N_13409,N_13170);
xor U13846 (N_13846,N_13102,N_13115);
or U13847 (N_13847,N_13284,N_13483);
nand U13848 (N_13848,N_13145,N_13019);
nor U13849 (N_13849,N_13442,N_13405);
nand U13850 (N_13850,N_13039,N_13279);
or U13851 (N_13851,N_13389,N_13204);
or U13852 (N_13852,N_13185,N_13428);
or U13853 (N_13853,N_13271,N_13195);
and U13854 (N_13854,N_13174,N_13374);
nor U13855 (N_13855,N_13319,N_13092);
nand U13856 (N_13856,N_13241,N_13100);
nor U13857 (N_13857,N_13195,N_13105);
nand U13858 (N_13858,N_13330,N_13024);
or U13859 (N_13859,N_13103,N_13455);
and U13860 (N_13860,N_13052,N_13004);
or U13861 (N_13861,N_13047,N_13393);
nor U13862 (N_13862,N_13495,N_13196);
nand U13863 (N_13863,N_13135,N_13063);
or U13864 (N_13864,N_13467,N_13390);
nand U13865 (N_13865,N_13488,N_13017);
nor U13866 (N_13866,N_13249,N_13203);
nor U13867 (N_13867,N_13238,N_13379);
or U13868 (N_13868,N_13459,N_13064);
nand U13869 (N_13869,N_13338,N_13025);
or U13870 (N_13870,N_13231,N_13425);
xor U13871 (N_13871,N_13326,N_13145);
nand U13872 (N_13872,N_13284,N_13323);
or U13873 (N_13873,N_13201,N_13158);
and U13874 (N_13874,N_13459,N_13139);
nand U13875 (N_13875,N_13322,N_13018);
and U13876 (N_13876,N_13226,N_13085);
or U13877 (N_13877,N_13270,N_13408);
nand U13878 (N_13878,N_13204,N_13145);
nor U13879 (N_13879,N_13123,N_13225);
xnor U13880 (N_13880,N_13346,N_13282);
xnor U13881 (N_13881,N_13314,N_13280);
nor U13882 (N_13882,N_13256,N_13302);
or U13883 (N_13883,N_13293,N_13163);
and U13884 (N_13884,N_13080,N_13070);
nor U13885 (N_13885,N_13253,N_13364);
nand U13886 (N_13886,N_13429,N_13373);
or U13887 (N_13887,N_13286,N_13384);
xor U13888 (N_13888,N_13491,N_13138);
or U13889 (N_13889,N_13014,N_13007);
nand U13890 (N_13890,N_13061,N_13341);
nor U13891 (N_13891,N_13358,N_13489);
or U13892 (N_13892,N_13128,N_13037);
xnor U13893 (N_13893,N_13422,N_13186);
or U13894 (N_13894,N_13166,N_13368);
nand U13895 (N_13895,N_13203,N_13413);
xnor U13896 (N_13896,N_13291,N_13177);
xor U13897 (N_13897,N_13485,N_13324);
or U13898 (N_13898,N_13358,N_13455);
nor U13899 (N_13899,N_13070,N_13078);
nand U13900 (N_13900,N_13240,N_13373);
nand U13901 (N_13901,N_13329,N_13471);
nor U13902 (N_13902,N_13400,N_13340);
and U13903 (N_13903,N_13122,N_13469);
or U13904 (N_13904,N_13441,N_13438);
and U13905 (N_13905,N_13074,N_13225);
xnor U13906 (N_13906,N_13102,N_13170);
nor U13907 (N_13907,N_13254,N_13497);
nor U13908 (N_13908,N_13030,N_13132);
nor U13909 (N_13909,N_13493,N_13017);
xnor U13910 (N_13910,N_13478,N_13101);
nand U13911 (N_13911,N_13242,N_13151);
xnor U13912 (N_13912,N_13017,N_13198);
nor U13913 (N_13913,N_13251,N_13386);
xnor U13914 (N_13914,N_13127,N_13336);
and U13915 (N_13915,N_13077,N_13127);
xor U13916 (N_13916,N_13224,N_13431);
xnor U13917 (N_13917,N_13006,N_13346);
xnor U13918 (N_13918,N_13287,N_13440);
nand U13919 (N_13919,N_13414,N_13485);
xor U13920 (N_13920,N_13185,N_13414);
xor U13921 (N_13921,N_13014,N_13416);
and U13922 (N_13922,N_13230,N_13378);
nand U13923 (N_13923,N_13063,N_13345);
nand U13924 (N_13924,N_13104,N_13276);
nor U13925 (N_13925,N_13155,N_13065);
nor U13926 (N_13926,N_13124,N_13237);
and U13927 (N_13927,N_13300,N_13057);
and U13928 (N_13928,N_13487,N_13095);
and U13929 (N_13929,N_13054,N_13155);
xnor U13930 (N_13930,N_13290,N_13191);
and U13931 (N_13931,N_13161,N_13045);
nand U13932 (N_13932,N_13446,N_13188);
xnor U13933 (N_13933,N_13004,N_13384);
nor U13934 (N_13934,N_13000,N_13024);
nor U13935 (N_13935,N_13098,N_13432);
xor U13936 (N_13936,N_13131,N_13006);
xnor U13937 (N_13937,N_13080,N_13472);
or U13938 (N_13938,N_13044,N_13260);
nor U13939 (N_13939,N_13271,N_13438);
or U13940 (N_13940,N_13478,N_13163);
or U13941 (N_13941,N_13210,N_13223);
xnor U13942 (N_13942,N_13363,N_13177);
nor U13943 (N_13943,N_13469,N_13456);
or U13944 (N_13944,N_13068,N_13376);
xnor U13945 (N_13945,N_13401,N_13402);
nand U13946 (N_13946,N_13346,N_13405);
or U13947 (N_13947,N_13425,N_13325);
and U13948 (N_13948,N_13260,N_13367);
xor U13949 (N_13949,N_13292,N_13275);
xnor U13950 (N_13950,N_13174,N_13080);
xor U13951 (N_13951,N_13013,N_13158);
xnor U13952 (N_13952,N_13326,N_13487);
nand U13953 (N_13953,N_13217,N_13410);
nor U13954 (N_13954,N_13465,N_13088);
nor U13955 (N_13955,N_13160,N_13013);
nand U13956 (N_13956,N_13209,N_13175);
nor U13957 (N_13957,N_13233,N_13137);
or U13958 (N_13958,N_13207,N_13469);
and U13959 (N_13959,N_13392,N_13154);
xnor U13960 (N_13960,N_13333,N_13300);
nor U13961 (N_13961,N_13446,N_13386);
nand U13962 (N_13962,N_13002,N_13246);
xnor U13963 (N_13963,N_13272,N_13253);
and U13964 (N_13964,N_13458,N_13284);
or U13965 (N_13965,N_13049,N_13133);
nand U13966 (N_13966,N_13494,N_13379);
nand U13967 (N_13967,N_13147,N_13353);
and U13968 (N_13968,N_13473,N_13289);
xnor U13969 (N_13969,N_13473,N_13385);
nor U13970 (N_13970,N_13403,N_13111);
and U13971 (N_13971,N_13017,N_13046);
and U13972 (N_13972,N_13196,N_13431);
and U13973 (N_13973,N_13322,N_13029);
xnor U13974 (N_13974,N_13230,N_13045);
nand U13975 (N_13975,N_13124,N_13026);
xnor U13976 (N_13976,N_13235,N_13281);
nand U13977 (N_13977,N_13051,N_13356);
nor U13978 (N_13978,N_13147,N_13161);
and U13979 (N_13979,N_13365,N_13238);
nand U13980 (N_13980,N_13013,N_13427);
and U13981 (N_13981,N_13193,N_13155);
or U13982 (N_13982,N_13352,N_13448);
nor U13983 (N_13983,N_13098,N_13451);
xnor U13984 (N_13984,N_13336,N_13251);
nand U13985 (N_13985,N_13042,N_13484);
nor U13986 (N_13986,N_13111,N_13485);
nor U13987 (N_13987,N_13004,N_13022);
nand U13988 (N_13988,N_13480,N_13155);
and U13989 (N_13989,N_13434,N_13013);
nand U13990 (N_13990,N_13191,N_13048);
nor U13991 (N_13991,N_13127,N_13098);
xnor U13992 (N_13992,N_13452,N_13256);
xor U13993 (N_13993,N_13480,N_13304);
xor U13994 (N_13994,N_13070,N_13184);
or U13995 (N_13995,N_13304,N_13162);
or U13996 (N_13996,N_13255,N_13229);
nand U13997 (N_13997,N_13310,N_13392);
and U13998 (N_13998,N_13176,N_13137);
or U13999 (N_13999,N_13018,N_13068);
or U14000 (N_14000,N_13824,N_13888);
or U14001 (N_14001,N_13954,N_13801);
or U14002 (N_14002,N_13791,N_13556);
or U14003 (N_14003,N_13544,N_13522);
xnor U14004 (N_14004,N_13618,N_13950);
nand U14005 (N_14005,N_13805,N_13973);
nor U14006 (N_14006,N_13899,N_13861);
nand U14007 (N_14007,N_13755,N_13662);
nand U14008 (N_14008,N_13847,N_13587);
nand U14009 (N_14009,N_13603,N_13518);
or U14010 (N_14010,N_13820,N_13822);
nor U14011 (N_14011,N_13844,N_13508);
xor U14012 (N_14012,N_13952,N_13978);
or U14013 (N_14013,N_13507,N_13584);
nor U14014 (N_14014,N_13945,N_13562);
and U14015 (N_14015,N_13878,N_13578);
and U14016 (N_14016,N_13609,N_13560);
or U14017 (N_14017,N_13632,N_13750);
nand U14018 (N_14018,N_13541,N_13761);
and U14019 (N_14019,N_13958,N_13616);
and U14020 (N_14020,N_13612,N_13961);
xnor U14021 (N_14021,N_13930,N_13887);
nor U14022 (N_14022,N_13933,N_13558);
or U14023 (N_14023,N_13826,N_13962);
and U14024 (N_14024,N_13811,N_13645);
and U14025 (N_14025,N_13848,N_13795);
or U14026 (N_14026,N_13994,N_13751);
and U14027 (N_14027,N_13714,N_13864);
xor U14028 (N_14028,N_13579,N_13604);
or U14029 (N_14029,N_13981,N_13817);
and U14030 (N_14030,N_13797,N_13884);
or U14031 (N_14031,N_13759,N_13707);
or U14032 (N_14032,N_13690,N_13920);
nor U14033 (N_14033,N_13652,N_13676);
and U14034 (N_14034,N_13535,N_13924);
nor U14035 (N_14035,N_13730,N_13925);
xnor U14036 (N_14036,N_13803,N_13914);
nand U14037 (N_14037,N_13784,N_13968);
xor U14038 (N_14038,N_13741,N_13533);
nor U14039 (N_14039,N_13553,N_13681);
nand U14040 (N_14040,N_13636,N_13992);
and U14041 (N_14041,N_13580,N_13849);
and U14042 (N_14042,N_13619,N_13561);
xor U14043 (N_14043,N_13571,N_13905);
nor U14044 (N_14044,N_13971,N_13724);
and U14045 (N_14045,N_13781,N_13531);
and U14046 (N_14046,N_13511,N_13519);
and U14047 (N_14047,N_13770,N_13926);
nand U14048 (N_14048,N_13787,N_13697);
nor U14049 (N_14049,N_13705,N_13794);
xor U14050 (N_14050,N_13935,N_13996);
nor U14051 (N_14051,N_13521,N_13732);
or U14052 (N_14052,N_13721,N_13540);
nor U14053 (N_14053,N_13881,N_13856);
or U14054 (N_14054,N_13734,N_13737);
or U14055 (N_14055,N_13532,N_13793);
xnor U14056 (N_14056,N_13753,N_13785);
and U14057 (N_14057,N_13680,N_13557);
nand U14058 (N_14058,N_13744,N_13995);
xnor U14059 (N_14059,N_13923,N_13859);
xnor U14060 (N_14060,N_13570,N_13912);
nand U14061 (N_14061,N_13775,N_13902);
or U14062 (N_14062,N_13964,N_13872);
nor U14063 (N_14063,N_13976,N_13733);
nand U14064 (N_14064,N_13726,N_13840);
nand U14065 (N_14065,N_13898,N_13665);
nor U14066 (N_14066,N_13895,N_13700);
nand U14067 (N_14067,N_13728,N_13673);
nor U14068 (N_14068,N_13740,N_13896);
nand U14069 (N_14069,N_13611,N_13804);
xor U14070 (N_14070,N_13808,N_13934);
xor U14071 (N_14071,N_13551,N_13957);
nand U14072 (N_14072,N_13543,N_13500);
xnor U14073 (N_14073,N_13910,N_13642);
xnor U14074 (N_14074,N_13670,N_13894);
or U14075 (N_14075,N_13688,N_13581);
and U14076 (N_14076,N_13524,N_13622);
nand U14077 (N_14077,N_13717,N_13893);
or U14078 (N_14078,N_13672,N_13788);
xnor U14079 (N_14079,N_13845,N_13526);
nor U14080 (N_14080,N_13701,N_13590);
xnor U14081 (N_14081,N_13615,N_13679);
or U14082 (N_14082,N_13509,N_13545);
xnor U14083 (N_14083,N_13602,N_13736);
nor U14084 (N_14084,N_13860,N_13566);
and U14085 (N_14085,N_13720,N_13746);
xor U14086 (N_14086,N_13598,N_13549);
and U14087 (N_14087,N_13815,N_13706);
nor U14088 (N_14088,N_13660,N_13823);
nor U14089 (N_14089,N_13646,N_13927);
nor U14090 (N_14090,N_13656,N_13539);
nor U14091 (N_14091,N_13982,N_13907);
and U14092 (N_14092,N_13627,N_13678);
and U14093 (N_14093,N_13985,N_13554);
or U14094 (N_14094,N_13932,N_13640);
or U14095 (N_14095,N_13832,N_13960);
and U14096 (N_14096,N_13542,N_13999);
nor U14097 (N_14097,N_13715,N_13747);
nand U14098 (N_14098,N_13668,N_13969);
xor U14099 (N_14099,N_13951,N_13825);
nor U14100 (N_14100,N_13589,N_13838);
nor U14101 (N_14101,N_13569,N_13601);
or U14102 (N_14102,N_13525,N_13798);
or U14103 (N_14103,N_13876,N_13591);
nand U14104 (N_14104,N_13889,N_13863);
and U14105 (N_14105,N_13727,N_13900);
or U14106 (N_14106,N_13503,N_13685);
nor U14107 (N_14107,N_13911,N_13937);
and U14108 (N_14108,N_13729,N_13537);
xnor U14109 (N_14109,N_13768,N_13648);
or U14110 (N_14110,N_13624,N_13550);
xnor U14111 (N_14111,N_13565,N_13644);
nand U14112 (N_14112,N_13936,N_13802);
xnor U14113 (N_14113,N_13588,N_13842);
or U14114 (N_14114,N_13599,N_13833);
and U14115 (N_14115,N_13818,N_13754);
xor U14116 (N_14116,N_13649,N_13693);
nand U14117 (N_14117,N_13830,N_13710);
and U14118 (N_14118,N_13821,N_13638);
xor U14119 (N_14119,N_13712,N_13988);
nor U14120 (N_14120,N_13564,N_13723);
nand U14121 (N_14121,N_13772,N_13790);
nand U14122 (N_14122,N_13866,N_13819);
xnor U14123 (N_14123,N_13684,N_13916);
or U14124 (N_14124,N_13666,N_13983);
xor U14125 (N_14125,N_13800,N_13689);
and U14126 (N_14126,N_13948,N_13719);
or U14127 (N_14127,N_13843,N_13943);
xor U14128 (N_14128,N_13594,N_13661);
nor U14129 (N_14129,N_13758,N_13659);
and U14130 (N_14130,N_13738,N_13850);
nand U14131 (N_14131,N_13628,N_13979);
nor U14132 (N_14132,N_13757,N_13870);
nor U14133 (N_14133,N_13629,N_13510);
nand U14134 (N_14134,N_13947,N_13959);
nand U14135 (N_14135,N_13711,N_13641);
and U14136 (N_14136,N_13585,N_13883);
nand U14137 (N_14137,N_13890,N_13546);
and U14138 (N_14138,N_13617,N_13575);
and U14139 (N_14139,N_13505,N_13931);
or U14140 (N_14140,N_13696,N_13839);
xnor U14141 (N_14141,N_13657,N_13941);
or U14142 (N_14142,N_13975,N_13913);
or U14143 (N_14143,N_13812,N_13658);
nor U14144 (N_14144,N_13852,N_13699);
or U14145 (N_14145,N_13674,N_13796);
or U14146 (N_14146,N_13997,N_13906);
and U14147 (N_14147,N_13865,N_13516);
nand U14148 (N_14148,N_13778,N_13692);
or U14149 (N_14149,N_13671,N_13596);
and U14150 (N_14150,N_13529,N_13536);
and U14151 (N_14151,N_13963,N_13742);
nand U14152 (N_14152,N_13610,N_13972);
nor U14153 (N_14153,N_13606,N_13908);
or U14154 (N_14154,N_13626,N_13669);
nor U14155 (N_14155,N_13527,N_13667);
xor U14156 (N_14156,N_13762,N_13663);
xor U14157 (N_14157,N_13873,N_13769);
and U14158 (N_14158,N_13514,N_13831);
nand U14159 (N_14159,N_13583,N_13538);
nor U14160 (N_14160,N_13909,N_13783);
nand U14161 (N_14161,N_13764,N_13828);
and U14162 (N_14162,N_13780,N_13980);
or U14163 (N_14163,N_13816,N_13592);
and U14164 (N_14164,N_13530,N_13875);
or U14165 (N_14165,N_13903,N_13846);
nor U14166 (N_14166,N_13809,N_13837);
or U14167 (N_14167,N_13749,N_13882);
and U14168 (N_14168,N_13760,N_13573);
or U14169 (N_14169,N_13630,N_13515);
or U14170 (N_14170,N_13970,N_13574);
or U14171 (N_14171,N_13917,N_13506);
nand U14172 (N_14172,N_13955,N_13694);
xnor U14173 (N_14173,N_13854,N_13748);
xor U14174 (N_14174,N_13608,N_13834);
or U14175 (N_14175,N_13886,N_13857);
nand U14176 (N_14176,N_13600,N_13965);
nand U14177 (N_14177,N_13998,N_13702);
xnor U14178 (N_14178,N_13739,N_13735);
and U14179 (N_14179,N_13568,N_13880);
or U14180 (N_14180,N_13634,N_13869);
or U14181 (N_14181,N_13792,N_13716);
nor U14182 (N_14182,N_13967,N_13523);
and U14183 (N_14183,N_13695,N_13841);
nor U14184 (N_14184,N_13835,N_13623);
nor U14185 (N_14185,N_13940,N_13752);
nand U14186 (N_14186,N_13938,N_13691);
xnor U14187 (N_14187,N_13766,N_13614);
or U14188 (N_14188,N_13779,N_13977);
nor U14189 (N_14189,N_13891,N_13984);
or U14190 (N_14190,N_13704,N_13974);
or U14191 (N_14191,N_13946,N_13725);
xnor U14192 (N_14192,N_13597,N_13577);
nand U14193 (N_14193,N_13765,N_13555);
or U14194 (N_14194,N_13966,N_13874);
xor U14195 (N_14195,N_13904,N_13501);
xor U14196 (N_14196,N_13677,N_13944);
xor U14197 (N_14197,N_13547,N_13918);
nor U14198 (N_14198,N_13621,N_13836);
nand U14199 (N_14199,N_13789,N_13885);
xor U14200 (N_14200,N_13512,N_13949);
nor U14201 (N_14201,N_13607,N_13855);
nor U14202 (N_14202,N_13922,N_13892);
nand U14203 (N_14203,N_13586,N_13813);
xor U14204 (N_14204,N_13552,N_13771);
xnor U14205 (N_14205,N_13991,N_13786);
nand U14206 (N_14206,N_13548,N_13582);
xor U14207 (N_14207,N_13743,N_13807);
or U14208 (N_14208,N_13713,N_13810);
nand U14209 (N_14209,N_13605,N_13633);
nor U14210 (N_14210,N_13877,N_13921);
nor U14211 (N_14211,N_13683,N_13853);
xor U14212 (N_14212,N_13576,N_13653);
nand U14213 (N_14213,N_13867,N_13986);
xnor U14214 (N_14214,N_13534,N_13520);
nand U14215 (N_14215,N_13647,N_13897);
nand U14216 (N_14216,N_13502,N_13643);
xnor U14217 (N_14217,N_13942,N_13682);
nand U14218 (N_14218,N_13595,N_13928);
nand U14219 (N_14219,N_13654,N_13953);
nor U14220 (N_14220,N_13698,N_13718);
or U14221 (N_14221,N_13709,N_13901);
nor U14222 (N_14222,N_13862,N_13773);
or U14223 (N_14223,N_13513,N_13620);
and U14224 (N_14224,N_13851,N_13708);
nor U14225 (N_14225,N_13929,N_13650);
and U14226 (N_14226,N_13799,N_13777);
xnor U14227 (N_14227,N_13528,N_13767);
nor U14228 (N_14228,N_13655,N_13919);
nor U14229 (N_14229,N_13703,N_13675);
and U14230 (N_14230,N_13858,N_13625);
and U14231 (N_14231,N_13990,N_13993);
and U14232 (N_14232,N_13756,N_13806);
and U14233 (N_14233,N_13829,N_13687);
xor U14234 (N_14234,N_13763,N_13868);
and U14235 (N_14235,N_13827,N_13731);
nor U14236 (N_14236,N_13989,N_13776);
nor U14237 (N_14237,N_13987,N_13517);
xnor U14238 (N_14238,N_13915,N_13686);
xnor U14239 (N_14239,N_13651,N_13639);
or U14240 (N_14240,N_13956,N_13559);
and U14241 (N_14241,N_13567,N_13814);
and U14242 (N_14242,N_13572,N_13637);
nand U14243 (N_14243,N_13613,N_13939);
xor U14244 (N_14244,N_13631,N_13879);
or U14245 (N_14245,N_13635,N_13782);
and U14246 (N_14246,N_13593,N_13722);
or U14247 (N_14247,N_13563,N_13664);
nor U14248 (N_14248,N_13504,N_13745);
xor U14249 (N_14249,N_13871,N_13774);
nor U14250 (N_14250,N_13626,N_13539);
nand U14251 (N_14251,N_13990,N_13526);
nor U14252 (N_14252,N_13675,N_13727);
and U14253 (N_14253,N_13607,N_13742);
or U14254 (N_14254,N_13862,N_13623);
xor U14255 (N_14255,N_13948,N_13918);
nor U14256 (N_14256,N_13916,N_13806);
or U14257 (N_14257,N_13656,N_13845);
nand U14258 (N_14258,N_13638,N_13786);
xor U14259 (N_14259,N_13680,N_13729);
nand U14260 (N_14260,N_13610,N_13622);
or U14261 (N_14261,N_13944,N_13568);
or U14262 (N_14262,N_13586,N_13989);
and U14263 (N_14263,N_13643,N_13875);
nand U14264 (N_14264,N_13781,N_13980);
xnor U14265 (N_14265,N_13734,N_13749);
and U14266 (N_14266,N_13796,N_13910);
nand U14267 (N_14267,N_13534,N_13697);
or U14268 (N_14268,N_13772,N_13819);
nand U14269 (N_14269,N_13633,N_13588);
xor U14270 (N_14270,N_13637,N_13924);
and U14271 (N_14271,N_13768,N_13569);
and U14272 (N_14272,N_13706,N_13856);
xnor U14273 (N_14273,N_13590,N_13565);
xnor U14274 (N_14274,N_13573,N_13870);
or U14275 (N_14275,N_13723,N_13618);
and U14276 (N_14276,N_13780,N_13846);
or U14277 (N_14277,N_13869,N_13857);
xor U14278 (N_14278,N_13883,N_13961);
nor U14279 (N_14279,N_13864,N_13821);
nand U14280 (N_14280,N_13779,N_13789);
and U14281 (N_14281,N_13506,N_13796);
nand U14282 (N_14282,N_13895,N_13704);
nand U14283 (N_14283,N_13832,N_13805);
and U14284 (N_14284,N_13545,N_13843);
xor U14285 (N_14285,N_13874,N_13834);
nand U14286 (N_14286,N_13648,N_13995);
xnor U14287 (N_14287,N_13908,N_13659);
xor U14288 (N_14288,N_13770,N_13854);
nor U14289 (N_14289,N_13569,N_13714);
and U14290 (N_14290,N_13686,N_13537);
xor U14291 (N_14291,N_13592,N_13547);
xnor U14292 (N_14292,N_13550,N_13732);
xnor U14293 (N_14293,N_13996,N_13713);
xor U14294 (N_14294,N_13628,N_13665);
nand U14295 (N_14295,N_13758,N_13982);
and U14296 (N_14296,N_13602,N_13635);
nand U14297 (N_14297,N_13598,N_13624);
nor U14298 (N_14298,N_13767,N_13682);
or U14299 (N_14299,N_13988,N_13622);
or U14300 (N_14300,N_13534,N_13730);
nand U14301 (N_14301,N_13929,N_13978);
nor U14302 (N_14302,N_13938,N_13588);
and U14303 (N_14303,N_13637,N_13804);
nor U14304 (N_14304,N_13902,N_13549);
and U14305 (N_14305,N_13680,N_13739);
nor U14306 (N_14306,N_13940,N_13675);
xor U14307 (N_14307,N_13644,N_13723);
and U14308 (N_14308,N_13938,N_13786);
nor U14309 (N_14309,N_13996,N_13798);
nand U14310 (N_14310,N_13877,N_13515);
and U14311 (N_14311,N_13707,N_13613);
or U14312 (N_14312,N_13519,N_13542);
or U14313 (N_14313,N_13850,N_13831);
xnor U14314 (N_14314,N_13723,N_13812);
nor U14315 (N_14315,N_13583,N_13998);
nor U14316 (N_14316,N_13722,N_13579);
or U14317 (N_14317,N_13994,N_13704);
nor U14318 (N_14318,N_13807,N_13818);
xnor U14319 (N_14319,N_13743,N_13591);
or U14320 (N_14320,N_13919,N_13687);
nor U14321 (N_14321,N_13582,N_13552);
nor U14322 (N_14322,N_13571,N_13807);
nand U14323 (N_14323,N_13757,N_13621);
nand U14324 (N_14324,N_13875,N_13873);
xnor U14325 (N_14325,N_13916,N_13780);
and U14326 (N_14326,N_13540,N_13863);
or U14327 (N_14327,N_13830,N_13699);
xnor U14328 (N_14328,N_13993,N_13582);
nand U14329 (N_14329,N_13659,N_13627);
nor U14330 (N_14330,N_13528,N_13647);
xnor U14331 (N_14331,N_13962,N_13526);
nor U14332 (N_14332,N_13524,N_13974);
and U14333 (N_14333,N_13983,N_13831);
nor U14334 (N_14334,N_13963,N_13525);
nand U14335 (N_14335,N_13624,N_13536);
and U14336 (N_14336,N_13575,N_13879);
or U14337 (N_14337,N_13975,N_13607);
xnor U14338 (N_14338,N_13739,N_13785);
or U14339 (N_14339,N_13707,N_13767);
xor U14340 (N_14340,N_13524,N_13731);
or U14341 (N_14341,N_13514,N_13885);
nand U14342 (N_14342,N_13868,N_13543);
nor U14343 (N_14343,N_13588,N_13816);
nor U14344 (N_14344,N_13823,N_13581);
nand U14345 (N_14345,N_13920,N_13596);
and U14346 (N_14346,N_13630,N_13642);
nand U14347 (N_14347,N_13769,N_13770);
and U14348 (N_14348,N_13975,N_13947);
xor U14349 (N_14349,N_13951,N_13676);
and U14350 (N_14350,N_13619,N_13502);
xor U14351 (N_14351,N_13555,N_13894);
nor U14352 (N_14352,N_13982,N_13724);
and U14353 (N_14353,N_13842,N_13915);
nand U14354 (N_14354,N_13647,N_13918);
xor U14355 (N_14355,N_13657,N_13559);
xnor U14356 (N_14356,N_13769,N_13723);
and U14357 (N_14357,N_13530,N_13766);
and U14358 (N_14358,N_13853,N_13906);
nand U14359 (N_14359,N_13731,N_13939);
xnor U14360 (N_14360,N_13500,N_13514);
nand U14361 (N_14361,N_13643,N_13551);
and U14362 (N_14362,N_13708,N_13747);
xor U14363 (N_14363,N_13842,N_13809);
or U14364 (N_14364,N_13814,N_13859);
xor U14365 (N_14365,N_13989,N_13618);
xor U14366 (N_14366,N_13510,N_13819);
and U14367 (N_14367,N_13567,N_13738);
nor U14368 (N_14368,N_13735,N_13899);
and U14369 (N_14369,N_13546,N_13601);
nor U14370 (N_14370,N_13611,N_13551);
xor U14371 (N_14371,N_13558,N_13598);
nand U14372 (N_14372,N_13569,N_13935);
xor U14373 (N_14373,N_13873,N_13729);
or U14374 (N_14374,N_13850,N_13686);
nor U14375 (N_14375,N_13580,N_13893);
nand U14376 (N_14376,N_13980,N_13993);
or U14377 (N_14377,N_13994,N_13643);
nor U14378 (N_14378,N_13551,N_13783);
nor U14379 (N_14379,N_13757,N_13787);
xnor U14380 (N_14380,N_13500,N_13616);
or U14381 (N_14381,N_13700,N_13870);
nor U14382 (N_14382,N_13798,N_13569);
xnor U14383 (N_14383,N_13663,N_13777);
and U14384 (N_14384,N_13995,N_13515);
nand U14385 (N_14385,N_13808,N_13817);
nand U14386 (N_14386,N_13528,N_13582);
or U14387 (N_14387,N_13930,N_13556);
xnor U14388 (N_14388,N_13867,N_13939);
xnor U14389 (N_14389,N_13927,N_13658);
nor U14390 (N_14390,N_13981,N_13619);
xnor U14391 (N_14391,N_13837,N_13841);
and U14392 (N_14392,N_13844,N_13731);
or U14393 (N_14393,N_13590,N_13724);
and U14394 (N_14394,N_13950,N_13754);
nor U14395 (N_14395,N_13809,N_13974);
or U14396 (N_14396,N_13549,N_13914);
xnor U14397 (N_14397,N_13533,N_13519);
and U14398 (N_14398,N_13963,N_13807);
nor U14399 (N_14399,N_13921,N_13558);
and U14400 (N_14400,N_13992,N_13549);
xnor U14401 (N_14401,N_13791,N_13877);
xor U14402 (N_14402,N_13617,N_13918);
xor U14403 (N_14403,N_13987,N_13889);
nor U14404 (N_14404,N_13916,N_13874);
nor U14405 (N_14405,N_13843,N_13945);
nand U14406 (N_14406,N_13834,N_13517);
xor U14407 (N_14407,N_13853,N_13505);
or U14408 (N_14408,N_13503,N_13978);
nand U14409 (N_14409,N_13692,N_13923);
and U14410 (N_14410,N_13750,N_13829);
and U14411 (N_14411,N_13704,N_13680);
nor U14412 (N_14412,N_13943,N_13523);
nor U14413 (N_14413,N_13732,N_13739);
nand U14414 (N_14414,N_13729,N_13853);
nand U14415 (N_14415,N_13704,N_13885);
nor U14416 (N_14416,N_13980,N_13819);
nor U14417 (N_14417,N_13547,N_13848);
and U14418 (N_14418,N_13800,N_13975);
or U14419 (N_14419,N_13609,N_13886);
or U14420 (N_14420,N_13665,N_13965);
nand U14421 (N_14421,N_13549,N_13788);
xor U14422 (N_14422,N_13707,N_13862);
xor U14423 (N_14423,N_13993,N_13997);
nand U14424 (N_14424,N_13722,N_13581);
nand U14425 (N_14425,N_13746,N_13971);
or U14426 (N_14426,N_13773,N_13514);
and U14427 (N_14427,N_13832,N_13689);
nor U14428 (N_14428,N_13766,N_13710);
xor U14429 (N_14429,N_13501,N_13847);
and U14430 (N_14430,N_13501,N_13703);
nand U14431 (N_14431,N_13958,N_13577);
nand U14432 (N_14432,N_13725,N_13835);
or U14433 (N_14433,N_13965,N_13812);
nor U14434 (N_14434,N_13889,N_13526);
or U14435 (N_14435,N_13544,N_13851);
and U14436 (N_14436,N_13743,N_13954);
nand U14437 (N_14437,N_13913,N_13630);
nand U14438 (N_14438,N_13582,N_13892);
or U14439 (N_14439,N_13756,N_13520);
or U14440 (N_14440,N_13923,N_13835);
nor U14441 (N_14441,N_13762,N_13625);
or U14442 (N_14442,N_13917,N_13883);
nor U14443 (N_14443,N_13896,N_13637);
nor U14444 (N_14444,N_13509,N_13757);
nor U14445 (N_14445,N_13578,N_13569);
nand U14446 (N_14446,N_13587,N_13732);
xor U14447 (N_14447,N_13597,N_13875);
and U14448 (N_14448,N_13668,N_13554);
nand U14449 (N_14449,N_13787,N_13921);
nor U14450 (N_14450,N_13710,N_13762);
nand U14451 (N_14451,N_13719,N_13967);
and U14452 (N_14452,N_13860,N_13975);
nor U14453 (N_14453,N_13858,N_13910);
nand U14454 (N_14454,N_13964,N_13555);
nand U14455 (N_14455,N_13629,N_13956);
nand U14456 (N_14456,N_13602,N_13611);
and U14457 (N_14457,N_13563,N_13609);
nor U14458 (N_14458,N_13821,N_13881);
or U14459 (N_14459,N_13846,N_13906);
and U14460 (N_14460,N_13572,N_13703);
xor U14461 (N_14461,N_13855,N_13903);
and U14462 (N_14462,N_13619,N_13853);
nand U14463 (N_14463,N_13901,N_13746);
nor U14464 (N_14464,N_13946,N_13793);
xor U14465 (N_14465,N_13698,N_13553);
nor U14466 (N_14466,N_13859,N_13631);
and U14467 (N_14467,N_13529,N_13819);
or U14468 (N_14468,N_13989,N_13619);
xnor U14469 (N_14469,N_13767,N_13966);
and U14470 (N_14470,N_13895,N_13940);
xor U14471 (N_14471,N_13747,N_13731);
and U14472 (N_14472,N_13839,N_13880);
or U14473 (N_14473,N_13849,N_13542);
and U14474 (N_14474,N_13753,N_13640);
xor U14475 (N_14475,N_13994,N_13802);
nor U14476 (N_14476,N_13703,N_13664);
xor U14477 (N_14477,N_13549,N_13630);
xnor U14478 (N_14478,N_13777,N_13572);
and U14479 (N_14479,N_13874,N_13949);
nor U14480 (N_14480,N_13714,N_13636);
nor U14481 (N_14481,N_13985,N_13576);
or U14482 (N_14482,N_13959,N_13948);
and U14483 (N_14483,N_13671,N_13763);
nand U14484 (N_14484,N_13567,N_13912);
and U14485 (N_14485,N_13583,N_13687);
nor U14486 (N_14486,N_13730,N_13767);
nand U14487 (N_14487,N_13599,N_13857);
nor U14488 (N_14488,N_13548,N_13603);
and U14489 (N_14489,N_13730,N_13742);
and U14490 (N_14490,N_13724,N_13668);
xnor U14491 (N_14491,N_13940,N_13727);
nor U14492 (N_14492,N_13726,N_13612);
or U14493 (N_14493,N_13661,N_13983);
nand U14494 (N_14494,N_13536,N_13561);
xnor U14495 (N_14495,N_13581,N_13638);
or U14496 (N_14496,N_13694,N_13813);
and U14497 (N_14497,N_13819,N_13816);
nor U14498 (N_14498,N_13560,N_13705);
nor U14499 (N_14499,N_13601,N_13828);
and U14500 (N_14500,N_14347,N_14415);
or U14501 (N_14501,N_14214,N_14029);
and U14502 (N_14502,N_14268,N_14438);
xor U14503 (N_14503,N_14264,N_14224);
or U14504 (N_14504,N_14297,N_14235);
or U14505 (N_14505,N_14336,N_14412);
nand U14506 (N_14506,N_14261,N_14435);
or U14507 (N_14507,N_14366,N_14309);
nand U14508 (N_14508,N_14335,N_14444);
nor U14509 (N_14509,N_14420,N_14094);
nand U14510 (N_14510,N_14051,N_14164);
or U14511 (N_14511,N_14463,N_14086);
and U14512 (N_14512,N_14240,N_14477);
nand U14513 (N_14513,N_14195,N_14315);
and U14514 (N_14514,N_14342,N_14471);
nor U14515 (N_14515,N_14220,N_14269);
and U14516 (N_14516,N_14197,N_14367);
nand U14517 (N_14517,N_14324,N_14166);
or U14518 (N_14518,N_14352,N_14329);
xnor U14519 (N_14519,N_14168,N_14263);
nor U14520 (N_14520,N_14497,N_14356);
nand U14521 (N_14521,N_14160,N_14149);
xor U14522 (N_14522,N_14408,N_14236);
or U14523 (N_14523,N_14440,N_14059);
and U14524 (N_14524,N_14380,N_14087);
nand U14525 (N_14525,N_14173,N_14428);
nand U14526 (N_14526,N_14486,N_14124);
or U14527 (N_14527,N_14141,N_14271);
or U14528 (N_14528,N_14256,N_14196);
xnor U14529 (N_14529,N_14257,N_14262);
or U14530 (N_14530,N_14354,N_14270);
nor U14531 (N_14531,N_14419,N_14301);
or U14532 (N_14532,N_14252,N_14016);
nor U14533 (N_14533,N_14298,N_14109);
nand U14534 (N_14534,N_14410,N_14212);
or U14535 (N_14535,N_14067,N_14012);
and U14536 (N_14536,N_14219,N_14439);
xor U14537 (N_14537,N_14260,N_14223);
or U14538 (N_14538,N_14392,N_14452);
nand U14539 (N_14539,N_14061,N_14243);
xor U14540 (N_14540,N_14343,N_14027);
nor U14541 (N_14541,N_14316,N_14221);
xnor U14542 (N_14542,N_14381,N_14421);
nand U14543 (N_14543,N_14348,N_14344);
or U14544 (N_14544,N_14484,N_14292);
nand U14545 (N_14545,N_14056,N_14206);
and U14546 (N_14546,N_14402,N_14165);
and U14547 (N_14547,N_14445,N_14287);
nand U14548 (N_14548,N_14038,N_14178);
and U14549 (N_14549,N_14281,N_14018);
nor U14550 (N_14550,N_14424,N_14154);
nand U14551 (N_14551,N_14093,N_14330);
nand U14552 (N_14552,N_14465,N_14098);
nand U14553 (N_14553,N_14218,N_14011);
and U14554 (N_14554,N_14288,N_14233);
nor U14555 (N_14555,N_14319,N_14377);
nand U14556 (N_14556,N_14110,N_14456);
nor U14557 (N_14557,N_14120,N_14009);
nand U14558 (N_14558,N_14142,N_14180);
xnor U14559 (N_14559,N_14250,N_14200);
nand U14560 (N_14560,N_14044,N_14395);
nor U14561 (N_14561,N_14085,N_14162);
nand U14562 (N_14562,N_14483,N_14429);
nor U14563 (N_14563,N_14215,N_14450);
or U14564 (N_14564,N_14161,N_14198);
nand U14565 (N_14565,N_14005,N_14425);
nand U14566 (N_14566,N_14432,N_14049);
xor U14567 (N_14567,N_14183,N_14474);
xnor U14568 (N_14568,N_14458,N_14186);
nor U14569 (N_14569,N_14308,N_14291);
nor U14570 (N_14570,N_14242,N_14095);
xor U14571 (N_14571,N_14290,N_14480);
nor U14572 (N_14572,N_14379,N_14313);
nor U14573 (N_14573,N_14090,N_14053);
xnor U14574 (N_14574,N_14418,N_14498);
xor U14575 (N_14575,N_14441,N_14157);
or U14576 (N_14576,N_14469,N_14464);
nor U14577 (N_14577,N_14394,N_14254);
or U14578 (N_14578,N_14184,N_14229);
xor U14579 (N_14579,N_14055,N_14150);
or U14580 (N_14580,N_14107,N_14487);
xnor U14581 (N_14581,N_14091,N_14000);
or U14582 (N_14582,N_14026,N_14286);
nor U14583 (N_14583,N_14489,N_14225);
nor U14584 (N_14584,N_14139,N_14265);
or U14585 (N_14585,N_14284,N_14013);
and U14586 (N_14586,N_14122,N_14131);
or U14587 (N_14587,N_14365,N_14217);
and U14588 (N_14588,N_14396,N_14404);
xnor U14589 (N_14589,N_14370,N_14430);
nand U14590 (N_14590,N_14072,N_14182);
and U14591 (N_14591,N_14436,N_14132);
nand U14592 (N_14592,N_14446,N_14117);
or U14593 (N_14593,N_14145,N_14070);
nand U14594 (N_14594,N_14434,N_14293);
nand U14595 (N_14595,N_14275,N_14378);
nor U14596 (N_14596,N_14064,N_14467);
nand U14597 (N_14597,N_14074,N_14314);
or U14598 (N_14598,N_14204,N_14478);
and U14599 (N_14599,N_14296,N_14159);
nand U14600 (N_14600,N_14065,N_14148);
and U14601 (N_14601,N_14023,N_14388);
nor U14602 (N_14602,N_14466,N_14244);
and U14603 (N_14603,N_14041,N_14353);
and U14604 (N_14604,N_14209,N_14391);
xnor U14605 (N_14605,N_14416,N_14062);
or U14606 (N_14606,N_14175,N_14136);
and U14607 (N_14607,N_14030,N_14099);
nand U14608 (N_14608,N_14128,N_14105);
nor U14609 (N_14609,N_14025,N_14312);
or U14610 (N_14610,N_14341,N_14205);
xnor U14611 (N_14611,N_14181,N_14285);
nor U14612 (N_14612,N_14040,N_14355);
nor U14613 (N_14613,N_14403,N_14066);
and U14614 (N_14614,N_14360,N_14177);
xor U14615 (N_14615,N_14002,N_14088);
xor U14616 (N_14616,N_14033,N_14024);
or U14617 (N_14617,N_14118,N_14202);
and U14618 (N_14618,N_14303,N_14100);
nor U14619 (N_14619,N_14376,N_14014);
nand U14620 (N_14620,N_14317,N_14406);
nand U14621 (N_14621,N_14082,N_14052);
nand U14622 (N_14622,N_14473,N_14310);
nand U14623 (N_14623,N_14143,N_14125);
or U14624 (N_14624,N_14102,N_14306);
xor U14625 (N_14625,N_14304,N_14300);
or U14626 (N_14626,N_14459,N_14192);
or U14627 (N_14627,N_14337,N_14171);
or U14628 (N_14628,N_14185,N_14389);
or U14629 (N_14629,N_14210,N_14199);
nor U14630 (N_14630,N_14302,N_14121);
and U14631 (N_14631,N_14442,N_14299);
nand U14632 (N_14632,N_14226,N_14147);
nand U14633 (N_14633,N_14008,N_14108);
xnor U14634 (N_14634,N_14015,N_14179);
and U14635 (N_14635,N_14328,N_14019);
or U14636 (N_14636,N_14111,N_14481);
xor U14637 (N_14637,N_14485,N_14476);
nand U14638 (N_14638,N_14273,N_14047);
nand U14639 (N_14639,N_14101,N_14375);
xnor U14640 (N_14640,N_14274,N_14211);
xnor U14641 (N_14641,N_14050,N_14039);
xnor U14642 (N_14642,N_14495,N_14045);
nor U14643 (N_14643,N_14151,N_14323);
and U14644 (N_14644,N_14282,N_14493);
nand U14645 (N_14645,N_14494,N_14208);
or U14646 (N_14646,N_14080,N_14021);
and U14647 (N_14647,N_14227,N_14228);
xnor U14648 (N_14648,N_14144,N_14321);
nand U14649 (N_14649,N_14248,N_14104);
nor U14650 (N_14650,N_14409,N_14455);
nand U14651 (N_14651,N_14077,N_14092);
xnor U14652 (N_14652,N_14245,N_14022);
nand U14653 (N_14653,N_14170,N_14081);
and U14654 (N_14654,N_14371,N_14449);
nor U14655 (N_14655,N_14462,N_14443);
and U14656 (N_14656,N_14238,N_14194);
and U14657 (N_14657,N_14345,N_14078);
nand U14658 (N_14658,N_14414,N_14373);
xor U14659 (N_14659,N_14350,N_14071);
and U14660 (N_14660,N_14239,N_14152);
and U14661 (N_14661,N_14411,N_14407);
nor U14662 (N_14662,N_14246,N_14326);
nor U14663 (N_14663,N_14318,N_14447);
nand U14664 (N_14664,N_14060,N_14325);
nor U14665 (N_14665,N_14037,N_14222);
nor U14666 (N_14666,N_14069,N_14032);
nand U14667 (N_14667,N_14338,N_14042);
nor U14668 (N_14668,N_14453,N_14133);
and U14669 (N_14669,N_14448,N_14167);
or U14670 (N_14670,N_14362,N_14174);
or U14671 (N_14671,N_14043,N_14358);
nor U14672 (N_14672,N_14004,N_14169);
nand U14673 (N_14673,N_14393,N_14451);
xor U14674 (N_14674,N_14028,N_14259);
and U14675 (N_14675,N_14126,N_14400);
nand U14676 (N_14676,N_14351,N_14340);
and U14677 (N_14677,N_14216,N_14146);
xnor U14678 (N_14678,N_14401,N_14470);
and U14679 (N_14679,N_14034,N_14433);
or U14680 (N_14680,N_14189,N_14073);
or U14681 (N_14681,N_14357,N_14106);
nand U14682 (N_14682,N_14007,N_14063);
nor U14683 (N_14683,N_14496,N_14334);
xnor U14684 (N_14684,N_14031,N_14390);
nand U14685 (N_14685,N_14305,N_14207);
or U14686 (N_14686,N_14491,N_14253);
nor U14687 (N_14687,N_14361,N_14156);
xnor U14688 (N_14688,N_14461,N_14279);
xnor U14689 (N_14689,N_14363,N_14413);
xor U14690 (N_14690,N_14158,N_14203);
nor U14691 (N_14691,N_14258,N_14490);
xnor U14692 (N_14692,N_14172,N_14454);
nand U14693 (N_14693,N_14331,N_14277);
nor U14694 (N_14694,N_14422,N_14475);
and U14695 (N_14695,N_14112,N_14488);
xor U14696 (N_14696,N_14127,N_14399);
xor U14697 (N_14697,N_14232,N_14193);
nand U14698 (N_14698,N_14096,N_14116);
and U14699 (N_14699,N_14255,N_14176);
nor U14700 (N_14700,N_14359,N_14083);
xor U14701 (N_14701,N_14398,N_14339);
nor U14702 (N_14702,N_14387,N_14384);
or U14703 (N_14703,N_14364,N_14048);
nor U14704 (N_14704,N_14247,N_14423);
and U14705 (N_14705,N_14130,N_14249);
nor U14706 (N_14706,N_14369,N_14190);
xor U14707 (N_14707,N_14084,N_14103);
or U14708 (N_14708,N_14266,N_14114);
or U14709 (N_14709,N_14213,N_14372);
xnor U14710 (N_14710,N_14427,N_14276);
xnor U14711 (N_14711,N_14006,N_14113);
and U14712 (N_14712,N_14251,N_14237);
and U14713 (N_14713,N_14138,N_14374);
or U14714 (N_14714,N_14241,N_14020);
nand U14715 (N_14715,N_14163,N_14322);
and U14716 (N_14716,N_14017,N_14472);
nor U14717 (N_14717,N_14135,N_14383);
and U14718 (N_14718,N_14346,N_14307);
nand U14719 (N_14719,N_14457,N_14129);
nor U14720 (N_14720,N_14385,N_14333);
xnor U14721 (N_14721,N_14230,N_14001);
or U14722 (N_14722,N_14320,N_14137);
or U14723 (N_14723,N_14003,N_14417);
and U14724 (N_14724,N_14283,N_14327);
or U14725 (N_14725,N_14231,N_14437);
nand U14726 (N_14726,N_14119,N_14057);
nor U14727 (N_14727,N_14123,N_14295);
and U14728 (N_14728,N_14035,N_14368);
xor U14729 (N_14729,N_14386,N_14115);
nand U14730 (N_14730,N_14201,N_14280);
or U14731 (N_14731,N_14479,N_14397);
nor U14732 (N_14732,N_14187,N_14332);
or U14733 (N_14733,N_14010,N_14294);
or U14734 (N_14734,N_14499,N_14153);
xor U14735 (N_14735,N_14405,N_14068);
nand U14736 (N_14736,N_14140,N_14482);
or U14737 (N_14737,N_14191,N_14089);
or U14738 (N_14738,N_14036,N_14054);
and U14739 (N_14739,N_14272,N_14058);
nand U14740 (N_14740,N_14075,N_14134);
nand U14741 (N_14741,N_14046,N_14076);
nor U14742 (N_14742,N_14234,N_14431);
or U14743 (N_14743,N_14492,N_14278);
and U14744 (N_14744,N_14188,N_14426);
and U14745 (N_14745,N_14289,N_14079);
or U14746 (N_14746,N_14382,N_14349);
and U14747 (N_14747,N_14155,N_14311);
or U14748 (N_14748,N_14468,N_14460);
nor U14749 (N_14749,N_14267,N_14097);
nand U14750 (N_14750,N_14219,N_14393);
nor U14751 (N_14751,N_14202,N_14182);
xnor U14752 (N_14752,N_14028,N_14108);
xor U14753 (N_14753,N_14257,N_14455);
or U14754 (N_14754,N_14043,N_14290);
nand U14755 (N_14755,N_14110,N_14170);
or U14756 (N_14756,N_14454,N_14315);
nor U14757 (N_14757,N_14425,N_14168);
nor U14758 (N_14758,N_14308,N_14079);
nand U14759 (N_14759,N_14285,N_14459);
nor U14760 (N_14760,N_14109,N_14320);
xnor U14761 (N_14761,N_14101,N_14341);
nor U14762 (N_14762,N_14137,N_14363);
nand U14763 (N_14763,N_14378,N_14442);
xnor U14764 (N_14764,N_14247,N_14443);
or U14765 (N_14765,N_14254,N_14113);
nand U14766 (N_14766,N_14401,N_14395);
xor U14767 (N_14767,N_14207,N_14131);
and U14768 (N_14768,N_14198,N_14115);
or U14769 (N_14769,N_14373,N_14407);
or U14770 (N_14770,N_14418,N_14392);
nor U14771 (N_14771,N_14436,N_14406);
and U14772 (N_14772,N_14039,N_14384);
nand U14773 (N_14773,N_14304,N_14114);
or U14774 (N_14774,N_14005,N_14378);
nand U14775 (N_14775,N_14481,N_14322);
or U14776 (N_14776,N_14214,N_14479);
nor U14777 (N_14777,N_14348,N_14309);
xor U14778 (N_14778,N_14024,N_14185);
nor U14779 (N_14779,N_14498,N_14401);
xnor U14780 (N_14780,N_14238,N_14042);
nor U14781 (N_14781,N_14127,N_14196);
and U14782 (N_14782,N_14139,N_14167);
xor U14783 (N_14783,N_14341,N_14137);
nor U14784 (N_14784,N_14172,N_14041);
or U14785 (N_14785,N_14023,N_14090);
and U14786 (N_14786,N_14337,N_14085);
nand U14787 (N_14787,N_14408,N_14133);
nor U14788 (N_14788,N_14005,N_14260);
nand U14789 (N_14789,N_14143,N_14124);
nor U14790 (N_14790,N_14252,N_14136);
and U14791 (N_14791,N_14224,N_14147);
or U14792 (N_14792,N_14219,N_14025);
nand U14793 (N_14793,N_14385,N_14325);
xnor U14794 (N_14794,N_14482,N_14042);
nand U14795 (N_14795,N_14121,N_14477);
or U14796 (N_14796,N_14128,N_14250);
nand U14797 (N_14797,N_14067,N_14453);
nand U14798 (N_14798,N_14142,N_14077);
xor U14799 (N_14799,N_14057,N_14349);
nand U14800 (N_14800,N_14272,N_14028);
xor U14801 (N_14801,N_14176,N_14031);
and U14802 (N_14802,N_14224,N_14498);
nand U14803 (N_14803,N_14456,N_14401);
nor U14804 (N_14804,N_14352,N_14290);
and U14805 (N_14805,N_14131,N_14381);
nand U14806 (N_14806,N_14087,N_14041);
xnor U14807 (N_14807,N_14049,N_14130);
xnor U14808 (N_14808,N_14186,N_14297);
and U14809 (N_14809,N_14480,N_14255);
nand U14810 (N_14810,N_14392,N_14168);
nor U14811 (N_14811,N_14202,N_14052);
nand U14812 (N_14812,N_14136,N_14176);
or U14813 (N_14813,N_14433,N_14088);
and U14814 (N_14814,N_14087,N_14385);
xnor U14815 (N_14815,N_14378,N_14206);
or U14816 (N_14816,N_14381,N_14150);
or U14817 (N_14817,N_14459,N_14165);
nand U14818 (N_14818,N_14263,N_14252);
nand U14819 (N_14819,N_14081,N_14320);
or U14820 (N_14820,N_14473,N_14097);
and U14821 (N_14821,N_14262,N_14188);
or U14822 (N_14822,N_14063,N_14144);
xor U14823 (N_14823,N_14428,N_14144);
or U14824 (N_14824,N_14395,N_14473);
nor U14825 (N_14825,N_14149,N_14013);
nor U14826 (N_14826,N_14477,N_14252);
or U14827 (N_14827,N_14310,N_14370);
nand U14828 (N_14828,N_14472,N_14492);
or U14829 (N_14829,N_14427,N_14210);
nor U14830 (N_14830,N_14303,N_14415);
and U14831 (N_14831,N_14276,N_14185);
and U14832 (N_14832,N_14489,N_14059);
nand U14833 (N_14833,N_14231,N_14052);
or U14834 (N_14834,N_14422,N_14061);
nand U14835 (N_14835,N_14102,N_14036);
or U14836 (N_14836,N_14309,N_14210);
xor U14837 (N_14837,N_14192,N_14396);
and U14838 (N_14838,N_14015,N_14476);
nor U14839 (N_14839,N_14456,N_14258);
nor U14840 (N_14840,N_14430,N_14067);
and U14841 (N_14841,N_14246,N_14134);
or U14842 (N_14842,N_14345,N_14390);
xnor U14843 (N_14843,N_14378,N_14306);
and U14844 (N_14844,N_14324,N_14413);
and U14845 (N_14845,N_14012,N_14268);
and U14846 (N_14846,N_14215,N_14386);
nor U14847 (N_14847,N_14409,N_14007);
nor U14848 (N_14848,N_14066,N_14057);
xnor U14849 (N_14849,N_14223,N_14251);
or U14850 (N_14850,N_14383,N_14032);
xor U14851 (N_14851,N_14139,N_14396);
or U14852 (N_14852,N_14210,N_14193);
nor U14853 (N_14853,N_14314,N_14272);
nand U14854 (N_14854,N_14463,N_14309);
and U14855 (N_14855,N_14349,N_14013);
nor U14856 (N_14856,N_14138,N_14451);
nand U14857 (N_14857,N_14357,N_14006);
xnor U14858 (N_14858,N_14345,N_14256);
xnor U14859 (N_14859,N_14025,N_14146);
xnor U14860 (N_14860,N_14440,N_14481);
xnor U14861 (N_14861,N_14266,N_14425);
and U14862 (N_14862,N_14234,N_14424);
nand U14863 (N_14863,N_14167,N_14148);
xor U14864 (N_14864,N_14440,N_14204);
or U14865 (N_14865,N_14166,N_14470);
nand U14866 (N_14866,N_14228,N_14117);
nor U14867 (N_14867,N_14081,N_14026);
nand U14868 (N_14868,N_14450,N_14276);
nand U14869 (N_14869,N_14112,N_14334);
or U14870 (N_14870,N_14014,N_14459);
and U14871 (N_14871,N_14187,N_14395);
xor U14872 (N_14872,N_14222,N_14418);
nor U14873 (N_14873,N_14486,N_14205);
or U14874 (N_14874,N_14059,N_14296);
nor U14875 (N_14875,N_14000,N_14194);
or U14876 (N_14876,N_14254,N_14333);
nand U14877 (N_14877,N_14419,N_14361);
xnor U14878 (N_14878,N_14323,N_14479);
or U14879 (N_14879,N_14169,N_14120);
nor U14880 (N_14880,N_14015,N_14359);
nor U14881 (N_14881,N_14243,N_14342);
or U14882 (N_14882,N_14152,N_14377);
and U14883 (N_14883,N_14248,N_14487);
nor U14884 (N_14884,N_14361,N_14340);
nor U14885 (N_14885,N_14314,N_14395);
xor U14886 (N_14886,N_14014,N_14434);
nand U14887 (N_14887,N_14449,N_14278);
nand U14888 (N_14888,N_14388,N_14256);
nor U14889 (N_14889,N_14306,N_14200);
nor U14890 (N_14890,N_14471,N_14415);
nand U14891 (N_14891,N_14052,N_14423);
nand U14892 (N_14892,N_14302,N_14143);
nor U14893 (N_14893,N_14468,N_14212);
and U14894 (N_14894,N_14485,N_14496);
nand U14895 (N_14895,N_14345,N_14392);
and U14896 (N_14896,N_14277,N_14149);
nor U14897 (N_14897,N_14065,N_14301);
nand U14898 (N_14898,N_14202,N_14249);
or U14899 (N_14899,N_14486,N_14405);
or U14900 (N_14900,N_14360,N_14062);
nor U14901 (N_14901,N_14463,N_14172);
or U14902 (N_14902,N_14170,N_14108);
or U14903 (N_14903,N_14329,N_14106);
and U14904 (N_14904,N_14081,N_14385);
and U14905 (N_14905,N_14491,N_14425);
nand U14906 (N_14906,N_14486,N_14406);
xnor U14907 (N_14907,N_14407,N_14083);
nand U14908 (N_14908,N_14281,N_14442);
nor U14909 (N_14909,N_14157,N_14108);
xnor U14910 (N_14910,N_14413,N_14247);
or U14911 (N_14911,N_14361,N_14468);
or U14912 (N_14912,N_14110,N_14338);
and U14913 (N_14913,N_14177,N_14421);
nor U14914 (N_14914,N_14369,N_14108);
or U14915 (N_14915,N_14029,N_14197);
nor U14916 (N_14916,N_14132,N_14195);
nand U14917 (N_14917,N_14337,N_14236);
and U14918 (N_14918,N_14337,N_14031);
nor U14919 (N_14919,N_14001,N_14014);
xor U14920 (N_14920,N_14116,N_14150);
xor U14921 (N_14921,N_14076,N_14490);
or U14922 (N_14922,N_14253,N_14278);
nand U14923 (N_14923,N_14201,N_14063);
xor U14924 (N_14924,N_14031,N_14053);
or U14925 (N_14925,N_14327,N_14133);
xnor U14926 (N_14926,N_14395,N_14128);
xor U14927 (N_14927,N_14287,N_14373);
nor U14928 (N_14928,N_14143,N_14343);
nor U14929 (N_14929,N_14295,N_14134);
nor U14930 (N_14930,N_14289,N_14150);
nor U14931 (N_14931,N_14125,N_14480);
and U14932 (N_14932,N_14153,N_14265);
xor U14933 (N_14933,N_14386,N_14307);
or U14934 (N_14934,N_14299,N_14199);
or U14935 (N_14935,N_14358,N_14445);
xor U14936 (N_14936,N_14161,N_14370);
nor U14937 (N_14937,N_14344,N_14144);
xor U14938 (N_14938,N_14093,N_14417);
or U14939 (N_14939,N_14189,N_14205);
nor U14940 (N_14940,N_14053,N_14202);
xor U14941 (N_14941,N_14207,N_14127);
or U14942 (N_14942,N_14358,N_14090);
or U14943 (N_14943,N_14114,N_14092);
nand U14944 (N_14944,N_14337,N_14207);
and U14945 (N_14945,N_14211,N_14270);
or U14946 (N_14946,N_14189,N_14484);
or U14947 (N_14947,N_14127,N_14380);
or U14948 (N_14948,N_14214,N_14224);
nor U14949 (N_14949,N_14016,N_14443);
nand U14950 (N_14950,N_14278,N_14277);
nor U14951 (N_14951,N_14069,N_14374);
and U14952 (N_14952,N_14036,N_14379);
nand U14953 (N_14953,N_14151,N_14427);
and U14954 (N_14954,N_14043,N_14231);
nand U14955 (N_14955,N_14460,N_14247);
or U14956 (N_14956,N_14050,N_14074);
nand U14957 (N_14957,N_14255,N_14192);
and U14958 (N_14958,N_14118,N_14435);
and U14959 (N_14959,N_14035,N_14011);
or U14960 (N_14960,N_14423,N_14132);
xor U14961 (N_14961,N_14491,N_14347);
nor U14962 (N_14962,N_14130,N_14258);
or U14963 (N_14963,N_14317,N_14277);
nor U14964 (N_14964,N_14293,N_14165);
xnor U14965 (N_14965,N_14416,N_14253);
or U14966 (N_14966,N_14451,N_14217);
nand U14967 (N_14967,N_14452,N_14474);
or U14968 (N_14968,N_14462,N_14010);
or U14969 (N_14969,N_14367,N_14271);
xor U14970 (N_14970,N_14441,N_14311);
and U14971 (N_14971,N_14272,N_14440);
xor U14972 (N_14972,N_14253,N_14296);
nand U14973 (N_14973,N_14048,N_14311);
or U14974 (N_14974,N_14282,N_14494);
nor U14975 (N_14975,N_14029,N_14069);
or U14976 (N_14976,N_14296,N_14094);
nand U14977 (N_14977,N_14456,N_14280);
xnor U14978 (N_14978,N_14312,N_14428);
and U14979 (N_14979,N_14056,N_14219);
nand U14980 (N_14980,N_14116,N_14115);
or U14981 (N_14981,N_14003,N_14013);
and U14982 (N_14982,N_14041,N_14363);
and U14983 (N_14983,N_14355,N_14372);
and U14984 (N_14984,N_14262,N_14316);
and U14985 (N_14985,N_14145,N_14316);
nand U14986 (N_14986,N_14191,N_14218);
nor U14987 (N_14987,N_14336,N_14425);
nor U14988 (N_14988,N_14161,N_14190);
nand U14989 (N_14989,N_14120,N_14306);
xor U14990 (N_14990,N_14175,N_14106);
xnor U14991 (N_14991,N_14496,N_14224);
and U14992 (N_14992,N_14367,N_14147);
nand U14993 (N_14993,N_14449,N_14221);
nand U14994 (N_14994,N_14380,N_14239);
or U14995 (N_14995,N_14432,N_14474);
xor U14996 (N_14996,N_14212,N_14495);
and U14997 (N_14997,N_14242,N_14267);
nor U14998 (N_14998,N_14066,N_14208);
xnor U14999 (N_14999,N_14130,N_14214);
or U15000 (N_15000,N_14617,N_14619);
and U15001 (N_15001,N_14995,N_14542);
and U15002 (N_15002,N_14695,N_14723);
and U15003 (N_15003,N_14680,N_14763);
nand U15004 (N_15004,N_14788,N_14981);
or U15005 (N_15005,N_14940,N_14814);
and U15006 (N_15006,N_14878,N_14669);
or U15007 (N_15007,N_14556,N_14861);
or U15008 (N_15008,N_14736,N_14716);
xnor U15009 (N_15009,N_14922,N_14785);
or U15010 (N_15010,N_14720,N_14510);
nor U15011 (N_15011,N_14694,N_14620);
nor U15012 (N_15012,N_14943,N_14744);
and U15013 (N_15013,N_14772,N_14590);
xor U15014 (N_15014,N_14708,N_14595);
nand U15015 (N_15015,N_14894,N_14836);
xor U15016 (N_15016,N_14851,N_14578);
xnor U15017 (N_15017,N_14954,N_14531);
nor U15018 (N_15018,N_14895,N_14982);
xnor U15019 (N_15019,N_14541,N_14855);
xor U15020 (N_15020,N_14914,N_14864);
nand U15021 (N_15021,N_14508,N_14874);
or U15022 (N_15022,N_14916,N_14656);
or U15023 (N_15023,N_14699,N_14593);
xor U15024 (N_15024,N_14516,N_14659);
xnor U15025 (N_15025,N_14948,N_14751);
and U15026 (N_15026,N_14887,N_14946);
nand U15027 (N_15027,N_14910,N_14777);
or U15028 (N_15028,N_14555,N_14920);
or U15029 (N_15029,N_14935,N_14858);
or U15030 (N_15030,N_14667,N_14997);
or U15031 (N_15031,N_14696,N_14882);
xnor U15032 (N_15032,N_14631,N_14759);
nand U15033 (N_15033,N_14765,N_14934);
and U15034 (N_15034,N_14719,N_14521);
and U15035 (N_15035,N_14950,N_14811);
or U15036 (N_15036,N_14726,N_14601);
xnor U15037 (N_15037,N_14615,N_14813);
nand U15038 (N_15038,N_14728,N_14762);
and U15039 (N_15039,N_14599,N_14947);
nand U15040 (N_15040,N_14626,N_14921);
xnor U15041 (N_15041,N_14580,N_14609);
xor U15042 (N_15042,N_14875,N_14941);
nor U15043 (N_15043,N_14579,N_14775);
xor U15044 (N_15044,N_14808,N_14640);
xnor U15045 (N_15045,N_14816,N_14803);
nand U15046 (N_15046,N_14819,N_14583);
nor U15047 (N_15047,N_14827,N_14953);
nor U15048 (N_15048,N_14526,N_14702);
nor U15049 (N_15049,N_14829,N_14919);
nor U15050 (N_15050,N_14789,N_14662);
nor U15051 (N_15051,N_14956,N_14932);
and U15052 (N_15052,N_14833,N_14629);
or U15053 (N_15053,N_14801,N_14884);
or U15054 (N_15054,N_14989,N_14581);
and U15055 (N_15055,N_14553,N_14831);
and U15056 (N_15056,N_14515,N_14890);
nor U15057 (N_15057,N_14797,N_14877);
nand U15058 (N_15058,N_14704,N_14820);
nor U15059 (N_15059,N_14928,N_14781);
nor U15060 (N_15060,N_14681,N_14905);
xor U15061 (N_15061,N_14652,N_14738);
or U15062 (N_15062,N_14577,N_14733);
and U15063 (N_15063,N_14976,N_14891);
or U15064 (N_15064,N_14650,N_14970);
nand U15065 (N_15065,N_14771,N_14821);
and U15066 (N_15066,N_14835,N_14859);
nand U15067 (N_15067,N_14929,N_14540);
nor U15068 (N_15068,N_14822,N_14588);
nand U15069 (N_15069,N_14944,N_14841);
or U15070 (N_15070,N_14984,N_14883);
and U15071 (N_15071,N_14826,N_14660);
nor U15072 (N_15072,N_14621,N_14769);
xor U15073 (N_15073,N_14565,N_14604);
xnor U15074 (N_15074,N_14800,N_14655);
nor U15075 (N_15075,N_14624,N_14679);
nor U15076 (N_15076,N_14727,N_14725);
or U15077 (N_15077,N_14994,N_14690);
xor U15078 (N_15078,N_14558,N_14548);
xnor U15079 (N_15079,N_14676,N_14721);
and U15080 (N_15080,N_14501,N_14697);
nand U15081 (N_15081,N_14589,N_14790);
nand U15082 (N_15082,N_14546,N_14575);
nand U15083 (N_15083,N_14828,N_14776);
xnor U15084 (N_15084,N_14670,N_14706);
nand U15085 (N_15085,N_14570,N_14915);
nand U15086 (N_15086,N_14730,N_14572);
nor U15087 (N_15087,N_14974,N_14825);
nand U15088 (N_15088,N_14533,N_14839);
xnor U15089 (N_15089,N_14886,N_14566);
nor U15090 (N_15090,N_14748,N_14684);
and U15091 (N_15091,N_14585,N_14661);
and U15092 (N_15092,N_14698,N_14938);
or U15093 (N_15093,N_14972,N_14709);
and U15094 (N_15094,N_14511,N_14608);
xor U15095 (N_15095,N_14627,N_14849);
xor U15096 (N_15096,N_14517,N_14605);
or U15097 (N_15097,N_14823,N_14668);
nand U15098 (N_15098,N_14830,N_14732);
nand U15099 (N_15099,N_14591,N_14971);
nor U15100 (N_15100,N_14688,N_14779);
and U15101 (N_15101,N_14795,N_14647);
or U15102 (N_15102,N_14646,N_14643);
or U15103 (N_15103,N_14966,N_14635);
or U15104 (N_15104,N_14991,N_14717);
nor U15105 (N_15105,N_14898,N_14587);
and U15106 (N_15106,N_14569,N_14793);
xor U15107 (N_15107,N_14806,N_14965);
and U15108 (N_15108,N_14529,N_14752);
nand U15109 (N_15109,N_14682,N_14610);
xor U15110 (N_15110,N_14628,N_14675);
nor U15111 (N_15111,N_14550,N_14737);
nor U15112 (N_15112,N_14507,N_14513);
nor U15113 (N_15113,N_14783,N_14852);
and U15114 (N_15114,N_14996,N_14923);
nor U15115 (N_15115,N_14912,N_14663);
xnor U15116 (N_15116,N_14975,N_14597);
xnor U15117 (N_15117,N_14959,N_14651);
nand U15118 (N_15118,N_14504,N_14623);
or U15119 (N_15119,N_14871,N_14584);
nand U15120 (N_15120,N_14798,N_14753);
xor U15121 (N_15121,N_14917,N_14774);
xor U15122 (N_15122,N_14952,N_14638);
nor U15123 (N_15123,N_14536,N_14764);
nor U15124 (N_15124,N_14700,N_14901);
or U15125 (N_15125,N_14527,N_14892);
nor U15126 (N_15126,N_14868,N_14547);
and U15127 (N_15127,N_14850,N_14936);
xnor U15128 (N_15128,N_14760,N_14881);
nand U15129 (N_15129,N_14809,N_14673);
nand U15130 (N_15130,N_14794,N_14707);
xor U15131 (N_15131,N_14685,N_14862);
xor U15132 (N_15132,N_14664,N_14523);
and U15133 (N_15133,N_14710,N_14909);
xor U15134 (N_15134,N_14955,N_14896);
or U15135 (N_15135,N_14576,N_14724);
nand U15136 (N_15136,N_14927,N_14973);
nor U15137 (N_15137,N_14987,N_14957);
and U15138 (N_15138,N_14666,N_14903);
xnor U15139 (N_15139,N_14714,N_14860);
nor U15140 (N_15140,N_14530,N_14622);
xor U15141 (N_15141,N_14741,N_14613);
xnor U15142 (N_15142,N_14552,N_14743);
nand U15143 (N_15143,N_14939,N_14644);
and U15144 (N_15144,N_14766,N_14693);
xnor U15145 (N_15145,N_14596,N_14543);
nor U15146 (N_15146,N_14722,N_14857);
nand U15147 (N_15147,N_14844,N_14761);
and U15148 (N_15148,N_14999,N_14992);
or U15149 (N_15149,N_14977,N_14782);
nor U15150 (N_15150,N_14592,N_14880);
or U15151 (N_15151,N_14930,N_14978);
xor U15152 (N_15152,N_14648,N_14888);
nor U15153 (N_15153,N_14554,N_14900);
nor U15154 (N_15154,N_14557,N_14602);
and U15155 (N_15155,N_14968,N_14879);
nor U15156 (N_15156,N_14600,N_14846);
and U15157 (N_15157,N_14799,N_14865);
and U15158 (N_15158,N_14632,N_14586);
and U15159 (N_15159,N_14757,N_14740);
or U15160 (N_15160,N_14747,N_14838);
xor U15161 (N_15161,N_14845,N_14606);
and U15162 (N_15162,N_14525,N_14870);
nor U15163 (N_15163,N_14969,N_14926);
or U15164 (N_15164,N_14869,N_14653);
nand U15165 (N_15165,N_14739,N_14678);
nand U15166 (N_15166,N_14742,N_14958);
xnor U15167 (N_15167,N_14840,N_14853);
xor U15168 (N_15168,N_14812,N_14848);
and U15169 (N_15169,N_14979,N_14949);
xnor U15170 (N_15170,N_14756,N_14746);
nor U15171 (N_15171,N_14689,N_14847);
nand U15172 (N_15172,N_14791,N_14674);
nor U15173 (N_15173,N_14594,N_14645);
and U15174 (N_15174,N_14522,N_14634);
nand U15175 (N_15175,N_14778,N_14780);
nand U15176 (N_15176,N_14711,N_14715);
nor U15177 (N_15177,N_14961,N_14642);
nand U15178 (N_15178,N_14832,N_14786);
nor U15179 (N_15179,N_14641,N_14639);
or U15180 (N_15180,N_14683,N_14654);
or U15181 (N_15181,N_14665,N_14918);
and U15182 (N_15182,N_14563,N_14734);
and U15183 (N_15183,N_14911,N_14990);
nor U15184 (N_15184,N_14983,N_14805);
xnor U15185 (N_15185,N_14562,N_14902);
xnor U15186 (N_15186,N_14560,N_14960);
and U15187 (N_15187,N_14962,N_14559);
and U15188 (N_15188,N_14537,N_14856);
or U15189 (N_15189,N_14993,N_14837);
or U15190 (N_15190,N_14768,N_14773);
or U15191 (N_15191,N_14512,N_14754);
xnor U15192 (N_15192,N_14749,N_14658);
or U15193 (N_15193,N_14503,N_14636);
nand U15194 (N_15194,N_14951,N_14770);
and U15195 (N_15195,N_14692,N_14571);
or U15196 (N_15196,N_14897,N_14872);
nor U15197 (N_15197,N_14863,N_14607);
xnor U15198 (N_15198,N_14933,N_14931);
nor U15199 (N_15199,N_14630,N_14866);
or U15200 (N_15200,N_14924,N_14582);
xnor U15201 (N_15201,N_14598,N_14980);
or U15202 (N_15202,N_14904,N_14899);
and U15203 (N_15203,N_14672,N_14637);
or U15204 (N_15204,N_14534,N_14514);
or U15205 (N_15205,N_14677,N_14535);
nor U15206 (N_15206,N_14889,N_14614);
and U15207 (N_15207,N_14500,N_14625);
nor U15208 (N_15208,N_14519,N_14810);
and U15209 (N_15209,N_14985,N_14561);
nor U15210 (N_15210,N_14731,N_14551);
nor U15211 (N_15211,N_14574,N_14701);
nand U15212 (N_15212,N_14854,N_14885);
or U15213 (N_15213,N_14796,N_14573);
or U15214 (N_15214,N_14817,N_14906);
nand U15215 (N_15215,N_14712,N_14925);
and U15216 (N_15216,N_14502,N_14568);
and U15217 (N_15217,N_14818,N_14611);
nor U15218 (N_15218,N_14633,N_14532);
or U15219 (N_15219,N_14815,N_14998);
and U15220 (N_15220,N_14942,N_14705);
or U15221 (N_15221,N_14967,N_14787);
or U15222 (N_15222,N_14767,N_14758);
nor U15223 (N_15223,N_14729,N_14755);
or U15224 (N_15224,N_14893,N_14691);
nand U15225 (N_15225,N_14657,N_14745);
xor U15226 (N_15226,N_14671,N_14509);
and U15227 (N_15227,N_14686,N_14687);
or U15228 (N_15228,N_14713,N_14528);
and U15229 (N_15229,N_14907,N_14544);
nor U15230 (N_15230,N_14567,N_14612);
or U15231 (N_15231,N_14802,N_14807);
or U15232 (N_15232,N_14986,N_14618);
and U15233 (N_15233,N_14518,N_14804);
or U15234 (N_15234,N_14538,N_14549);
nand U15235 (N_15235,N_14988,N_14718);
or U15236 (N_15236,N_14735,N_14964);
and U15237 (N_15237,N_14703,N_14524);
nor U15238 (N_15238,N_14963,N_14792);
or U15239 (N_15239,N_14505,N_14616);
and U15240 (N_15240,N_14750,N_14843);
or U15241 (N_15241,N_14564,N_14603);
or U15242 (N_15242,N_14908,N_14867);
and U15243 (N_15243,N_14937,N_14506);
nor U15244 (N_15244,N_14545,N_14873);
or U15245 (N_15245,N_14539,N_14876);
nor U15246 (N_15246,N_14945,N_14913);
and U15247 (N_15247,N_14649,N_14520);
xor U15248 (N_15248,N_14842,N_14784);
nor U15249 (N_15249,N_14824,N_14834);
nor U15250 (N_15250,N_14891,N_14596);
nand U15251 (N_15251,N_14530,N_14705);
and U15252 (N_15252,N_14544,N_14913);
xor U15253 (N_15253,N_14504,N_14712);
nor U15254 (N_15254,N_14539,N_14579);
and U15255 (N_15255,N_14749,N_14763);
nor U15256 (N_15256,N_14689,N_14970);
nand U15257 (N_15257,N_14642,N_14648);
nor U15258 (N_15258,N_14531,N_14781);
nor U15259 (N_15259,N_14791,N_14789);
nand U15260 (N_15260,N_14539,N_14849);
xnor U15261 (N_15261,N_14893,N_14703);
nor U15262 (N_15262,N_14836,N_14739);
or U15263 (N_15263,N_14847,N_14812);
or U15264 (N_15264,N_14590,N_14578);
nand U15265 (N_15265,N_14617,N_14643);
nor U15266 (N_15266,N_14678,N_14633);
and U15267 (N_15267,N_14936,N_14700);
or U15268 (N_15268,N_14624,N_14585);
nor U15269 (N_15269,N_14871,N_14617);
nor U15270 (N_15270,N_14788,N_14724);
or U15271 (N_15271,N_14765,N_14939);
or U15272 (N_15272,N_14984,N_14973);
xnor U15273 (N_15273,N_14718,N_14531);
nand U15274 (N_15274,N_14689,N_14619);
or U15275 (N_15275,N_14648,N_14685);
nand U15276 (N_15276,N_14579,N_14748);
and U15277 (N_15277,N_14664,N_14634);
or U15278 (N_15278,N_14834,N_14731);
xnor U15279 (N_15279,N_14526,N_14753);
xnor U15280 (N_15280,N_14634,N_14586);
and U15281 (N_15281,N_14660,N_14514);
nor U15282 (N_15282,N_14537,N_14556);
xnor U15283 (N_15283,N_14997,N_14625);
nor U15284 (N_15284,N_14852,N_14693);
nor U15285 (N_15285,N_14942,N_14917);
nand U15286 (N_15286,N_14890,N_14989);
or U15287 (N_15287,N_14654,N_14575);
or U15288 (N_15288,N_14567,N_14930);
xnor U15289 (N_15289,N_14827,N_14742);
and U15290 (N_15290,N_14916,N_14698);
and U15291 (N_15291,N_14588,N_14961);
xnor U15292 (N_15292,N_14868,N_14789);
nand U15293 (N_15293,N_14948,N_14718);
nor U15294 (N_15294,N_14665,N_14797);
or U15295 (N_15295,N_14945,N_14527);
nand U15296 (N_15296,N_14883,N_14943);
and U15297 (N_15297,N_14770,N_14847);
xor U15298 (N_15298,N_14717,N_14736);
and U15299 (N_15299,N_14604,N_14721);
and U15300 (N_15300,N_14845,N_14683);
nand U15301 (N_15301,N_14711,N_14598);
nand U15302 (N_15302,N_14732,N_14507);
and U15303 (N_15303,N_14839,N_14920);
nor U15304 (N_15304,N_14668,N_14667);
or U15305 (N_15305,N_14589,N_14629);
nand U15306 (N_15306,N_14719,N_14850);
xor U15307 (N_15307,N_14953,N_14845);
xor U15308 (N_15308,N_14619,N_14741);
nor U15309 (N_15309,N_14575,N_14925);
nor U15310 (N_15310,N_14597,N_14910);
and U15311 (N_15311,N_14903,N_14956);
nand U15312 (N_15312,N_14509,N_14912);
nor U15313 (N_15313,N_14718,N_14605);
xor U15314 (N_15314,N_14600,N_14576);
nor U15315 (N_15315,N_14692,N_14579);
nand U15316 (N_15316,N_14597,N_14911);
nor U15317 (N_15317,N_14857,N_14840);
nand U15318 (N_15318,N_14701,N_14507);
or U15319 (N_15319,N_14649,N_14604);
or U15320 (N_15320,N_14938,N_14726);
nor U15321 (N_15321,N_14596,N_14892);
xor U15322 (N_15322,N_14536,N_14703);
or U15323 (N_15323,N_14536,N_14561);
and U15324 (N_15324,N_14737,N_14908);
or U15325 (N_15325,N_14538,N_14859);
and U15326 (N_15326,N_14789,N_14792);
xnor U15327 (N_15327,N_14520,N_14928);
nor U15328 (N_15328,N_14843,N_14880);
nand U15329 (N_15329,N_14593,N_14980);
nand U15330 (N_15330,N_14553,N_14963);
nand U15331 (N_15331,N_14516,N_14673);
and U15332 (N_15332,N_14606,N_14583);
and U15333 (N_15333,N_14668,N_14530);
xnor U15334 (N_15334,N_14847,N_14995);
xnor U15335 (N_15335,N_14680,N_14729);
nor U15336 (N_15336,N_14667,N_14569);
xor U15337 (N_15337,N_14922,N_14835);
xor U15338 (N_15338,N_14630,N_14796);
xnor U15339 (N_15339,N_14988,N_14539);
xor U15340 (N_15340,N_14949,N_14640);
nand U15341 (N_15341,N_14665,N_14822);
or U15342 (N_15342,N_14830,N_14851);
nor U15343 (N_15343,N_14599,N_14830);
or U15344 (N_15344,N_14789,N_14586);
and U15345 (N_15345,N_14790,N_14713);
and U15346 (N_15346,N_14942,N_14627);
and U15347 (N_15347,N_14908,N_14583);
nand U15348 (N_15348,N_14932,N_14850);
and U15349 (N_15349,N_14640,N_14711);
nand U15350 (N_15350,N_14651,N_14687);
nand U15351 (N_15351,N_14731,N_14873);
nand U15352 (N_15352,N_14662,N_14841);
nand U15353 (N_15353,N_14599,N_14913);
xor U15354 (N_15354,N_14922,N_14665);
nor U15355 (N_15355,N_14832,N_14637);
nand U15356 (N_15356,N_14987,N_14677);
nor U15357 (N_15357,N_14824,N_14531);
or U15358 (N_15358,N_14607,N_14803);
or U15359 (N_15359,N_14676,N_14870);
nor U15360 (N_15360,N_14604,N_14970);
nand U15361 (N_15361,N_14627,N_14917);
or U15362 (N_15362,N_14581,N_14654);
or U15363 (N_15363,N_14580,N_14799);
nand U15364 (N_15364,N_14667,N_14930);
nor U15365 (N_15365,N_14931,N_14786);
xnor U15366 (N_15366,N_14753,N_14861);
or U15367 (N_15367,N_14712,N_14645);
or U15368 (N_15368,N_14813,N_14816);
nor U15369 (N_15369,N_14876,N_14566);
and U15370 (N_15370,N_14616,N_14911);
xnor U15371 (N_15371,N_14990,N_14935);
and U15372 (N_15372,N_14631,N_14666);
and U15373 (N_15373,N_14878,N_14890);
or U15374 (N_15374,N_14604,N_14939);
xor U15375 (N_15375,N_14715,N_14782);
and U15376 (N_15376,N_14970,N_14547);
nand U15377 (N_15377,N_14540,N_14571);
nand U15378 (N_15378,N_14722,N_14509);
nor U15379 (N_15379,N_14796,N_14883);
nor U15380 (N_15380,N_14871,N_14697);
nor U15381 (N_15381,N_14897,N_14573);
and U15382 (N_15382,N_14672,N_14633);
xnor U15383 (N_15383,N_14956,N_14920);
or U15384 (N_15384,N_14662,N_14553);
and U15385 (N_15385,N_14779,N_14570);
nor U15386 (N_15386,N_14949,N_14772);
or U15387 (N_15387,N_14941,N_14510);
or U15388 (N_15388,N_14603,N_14771);
and U15389 (N_15389,N_14640,N_14953);
nand U15390 (N_15390,N_14824,N_14783);
xor U15391 (N_15391,N_14650,N_14666);
or U15392 (N_15392,N_14930,N_14620);
nand U15393 (N_15393,N_14926,N_14797);
nand U15394 (N_15394,N_14926,N_14826);
xor U15395 (N_15395,N_14982,N_14994);
nor U15396 (N_15396,N_14839,N_14802);
nand U15397 (N_15397,N_14621,N_14505);
nor U15398 (N_15398,N_14667,N_14916);
nand U15399 (N_15399,N_14646,N_14832);
xor U15400 (N_15400,N_14538,N_14664);
and U15401 (N_15401,N_14533,N_14673);
or U15402 (N_15402,N_14714,N_14984);
nor U15403 (N_15403,N_14792,N_14689);
and U15404 (N_15404,N_14717,N_14879);
nand U15405 (N_15405,N_14577,N_14967);
nor U15406 (N_15406,N_14695,N_14522);
nor U15407 (N_15407,N_14813,N_14679);
nor U15408 (N_15408,N_14645,N_14723);
nand U15409 (N_15409,N_14922,N_14858);
nor U15410 (N_15410,N_14971,N_14539);
or U15411 (N_15411,N_14556,N_14708);
and U15412 (N_15412,N_14704,N_14963);
xor U15413 (N_15413,N_14848,N_14627);
and U15414 (N_15414,N_14523,N_14710);
nand U15415 (N_15415,N_14968,N_14785);
nand U15416 (N_15416,N_14912,N_14856);
or U15417 (N_15417,N_14848,N_14781);
xor U15418 (N_15418,N_14670,N_14896);
nand U15419 (N_15419,N_14940,N_14596);
xor U15420 (N_15420,N_14839,N_14503);
nor U15421 (N_15421,N_14871,N_14785);
nand U15422 (N_15422,N_14538,N_14552);
nand U15423 (N_15423,N_14753,N_14949);
and U15424 (N_15424,N_14687,N_14520);
or U15425 (N_15425,N_14605,N_14585);
nand U15426 (N_15426,N_14752,N_14590);
nand U15427 (N_15427,N_14967,N_14944);
xnor U15428 (N_15428,N_14981,N_14586);
and U15429 (N_15429,N_14924,N_14896);
or U15430 (N_15430,N_14918,N_14644);
nand U15431 (N_15431,N_14820,N_14594);
nor U15432 (N_15432,N_14847,N_14889);
or U15433 (N_15433,N_14588,N_14754);
and U15434 (N_15434,N_14931,N_14725);
or U15435 (N_15435,N_14632,N_14557);
or U15436 (N_15436,N_14580,N_14952);
xnor U15437 (N_15437,N_14726,N_14840);
or U15438 (N_15438,N_14680,N_14689);
or U15439 (N_15439,N_14746,N_14720);
xor U15440 (N_15440,N_14642,N_14617);
and U15441 (N_15441,N_14707,N_14688);
or U15442 (N_15442,N_14507,N_14823);
and U15443 (N_15443,N_14924,N_14929);
or U15444 (N_15444,N_14990,N_14522);
or U15445 (N_15445,N_14624,N_14517);
xnor U15446 (N_15446,N_14929,N_14953);
or U15447 (N_15447,N_14519,N_14511);
and U15448 (N_15448,N_14849,N_14598);
xnor U15449 (N_15449,N_14893,N_14775);
xnor U15450 (N_15450,N_14755,N_14510);
or U15451 (N_15451,N_14928,N_14972);
or U15452 (N_15452,N_14518,N_14814);
xor U15453 (N_15453,N_14538,N_14663);
and U15454 (N_15454,N_14664,N_14539);
and U15455 (N_15455,N_14553,N_14630);
and U15456 (N_15456,N_14745,N_14783);
nand U15457 (N_15457,N_14589,N_14769);
nor U15458 (N_15458,N_14897,N_14787);
nand U15459 (N_15459,N_14847,N_14693);
or U15460 (N_15460,N_14969,N_14526);
nand U15461 (N_15461,N_14944,N_14559);
and U15462 (N_15462,N_14765,N_14692);
and U15463 (N_15463,N_14969,N_14906);
and U15464 (N_15464,N_14634,N_14841);
and U15465 (N_15465,N_14678,N_14773);
or U15466 (N_15466,N_14741,N_14852);
nor U15467 (N_15467,N_14574,N_14860);
nand U15468 (N_15468,N_14621,N_14645);
xor U15469 (N_15469,N_14616,N_14636);
xnor U15470 (N_15470,N_14812,N_14609);
xor U15471 (N_15471,N_14742,N_14679);
or U15472 (N_15472,N_14871,N_14642);
nor U15473 (N_15473,N_14552,N_14726);
or U15474 (N_15474,N_14601,N_14543);
xor U15475 (N_15475,N_14595,N_14787);
or U15476 (N_15476,N_14693,N_14664);
and U15477 (N_15477,N_14754,N_14971);
or U15478 (N_15478,N_14963,N_14752);
xor U15479 (N_15479,N_14551,N_14523);
or U15480 (N_15480,N_14895,N_14578);
nor U15481 (N_15481,N_14639,N_14791);
or U15482 (N_15482,N_14567,N_14749);
nand U15483 (N_15483,N_14624,N_14560);
and U15484 (N_15484,N_14811,N_14778);
and U15485 (N_15485,N_14685,N_14878);
and U15486 (N_15486,N_14914,N_14614);
nand U15487 (N_15487,N_14861,N_14647);
xnor U15488 (N_15488,N_14645,N_14557);
xnor U15489 (N_15489,N_14524,N_14615);
nand U15490 (N_15490,N_14514,N_14793);
or U15491 (N_15491,N_14581,N_14835);
xnor U15492 (N_15492,N_14698,N_14784);
or U15493 (N_15493,N_14731,N_14618);
or U15494 (N_15494,N_14828,N_14623);
and U15495 (N_15495,N_14596,N_14536);
or U15496 (N_15496,N_14519,N_14722);
xor U15497 (N_15497,N_14549,N_14502);
nand U15498 (N_15498,N_14807,N_14754);
or U15499 (N_15499,N_14518,N_14963);
and U15500 (N_15500,N_15037,N_15492);
or U15501 (N_15501,N_15407,N_15482);
xnor U15502 (N_15502,N_15024,N_15113);
and U15503 (N_15503,N_15493,N_15063);
xor U15504 (N_15504,N_15296,N_15123);
nand U15505 (N_15505,N_15404,N_15405);
xor U15506 (N_15506,N_15495,N_15274);
nor U15507 (N_15507,N_15322,N_15246);
and U15508 (N_15508,N_15109,N_15031);
nor U15509 (N_15509,N_15114,N_15145);
or U15510 (N_15510,N_15272,N_15427);
and U15511 (N_15511,N_15172,N_15294);
nand U15512 (N_15512,N_15429,N_15267);
and U15513 (N_15513,N_15039,N_15112);
nand U15514 (N_15514,N_15140,N_15319);
nand U15515 (N_15515,N_15364,N_15009);
and U15516 (N_15516,N_15257,N_15194);
nand U15517 (N_15517,N_15342,N_15350);
or U15518 (N_15518,N_15305,N_15491);
nor U15519 (N_15519,N_15196,N_15358);
nand U15520 (N_15520,N_15215,N_15415);
xnor U15521 (N_15521,N_15012,N_15264);
or U15522 (N_15522,N_15268,N_15078);
nor U15523 (N_15523,N_15291,N_15421);
nor U15524 (N_15524,N_15248,N_15065);
nor U15525 (N_15525,N_15046,N_15420);
or U15526 (N_15526,N_15461,N_15304);
xor U15527 (N_15527,N_15391,N_15459);
xnor U15528 (N_15528,N_15001,N_15088);
nor U15529 (N_15529,N_15390,N_15019);
or U15530 (N_15530,N_15173,N_15227);
nor U15531 (N_15531,N_15048,N_15105);
and U15532 (N_15532,N_15398,N_15155);
xnor U15533 (N_15533,N_15126,N_15101);
nand U15534 (N_15534,N_15275,N_15022);
nand U15535 (N_15535,N_15410,N_15211);
nor U15536 (N_15536,N_15265,N_15058);
nand U15537 (N_15537,N_15213,N_15047);
nor U15538 (N_15538,N_15212,N_15277);
or U15539 (N_15539,N_15150,N_15070);
and U15540 (N_15540,N_15130,N_15157);
nand U15541 (N_15541,N_15317,N_15284);
or U15542 (N_15542,N_15355,N_15445);
nand U15543 (N_15543,N_15422,N_15146);
xor U15544 (N_15544,N_15242,N_15326);
and U15545 (N_15545,N_15283,N_15362);
xor U15546 (N_15546,N_15111,N_15159);
or U15547 (N_15547,N_15321,N_15318);
or U15548 (N_15548,N_15367,N_15383);
nor U15549 (N_15549,N_15399,N_15219);
nor U15550 (N_15550,N_15380,N_15018);
xor U15551 (N_15551,N_15426,N_15360);
nand U15552 (N_15552,N_15258,N_15247);
and U15553 (N_15553,N_15125,N_15076);
or U15554 (N_15554,N_15216,N_15440);
or U15555 (N_15555,N_15214,N_15385);
xnor U15556 (N_15556,N_15132,N_15210);
nand U15557 (N_15557,N_15457,N_15306);
and U15558 (N_15558,N_15189,N_15004);
and U15559 (N_15559,N_15151,N_15148);
nor U15560 (N_15560,N_15122,N_15300);
or U15561 (N_15561,N_15201,N_15128);
and U15562 (N_15562,N_15338,N_15016);
nor U15563 (N_15563,N_15167,N_15010);
or U15564 (N_15564,N_15480,N_15494);
or U15565 (N_15565,N_15424,N_15261);
or U15566 (N_15566,N_15456,N_15449);
xor U15567 (N_15567,N_15202,N_15307);
xnor U15568 (N_15568,N_15137,N_15477);
or U15569 (N_15569,N_15345,N_15439);
and U15570 (N_15570,N_15443,N_15066);
nor U15571 (N_15571,N_15107,N_15086);
nand U15572 (N_15572,N_15286,N_15182);
or U15573 (N_15573,N_15073,N_15053);
or U15574 (N_15574,N_15365,N_15147);
xor U15575 (N_15575,N_15329,N_15327);
nand U15576 (N_15576,N_15181,N_15093);
or U15577 (N_15577,N_15255,N_15206);
nor U15578 (N_15578,N_15092,N_15463);
nor U15579 (N_15579,N_15400,N_15428);
and U15580 (N_15580,N_15320,N_15425);
and U15581 (N_15581,N_15185,N_15199);
nor U15582 (N_15582,N_15045,N_15143);
nor U15583 (N_15583,N_15171,N_15115);
or U15584 (N_15584,N_15444,N_15310);
nand U15585 (N_15585,N_15131,N_15042);
or U15586 (N_15586,N_15301,N_15295);
nand U15587 (N_15587,N_15003,N_15470);
nand U15588 (N_15588,N_15079,N_15149);
nor U15589 (N_15589,N_15026,N_15187);
xor U15590 (N_15590,N_15292,N_15351);
xnor U15591 (N_15591,N_15486,N_15489);
and U15592 (N_15592,N_15401,N_15176);
xor U15593 (N_15593,N_15288,N_15020);
xor U15594 (N_15594,N_15209,N_15334);
and U15595 (N_15595,N_15077,N_15336);
or U15596 (N_15596,N_15082,N_15160);
nor U15597 (N_15597,N_15040,N_15230);
or U15598 (N_15598,N_15184,N_15223);
nand U15599 (N_15599,N_15027,N_15029);
or U15600 (N_15600,N_15376,N_15084);
or U15601 (N_15601,N_15472,N_15281);
nor U15602 (N_15602,N_15054,N_15423);
nor U15603 (N_15603,N_15005,N_15134);
or U15604 (N_15604,N_15237,N_15441);
or U15605 (N_15605,N_15475,N_15303);
xnor U15606 (N_15606,N_15110,N_15233);
xor U15607 (N_15607,N_15348,N_15080);
or U15608 (N_15608,N_15437,N_15235);
and U15609 (N_15609,N_15413,N_15013);
xor U15610 (N_15610,N_15190,N_15166);
nor U15611 (N_15611,N_15386,N_15169);
xnor U15612 (N_15612,N_15431,N_15144);
nor U15613 (N_15613,N_15200,N_15259);
xnor U15614 (N_15614,N_15344,N_15314);
nor U15615 (N_15615,N_15299,N_15118);
xnor U15616 (N_15616,N_15282,N_15468);
or U15617 (N_15617,N_15007,N_15361);
and U15618 (N_15618,N_15442,N_15384);
and U15619 (N_15619,N_15389,N_15488);
nor U15620 (N_15620,N_15256,N_15059);
xnor U15621 (N_15621,N_15085,N_15225);
or U15622 (N_15622,N_15438,N_15354);
or U15623 (N_15623,N_15096,N_15074);
or U15624 (N_15624,N_15158,N_15290);
or U15625 (N_15625,N_15394,N_15412);
and U15626 (N_15626,N_15240,N_15411);
or U15627 (N_15627,N_15363,N_15030);
and U15628 (N_15628,N_15094,N_15152);
and U15629 (N_15629,N_15451,N_15108);
nand U15630 (N_15630,N_15032,N_15381);
xor U15631 (N_15631,N_15083,N_15309);
nor U15632 (N_15632,N_15392,N_15249);
xnor U15633 (N_15633,N_15117,N_15239);
xnor U15634 (N_15634,N_15120,N_15232);
nor U15635 (N_15635,N_15081,N_15408);
nand U15636 (N_15636,N_15104,N_15174);
or U15637 (N_15637,N_15186,N_15287);
nor U15638 (N_15638,N_15378,N_15238);
nand U15639 (N_15639,N_15197,N_15496);
or U15640 (N_15640,N_15397,N_15373);
nor U15641 (N_15641,N_15460,N_15406);
or U15642 (N_15642,N_15476,N_15006);
nand U15643 (N_15643,N_15121,N_15331);
nor U15644 (N_15644,N_15098,N_15285);
xor U15645 (N_15645,N_15231,N_15067);
nor U15646 (N_15646,N_15293,N_15395);
or U15647 (N_15647,N_15091,N_15436);
xnor U15648 (N_15648,N_15485,N_15154);
and U15649 (N_15649,N_15127,N_15271);
or U15650 (N_15650,N_15244,N_15313);
nor U15651 (N_15651,N_15497,N_15356);
nor U15652 (N_15652,N_15183,N_15087);
nor U15653 (N_15653,N_15462,N_15435);
xor U15654 (N_15654,N_15332,N_15490);
xnor U15655 (N_15655,N_15162,N_15023);
nor U15656 (N_15656,N_15372,N_15419);
and U15657 (N_15657,N_15165,N_15450);
or U15658 (N_15658,N_15382,N_15266);
and U15659 (N_15659,N_15430,N_15498);
xor U15660 (N_15660,N_15052,N_15141);
xnor U15661 (N_15661,N_15368,N_15308);
nand U15662 (N_15662,N_15036,N_15370);
or U15663 (N_15663,N_15208,N_15139);
or U15664 (N_15664,N_15116,N_15388);
xor U15665 (N_15665,N_15017,N_15323);
or U15666 (N_15666,N_15038,N_15254);
or U15667 (N_15667,N_15467,N_15124);
nor U15668 (N_15668,N_15234,N_15015);
nor U15669 (N_15669,N_15479,N_15218);
xnor U15670 (N_15670,N_15222,N_15056);
or U15671 (N_15671,N_15434,N_15260);
nor U15672 (N_15672,N_15068,N_15033);
xnor U15673 (N_15673,N_15224,N_15371);
and U15674 (N_15674,N_15335,N_15057);
nor U15675 (N_15675,N_15416,N_15262);
nor U15676 (N_15676,N_15481,N_15156);
nor U15677 (N_15677,N_15474,N_15387);
nor U15678 (N_15678,N_15192,N_15180);
and U15679 (N_15679,N_15191,N_15102);
xor U15680 (N_15680,N_15178,N_15417);
nor U15681 (N_15681,N_15478,N_15458);
nand U15682 (N_15682,N_15236,N_15253);
and U15683 (N_15683,N_15312,N_15204);
nor U15684 (N_15684,N_15071,N_15049);
and U15685 (N_15685,N_15366,N_15168);
nor U15686 (N_15686,N_15353,N_15269);
nand U15687 (N_15687,N_15278,N_15175);
and U15688 (N_15688,N_15433,N_15369);
xnor U15689 (N_15689,N_15043,N_15100);
nor U15690 (N_15690,N_15455,N_15349);
or U15691 (N_15691,N_15316,N_15008);
and U15692 (N_15692,N_15044,N_15393);
or U15693 (N_15693,N_15464,N_15099);
xnor U15694 (N_15694,N_15055,N_15465);
nand U15695 (N_15695,N_15379,N_15446);
nand U15696 (N_15696,N_15346,N_15324);
or U15697 (N_15697,N_15357,N_15025);
nor U15698 (N_15698,N_15089,N_15095);
xnor U15699 (N_15699,N_15302,N_15403);
and U15700 (N_15700,N_15179,N_15409);
nand U15701 (N_15701,N_15297,N_15251);
nand U15702 (N_15702,N_15136,N_15339);
or U15703 (N_15703,N_15447,N_15414);
xnor U15704 (N_15704,N_15245,N_15163);
or U15705 (N_15705,N_15337,N_15289);
xnor U15706 (N_15706,N_15374,N_15452);
nor U15707 (N_15707,N_15483,N_15028);
xor U15708 (N_15708,N_15069,N_15311);
or U15709 (N_15709,N_15243,N_15375);
or U15710 (N_15710,N_15343,N_15203);
nor U15711 (N_15711,N_15135,N_15341);
nor U15712 (N_15712,N_15075,N_15333);
xor U15713 (N_15713,N_15220,N_15161);
nand U15714 (N_15714,N_15325,N_15198);
nor U15715 (N_15715,N_15448,N_15072);
xor U15716 (N_15716,N_15226,N_15432);
nor U15717 (N_15717,N_15241,N_15499);
xnor U15718 (N_15718,N_15035,N_15279);
nand U15719 (N_15719,N_15250,N_15119);
and U15720 (N_15720,N_15402,N_15164);
xor U15721 (N_15721,N_15207,N_15484);
nor U15722 (N_15722,N_15229,N_15473);
nor U15723 (N_15723,N_15377,N_15263);
xnor U15724 (N_15724,N_15315,N_15097);
nor U15725 (N_15725,N_15170,N_15273);
xnor U15726 (N_15726,N_15276,N_15352);
nor U15727 (N_15727,N_15064,N_15106);
or U15728 (N_15728,N_15142,N_15340);
and U15729 (N_15729,N_15217,N_15188);
or U15730 (N_15730,N_15205,N_15133);
and U15731 (N_15731,N_15469,N_15050);
and U15732 (N_15732,N_15041,N_15034);
nor U15733 (N_15733,N_15177,N_15051);
and U15734 (N_15734,N_15138,N_15418);
and U15735 (N_15735,N_15471,N_15011);
nand U15736 (N_15736,N_15328,N_15466);
nor U15737 (N_15737,N_15021,N_15014);
and U15738 (N_15738,N_15103,N_15060);
nor U15739 (N_15739,N_15487,N_15061);
xnor U15740 (N_15740,N_15000,N_15062);
or U15741 (N_15741,N_15153,N_15195);
nor U15742 (N_15742,N_15454,N_15453);
nand U15743 (N_15743,N_15090,N_15298);
nor U15744 (N_15744,N_15280,N_15252);
and U15745 (N_15745,N_15359,N_15129);
xnor U15746 (N_15746,N_15228,N_15270);
or U15747 (N_15747,N_15396,N_15347);
and U15748 (N_15748,N_15330,N_15193);
or U15749 (N_15749,N_15221,N_15002);
xnor U15750 (N_15750,N_15454,N_15320);
xnor U15751 (N_15751,N_15193,N_15189);
nor U15752 (N_15752,N_15076,N_15238);
nand U15753 (N_15753,N_15493,N_15131);
and U15754 (N_15754,N_15056,N_15137);
nor U15755 (N_15755,N_15305,N_15325);
and U15756 (N_15756,N_15183,N_15224);
or U15757 (N_15757,N_15416,N_15434);
xnor U15758 (N_15758,N_15320,N_15361);
xor U15759 (N_15759,N_15384,N_15387);
and U15760 (N_15760,N_15142,N_15443);
xor U15761 (N_15761,N_15077,N_15295);
and U15762 (N_15762,N_15126,N_15453);
nor U15763 (N_15763,N_15320,N_15351);
xor U15764 (N_15764,N_15365,N_15210);
xnor U15765 (N_15765,N_15290,N_15143);
and U15766 (N_15766,N_15456,N_15376);
and U15767 (N_15767,N_15113,N_15096);
or U15768 (N_15768,N_15414,N_15448);
nor U15769 (N_15769,N_15202,N_15462);
or U15770 (N_15770,N_15336,N_15098);
nor U15771 (N_15771,N_15410,N_15166);
or U15772 (N_15772,N_15289,N_15346);
nor U15773 (N_15773,N_15224,N_15109);
and U15774 (N_15774,N_15415,N_15410);
or U15775 (N_15775,N_15289,N_15396);
xnor U15776 (N_15776,N_15293,N_15400);
nand U15777 (N_15777,N_15320,N_15445);
nand U15778 (N_15778,N_15013,N_15479);
nor U15779 (N_15779,N_15199,N_15382);
nor U15780 (N_15780,N_15209,N_15149);
and U15781 (N_15781,N_15339,N_15412);
nor U15782 (N_15782,N_15200,N_15068);
nor U15783 (N_15783,N_15335,N_15065);
nand U15784 (N_15784,N_15158,N_15219);
nand U15785 (N_15785,N_15359,N_15164);
and U15786 (N_15786,N_15096,N_15176);
and U15787 (N_15787,N_15063,N_15170);
xnor U15788 (N_15788,N_15312,N_15457);
nor U15789 (N_15789,N_15184,N_15194);
nand U15790 (N_15790,N_15053,N_15203);
or U15791 (N_15791,N_15290,N_15212);
nor U15792 (N_15792,N_15356,N_15015);
xnor U15793 (N_15793,N_15328,N_15490);
or U15794 (N_15794,N_15133,N_15070);
and U15795 (N_15795,N_15342,N_15086);
nor U15796 (N_15796,N_15020,N_15106);
nor U15797 (N_15797,N_15238,N_15256);
nand U15798 (N_15798,N_15350,N_15192);
nand U15799 (N_15799,N_15401,N_15216);
nand U15800 (N_15800,N_15490,N_15290);
and U15801 (N_15801,N_15086,N_15406);
or U15802 (N_15802,N_15388,N_15435);
xnor U15803 (N_15803,N_15497,N_15286);
or U15804 (N_15804,N_15012,N_15118);
nor U15805 (N_15805,N_15281,N_15100);
nor U15806 (N_15806,N_15429,N_15468);
nor U15807 (N_15807,N_15427,N_15444);
and U15808 (N_15808,N_15196,N_15272);
and U15809 (N_15809,N_15310,N_15129);
nand U15810 (N_15810,N_15273,N_15496);
nor U15811 (N_15811,N_15380,N_15196);
and U15812 (N_15812,N_15140,N_15019);
nand U15813 (N_15813,N_15046,N_15457);
nor U15814 (N_15814,N_15046,N_15438);
nor U15815 (N_15815,N_15419,N_15352);
nor U15816 (N_15816,N_15401,N_15465);
or U15817 (N_15817,N_15221,N_15032);
or U15818 (N_15818,N_15413,N_15141);
nand U15819 (N_15819,N_15478,N_15033);
or U15820 (N_15820,N_15261,N_15224);
or U15821 (N_15821,N_15072,N_15283);
or U15822 (N_15822,N_15341,N_15186);
nand U15823 (N_15823,N_15048,N_15023);
or U15824 (N_15824,N_15358,N_15073);
nand U15825 (N_15825,N_15131,N_15225);
nor U15826 (N_15826,N_15460,N_15334);
xnor U15827 (N_15827,N_15368,N_15145);
and U15828 (N_15828,N_15440,N_15162);
nor U15829 (N_15829,N_15079,N_15090);
nand U15830 (N_15830,N_15413,N_15062);
or U15831 (N_15831,N_15152,N_15366);
nand U15832 (N_15832,N_15106,N_15138);
nor U15833 (N_15833,N_15497,N_15059);
xnor U15834 (N_15834,N_15091,N_15133);
xor U15835 (N_15835,N_15173,N_15239);
or U15836 (N_15836,N_15051,N_15211);
and U15837 (N_15837,N_15368,N_15126);
nand U15838 (N_15838,N_15450,N_15030);
or U15839 (N_15839,N_15374,N_15330);
nor U15840 (N_15840,N_15491,N_15000);
xnor U15841 (N_15841,N_15353,N_15187);
and U15842 (N_15842,N_15396,N_15485);
or U15843 (N_15843,N_15494,N_15387);
nor U15844 (N_15844,N_15374,N_15041);
or U15845 (N_15845,N_15306,N_15150);
nand U15846 (N_15846,N_15119,N_15111);
xor U15847 (N_15847,N_15237,N_15072);
xor U15848 (N_15848,N_15350,N_15395);
nand U15849 (N_15849,N_15234,N_15323);
xor U15850 (N_15850,N_15174,N_15219);
nand U15851 (N_15851,N_15420,N_15251);
xor U15852 (N_15852,N_15356,N_15265);
and U15853 (N_15853,N_15005,N_15184);
nor U15854 (N_15854,N_15450,N_15092);
xnor U15855 (N_15855,N_15248,N_15470);
nand U15856 (N_15856,N_15095,N_15034);
nor U15857 (N_15857,N_15158,N_15478);
and U15858 (N_15858,N_15232,N_15033);
nand U15859 (N_15859,N_15450,N_15020);
or U15860 (N_15860,N_15415,N_15255);
or U15861 (N_15861,N_15492,N_15377);
and U15862 (N_15862,N_15166,N_15145);
nand U15863 (N_15863,N_15038,N_15289);
or U15864 (N_15864,N_15025,N_15245);
or U15865 (N_15865,N_15224,N_15191);
and U15866 (N_15866,N_15422,N_15358);
nand U15867 (N_15867,N_15358,N_15360);
and U15868 (N_15868,N_15189,N_15345);
nand U15869 (N_15869,N_15336,N_15327);
or U15870 (N_15870,N_15406,N_15204);
and U15871 (N_15871,N_15310,N_15219);
nor U15872 (N_15872,N_15105,N_15323);
xor U15873 (N_15873,N_15447,N_15010);
nor U15874 (N_15874,N_15032,N_15465);
xor U15875 (N_15875,N_15449,N_15030);
or U15876 (N_15876,N_15159,N_15041);
and U15877 (N_15877,N_15063,N_15278);
or U15878 (N_15878,N_15115,N_15108);
nand U15879 (N_15879,N_15429,N_15129);
or U15880 (N_15880,N_15415,N_15115);
nand U15881 (N_15881,N_15475,N_15272);
xor U15882 (N_15882,N_15218,N_15162);
xnor U15883 (N_15883,N_15004,N_15361);
or U15884 (N_15884,N_15268,N_15230);
nand U15885 (N_15885,N_15295,N_15209);
nand U15886 (N_15886,N_15137,N_15383);
xnor U15887 (N_15887,N_15317,N_15156);
and U15888 (N_15888,N_15187,N_15256);
xnor U15889 (N_15889,N_15410,N_15103);
xnor U15890 (N_15890,N_15445,N_15153);
and U15891 (N_15891,N_15209,N_15038);
nor U15892 (N_15892,N_15344,N_15363);
nor U15893 (N_15893,N_15473,N_15224);
xnor U15894 (N_15894,N_15309,N_15247);
or U15895 (N_15895,N_15095,N_15062);
or U15896 (N_15896,N_15388,N_15231);
xnor U15897 (N_15897,N_15023,N_15139);
nand U15898 (N_15898,N_15484,N_15462);
xnor U15899 (N_15899,N_15031,N_15336);
and U15900 (N_15900,N_15237,N_15052);
xnor U15901 (N_15901,N_15373,N_15457);
or U15902 (N_15902,N_15333,N_15220);
nor U15903 (N_15903,N_15320,N_15095);
and U15904 (N_15904,N_15235,N_15166);
xor U15905 (N_15905,N_15191,N_15040);
or U15906 (N_15906,N_15179,N_15086);
nand U15907 (N_15907,N_15190,N_15398);
nand U15908 (N_15908,N_15007,N_15207);
and U15909 (N_15909,N_15380,N_15470);
nor U15910 (N_15910,N_15095,N_15149);
and U15911 (N_15911,N_15440,N_15374);
nand U15912 (N_15912,N_15466,N_15166);
nor U15913 (N_15913,N_15264,N_15343);
nand U15914 (N_15914,N_15062,N_15447);
or U15915 (N_15915,N_15334,N_15044);
xor U15916 (N_15916,N_15240,N_15285);
or U15917 (N_15917,N_15447,N_15448);
and U15918 (N_15918,N_15120,N_15038);
or U15919 (N_15919,N_15424,N_15415);
or U15920 (N_15920,N_15497,N_15204);
or U15921 (N_15921,N_15387,N_15018);
xor U15922 (N_15922,N_15288,N_15450);
and U15923 (N_15923,N_15055,N_15062);
or U15924 (N_15924,N_15126,N_15046);
nand U15925 (N_15925,N_15116,N_15342);
nor U15926 (N_15926,N_15030,N_15361);
or U15927 (N_15927,N_15069,N_15078);
or U15928 (N_15928,N_15152,N_15265);
nand U15929 (N_15929,N_15403,N_15169);
nand U15930 (N_15930,N_15162,N_15435);
and U15931 (N_15931,N_15467,N_15477);
and U15932 (N_15932,N_15049,N_15080);
nor U15933 (N_15933,N_15108,N_15135);
xor U15934 (N_15934,N_15088,N_15077);
nor U15935 (N_15935,N_15409,N_15336);
xor U15936 (N_15936,N_15202,N_15461);
and U15937 (N_15937,N_15429,N_15006);
and U15938 (N_15938,N_15064,N_15045);
and U15939 (N_15939,N_15243,N_15191);
xor U15940 (N_15940,N_15264,N_15099);
or U15941 (N_15941,N_15472,N_15271);
or U15942 (N_15942,N_15385,N_15158);
nor U15943 (N_15943,N_15204,N_15445);
nor U15944 (N_15944,N_15166,N_15388);
or U15945 (N_15945,N_15174,N_15208);
nor U15946 (N_15946,N_15042,N_15002);
nor U15947 (N_15947,N_15314,N_15030);
or U15948 (N_15948,N_15152,N_15463);
and U15949 (N_15949,N_15221,N_15425);
xor U15950 (N_15950,N_15374,N_15469);
nor U15951 (N_15951,N_15101,N_15196);
nand U15952 (N_15952,N_15401,N_15324);
nand U15953 (N_15953,N_15283,N_15497);
and U15954 (N_15954,N_15326,N_15205);
or U15955 (N_15955,N_15406,N_15015);
and U15956 (N_15956,N_15005,N_15116);
nor U15957 (N_15957,N_15484,N_15273);
and U15958 (N_15958,N_15300,N_15218);
or U15959 (N_15959,N_15190,N_15140);
or U15960 (N_15960,N_15406,N_15057);
or U15961 (N_15961,N_15110,N_15311);
xor U15962 (N_15962,N_15267,N_15303);
or U15963 (N_15963,N_15420,N_15237);
and U15964 (N_15964,N_15086,N_15106);
nor U15965 (N_15965,N_15066,N_15135);
or U15966 (N_15966,N_15459,N_15446);
or U15967 (N_15967,N_15178,N_15293);
and U15968 (N_15968,N_15288,N_15331);
xor U15969 (N_15969,N_15109,N_15084);
or U15970 (N_15970,N_15346,N_15081);
nand U15971 (N_15971,N_15162,N_15357);
nor U15972 (N_15972,N_15444,N_15205);
nor U15973 (N_15973,N_15238,N_15244);
or U15974 (N_15974,N_15243,N_15091);
and U15975 (N_15975,N_15337,N_15312);
or U15976 (N_15976,N_15301,N_15428);
or U15977 (N_15977,N_15267,N_15205);
nand U15978 (N_15978,N_15001,N_15338);
nand U15979 (N_15979,N_15074,N_15310);
xor U15980 (N_15980,N_15108,N_15068);
xor U15981 (N_15981,N_15333,N_15178);
nor U15982 (N_15982,N_15161,N_15448);
nor U15983 (N_15983,N_15314,N_15299);
nor U15984 (N_15984,N_15476,N_15470);
nand U15985 (N_15985,N_15251,N_15397);
xor U15986 (N_15986,N_15037,N_15389);
nor U15987 (N_15987,N_15210,N_15056);
nor U15988 (N_15988,N_15476,N_15129);
or U15989 (N_15989,N_15148,N_15087);
xnor U15990 (N_15990,N_15083,N_15310);
nand U15991 (N_15991,N_15131,N_15445);
xor U15992 (N_15992,N_15470,N_15113);
nand U15993 (N_15993,N_15084,N_15244);
nand U15994 (N_15994,N_15069,N_15219);
xnor U15995 (N_15995,N_15184,N_15471);
nor U15996 (N_15996,N_15071,N_15199);
and U15997 (N_15997,N_15228,N_15229);
xor U15998 (N_15998,N_15177,N_15409);
nand U15999 (N_15999,N_15458,N_15260);
and U16000 (N_16000,N_15559,N_15746);
and U16001 (N_16001,N_15954,N_15884);
xnor U16002 (N_16002,N_15546,N_15531);
nor U16003 (N_16003,N_15990,N_15805);
and U16004 (N_16004,N_15636,N_15569);
xnor U16005 (N_16005,N_15796,N_15577);
xor U16006 (N_16006,N_15725,N_15873);
nor U16007 (N_16007,N_15795,N_15517);
nor U16008 (N_16008,N_15631,N_15993);
nor U16009 (N_16009,N_15637,N_15629);
xor U16010 (N_16010,N_15513,N_15509);
nor U16011 (N_16011,N_15832,N_15802);
or U16012 (N_16012,N_15789,N_15558);
nor U16013 (N_16013,N_15890,N_15861);
nand U16014 (N_16014,N_15753,N_15868);
nand U16015 (N_16015,N_15682,N_15843);
nand U16016 (N_16016,N_15688,N_15984);
and U16017 (N_16017,N_15889,N_15625);
and U16018 (N_16018,N_15968,N_15800);
xnor U16019 (N_16019,N_15952,N_15925);
or U16020 (N_16020,N_15595,N_15827);
nand U16021 (N_16021,N_15582,N_15869);
xor U16022 (N_16022,N_15891,N_15865);
and U16023 (N_16023,N_15914,N_15886);
nor U16024 (N_16024,N_15912,N_15689);
xnor U16025 (N_16025,N_15534,N_15609);
xor U16026 (N_16026,N_15537,N_15812);
and U16027 (N_16027,N_15672,N_15542);
or U16028 (N_16028,N_15634,N_15658);
or U16029 (N_16029,N_15982,N_15573);
nor U16030 (N_16030,N_15944,N_15511);
xor U16031 (N_16031,N_15960,N_15806);
and U16032 (N_16032,N_15817,N_15823);
and U16033 (N_16033,N_15966,N_15856);
or U16034 (N_16034,N_15848,N_15878);
xnor U16035 (N_16035,N_15696,N_15600);
xor U16036 (N_16036,N_15521,N_15854);
nor U16037 (N_16037,N_15719,N_15663);
nand U16038 (N_16038,N_15533,N_15695);
nor U16039 (N_16039,N_15557,N_15726);
nand U16040 (N_16040,N_15583,N_15524);
or U16041 (N_16041,N_15760,N_15662);
xnor U16042 (N_16042,N_15505,N_15586);
nor U16043 (N_16043,N_15602,N_15681);
or U16044 (N_16044,N_15840,N_15700);
nand U16045 (N_16045,N_15540,N_15530);
xnor U16046 (N_16046,N_15860,N_15736);
nand U16047 (N_16047,N_15526,N_15617);
and U16048 (N_16048,N_15971,N_15642);
nand U16049 (N_16049,N_15898,N_15776);
or U16050 (N_16050,N_15942,N_15846);
nand U16051 (N_16051,N_15774,N_15626);
or U16052 (N_16052,N_15815,N_15938);
or U16053 (N_16053,N_15959,N_15732);
nor U16054 (N_16054,N_15887,N_15562);
and U16055 (N_16055,N_15734,N_15677);
nor U16056 (N_16056,N_15826,N_15633);
or U16057 (N_16057,N_15824,N_15568);
xnor U16058 (N_16058,N_15702,N_15855);
and U16059 (N_16059,N_15527,N_15933);
nand U16060 (N_16060,N_15772,N_15989);
nor U16061 (N_16061,N_15581,N_15980);
and U16062 (N_16062,N_15652,N_15893);
xnor U16063 (N_16063,N_15644,N_15782);
or U16064 (N_16064,N_15769,N_15512);
xnor U16065 (N_16065,N_15956,N_15588);
or U16066 (N_16066,N_15948,N_15991);
xnor U16067 (N_16067,N_15838,N_15999);
and U16068 (N_16068,N_15563,N_15572);
or U16069 (N_16069,N_15678,N_15836);
nor U16070 (N_16070,N_15913,N_15766);
and U16071 (N_16071,N_15937,N_15754);
or U16072 (N_16072,N_15945,N_15941);
xor U16073 (N_16073,N_15804,N_15510);
and U16074 (N_16074,N_15685,N_15750);
nand U16075 (N_16075,N_15965,N_15833);
nand U16076 (N_16076,N_15645,N_15679);
xnor U16077 (N_16077,N_15829,N_15545);
and U16078 (N_16078,N_15523,N_15738);
xor U16079 (N_16079,N_15741,N_15798);
nor U16080 (N_16080,N_15905,N_15541);
nor U16081 (N_16081,N_15946,N_15713);
and U16082 (N_16082,N_15538,N_15601);
xnor U16083 (N_16083,N_15655,N_15716);
or U16084 (N_16084,N_15867,N_15503);
and U16085 (N_16085,N_15651,N_15504);
and U16086 (N_16086,N_15718,N_15668);
nand U16087 (N_16087,N_15666,N_15697);
xnor U16088 (N_16088,N_15618,N_15904);
xnor U16089 (N_16089,N_15686,N_15759);
or U16090 (N_16090,N_15529,N_15711);
xnor U16091 (N_16091,N_15687,N_15632);
and U16092 (N_16092,N_15790,N_15923);
xnor U16093 (N_16093,N_15995,N_15849);
and U16094 (N_16094,N_15751,N_15997);
nor U16095 (N_16095,N_15698,N_15724);
nor U16096 (N_16096,N_15828,N_15731);
or U16097 (N_16097,N_15680,N_15947);
and U16098 (N_16098,N_15596,N_15566);
nand U16099 (N_16099,N_15797,N_15972);
and U16100 (N_16100,N_15811,N_15575);
and U16101 (N_16101,N_15919,N_15837);
nor U16102 (N_16102,N_15799,N_15665);
nor U16103 (N_16103,N_15974,N_15901);
nor U16104 (N_16104,N_15996,N_15684);
and U16105 (N_16105,N_15727,N_15528);
and U16106 (N_16106,N_15770,N_15940);
or U16107 (N_16107,N_15756,N_15957);
nand U16108 (N_16108,N_15788,N_15951);
and U16109 (N_16109,N_15821,N_15987);
nand U16110 (N_16110,N_15561,N_15714);
or U16111 (N_16111,N_15851,N_15585);
xor U16112 (N_16112,N_15871,N_15749);
or U16113 (N_16113,N_15640,N_15660);
and U16114 (N_16114,N_15560,N_15519);
nand U16115 (N_16115,N_15794,N_15844);
nand U16116 (N_16116,N_15622,N_15742);
and U16117 (N_16117,N_15525,N_15858);
xnor U16118 (N_16118,N_15842,N_15669);
xnor U16119 (N_16119,N_15579,N_15692);
or U16120 (N_16120,N_15608,N_15780);
nand U16121 (N_16121,N_15864,N_15648);
xnor U16122 (N_16122,N_15615,N_15639);
nor U16123 (N_16123,N_15986,N_15721);
nand U16124 (N_16124,N_15978,N_15690);
nand U16125 (N_16125,N_15894,N_15704);
nor U16126 (N_16126,N_15584,N_15627);
or U16127 (N_16127,N_15612,N_15535);
xor U16128 (N_16128,N_15786,N_15973);
xor U16129 (N_16129,N_15740,N_15853);
and U16130 (N_16130,N_15703,N_15981);
and U16131 (N_16131,N_15675,N_15730);
nor U16132 (N_16132,N_15603,N_15580);
and U16133 (N_16133,N_15723,N_15813);
nand U16134 (N_16134,N_15939,N_15735);
and U16135 (N_16135,N_15863,N_15808);
and U16136 (N_16136,N_15880,N_15623);
or U16137 (N_16137,N_15587,N_15818);
or U16138 (N_16138,N_15928,N_15653);
or U16139 (N_16139,N_15908,N_15694);
nand U16140 (N_16140,N_15915,N_15881);
and U16141 (N_16141,N_15775,N_15641);
xnor U16142 (N_16142,N_15619,N_15819);
or U16143 (N_16143,N_15847,N_15816);
xnor U16144 (N_16144,N_15969,N_15879);
xnor U16145 (N_16145,N_15547,N_15850);
or U16146 (N_16146,N_15934,N_15988);
xnor U16147 (N_16147,N_15606,N_15520);
nand U16148 (N_16148,N_15656,N_15610);
nor U16149 (N_16149,N_15709,N_15729);
or U16150 (N_16150,N_15551,N_15657);
or U16151 (N_16151,N_15773,N_15779);
or U16152 (N_16152,N_15825,N_15571);
xnor U16153 (N_16153,N_15752,N_15717);
xnor U16154 (N_16154,N_15565,N_15744);
and U16155 (N_16155,N_15638,N_15930);
nor U16156 (N_16156,N_15907,N_15674);
xor U16157 (N_16157,N_15883,N_15768);
nor U16158 (N_16158,N_15983,N_15543);
or U16159 (N_16159,N_15892,N_15979);
nor U16160 (N_16160,N_15567,N_15916);
nand U16161 (N_16161,N_15593,N_15548);
and U16162 (N_16162,N_15500,N_15589);
nor U16163 (N_16163,N_15624,N_15874);
nand U16164 (N_16164,N_15594,N_15918);
or U16165 (N_16165,N_15943,N_15955);
nand U16166 (N_16166,N_15607,N_15970);
and U16167 (N_16167,N_15683,N_15616);
or U16168 (N_16168,N_15807,N_15791);
nand U16169 (N_16169,N_15862,N_15762);
and U16170 (N_16170,N_15781,N_15708);
nor U16171 (N_16171,N_15764,N_15936);
and U16172 (N_16172,N_15699,N_15508);
nand U16173 (N_16173,N_15720,N_15733);
nand U16174 (N_16174,N_15920,N_15778);
nor U16175 (N_16175,N_15630,N_15924);
or U16176 (N_16176,N_15613,N_15872);
and U16177 (N_16177,N_15755,N_15643);
or U16178 (N_16178,N_15536,N_15705);
or U16179 (N_16179,N_15897,N_15701);
or U16180 (N_16180,N_15831,N_15953);
and U16181 (N_16181,N_15830,N_15555);
xnor U16182 (N_16182,N_15992,N_15591);
xor U16183 (N_16183,N_15516,N_15757);
and U16184 (N_16184,N_15932,N_15809);
nand U16185 (N_16185,N_15654,N_15590);
or U16186 (N_16186,N_15927,N_15877);
nand U16187 (N_16187,N_15964,N_15673);
nor U16188 (N_16188,N_15985,N_15765);
xnor U16189 (N_16189,N_15650,N_15539);
nand U16190 (N_16190,N_15635,N_15707);
nor U16191 (N_16191,N_15949,N_15605);
or U16192 (N_16192,N_15801,N_15906);
nor U16193 (N_16193,N_15552,N_15659);
nor U16194 (N_16194,N_15564,N_15739);
xnor U16195 (N_16195,N_15763,N_15922);
nor U16196 (N_16196,N_15870,N_15506);
nor U16197 (N_16197,N_15921,N_15777);
nand U16198 (N_16198,N_15611,N_15646);
xor U16199 (N_16199,N_15670,N_15761);
xnor U16200 (N_16200,N_15522,N_15785);
xor U16201 (N_16201,N_15554,N_15614);
xor U16202 (N_16202,N_15574,N_15661);
nor U16203 (N_16203,N_15822,N_15501);
nand U16204 (N_16204,N_15747,N_15866);
nor U16205 (N_16205,N_15803,N_15628);
or U16206 (N_16206,N_15647,N_15621);
and U16207 (N_16207,N_15792,N_15793);
xor U16208 (N_16208,N_15758,N_15706);
xor U16209 (N_16209,N_15902,N_15620);
nor U16210 (N_16210,N_15814,N_15909);
and U16211 (N_16211,N_15578,N_15931);
nor U16212 (N_16212,N_15911,N_15876);
nand U16213 (N_16213,N_15903,N_15783);
nor U16214 (N_16214,N_15728,N_15929);
and U16215 (N_16215,N_15845,N_15745);
nor U16216 (N_16216,N_15570,N_15507);
xor U16217 (N_16217,N_15691,N_15502);
xnor U16218 (N_16218,N_15532,N_15715);
and U16219 (N_16219,N_15839,N_15841);
or U16220 (N_16220,N_15693,N_15671);
or U16221 (N_16221,N_15958,N_15676);
xnor U16222 (N_16222,N_15599,N_15515);
and U16223 (N_16223,N_15664,N_15899);
or U16224 (N_16224,N_15976,N_15712);
and U16225 (N_16225,N_15962,N_15885);
nor U16226 (N_16226,N_15592,N_15859);
nor U16227 (N_16227,N_15820,N_15998);
or U16228 (N_16228,N_15710,N_15888);
and U16229 (N_16229,N_15722,N_15784);
xnor U16230 (N_16230,N_15748,N_15935);
nand U16231 (N_16231,N_15649,N_15598);
nand U16232 (N_16232,N_15553,N_15994);
or U16233 (N_16233,N_15852,N_15544);
nand U16234 (N_16234,N_15834,N_15857);
nor U16235 (N_16235,N_15896,N_15576);
or U16236 (N_16236,N_15975,N_15743);
or U16237 (N_16237,N_15910,N_15549);
nand U16238 (N_16238,N_15963,N_15882);
or U16239 (N_16239,N_15667,N_15967);
xnor U16240 (N_16240,N_15926,N_15977);
nor U16241 (N_16241,N_15835,N_15556);
nor U16242 (N_16242,N_15597,N_15604);
and U16243 (N_16243,N_15810,N_15961);
nand U16244 (N_16244,N_15895,N_15518);
nand U16245 (N_16245,N_15737,N_15917);
nand U16246 (N_16246,N_15550,N_15950);
xor U16247 (N_16247,N_15767,N_15771);
xor U16248 (N_16248,N_15787,N_15900);
nor U16249 (N_16249,N_15875,N_15514);
xnor U16250 (N_16250,N_15834,N_15946);
nand U16251 (N_16251,N_15680,N_15502);
nor U16252 (N_16252,N_15761,N_15765);
nor U16253 (N_16253,N_15988,N_15551);
and U16254 (N_16254,N_15839,N_15618);
xor U16255 (N_16255,N_15721,N_15575);
nand U16256 (N_16256,N_15627,N_15937);
or U16257 (N_16257,N_15526,N_15580);
nor U16258 (N_16258,N_15679,N_15584);
and U16259 (N_16259,N_15635,N_15692);
xor U16260 (N_16260,N_15887,N_15742);
or U16261 (N_16261,N_15865,N_15875);
nand U16262 (N_16262,N_15659,N_15539);
nor U16263 (N_16263,N_15586,N_15943);
or U16264 (N_16264,N_15949,N_15946);
or U16265 (N_16265,N_15967,N_15550);
nand U16266 (N_16266,N_15516,N_15904);
nand U16267 (N_16267,N_15531,N_15595);
and U16268 (N_16268,N_15989,N_15774);
and U16269 (N_16269,N_15855,N_15693);
nor U16270 (N_16270,N_15888,N_15503);
nand U16271 (N_16271,N_15640,N_15562);
or U16272 (N_16272,N_15959,N_15664);
nand U16273 (N_16273,N_15837,N_15898);
nor U16274 (N_16274,N_15516,N_15533);
nor U16275 (N_16275,N_15918,N_15728);
xor U16276 (N_16276,N_15628,N_15855);
or U16277 (N_16277,N_15725,N_15736);
and U16278 (N_16278,N_15678,N_15509);
nor U16279 (N_16279,N_15600,N_15605);
nand U16280 (N_16280,N_15711,N_15536);
and U16281 (N_16281,N_15930,N_15945);
or U16282 (N_16282,N_15844,N_15608);
xor U16283 (N_16283,N_15681,N_15776);
and U16284 (N_16284,N_15878,N_15897);
or U16285 (N_16285,N_15676,N_15600);
xnor U16286 (N_16286,N_15736,N_15718);
or U16287 (N_16287,N_15965,N_15673);
xnor U16288 (N_16288,N_15830,N_15576);
nand U16289 (N_16289,N_15720,N_15559);
xor U16290 (N_16290,N_15605,N_15510);
or U16291 (N_16291,N_15809,N_15815);
or U16292 (N_16292,N_15776,N_15896);
nand U16293 (N_16293,N_15669,N_15504);
xnor U16294 (N_16294,N_15731,N_15513);
or U16295 (N_16295,N_15809,N_15713);
xor U16296 (N_16296,N_15859,N_15507);
nand U16297 (N_16297,N_15948,N_15759);
or U16298 (N_16298,N_15526,N_15509);
and U16299 (N_16299,N_15521,N_15892);
and U16300 (N_16300,N_15931,N_15536);
and U16301 (N_16301,N_15516,N_15811);
nand U16302 (N_16302,N_15858,N_15886);
nand U16303 (N_16303,N_15998,N_15794);
xnor U16304 (N_16304,N_15994,N_15862);
nor U16305 (N_16305,N_15888,N_15661);
nand U16306 (N_16306,N_15793,N_15962);
and U16307 (N_16307,N_15771,N_15790);
and U16308 (N_16308,N_15518,N_15710);
nand U16309 (N_16309,N_15567,N_15911);
and U16310 (N_16310,N_15673,N_15885);
xnor U16311 (N_16311,N_15889,N_15907);
nor U16312 (N_16312,N_15674,N_15946);
xnor U16313 (N_16313,N_15958,N_15760);
and U16314 (N_16314,N_15893,N_15574);
and U16315 (N_16315,N_15585,N_15641);
and U16316 (N_16316,N_15728,N_15958);
or U16317 (N_16317,N_15744,N_15667);
or U16318 (N_16318,N_15711,N_15808);
nor U16319 (N_16319,N_15788,N_15879);
xnor U16320 (N_16320,N_15638,N_15553);
nor U16321 (N_16321,N_15829,N_15657);
nand U16322 (N_16322,N_15560,N_15797);
xor U16323 (N_16323,N_15937,N_15580);
xor U16324 (N_16324,N_15850,N_15949);
and U16325 (N_16325,N_15750,N_15654);
and U16326 (N_16326,N_15773,N_15591);
xnor U16327 (N_16327,N_15742,N_15713);
nor U16328 (N_16328,N_15737,N_15818);
nor U16329 (N_16329,N_15734,N_15946);
nor U16330 (N_16330,N_15668,N_15958);
and U16331 (N_16331,N_15635,N_15903);
nor U16332 (N_16332,N_15613,N_15999);
nor U16333 (N_16333,N_15785,N_15720);
nor U16334 (N_16334,N_15566,N_15600);
nor U16335 (N_16335,N_15686,N_15705);
and U16336 (N_16336,N_15532,N_15632);
nand U16337 (N_16337,N_15551,N_15993);
nor U16338 (N_16338,N_15607,N_15766);
nor U16339 (N_16339,N_15511,N_15591);
or U16340 (N_16340,N_15515,N_15952);
or U16341 (N_16341,N_15815,N_15882);
nor U16342 (N_16342,N_15858,N_15801);
nand U16343 (N_16343,N_15869,N_15709);
xnor U16344 (N_16344,N_15835,N_15944);
nand U16345 (N_16345,N_15621,N_15685);
xnor U16346 (N_16346,N_15949,N_15794);
nor U16347 (N_16347,N_15784,N_15680);
and U16348 (N_16348,N_15517,N_15707);
xnor U16349 (N_16349,N_15648,N_15632);
or U16350 (N_16350,N_15727,N_15603);
or U16351 (N_16351,N_15722,N_15719);
or U16352 (N_16352,N_15714,N_15591);
or U16353 (N_16353,N_15516,N_15520);
nor U16354 (N_16354,N_15765,N_15530);
nand U16355 (N_16355,N_15850,N_15931);
xnor U16356 (N_16356,N_15867,N_15986);
or U16357 (N_16357,N_15864,N_15898);
and U16358 (N_16358,N_15947,N_15678);
nor U16359 (N_16359,N_15718,N_15618);
xnor U16360 (N_16360,N_15890,N_15880);
and U16361 (N_16361,N_15676,N_15694);
xor U16362 (N_16362,N_15535,N_15977);
or U16363 (N_16363,N_15725,N_15546);
or U16364 (N_16364,N_15930,N_15812);
xor U16365 (N_16365,N_15509,N_15762);
nor U16366 (N_16366,N_15999,N_15974);
and U16367 (N_16367,N_15709,N_15917);
or U16368 (N_16368,N_15713,N_15703);
xor U16369 (N_16369,N_15701,N_15963);
and U16370 (N_16370,N_15963,N_15985);
xor U16371 (N_16371,N_15913,N_15908);
xnor U16372 (N_16372,N_15789,N_15751);
and U16373 (N_16373,N_15930,N_15591);
and U16374 (N_16374,N_15528,N_15684);
xnor U16375 (N_16375,N_15916,N_15597);
xor U16376 (N_16376,N_15588,N_15600);
and U16377 (N_16377,N_15904,N_15684);
xnor U16378 (N_16378,N_15689,N_15727);
nor U16379 (N_16379,N_15914,N_15510);
and U16380 (N_16380,N_15619,N_15814);
nand U16381 (N_16381,N_15882,N_15673);
or U16382 (N_16382,N_15535,N_15570);
or U16383 (N_16383,N_15622,N_15568);
xor U16384 (N_16384,N_15802,N_15827);
nand U16385 (N_16385,N_15554,N_15963);
xor U16386 (N_16386,N_15513,N_15522);
or U16387 (N_16387,N_15742,N_15931);
nand U16388 (N_16388,N_15992,N_15921);
or U16389 (N_16389,N_15791,N_15689);
nand U16390 (N_16390,N_15765,N_15974);
nand U16391 (N_16391,N_15985,N_15611);
or U16392 (N_16392,N_15570,N_15575);
and U16393 (N_16393,N_15746,N_15856);
xnor U16394 (N_16394,N_15791,N_15790);
nor U16395 (N_16395,N_15525,N_15828);
and U16396 (N_16396,N_15696,N_15501);
nor U16397 (N_16397,N_15796,N_15992);
xor U16398 (N_16398,N_15795,N_15575);
and U16399 (N_16399,N_15893,N_15526);
and U16400 (N_16400,N_15586,N_15587);
nor U16401 (N_16401,N_15594,N_15940);
xor U16402 (N_16402,N_15588,N_15858);
nor U16403 (N_16403,N_15974,N_15937);
and U16404 (N_16404,N_15906,N_15972);
and U16405 (N_16405,N_15766,N_15877);
nand U16406 (N_16406,N_15744,N_15658);
xnor U16407 (N_16407,N_15624,N_15934);
xor U16408 (N_16408,N_15672,N_15893);
and U16409 (N_16409,N_15583,N_15945);
nor U16410 (N_16410,N_15710,N_15872);
or U16411 (N_16411,N_15750,N_15993);
xor U16412 (N_16412,N_15632,N_15986);
xor U16413 (N_16413,N_15747,N_15767);
xnor U16414 (N_16414,N_15526,N_15586);
xor U16415 (N_16415,N_15658,N_15725);
nor U16416 (N_16416,N_15965,N_15728);
or U16417 (N_16417,N_15765,N_15870);
xor U16418 (N_16418,N_15709,N_15511);
and U16419 (N_16419,N_15730,N_15630);
nor U16420 (N_16420,N_15768,N_15965);
or U16421 (N_16421,N_15697,N_15892);
nor U16422 (N_16422,N_15798,N_15863);
xnor U16423 (N_16423,N_15698,N_15979);
or U16424 (N_16424,N_15595,N_15686);
nor U16425 (N_16425,N_15827,N_15853);
xnor U16426 (N_16426,N_15791,N_15671);
nor U16427 (N_16427,N_15824,N_15957);
nor U16428 (N_16428,N_15833,N_15853);
and U16429 (N_16429,N_15520,N_15593);
or U16430 (N_16430,N_15988,N_15671);
nor U16431 (N_16431,N_15670,N_15826);
nor U16432 (N_16432,N_15562,N_15848);
or U16433 (N_16433,N_15649,N_15676);
or U16434 (N_16434,N_15619,N_15620);
or U16435 (N_16435,N_15805,N_15929);
or U16436 (N_16436,N_15963,N_15653);
nor U16437 (N_16437,N_15677,N_15649);
nand U16438 (N_16438,N_15953,N_15607);
and U16439 (N_16439,N_15750,N_15630);
and U16440 (N_16440,N_15828,N_15638);
nand U16441 (N_16441,N_15775,N_15801);
and U16442 (N_16442,N_15741,N_15593);
or U16443 (N_16443,N_15962,N_15792);
nor U16444 (N_16444,N_15711,N_15658);
nand U16445 (N_16445,N_15786,N_15760);
nand U16446 (N_16446,N_15647,N_15641);
nor U16447 (N_16447,N_15762,N_15542);
xnor U16448 (N_16448,N_15623,N_15613);
nor U16449 (N_16449,N_15968,N_15716);
nand U16450 (N_16450,N_15632,N_15604);
xor U16451 (N_16451,N_15603,N_15917);
or U16452 (N_16452,N_15569,N_15763);
nor U16453 (N_16453,N_15890,N_15544);
xnor U16454 (N_16454,N_15730,N_15626);
nor U16455 (N_16455,N_15679,N_15840);
and U16456 (N_16456,N_15531,N_15633);
nor U16457 (N_16457,N_15510,N_15811);
and U16458 (N_16458,N_15892,N_15610);
nand U16459 (N_16459,N_15804,N_15759);
nor U16460 (N_16460,N_15624,N_15954);
xnor U16461 (N_16461,N_15958,N_15881);
nor U16462 (N_16462,N_15889,N_15791);
nor U16463 (N_16463,N_15819,N_15575);
xnor U16464 (N_16464,N_15779,N_15610);
xor U16465 (N_16465,N_15971,N_15952);
xnor U16466 (N_16466,N_15825,N_15897);
xnor U16467 (N_16467,N_15887,N_15970);
xor U16468 (N_16468,N_15521,N_15620);
xnor U16469 (N_16469,N_15788,N_15666);
xnor U16470 (N_16470,N_15749,N_15587);
nor U16471 (N_16471,N_15909,N_15696);
xor U16472 (N_16472,N_15786,N_15989);
and U16473 (N_16473,N_15584,N_15662);
or U16474 (N_16474,N_15673,N_15609);
or U16475 (N_16475,N_15971,N_15938);
nand U16476 (N_16476,N_15925,N_15820);
or U16477 (N_16477,N_15694,N_15567);
xor U16478 (N_16478,N_15884,N_15685);
and U16479 (N_16479,N_15694,N_15864);
nor U16480 (N_16480,N_15824,N_15742);
nor U16481 (N_16481,N_15752,N_15915);
xnor U16482 (N_16482,N_15983,N_15839);
nor U16483 (N_16483,N_15967,N_15995);
nand U16484 (N_16484,N_15880,N_15570);
or U16485 (N_16485,N_15964,N_15814);
or U16486 (N_16486,N_15942,N_15978);
nor U16487 (N_16487,N_15733,N_15880);
and U16488 (N_16488,N_15621,N_15582);
nor U16489 (N_16489,N_15600,N_15615);
nand U16490 (N_16490,N_15977,N_15972);
nor U16491 (N_16491,N_15597,N_15896);
nor U16492 (N_16492,N_15952,N_15961);
xor U16493 (N_16493,N_15849,N_15754);
nor U16494 (N_16494,N_15867,N_15964);
or U16495 (N_16495,N_15672,N_15617);
nor U16496 (N_16496,N_15996,N_15876);
or U16497 (N_16497,N_15558,N_15622);
nand U16498 (N_16498,N_15814,N_15611);
nor U16499 (N_16499,N_15740,N_15781);
xor U16500 (N_16500,N_16498,N_16394);
and U16501 (N_16501,N_16410,N_16411);
nand U16502 (N_16502,N_16441,N_16357);
nor U16503 (N_16503,N_16323,N_16261);
nand U16504 (N_16504,N_16073,N_16131);
or U16505 (N_16505,N_16472,N_16107);
or U16506 (N_16506,N_16072,N_16316);
and U16507 (N_16507,N_16326,N_16228);
and U16508 (N_16508,N_16351,N_16343);
and U16509 (N_16509,N_16454,N_16226);
nor U16510 (N_16510,N_16079,N_16208);
xor U16511 (N_16511,N_16439,N_16081);
or U16512 (N_16512,N_16379,N_16287);
and U16513 (N_16513,N_16245,N_16309);
or U16514 (N_16514,N_16295,N_16429);
nand U16515 (N_16515,N_16041,N_16056);
or U16516 (N_16516,N_16468,N_16018);
or U16517 (N_16517,N_16005,N_16345);
xnor U16518 (N_16518,N_16012,N_16354);
xnor U16519 (N_16519,N_16404,N_16001);
xor U16520 (N_16520,N_16301,N_16390);
nor U16521 (N_16521,N_16098,N_16042);
and U16522 (N_16522,N_16252,N_16258);
xor U16523 (N_16523,N_16415,N_16127);
and U16524 (N_16524,N_16482,N_16060);
xnor U16525 (N_16525,N_16134,N_16125);
and U16526 (N_16526,N_16263,N_16090);
xor U16527 (N_16527,N_16270,N_16217);
or U16528 (N_16528,N_16064,N_16015);
nand U16529 (N_16529,N_16337,N_16484);
or U16530 (N_16530,N_16218,N_16160);
xnor U16531 (N_16531,N_16046,N_16278);
nor U16532 (N_16532,N_16008,N_16488);
xor U16533 (N_16533,N_16077,N_16111);
xor U16534 (N_16534,N_16413,N_16052);
nand U16535 (N_16535,N_16348,N_16367);
xor U16536 (N_16536,N_16207,N_16414);
nor U16537 (N_16537,N_16066,N_16310);
or U16538 (N_16538,N_16092,N_16435);
and U16539 (N_16539,N_16391,N_16007);
nor U16540 (N_16540,N_16034,N_16055);
or U16541 (N_16541,N_16334,N_16458);
and U16542 (N_16542,N_16496,N_16062);
or U16543 (N_16543,N_16045,N_16084);
nand U16544 (N_16544,N_16068,N_16196);
or U16545 (N_16545,N_16232,N_16133);
or U16546 (N_16546,N_16342,N_16256);
xnor U16547 (N_16547,N_16373,N_16115);
nand U16548 (N_16548,N_16445,N_16028);
nor U16549 (N_16549,N_16393,N_16156);
nand U16550 (N_16550,N_16225,N_16204);
nand U16551 (N_16551,N_16311,N_16286);
or U16552 (N_16552,N_16327,N_16304);
and U16553 (N_16553,N_16412,N_16233);
or U16554 (N_16554,N_16176,N_16402);
nor U16555 (N_16555,N_16387,N_16416);
or U16556 (N_16556,N_16210,N_16293);
nor U16557 (N_16557,N_16030,N_16014);
and U16558 (N_16558,N_16239,N_16124);
nor U16559 (N_16559,N_16102,N_16364);
and U16560 (N_16560,N_16112,N_16025);
and U16561 (N_16561,N_16251,N_16230);
or U16562 (N_16562,N_16384,N_16299);
nand U16563 (N_16563,N_16450,N_16019);
or U16564 (N_16564,N_16070,N_16231);
or U16565 (N_16565,N_16080,N_16267);
xor U16566 (N_16566,N_16021,N_16451);
or U16567 (N_16567,N_16213,N_16476);
nand U16568 (N_16568,N_16303,N_16223);
and U16569 (N_16569,N_16024,N_16183);
or U16570 (N_16570,N_16449,N_16273);
or U16571 (N_16571,N_16248,N_16362);
or U16572 (N_16572,N_16478,N_16063);
or U16573 (N_16573,N_16358,N_16203);
nand U16574 (N_16574,N_16318,N_16395);
nor U16575 (N_16575,N_16378,N_16499);
and U16576 (N_16576,N_16082,N_16117);
nor U16577 (N_16577,N_16071,N_16150);
or U16578 (N_16578,N_16474,N_16057);
xnor U16579 (N_16579,N_16162,N_16101);
nor U16580 (N_16580,N_16452,N_16302);
nor U16581 (N_16581,N_16419,N_16214);
nand U16582 (N_16582,N_16355,N_16164);
and U16583 (N_16583,N_16148,N_16200);
xnor U16584 (N_16584,N_16006,N_16136);
or U16585 (N_16585,N_16154,N_16386);
nor U16586 (N_16586,N_16308,N_16181);
and U16587 (N_16587,N_16189,N_16132);
or U16588 (N_16588,N_16175,N_16398);
or U16589 (N_16589,N_16087,N_16193);
or U16590 (N_16590,N_16365,N_16027);
nand U16591 (N_16591,N_16241,N_16460);
xor U16592 (N_16592,N_16473,N_16464);
and U16593 (N_16593,N_16209,N_16195);
and U16594 (N_16594,N_16331,N_16288);
xor U16595 (N_16595,N_16184,N_16088);
xnor U16596 (N_16596,N_16246,N_16255);
or U16597 (N_16597,N_16022,N_16141);
and U16598 (N_16598,N_16321,N_16061);
nor U16599 (N_16599,N_16177,N_16383);
nand U16600 (N_16600,N_16380,N_16469);
xnor U16601 (N_16601,N_16491,N_16155);
xnor U16602 (N_16602,N_16202,N_16433);
nor U16603 (N_16603,N_16140,N_16338);
nand U16604 (N_16604,N_16485,N_16244);
or U16605 (N_16605,N_16418,N_16423);
nand U16606 (N_16606,N_16157,N_16428);
or U16607 (N_16607,N_16280,N_16172);
and U16608 (N_16608,N_16455,N_16216);
and U16609 (N_16609,N_16249,N_16047);
nor U16610 (N_16610,N_16347,N_16237);
nand U16611 (N_16611,N_16039,N_16352);
nand U16612 (N_16612,N_16329,N_16269);
nand U16613 (N_16613,N_16040,N_16100);
xor U16614 (N_16614,N_16163,N_16053);
or U16615 (N_16615,N_16330,N_16312);
xor U16616 (N_16616,N_16099,N_16199);
and U16617 (N_16617,N_16179,N_16314);
or U16618 (N_16618,N_16294,N_16319);
xnor U16619 (N_16619,N_16477,N_16178);
nor U16620 (N_16620,N_16235,N_16322);
xnor U16621 (N_16621,N_16211,N_16389);
nor U16622 (N_16622,N_16279,N_16408);
xor U16623 (N_16623,N_16290,N_16094);
xor U16624 (N_16624,N_16283,N_16149);
or U16625 (N_16625,N_16159,N_16421);
and U16626 (N_16626,N_16197,N_16126);
xnor U16627 (N_16627,N_16422,N_16253);
or U16628 (N_16628,N_16446,N_16264);
nand U16629 (N_16629,N_16467,N_16260);
nor U16630 (N_16630,N_16424,N_16272);
and U16631 (N_16631,N_16229,N_16086);
or U16632 (N_16632,N_16259,N_16430);
xor U16633 (N_16633,N_16031,N_16250);
and U16634 (N_16634,N_16242,N_16463);
and U16635 (N_16635,N_16361,N_16443);
nor U16636 (N_16636,N_16339,N_16324);
nor U16637 (N_16637,N_16447,N_16166);
nor U16638 (N_16638,N_16281,N_16038);
nor U16639 (N_16639,N_16002,N_16085);
xnor U16640 (N_16640,N_16417,N_16219);
and U16641 (N_16641,N_16033,N_16453);
and U16642 (N_16642,N_16146,N_16145);
or U16643 (N_16643,N_16017,N_16103);
xnor U16644 (N_16644,N_16097,N_16448);
and U16645 (N_16645,N_16497,N_16276);
and U16646 (N_16646,N_16289,N_16377);
nor U16647 (N_16647,N_16201,N_16298);
or U16648 (N_16648,N_16236,N_16004);
nor U16649 (N_16649,N_16128,N_16013);
nand U16650 (N_16650,N_16392,N_16048);
nand U16651 (N_16651,N_16444,N_16492);
and U16652 (N_16652,N_16078,N_16067);
and U16653 (N_16653,N_16108,N_16003);
nor U16654 (N_16654,N_16116,N_16049);
nand U16655 (N_16655,N_16481,N_16461);
or U16656 (N_16656,N_16284,N_16059);
or U16657 (N_16657,N_16265,N_16407);
xnor U16658 (N_16658,N_16268,N_16471);
xor U16659 (N_16659,N_16396,N_16247);
or U16660 (N_16660,N_16317,N_16306);
nand U16661 (N_16661,N_16009,N_16143);
nand U16662 (N_16662,N_16296,N_16091);
and U16663 (N_16663,N_16307,N_16371);
or U16664 (N_16664,N_16029,N_16050);
nand U16665 (N_16665,N_16313,N_16328);
nor U16666 (N_16666,N_16370,N_16388);
nand U16667 (N_16667,N_16074,N_16336);
nor U16668 (N_16668,N_16401,N_16405);
and U16669 (N_16669,N_16020,N_16479);
xor U16670 (N_16670,N_16069,N_16212);
or U16671 (N_16671,N_16432,N_16147);
xnor U16672 (N_16672,N_16138,N_16425);
or U16673 (N_16673,N_16180,N_16360);
or U16674 (N_16674,N_16104,N_16043);
xor U16675 (N_16675,N_16121,N_16480);
or U16676 (N_16676,N_16490,N_16010);
or U16677 (N_16677,N_16105,N_16483);
nand U16678 (N_16678,N_16106,N_16266);
nand U16679 (N_16679,N_16332,N_16486);
and U16680 (N_16680,N_16168,N_16438);
nor U16681 (N_16681,N_16120,N_16152);
nor U16682 (N_16682,N_16493,N_16385);
xor U16683 (N_16683,N_16494,N_16442);
and U16684 (N_16684,N_16076,N_16349);
and U16685 (N_16685,N_16431,N_16167);
and U16686 (N_16686,N_16489,N_16220);
or U16687 (N_16687,N_16277,N_16016);
and U16688 (N_16688,N_16165,N_16096);
and U16689 (N_16689,N_16173,N_16054);
nand U16690 (N_16690,N_16194,N_16151);
or U16691 (N_16691,N_16400,N_16083);
or U16692 (N_16692,N_16320,N_16109);
nor U16693 (N_16693,N_16129,N_16254);
nor U16694 (N_16694,N_16275,N_16466);
nand U16695 (N_16695,N_16135,N_16426);
and U16696 (N_16696,N_16037,N_16240);
xor U16697 (N_16697,N_16114,N_16409);
nor U16698 (N_16698,N_16243,N_16036);
and U16699 (N_16699,N_16427,N_16187);
or U16700 (N_16700,N_16185,N_16325);
and U16701 (N_16701,N_16356,N_16359);
xnor U16702 (N_16702,N_16300,N_16113);
xor U16703 (N_16703,N_16182,N_16353);
xnor U16704 (N_16704,N_16089,N_16174);
nand U16705 (N_16705,N_16374,N_16274);
or U16706 (N_16706,N_16291,N_16170);
and U16707 (N_16707,N_16495,N_16344);
xnor U16708 (N_16708,N_16191,N_16462);
nor U16709 (N_16709,N_16363,N_16095);
xnor U16710 (N_16710,N_16487,N_16171);
nor U16711 (N_16711,N_16381,N_16224);
or U16712 (N_16712,N_16257,N_16198);
nor U16713 (N_16713,N_16139,N_16123);
nor U16714 (N_16714,N_16369,N_16142);
nand U16715 (N_16715,N_16333,N_16457);
or U16716 (N_16716,N_16205,N_16075);
and U16717 (N_16717,N_16023,N_16065);
nand U16718 (N_16718,N_16110,N_16305);
or U16719 (N_16719,N_16285,N_16227);
nor U16720 (N_16720,N_16222,N_16188);
nor U16721 (N_16721,N_16459,N_16119);
nor U16722 (N_16722,N_16350,N_16011);
nand U16723 (N_16723,N_16292,N_16032);
and U16724 (N_16724,N_16035,N_16420);
xnor U16725 (N_16725,N_16161,N_16058);
and U16726 (N_16726,N_16238,N_16215);
nor U16727 (N_16727,N_16169,N_16234);
or U16728 (N_16728,N_16153,N_16340);
nor U16729 (N_16729,N_16206,N_16406);
nand U16730 (N_16730,N_16366,N_16399);
or U16731 (N_16731,N_16144,N_16382);
nand U16732 (N_16732,N_16130,N_16437);
or U16733 (N_16733,N_16158,N_16190);
nor U16734 (N_16734,N_16470,N_16375);
xor U16735 (N_16735,N_16456,N_16026);
or U16736 (N_16736,N_16475,N_16000);
nor U16737 (N_16737,N_16346,N_16341);
xor U16738 (N_16738,N_16335,N_16192);
nor U16739 (N_16739,N_16271,N_16282);
xor U16740 (N_16740,N_16315,N_16093);
nor U16741 (N_16741,N_16368,N_16051);
nand U16742 (N_16742,N_16372,N_16297);
or U16743 (N_16743,N_16434,N_16465);
xnor U16744 (N_16744,N_16137,N_16122);
or U16745 (N_16745,N_16221,N_16262);
and U16746 (N_16746,N_16186,N_16044);
and U16747 (N_16747,N_16403,N_16397);
nand U16748 (N_16748,N_16440,N_16436);
nand U16749 (N_16749,N_16376,N_16118);
nor U16750 (N_16750,N_16191,N_16027);
or U16751 (N_16751,N_16250,N_16435);
nor U16752 (N_16752,N_16088,N_16400);
nand U16753 (N_16753,N_16302,N_16195);
nand U16754 (N_16754,N_16391,N_16444);
xnor U16755 (N_16755,N_16199,N_16345);
and U16756 (N_16756,N_16263,N_16145);
and U16757 (N_16757,N_16047,N_16111);
xor U16758 (N_16758,N_16237,N_16145);
nand U16759 (N_16759,N_16042,N_16266);
nand U16760 (N_16760,N_16057,N_16483);
xnor U16761 (N_16761,N_16001,N_16327);
nand U16762 (N_16762,N_16423,N_16014);
xnor U16763 (N_16763,N_16349,N_16246);
and U16764 (N_16764,N_16042,N_16167);
xnor U16765 (N_16765,N_16159,N_16152);
nand U16766 (N_16766,N_16459,N_16362);
or U16767 (N_16767,N_16451,N_16467);
or U16768 (N_16768,N_16479,N_16437);
and U16769 (N_16769,N_16490,N_16244);
or U16770 (N_16770,N_16255,N_16199);
and U16771 (N_16771,N_16309,N_16332);
and U16772 (N_16772,N_16047,N_16415);
nor U16773 (N_16773,N_16387,N_16080);
or U16774 (N_16774,N_16393,N_16187);
or U16775 (N_16775,N_16040,N_16142);
and U16776 (N_16776,N_16085,N_16489);
nand U16777 (N_16777,N_16475,N_16050);
nand U16778 (N_16778,N_16493,N_16006);
nor U16779 (N_16779,N_16445,N_16413);
nor U16780 (N_16780,N_16407,N_16003);
xnor U16781 (N_16781,N_16458,N_16379);
or U16782 (N_16782,N_16487,N_16441);
and U16783 (N_16783,N_16037,N_16232);
or U16784 (N_16784,N_16281,N_16143);
and U16785 (N_16785,N_16464,N_16274);
and U16786 (N_16786,N_16360,N_16355);
or U16787 (N_16787,N_16169,N_16427);
xor U16788 (N_16788,N_16473,N_16366);
or U16789 (N_16789,N_16445,N_16487);
or U16790 (N_16790,N_16495,N_16389);
and U16791 (N_16791,N_16201,N_16127);
and U16792 (N_16792,N_16466,N_16022);
and U16793 (N_16793,N_16182,N_16358);
nor U16794 (N_16794,N_16366,N_16088);
xor U16795 (N_16795,N_16097,N_16477);
and U16796 (N_16796,N_16290,N_16451);
and U16797 (N_16797,N_16018,N_16100);
or U16798 (N_16798,N_16339,N_16361);
and U16799 (N_16799,N_16006,N_16065);
or U16800 (N_16800,N_16095,N_16255);
or U16801 (N_16801,N_16348,N_16295);
and U16802 (N_16802,N_16170,N_16355);
nand U16803 (N_16803,N_16334,N_16034);
nand U16804 (N_16804,N_16375,N_16136);
nor U16805 (N_16805,N_16491,N_16277);
nor U16806 (N_16806,N_16157,N_16398);
and U16807 (N_16807,N_16370,N_16480);
or U16808 (N_16808,N_16317,N_16180);
or U16809 (N_16809,N_16246,N_16085);
xor U16810 (N_16810,N_16365,N_16292);
nand U16811 (N_16811,N_16282,N_16103);
nand U16812 (N_16812,N_16466,N_16432);
xor U16813 (N_16813,N_16366,N_16498);
xor U16814 (N_16814,N_16211,N_16314);
and U16815 (N_16815,N_16229,N_16394);
nand U16816 (N_16816,N_16402,N_16022);
nor U16817 (N_16817,N_16114,N_16127);
nand U16818 (N_16818,N_16335,N_16071);
nand U16819 (N_16819,N_16460,N_16184);
nor U16820 (N_16820,N_16250,N_16007);
or U16821 (N_16821,N_16493,N_16322);
nand U16822 (N_16822,N_16054,N_16006);
or U16823 (N_16823,N_16081,N_16464);
and U16824 (N_16824,N_16325,N_16160);
or U16825 (N_16825,N_16396,N_16239);
xor U16826 (N_16826,N_16153,N_16215);
and U16827 (N_16827,N_16158,N_16286);
or U16828 (N_16828,N_16466,N_16179);
xor U16829 (N_16829,N_16414,N_16060);
nand U16830 (N_16830,N_16471,N_16338);
or U16831 (N_16831,N_16238,N_16096);
and U16832 (N_16832,N_16476,N_16224);
xor U16833 (N_16833,N_16252,N_16403);
nand U16834 (N_16834,N_16100,N_16412);
nor U16835 (N_16835,N_16213,N_16353);
xnor U16836 (N_16836,N_16036,N_16410);
nor U16837 (N_16837,N_16464,N_16032);
nand U16838 (N_16838,N_16274,N_16399);
and U16839 (N_16839,N_16144,N_16295);
nand U16840 (N_16840,N_16140,N_16364);
nor U16841 (N_16841,N_16202,N_16316);
and U16842 (N_16842,N_16249,N_16073);
nor U16843 (N_16843,N_16305,N_16380);
and U16844 (N_16844,N_16470,N_16431);
or U16845 (N_16845,N_16089,N_16384);
nand U16846 (N_16846,N_16397,N_16244);
nand U16847 (N_16847,N_16357,N_16370);
and U16848 (N_16848,N_16087,N_16195);
nor U16849 (N_16849,N_16004,N_16481);
or U16850 (N_16850,N_16062,N_16066);
or U16851 (N_16851,N_16034,N_16218);
xor U16852 (N_16852,N_16188,N_16441);
or U16853 (N_16853,N_16131,N_16050);
nand U16854 (N_16854,N_16126,N_16252);
nor U16855 (N_16855,N_16291,N_16111);
xnor U16856 (N_16856,N_16246,N_16199);
xor U16857 (N_16857,N_16334,N_16046);
or U16858 (N_16858,N_16483,N_16300);
nor U16859 (N_16859,N_16399,N_16152);
xnor U16860 (N_16860,N_16362,N_16415);
and U16861 (N_16861,N_16154,N_16135);
nand U16862 (N_16862,N_16125,N_16189);
nand U16863 (N_16863,N_16459,N_16487);
xnor U16864 (N_16864,N_16164,N_16197);
and U16865 (N_16865,N_16292,N_16310);
and U16866 (N_16866,N_16347,N_16205);
or U16867 (N_16867,N_16171,N_16320);
xor U16868 (N_16868,N_16300,N_16138);
nand U16869 (N_16869,N_16055,N_16423);
and U16870 (N_16870,N_16454,N_16371);
nand U16871 (N_16871,N_16118,N_16462);
nand U16872 (N_16872,N_16152,N_16369);
xor U16873 (N_16873,N_16344,N_16220);
and U16874 (N_16874,N_16082,N_16221);
or U16875 (N_16875,N_16056,N_16126);
nand U16876 (N_16876,N_16317,N_16029);
xor U16877 (N_16877,N_16341,N_16289);
or U16878 (N_16878,N_16437,N_16089);
or U16879 (N_16879,N_16241,N_16195);
nand U16880 (N_16880,N_16244,N_16467);
nor U16881 (N_16881,N_16258,N_16281);
and U16882 (N_16882,N_16125,N_16190);
or U16883 (N_16883,N_16007,N_16312);
or U16884 (N_16884,N_16329,N_16331);
or U16885 (N_16885,N_16388,N_16033);
nor U16886 (N_16886,N_16311,N_16470);
xor U16887 (N_16887,N_16445,N_16023);
or U16888 (N_16888,N_16385,N_16024);
xnor U16889 (N_16889,N_16456,N_16260);
xnor U16890 (N_16890,N_16436,N_16200);
xor U16891 (N_16891,N_16286,N_16241);
and U16892 (N_16892,N_16306,N_16008);
nand U16893 (N_16893,N_16190,N_16169);
nor U16894 (N_16894,N_16288,N_16272);
nor U16895 (N_16895,N_16317,N_16291);
nand U16896 (N_16896,N_16455,N_16251);
or U16897 (N_16897,N_16203,N_16005);
nor U16898 (N_16898,N_16385,N_16092);
nand U16899 (N_16899,N_16191,N_16303);
and U16900 (N_16900,N_16339,N_16332);
nor U16901 (N_16901,N_16117,N_16262);
and U16902 (N_16902,N_16118,N_16062);
and U16903 (N_16903,N_16150,N_16355);
and U16904 (N_16904,N_16026,N_16454);
xnor U16905 (N_16905,N_16020,N_16090);
and U16906 (N_16906,N_16354,N_16246);
or U16907 (N_16907,N_16116,N_16244);
and U16908 (N_16908,N_16053,N_16180);
or U16909 (N_16909,N_16306,N_16121);
or U16910 (N_16910,N_16233,N_16140);
nor U16911 (N_16911,N_16177,N_16083);
xor U16912 (N_16912,N_16047,N_16446);
and U16913 (N_16913,N_16109,N_16317);
nor U16914 (N_16914,N_16035,N_16250);
or U16915 (N_16915,N_16198,N_16139);
nand U16916 (N_16916,N_16314,N_16197);
nor U16917 (N_16917,N_16406,N_16494);
nand U16918 (N_16918,N_16432,N_16465);
nor U16919 (N_16919,N_16023,N_16028);
or U16920 (N_16920,N_16352,N_16435);
or U16921 (N_16921,N_16198,N_16433);
xnor U16922 (N_16922,N_16315,N_16270);
xor U16923 (N_16923,N_16086,N_16452);
or U16924 (N_16924,N_16060,N_16252);
nand U16925 (N_16925,N_16102,N_16173);
and U16926 (N_16926,N_16121,N_16106);
xor U16927 (N_16927,N_16429,N_16239);
and U16928 (N_16928,N_16277,N_16387);
xor U16929 (N_16929,N_16017,N_16384);
nor U16930 (N_16930,N_16335,N_16134);
and U16931 (N_16931,N_16116,N_16272);
nand U16932 (N_16932,N_16145,N_16346);
nand U16933 (N_16933,N_16387,N_16454);
xnor U16934 (N_16934,N_16466,N_16067);
nand U16935 (N_16935,N_16142,N_16350);
and U16936 (N_16936,N_16041,N_16348);
or U16937 (N_16937,N_16277,N_16157);
nand U16938 (N_16938,N_16422,N_16488);
and U16939 (N_16939,N_16206,N_16470);
nor U16940 (N_16940,N_16382,N_16414);
nor U16941 (N_16941,N_16475,N_16398);
xor U16942 (N_16942,N_16334,N_16141);
and U16943 (N_16943,N_16409,N_16337);
or U16944 (N_16944,N_16042,N_16212);
or U16945 (N_16945,N_16418,N_16347);
nand U16946 (N_16946,N_16445,N_16235);
or U16947 (N_16947,N_16324,N_16443);
nor U16948 (N_16948,N_16223,N_16413);
or U16949 (N_16949,N_16115,N_16103);
or U16950 (N_16950,N_16208,N_16461);
or U16951 (N_16951,N_16159,N_16165);
xor U16952 (N_16952,N_16229,N_16401);
nand U16953 (N_16953,N_16338,N_16037);
nand U16954 (N_16954,N_16458,N_16269);
nor U16955 (N_16955,N_16321,N_16456);
nand U16956 (N_16956,N_16131,N_16299);
or U16957 (N_16957,N_16469,N_16309);
and U16958 (N_16958,N_16199,N_16127);
or U16959 (N_16959,N_16190,N_16239);
xnor U16960 (N_16960,N_16008,N_16314);
or U16961 (N_16961,N_16321,N_16178);
xnor U16962 (N_16962,N_16104,N_16210);
and U16963 (N_16963,N_16140,N_16431);
or U16964 (N_16964,N_16442,N_16169);
xnor U16965 (N_16965,N_16234,N_16079);
and U16966 (N_16966,N_16342,N_16314);
nor U16967 (N_16967,N_16261,N_16335);
or U16968 (N_16968,N_16151,N_16088);
or U16969 (N_16969,N_16330,N_16070);
nor U16970 (N_16970,N_16008,N_16186);
xnor U16971 (N_16971,N_16126,N_16091);
or U16972 (N_16972,N_16226,N_16130);
nor U16973 (N_16973,N_16348,N_16384);
nor U16974 (N_16974,N_16497,N_16189);
or U16975 (N_16975,N_16367,N_16241);
and U16976 (N_16976,N_16361,N_16101);
and U16977 (N_16977,N_16002,N_16334);
or U16978 (N_16978,N_16145,N_16168);
or U16979 (N_16979,N_16190,N_16482);
nor U16980 (N_16980,N_16062,N_16191);
or U16981 (N_16981,N_16062,N_16279);
xor U16982 (N_16982,N_16038,N_16156);
xor U16983 (N_16983,N_16346,N_16403);
xnor U16984 (N_16984,N_16330,N_16031);
nand U16985 (N_16985,N_16275,N_16087);
and U16986 (N_16986,N_16308,N_16015);
or U16987 (N_16987,N_16402,N_16268);
nand U16988 (N_16988,N_16149,N_16249);
xnor U16989 (N_16989,N_16041,N_16367);
nand U16990 (N_16990,N_16386,N_16369);
xor U16991 (N_16991,N_16148,N_16186);
nand U16992 (N_16992,N_16349,N_16127);
xor U16993 (N_16993,N_16195,N_16490);
xnor U16994 (N_16994,N_16350,N_16257);
xnor U16995 (N_16995,N_16234,N_16267);
nand U16996 (N_16996,N_16478,N_16267);
or U16997 (N_16997,N_16359,N_16414);
or U16998 (N_16998,N_16222,N_16290);
nor U16999 (N_16999,N_16141,N_16008);
nor U17000 (N_17000,N_16778,N_16744);
nand U17001 (N_17001,N_16645,N_16836);
and U17002 (N_17002,N_16956,N_16805);
nand U17003 (N_17003,N_16603,N_16804);
or U17004 (N_17004,N_16726,N_16987);
nand U17005 (N_17005,N_16661,N_16644);
and U17006 (N_17006,N_16742,N_16948);
or U17007 (N_17007,N_16602,N_16528);
nand U17008 (N_17008,N_16981,N_16894);
nand U17009 (N_17009,N_16860,N_16776);
and U17010 (N_17010,N_16574,N_16738);
nor U17011 (N_17011,N_16656,N_16908);
and U17012 (N_17012,N_16830,N_16994);
and U17013 (N_17013,N_16713,N_16789);
and U17014 (N_17014,N_16608,N_16712);
nand U17015 (N_17015,N_16698,N_16692);
nand U17016 (N_17016,N_16695,N_16892);
nor U17017 (N_17017,N_16677,N_16861);
nor U17018 (N_17018,N_16967,N_16785);
nor U17019 (N_17019,N_16732,N_16501);
or U17020 (N_17020,N_16992,N_16588);
and U17021 (N_17021,N_16506,N_16817);
or U17022 (N_17022,N_16901,N_16984);
nand U17023 (N_17023,N_16708,N_16990);
nand U17024 (N_17024,N_16592,N_16702);
or U17025 (N_17025,N_16769,N_16910);
xnor U17026 (N_17026,N_16885,N_16735);
or U17027 (N_17027,N_16845,N_16676);
nand U17028 (N_17028,N_16896,N_16569);
nand U17029 (N_17029,N_16583,N_16640);
or U17030 (N_17030,N_16549,N_16826);
nand U17031 (N_17031,N_16965,N_16904);
or U17032 (N_17032,N_16853,N_16686);
xor U17033 (N_17033,N_16977,N_16669);
xor U17034 (N_17034,N_16774,N_16566);
nor U17035 (N_17035,N_16810,N_16706);
nor U17036 (N_17036,N_16689,N_16673);
xor U17037 (N_17037,N_16754,N_16643);
or U17038 (N_17038,N_16560,N_16950);
nor U17039 (N_17039,N_16564,N_16606);
nand U17040 (N_17040,N_16832,N_16957);
nand U17041 (N_17041,N_16516,N_16972);
and U17042 (N_17042,N_16944,N_16850);
xnor U17043 (N_17043,N_16936,N_16511);
xor U17044 (N_17044,N_16868,N_16631);
nand U17045 (N_17045,N_16898,N_16837);
nor U17046 (N_17046,N_16554,N_16615);
or U17047 (N_17047,N_16775,N_16895);
nor U17048 (N_17048,N_16642,N_16862);
xor U17049 (N_17049,N_16970,N_16522);
nand U17050 (N_17050,N_16607,N_16681);
xor U17051 (N_17051,N_16581,N_16833);
and U17052 (N_17052,N_16865,N_16985);
xnor U17053 (N_17053,N_16856,N_16544);
and U17054 (N_17054,N_16703,N_16768);
and U17055 (N_17055,N_16991,N_16730);
xnor U17056 (N_17056,N_16829,N_16928);
and U17057 (N_17057,N_16838,N_16548);
nor U17058 (N_17058,N_16650,N_16601);
and U17059 (N_17059,N_16932,N_16843);
nor U17060 (N_17060,N_16568,N_16727);
nand U17061 (N_17061,N_16524,N_16561);
nor U17062 (N_17062,N_16858,N_16940);
xor U17063 (N_17063,N_16973,N_16873);
xor U17064 (N_17064,N_16664,N_16530);
nor U17065 (N_17065,N_16866,N_16960);
nor U17066 (N_17066,N_16534,N_16556);
or U17067 (N_17067,N_16619,N_16777);
nor U17068 (N_17068,N_16504,N_16889);
xnor U17069 (N_17069,N_16629,N_16515);
or U17070 (N_17070,N_16959,N_16941);
nand U17071 (N_17071,N_16827,N_16694);
and U17072 (N_17072,N_16551,N_16532);
xnor U17073 (N_17073,N_16766,N_16546);
nand U17074 (N_17074,N_16864,N_16600);
xnor U17075 (N_17075,N_16998,N_16938);
and U17076 (N_17076,N_16596,N_16507);
and U17077 (N_17077,N_16872,N_16880);
nand U17078 (N_17078,N_16668,N_16540);
or U17079 (N_17079,N_16671,N_16746);
xnor U17080 (N_17080,N_16797,N_16926);
xnor U17081 (N_17081,N_16584,N_16796);
nor U17082 (N_17082,N_16764,N_16809);
nand U17083 (N_17083,N_16709,N_16573);
and U17084 (N_17084,N_16680,N_16711);
or U17085 (N_17085,N_16597,N_16610);
nand U17086 (N_17086,N_16899,N_16510);
nand U17087 (N_17087,N_16587,N_16812);
or U17088 (N_17088,N_16691,N_16842);
and U17089 (N_17089,N_16787,N_16783);
nand U17090 (N_17090,N_16772,N_16638);
or U17091 (N_17091,N_16930,N_16997);
or U17092 (N_17092,N_16575,N_16514);
nor U17093 (N_17093,N_16578,N_16792);
and U17094 (N_17094,N_16627,N_16937);
xor U17095 (N_17095,N_16788,N_16718);
or U17096 (N_17096,N_16536,N_16943);
or U17097 (N_17097,N_16927,N_16923);
and U17098 (N_17098,N_16893,N_16751);
xor U17099 (N_17099,N_16969,N_16846);
nor U17100 (N_17100,N_16550,N_16803);
and U17101 (N_17101,N_16799,N_16869);
xor U17102 (N_17102,N_16814,N_16533);
and U17103 (N_17103,N_16633,N_16626);
or U17104 (N_17104,N_16877,N_16793);
nor U17105 (N_17105,N_16700,N_16641);
or U17106 (N_17106,N_16798,N_16527);
and U17107 (N_17107,N_16974,N_16502);
nor U17108 (N_17108,N_16781,N_16834);
xnor U17109 (N_17109,N_16586,N_16825);
or U17110 (N_17110,N_16674,N_16882);
nand U17111 (N_17111,N_16841,N_16848);
and U17112 (N_17112,N_16637,N_16851);
or U17113 (N_17113,N_16500,N_16818);
nand U17114 (N_17114,N_16745,N_16667);
nor U17115 (N_17115,N_16947,N_16958);
and U17116 (N_17116,N_16741,N_16765);
and U17117 (N_17117,N_16594,N_16929);
or U17118 (N_17118,N_16962,N_16897);
nor U17119 (N_17119,N_16807,N_16949);
nor U17120 (N_17120,N_16852,N_16808);
xor U17121 (N_17121,N_16525,N_16755);
nand U17122 (N_17122,N_16963,N_16978);
xnor U17123 (N_17123,N_16690,N_16599);
nand U17124 (N_17124,N_16675,N_16704);
nand U17125 (N_17125,N_16729,N_16593);
nand U17126 (N_17126,N_16577,N_16784);
nand U17127 (N_17127,N_16687,N_16685);
nor U17128 (N_17128,N_16934,N_16911);
nand U17129 (N_17129,N_16771,N_16802);
nor U17130 (N_17130,N_16721,N_16635);
nor U17131 (N_17131,N_16773,N_16859);
nand U17132 (N_17132,N_16678,N_16646);
or U17133 (N_17133,N_16761,N_16535);
nor U17134 (N_17134,N_16995,N_16790);
nand U17135 (N_17135,N_16870,N_16683);
or U17136 (N_17136,N_16747,N_16800);
and U17137 (N_17137,N_16905,N_16662);
and U17138 (N_17138,N_16831,N_16907);
nand U17139 (N_17139,N_16717,N_16562);
nand U17140 (N_17140,N_16922,N_16756);
nand U17141 (N_17141,N_16611,N_16734);
xnor U17142 (N_17142,N_16557,N_16740);
xnor U17143 (N_17143,N_16519,N_16714);
xnor U17144 (N_17144,N_16770,N_16719);
nand U17145 (N_17145,N_16913,N_16579);
nor U17146 (N_17146,N_16531,N_16736);
or U17147 (N_17147,N_16979,N_16925);
and U17148 (N_17148,N_16688,N_16613);
or U17149 (N_17149,N_16902,N_16705);
nand U17150 (N_17150,N_16976,N_16921);
or U17151 (N_17151,N_16720,N_16945);
or U17152 (N_17152,N_16612,N_16743);
nand U17153 (N_17153,N_16563,N_16855);
and U17154 (N_17154,N_16975,N_16565);
nand U17155 (N_17155,N_16854,N_16822);
and U17156 (N_17156,N_16715,N_16779);
nor U17157 (N_17157,N_16996,N_16699);
xor U17158 (N_17158,N_16946,N_16980);
xor U17159 (N_17159,N_16903,N_16659);
or U17160 (N_17160,N_16966,N_16555);
xor U17161 (N_17161,N_16657,N_16823);
and U17162 (N_17162,N_16537,N_16986);
xor U17163 (N_17163,N_16780,N_16820);
xor U17164 (N_17164,N_16933,N_16993);
xnor U17165 (N_17165,N_16670,N_16508);
and U17166 (N_17166,N_16585,N_16939);
and U17167 (N_17167,N_16538,N_16666);
or U17168 (N_17168,N_16722,N_16795);
or U17169 (N_17169,N_16849,N_16647);
nand U17170 (N_17170,N_16665,N_16867);
xor U17171 (N_17171,N_16914,N_16697);
or U17172 (N_17172,N_16623,N_16900);
nand U17173 (N_17173,N_16821,N_16813);
nor U17174 (N_17174,N_16758,N_16636);
nand U17175 (N_17175,N_16503,N_16884);
or U17176 (N_17176,N_16570,N_16652);
and U17177 (N_17177,N_16824,N_16876);
nor U17178 (N_17178,N_16580,N_16693);
nor U17179 (N_17179,N_16886,N_16786);
nor U17180 (N_17180,N_16542,N_16526);
and U17181 (N_17181,N_16649,N_16559);
nand U17182 (N_17182,N_16521,N_16553);
and U17183 (N_17183,N_16663,N_16589);
or U17184 (N_17184,N_16935,N_16624);
or U17185 (N_17185,N_16890,N_16881);
nand U17186 (N_17186,N_16888,N_16816);
nand U17187 (N_17187,N_16828,N_16920);
and U17188 (N_17188,N_16547,N_16763);
xor U17189 (N_17189,N_16748,N_16598);
nand U17190 (N_17190,N_16582,N_16952);
nor U17191 (N_17191,N_16955,N_16523);
and U17192 (N_17192,N_16794,N_16942);
nor U17193 (N_17193,N_16621,N_16961);
nor U17194 (N_17194,N_16614,N_16953);
and U17195 (N_17195,N_16634,N_16628);
nor U17196 (N_17196,N_16819,N_16620);
nand U17197 (N_17197,N_16616,N_16716);
and U17198 (N_17198,N_16639,N_16617);
and U17199 (N_17199,N_16767,N_16707);
xor U17200 (N_17200,N_16604,N_16847);
and U17201 (N_17201,N_16815,N_16753);
nand U17202 (N_17202,N_16571,N_16924);
or U17203 (N_17203,N_16558,N_16917);
or U17204 (N_17204,N_16840,N_16622);
or U17205 (N_17205,N_16999,N_16739);
and U17206 (N_17206,N_16931,N_16609);
xnor U17207 (N_17207,N_16916,N_16505);
and U17208 (N_17208,N_16918,N_16811);
nand U17209 (N_17209,N_16682,N_16543);
xnor U17210 (N_17210,N_16863,N_16724);
xnor U17211 (N_17211,N_16839,N_16909);
nor U17212 (N_17212,N_16791,N_16954);
nor U17213 (N_17213,N_16982,N_16518);
and U17214 (N_17214,N_16731,N_16517);
and U17215 (N_17215,N_16857,N_16879);
or U17216 (N_17216,N_16968,N_16590);
xnor U17217 (N_17217,N_16725,N_16964);
xor U17218 (N_17218,N_16757,N_16513);
and U17219 (N_17219,N_16572,N_16749);
and U17220 (N_17220,N_16660,N_16632);
and U17221 (N_17221,N_16576,N_16651);
xnor U17222 (N_17222,N_16915,N_16567);
nor U17223 (N_17223,N_16762,N_16520);
nand U17224 (N_17224,N_16541,N_16529);
nor U17225 (N_17225,N_16723,N_16906);
nor U17226 (N_17226,N_16728,N_16625);
xor U17227 (N_17227,N_16883,N_16801);
or U17228 (N_17228,N_16835,N_16887);
nand U17229 (N_17229,N_16733,N_16684);
nor U17230 (N_17230,N_16654,N_16679);
nor U17231 (N_17231,N_16750,N_16710);
nand U17232 (N_17232,N_16988,N_16509);
and U17233 (N_17233,N_16591,N_16891);
and U17234 (N_17234,N_16759,N_16545);
nand U17235 (N_17235,N_16648,N_16875);
xnor U17236 (N_17236,N_16595,N_16512);
nand U17237 (N_17237,N_16658,N_16983);
xnor U17238 (N_17238,N_16806,N_16878);
nor U17239 (N_17239,N_16696,N_16951);
or U17240 (N_17240,N_16919,N_16971);
nand U17241 (N_17241,N_16874,N_16871);
or U17242 (N_17242,N_16630,N_16737);
xor U17243 (N_17243,N_16672,N_16782);
nor U17244 (N_17244,N_16844,N_16539);
nor U17245 (N_17245,N_16760,N_16655);
xor U17246 (N_17246,N_16653,N_16618);
xor U17247 (N_17247,N_16752,N_16912);
and U17248 (N_17248,N_16552,N_16701);
or U17249 (N_17249,N_16605,N_16989);
and U17250 (N_17250,N_16937,N_16905);
nor U17251 (N_17251,N_16649,N_16576);
nor U17252 (N_17252,N_16500,N_16904);
nor U17253 (N_17253,N_16847,N_16556);
xnor U17254 (N_17254,N_16619,N_16540);
nor U17255 (N_17255,N_16772,N_16531);
or U17256 (N_17256,N_16893,N_16948);
and U17257 (N_17257,N_16801,N_16503);
xor U17258 (N_17258,N_16717,N_16803);
nor U17259 (N_17259,N_16640,N_16814);
and U17260 (N_17260,N_16999,N_16546);
nand U17261 (N_17261,N_16873,N_16551);
and U17262 (N_17262,N_16627,N_16543);
xor U17263 (N_17263,N_16551,N_16755);
nor U17264 (N_17264,N_16878,N_16694);
nor U17265 (N_17265,N_16859,N_16813);
nand U17266 (N_17266,N_16625,N_16887);
nand U17267 (N_17267,N_16803,N_16640);
and U17268 (N_17268,N_16731,N_16891);
nand U17269 (N_17269,N_16976,N_16960);
nand U17270 (N_17270,N_16736,N_16622);
xnor U17271 (N_17271,N_16982,N_16988);
nor U17272 (N_17272,N_16658,N_16500);
nand U17273 (N_17273,N_16644,N_16870);
and U17274 (N_17274,N_16703,N_16807);
nor U17275 (N_17275,N_16951,N_16645);
nor U17276 (N_17276,N_16645,N_16827);
nand U17277 (N_17277,N_16910,N_16966);
nand U17278 (N_17278,N_16534,N_16632);
nand U17279 (N_17279,N_16638,N_16758);
and U17280 (N_17280,N_16795,N_16556);
and U17281 (N_17281,N_16918,N_16770);
nand U17282 (N_17282,N_16844,N_16901);
nand U17283 (N_17283,N_16708,N_16950);
nand U17284 (N_17284,N_16691,N_16806);
nand U17285 (N_17285,N_16617,N_16637);
nand U17286 (N_17286,N_16702,N_16679);
nor U17287 (N_17287,N_16857,N_16513);
or U17288 (N_17288,N_16875,N_16868);
or U17289 (N_17289,N_16830,N_16636);
or U17290 (N_17290,N_16814,N_16969);
and U17291 (N_17291,N_16862,N_16986);
and U17292 (N_17292,N_16681,N_16537);
nor U17293 (N_17293,N_16765,N_16641);
or U17294 (N_17294,N_16564,N_16835);
xnor U17295 (N_17295,N_16804,N_16543);
nor U17296 (N_17296,N_16773,N_16883);
xor U17297 (N_17297,N_16863,N_16994);
or U17298 (N_17298,N_16776,N_16584);
nor U17299 (N_17299,N_16622,N_16831);
xor U17300 (N_17300,N_16725,N_16550);
and U17301 (N_17301,N_16513,N_16937);
or U17302 (N_17302,N_16841,N_16769);
xnor U17303 (N_17303,N_16835,N_16686);
nor U17304 (N_17304,N_16981,N_16756);
nor U17305 (N_17305,N_16665,N_16790);
xnor U17306 (N_17306,N_16699,N_16669);
nand U17307 (N_17307,N_16666,N_16876);
xor U17308 (N_17308,N_16617,N_16560);
or U17309 (N_17309,N_16517,N_16641);
xor U17310 (N_17310,N_16657,N_16559);
and U17311 (N_17311,N_16944,N_16955);
and U17312 (N_17312,N_16777,N_16964);
xor U17313 (N_17313,N_16952,N_16817);
xor U17314 (N_17314,N_16921,N_16707);
nor U17315 (N_17315,N_16757,N_16681);
nor U17316 (N_17316,N_16694,N_16519);
nand U17317 (N_17317,N_16753,N_16898);
xnor U17318 (N_17318,N_16650,N_16540);
and U17319 (N_17319,N_16642,N_16744);
nor U17320 (N_17320,N_16963,N_16733);
nor U17321 (N_17321,N_16768,N_16686);
and U17322 (N_17322,N_16997,N_16874);
nand U17323 (N_17323,N_16680,N_16671);
xnor U17324 (N_17324,N_16707,N_16636);
and U17325 (N_17325,N_16867,N_16908);
xnor U17326 (N_17326,N_16756,N_16685);
and U17327 (N_17327,N_16905,N_16598);
xnor U17328 (N_17328,N_16592,N_16682);
nor U17329 (N_17329,N_16748,N_16953);
xnor U17330 (N_17330,N_16817,N_16681);
and U17331 (N_17331,N_16503,N_16952);
or U17332 (N_17332,N_16862,N_16654);
xnor U17333 (N_17333,N_16677,N_16680);
nand U17334 (N_17334,N_16618,N_16609);
nor U17335 (N_17335,N_16604,N_16677);
xnor U17336 (N_17336,N_16978,N_16819);
nor U17337 (N_17337,N_16849,N_16593);
and U17338 (N_17338,N_16577,N_16974);
xor U17339 (N_17339,N_16653,N_16759);
or U17340 (N_17340,N_16662,N_16788);
or U17341 (N_17341,N_16995,N_16567);
nor U17342 (N_17342,N_16748,N_16629);
nand U17343 (N_17343,N_16805,N_16560);
nor U17344 (N_17344,N_16806,N_16957);
or U17345 (N_17345,N_16887,N_16863);
and U17346 (N_17346,N_16804,N_16684);
nand U17347 (N_17347,N_16926,N_16613);
nand U17348 (N_17348,N_16896,N_16988);
nand U17349 (N_17349,N_16670,N_16718);
nand U17350 (N_17350,N_16784,N_16637);
xnor U17351 (N_17351,N_16735,N_16647);
nor U17352 (N_17352,N_16895,N_16670);
xor U17353 (N_17353,N_16618,N_16874);
and U17354 (N_17354,N_16530,N_16888);
xnor U17355 (N_17355,N_16836,N_16537);
nor U17356 (N_17356,N_16501,N_16787);
and U17357 (N_17357,N_16831,N_16864);
xnor U17358 (N_17358,N_16862,N_16949);
or U17359 (N_17359,N_16984,N_16648);
xnor U17360 (N_17360,N_16522,N_16824);
nand U17361 (N_17361,N_16609,N_16624);
and U17362 (N_17362,N_16585,N_16922);
and U17363 (N_17363,N_16973,N_16764);
or U17364 (N_17364,N_16581,N_16788);
nand U17365 (N_17365,N_16931,N_16677);
xnor U17366 (N_17366,N_16914,N_16625);
xor U17367 (N_17367,N_16632,N_16552);
and U17368 (N_17368,N_16504,N_16971);
and U17369 (N_17369,N_16624,N_16560);
nor U17370 (N_17370,N_16799,N_16638);
nand U17371 (N_17371,N_16807,N_16547);
and U17372 (N_17372,N_16838,N_16644);
nor U17373 (N_17373,N_16788,N_16806);
or U17374 (N_17374,N_16833,N_16712);
xnor U17375 (N_17375,N_16774,N_16925);
nor U17376 (N_17376,N_16557,N_16870);
and U17377 (N_17377,N_16769,N_16688);
and U17378 (N_17378,N_16554,N_16582);
xor U17379 (N_17379,N_16748,N_16607);
or U17380 (N_17380,N_16618,N_16763);
and U17381 (N_17381,N_16997,N_16595);
nor U17382 (N_17382,N_16705,N_16725);
nand U17383 (N_17383,N_16530,N_16821);
nor U17384 (N_17384,N_16655,N_16862);
or U17385 (N_17385,N_16602,N_16578);
xnor U17386 (N_17386,N_16874,N_16980);
nor U17387 (N_17387,N_16991,N_16788);
nor U17388 (N_17388,N_16548,N_16788);
and U17389 (N_17389,N_16856,N_16909);
nand U17390 (N_17390,N_16615,N_16972);
nor U17391 (N_17391,N_16701,N_16823);
nand U17392 (N_17392,N_16692,N_16820);
nand U17393 (N_17393,N_16761,N_16644);
nor U17394 (N_17394,N_16618,N_16775);
nand U17395 (N_17395,N_16864,N_16905);
nor U17396 (N_17396,N_16986,N_16767);
xnor U17397 (N_17397,N_16521,N_16919);
xnor U17398 (N_17398,N_16716,N_16758);
or U17399 (N_17399,N_16831,N_16899);
or U17400 (N_17400,N_16957,N_16700);
nand U17401 (N_17401,N_16965,N_16524);
nand U17402 (N_17402,N_16553,N_16717);
and U17403 (N_17403,N_16883,N_16907);
nor U17404 (N_17404,N_16525,N_16585);
and U17405 (N_17405,N_16811,N_16636);
xor U17406 (N_17406,N_16822,N_16552);
nand U17407 (N_17407,N_16694,N_16868);
nor U17408 (N_17408,N_16754,N_16666);
nor U17409 (N_17409,N_16777,N_16904);
or U17410 (N_17410,N_16789,N_16739);
xor U17411 (N_17411,N_16581,N_16991);
or U17412 (N_17412,N_16515,N_16980);
nand U17413 (N_17413,N_16664,N_16755);
or U17414 (N_17414,N_16886,N_16654);
or U17415 (N_17415,N_16799,N_16867);
xor U17416 (N_17416,N_16760,N_16618);
nor U17417 (N_17417,N_16769,N_16870);
or U17418 (N_17418,N_16755,N_16579);
nand U17419 (N_17419,N_16637,N_16628);
and U17420 (N_17420,N_16803,N_16993);
xor U17421 (N_17421,N_16646,N_16991);
or U17422 (N_17422,N_16925,N_16760);
and U17423 (N_17423,N_16875,N_16903);
and U17424 (N_17424,N_16861,N_16814);
or U17425 (N_17425,N_16705,N_16962);
and U17426 (N_17426,N_16694,N_16776);
nand U17427 (N_17427,N_16556,N_16530);
nand U17428 (N_17428,N_16868,N_16726);
and U17429 (N_17429,N_16633,N_16927);
and U17430 (N_17430,N_16974,N_16911);
and U17431 (N_17431,N_16652,N_16862);
xor U17432 (N_17432,N_16842,N_16938);
or U17433 (N_17433,N_16862,N_16821);
nor U17434 (N_17434,N_16701,N_16561);
and U17435 (N_17435,N_16937,N_16758);
xor U17436 (N_17436,N_16992,N_16912);
or U17437 (N_17437,N_16779,N_16510);
and U17438 (N_17438,N_16617,N_16906);
or U17439 (N_17439,N_16576,N_16742);
nor U17440 (N_17440,N_16579,N_16894);
or U17441 (N_17441,N_16598,N_16719);
or U17442 (N_17442,N_16998,N_16873);
xor U17443 (N_17443,N_16688,N_16985);
nor U17444 (N_17444,N_16628,N_16760);
nand U17445 (N_17445,N_16890,N_16670);
and U17446 (N_17446,N_16510,N_16728);
nor U17447 (N_17447,N_16809,N_16939);
xnor U17448 (N_17448,N_16647,N_16973);
and U17449 (N_17449,N_16555,N_16900);
xor U17450 (N_17450,N_16819,N_16751);
nand U17451 (N_17451,N_16736,N_16733);
nor U17452 (N_17452,N_16891,N_16615);
nor U17453 (N_17453,N_16829,N_16525);
nor U17454 (N_17454,N_16508,N_16931);
nand U17455 (N_17455,N_16700,N_16529);
xor U17456 (N_17456,N_16770,N_16549);
nor U17457 (N_17457,N_16648,N_16609);
nand U17458 (N_17458,N_16730,N_16510);
and U17459 (N_17459,N_16681,N_16911);
nand U17460 (N_17460,N_16767,N_16755);
or U17461 (N_17461,N_16737,N_16560);
nor U17462 (N_17462,N_16910,N_16821);
and U17463 (N_17463,N_16715,N_16620);
xor U17464 (N_17464,N_16709,N_16879);
xor U17465 (N_17465,N_16860,N_16798);
nor U17466 (N_17466,N_16682,N_16996);
and U17467 (N_17467,N_16579,N_16961);
xnor U17468 (N_17468,N_16933,N_16877);
nor U17469 (N_17469,N_16842,N_16682);
nand U17470 (N_17470,N_16806,N_16654);
nand U17471 (N_17471,N_16967,N_16922);
or U17472 (N_17472,N_16983,N_16998);
and U17473 (N_17473,N_16677,N_16744);
and U17474 (N_17474,N_16539,N_16935);
xnor U17475 (N_17475,N_16856,N_16560);
nand U17476 (N_17476,N_16948,N_16878);
nor U17477 (N_17477,N_16785,N_16602);
nand U17478 (N_17478,N_16865,N_16775);
or U17479 (N_17479,N_16710,N_16876);
or U17480 (N_17480,N_16757,N_16945);
and U17481 (N_17481,N_16774,N_16928);
or U17482 (N_17482,N_16545,N_16871);
or U17483 (N_17483,N_16516,N_16806);
nor U17484 (N_17484,N_16896,N_16728);
or U17485 (N_17485,N_16878,N_16906);
xor U17486 (N_17486,N_16848,N_16872);
nand U17487 (N_17487,N_16620,N_16774);
nand U17488 (N_17488,N_16813,N_16650);
nand U17489 (N_17489,N_16937,N_16571);
xor U17490 (N_17490,N_16933,N_16873);
and U17491 (N_17491,N_16819,N_16873);
and U17492 (N_17492,N_16542,N_16948);
or U17493 (N_17493,N_16573,N_16773);
and U17494 (N_17494,N_16978,N_16575);
nor U17495 (N_17495,N_16778,N_16896);
nor U17496 (N_17496,N_16668,N_16535);
and U17497 (N_17497,N_16960,N_16861);
and U17498 (N_17498,N_16923,N_16989);
nand U17499 (N_17499,N_16994,N_16676);
and U17500 (N_17500,N_17465,N_17177);
nand U17501 (N_17501,N_17195,N_17227);
and U17502 (N_17502,N_17176,N_17114);
nor U17503 (N_17503,N_17228,N_17394);
or U17504 (N_17504,N_17271,N_17382);
nor U17505 (N_17505,N_17373,N_17010);
nor U17506 (N_17506,N_17357,N_17030);
xnor U17507 (N_17507,N_17398,N_17341);
or U17508 (N_17508,N_17024,N_17063);
xnor U17509 (N_17509,N_17043,N_17081);
and U17510 (N_17510,N_17255,N_17348);
xor U17511 (N_17511,N_17250,N_17276);
nor U17512 (N_17512,N_17131,N_17327);
and U17513 (N_17513,N_17069,N_17455);
xor U17514 (N_17514,N_17428,N_17111);
or U17515 (N_17515,N_17236,N_17193);
nand U17516 (N_17516,N_17129,N_17481);
and U17517 (N_17517,N_17226,N_17256);
or U17518 (N_17518,N_17216,N_17174);
or U17519 (N_17519,N_17007,N_17196);
xnor U17520 (N_17520,N_17170,N_17393);
nand U17521 (N_17521,N_17082,N_17208);
and U17522 (N_17522,N_17288,N_17108);
xnor U17523 (N_17523,N_17380,N_17054);
or U17524 (N_17524,N_17060,N_17378);
and U17525 (N_17525,N_17138,N_17302);
xnor U17526 (N_17526,N_17212,N_17299);
nand U17527 (N_17527,N_17312,N_17166);
nor U17528 (N_17528,N_17157,N_17161);
nand U17529 (N_17529,N_17261,N_17223);
xor U17530 (N_17530,N_17353,N_17339);
nor U17531 (N_17531,N_17077,N_17301);
or U17532 (N_17532,N_17427,N_17396);
xor U17533 (N_17533,N_17025,N_17445);
nand U17534 (N_17534,N_17416,N_17337);
nand U17535 (N_17535,N_17232,N_17184);
or U17536 (N_17536,N_17233,N_17057);
and U17537 (N_17537,N_17061,N_17038);
and U17538 (N_17538,N_17086,N_17046);
xor U17539 (N_17539,N_17135,N_17376);
nand U17540 (N_17540,N_17149,N_17004);
or U17541 (N_17541,N_17031,N_17207);
nor U17542 (N_17542,N_17485,N_17359);
xnor U17543 (N_17543,N_17486,N_17005);
and U17544 (N_17544,N_17319,N_17065);
nand U17545 (N_17545,N_17464,N_17365);
nor U17546 (N_17546,N_17266,N_17286);
nor U17547 (N_17547,N_17009,N_17355);
nor U17548 (N_17548,N_17461,N_17080);
xnor U17549 (N_17549,N_17214,N_17423);
nand U17550 (N_17550,N_17285,N_17435);
xnor U17551 (N_17551,N_17265,N_17039);
xnor U17552 (N_17552,N_17473,N_17167);
nor U17553 (N_17553,N_17493,N_17400);
xor U17554 (N_17554,N_17076,N_17451);
nand U17555 (N_17555,N_17370,N_17338);
nand U17556 (N_17556,N_17156,N_17071);
nor U17557 (N_17557,N_17075,N_17412);
and U17558 (N_17558,N_17342,N_17397);
and U17559 (N_17559,N_17107,N_17418);
or U17560 (N_17560,N_17016,N_17254);
nand U17561 (N_17561,N_17383,N_17122);
nor U17562 (N_17562,N_17048,N_17127);
nor U17563 (N_17563,N_17116,N_17333);
nand U17564 (N_17564,N_17309,N_17409);
nand U17565 (N_17565,N_17124,N_17316);
or U17566 (N_17566,N_17109,N_17320);
nor U17567 (N_17567,N_17387,N_17126);
xor U17568 (N_17568,N_17115,N_17173);
and U17569 (N_17569,N_17282,N_17033);
nand U17570 (N_17570,N_17117,N_17251);
nor U17571 (N_17571,N_17145,N_17438);
xor U17572 (N_17572,N_17499,N_17148);
xor U17573 (N_17573,N_17392,N_17460);
and U17574 (N_17574,N_17183,N_17186);
xor U17575 (N_17575,N_17289,N_17110);
nand U17576 (N_17576,N_17091,N_17468);
and U17577 (N_17577,N_17487,N_17344);
xor U17578 (N_17578,N_17347,N_17123);
or U17579 (N_17579,N_17273,N_17308);
or U17580 (N_17580,N_17495,N_17277);
nand U17581 (N_17581,N_17477,N_17225);
nand U17582 (N_17582,N_17315,N_17034);
nand U17583 (N_17583,N_17022,N_17243);
and U17584 (N_17584,N_17420,N_17128);
nor U17585 (N_17585,N_17200,N_17492);
and U17586 (N_17586,N_17087,N_17406);
nor U17587 (N_17587,N_17484,N_17047);
or U17588 (N_17588,N_17346,N_17084);
nand U17589 (N_17589,N_17479,N_17472);
nand U17590 (N_17590,N_17475,N_17293);
nor U17591 (N_17591,N_17152,N_17379);
nor U17592 (N_17592,N_17402,N_17326);
nor U17593 (N_17593,N_17407,N_17112);
or U17594 (N_17594,N_17074,N_17163);
and U17595 (N_17595,N_17323,N_17313);
nand U17596 (N_17596,N_17272,N_17137);
nand U17597 (N_17597,N_17280,N_17098);
nor U17598 (N_17598,N_17015,N_17292);
nor U17599 (N_17599,N_17300,N_17188);
and U17600 (N_17600,N_17494,N_17062);
and U17601 (N_17601,N_17147,N_17028);
xor U17602 (N_17602,N_17011,N_17281);
and U17603 (N_17603,N_17369,N_17044);
and U17604 (N_17604,N_17229,N_17066);
xnor U17605 (N_17605,N_17260,N_17410);
nor U17606 (N_17606,N_17432,N_17317);
nor U17607 (N_17607,N_17310,N_17203);
and U17608 (N_17608,N_17095,N_17390);
nor U17609 (N_17609,N_17434,N_17252);
and U17610 (N_17610,N_17142,N_17458);
and U17611 (N_17611,N_17205,N_17073);
nand U17612 (N_17612,N_17118,N_17094);
xnor U17613 (N_17613,N_17377,N_17097);
nor U17614 (N_17614,N_17498,N_17058);
nand U17615 (N_17615,N_17431,N_17235);
and U17616 (N_17616,N_17325,N_17204);
nand U17617 (N_17617,N_17399,N_17248);
nand U17618 (N_17618,N_17102,N_17388);
xor U17619 (N_17619,N_17478,N_17191);
or U17620 (N_17620,N_17245,N_17335);
xnor U17621 (N_17621,N_17329,N_17153);
or U17622 (N_17622,N_17303,N_17106);
or U17623 (N_17623,N_17351,N_17017);
or U17624 (N_17624,N_17356,N_17125);
xor U17625 (N_17625,N_17040,N_17422);
or U17626 (N_17626,N_17158,N_17140);
nor U17627 (N_17627,N_17291,N_17162);
and U17628 (N_17628,N_17104,N_17314);
nand U17629 (N_17629,N_17070,N_17413);
or U17630 (N_17630,N_17072,N_17417);
and U17631 (N_17631,N_17194,N_17491);
or U17632 (N_17632,N_17018,N_17241);
or U17633 (N_17633,N_17036,N_17381);
nor U17634 (N_17634,N_17113,N_17059);
xor U17635 (N_17635,N_17429,N_17056);
and U17636 (N_17636,N_17470,N_17083);
xnor U17637 (N_17637,N_17283,N_17463);
xor U17638 (N_17638,N_17437,N_17467);
xor U17639 (N_17639,N_17295,N_17322);
nor U17640 (N_17640,N_17363,N_17278);
nor U17641 (N_17641,N_17002,N_17190);
nand U17642 (N_17642,N_17426,N_17234);
nand U17643 (N_17643,N_17192,N_17055);
and U17644 (N_17644,N_17441,N_17297);
xnor U17645 (N_17645,N_17240,N_17414);
nand U17646 (N_17646,N_17332,N_17134);
nor U17647 (N_17647,N_17103,N_17244);
or U17648 (N_17648,N_17405,N_17480);
or U17649 (N_17649,N_17143,N_17222);
or U17650 (N_17650,N_17328,N_17202);
nand U17651 (N_17651,N_17362,N_17476);
or U17652 (N_17652,N_17318,N_17268);
nor U17653 (N_17653,N_17052,N_17237);
and U17654 (N_17654,N_17139,N_17389);
or U17655 (N_17655,N_17171,N_17012);
nor U17656 (N_17656,N_17199,N_17053);
nor U17657 (N_17657,N_17133,N_17321);
xnor U17658 (N_17658,N_17466,N_17239);
nand U17659 (N_17659,N_17224,N_17275);
xor U17660 (N_17660,N_17221,N_17085);
nor U17661 (N_17661,N_17021,N_17185);
nor U17662 (N_17662,N_17041,N_17096);
xnor U17663 (N_17663,N_17258,N_17067);
or U17664 (N_17664,N_17154,N_17037);
nor U17665 (N_17665,N_17456,N_17014);
xor U17666 (N_17666,N_17311,N_17403);
nor U17667 (N_17667,N_17367,N_17262);
and U17668 (N_17668,N_17349,N_17415);
nand U17669 (N_17669,N_17159,N_17064);
xnor U17670 (N_17670,N_17209,N_17386);
and U17671 (N_17671,N_17187,N_17092);
xor U17672 (N_17672,N_17454,N_17408);
and U17673 (N_17673,N_17179,N_17334);
xor U17674 (N_17674,N_17001,N_17459);
xnor U17675 (N_17675,N_17345,N_17247);
or U17676 (N_17676,N_17453,N_17093);
xnor U17677 (N_17677,N_17264,N_17090);
nand U17678 (N_17678,N_17100,N_17457);
xor U17679 (N_17679,N_17197,N_17385);
or U17680 (N_17680,N_17160,N_17439);
nor U17681 (N_17681,N_17136,N_17462);
nor U17682 (N_17682,N_17032,N_17105);
nand U17683 (N_17683,N_17471,N_17088);
and U17684 (N_17684,N_17249,N_17444);
nor U17685 (N_17685,N_17121,N_17217);
nor U17686 (N_17686,N_17364,N_17488);
and U17687 (N_17687,N_17290,N_17401);
xor U17688 (N_17688,N_17068,N_17284);
and U17689 (N_17689,N_17331,N_17433);
nor U17690 (N_17690,N_17482,N_17474);
and U17691 (N_17691,N_17340,N_17099);
nor U17692 (N_17692,N_17026,N_17042);
nor U17693 (N_17693,N_17452,N_17440);
xnor U17694 (N_17694,N_17242,N_17371);
and U17695 (N_17695,N_17330,N_17307);
and U17696 (N_17696,N_17490,N_17019);
or U17697 (N_17697,N_17424,N_17013);
or U17698 (N_17698,N_17425,N_17172);
nand U17699 (N_17699,N_17219,N_17051);
xnor U17700 (N_17700,N_17175,N_17220);
nand U17701 (N_17701,N_17375,N_17469);
nor U17702 (N_17702,N_17050,N_17336);
and U17703 (N_17703,N_17215,N_17384);
nor U17704 (N_17704,N_17180,N_17287);
xor U17705 (N_17705,N_17049,N_17035);
nand U17706 (N_17706,N_17360,N_17029);
nand U17707 (N_17707,N_17449,N_17201);
nor U17708 (N_17708,N_17446,N_17213);
nor U17709 (N_17709,N_17189,N_17366);
nand U17710 (N_17710,N_17489,N_17298);
or U17711 (N_17711,N_17274,N_17436);
and U17712 (N_17712,N_17497,N_17000);
or U17713 (N_17713,N_17305,N_17150);
and U17714 (N_17714,N_17101,N_17404);
or U17715 (N_17715,N_17246,N_17132);
nor U17716 (N_17716,N_17395,N_17020);
nand U17717 (N_17717,N_17164,N_17206);
or U17718 (N_17718,N_17294,N_17198);
xor U17719 (N_17719,N_17391,N_17210);
or U17720 (N_17720,N_17006,N_17144);
or U17721 (N_17721,N_17231,N_17419);
and U17722 (N_17722,N_17304,N_17448);
or U17723 (N_17723,N_17306,N_17211);
and U17724 (N_17724,N_17181,N_17270);
xor U17725 (N_17725,N_17008,N_17141);
or U17726 (N_17726,N_17257,N_17259);
xor U17727 (N_17727,N_17023,N_17182);
nor U17728 (N_17728,N_17421,N_17269);
xor U17729 (N_17729,N_17146,N_17442);
nand U17730 (N_17730,N_17169,N_17003);
nand U17731 (N_17731,N_17483,N_17151);
xnor U17732 (N_17732,N_17165,N_17263);
xnor U17733 (N_17733,N_17350,N_17296);
nor U17734 (N_17734,N_17411,N_17324);
nor U17735 (N_17735,N_17238,N_17374);
xnor U17736 (N_17736,N_17352,N_17089);
xor U17737 (N_17737,N_17078,N_17430);
nand U17738 (N_17738,N_17358,N_17178);
and U17739 (N_17739,N_17079,N_17343);
and U17740 (N_17740,N_17361,N_17368);
nand U17741 (N_17741,N_17443,N_17027);
and U17742 (N_17742,N_17450,N_17168);
xnor U17743 (N_17743,N_17120,N_17279);
nand U17744 (N_17744,N_17155,N_17253);
or U17745 (N_17745,N_17218,N_17354);
and U17746 (N_17746,N_17045,N_17372);
xnor U17747 (N_17747,N_17447,N_17130);
and U17748 (N_17748,N_17230,N_17267);
nand U17749 (N_17749,N_17119,N_17496);
and U17750 (N_17750,N_17334,N_17126);
or U17751 (N_17751,N_17005,N_17464);
or U17752 (N_17752,N_17068,N_17372);
or U17753 (N_17753,N_17473,N_17213);
and U17754 (N_17754,N_17413,N_17353);
and U17755 (N_17755,N_17267,N_17146);
nand U17756 (N_17756,N_17130,N_17494);
xnor U17757 (N_17757,N_17280,N_17449);
nand U17758 (N_17758,N_17010,N_17424);
nor U17759 (N_17759,N_17143,N_17253);
xnor U17760 (N_17760,N_17370,N_17161);
nor U17761 (N_17761,N_17370,N_17201);
and U17762 (N_17762,N_17235,N_17383);
and U17763 (N_17763,N_17303,N_17250);
and U17764 (N_17764,N_17340,N_17488);
and U17765 (N_17765,N_17453,N_17472);
nor U17766 (N_17766,N_17423,N_17339);
or U17767 (N_17767,N_17137,N_17186);
nor U17768 (N_17768,N_17189,N_17348);
and U17769 (N_17769,N_17408,N_17099);
nand U17770 (N_17770,N_17025,N_17437);
or U17771 (N_17771,N_17182,N_17405);
or U17772 (N_17772,N_17131,N_17494);
nand U17773 (N_17773,N_17479,N_17000);
nand U17774 (N_17774,N_17355,N_17249);
xnor U17775 (N_17775,N_17123,N_17288);
or U17776 (N_17776,N_17459,N_17177);
nor U17777 (N_17777,N_17401,N_17166);
nor U17778 (N_17778,N_17063,N_17157);
nor U17779 (N_17779,N_17369,N_17088);
nor U17780 (N_17780,N_17044,N_17440);
xor U17781 (N_17781,N_17142,N_17413);
and U17782 (N_17782,N_17343,N_17418);
or U17783 (N_17783,N_17039,N_17027);
nor U17784 (N_17784,N_17302,N_17441);
or U17785 (N_17785,N_17369,N_17216);
xnor U17786 (N_17786,N_17068,N_17219);
nor U17787 (N_17787,N_17256,N_17143);
xor U17788 (N_17788,N_17238,N_17203);
and U17789 (N_17789,N_17318,N_17363);
and U17790 (N_17790,N_17114,N_17430);
nor U17791 (N_17791,N_17127,N_17350);
and U17792 (N_17792,N_17322,N_17477);
xnor U17793 (N_17793,N_17205,N_17432);
or U17794 (N_17794,N_17312,N_17081);
nand U17795 (N_17795,N_17279,N_17357);
nand U17796 (N_17796,N_17481,N_17399);
nand U17797 (N_17797,N_17315,N_17383);
or U17798 (N_17798,N_17144,N_17107);
nor U17799 (N_17799,N_17158,N_17237);
nor U17800 (N_17800,N_17264,N_17359);
nor U17801 (N_17801,N_17177,N_17021);
nand U17802 (N_17802,N_17240,N_17068);
xnor U17803 (N_17803,N_17497,N_17274);
xnor U17804 (N_17804,N_17014,N_17001);
xor U17805 (N_17805,N_17285,N_17143);
nor U17806 (N_17806,N_17221,N_17484);
xnor U17807 (N_17807,N_17231,N_17216);
and U17808 (N_17808,N_17214,N_17422);
nor U17809 (N_17809,N_17454,N_17182);
or U17810 (N_17810,N_17289,N_17311);
xor U17811 (N_17811,N_17478,N_17245);
nand U17812 (N_17812,N_17045,N_17240);
xor U17813 (N_17813,N_17492,N_17211);
nand U17814 (N_17814,N_17198,N_17494);
or U17815 (N_17815,N_17292,N_17107);
or U17816 (N_17816,N_17458,N_17012);
and U17817 (N_17817,N_17021,N_17402);
nor U17818 (N_17818,N_17297,N_17012);
or U17819 (N_17819,N_17354,N_17289);
xor U17820 (N_17820,N_17408,N_17488);
or U17821 (N_17821,N_17438,N_17070);
xnor U17822 (N_17822,N_17202,N_17082);
and U17823 (N_17823,N_17040,N_17093);
or U17824 (N_17824,N_17367,N_17164);
or U17825 (N_17825,N_17152,N_17338);
and U17826 (N_17826,N_17042,N_17040);
or U17827 (N_17827,N_17137,N_17187);
xor U17828 (N_17828,N_17197,N_17283);
nand U17829 (N_17829,N_17216,N_17271);
nor U17830 (N_17830,N_17179,N_17294);
and U17831 (N_17831,N_17041,N_17167);
nor U17832 (N_17832,N_17109,N_17421);
xor U17833 (N_17833,N_17095,N_17205);
and U17834 (N_17834,N_17387,N_17055);
and U17835 (N_17835,N_17479,N_17054);
or U17836 (N_17836,N_17216,N_17361);
or U17837 (N_17837,N_17035,N_17493);
nand U17838 (N_17838,N_17140,N_17471);
and U17839 (N_17839,N_17328,N_17166);
and U17840 (N_17840,N_17105,N_17135);
or U17841 (N_17841,N_17010,N_17136);
or U17842 (N_17842,N_17014,N_17443);
xor U17843 (N_17843,N_17244,N_17196);
or U17844 (N_17844,N_17053,N_17437);
nand U17845 (N_17845,N_17438,N_17051);
and U17846 (N_17846,N_17205,N_17101);
nor U17847 (N_17847,N_17373,N_17074);
or U17848 (N_17848,N_17036,N_17300);
nor U17849 (N_17849,N_17352,N_17159);
and U17850 (N_17850,N_17225,N_17492);
or U17851 (N_17851,N_17393,N_17139);
and U17852 (N_17852,N_17207,N_17210);
or U17853 (N_17853,N_17134,N_17461);
nor U17854 (N_17854,N_17405,N_17104);
and U17855 (N_17855,N_17057,N_17331);
xor U17856 (N_17856,N_17009,N_17440);
nand U17857 (N_17857,N_17328,N_17027);
nand U17858 (N_17858,N_17081,N_17259);
xnor U17859 (N_17859,N_17174,N_17400);
and U17860 (N_17860,N_17382,N_17428);
nand U17861 (N_17861,N_17157,N_17151);
and U17862 (N_17862,N_17161,N_17432);
and U17863 (N_17863,N_17187,N_17001);
or U17864 (N_17864,N_17233,N_17362);
and U17865 (N_17865,N_17206,N_17301);
xor U17866 (N_17866,N_17171,N_17394);
nand U17867 (N_17867,N_17053,N_17141);
nor U17868 (N_17868,N_17304,N_17314);
and U17869 (N_17869,N_17343,N_17372);
nand U17870 (N_17870,N_17419,N_17185);
and U17871 (N_17871,N_17119,N_17382);
xnor U17872 (N_17872,N_17000,N_17491);
nand U17873 (N_17873,N_17283,N_17467);
xor U17874 (N_17874,N_17480,N_17482);
xnor U17875 (N_17875,N_17415,N_17437);
or U17876 (N_17876,N_17225,N_17033);
or U17877 (N_17877,N_17195,N_17229);
or U17878 (N_17878,N_17126,N_17273);
or U17879 (N_17879,N_17374,N_17132);
nand U17880 (N_17880,N_17412,N_17114);
and U17881 (N_17881,N_17120,N_17409);
nor U17882 (N_17882,N_17276,N_17427);
and U17883 (N_17883,N_17408,N_17195);
nor U17884 (N_17884,N_17216,N_17099);
xor U17885 (N_17885,N_17302,N_17391);
nand U17886 (N_17886,N_17324,N_17368);
or U17887 (N_17887,N_17160,N_17206);
xnor U17888 (N_17888,N_17100,N_17294);
nand U17889 (N_17889,N_17024,N_17000);
or U17890 (N_17890,N_17189,N_17283);
or U17891 (N_17891,N_17023,N_17492);
nand U17892 (N_17892,N_17391,N_17371);
nand U17893 (N_17893,N_17294,N_17024);
and U17894 (N_17894,N_17207,N_17320);
or U17895 (N_17895,N_17289,N_17286);
nand U17896 (N_17896,N_17110,N_17054);
nor U17897 (N_17897,N_17223,N_17032);
xnor U17898 (N_17898,N_17329,N_17350);
nor U17899 (N_17899,N_17440,N_17194);
xnor U17900 (N_17900,N_17154,N_17444);
and U17901 (N_17901,N_17442,N_17262);
and U17902 (N_17902,N_17123,N_17318);
nand U17903 (N_17903,N_17322,N_17124);
nor U17904 (N_17904,N_17403,N_17446);
and U17905 (N_17905,N_17119,N_17459);
and U17906 (N_17906,N_17395,N_17233);
or U17907 (N_17907,N_17149,N_17257);
and U17908 (N_17908,N_17372,N_17266);
nor U17909 (N_17909,N_17168,N_17251);
or U17910 (N_17910,N_17388,N_17216);
or U17911 (N_17911,N_17062,N_17418);
nor U17912 (N_17912,N_17331,N_17093);
and U17913 (N_17913,N_17260,N_17342);
and U17914 (N_17914,N_17300,N_17242);
nand U17915 (N_17915,N_17345,N_17092);
nor U17916 (N_17916,N_17206,N_17201);
and U17917 (N_17917,N_17445,N_17299);
nand U17918 (N_17918,N_17231,N_17009);
and U17919 (N_17919,N_17093,N_17259);
nor U17920 (N_17920,N_17334,N_17473);
xnor U17921 (N_17921,N_17162,N_17295);
and U17922 (N_17922,N_17187,N_17053);
nor U17923 (N_17923,N_17173,N_17276);
or U17924 (N_17924,N_17346,N_17091);
and U17925 (N_17925,N_17444,N_17399);
xnor U17926 (N_17926,N_17400,N_17484);
nand U17927 (N_17927,N_17079,N_17325);
and U17928 (N_17928,N_17313,N_17192);
and U17929 (N_17929,N_17423,N_17120);
nand U17930 (N_17930,N_17474,N_17339);
and U17931 (N_17931,N_17093,N_17176);
nand U17932 (N_17932,N_17488,N_17076);
or U17933 (N_17933,N_17402,N_17096);
xor U17934 (N_17934,N_17027,N_17296);
xnor U17935 (N_17935,N_17007,N_17194);
nand U17936 (N_17936,N_17436,N_17496);
xnor U17937 (N_17937,N_17235,N_17294);
or U17938 (N_17938,N_17001,N_17097);
nor U17939 (N_17939,N_17236,N_17341);
nand U17940 (N_17940,N_17322,N_17060);
nor U17941 (N_17941,N_17158,N_17115);
nor U17942 (N_17942,N_17084,N_17206);
nand U17943 (N_17943,N_17215,N_17083);
nor U17944 (N_17944,N_17046,N_17281);
or U17945 (N_17945,N_17231,N_17182);
or U17946 (N_17946,N_17477,N_17312);
nor U17947 (N_17947,N_17458,N_17468);
nand U17948 (N_17948,N_17214,N_17094);
nor U17949 (N_17949,N_17430,N_17459);
and U17950 (N_17950,N_17076,N_17345);
nand U17951 (N_17951,N_17337,N_17237);
and U17952 (N_17952,N_17195,N_17224);
or U17953 (N_17953,N_17341,N_17390);
or U17954 (N_17954,N_17415,N_17441);
nand U17955 (N_17955,N_17122,N_17278);
or U17956 (N_17956,N_17200,N_17160);
nor U17957 (N_17957,N_17167,N_17026);
nand U17958 (N_17958,N_17063,N_17356);
nor U17959 (N_17959,N_17407,N_17169);
and U17960 (N_17960,N_17406,N_17477);
nor U17961 (N_17961,N_17247,N_17277);
or U17962 (N_17962,N_17298,N_17090);
or U17963 (N_17963,N_17114,N_17034);
or U17964 (N_17964,N_17336,N_17267);
nand U17965 (N_17965,N_17083,N_17411);
nor U17966 (N_17966,N_17325,N_17064);
xor U17967 (N_17967,N_17223,N_17409);
or U17968 (N_17968,N_17093,N_17092);
nand U17969 (N_17969,N_17076,N_17128);
xnor U17970 (N_17970,N_17241,N_17308);
xor U17971 (N_17971,N_17254,N_17223);
nand U17972 (N_17972,N_17377,N_17107);
nor U17973 (N_17973,N_17164,N_17305);
and U17974 (N_17974,N_17495,N_17331);
nor U17975 (N_17975,N_17162,N_17400);
nand U17976 (N_17976,N_17341,N_17308);
nor U17977 (N_17977,N_17429,N_17011);
and U17978 (N_17978,N_17102,N_17336);
xor U17979 (N_17979,N_17413,N_17056);
or U17980 (N_17980,N_17286,N_17332);
xor U17981 (N_17981,N_17101,N_17239);
nor U17982 (N_17982,N_17205,N_17142);
nor U17983 (N_17983,N_17136,N_17002);
and U17984 (N_17984,N_17142,N_17073);
or U17985 (N_17985,N_17451,N_17440);
nand U17986 (N_17986,N_17347,N_17362);
xnor U17987 (N_17987,N_17121,N_17392);
nor U17988 (N_17988,N_17238,N_17272);
nor U17989 (N_17989,N_17305,N_17436);
or U17990 (N_17990,N_17232,N_17057);
nand U17991 (N_17991,N_17407,N_17103);
nor U17992 (N_17992,N_17112,N_17221);
nand U17993 (N_17993,N_17493,N_17079);
nor U17994 (N_17994,N_17105,N_17294);
nand U17995 (N_17995,N_17247,N_17447);
nor U17996 (N_17996,N_17190,N_17486);
xnor U17997 (N_17997,N_17390,N_17013);
or U17998 (N_17998,N_17448,N_17274);
nor U17999 (N_17999,N_17098,N_17120);
or U18000 (N_18000,N_17834,N_17971);
xor U18001 (N_18001,N_17667,N_17908);
nor U18002 (N_18002,N_17552,N_17725);
nor U18003 (N_18003,N_17697,N_17679);
nand U18004 (N_18004,N_17519,N_17561);
or U18005 (N_18005,N_17629,N_17735);
and U18006 (N_18006,N_17965,N_17674);
nor U18007 (N_18007,N_17822,N_17938);
or U18008 (N_18008,N_17538,N_17878);
nand U18009 (N_18009,N_17956,N_17584);
nand U18010 (N_18010,N_17569,N_17568);
nor U18011 (N_18011,N_17779,N_17580);
or U18012 (N_18012,N_17591,N_17645);
and U18013 (N_18013,N_17719,N_17846);
and U18014 (N_18014,N_17879,N_17869);
nor U18015 (N_18015,N_17848,N_17778);
xor U18016 (N_18016,N_17880,N_17788);
xor U18017 (N_18017,N_17508,N_17939);
and U18018 (N_18018,N_17798,N_17505);
nor U18019 (N_18019,N_17644,N_17632);
xor U18020 (N_18020,N_17706,N_17922);
nand U18021 (N_18021,N_17600,N_17671);
or U18022 (N_18022,N_17795,N_17741);
and U18023 (N_18023,N_17703,N_17998);
nor U18024 (N_18024,N_17658,N_17889);
xor U18025 (N_18025,N_17883,N_17692);
or U18026 (N_18026,N_17736,N_17919);
nor U18027 (N_18027,N_17571,N_17760);
or U18028 (N_18028,N_17825,N_17770);
nand U18029 (N_18029,N_17663,N_17813);
or U18030 (N_18030,N_17817,N_17710);
nand U18031 (N_18031,N_17799,N_17759);
or U18032 (N_18032,N_17581,N_17729);
and U18033 (N_18033,N_17718,N_17689);
nand U18034 (N_18034,N_17946,N_17844);
and U18035 (N_18035,N_17756,N_17755);
or U18036 (N_18036,N_17690,N_17953);
nand U18037 (N_18037,N_17514,N_17651);
nor U18038 (N_18038,N_17738,N_17852);
nand U18039 (N_18039,N_17954,N_17827);
or U18040 (N_18040,N_17854,N_17959);
and U18041 (N_18041,N_17804,N_17583);
or U18042 (N_18042,N_17837,N_17542);
nand U18043 (N_18043,N_17579,N_17857);
nor U18044 (N_18044,N_17536,N_17979);
and U18045 (N_18045,N_17700,N_17960);
xor U18046 (N_18046,N_17557,N_17943);
nand U18047 (N_18047,N_17845,N_17626);
or U18048 (N_18048,N_17850,N_17596);
nand U18049 (N_18049,N_17944,N_17912);
or U18050 (N_18050,N_17859,N_17546);
nor U18051 (N_18051,N_17999,N_17726);
xnor U18052 (N_18052,N_17618,N_17665);
and U18053 (N_18053,N_17733,N_17945);
and U18054 (N_18054,N_17796,N_17649);
or U18055 (N_18055,N_17661,N_17809);
xnor U18056 (N_18056,N_17526,N_17819);
or U18057 (N_18057,N_17918,N_17709);
xnor U18058 (N_18058,N_17962,N_17957);
or U18059 (N_18059,N_17826,N_17533);
nand U18060 (N_18060,N_17717,N_17951);
and U18061 (N_18061,N_17550,N_17896);
or U18062 (N_18062,N_17720,N_17914);
nor U18063 (N_18063,N_17611,N_17517);
and U18064 (N_18064,N_17818,N_17592);
or U18065 (N_18065,N_17545,N_17680);
nor U18066 (N_18066,N_17868,N_17551);
nor U18067 (N_18067,N_17932,N_17976);
and U18068 (N_18068,N_17814,N_17807);
and U18069 (N_18069,N_17847,N_17750);
and U18070 (N_18070,N_17647,N_17802);
xnor U18071 (N_18071,N_17660,N_17572);
or U18072 (N_18072,N_17888,N_17636);
nor U18073 (N_18073,N_17547,N_17702);
or U18074 (N_18074,N_17686,N_17820);
xor U18075 (N_18075,N_17642,N_17881);
or U18076 (N_18076,N_17502,N_17673);
nand U18077 (N_18077,N_17753,N_17664);
or U18078 (N_18078,N_17531,N_17511);
nor U18079 (N_18079,N_17512,N_17603);
nor U18080 (N_18080,N_17929,N_17641);
and U18081 (N_18081,N_17593,N_17539);
nand U18082 (N_18082,N_17865,N_17899);
and U18083 (N_18083,N_17926,N_17566);
nor U18084 (N_18084,N_17993,N_17904);
xor U18085 (N_18085,N_17874,N_17556);
or U18086 (N_18086,N_17708,N_17563);
nor U18087 (N_18087,N_17500,N_17609);
nand U18088 (N_18088,N_17876,N_17935);
nand U18089 (N_18089,N_17801,N_17616);
xnor U18090 (N_18090,N_17861,N_17555);
and U18091 (N_18091,N_17964,N_17527);
or U18092 (N_18092,N_17737,N_17782);
and U18093 (N_18093,N_17521,N_17763);
and U18094 (N_18094,N_17675,N_17685);
nor U18095 (N_18095,N_17607,N_17676);
nand U18096 (N_18096,N_17585,N_17530);
nor U18097 (N_18097,N_17564,N_17775);
nor U18098 (N_18098,N_17875,N_17503);
xor U18099 (N_18099,N_17537,N_17604);
xnor U18100 (N_18100,N_17523,N_17828);
nand U18101 (N_18101,N_17842,N_17969);
nand U18102 (N_18102,N_17885,N_17507);
xor U18103 (N_18103,N_17748,N_17967);
nor U18104 (N_18104,N_17839,N_17501);
and U18105 (N_18105,N_17786,N_17829);
and U18106 (N_18106,N_17974,N_17921);
or U18107 (N_18107,N_17648,N_17744);
and U18108 (N_18108,N_17518,N_17713);
or U18109 (N_18109,N_17623,N_17723);
xor U18110 (N_18110,N_17890,N_17747);
nand U18111 (N_18111,N_17524,N_17942);
nor U18112 (N_18112,N_17949,N_17696);
and U18113 (N_18113,N_17906,N_17787);
nor U18114 (N_18114,N_17877,N_17586);
or U18115 (N_18115,N_17900,N_17994);
xnor U18116 (N_18116,N_17785,N_17646);
xor U18117 (N_18117,N_17529,N_17762);
xnor U18118 (N_18118,N_17833,N_17606);
xor U18119 (N_18119,N_17767,N_17996);
or U18120 (N_18120,N_17619,N_17990);
nand U18121 (N_18121,N_17892,N_17669);
nor U18122 (N_18122,N_17920,N_17821);
nand U18123 (N_18123,N_17522,N_17856);
xor U18124 (N_18124,N_17811,N_17727);
and U18125 (N_18125,N_17769,N_17554);
nand U18126 (N_18126,N_17650,N_17952);
nand U18127 (N_18127,N_17752,N_17652);
nand U18128 (N_18128,N_17950,N_17862);
xnor U18129 (N_18129,N_17984,N_17602);
nor U18130 (N_18130,N_17955,N_17764);
xnor U18131 (N_18131,N_17504,N_17815);
xnor U18132 (N_18132,N_17622,N_17902);
or U18133 (N_18133,N_17858,N_17631);
or U18134 (N_18134,N_17575,N_17608);
nor U18135 (N_18135,N_17614,N_17630);
xor U18136 (N_18136,N_17758,N_17863);
nand U18137 (N_18137,N_17525,N_17958);
nor U18138 (N_18138,N_17528,N_17831);
or U18139 (N_18139,N_17541,N_17615);
nor U18140 (N_18140,N_17988,N_17898);
nor U18141 (N_18141,N_17694,N_17768);
and U18142 (N_18142,N_17633,N_17610);
and U18143 (N_18143,N_17670,N_17937);
nor U18144 (N_18144,N_17916,N_17698);
xnor U18145 (N_18145,N_17684,N_17800);
or U18146 (N_18146,N_17903,N_17659);
xnor U18147 (N_18147,N_17925,N_17978);
xnor U18148 (N_18148,N_17757,N_17995);
nand U18149 (N_18149,N_17510,N_17792);
or U18150 (N_18150,N_17662,N_17816);
nand U18151 (N_18151,N_17980,N_17989);
nand U18152 (N_18152,N_17628,N_17695);
and U18153 (N_18153,N_17621,N_17516);
or U18154 (N_18154,N_17771,N_17715);
xor U18155 (N_18155,N_17884,N_17655);
xnor U18156 (N_18156,N_17617,N_17506);
and U18157 (N_18157,N_17843,N_17640);
nand U18158 (N_18158,N_17761,N_17987);
xor U18159 (N_18159,N_17893,N_17543);
and U18160 (N_18160,N_17553,N_17866);
nand U18161 (N_18161,N_17559,N_17509);
and U18162 (N_18162,N_17936,N_17578);
or U18163 (N_18163,N_17928,N_17535);
nor U18164 (N_18164,N_17605,N_17751);
and U18165 (N_18165,N_17982,N_17595);
nor U18166 (N_18166,N_17773,N_17794);
or U18167 (N_18167,N_17823,N_17907);
or U18168 (N_18168,N_17643,N_17520);
and U18169 (N_18169,N_17532,N_17840);
xnor U18170 (N_18170,N_17743,N_17793);
xor U18171 (N_18171,N_17590,N_17613);
nor U18172 (N_18172,N_17891,N_17886);
nand U18173 (N_18173,N_17849,N_17991);
nand U18174 (N_18174,N_17887,N_17997);
nor U18175 (N_18175,N_17961,N_17594);
nor U18176 (N_18176,N_17973,N_17625);
and U18177 (N_18177,N_17797,N_17732);
and U18178 (N_18178,N_17772,N_17734);
and U18179 (N_18179,N_17704,N_17765);
or U18180 (N_18180,N_17812,N_17707);
or U18181 (N_18181,N_17774,N_17599);
nand U18182 (N_18182,N_17573,N_17992);
and U18183 (N_18183,N_17851,N_17927);
or U18184 (N_18184,N_17913,N_17784);
xnor U18185 (N_18185,N_17860,N_17940);
nand U18186 (N_18186,N_17540,N_17570);
and U18187 (N_18187,N_17634,N_17567);
or U18188 (N_18188,N_17931,N_17830);
xnor U18189 (N_18189,N_17588,N_17832);
nor U18190 (N_18190,N_17597,N_17871);
or U18191 (N_18191,N_17972,N_17612);
nor U18192 (N_18192,N_17601,N_17565);
or U18193 (N_18193,N_17678,N_17677);
and U18194 (N_18194,N_17699,N_17970);
nand U18195 (N_18195,N_17742,N_17790);
nor U18196 (N_18196,N_17560,N_17895);
xor U18197 (N_18197,N_17824,N_17911);
nor U18198 (N_18198,N_17745,N_17534);
and U18199 (N_18199,N_17910,N_17808);
nand U18200 (N_18200,N_17882,N_17855);
or U18201 (N_18201,N_17909,N_17688);
or U18202 (N_18202,N_17730,N_17924);
nor U18203 (N_18203,N_17835,N_17836);
nor U18204 (N_18204,N_17934,N_17624);
and U18205 (N_18205,N_17985,N_17805);
nor U18206 (N_18206,N_17791,N_17754);
and U18207 (N_18207,N_17986,N_17653);
or U18208 (N_18208,N_17682,N_17873);
or U18209 (N_18209,N_17687,N_17666);
nor U18210 (N_18210,N_17716,N_17576);
nand U18211 (N_18211,N_17963,N_17766);
nor U18212 (N_18212,N_17574,N_17975);
nand U18213 (N_18213,N_17724,N_17701);
nor U18214 (N_18214,N_17668,N_17905);
or U18215 (N_18215,N_17683,N_17721);
nor U18216 (N_18216,N_17712,N_17513);
xor U18217 (N_18217,N_17941,N_17549);
or U18218 (N_18218,N_17598,N_17948);
nor U18219 (N_18219,N_17639,N_17981);
nor U18220 (N_18220,N_17853,N_17587);
or U18221 (N_18221,N_17872,N_17637);
and U18222 (N_18222,N_17806,N_17722);
or U18223 (N_18223,N_17544,N_17966);
and U18224 (N_18224,N_17562,N_17776);
nand U18225 (N_18225,N_17638,N_17627);
or U18226 (N_18226,N_17705,N_17894);
or U18227 (N_18227,N_17864,N_17870);
nand U18228 (N_18228,N_17731,N_17515);
nor U18229 (N_18229,N_17740,N_17558);
or U18230 (N_18230,N_17838,N_17789);
and U18231 (N_18231,N_17681,N_17810);
nand U18232 (N_18232,N_17657,N_17746);
or U18233 (N_18233,N_17620,N_17589);
nand U18234 (N_18234,N_17803,N_17577);
or U18235 (N_18235,N_17714,N_17781);
nand U18236 (N_18236,N_17867,N_17933);
xor U18237 (N_18237,N_17915,N_17930);
nor U18238 (N_18238,N_17947,N_17783);
nand U18239 (N_18239,N_17548,N_17923);
nor U18240 (N_18240,N_17711,N_17656);
or U18241 (N_18241,N_17977,N_17728);
nor U18242 (N_18242,N_17654,N_17968);
and U18243 (N_18243,N_17983,N_17897);
nand U18244 (N_18244,N_17777,N_17780);
xnor U18245 (N_18245,N_17917,N_17901);
nand U18246 (N_18246,N_17841,N_17693);
and U18247 (N_18247,N_17582,N_17672);
nor U18248 (N_18248,N_17635,N_17749);
or U18249 (N_18249,N_17691,N_17739);
and U18250 (N_18250,N_17608,N_17912);
nand U18251 (N_18251,N_17627,N_17873);
and U18252 (N_18252,N_17778,N_17563);
nand U18253 (N_18253,N_17732,N_17664);
and U18254 (N_18254,N_17841,N_17617);
or U18255 (N_18255,N_17765,N_17715);
or U18256 (N_18256,N_17752,N_17558);
nor U18257 (N_18257,N_17969,N_17598);
nand U18258 (N_18258,N_17917,N_17985);
and U18259 (N_18259,N_17706,N_17872);
nor U18260 (N_18260,N_17627,N_17514);
nor U18261 (N_18261,N_17942,N_17660);
xor U18262 (N_18262,N_17832,N_17694);
xnor U18263 (N_18263,N_17844,N_17707);
or U18264 (N_18264,N_17649,N_17546);
or U18265 (N_18265,N_17740,N_17653);
xor U18266 (N_18266,N_17772,N_17898);
and U18267 (N_18267,N_17973,N_17776);
and U18268 (N_18268,N_17631,N_17594);
nand U18269 (N_18269,N_17837,N_17940);
nand U18270 (N_18270,N_17528,N_17774);
and U18271 (N_18271,N_17520,N_17760);
nand U18272 (N_18272,N_17725,N_17998);
xnor U18273 (N_18273,N_17741,N_17760);
xor U18274 (N_18274,N_17578,N_17817);
xnor U18275 (N_18275,N_17593,N_17690);
nand U18276 (N_18276,N_17965,N_17635);
nor U18277 (N_18277,N_17966,N_17566);
nand U18278 (N_18278,N_17732,N_17787);
nor U18279 (N_18279,N_17783,N_17918);
or U18280 (N_18280,N_17809,N_17505);
xnor U18281 (N_18281,N_17738,N_17903);
or U18282 (N_18282,N_17920,N_17935);
nand U18283 (N_18283,N_17750,N_17786);
nand U18284 (N_18284,N_17712,N_17888);
xnor U18285 (N_18285,N_17972,N_17981);
xnor U18286 (N_18286,N_17656,N_17865);
xnor U18287 (N_18287,N_17841,N_17511);
or U18288 (N_18288,N_17913,N_17848);
or U18289 (N_18289,N_17563,N_17990);
and U18290 (N_18290,N_17986,N_17836);
nand U18291 (N_18291,N_17722,N_17779);
nor U18292 (N_18292,N_17887,N_17575);
nor U18293 (N_18293,N_17660,N_17883);
nor U18294 (N_18294,N_17701,N_17928);
nor U18295 (N_18295,N_17660,N_17596);
nor U18296 (N_18296,N_17778,N_17804);
nor U18297 (N_18297,N_17941,N_17634);
or U18298 (N_18298,N_17970,N_17673);
nor U18299 (N_18299,N_17560,N_17861);
nor U18300 (N_18300,N_17928,N_17839);
xor U18301 (N_18301,N_17540,N_17990);
nand U18302 (N_18302,N_17688,N_17762);
and U18303 (N_18303,N_17972,N_17531);
nand U18304 (N_18304,N_17835,N_17859);
nor U18305 (N_18305,N_17784,N_17928);
nor U18306 (N_18306,N_17638,N_17755);
nor U18307 (N_18307,N_17692,N_17749);
and U18308 (N_18308,N_17799,N_17700);
and U18309 (N_18309,N_17932,N_17687);
nor U18310 (N_18310,N_17894,N_17611);
xnor U18311 (N_18311,N_17927,N_17580);
nor U18312 (N_18312,N_17875,N_17974);
nand U18313 (N_18313,N_17769,N_17990);
xnor U18314 (N_18314,N_17743,N_17724);
and U18315 (N_18315,N_17579,N_17670);
xnor U18316 (N_18316,N_17889,N_17618);
xnor U18317 (N_18317,N_17577,N_17593);
and U18318 (N_18318,N_17983,N_17841);
nor U18319 (N_18319,N_17841,N_17722);
xnor U18320 (N_18320,N_17920,N_17861);
and U18321 (N_18321,N_17564,N_17702);
or U18322 (N_18322,N_17756,N_17854);
nor U18323 (N_18323,N_17622,N_17896);
and U18324 (N_18324,N_17725,N_17578);
or U18325 (N_18325,N_17737,N_17723);
or U18326 (N_18326,N_17722,N_17687);
nor U18327 (N_18327,N_17988,N_17564);
nand U18328 (N_18328,N_17850,N_17592);
nor U18329 (N_18329,N_17929,N_17747);
xnor U18330 (N_18330,N_17570,N_17842);
or U18331 (N_18331,N_17791,N_17550);
and U18332 (N_18332,N_17902,N_17684);
nand U18333 (N_18333,N_17745,N_17778);
xnor U18334 (N_18334,N_17557,N_17793);
nand U18335 (N_18335,N_17781,N_17500);
and U18336 (N_18336,N_17591,N_17813);
nand U18337 (N_18337,N_17792,N_17684);
or U18338 (N_18338,N_17857,N_17611);
xnor U18339 (N_18339,N_17630,N_17733);
and U18340 (N_18340,N_17878,N_17982);
and U18341 (N_18341,N_17920,N_17528);
and U18342 (N_18342,N_17645,N_17751);
nand U18343 (N_18343,N_17804,N_17624);
nor U18344 (N_18344,N_17717,N_17580);
nand U18345 (N_18345,N_17837,N_17767);
xnor U18346 (N_18346,N_17535,N_17687);
xnor U18347 (N_18347,N_17815,N_17844);
and U18348 (N_18348,N_17747,N_17623);
nand U18349 (N_18349,N_17993,N_17743);
or U18350 (N_18350,N_17756,N_17787);
nor U18351 (N_18351,N_17989,N_17678);
nor U18352 (N_18352,N_17807,N_17990);
nor U18353 (N_18353,N_17691,N_17620);
or U18354 (N_18354,N_17944,N_17554);
nor U18355 (N_18355,N_17869,N_17630);
xor U18356 (N_18356,N_17616,N_17569);
nand U18357 (N_18357,N_17523,N_17871);
and U18358 (N_18358,N_17589,N_17954);
xor U18359 (N_18359,N_17515,N_17875);
and U18360 (N_18360,N_17897,N_17995);
or U18361 (N_18361,N_17742,N_17905);
nand U18362 (N_18362,N_17623,N_17922);
nor U18363 (N_18363,N_17861,N_17585);
nand U18364 (N_18364,N_17672,N_17804);
xnor U18365 (N_18365,N_17624,N_17832);
nor U18366 (N_18366,N_17766,N_17889);
and U18367 (N_18367,N_17903,N_17736);
or U18368 (N_18368,N_17823,N_17588);
nand U18369 (N_18369,N_17794,N_17807);
xor U18370 (N_18370,N_17854,N_17830);
nor U18371 (N_18371,N_17535,N_17591);
nor U18372 (N_18372,N_17604,N_17672);
or U18373 (N_18373,N_17768,N_17715);
nand U18374 (N_18374,N_17834,N_17907);
and U18375 (N_18375,N_17788,N_17744);
xor U18376 (N_18376,N_17772,N_17622);
and U18377 (N_18377,N_17839,N_17524);
or U18378 (N_18378,N_17897,N_17949);
and U18379 (N_18379,N_17845,N_17929);
or U18380 (N_18380,N_17908,N_17925);
nand U18381 (N_18381,N_17510,N_17629);
or U18382 (N_18382,N_17851,N_17797);
or U18383 (N_18383,N_17824,N_17666);
and U18384 (N_18384,N_17703,N_17817);
xnor U18385 (N_18385,N_17945,N_17685);
nor U18386 (N_18386,N_17537,N_17544);
or U18387 (N_18387,N_17633,N_17631);
or U18388 (N_18388,N_17993,N_17837);
nor U18389 (N_18389,N_17981,N_17935);
xor U18390 (N_18390,N_17660,N_17714);
and U18391 (N_18391,N_17845,N_17939);
xor U18392 (N_18392,N_17533,N_17978);
or U18393 (N_18393,N_17940,N_17519);
xnor U18394 (N_18394,N_17976,N_17672);
nor U18395 (N_18395,N_17912,N_17674);
nand U18396 (N_18396,N_17574,N_17969);
nand U18397 (N_18397,N_17997,N_17971);
and U18398 (N_18398,N_17542,N_17564);
or U18399 (N_18399,N_17685,N_17550);
xor U18400 (N_18400,N_17992,N_17753);
nand U18401 (N_18401,N_17535,N_17877);
nor U18402 (N_18402,N_17705,N_17946);
nor U18403 (N_18403,N_17979,N_17836);
nand U18404 (N_18404,N_17878,N_17555);
or U18405 (N_18405,N_17961,N_17733);
or U18406 (N_18406,N_17563,N_17892);
nor U18407 (N_18407,N_17738,N_17666);
xnor U18408 (N_18408,N_17512,N_17903);
and U18409 (N_18409,N_17693,N_17890);
and U18410 (N_18410,N_17733,N_17568);
or U18411 (N_18411,N_17590,N_17938);
xnor U18412 (N_18412,N_17743,N_17668);
or U18413 (N_18413,N_17746,N_17720);
xor U18414 (N_18414,N_17854,N_17728);
nor U18415 (N_18415,N_17872,N_17622);
or U18416 (N_18416,N_17710,N_17863);
or U18417 (N_18417,N_17550,N_17613);
and U18418 (N_18418,N_17822,N_17574);
nand U18419 (N_18419,N_17983,N_17517);
or U18420 (N_18420,N_17865,N_17866);
and U18421 (N_18421,N_17990,N_17979);
or U18422 (N_18422,N_17759,N_17596);
xnor U18423 (N_18423,N_17828,N_17790);
xnor U18424 (N_18424,N_17871,N_17685);
nor U18425 (N_18425,N_17823,N_17598);
nor U18426 (N_18426,N_17734,N_17797);
nor U18427 (N_18427,N_17504,N_17968);
and U18428 (N_18428,N_17879,N_17902);
nand U18429 (N_18429,N_17683,N_17872);
xnor U18430 (N_18430,N_17508,N_17784);
or U18431 (N_18431,N_17901,N_17910);
xnor U18432 (N_18432,N_17567,N_17855);
or U18433 (N_18433,N_17531,N_17719);
or U18434 (N_18434,N_17600,N_17998);
nand U18435 (N_18435,N_17617,N_17648);
xor U18436 (N_18436,N_17986,N_17705);
nor U18437 (N_18437,N_17588,N_17595);
or U18438 (N_18438,N_17808,N_17837);
and U18439 (N_18439,N_17611,N_17778);
xor U18440 (N_18440,N_17720,N_17705);
nor U18441 (N_18441,N_17536,N_17949);
or U18442 (N_18442,N_17986,N_17807);
xnor U18443 (N_18443,N_17939,N_17925);
xor U18444 (N_18444,N_17650,N_17817);
xnor U18445 (N_18445,N_17985,N_17992);
xor U18446 (N_18446,N_17584,N_17715);
or U18447 (N_18447,N_17527,N_17594);
nand U18448 (N_18448,N_17832,N_17988);
nor U18449 (N_18449,N_17676,N_17803);
nor U18450 (N_18450,N_17713,N_17703);
nor U18451 (N_18451,N_17999,N_17612);
and U18452 (N_18452,N_17704,N_17856);
xor U18453 (N_18453,N_17515,N_17956);
xor U18454 (N_18454,N_17791,N_17972);
or U18455 (N_18455,N_17983,N_17700);
nand U18456 (N_18456,N_17642,N_17705);
nand U18457 (N_18457,N_17952,N_17687);
nand U18458 (N_18458,N_17927,N_17842);
or U18459 (N_18459,N_17560,N_17653);
or U18460 (N_18460,N_17847,N_17846);
xnor U18461 (N_18461,N_17879,N_17982);
nor U18462 (N_18462,N_17998,N_17524);
nor U18463 (N_18463,N_17639,N_17834);
nor U18464 (N_18464,N_17809,N_17683);
nor U18465 (N_18465,N_17814,N_17881);
or U18466 (N_18466,N_17717,N_17964);
nor U18467 (N_18467,N_17591,N_17719);
nor U18468 (N_18468,N_17893,N_17912);
or U18469 (N_18469,N_17537,N_17815);
nand U18470 (N_18470,N_17706,N_17643);
nand U18471 (N_18471,N_17537,N_17586);
xnor U18472 (N_18472,N_17826,N_17680);
and U18473 (N_18473,N_17566,N_17536);
nand U18474 (N_18474,N_17781,N_17705);
xnor U18475 (N_18475,N_17500,N_17663);
nor U18476 (N_18476,N_17725,N_17641);
nand U18477 (N_18477,N_17733,N_17704);
xor U18478 (N_18478,N_17978,N_17579);
nand U18479 (N_18479,N_17714,N_17567);
nand U18480 (N_18480,N_17856,N_17592);
or U18481 (N_18481,N_17932,N_17887);
xor U18482 (N_18482,N_17995,N_17919);
nor U18483 (N_18483,N_17655,N_17532);
or U18484 (N_18484,N_17660,N_17688);
nor U18485 (N_18485,N_17599,N_17574);
or U18486 (N_18486,N_17652,N_17824);
or U18487 (N_18487,N_17861,N_17568);
xnor U18488 (N_18488,N_17867,N_17713);
and U18489 (N_18489,N_17944,N_17961);
and U18490 (N_18490,N_17691,N_17594);
nand U18491 (N_18491,N_17507,N_17616);
or U18492 (N_18492,N_17965,N_17990);
nand U18493 (N_18493,N_17953,N_17807);
nor U18494 (N_18494,N_17658,N_17606);
or U18495 (N_18495,N_17585,N_17965);
xnor U18496 (N_18496,N_17756,N_17934);
xnor U18497 (N_18497,N_17675,N_17537);
nor U18498 (N_18498,N_17772,N_17756);
or U18499 (N_18499,N_17917,N_17957);
or U18500 (N_18500,N_18284,N_18455);
nor U18501 (N_18501,N_18396,N_18457);
or U18502 (N_18502,N_18494,N_18395);
nand U18503 (N_18503,N_18064,N_18282);
or U18504 (N_18504,N_18382,N_18281);
and U18505 (N_18505,N_18491,N_18175);
and U18506 (N_18506,N_18480,N_18076);
nand U18507 (N_18507,N_18373,N_18213);
or U18508 (N_18508,N_18366,N_18136);
and U18509 (N_18509,N_18309,N_18279);
and U18510 (N_18510,N_18075,N_18238);
nand U18511 (N_18511,N_18258,N_18454);
nand U18512 (N_18512,N_18351,N_18036);
or U18513 (N_18513,N_18115,N_18318);
and U18514 (N_18514,N_18095,N_18011);
nor U18515 (N_18515,N_18026,N_18287);
xnor U18516 (N_18516,N_18296,N_18211);
xor U18517 (N_18517,N_18021,N_18404);
xnor U18518 (N_18518,N_18320,N_18051);
and U18519 (N_18519,N_18161,N_18473);
nor U18520 (N_18520,N_18363,N_18090);
or U18521 (N_18521,N_18035,N_18140);
and U18522 (N_18522,N_18183,N_18359);
nor U18523 (N_18523,N_18171,N_18354);
nand U18524 (N_18524,N_18121,N_18102);
and U18525 (N_18525,N_18106,N_18241);
or U18526 (N_18526,N_18043,N_18113);
nor U18527 (N_18527,N_18418,N_18391);
nand U18528 (N_18528,N_18149,N_18104);
or U18529 (N_18529,N_18132,N_18409);
or U18530 (N_18530,N_18264,N_18014);
nand U18531 (N_18531,N_18361,N_18466);
or U18532 (N_18532,N_18135,N_18180);
nor U18533 (N_18533,N_18001,N_18493);
nand U18534 (N_18534,N_18402,N_18044);
xor U18535 (N_18535,N_18177,N_18294);
nor U18536 (N_18536,N_18156,N_18393);
and U18537 (N_18537,N_18224,N_18255);
or U18538 (N_18538,N_18059,N_18267);
xor U18539 (N_18539,N_18441,N_18440);
nand U18540 (N_18540,N_18429,N_18338);
or U18541 (N_18541,N_18192,N_18375);
nand U18542 (N_18542,N_18147,N_18070);
and U18543 (N_18543,N_18196,N_18461);
xor U18544 (N_18544,N_18303,N_18145);
xnor U18545 (N_18545,N_18399,N_18487);
nor U18546 (N_18546,N_18029,N_18484);
or U18547 (N_18547,N_18261,N_18197);
or U18548 (N_18548,N_18253,N_18041);
nor U18549 (N_18549,N_18385,N_18206);
xor U18550 (N_18550,N_18214,N_18462);
nand U18551 (N_18551,N_18005,N_18308);
and U18552 (N_18552,N_18277,N_18038);
xor U18553 (N_18553,N_18424,N_18207);
nand U18554 (N_18554,N_18388,N_18439);
nand U18555 (N_18555,N_18293,N_18420);
and U18556 (N_18556,N_18364,N_18194);
nand U18557 (N_18557,N_18017,N_18269);
and U18558 (N_18558,N_18299,N_18371);
nor U18559 (N_18559,N_18481,N_18278);
nor U18560 (N_18560,N_18155,N_18406);
nor U18561 (N_18561,N_18428,N_18356);
nand U18562 (N_18562,N_18355,N_18478);
and U18563 (N_18563,N_18340,N_18127);
and U18564 (N_18564,N_18200,N_18431);
xnor U18565 (N_18565,N_18100,N_18226);
nor U18566 (N_18566,N_18419,N_18368);
xor U18567 (N_18567,N_18474,N_18326);
xnor U18568 (N_18568,N_18223,N_18436);
nand U18569 (N_18569,N_18144,N_18122);
or U18570 (N_18570,N_18025,N_18015);
nor U18571 (N_18571,N_18082,N_18448);
nor U18572 (N_18572,N_18221,N_18107);
xnor U18573 (N_18573,N_18413,N_18407);
nand U18574 (N_18574,N_18010,N_18479);
xnor U18575 (N_18575,N_18311,N_18425);
nor U18576 (N_18576,N_18463,N_18446);
nor U18577 (N_18577,N_18062,N_18381);
nand U18578 (N_18578,N_18182,N_18272);
or U18579 (N_18579,N_18482,N_18073);
nand U18580 (N_18580,N_18138,N_18445);
xor U18581 (N_18581,N_18344,N_18327);
nand U18582 (N_18582,N_18159,N_18004);
nor U18583 (N_18583,N_18112,N_18348);
nand U18584 (N_18584,N_18416,N_18316);
nor U18585 (N_18585,N_18237,N_18204);
nor U18586 (N_18586,N_18307,N_18378);
xor U18587 (N_18587,N_18114,N_18216);
or U18588 (N_18588,N_18153,N_18266);
and U18589 (N_18589,N_18151,N_18083);
and U18590 (N_18590,N_18165,N_18063);
and U18591 (N_18591,N_18489,N_18018);
nor U18592 (N_18592,N_18250,N_18016);
nor U18593 (N_18593,N_18442,N_18490);
xor U18594 (N_18594,N_18343,N_18154);
and U18595 (N_18595,N_18235,N_18139);
xnor U18596 (N_18596,N_18280,N_18372);
nor U18597 (N_18597,N_18242,N_18220);
nor U18598 (N_18598,N_18443,N_18067);
xnor U18599 (N_18599,N_18124,N_18110);
or U18600 (N_18600,N_18212,N_18485);
and U18601 (N_18601,N_18006,N_18398);
nand U18602 (N_18602,N_18084,N_18251);
nand U18603 (N_18603,N_18047,N_18077);
or U18604 (N_18604,N_18260,N_18290);
and U18605 (N_18605,N_18379,N_18142);
nand U18606 (N_18606,N_18225,N_18256);
nor U18607 (N_18607,N_18336,N_18450);
and U18608 (N_18608,N_18126,N_18332);
nand U18609 (N_18609,N_18012,N_18410);
or U18610 (N_18610,N_18358,N_18325);
nor U18611 (N_18611,N_18288,N_18158);
and U18612 (N_18612,N_18392,N_18013);
nand U18613 (N_18613,N_18360,N_18049);
nor U18614 (N_18614,N_18297,N_18060);
xnor U18615 (N_18615,N_18032,N_18345);
nand U18616 (N_18616,N_18313,N_18205);
and U18617 (N_18617,N_18133,N_18168);
nor U18618 (N_18618,N_18160,N_18000);
xor U18619 (N_18619,N_18117,N_18085);
nand U18620 (N_18620,N_18414,N_18471);
and U18621 (N_18621,N_18184,N_18056);
nand U18622 (N_18622,N_18169,N_18401);
and U18623 (N_18623,N_18486,N_18247);
and U18624 (N_18624,N_18289,N_18178);
nor U18625 (N_18625,N_18435,N_18459);
nand U18626 (N_18626,N_18315,N_18209);
xor U18627 (N_18627,N_18475,N_18065);
or U18628 (N_18628,N_18210,N_18141);
nand U18629 (N_18629,N_18191,N_18150);
nand U18630 (N_18630,N_18199,N_18098);
nor U18631 (N_18631,N_18397,N_18451);
nand U18632 (N_18632,N_18131,N_18053);
or U18633 (N_18633,N_18087,N_18497);
and U18634 (N_18634,N_18469,N_18152);
nor U18635 (N_18635,N_18331,N_18119);
or U18636 (N_18636,N_18239,N_18019);
or U18637 (N_18637,N_18219,N_18456);
nor U18638 (N_18638,N_18499,N_18426);
xor U18639 (N_18639,N_18302,N_18061);
xnor U18640 (N_18640,N_18190,N_18321);
nand U18641 (N_18641,N_18003,N_18086);
xor U18642 (N_18642,N_18476,N_18349);
nor U18643 (N_18643,N_18460,N_18262);
nand U18644 (N_18644,N_18066,N_18350);
xor U18645 (N_18645,N_18002,N_18329);
and U18646 (N_18646,N_18109,N_18097);
xnor U18647 (N_18647,N_18286,N_18042);
and U18648 (N_18648,N_18055,N_18233);
and U18649 (N_18649,N_18186,N_18317);
nand U18650 (N_18650,N_18408,N_18228);
nor U18651 (N_18651,N_18285,N_18034);
xnor U18652 (N_18652,N_18037,N_18477);
xnor U18653 (N_18653,N_18447,N_18230);
xor U18654 (N_18654,N_18273,N_18423);
xnor U18655 (N_18655,N_18172,N_18265);
nand U18656 (N_18656,N_18046,N_18328);
and U18657 (N_18657,N_18222,N_18008);
or U18658 (N_18658,N_18215,N_18157);
xor U18659 (N_18659,N_18217,N_18352);
xnor U18660 (N_18660,N_18092,N_18146);
xnor U18661 (N_18661,N_18434,N_18088);
nand U18662 (N_18662,N_18376,N_18495);
xnor U18663 (N_18663,N_18218,N_18128);
nor U18664 (N_18664,N_18301,N_18208);
and U18665 (N_18665,N_18292,N_18400);
and U18666 (N_18666,N_18458,N_18417);
or U18667 (N_18667,N_18319,N_18202);
xor U18668 (N_18668,N_18058,N_18257);
and U18669 (N_18669,N_18123,N_18283);
nand U18670 (N_18670,N_18118,N_18310);
nand U18671 (N_18671,N_18362,N_18027);
and U18672 (N_18672,N_18081,N_18470);
or U18673 (N_18673,N_18229,N_18148);
and U18674 (N_18674,N_18342,N_18452);
xor U18675 (N_18675,N_18488,N_18300);
xnor U18676 (N_18676,N_18185,N_18427);
and U18677 (N_18677,N_18129,N_18068);
nand U18678 (N_18678,N_18166,N_18120);
nand U18679 (N_18679,N_18020,N_18137);
and U18680 (N_18680,N_18181,N_18022);
or U18681 (N_18681,N_18268,N_18164);
and U18682 (N_18682,N_18449,N_18187);
or U18683 (N_18683,N_18023,N_18080);
and U18684 (N_18684,N_18162,N_18093);
xor U18685 (N_18685,N_18116,N_18498);
and U18686 (N_18686,N_18227,N_18305);
and U18687 (N_18687,N_18232,N_18105);
xor U18688 (N_18688,N_18339,N_18173);
and U18689 (N_18689,N_18089,N_18099);
nor U18690 (N_18690,N_18383,N_18333);
nor U18691 (N_18691,N_18030,N_18341);
or U18692 (N_18692,N_18031,N_18054);
or U18693 (N_18693,N_18403,N_18094);
nand U18694 (N_18694,N_18324,N_18271);
nor U18695 (N_18695,N_18415,N_18111);
xor U18696 (N_18696,N_18334,N_18143);
and U18697 (N_18697,N_18091,N_18048);
xor U18698 (N_18698,N_18130,N_18467);
nor U18699 (N_18699,N_18203,N_18078);
and U18700 (N_18700,N_18384,N_18353);
nand U18701 (N_18701,N_18050,N_18276);
nand U18702 (N_18702,N_18394,N_18453);
nor U18703 (N_18703,N_18179,N_18028);
nand U18704 (N_18704,N_18174,N_18421);
or U18705 (N_18705,N_18330,N_18430);
nor U18706 (N_18706,N_18347,N_18236);
xnor U18707 (N_18707,N_18198,N_18074);
nor U18708 (N_18708,N_18275,N_18437);
and U18709 (N_18709,N_18370,N_18433);
nor U18710 (N_18710,N_18306,N_18079);
nor U18711 (N_18711,N_18163,N_18411);
or U18712 (N_18712,N_18246,N_18422);
or U18713 (N_18713,N_18312,N_18007);
or U18714 (N_18714,N_18033,N_18374);
and U18715 (N_18715,N_18298,N_18270);
or U18716 (N_18716,N_18263,N_18464);
nand U18717 (N_18717,N_18380,N_18335);
and U18718 (N_18718,N_18314,N_18337);
or U18719 (N_18719,N_18252,N_18249);
xnor U18720 (N_18720,N_18259,N_18304);
or U18721 (N_18721,N_18483,N_18195);
nand U18722 (N_18722,N_18438,N_18492);
or U18723 (N_18723,N_18009,N_18322);
nand U18724 (N_18724,N_18248,N_18357);
nand U18725 (N_18725,N_18108,N_18295);
nor U18726 (N_18726,N_18365,N_18244);
or U18727 (N_18727,N_18103,N_18405);
nand U18728 (N_18728,N_18057,N_18369);
or U18729 (N_18729,N_18412,N_18496);
xor U18730 (N_18730,N_18254,N_18189);
or U18731 (N_18731,N_18193,N_18096);
xnor U18732 (N_18732,N_18052,N_18176);
and U18733 (N_18733,N_18274,N_18170);
xnor U18734 (N_18734,N_18346,N_18240);
nor U18735 (N_18735,N_18201,N_18071);
nand U18736 (N_18736,N_18125,N_18167);
nand U18737 (N_18737,N_18231,N_18188);
or U18738 (N_18738,N_18468,N_18072);
xnor U18739 (N_18739,N_18377,N_18387);
nand U18740 (N_18740,N_18024,N_18444);
xnor U18741 (N_18741,N_18390,N_18386);
xor U18742 (N_18742,N_18134,N_18045);
nand U18743 (N_18743,N_18291,N_18040);
nand U18744 (N_18744,N_18101,N_18069);
nand U18745 (N_18745,N_18039,N_18389);
xor U18746 (N_18746,N_18323,N_18465);
nand U18747 (N_18747,N_18432,N_18243);
or U18748 (N_18748,N_18367,N_18245);
and U18749 (N_18749,N_18472,N_18234);
nor U18750 (N_18750,N_18331,N_18047);
or U18751 (N_18751,N_18272,N_18469);
nor U18752 (N_18752,N_18047,N_18078);
nand U18753 (N_18753,N_18344,N_18020);
or U18754 (N_18754,N_18113,N_18339);
nand U18755 (N_18755,N_18072,N_18041);
nor U18756 (N_18756,N_18473,N_18450);
and U18757 (N_18757,N_18045,N_18307);
nand U18758 (N_18758,N_18436,N_18362);
or U18759 (N_18759,N_18166,N_18324);
nor U18760 (N_18760,N_18117,N_18198);
and U18761 (N_18761,N_18226,N_18327);
or U18762 (N_18762,N_18169,N_18303);
xnor U18763 (N_18763,N_18441,N_18265);
xnor U18764 (N_18764,N_18039,N_18494);
nor U18765 (N_18765,N_18146,N_18049);
or U18766 (N_18766,N_18035,N_18003);
nand U18767 (N_18767,N_18453,N_18116);
nor U18768 (N_18768,N_18172,N_18087);
nor U18769 (N_18769,N_18246,N_18184);
nor U18770 (N_18770,N_18164,N_18295);
nand U18771 (N_18771,N_18383,N_18355);
and U18772 (N_18772,N_18147,N_18469);
nand U18773 (N_18773,N_18298,N_18446);
xnor U18774 (N_18774,N_18416,N_18438);
nor U18775 (N_18775,N_18075,N_18490);
and U18776 (N_18776,N_18038,N_18279);
xor U18777 (N_18777,N_18129,N_18405);
nor U18778 (N_18778,N_18189,N_18391);
nand U18779 (N_18779,N_18078,N_18169);
and U18780 (N_18780,N_18293,N_18302);
nor U18781 (N_18781,N_18031,N_18406);
nor U18782 (N_18782,N_18197,N_18027);
nor U18783 (N_18783,N_18120,N_18088);
nand U18784 (N_18784,N_18208,N_18097);
xnor U18785 (N_18785,N_18259,N_18032);
or U18786 (N_18786,N_18215,N_18373);
or U18787 (N_18787,N_18496,N_18374);
and U18788 (N_18788,N_18209,N_18226);
nand U18789 (N_18789,N_18208,N_18165);
and U18790 (N_18790,N_18493,N_18265);
nand U18791 (N_18791,N_18194,N_18234);
nand U18792 (N_18792,N_18421,N_18406);
or U18793 (N_18793,N_18364,N_18164);
nor U18794 (N_18794,N_18491,N_18359);
and U18795 (N_18795,N_18332,N_18148);
xnor U18796 (N_18796,N_18099,N_18239);
and U18797 (N_18797,N_18218,N_18304);
nor U18798 (N_18798,N_18156,N_18137);
xor U18799 (N_18799,N_18402,N_18283);
and U18800 (N_18800,N_18242,N_18208);
or U18801 (N_18801,N_18310,N_18164);
xor U18802 (N_18802,N_18057,N_18496);
nand U18803 (N_18803,N_18452,N_18261);
nand U18804 (N_18804,N_18137,N_18087);
or U18805 (N_18805,N_18310,N_18197);
nand U18806 (N_18806,N_18444,N_18343);
and U18807 (N_18807,N_18341,N_18155);
and U18808 (N_18808,N_18049,N_18344);
and U18809 (N_18809,N_18005,N_18408);
nor U18810 (N_18810,N_18318,N_18214);
nand U18811 (N_18811,N_18055,N_18473);
and U18812 (N_18812,N_18047,N_18355);
xor U18813 (N_18813,N_18401,N_18054);
nor U18814 (N_18814,N_18346,N_18353);
and U18815 (N_18815,N_18354,N_18258);
and U18816 (N_18816,N_18284,N_18064);
or U18817 (N_18817,N_18060,N_18145);
or U18818 (N_18818,N_18473,N_18487);
nand U18819 (N_18819,N_18059,N_18287);
and U18820 (N_18820,N_18302,N_18073);
xnor U18821 (N_18821,N_18063,N_18425);
and U18822 (N_18822,N_18128,N_18493);
xnor U18823 (N_18823,N_18222,N_18447);
nand U18824 (N_18824,N_18424,N_18090);
and U18825 (N_18825,N_18192,N_18413);
nand U18826 (N_18826,N_18399,N_18076);
or U18827 (N_18827,N_18157,N_18427);
or U18828 (N_18828,N_18045,N_18259);
or U18829 (N_18829,N_18159,N_18206);
or U18830 (N_18830,N_18150,N_18080);
xor U18831 (N_18831,N_18112,N_18481);
xor U18832 (N_18832,N_18085,N_18438);
or U18833 (N_18833,N_18482,N_18240);
and U18834 (N_18834,N_18324,N_18242);
and U18835 (N_18835,N_18395,N_18246);
nand U18836 (N_18836,N_18200,N_18024);
nand U18837 (N_18837,N_18471,N_18115);
nand U18838 (N_18838,N_18038,N_18480);
and U18839 (N_18839,N_18331,N_18144);
or U18840 (N_18840,N_18274,N_18077);
nor U18841 (N_18841,N_18199,N_18479);
nand U18842 (N_18842,N_18008,N_18387);
xor U18843 (N_18843,N_18362,N_18120);
or U18844 (N_18844,N_18377,N_18266);
or U18845 (N_18845,N_18005,N_18042);
and U18846 (N_18846,N_18254,N_18158);
xor U18847 (N_18847,N_18073,N_18483);
nor U18848 (N_18848,N_18394,N_18373);
xor U18849 (N_18849,N_18305,N_18352);
xor U18850 (N_18850,N_18349,N_18140);
nand U18851 (N_18851,N_18421,N_18420);
xnor U18852 (N_18852,N_18331,N_18269);
xnor U18853 (N_18853,N_18070,N_18237);
xor U18854 (N_18854,N_18380,N_18341);
and U18855 (N_18855,N_18317,N_18497);
and U18856 (N_18856,N_18498,N_18397);
xor U18857 (N_18857,N_18303,N_18168);
nor U18858 (N_18858,N_18166,N_18383);
xnor U18859 (N_18859,N_18044,N_18273);
or U18860 (N_18860,N_18103,N_18158);
and U18861 (N_18861,N_18006,N_18428);
xnor U18862 (N_18862,N_18415,N_18050);
nor U18863 (N_18863,N_18138,N_18047);
and U18864 (N_18864,N_18180,N_18013);
xnor U18865 (N_18865,N_18322,N_18250);
nor U18866 (N_18866,N_18427,N_18496);
xor U18867 (N_18867,N_18485,N_18355);
nand U18868 (N_18868,N_18018,N_18280);
xor U18869 (N_18869,N_18452,N_18271);
nor U18870 (N_18870,N_18063,N_18420);
xnor U18871 (N_18871,N_18286,N_18188);
nand U18872 (N_18872,N_18009,N_18022);
and U18873 (N_18873,N_18484,N_18054);
nor U18874 (N_18874,N_18297,N_18427);
nor U18875 (N_18875,N_18236,N_18383);
nand U18876 (N_18876,N_18326,N_18251);
nand U18877 (N_18877,N_18133,N_18188);
nor U18878 (N_18878,N_18274,N_18292);
or U18879 (N_18879,N_18363,N_18378);
or U18880 (N_18880,N_18029,N_18240);
or U18881 (N_18881,N_18427,N_18198);
nand U18882 (N_18882,N_18323,N_18399);
nor U18883 (N_18883,N_18052,N_18249);
and U18884 (N_18884,N_18152,N_18413);
xnor U18885 (N_18885,N_18113,N_18147);
nor U18886 (N_18886,N_18013,N_18075);
and U18887 (N_18887,N_18074,N_18488);
nor U18888 (N_18888,N_18006,N_18141);
nor U18889 (N_18889,N_18231,N_18386);
and U18890 (N_18890,N_18052,N_18068);
or U18891 (N_18891,N_18298,N_18384);
or U18892 (N_18892,N_18299,N_18100);
and U18893 (N_18893,N_18258,N_18189);
nand U18894 (N_18894,N_18142,N_18329);
and U18895 (N_18895,N_18390,N_18186);
and U18896 (N_18896,N_18266,N_18386);
nand U18897 (N_18897,N_18168,N_18062);
nor U18898 (N_18898,N_18120,N_18128);
and U18899 (N_18899,N_18219,N_18429);
xnor U18900 (N_18900,N_18031,N_18189);
xor U18901 (N_18901,N_18384,N_18379);
and U18902 (N_18902,N_18117,N_18235);
or U18903 (N_18903,N_18003,N_18016);
xnor U18904 (N_18904,N_18328,N_18027);
xor U18905 (N_18905,N_18118,N_18303);
nor U18906 (N_18906,N_18451,N_18124);
nand U18907 (N_18907,N_18212,N_18058);
and U18908 (N_18908,N_18407,N_18189);
and U18909 (N_18909,N_18436,N_18094);
or U18910 (N_18910,N_18316,N_18160);
nand U18911 (N_18911,N_18424,N_18238);
nor U18912 (N_18912,N_18301,N_18257);
xnor U18913 (N_18913,N_18443,N_18485);
and U18914 (N_18914,N_18382,N_18033);
xnor U18915 (N_18915,N_18029,N_18230);
or U18916 (N_18916,N_18223,N_18414);
nand U18917 (N_18917,N_18350,N_18479);
and U18918 (N_18918,N_18242,N_18301);
nand U18919 (N_18919,N_18131,N_18181);
nor U18920 (N_18920,N_18452,N_18017);
and U18921 (N_18921,N_18141,N_18118);
and U18922 (N_18922,N_18178,N_18120);
xnor U18923 (N_18923,N_18287,N_18387);
nor U18924 (N_18924,N_18235,N_18043);
and U18925 (N_18925,N_18209,N_18050);
xor U18926 (N_18926,N_18050,N_18259);
xnor U18927 (N_18927,N_18246,N_18457);
xnor U18928 (N_18928,N_18082,N_18426);
nand U18929 (N_18929,N_18361,N_18322);
xor U18930 (N_18930,N_18051,N_18344);
nand U18931 (N_18931,N_18206,N_18425);
or U18932 (N_18932,N_18250,N_18227);
nor U18933 (N_18933,N_18281,N_18368);
nand U18934 (N_18934,N_18091,N_18322);
xor U18935 (N_18935,N_18445,N_18437);
nand U18936 (N_18936,N_18367,N_18112);
and U18937 (N_18937,N_18271,N_18096);
nand U18938 (N_18938,N_18343,N_18488);
nand U18939 (N_18939,N_18249,N_18138);
nor U18940 (N_18940,N_18286,N_18232);
or U18941 (N_18941,N_18267,N_18219);
nand U18942 (N_18942,N_18390,N_18339);
xor U18943 (N_18943,N_18325,N_18291);
nor U18944 (N_18944,N_18081,N_18475);
and U18945 (N_18945,N_18079,N_18014);
xnor U18946 (N_18946,N_18416,N_18406);
or U18947 (N_18947,N_18235,N_18250);
nand U18948 (N_18948,N_18478,N_18439);
nand U18949 (N_18949,N_18050,N_18142);
and U18950 (N_18950,N_18311,N_18072);
xor U18951 (N_18951,N_18050,N_18041);
xnor U18952 (N_18952,N_18377,N_18162);
or U18953 (N_18953,N_18297,N_18434);
or U18954 (N_18954,N_18027,N_18274);
nand U18955 (N_18955,N_18420,N_18004);
nor U18956 (N_18956,N_18431,N_18031);
and U18957 (N_18957,N_18469,N_18173);
and U18958 (N_18958,N_18317,N_18121);
nor U18959 (N_18959,N_18297,N_18189);
nand U18960 (N_18960,N_18292,N_18095);
or U18961 (N_18961,N_18394,N_18372);
or U18962 (N_18962,N_18215,N_18340);
nand U18963 (N_18963,N_18299,N_18108);
nor U18964 (N_18964,N_18466,N_18449);
xnor U18965 (N_18965,N_18432,N_18395);
or U18966 (N_18966,N_18134,N_18057);
nor U18967 (N_18967,N_18425,N_18336);
nor U18968 (N_18968,N_18004,N_18202);
xor U18969 (N_18969,N_18188,N_18343);
nor U18970 (N_18970,N_18336,N_18086);
and U18971 (N_18971,N_18046,N_18305);
nand U18972 (N_18972,N_18410,N_18378);
nand U18973 (N_18973,N_18251,N_18441);
and U18974 (N_18974,N_18476,N_18488);
nor U18975 (N_18975,N_18120,N_18052);
xnor U18976 (N_18976,N_18184,N_18283);
nand U18977 (N_18977,N_18085,N_18430);
and U18978 (N_18978,N_18192,N_18391);
and U18979 (N_18979,N_18149,N_18483);
nand U18980 (N_18980,N_18408,N_18038);
nand U18981 (N_18981,N_18448,N_18221);
nor U18982 (N_18982,N_18384,N_18184);
xnor U18983 (N_18983,N_18190,N_18470);
xnor U18984 (N_18984,N_18132,N_18008);
nand U18985 (N_18985,N_18325,N_18019);
and U18986 (N_18986,N_18393,N_18387);
nor U18987 (N_18987,N_18200,N_18414);
and U18988 (N_18988,N_18032,N_18076);
and U18989 (N_18989,N_18248,N_18493);
xor U18990 (N_18990,N_18191,N_18220);
and U18991 (N_18991,N_18286,N_18225);
or U18992 (N_18992,N_18022,N_18218);
or U18993 (N_18993,N_18349,N_18384);
or U18994 (N_18994,N_18409,N_18121);
and U18995 (N_18995,N_18077,N_18288);
or U18996 (N_18996,N_18429,N_18163);
or U18997 (N_18997,N_18170,N_18260);
or U18998 (N_18998,N_18116,N_18253);
and U18999 (N_18999,N_18379,N_18458);
nand U19000 (N_19000,N_18725,N_18568);
or U19001 (N_19001,N_18831,N_18686);
and U19002 (N_19002,N_18965,N_18892);
and U19003 (N_19003,N_18997,N_18878);
nor U19004 (N_19004,N_18757,N_18847);
nand U19005 (N_19005,N_18719,N_18896);
nand U19006 (N_19006,N_18631,N_18730);
xnor U19007 (N_19007,N_18870,N_18503);
nor U19008 (N_19008,N_18977,N_18671);
and U19009 (N_19009,N_18779,N_18880);
or U19010 (N_19010,N_18673,N_18639);
and U19011 (N_19011,N_18800,N_18993);
nand U19012 (N_19012,N_18821,N_18538);
nand U19013 (N_19013,N_18511,N_18844);
nor U19014 (N_19014,N_18634,N_18843);
and U19015 (N_19015,N_18565,N_18752);
or U19016 (N_19016,N_18708,N_18990);
nand U19017 (N_19017,N_18901,N_18760);
xor U19018 (N_19018,N_18682,N_18798);
and U19019 (N_19019,N_18845,N_18717);
nor U19020 (N_19020,N_18664,N_18992);
xor U19021 (N_19021,N_18987,N_18547);
nand U19022 (N_19022,N_18807,N_18777);
nor U19023 (N_19023,N_18562,N_18942);
nor U19024 (N_19024,N_18726,N_18913);
and U19025 (N_19025,N_18791,N_18999);
nand U19026 (N_19026,N_18533,N_18567);
and U19027 (N_19027,N_18770,N_18933);
nor U19028 (N_19028,N_18549,N_18552);
and U19029 (N_19029,N_18638,N_18665);
nand U19030 (N_19030,N_18700,N_18976);
or U19031 (N_19031,N_18830,N_18668);
or U19032 (N_19032,N_18893,N_18571);
and U19033 (N_19033,N_18619,N_18616);
nand U19034 (N_19034,N_18623,N_18528);
nand U19035 (N_19035,N_18863,N_18857);
nand U19036 (N_19036,N_18731,N_18524);
nand U19037 (N_19037,N_18795,N_18996);
and U19038 (N_19038,N_18529,N_18888);
or U19039 (N_19039,N_18615,N_18507);
nor U19040 (N_19040,N_18522,N_18756);
nor U19041 (N_19041,N_18501,N_18799);
xnor U19042 (N_19042,N_18793,N_18628);
and U19043 (N_19043,N_18903,N_18747);
or U19044 (N_19044,N_18781,N_18832);
xor U19045 (N_19045,N_18774,N_18763);
or U19046 (N_19046,N_18691,N_18755);
nor U19047 (N_19047,N_18923,N_18521);
and U19048 (N_19048,N_18908,N_18625);
nor U19049 (N_19049,N_18883,N_18932);
or U19050 (N_19050,N_18835,N_18972);
and U19051 (N_19051,N_18575,N_18978);
and U19052 (N_19052,N_18827,N_18504);
and U19053 (N_19053,N_18598,N_18592);
or U19054 (N_19054,N_18558,N_18710);
xor U19055 (N_19055,N_18729,N_18502);
nand U19056 (N_19056,N_18981,N_18829);
nor U19057 (N_19057,N_18527,N_18738);
nand U19058 (N_19058,N_18566,N_18998);
xor U19059 (N_19059,N_18956,N_18605);
nor U19060 (N_19060,N_18722,N_18563);
nor U19061 (N_19061,N_18946,N_18850);
nor U19062 (N_19062,N_18868,N_18825);
and U19063 (N_19063,N_18769,N_18890);
or U19064 (N_19064,N_18629,N_18810);
nand U19065 (N_19065,N_18657,N_18873);
and U19066 (N_19066,N_18654,N_18588);
or U19067 (N_19067,N_18790,N_18785);
nand U19068 (N_19068,N_18594,N_18787);
or U19069 (N_19069,N_18937,N_18662);
or U19070 (N_19070,N_18675,N_18739);
nand U19071 (N_19071,N_18822,N_18572);
or U19072 (N_19072,N_18688,N_18819);
xnor U19073 (N_19073,N_18559,N_18573);
xnor U19074 (N_19074,N_18804,N_18599);
nor U19075 (N_19075,N_18602,N_18927);
nand U19076 (N_19076,N_18906,N_18570);
xor U19077 (N_19077,N_18741,N_18669);
xor U19078 (N_19078,N_18643,N_18676);
and U19079 (N_19079,N_18612,N_18809);
and U19080 (N_19080,N_18737,N_18744);
xnor U19081 (N_19081,N_18805,N_18811);
nor U19082 (N_19082,N_18548,N_18525);
nor U19083 (N_19083,N_18564,N_18887);
or U19084 (N_19084,N_18649,N_18745);
and U19085 (N_19085,N_18814,N_18967);
nor U19086 (N_19086,N_18580,N_18620);
or U19087 (N_19087,N_18505,N_18553);
xor U19088 (N_19088,N_18792,N_18974);
and U19089 (N_19089,N_18980,N_18921);
or U19090 (N_19090,N_18532,N_18855);
and U19091 (N_19091,N_18622,N_18579);
nand U19092 (N_19092,N_18907,N_18551);
nand U19093 (N_19093,N_18578,N_18899);
nand U19094 (N_19094,N_18569,N_18900);
xnor U19095 (N_19095,N_18693,N_18627);
xnor U19096 (N_19096,N_18928,N_18584);
xnor U19097 (N_19097,N_18852,N_18544);
xnor U19098 (N_19098,N_18698,N_18851);
or U19099 (N_19099,N_18773,N_18585);
or U19100 (N_19100,N_18513,N_18876);
or U19101 (N_19101,N_18938,N_18866);
nor U19102 (N_19102,N_18824,N_18861);
and U19103 (N_19103,N_18670,N_18642);
nand U19104 (N_19104,N_18636,N_18886);
nand U19105 (N_19105,N_18754,N_18609);
nor U19106 (N_19106,N_18557,N_18969);
and U19107 (N_19107,N_18721,N_18540);
and U19108 (N_19108,N_18604,N_18608);
or U19109 (N_19109,N_18879,N_18813);
nand U19110 (N_19110,N_18838,N_18581);
and U19111 (N_19111,N_18839,N_18914);
xor U19112 (N_19112,N_18920,N_18771);
nand U19113 (N_19113,N_18661,N_18658);
nand U19114 (N_19114,N_18704,N_18746);
and U19115 (N_19115,N_18617,N_18836);
or U19116 (N_19116,N_18794,N_18520);
nor U19117 (N_19117,N_18561,N_18606);
nand U19118 (N_19118,N_18841,N_18954);
nand U19119 (N_19119,N_18542,N_18926);
or U19120 (N_19120,N_18645,N_18930);
xor U19121 (N_19121,N_18780,N_18950);
and U19122 (N_19122,N_18758,N_18591);
nand U19123 (N_19123,N_18797,N_18742);
xor U19124 (N_19124,N_18632,N_18699);
nor U19125 (N_19125,N_18711,N_18556);
nand U19126 (N_19126,N_18709,N_18788);
nand U19127 (N_19127,N_18621,N_18834);
xnor U19128 (N_19128,N_18646,N_18626);
nor U19129 (N_19129,N_18713,N_18947);
or U19130 (N_19130,N_18917,N_18840);
nand U19131 (N_19131,N_18782,N_18534);
nand U19132 (N_19132,N_18966,N_18775);
nor U19133 (N_19133,N_18940,N_18537);
nor U19134 (N_19134,N_18833,N_18812);
xor U19135 (N_19135,N_18768,N_18885);
nor U19136 (N_19136,N_18909,N_18948);
or U19137 (N_19137,N_18740,N_18536);
nand U19138 (N_19138,N_18955,N_18655);
nand U19139 (N_19139,N_18597,N_18510);
and U19140 (N_19140,N_18672,N_18970);
nor U19141 (N_19141,N_18881,N_18539);
nor U19142 (N_19142,N_18500,N_18724);
or U19143 (N_19143,N_18614,N_18595);
xor U19144 (N_19144,N_18714,N_18706);
xor U19145 (N_19145,N_18818,N_18678);
nor U19146 (N_19146,N_18973,N_18952);
nor U19147 (N_19147,N_18697,N_18867);
xor U19148 (N_19148,N_18647,N_18929);
nand U19149 (N_19149,N_18679,N_18960);
nor U19150 (N_19150,N_18541,N_18716);
nor U19151 (N_19151,N_18944,N_18856);
or U19152 (N_19152,N_18554,N_18786);
nand U19153 (N_19153,N_18660,N_18610);
nand U19154 (N_19154,N_18817,N_18743);
and U19155 (N_19155,N_18687,N_18733);
and U19156 (N_19156,N_18875,N_18535);
xor U19157 (N_19157,N_18509,N_18633);
nor U19158 (N_19158,N_18986,N_18667);
nand U19159 (N_19159,N_18858,N_18964);
nand U19160 (N_19160,N_18802,N_18968);
or U19161 (N_19161,N_18939,N_18694);
nor U19162 (N_19162,N_18689,N_18749);
nor U19163 (N_19163,N_18941,N_18518);
nand U19164 (N_19164,N_18652,N_18935);
xor U19165 (N_19165,N_18685,N_18640);
nor U19166 (N_19166,N_18842,N_18677);
nor U19167 (N_19167,N_18874,N_18583);
and U19168 (N_19168,N_18630,N_18806);
and U19169 (N_19169,N_18506,N_18849);
nor U19170 (N_19170,N_18653,N_18531);
nand U19171 (N_19171,N_18601,N_18959);
nand U19172 (N_19172,N_18735,N_18925);
xnor U19173 (N_19173,N_18732,N_18663);
xor U19174 (N_19174,N_18736,N_18936);
or U19175 (N_19175,N_18590,N_18512);
nand U19176 (N_19176,N_18848,N_18982);
xnor U19177 (N_19177,N_18611,N_18971);
nand U19178 (N_19178,N_18577,N_18593);
nand U19179 (N_19179,N_18764,N_18789);
nand U19180 (N_19180,N_18574,N_18681);
nor U19181 (N_19181,N_18707,N_18983);
nand U19182 (N_19182,N_18816,N_18712);
nor U19183 (N_19183,N_18703,N_18656);
nor U19184 (N_19184,N_18934,N_18778);
nor U19185 (N_19185,N_18924,N_18603);
xor U19186 (N_19186,N_18530,N_18526);
nand U19187 (N_19187,N_18674,N_18891);
xor U19188 (N_19188,N_18985,N_18820);
nor U19189 (N_19189,N_18905,N_18979);
or U19190 (N_19190,N_18916,N_18989);
nand U19191 (N_19191,N_18582,N_18823);
xor U19192 (N_19192,N_18963,N_18651);
nor U19193 (N_19193,N_18991,N_18796);
and U19194 (N_19194,N_18753,N_18696);
nand U19195 (N_19195,N_18803,N_18958);
xor U19196 (N_19196,N_18508,N_18666);
or U19197 (N_19197,N_18872,N_18589);
nand U19198 (N_19198,N_18895,N_18864);
nor U19199 (N_19199,N_18894,N_18680);
nand U19200 (N_19200,N_18750,N_18515);
or U19201 (N_19201,N_18600,N_18837);
xor U19202 (N_19202,N_18514,N_18846);
and U19203 (N_19203,N_18902,N_18587);
nand U19204 (N_19204,N_18692,N_18765);
and U19205 (N_19205,N_18523,N_18957);
nand U19206 (N_19206,N_18550,N_18545);
nor U19207 (N_19207,N_18826,N_18808);
and U19208 (N_19208,N_18869,N_18543);
xor U19209 (N_19209,N_18728,N_18659);
or U19210 (N_19210,N_18911,N_18854);
nor U19211 (N_19211,N_18723,N_18953);
xor U19212 (N_19212,N_18776,N_18884);
nor U19213 (N_19213,N_18690,N_18898);
or U19214 (N_19214,N_18727,N_18897);
xnor U19215 (N_19215,N_18975,N_18715);
nor U19216 (N_19216,N_18860,N_18871);
nand U19217 (N_19217,N_18949,N_18761);
xor U19218 (N_19218,N_18912,N_18718);
nor U19219 (N_19219,N_18815,N_18995);
and U19220 (N_19220,N_18931,N_18877);
and U19221 (N_19221,N_18734,N_18865);
nand U19222 (N_19222,N_18618,N_18984);
or U19223 (N_19223,N_18943,N_18882);
and U19224 (N_19224,N_18684,N_18919);
xor U19225 (N_19225,N_18546,N_18762);
xor U19226 (N_19226,N_18988,N_18945);
nor U19227 (N_19227,N_18720,N_18683);
nand U19228 (N_19228,N_18519,N_18889);
xnor U19229 (N_19229,N_18918,N_18859);
nor U19230 (N_19230,N_18759,N_18516);
and U19231 (N_19231,N_18904,N_18705);
nor U19232 (N_19232,N_18702,N_18650);
nand U19233 (N_19233,N_18517,N_18748);
and U19234 (N_19234,N_18862,N_18772);
or U19235 (N_19235,N_18560,N_18853);
or U19236 (N_19236,N_18751,N_18555);
or U19237 (N_19237,N_18994,N_18828);
xnor U19238 (N_19238,N_18951,N_18586);
or U19239 (N_19239,N_18607,N_18766);
nor U19240 (N_19240,N_18613,N_18637);
and U19241 (N_19241,N_18961,N_18801);
nand U19242 (N_19242,N_18648,N_18910);
or U19243 (N_19243,N_18641,N_18783);
xnor U19244 (N_19244,N_18635,N_18767);
xor U19245 (N_19245,N_18596,N_18695);
xnor U19246 (N_19246,N_18701,N_18784);
or U19247 (N_19247,N_18644,N_18922);
or U19248 (N_19248,N_18624,N_18915);
nand U19249 (N_19249,N_18962,N_18576);
nor U19250 (N_19250,N_18642,N_18516);
or U19251 (N_19251,N_18940,N_18617);
and U19252 (N_19252,N_18547,N_18582);
nor U19253 (N_19253,N_18958,N_18802);
xnor U19254 (N_19254,N_18762,N_18550);
and U19255 (N_19255,N_18677,N_18927);
nor U19256 (N_19256,N_18579,N_18819);
and U19257 (N_19257,N_18649,N_18848);
and U19258 (N_19258,N_18906,N_18834);
nand U19259 (N_19259,N_18866,N_18959);
xnor U19260 (N_19260,N_18946,N_18641);
and U19261 (N_19261,N_18598,N_18687);
and U19262 (N_19262,N_18684,N_18733);
or U19263 (N_19263,N_18612,N_18654);
or U19264 (N_19264,N_18916,N_18863);
nand U19265 (N_19265,N_18723,N_18973);
nand U19266 (N_19266,N_18821,N_18622);
nand U19267 (N_19267,N_18703,N_18878);
or U19268 (N_19268,N_18678,N_18993);
nor U19269 (N_19269,N_18551,N_18902);
nand U19270 (N_19270,N_18900,N_18707);
and U19271 (N_19271,N_18796,N_18677);
and U19272 (N_19272,N_18808,N_18750);
nor U19273 (N_19273,N_18930,N_18662);
and U19274 (N_19274,N_18561,N_18823);
nor U19275 (N_19275,N_18502,N_18631);
or U19276 (N_19276,N_18866,N_18963);
and U19277 (N_19277,N_18886,N_18525);
nor U19278 (N_19278,N_18939,N_18820);
nand U19279 (N_19279,N_18825,N_18583);
and U19280 (N_19280,N_18573,N_18649);
nand U19281 (N_19281,N_18736,N_18889);
and U19282 (N_19282,N_18968,N_18595);
nand U19283 (N_19283,N_18919,N_18541);
xnor U19284 (N_19284,N_18566,N_18786);
and U19285 (N_19285,N_18811,N_18504);
and U19286 (N_19286,N_18986,N_18681);
nor U19287 (N_19287,N_18946,N_18806);
xnor U19288 (N_19288,N_18748,N_18833);
xnor U19289 (N_19289,N_18950,N_18740);
xnor U19290 (N_19290,N_18813,N_18673);
xnor U19291 (N_19291,N_18836,N_18550);
xor U19292 (N_19292,N_18950,N_18753);
and U19293 (N_19293,N_18602,N_18632);
nand U19294 (N_19294,N_18850,N_18810);
nand U19295 (N_19295,N_18912,N_18772);
and U19296 (N_19296,N_18904,N_18628);
or U19297 (N_19297,N_18754,N_18914);
and U19298 (N_19298,N_18990,N_18636);
or U19299 (N_19299,N_18887,N_18934);
and U19300 (N_19300,N_18961,N_18815);
nand U19301 (N_19301,N_18527,N_18717);
nand U19302 (N_19302,N_18901,N_18950);
nor U19303 (N_19303,N_18712,N_18576);
nor U19304 (N_19304,N_18501,N_18510);
nand U19305 (N_19305,N_18681,N_18558);
or U19306 (N_19306,N_18511,N_18847);
or U19307 (N_19307,N_18928,N_18645);
or U19308 (N_19308,N_18722,N_18984);
nand U19309 (N_19309,N_18984,N_18798);
xor U19310 (N_19310,N_18685,N_18798);
xor U19311 (N_19311,N_18807,N_18507);
nand U19312 (N_19312,N_18579,N_18880);
xor U19313 (N_19313,N_18729,N_18897);
xor U19314 (N_19314,N_18785,N_18745);
nand U19315 (N_19315,N_18966,N_18529);
nor U19316 (N_19316,N_18581,N_18758);
and U19317 (N_19317,N_18629,N_18891);
nand U19318 (N_19318,N_18880,N_18680);
nand U19319 (N_19319,N_18784,N_18591);
xnor U19320 (N_19320,N_18568,N_18519);
or U19321 (N_19321,N_18908,N_18515);
xnor U19322 (N_19322,N_18678,N_18911);
and U19323 (N_19323,N_18533,N_18693);
or U19324 (N_19324,N_18830,N_18848);
nor U19325 (N_19325,N_18636,N_18780);
nor U19326 (N_19326,N_18562,N_18638);
nand U19327 (N_19327,N_18638,N_18644);
or U19328 (N_19328,N_18875,N_18753);
nor U19329 (N_19329,N_18617,N_18604);
and U19330 (N_19330,N_18685,N_18949);
or U19331 (N_19331,N_18724,N_18630);
or U19332 (N_19332,N_18757,N_18752);
nand U19333 (N_19333,N_18580,N_18604);
or U19334 (N_19334,N_18770,N_18600);
xor U19335 (N_19335,N_18878,N_18669);
or U19336 (N_19336,N_18897,N_18537);
nor U19337 (N_19337,N_18836,N_18866);
xnor U19338 (N_19338,N_18734,N_18670);
xor U19339 (N_19339,N_18538,N_18820);
nand U19340 (N_19340,N_18742,N_18583);
nor U19341 (N_19341,N_18580,N_18744);
xnor U19342 (N_19342,N_18869,N_18989);
or U19343 (N_19343,N_18773,N_18636);
xor U19344 (N_19344,N_18722,N_18549);
xor U19345 (N_19345,N_18847,N_18610);
nor U19346 (N_19346,N_18599,N_18944);
nand U19347 (N_19347,N_18646,N_18673);
nor U19348 (N_19348,N_18977,N_18867);
or U19349 (N_19349,N_18980,N_18743);
xor U19350 (N_19350,N_18713,N_18806);
nor U19351 (N_19351,N_18530,N_18689);
nor U19352 (N_19352,N_18862,N_18694);
or U19353 (N_19353,N_18870,N_18694);
nand U19354 (N_19354,N_18551,N_18632);
and U19355 (N_19355,N_18961,N_18838);
nand U19356 (N_19356,N_18902,N_18628);
xnor U19357 (N_19357,N_18961,N_18745);
nor U19358 (N_19358,N_18510,N_18974);
nand U19359 (N_19359,N_18541,N_18759);
or U19360 (N_19360,N_18617,N_18702);
nor U19361 (N_19361,N_18945,N_18729);
nand U19362 (N_19362,N_18527,N_18706);
and U19363 (N_19363,N_18824,N_18649);
nand U19364 (N_19364,N_18823,N_18962);
xnor U19365 (N_19365,N_18653,N_18674);
and U19366 (N_19366,N_18719,N_18932);
or U19367 (N_19367,N_18948,N_18726);
and U19368 (N_19368,N_18743,N_18841);
or U19369 (N_19369,N_18968,N_18989);
nor U19370 (N_19370,N_18943,N_18895);
or U19371 (N_19371,N_18533,N_18862);
or U19372 (N_19372,N_18893,N_18705);
or U19373 (N_19373,N_18991,N_18735);
or U19374 (N_19374,N_18933,N_18624);
nand U19375 (N_19375,N_18812,N_18605);
nand U19376 (N_19376,N_18589,N_18863);
nor U19377 (N_19377,N_18843,N_18509);
nand U19378 (N_19378,N_18930,N_18570);
xnor U19379 (N_19379,N_18825,N_18684);
and U19380 (N_19380,N_18514,N_18730);
nor U19381 (N_19381,N_18776,N_18942);
nand U19382 (N_19382,N_18715,N_18909);
nand U19383 (N_19383,N_18864,N_18555);
and U19384 (N_19384,N_18679,N_18957);
nand U19385 (N_19385,N_18716,N_18777);
nor U19386 (N_19386,N_18500,N_18718);
or U19387 (N_19387,N_18637,N_18726);
and U19388 (N_19388,N_18704,N_18694);
nand U19389 (N_19389,N_18693,N_18768);
xor U19390 (N_19390,N_18960,N_18927);
nand U19391 (N_19391,N_18610,N_18830);
or U19392 (N_19392,N_18655,N_18857);
nand U19393 (N_19393,N_18870,N_18922);
and U19394 (N_19394,N_18514,N_18879);
or U19395 (N_19395,N_18741,N_18958);
xor U19396 (N_19396,N_18991,N_18510);
xor U19397 (N_19397,N_18856,N_18958);
and U19398 (N_19398,N_18690,N_18572);
nand U19399 (N_19399,N_18512,N_18903);
and U19400 (N_19400,N_18558,N_18778);
and U19401 (N_19401,N_18931,N_18691);
or U19402 (N_19402,N_18810,N_18556);
nor U19403 (N_19403,N_18823,N_18616);
nand U19404 (N_19404,N_18905,N_18723);
nor U19405 (N_19405,N_18697,N_18792);
nand U19406 (N_19406,N_18701,N_18942);
xor U19407 (N_19407,N_18558,N_18981);
and U19408 (N_19408,N_18694,N_18986);
nor U19409 (N_19409,N_18512,N_18892);
and U19410 (N_19410,N_18888,N_18699);
xor U19411 (N_19411,N_18916,N_18900);
xor U19412 (N_19412,N_18761,N_18998);
nor U19413 (N_19413,N_18620,N_18715);
nand U19414 (N_19414,N_18952,N_18926);
and U19415 (N_19415,N_18763,N_18750);
nand U19416 (N_19416,N_18574,N_18921);
xnor U19417 (N_19417,N_18665,N_18733);
and U19418 (N_19418,N_18775,N_18507);
xnor U19419 (N_19419,N_18940,N_18803);
xnor U19420 (N_19420,N_18620,N_18829);
and U19421 (N_19421,N_18853,N_18688);
xnor U19422 (N_19422,N_18621,N_18564);
xnor U19423 (N_19423,N_18729,N_18529);
xor U19424 (N_19424,N_18943,N_18824);
xnor U19425 (N_19425,N_18529,N_18797);
and U19426 (N_19426,N_18937,N_18800);
and U19427 (N_19427,N_18939,N_18623);
and U19428 (N_19428,N_18509,N_18569);
nor U19429 (N_19429,N_18823,N_18554);
nand U19430 (N_19430,N_18761,N_18763);
nand U19431 (N_19431,N_18708,N_18770);
nor U19432 (N_19432,N_18642,N_18748);
and U19433 (N_19433,N_18990,N_18663);
and U19434 (N_19434,N_18680,N_18993);
nor U19435 (N_19435,N_18875,N_18928);
and U19436 (N_19436,N_18555,N_18716);
and U19437 (N_19437,N_18816,N_18606);
nor U19438 (N_19438,N_18684,N_18731);
xor U19439 (N_19439,N_18520,N_18610);
nor U19440 (N_19440,N_18669,N_18782);
and U19441 (N_19441,N_18924,N_18743);
and U19442 (N_19442,N_18764,N_18579);
and U19443 (N_19443,N_18912,N_18832);
nand U19444 (N_19444,N_18809,N_18964);
nor U19445 (N_19445,N_18779,N_18793);
nand U19446 (N_19446,N_18517,N_18793);
and U19447 (N_19447,N_18500,N_18630);
xnor U19448 (N_19448,N_18751,N_18617);
or U19449 (N_19449,N_18648,N_18840);
and U19450 (N_19450,N_18633,N_18942);
and U19451 (N_19451,N_18657,N_18817);
and U19452 (N_19452,N_18848,N_18760);
and U19453 (N_19453,N_18749,N_18649);
or U19454 (N_19454,N_18605,N_18614);
nand U19455 (N_19455,N_18726,N_18785);
xnor U19456 (N_19456,N_18547,N_18513);
nand U19457 (N_19457,N_18626,N_18515);
and U19458 (N_19458,N_18978,N_18833);
nor U19459 (N_19459,N_18781,N_18788);
nor U19460 (N_19460,N_18886,N_18683);
xor U19461 (N_19461,N_18918,N_18793);
and U19462 (N_19462,N_18628,N_18869);
and U19463 (N_19463,N_18682,N_18884);
xnor U19464 (N_19464,N_18918,N_18879);
nand U19465 (N_19465,N_18921,N_18501);
nand U19466 (N_19466,N_18930,N_18981);
nand U19467 (N_19467,N_18644,N_18800);
or U19468 (N_19468,N_18912,N_18530);
xor U19469 (N_19469,N_18956,N_18975);
xnor U19470 (N_19470,N_18988,N_18861);
and U19471 (N_19471,N_18808,N_18963);
nand U19472 (N_19472,N_18547,N_18781);
nor U19473 (N_19473,N_18802,N_18831);
xnor U19474 (N_19474,N_18858,N_18607);
nor U19475 (N_19475,N_18619,N_18888);
xor U19476 (N_19476,N_18838,N_18557);
nand U19477 (N_19477,N_18620,N_18565);
nor U19478 (N_19478,N_18744,N_18658);
nor U19479 (N_19479,N_18594,N_18873);
nor U19480 (N_19480,N_18685,N_18636);
and U19481 (N_19481,N_18967,N_18556);
or U19482 (N_19482,N_18543,N_18877);
xnor U19483 (N_19483,N_18712,N_18534);
nor U19484 (N_19484,N_18918,N_18515);
or U19485 (N_19485,N_18916,N_18545);
and U19486 (N_19486,N_18696,N_18514);
and U19487 (N_19487,N_18701,N_18774);
nand U19488 (N_19488,N_18693,N_18513);
nor U19489 (N_19489,N_18745,N_18860);
and U19490 (N_19490,N_18729,N_18619);
or U19491 (N_19491,N_18833,N_18822);
nor U19492 (N_19492,N_18932,N_18529);
nor U19493 (N_19493,N_18562,N_18570);
nand U19494 (N_19494,N_18793,N_18584);
nand U19495 (N_19495,N_18831,N_18570);
nor U19496 (N_19496,N_18909,N_18896);
and U19497 (N_19497,N_18710,N_18954);
and U19498 (N_19498,N_18607,N_18810);
nor U19499 (N_19499,N_18741,N_18680);
or U19500 (N_19500,N_19160,N_19141);
nor U19501 (N_19501,N_19067,N_19345);
and U19502 (N_19502,N_19153,N_19177);
nand U19503 (N_19503,N_19365,N_19033);
nand U19504 (N_19504,N_19037,N_19253);
nor U19505 (N_19505,N_19127,N_19169);
xnor U19506 (N_19506,N_19464,N_19405);
or U19507 (N_19507,N_19489,N_19439);
nand U19508 (N_19508,N_19041,N_19254);
and U19509 (N_19509,N_19247,N_19011);
nand U19510 (N_19510,N_19029,N_19392);
nor U19511 (N_19511,N_19337,N_19239);
and U19512 (N_19512,N_19133,N_19055);
or U19513 (N_19513,N_19204,N_19143);
nor U19514 (N_19514,N_19475,N_19425);
nand U19515 (N_19515,N_19105,N_19452);
nand U19516 (N_19516,N_19137,N_19236);
nand U19517 (N_19517,N_19146,N_19013);
and U19518 (N_19518,N_19447,N_19002);
and U19519 (N_19519,N_19463,N_19344);
or U19520 (N_19520,N_19458,N_19301);
or U19521 (N_19521,N_19049,N_19418);
nand U19522 (N_19522,N_19008,N_19496);
nand U19523 (N_19523,N_19080,N_19082);
nor U19524 (N_19524,N_19052,N_19191);
and U19525 (N_19525,N_19035,N_19100);
nand U19526 (N_19526,N_19310,N_19183);
or U19527 (N_19527,N_19111,N_19370);
xor U19528 (N_19528,N_19385,N_19390);
and U19529 (N_19529,N_19134,N_19139);
and U19530 (N_19530,N_19097,N_19075);
nand U19531 (N_19531,N_19154,N_19042);
or U19532 (N_19532,N_19380,N_19271);
and U19533 (N_19533,N_19226,N_19393);
xor U19534 (N_19534,N_19443,N_19218);
nand U19535 (N_19535,N_19409,N_19259);
nor U19536 (N_19536,N_19479,N_19126);
xor U19537 (N_19537,N_19015,N_19469);
xnor U19538 (N_19538,N_19286,N_19106);
or U19539 (N_19539,N_19039,N_19113);
or U19540 (N_19540,N_19244,N_19468);
and U19541 (N_19541,N_19058,N_19459);
and U19542 (N_19542,N_19145,N_19031);
nor U19543 (N_19543,N_19270,N_19394);
and U19544 (N_19544,N_19158,N_19077);
nand U19545 (N_19545,N_19197,N_19320);
nor U19546 (N_19546,N_19240,N_19351);
and U19547 (N_19547,N_19352,N_19114);
xor U19548 (N_19548,N_19428,N_19006);
nand U19549 (N_19549,N_19168,N_19482);
and U19550 (N_19550,N_19026,N_19333);
nand U19551 (N_19551,N_19446,N_19328);
xnor U19552 (N_19552,N_19068,N_19233);
nand U19553 (N_19553,N_19257,N_19147);
or U19554 (N_19554,N_19156,N_19148);
nand U19555 (N_19555,N_19359,N_19074);
nor U19556 (N_19556,N_19076,N_19431);
and U19557 (N_19557,N_19000,N_19451);
xor U19558 (N_19558,N_19429,N_19317);
nor U19559 (N_19559,N_19493,N_19305);
nand U19560 (N_19560,N_19064,N_19379);
or U19561 (N_19561,N_19422,N_19216);
xnor U19562 (N_19562,N_19420,N_19151);
nand U19563 (N_19563,N_19339,N_19432);
and U19564 (N_19564,N_19349,N_19223);
nand U19565 (N_19565,N_19371,N_19047);
or U19566 (N_19566,N_19028,N_19121);
nand U19567 (N_19567,N_19262,N_19250);
and U19568 (N_19568,N_19099,N_19228);
xor U19569 (N_19569,N_19001,N_19030);
nor U19570 (N_19570,N_19258,N_19263);
nor U19571 (N_19571,N_19481,N_19036);
nand U19572 (N_19572,N_19378,N_19059);
nand U19573 (N_19573,N_19265,N_19167);
nand U19574 (N_19574,N_19086,N_19484);
nor U19575 (N_19575,N_19264,N_19119);
and U19576 (N_19576,N_19492,N_19499);
or U19577 (N_19577,N_19088,N_19315);
or U19578 (N_19578,N_19051,N_19162);
nand U19579 (N_19579,N_19377,N_19275);
nor U19580 (N_19580,N_19303,N_19172);
nand U19581 (N_19581,N_19255,N_19292);
xor U19582 (N_19582,N_19066,N_19101);
xor U19583 (N_19583,N_19136,N_19347);
xor U19584 (N_19584,N_19291,N_19159);
or U19585 (N_19585,N_19391,N_19338);
and U19586 (N_19586,N_19020,N_19217);
nand U19587 (N_19587,N_19161,N_19355);
nand U19588 (N_19588,N_19222,N_19408);
xor U19589 (N_19589,N_19190,N_19060);
nand U19590 (N_19590,N_19282,N_19232);
nand U19591 (N_19591,N_19297,N_19112);
nand U19592 (N_19592,N_19381,N_19415);
nor U19593 (N_19593,N_19230,N_19063);
nor U19594 (N_19594,N_19289,N_19318);
nor U19595 (N_19595,N_19323,N_19166);
or U19596 (N_19596,N_19384,N_19465);
or U19597 (N_19597,N_19280,N_19186);
xnor U19598 (N_19598,N_19382,N_19205);
and U19599 (N_19599,N_19092,N_19497);
nor U19600 (N_19600,N_19219,N_19235);
nor U19601 (N_19601,N_19144,N_19331);
nor U19602 (N_19602,N_19046,N_19322);
xnor U19603 (N_19603,N_19477,N_19329);
nand U19604 (N_19604,N_19098,N_19246);
nor U19605 (N_19605,N_19478,N_19043);
nor U19606 (N_19606,N_19430,N_19470);
nor U19607 (N_19607,N_19399,N_19056);
or U19608 (N_19608,N_19438,N_19192);
or U19609 (N_19609,N_19313,N_19107);
nand U19610 (N_19610,N_19367,N_19116);
and U19611 (N_19611,N_19495,N_19407);
nor U19612 (N_19612,N_19241,N_19442);
nand U19613 (N_19613,N_19061,N_19403);
and U19614 (N_19614,N_19248,N_19188);
nand U19615 (N_19615,N_19091,N_19335);
nand U19616 (N_19616,N_19357,N_19319);
xor U19617 (N_19617,N_19312,N_19473);
and U19618 (N_19618,N_19308,N_19184);
or U19619 (N_19619,N_19461,N_19096);
nand U19620 (N_19620,N_19109,N_19069);
nor U19621 (N_19621,N_19135,N_19251);
xor U19622 (N_19622,N_19368,N_19453);
and U19623 (N_19623,N_19003,N_19087);
and U19624 (N_19624,N_19395,N_19332);
or U19625 (N_19625,N_19314,N_19130);
and U19626 (N_19626,N_19129,N_19140);
nand U19627 (N_19627,N_19449,N_19157);
nand U19628 (N_19628,N_19366,N_19256);
or U19629 (N_19629,N_19454,N_19103);
xnor U19630 (N_19630,N_19456,N_19071);
nand U19631 (N_19631,N_19180,N_19007);
nor U19632 (N_19632,N_19362,N_19155);
or U19633 (N_19633,N_19138,N_19325);
nand U19634 (N_19634,N_19016,N_19072);
nor U19635 (N_19635,N_19245,N_19388);
nor U19636 (N_19636,N_19181,N_19152);
nand U19637 (N_19637,N_19298,N_19027);
xnor U19638 (N_19638,N_19182,N_19488);
or U19639 (N_19639,N_19083,N_19490);
xor U19640 (N_19640,N_19120,N_19336);
xnor U19641 (N_19641,N_19372,N_19227);
or U19642 (N_19642,N_19110,N_19242);
or U19643 (N_19643,N_19118,N_19348);
or U19644 (N_19644,N_19079,N_19173);
or U19645 (N_19645,N_19455,N_19040);
nand U19646 (N_19646,N_19022,N_19081);
xnor U19647 (N_19647,N_19423,N_19293);
nand U19648 (N_19648,N_19164,N_19476);
or U19649 (N_19649,N_19045,N_19462);
nand U19650 (N_19650,N_19194,N_19207);
nand U19651 (N_19651,N_19402,N_19448);
or U19652 (N_19652,N_19278,N_19386);
xnor U19653 (N_19653,N_19108,N_19005);
and U19654 (N_19654,N_19050,N_19221);
or U19655 (N_19655,N_19165,N_19234);
xnor U19656 (N_19656,N_19273,N_19125);
nor U19657 (N_19657,N_19413,N_19122);
nand U19658 (N_19658,N_19324,N_19179);
xor U19659 (N_19659,N_19341,N_19436);
nand U19660 (N_19660,N_19023,N_19261);
and U19661 (N_19661,N_19417,N_19426);
nor U19662 (N_19662,N_19363,N_19062);
nor U19663 (N_19663,N_19201,N_19414);
xor U19664 (N_19664,N_19406,N_19124);
nand U19665 (N_19665,N_19123,N_19311);
or U19666 (N_19666,N_19326,N_19018);
xor U19667 (N_19667,N_19200,N_19485);
or U19668 (N_19668,N_19342,N_19229);
nand U19669 (N_19669,N_19334,N_19435);
or U19670 (N_19670,N_19149,N_19327);
nand U19671 (N_19671,N_19210,N_19471);
or U19672 (N_19672,N_19203,N_19296);
xnor U19673 (N_19673,N_19460,N_19330);
nor U19674 (N_19674,N_19316,N_19078);
nand U19675 (N_19675,N_19411,N_19225);
nand U19676 (N_19676,N_19131,N_19009);
or U19677 (N_19677,N_19486,N_19350);
nor U19678 (N_19678,N_19434,N_19400);
nand U19679 (N_19679,N_19376,N_19032);
nand U19680 (N_19680,N_19014,N_19252);
nor U19681 (N_19681,N_19224,N_19437);
nor U19682 (N_19682,N_19290,N_19171);
nand U19683 (N_19683,N_19176,N_19054);
nor U19684 (N_19684,N_19266,N_19208);
xor U19685 (N_19685,N_19354,N_19187);
xor U19686 (N_19686,N_19170,N_19364);
xnor U19687 (N_19687,N_19279,N_19057);
nor U19688 (N_19688,N_19189,N_19277);
or U19689 (N_19689,N_19211,N_19206);
nor U19690 (N_19690,N_19024,N_19281);
nand U19691 (N_19691,N_19412,N_19053);
and U19692 (N_19692,N_19093,N_19285);
nor U19693 (N_19693,N_19466,N_19094);
and U19694 (N_19694,N_19295,N_19360);
xor U19695 (N_19695,N_19260,N_19498);
or U19696 (N_19696,N_19450,N_19025);
nand U19697 (N_19697,N_19491,N_19034);
nor U19698 (N_19698,N_19410,N_19202);
or U19699 (N_19699,N_19012,N_19472);
nor U19700 (N_19700,N_19195,N_19142);
nor U19701 (N_19701,N_19215,N_19175);
or U19702 (N_19702,N_19115,N_19284);
nand U19703 (N_19703,N_19268,N_19369);
and U19704 (N_19704,N_19433,N_19150);
nand U19705 (N_19705,N_19174,N_19231);
xnor U19706 (N_19706,N_19356,N_19283);
xor U19707 (N_19707,N_19358,N_19300);
nor U19708 (N_19708,N_19019,N_19209);
nor U19709 (N_19709,N_19073,N_19214);
xor U19710 (N_19710,N_19220,N_19445);
and U19711 (N_19711,N_19361,N_19272);
or U19712 (N_19712,N_19383,N_19404);
xnor U19713 (N_19713,N_19084,N_19274);
nor U19714 (N_19714,N_19419,N_19102);
nand U19715 (N_19715,N_19196,N_19421);
nor U19716 (N_19716,N_19474,N_19185);
or U19717 (N_19717,N_19427,N_19237);
xor U19718 (N_19718,N_19267,N_19243);
nor U19719 (N_19719,N_19401,N_19276);
xor U19720 (N_19720,N_19387,N_19494);
nor U19721 (N_19721,N_19269,N_19128);
xnor U19722 (N_19722,N_19457,N_19398);
nand U19723 (N_19723,N_19480,N_19212);
and U19724 (N_19724,N_19375,N_19302);
xnor U19725 (N_19725,N_19441,N_19090);
or U19726 (N_19726,N_19089,N_19010);
nor U19727 (N_19727,N_19321,N_19085);
nand U19728 (N_19728,N_19104,N_19070);
or U19729 (N_19729,N_19017,N_19340);
or U19730 (N_19730,N_19444,N_19178);
or U19731 (N_19731,N_19021,N_19343);
nor U19732 (N_19732,N_19346,N_19396);
and U19733 (N_19733,N_19353,N_19287);
nand U19734 (N_19734,N_19048,N_19373);
nand U19735 (N_19735,N_19044,N_19416);
and U19736 (N_19736,N_19424,N_19065);
or U19737 (N_19737,N_19307,N_19304);
and U19738 (N_19738,N_19299,N_19306);
nand U19739 (N_19739,N_19483,N_19038);
xor U19740 (N_19740,N_19117,N_19238);
and U19741 (N_19741,N_19389,N_19440);
and U19742 (N_19742,N_19213,N_19309);
or U19743 (N_19743,N_19198,N_19132);
nand U19744 (N_19744,N_19294,N_19397);
or U19745 (N_19745,N_19095,N_19374);
nand U19746 (N_19746,N_19467,N_19193);
nor U19747 (N_19747,N_19487,N_19004);
and U19748 (N_19748,N_19199,N_19163);
or U19749 (N_19749,N_19288,N_19249);
nand U19750 (N_19750,N_19188,N_19023);
nor U19751 (N_19751,N_19181,N_19149);
or U19752 (N_19752,N_19256,N_19374);
xor U19753 (N_19753,N_19036,N_19021);
nor U19754 (N_19754,N_19347,N_19359);
xor U19755 (N_19755,N_19072,N_19183);
nor U19756 (N_19756,N_19402,N_19366);
or U19757 (N_19757,N_19108,N_19467);
xor U19758 (N_19758,N_19380,N_19128);
or U19759 (N_19759,N_19357,N_19329);
or U19760 (N_19760,N_19096,N_19042);
and U19761 (N_19761,N_19392,N_19451);
xnor U19762 (N_19762,N_19153,N_19067);
nand U19763 (N_19763,N_19347,N_19371);
nor U19764 (N_19764,N_19411,N_19067);
xor U19765 (N_19765,N_19160,N_19304);
and U19766 (N_19766,N_19392,N_19477);
nor U19767 (N_19767,N_19416,N_19329);
nor U19768 (N_19768,N_19065,N_19203);
and U19769 (N_19769,N_19478,N_19335);
nor U19770 (N_19770,N_19293,N_19369);
nor U19771 (N_19771,N_19388,N_19483);
and U19772 (N_19772,N_19464,N_19248);
nand U19773 (N_19773,N_19449,N_19366);
or U19774 (N_19774,N_19453,N_19265);
nand U19775 (N_19775,N_19067,N_19454);
or U19776 (N_19776,N_19248,N_19376);
or U19777 (N_19777,N_19130,N_19423);
nand U19778 (N_19778,N_19269,N_19310);
and U19779 (N_19779,N_19128,N_19222);
or U19780 (N_19780,N_19203,N_19305);
or U19781 (N_19781,N_19025,N_19428);
or U19782 (N_19782,N_19372,N_19275);
xnor U19783 (N_19783,N_19109,N_19250);
xnor U19784 (N_19784,N_19285,N_19234);
nand U19785 (N_19785,N_19475,N_19413);
nand U19786 (N_19786,N_19250,N_19101);
nor U19787 (N_19787,N_19044,N_19117);
or U19788 (N_19788,N_19090,N_19344);
xnor U19789 (N_19789,N_19286,N_19137);
nand U19790 (N_19790,N_19227,N_19354);
or U19791 (N_19791,N_19309,N_19153);
nand U19792 (N_19792,N_19298,N_19271);
and U19793 (N_19793,N_19378,N_19225);
nand U19794 (N_19794,N_19284,N_19312);
xor U19795 (N_19795,N_19490,N_19223);
xnor U19796 (N_19796,N_19342,N_19259);
and U19797 (N_19797,N_19325,N_19450);
and U19798 (N_19798,N_19265,N_19009);
and U19799 (N_19799,N_19146,N_19001);
nand U19800 (N_19800,N_19476,N_19323);
nand U19801 (N_19801,N_19096,N_19013);
or U19802 (N_19802,N_19203,N_19324);
and U19803 (N_19803,N_19300,N_19027);
nor U19804 (N_19804,N_19297,N_19373);
xnor U19805 (N_19805,N_19360,N_19078);
and U19806 (N_19806,N_19330,N_19025);
nand U19807 (N_19807,N_19361,N_19026);
nand U19808 (N_19808,N_19164,N_19349);
xor U19809 (N_19809,N_19335,N_19359);
nor U19810 (N_19810,N_19460,N_19377);
and U19811 (N_19811,N_19283,N_19451);
and U19812 (N_19812,N_19265,N_19341);
and U19813 (N_19813,N_19306,N_19212);
xnor U19814 (N_19814,N_19020,N_19183);
nand U19815 (N_19815,N_19099,N_19072);
and U19816 (N_19816,N_19131,N_19418);
and U19817 (N_19817,N_19268,N_19068);
and U19818 (N_19818,N_19149,N_19210);
xor U19819 (N_19819,N_19108,N_19371);
and U19820 (N_19820,N_19053,N_19028);
and U19821 (N_19821,N_19374,N_19312);
or U19822 (N_19822,N_19057,N_19482);
and U19823 (N_19823,N_19247,N_19485);
nor U19824 (N_19824,N_19341,N_19095);
xor U19825 (N_19825,N_19039,N_19071);
xnor U19826 (N_19826,N_19030,N_19171);
nor U19827 (N_19827,N_19335,N_19125);
or U19828 (N_19828,N_19190,N_19354);
nor U19829 (N_19829,N_19200,N_19150);
xnor U19830 (N_19830,N_19281,N_19176);
and U19831 (N_19831,N_19267,N_19219);
or U19832 (N_19832,N_19200,N_19223);
nor U19833 (N_19833,N_19133,N_19484);
nor U19834 (N_19834,N_19482,N_19065);
and U19835 (N_19835,N_19127,N_19081);
or U19836 (N_19836,N_19105,N_19044);
xor U19837 (N_19837,N_19082,N_19372);
xnor U19838 (N_19838,N_19176,N_19244);
xor U19839 (N_19839,N_19105,N_19232);
nand U19840 (N_19840,N_19226,N_19070);
and U19841 (N_19841,N_19179,N_19183);
nand U19842 (N_19842,N_19453,N_19318);
or U19843 (N_19843,N_19058,N_19302);
nor U19844 (N_19844,N_19032,N_19444);
nand U19845 (N_19845,N_19167,N_19257);
nand U19846 (N_19846,N_19383,N_19189);
xor U19847 (N_19847,N_19251,N_19379);
and U19848 (N_19848,N_19461,N_19451);
or U19849 (N_19849,N_19364,N_19109);
nand U19850 (N_19850,N_19357,N_19371);
and U19851 (N_19851,N_19027,N_19144);
nand U19852 (N_19852,N_19220,N_19182);
or U19853 (N_19853,N_19089,N_19302);
and U19854 (N_19854,N_19468,N_19011);
xnor U19855 (N_19855,N_19301,N_19076);
or U19856 (N_19856,N_19378,N_19158);
or U19857 (N_19857,N_19201,N_19022);
nand U19858 (N_19858,N_19201,N_19053);
xnor U19859 (N_19859,N_19369,N_19385);
nand U19860 (N_19860,N_19211,N_19178);
nand U19861 (N_19861,N_19268,N_19212);
or U19862 (N_19862,N_19165,N_19408);
and U19863 (N_19863,N_19181,N_19258);
and U19864 (N_19864,N_19184,N_19220);
and U19865 (N_19865,N_19120,N_19308);
and U19866 (N_19866,N_19464,N_19424);
and U19867 (N_19867,N_19423,N_19171);
or U19868 (N_19868,N_19241,N_19475);
nor U19869 (N_19869,N_19070,N_19367);
nor U19870 (N_19870,N_19477,N_19159);
and U19871 (N_19871,N_19334,N_19317);
xor U19872 (N_19872,N_19212,N_19419);
nor U19873 (N_19873,N_19471,N_19337);
nor U19874 (N_19874,N_19341,N_19044);
nor U19875 (N_19875,N_19038,N_19008);
xor U19876 (N_19876,N_19176,N_19042);
xnor U19877 (N_19877,N_19388,N_19277);
or U19878 (N_19878,N_19411,N_19444);
or U19879 (N_19879,N_19265,N_19155);
nand U19880 (N_19880,N_19157,N_19113);
xor U19881 (N_19881,N_19164,N_19405);
or U19882 (N_19882,N_19429,N_19411);
nor U19883 (N_19883,N_19256,N_19219);
or U19884 (N_19884,N_19016,N_19494);
nor U19885 (N_19885,N_19471,N_19057);
nand U19886 (N_19886,N_19280,N_19334);
or U19887 (N_19887,N_19259,N_19170);
nor U19888 (N_19888,N_19018,N_19065);
nor U19889 (N_19889,N_19308,N_19108);
xor U19890 (N_19890,N_19058,N_19168);
xor U19891 (N_19891,N_19448,N_19262);
nor U19892 (N_19892,N_19085,N_19367);
and U19893 (N_19893,N_19418,N_19112);
xor U19894 (N_19894,N_19170,N_19256);
and U19895 (N_19895,N_19122,N_19163);
or U19896 (N_19896,N_19131,N_19492);
nand U19897 (N_19897,N_19057,N_19434);
nand U19898 (N_19898,N_19137,N_19232);
nand U19899 (N_19899,N_19085,N_19043);
and U19900 (N_19900,N_19311,N_19039);
and U19901 (N_19901,N_19476,N_19238);
nand U19902 (N_19902,N_19260,N_19148);
nor U19903 (N_19903,N_19134,N_19169);
or U19904 (N_19904,N_19427,N_19368);
nand U19905 (N_19905,N_19037,N_19314);
nand U19906 (N_19906,N_19375,N_19323);
nor U19907 (N_19907,N_19056,N_19111);
nand U19908 (N_19908,N_19104,N_19020);
nor U19909 (N_19909,N_19279,N_19204);
and U19910 (N_19910,N_19281,N_19240);
or U19911 (N_19911,N_19218,N_19120);
xnor U19912 (N_19912,N_19115,N_19292);
xor U19913 (N_19913,N_19303,N_19218);
or U19914 (N_19914,N_19499,N_19448);
and U19915 (N_19915,N_19427,N_19424);
and U19916 (N_19916,N_19136,N_19266);
nor U19917 (N_19917,N_19023,N_19471);
xor U19918 (N_19918,N_19243,N_19085);
or U19919 (N_19919,N_19445,N_19338);
and U19920 (N_19920,N_19189,N_19282);
or U19921 (N_19921,N_19335,N_19399);
and U19922 (N_19922,N_19324,N_19370);
and U19923 (N_19923,N_19301,N_19007);
or U19924 (N_19924,N_19395,N_19293);
and U19925 (N_19925,N_19425,N_19324);
xnor U19926 (N_19926,N_19460,N_19384);
or U19927 (N_19927,N_19061,N_19456);
nand U19928 (N_19928,N_19444,N_19110);
and U19929 (N_19929,N_19319,N_19293);
nand U19930 (N_19930,N_19310,N_19313);
nand U19931 (N_19931,N_19379,N_19145);
or U19932 (N_19932,N_19363,N_19436);
and U19933 (N_19933,N_19391,N_19021);
or U19934 (N_19934,N_19042,N_19471);
nor U19935 (N_19935,N_19308,N_19252);
xor U19936 (N_19936,N_19390,N_19021);
nor U19937 (N_19937,N_19032,N_19035);
nand U19938 (N_19938,N_19496,N_19037);
or U19939 (N_19939,N_19324,N_19267);
and U19940 (N_19940,N_19414,N_19135);
nand U19941 (N_19941,N_19125,N_19466);
nand U19942 (N_19942,N_19146,N_19257);
nor U19943 (N_19943,N_19375,N_19069);
nor U19944 (N_19944,N_19262,N_19073);
and U19945 (N_19945,N_19058,N_19167);
or U19946 (N_19946,N_19278,N_19042);
or U19947 (N_19947,N_19311,N_19351);
and U19948 (N_19948,N_19212,N_19026);
nor U19949 (N_19949,N_19196,N_19496);
nand U19950 (N_19950,N_19046,N_19283);
xnor U19951 (N_19951,N_19067,N_19127);
nor U19952 (N_19952,N_19357,N_19192);
nand U19953 (N_19953,N_19201,N_19359);
or U19954 (N_19954,N_19060,N_19129);
nor U19955 (N_19955,N_19153,N_19436);
xnor U19956 (N_19956,N_19336,N_19327);
nor U19957 (N_19957,N_19013,N_19236);
or U19958 (N_19958,N_19485,N_19017);
or U19959 (N_19959,N_19388,N_19332);
nand U19960 (N_19960,N_19245,N_19012);
or U19961 (N_19961,N_19240,N_19365);
nand U19962 (N_19962,N_19080,N_19408);
or U19963 (N_19963,N_19427,N_19474);
nand U19964 (N_19964,N_19472,N_19060);
or U19965 (N_19965,N_19342,N_19215);
and U19966 (N_19966,N_19469,N_19125);
or U19967 (N_19967,N_19175,N_19140);
or U19968 (N_19968,N_19351,N_19374);
nand U19969 (N_19969,N_19001,N_19322);
and U19970 (N_19970,N_19371,N_19376);
xor U19971 (N_19971,N_19098,N_19065);
nor U19972 (N_19972,N_19364,N_19203);
or U19973 (N_19973,N_19197,N_19351);
or U19974 (N_19974,N_19059,N_19065);
or U19975 (N_19975,N_19358,N_19266);
and U19976 (N_19976,N_19062,N_19186);
nor U19977 (N_19977,N_19208,N_19435);
xor U19978 (N_19978,N_19358,N_19243);
nor U19979 (N_19979,N_19462,N_19472);
nor U19980 (N_19980,N_19448,N_19111);
nand U19981 (N_19981,N_19466,N_19068);
nor U19982 (N_19982,N_19006,N_19379);
nand U19983 (N_19983,N_19169,N_19073);
xor U19984 (N_19984,N_19048,N_19463);
nand U19985 (N_19985,N_19180,N_19399);
nor U19986 (N_19986,N_19446,N_19168);
xnor U19987 (N_19987,N_19018,N_19409);
nor U19988 (N_19988,N_19444,N_19062);
nor U19989 (N_19989,N_19281,N_19236);
or U19990 (N_19990,N_19153,N_19249);
nand U19991 (N_19991,N_19066,N_19289);
and U19992 (N_19992,N_19409,N_19304);
nand U19993 (N_19993,N_19498,N_19028);
or U19994 (N_19994,N_19263,N_19364);
nor U19995 (N_19995,N_19118,N_19045);
and U19996 (N_19996,N_19060,N_19442);
nand U19997 (N_19997,N_19496,N_19129);
nand U19998 (N_19998,N_19433,N_19121);
or U19999 (N_19999,N_19200,N_19084);
or U20000 (N_20000,N_19991,N_19866);
or U20001 (N_20001,N_19590,N_19778);
and U20002 (N_20002,N_19619,N_19714);
and U20003 (N_20003,N_19622,N_19754);
and U20004 (N_20004,N_19730,N_19629);
nor U20005 (N_20005,N_19728,N_19820);
nor U20006 (N_20006,N_19566,N_19620);
nand U20007 (N_20007,N_19780,N_19831);
xor U20008 (N_20008,N_19797,N_19539);
or U20009 (N_20009,N_19654,N_19633);
nor U20010 (N_20010,N_19685,N_19844);
and U20011 (N_20011,N_19549,N_19751);
nand U20012 (N_20012,N_19857,N_19960);
nor U20013 (N_20013,N_19740,N_19998);
xor U20014 (N_20014,N_19707,N_19735);
or U20015 (N_20015,N_19738,N_19529);
xor U20016 (N_20016,N_19647,N_19547);
and U20017 (N_20017,N_19704,N_19631);
nand U20018 (N_20018,N_19625,N_19542);
or U20019 (N_20019,N_19899,N_19979);
and U20020 (N_20020,N_19775,N_19605);
xor U20021 (N_20021,N_19776,N_19750);
and U20022 (N_20022,N_19601,N_19937);
xor U20023 (N_20023,N_19906,N_19962);
nand U20024 (N_20024,N_19944,N_19657);
xor U20025 (N_20025,N_19987,N_19663);
nand U20026 (N_20026,N_19548,N_19798);
and U20027 (N_20027,N_19974,N_19638);
xnor U20028 (N_20028,N_19925,N_19816);
and U20029 (N_20029,N_19560,N_19587);
nor U20030 (N_20030,N_19719,N_19951);
or U20031 (N_20031,N_19992,N_19939);
xnor U20032 (N_20032,N_19867,N_19957);
and U20033 (N_20033,N_19502,N_19597);
nand U20034 (N_20034,N_19881,N_19723);
and U20035 (N_20035,N_19860,N_19990);
or U20036 (N_20036,N_19713,N_19733);
and U20037 (N_20037,N_19655,N_19612);
nand U20038 (N_20038,N_19766,N_19783);
nand U20039 (N_20039,N_19842,N_19912);
or U20040 (N_20040,N_19852,N_19532);
nor U20041 (N_20041,N_19513,N_19642);
or U20042 (N_20042,N_19940,N_19973);
nor U20043 (N_20043,N_19869,N_19941);
nand U20044 (N_20044,N_19607,N_19804);
or U20045 (N_20045,N_19970,N_19569);
nand U20046 (N_20046,N_19986,N_19902);
and U20047 (N_20047,N_19676,N_19672);
and U20048 (N_20048,N_19554,N_19594);
nand U20049 (N_20049,N_19774,N_19661);
and U20050 (N_20050,N_19571,N_19604);
or U20051 (N_20051,N_19829,N_19926);
and U20052 (N_20052,N_19935,N_19512);
xor U20053 (N_20053,N_19561,N_19598);
and U20054 (N_20054,N_19817,N_19834);
or U20055 (N_20055,N_19865,N_19884);
nand U20056 (N_20056,N_19716,N_19602);
xor U20057 (N_20057,N_19916,N_19764);
and U20058 (N_20058,N_19807,N_19706);
or U20059 (N_20059,N_19878,N_19995);
nand U20060 (N_20060,N_19679,N_19737);
xnor U20061 (N_20061,N_19721,N_19837);
and U20062 (N_20062,N_19938,N_19889);
nand U20063 (N_20063,N_19969,N_19507);
nor U20064 (N_20064,N_19755,N_19586);
xnor U20065 (N_20065,N_19806,N_19551);
xor U20066 (N_20066,N_19717,N_19833);
nand U20067 (N_20067,N_19964,N_19989);
or U20068 (N_20068,N_19558,N_19589);
xnor U20069 (N_20069,N_19903,N_19579);
or U20070 (N_20070,N_19967,N_19684);
and U20071 (N_20071,N_19634,N_19680);
nor U20072 (N_20072,N_19736,N_19983);
nor U20073 (N_20073,N_19623,N_19915);
xor U20074 (N_20074,N_19515,N_19825);
or U20075 (N_20075,N_19943,N_19644);
xor U20076 (N_20076,N_19643,N_19729);
or U20077 (N_20077,N_19863,N_19892);
nor U20078 (N_20078,N_19904,N_19870);
xor U20079 (N_20079,N_19799,N_19782);
nor U20080 (N_20080,N_19621,N_19762);
xnor U20081 (N_20081,N_19808,N_19965);
and U20082 (N_20082,N_19699,N_19683);
nor U20083 (N_20083,N_19827,N_19596);
nor U20084 (N_20084,N_19789,N_19653);
or U20085 (N_20085,N_19667,N_19627);
nand U20086 (N_20086,N_19779,N_19618);
xnor U20087 (N_20087,N_19862,N_19763);
nand U20088 (N_20088,N_19841,N_19793);
and U20089 (N_20089,N_19744,N_19811);
xor U20090 (N_20090,N_19993,N_19541);
xor U20091 (N_20091,N_19972,N_19521);
nor U20092 (N_20092,N_19914,N_19896);
xnor U20093 (N_20093,N_19696,N_19981);
or U20094 (N_20094,N_19659,N_19952);
or U20095 (N_20095,N_19947,N_19503);
and U20096 (N_20096,N_19756,N_19879);
nor U20097 (N_20097,N_19978,N_19890);
or U20098 (N_20098,N_19930,N_19765);
nor U20099 (N_20099,N_19709,N_19666);
xor U20100 (N_20100,N_19658,N_19905);
xor U20101 (N_20101,N_19636,N_19800);
and U20102 (N_20102,N_19961,N_19769);
xnor U20103 (N_20103,N_19897,N_19656);
xor U20104 (N_20104,N_19514,N_19574);
xnor U20105 (N_20105,N_19552,N_19641);
xor U20106 (N_20106,N_19767,N_19823);
xnor U20107 (N_20107,N_19877,N_19509);
nand U20108 (N_20108,N_19525,N_19510);
xor U20109 (N_20109,N_19924,N_19985);
or U20110 (N_20110,N_19872,N_19747);
nand U20111 (N_20111,N_19669,N_19893);
nand U20112 (N_20112,N_19847,N_19977);
nand U20113 (N_20113,N_19575,N_19648);
and U20114 (N_20114,N_19535,N_19572);
nand U20115 (N_20115,N_19553,N_19801);
nand U20116 (N_20116,N_19673,N_19523);
xor U20117 (N_20117,N_19874,N_19578);
or U20118 (N_20118,N_19573,N_19888);
or U20119 (N_20119,N_19703,N_19945);
or U20120 (N_20120,N_19805,N_19950);
and U20121 (N_20121,N_19691,N_19843);
nand U20122 (N_20122,N_19570,N_19871);
xnor U20123 (N_20123,N_19649,N_19722);
or U20124 (N_20124,N_19585,N_19745);
and U20125 (N_20125,N_19880,N_19853);
xor U20126 (N_20126,N_19876,N_19671);
xnor U20127 (N_20127,N_19564,N_19791);
and U20128 (N_20128,N_19614,N_19855);
or U20129 (N_20129,N_19505,N_19898);
xnor U20130 (N_20130,N_19997,N_19856);
nand U20131 (N_20131,N_19787,N_19506);
or U20132 (N_20132,N_19908,N_19688);
nand U20133 (N_20133,N_19813,N_19686);
and U20134 (N_20134,N_19556,N_19690);
nor U20135 (N_20135,N_19645,N_19710);
or U20136 (N_20136,N_19768,N_19836);
nor U20137 (N_20137,N_19932,N_19900);
and U20138 (N_20138,N_19694,N_19999);
nand U20139 (N_20139,N_19757,N_19624);
nand U20140 (N_20140,N_19790,N_19803);
nand U20141 (N_20141,N_19581,N_19533);
nor U20142 (N_20142,N_19591,N_19522);
nor U20143 (N_20143,N_19784,N_19753);
or U20144 (N_20144,N_19946,N_19637);
nand U20145 (N_20145,N_19794,N_19785);
xnor U20146 (N_20146,N_19772,N_19527);
nor U20147 (N_20147,N_19802,N_19907);
nor U20148 (N_20148,N_19689,N_19795);
xnor U20149 (N_20149,N_19963,N_19919);
nor U20150 (N_20150,N_19821,N_19859);
or U20151 (N_20151,N_19702,N_19603);
nand U20152 (N_20152,N_19720,N_19832);
nand U20153 (N_20153,N_19885,N_19773);
xnor U20154 (N_20154,N_19557,N_19595);
and U20155 (N_20155,N_19500,N_19968);
nor U20156 (N_20156,N_19909,N_19588);
or U20157 (N_20157,N_19531,N_19749);
nand U20158 (N_20158,N_19913,N_19519);
nand U20159 (N_20159,N_19678,N_19504);
xor U20160 (N_20160,N_19921,N_19718);
xor U20161 (N_20161,N_19727,N_19600);
nor U20162 (N_20162,N_19922,N_19858);
nand U20163 (N_20163,N_19545,N_19695);
nand U20164 (N_20164,N_19501,N_19948);
nand U20165 (N_20165,N_19609,N_19956);
xnor U20166 (N_20166,N_19664,N_19982);
or U20167 (N_20167,N_19810,N_19536);
nand U20168 (N_20168,N_19517,N_19984);
xor U20169 (N_20169,N_19692,N_19777);
or U20170 (N_20170,N_19942,N_19839);
nand U20171 (N_20171,N_19608,N_19838);
or U20172 (N_20172,N_19927,N_19626);
nor U20173 (N_20173,N_19565,N_19910);
nor U20174 (N_20174,N_19819,N_19901);
nand U20175 (N_20175,N_19660,N_19883);
nor U20176 (N_20176,N_19526,N_19953);
and U20177 (N_20177,N_19917,N_19518);
or U20178 (N_20178,N_19891,N_19610);
xor U20179 (N_20179,N_19911,N_19894);
and U20180 (N_20180,N_19534,N_19538);
nor U20181 (N_20181,N_19954,N_19796);
nor U20182 (N_20182,N_19543,N_19611);
xnor U20183 (N_20183,N_19976,N_19630);
nor U20184 (N_20184,N_19849,N_19955);
nand U20185 (N_20185,N_19812,N_19781);
nor U20186 (N_20186,N_19563,N_19725);
xor U20187 (N_20187,N_19786,N_19700);
nor U20188 (N_20188,N_19936,N_19546);
xnor U20189 (N_20189,N_19559,N_19850);
or U20190 (N_20190,N_19818,N_19583);
or U20191 (N_20191,N_19966,N_19923);
nand U20192 (N_20192,N_19606,N_19516);
nor U20193 (N_20193,N_19520,N_19854);
nand U20194 (N_20194,N_19732,N_19652);
or U20195 (N_20195,N_19988,N_19815);
xnor U20196 (N_20196,N_19840,N_19511);
xnor U20197 (N_20197,N_19555,N_19635);
nor U20198 (N_20198,N_19851,N_19712);
xor U20199 (N_20199,N_19931,N_19994);
xnor U20200 (N_20200,N_19741,N_19864);
or U20201 (N_20201,N_19593,N_19846);
or U20202 (N_20202,N_19934,N_19975);
xor U20203 (N_20203,N_19701,N_19592);
or U20204 (N_20204,N_19770,N_19693);
or U20205 (N_20205,N_19668,N_19882);
nor U20206 (N_20206,N_19873,N_19697);
xnor U20207 (N_20207,N_19828,N_19746);
xnor U20208 (N_20208,N_19743,N_19886);
nand U20209 (N_20209,N_19824,N_19996);
and U20210 (N_20210,N_19550,N_19980);
or U20211 (N_20211,N_19698,N_19651);
nand U20212 (N_20212,N_19759,N_19528);
or U20213 (N_20213,N_19567,N_19674);
nor U20214 (N_20214,N_19687,N_19771);
xor U20215 (N_20215,N_19933,N_19662);
nor U20216 (N_20216,N_19568,N_19971);
or U20217 (N_20217,N_19650,N_19675);
or U20218 (N_20218,N_19708,N_19758);
or U20219 (N_20219,N_19848,N_19639);
nor U20220 (N_20220,N_19835,N_19826);
and U20221 (N_20221,N_19734,N_19726);
or U20222 (N_20222,N_19562,N_19613);
or U20223 (N_20223,N_19809,N_19632);
or U20224 (N_20224,N_19949,N_19928);
nor U20225 (N_20225,N_19584,N_19508);
or U20226 (N_20226,N_19616,N_19822);
xnor U20227 (N_20227,N_19861,N_19868);
xor U20228 (N_20228,N_19640,N_19715);
or U20229 (N_20229,N_19761,N_19524);
xor U20230 (N_20230,N_19711,N_19760);
or U20231 (N_20231,N_19918,N_19530);
nand U20232 (N_20232,N_19577,N_19537);
nand U20233 (N_20233,N_19788,N_19959);
xnor U20234 (N_20234,N_19958,N_19544);
nor U20235 (N_20235,N_19929,N_19615);
nor U20236 (N_20236,N_19887,N_19739);
nand U20237 (N_20237,N_19875,N_19731);
xnor U20238 (N_20238,N_19582,N_19895);
nor U20239 (N_20239,N_19599,N_19748);
or U20240 (N_20240,N_19617,N_19540);
nor U20241 (N_20241,N_19742,N_19724);
or U20242 (N_20242,N_19682,N_19580);
nand U20243 (N_20243,N_19830,N_19792);
nor U20244 (N_20244,N_19646,N_19576);
or U20245 (N_20245,N_19665,N_19628);
or U20246 (N_20246,N_19677,N_19845);
xnor U20247 (N_20247,N_19670,N_19752);
nor U20248 (N_20248,N_19920,N_19814);
or U20249 (N_20249,N_19681,N_19705);
and U20250 (N_20250,N_19662,N_19961);
or U20251 (N_20251,N_19771,N_19929);
and U20252 (N_20252,N_19693,N_19730);
and U20253 (N_20253,N_19896,N_19985);
nand U20254 (N_20254,N_19946,N_19511);
nor U20255 (N_20255,N_19513,N_19695);
xnor U20256 (N_20256,N_19757,N_19983);
nand U20257 (N_20257,N_19611,N_19625);
nand U20258 (N_20258,N_19907,N_19752);
xor U20259 (N_20259,N_19804,N_19836);
and U20260 (N_20260,N_19528,N_19649);
or U20261 (N_20261,N_19897,N_19960);
nor U20262 (N_20262,N_19557,N_19797);
nand U20263 (N_20263,N_19774,N_19625);
nor U20264 (N_20264,N_19975,N_19540);
nor U20265 (N_20265,N_19892,N_19843);
nor U20266 (N_20266,N_19838,N_19960);
and U20267 (N_20267,N_19629,N_19676);
nand U20268 (N_20268,N_19635,N_19865);
xor U20269 (N_20269,N_19784,N_19846);
and U20270 (N_20270,N_19509,N_19850);
nor U20271 (N_20271,N_19921,N_19686);
or U20272 (N_20272,N_19811,N_19749);
nand U20273 (N_20273,N_19536,N_19997);
or U20274 (N_20274,N_19569,N_19665);
nor U20275 (N_20275,N_19586,N_19927);
and U20276 (N_20276,N_19717,N_19787);
xor U20277 (N_20277,N_19765,N_19870);
xnor U20278 (N_20278,N_19665,N_19832);
nand U20279 (N_20279,N_19655,N_19638);
nor U20280 (N_20280,N_19940,N_19606);
or U20281 (N_20281,N_19510,N_19537);
xnor U20282 (N_20282,N_19882,N_19822);
xnor U20283 (N_20283,N_19957,N_19967);
nand U20284 (N_20284,N_19686,N_19740);
nor U20285 (N_20285,N_19978,N_19581);
or U20286 (N_20286,N_19685,N_19849);
xnor U20287 (N_20287,N_19647,N_19986);
or U20288 (N_20288,N_19910,N_19728);
nor U20289 (N_20289,N_19627,N_19707);
nor U20290 (N_20290,N_19620,N_19610);
and U20291 (N_20291,N_19639,N_19624);
nand U20292 (N_20292,N_19753,N_19966);
nor U20293 (N_20293,N_19701,N_19833);
nand U20294 (N_20294,N_19875,N_19529);
nor U20295 (N_20295,N_19841,N_19914);
and U20296 (N_20296,N_19575,N_19889);
xnor U20297 (N_20297,N_19630,N_19900);
nor U20298 (N_20298,N_19756,N_19967);
xor U20299 (N_20299,N_19983,N_19651);
nand U20300 (N_20300,N_19868,N_19621);
nor U20301 (N_20301,N_19791,N_19858);
and U20302 (N_20302,N_19762,N_19714);
xor U20303 (N_20303,N_19550,N_19889);
and U20304 (N_20304,N_19511,N_19563);
and U20305 (N_20305,N_19959,N_19587);
or U20306 (N_20306,N_19598,N_19545);
nor U20307 (N_20307,N_19575,N_19607);
nand U20308 (N_20308,N_19784,N_19718);
and U20309 (N_20309,N_19686,N_19587);
nand U20310 (N_20310,N_19585,N_19536);
xnor U20311 (N_20311,N_19602,N_19880);
nand U20312 (N_20312,N_19555,N_19981);
and U20313 (N_20313,N_19794,N_19717);
and U20314 (N_20314,N_19613,N_19620);
or U20315 (N_20315,N_19985,N_19667);
and U20316 (N_20316,N_19969,N_19889);
xor U20317 (N_20317,N_19936,N_19885);
nand U20318 (N_20318,N_19850,N_19746);
nor U20319 (N_20319,N_19732,N_19895);
nand U20320 (N_20320,N_19775,N_19591);
and U20321 (N_20321,N_19632,N_19795);
nand U20322 (N_20322,N_19880,N_19894);
xor U20323 (N_20323,N_19657,N_19683);
and U20324 (N_20324,N_19820,N_19887);
and U20325 (N_20325,N_19748,N_19645);
or U20326 (N_20326,N_19570,N_19948);
nor U20327 (N_20327,N_19652,N_19881);
or U20328 (N_20328,N_19921,N_19907);
xor U20329 (N_20329,N_19577,N_19508);
xor U20330 (N_20330,N_19736,N_19740);
or U20331 (N_20331,N_19734,N_19534);
xnor U20332 (N_20332,N_19527,N_19784);
nor U20333 (N_20333,N_19896,N_19527);
xor U20334 (N_20334,N_19684,N_19971);
and U20335 (N_20335,N_19818,N_19753);
and U20336 (N_20336,N_19926,N_19522);
and U20337 (N_20337,N_19882,N_19933);
or U20338 (N_20338,N_19522,N_19753);
nand U20339 (N_20339,N_19674,N_19960);
and U20340 (N_20340,N_19791,N_19958);
xor U20341 (N_20341,N_19664,N_19870);
nor U20342 (N_20342,N_19670,N_19502);
and U20343 (N_20343,N_19621,N_19708);
nor U20344 (N_20344,N_19625,N_19906);
and U20345 (N_20345,N_19845,N_19821);
nand U20346 (N_20346,N_19762,N_19772);
xnor U20347 (N_20347,N_19889,N_19845);
xnor U20348 (N_20348,N_19604,N_19970);
or U20349 (N_20349,N_19612,N_19921);
xor U20350 (N_20350,N_19649,N_19936);
or U20351 (N_20351,N_19775,N_19978);
and U20352 (N_20352,N_19818,N_19910);
or U20353 (N_20353,N_19968,N_19567);
or U20354 (N_20354,N_19918,N_19609);
or U20355 (N_20355,N_19836,N_19689);
nor U20356 (N_20356,N_19856,N_19557);
or U20357 (N_20357,N_19788,N_19743);
nand U20358 (N_20358,N_19900,N_19689);
nand U20359 (N_20359,N_19527,N_19775);
xor U20360 (N_20360,N_19973,N_19879);
and U20361 (N_20361,N_19570,N_19872);
or U20362 (N_20362,N_19501,N_19560);
xor U20363 (N_20363,N_19732,N_19859);
nor U20364 (N_20364,N_19848,N_19998);
or U20365 (N_20365,N_19682,N_19810);
and U20366 (N_20366,N_19992,N_19949);
xnor U20367 (N_20367,N_19799,N_19577);
nand U20368 (N_20368,N_19521,N_19587);
xnor U20369 (N_20369,N_19716,N_19950);
nand U20370 (N_20370,N_19669,N_19616);
nor U20371 (N_20371,N_19782,N_19670);
or U20372 (N_20372,N_19905,N_19698);
xnor U20373 (N_20373,N_19841,N_19743);
or U20374 (N_20374,N_19595,N_19964);
and U20375 (N_20375,N_19577,N_19886);
and U20376 (N_20376,N_19843,N_19720);
nand U20377 (N_20377,N_19836,N_19520);
or U20378 (N_20378,N_19799,N_19559);
or U20379 (N_20379,N_19878,N_19845);
or U20380 (N_20380,N_19562,N_19568);
nor U20381 (N_20381,N_19804,N_19588);
or U20382 (N_20382,N_19757,N_19878);
and U20383 (N_20383,N_19823,N_19685);
or U20384 (N_20384,N_19634,N_19878);
xnor U20385 (N_20385,N_19762,N_19541);
nand U20386 (N_20386,N_19875,N_19902);
and U20387 (N_20387,N_19884,N_19604);
nand U20388 (N_20388,N_19502,N_19775);
and U20389 (N_20389,N_19631,N_19966);
nand U20390 (N_20390,N_19764,N_19813);
nand U20391 (N_20391,N_19617,N_19837);
or U20392 (N_20392,N_19732,N_19919);
or U20393 (N_20393,N_19819,N_19909);
nand U20394 (N_20394,N_19630,N_19868);
and U20395 (N_20395,N_19952,N_19760);
nor U20396 (N_20396,N_19528,N_19633);
nor U20397 (N_20397,N_19944,N_19809);
xor U20398 (N_20398,N_19855,N_19749);
and U20399 (N_20399,N_19878,N_19893);
nand U20400 (N_20400,N_19805,N_19940);
nor U20401 (N_20401,N_19658,N_19618);
and U20402 (N_20402,N_19506,N_19694);
or U20403 (N_20403,N_19745,N_19917);
nor U20404 (N_20404,N_19617,N_19577);
and U20405 (N_20405,N_19836,N_19941);
nor U20406 (N_20406,N_19975,N_19547);
nor U20407 (N_20407,N_19551,N_19529);
or U20408 (N_20408,N_19806,N_19566);
or U20409 (N_20409,N_19787,N_19619);
xor U20410 (N_20410,N_19607,N_19742);
xor U20411 (N_20411,N_19958,N_19899);
nand U20412 (N_20412,N_19505,N_19652);
nand U20413 (N_20413,N_19504,N_19953);
and U20414 (N_20414,N_19655,N_19639);
nor U20415 (N_20415,N_19877,N_19809);
xor U20416 (N_20416,N_19877,N_19766);
nand U20417 (N_20417,N_19910,N_19556);
and U20418 (N_20418,N_19678,N_19505);
and U20419 (N_20419,N_19683,N_19506);
nor U20420 (N_20420,N_19769,N_19621);
nor U20421 (N_20421,N_19905,N_19662);
or U20422 (N_20422,N_19725,N_19635);
and U20423 (N_20423,N_19856,N_19797);
nor U20424 (N_20424,N_19805,N_19749);
and U20425 (N_20425,N_19697,N_19711);
nor U20426 (N_20426,N_19993,N_19801);
nand U20427 (N_20427,N_19881,N_19859);
and U20428 (N_20428,N_19502,N_19814);
or U20429 (N_20429,N_19570,N_19848);
nor U20430 (N_20430,N_19951,N_19864);
nand U20431 (N_20431,N_19953,N_19981);
or U20432 (N_20432,N_19742,N_19894);
nand U20433 (N_20433,N_19722,N_19787);
nand U20434 (N_20434,N_19571,N_19988);
nor U20435 (N_20435,N_19856,N_19835);
xor U20436 (N_20436,N_19557,N_19605);
nor U20437 (N_20437,N_19932,N_19728);
xor U20438 (N_20438,N_19714,N_19505);
and U20439 (N_20439,N_19649,N_19790);
nor U20440 (N_20440,N_19791,N_19658);
nor U20441 (N_20441,N_19537,N_19966);
nand U20442 (N_20442,N_19830,N_19873);
nand U20443 (N_20443,N_19950,N_19545);
xor U20444 (N_20444,N_19894,N_19750);
nor U20445 (N_20445,N_19970,N_19849);
xor U20446 (N_20446,N_19908,N_19580);
xor U20447 (N_20447,N_19739,N_19904);
nor U20448 (N_20448,N_19818,N_19511);
or U20449 (N_20449,N_19678,N_19704);
xnor U20450 (N_20450,N_19890,N_19583);
nand U20451 (N_20451,N_19823,N_19922);
or U20452 (N_20452,N_19592,N_19872);
or U20453 (N_20453,N_19777,N_19924);
nand U20454 (N_20454,N_19690,N_19589);
or U20455 (N_20455,N_19796,N_19724);
nor U20456 (N_20456,N_19943,N_19511);
xnor U20457 (N_20457,N_19962,N_19827);
and U20458 (N_20458,N_19867,N_19690);
and U20459 (N_20459,N_19847,N_19848);
xor U20460 (N_20460,N_19766,N_19661);
or U20461 (N_20461,N_19598,N_19992);
and U20462 (N_20462,N_19741,N_19899);
xor U20463 (N_20463,N_19671,N_19574);
or U20464 (N_20464,N_19644,N_19992);
nor U20465 (N_20465,N_19712,N_19998);
nand U20466 (N_20466,N_19615,N_19921);
and U20467 (N_20467,N_19944,N_19503);
xor U20468 (N_20468,N_19797,N_19741);
nand U20469 (N_20469,N_19641,N_19989);
nand U20470 (N_20470,N_19978,N_19553);
or U20471 (N_20471,N_19871,N_19699);
or U20472 (N_20472,N_19843,N_19870);
xor U20473 (N_20473,N_19895,N_19654);
and U20474 (N_20474,N_19834,N_19607);
xor U20475 (N_20475,N_19956,N_19514);
or U20476 (N_20476,N_19907,N_19596);
and U20477 (N_20477,N_19970,N_19750);
and U20478 (N_20478,N_19674,N_19506);
nand U20479 (N_20479,N_19542,N_19937);
nand U20480 (N_20480,N_19577,N_19549);
or U20481 (N_20481,N_19508,N_19932);
or U20482 (N_20482,N_19790,N_19727);
nor U20483 (N_20483,N_19546,N_19966);
or U20484 (N_20484,N_19820,N_19513);
xor U20485 (N_20485,N_19808,N_19730);
and U20486 (N_20486,N_19542,N_19629);
nand U20487 (N_20487,N_19928,N_19881);
and U20488 (N_20488,N_19624,N_19593);
xor U20489 (N_20489,N_19796,N_19725);
nor U20490 (N_20490,N_19921,N_19926);
nand U20491 (N_20491,N_19942,N_19781);
xnor U20492 (N_20492,N_19706,N_19673);
and U20493 (N_20493,N_19637,N_19630);
xor U20494 (N_20494,N_19936,N_19679);
nor U20495 (N_20495,N_19523,N_19833);
nand U20496 (N_20496,N_19996,N_19950);
and U20497 (N_20497,N_19856,N_19673);
or U20498 (N_20498,N_19874,N_19774);
nand U20499 (N_20499,N_19979,N_19985);
xor U20500 (N_20500,N_20482,N_20377);
or U20501 (N_20501,N_20126,N_20316);
nor U20502 (N_20502,N_20157,N_20067);
xor U20503 (N_20503,N_20446,N_20308);
or U20504 (N_20504,N_20251,N_20434);
nor U20505 (N_20505,N_20436,N_20419);
xor U20506 (N_20506,N_20116,N_20256);
or U20507 (N_20507,N_20042,N_20315);
nand U20508 (N_20508,N_20101,N_20100);
xor U20509 (N_20509,N_20132,N_20337);
nand U20510 (N_20510,N_20295,N_20466);
nor U20511 (N_20511,N_20254,N_20303);
or U20512 (N_20512,N_20069,N_20203);
or U20513 (N_20513,N_20387,N_20223);
xor U20514 (N_20514,N_20052,N_20189);
nor U20515 (N_20515,N_20476,N_20334);
and U20516 (N_20516,N_20089,N_20168);
and U20517 (N_20517,N_20006,N_20452);
nor U20518 (N_20518,N_20267,N_20495);
and U20519 (N_20519,N_20394,N_20141);
and U20520 (N_20520,N_20226,N_20428);
nor U20521 (N_20521,N_20172,N_20301);
or U20522 (N_20522,N_20230,N_20079);
and U20523 (N_20523,N_20487,N_20087);
xor U20524 (N_20524,N_20348,N_20444);
xor U20525 (N_20525,N_20182,N_20139);
and U20526 (N_20526,N_20043,N_20094);
nor U20527 (N_20527,N_20276,N_20453);
xor U20528 (N_20528,N_20137,N_20237);
and U20529 (N_20529,N_20107,N_20265);
nor U20530 (N_20530,N_20386,N_20218);
and U20531 (N_20531,N_20460,N_20366);
nor U20532 (N_20532,N_20361,N_20411);
nor U20533 (N_20533,N_20481,N_20472);
nand U20534 (N_20534,N_20369,N_20117);
xor U20535 (N_20535,N_20022,N_20349);
or U20536 (N_20536,N_20469,N_20364);
nor U20537 (N_20537,N_20028,N_20129);
and U20538 (N_20538,N_20260,N_20128);
and U20539 (N_20539,N_20220,N_20017);
and U20540 (N_20540,N_20246,N_20153);
or U20541 (N_20541,N_20216,N_20156);
and U20542 (N_20542,N_20441,N_20065);
nor U20543 (N_20543,N_20140,N_20282);
xnor U20544 (N_20544,N_20414,N_20468);
xor U20545 (N_20545,N_20484,N_20373);
nor U20546 (N_20546,N_20328,N_20071);
nor U20547 (N_20547,N_20410,N_20447);
xor U20548 (N_20548,N_20335,N_20143);
xor U20549 (N_20549,N_20241,N_20381);
xnor U20550 (N_20550,N_20380,N_20086);
nor U20551 (N_20551,N_20025,N_20463);
xor U20552 (N_20552,N_20073,N_20102);
or U20553 (N_20553,N_20440,N_20014);
and U20554 (N_20554,N_20290,N_20286);
and U20555 (N_20555,N_20329,N_20109);
or U20556 (N_20556,N_20376,N_20046);
nor U20557 (N_20557,N_20471,N_20355);
or U20558 (N_20558,N_20291,N_20059);
xor U20559 (N_20559,N_20106,N_20161);
or U20560 (N_20560,N_20357,N_20420);
and U20561 (N_20561,N_20180,N_20389);
xor U20562 (N_20562,N_20352,N_20345);
and U20563 (N_20563,N_20339,N_20114);
and U20564 (N_20564,N_20062,N_20397);
nand U20565 (N_20565,N_20298,N_20279);
nand U20566 (N_20566,N_20047,N_20407);
xor U20567 (N_20567,N_20125,N_20497);
nand U20568 (N_20568,N_20217,N_20206);
nor U20569 (N_20569,N_20375,N_20347);
nand U20570 (N_20570,N_20383,N_20098);
and U20571 (N_20571,N_20091,N_20020);
nor U20572 (N_20572,N_20127,N_20204);
xnor U20573 (N_20573,N_20242,N_20494);
nor U20574 (N_20574,N_20437,N_20296);
xor U20575 (N_20575,N_20036,N_20270);
and U20576 (N_20576,N_20198,N_20031);
nor U20577 (N_20577,N_20038,N_20093);
nor U20578 (N_20578,N_20372,N_20451);
xor U20579 (N_20579,N_20273,N_20278);
and U20580 (N_20580,N_20297,N_20262);
and U20581 (N_20581,N_20430,N_20341);
xor U20582 (N_20582,N_20388,N_20259);
and U20583 (N_20583,N_20008,N_20148);
xnor U20584 (N_20584,N_20121,N_20370);
or U20585 (N_20585,N_20338,N_20299);
and U20586 (N_20586,N_20418,N_20310);
and U20587 (N_20587,N_20110,N_20219);
and U20588 (N_20588,N_20099,N_20177);
nand U20589 (N_20589,N_20231,N_20212);
nor U20590 (N_20590,N_20443,N_20393);
nor U20591 (N_20591,N_20056,N_20200);
and U20592 (N_20592,N_20272,N_20408);
nor U20593 (N_20593,N_20285,N_20435);
xor U20594 (N_20594,N_20039,N_20225);
nand U20595 (N_20595,N_20068,N_20354);
or U20596 (N_20596,N_20123,N_20274);
nand U20597 (N_20597,N_20084,N_20283);
and U20598 (N_20598,N_20258,N_20379);
nand U20599 (N_20599,N_20007,N_20331);
nor U20600 (N_20600,N_20240,N_20118);
xnor U20601 (N_20601,N_20485,N_20187);
or U20602 (N_20602,N_20247,N_20122);
nor U20603 (N_20603,N_20064,N_20045);
nand U20604 (N_20604,N_20088,N_20188);
and U20605 (N_20605,N_20488,N_20422);
and U20606 (N_20606,N_20350,N_20384);
or U20607 (N_20607,N_20374,N_20176);
nor U20608 (N_20608,N_20314,N_20077);
and U20609 (N_20609,N_20277,N_20103);
nand U20610 (N_20610,N_20261,N_20238);
or U20611 (N_20611,N_20300,N_20095);
nor U20612 (N_20612,N_20013,N_20306);
and U20613 (N_20613,N_20417,N_20433);
nand U20614 (N_20614,N_20210,N_20054);
xor U20615 (N_20615,N_20367,N_20213);
or U20616 (N_20616,N_20183,N_20409);
nand U20617 (N_20617,N_20281,N_20326);
nand U20618 (N_20618,N_20015,N_20343);
nand U20619 (N_20619,N_20138,N_20191);
xnor U20620 (N_20620,N_20236,N_20131);
nand U20621 (N_20621,N_20147,N_20021);
or U20622 (N_20622,N_20060,N_20235);
nand U20623 (N_20623,N_20169,N_20197);
or U20624 (N_20624,N_20458,N_20112);
or U20625 (N_20625,N_20181,N_20185);
and U20626 (N_20626,N_20423,N_20294);
and U20627 (N_20627,N_20150,N_20351);
or U20628 (N_20628,N_20074,N_20319);
or U20629 (N_20629,N_20465,N_20461);
or U20630 (N_20630,N_20392,N_20493);
nand U20631 (N_20631,N_20082,N_20224);
or U20632 (N_20632,N_20041,N_20229);
xor U20633 (N_20633,N_20416,N_20199);
nor U20634 (N_20634,N_20317,N_20269);
or U20635 (N_20635,N_20280,N_20111);
nor U20636 (N_20636,N_20255,N_20403);
or U20637 (N_20637,N_20234,N_20429);
or U20638 (N_20638,N_20340,N_20201);
and U20639 (N_20639,N_20450,N_20344);
and U20640 (N_20640,N_20405,N_20080);
xnor U20641 (N_20641,N_20134,N_20214);
nor U20642 (N_20642,N_20413,N_20108);
nor U20643 (N_20643,N_20104,N_20195);
nand U20644 (N_20644,N_20426,N_20336);
and U20645 (N_20645,N_20005,N_20342);
xor U20646 (N_20646,N_20479,N_20034);
and U20647 (N_20647,N_20090,N_20402);
or U20648 (N_20648,N_20412,N_20467);
and U20649 (N_20649,N_20268,N_20391);
xnor U20650 (N_20650,N_20215,N_20368);
or U20651 (N_20651,N_20164,N_20400);
nand U20652 (N_20652,N_20385,N_20478);
xnor U20653 (N_20653,N_20167,N_20390);
xor U20654 (N_20654,N_20012,N_20371);
nor U20655 (N_20655,N_20055,N_20002);
or U20656 (N_20656,N_20033,N_20320);
or U20657 (N_20657,N_20119,N_20211);
nor U20658 (N_20658,N_20027,N_20486);
nand U20659 (N_20659,N_20026,N_20072);
nor U20660 (N_20660,N_20232,N_20162);
nand U20661 (N_20661,N_20222,N_20186);
nand U20662 (N_20662,N_20442,N_20154);
or U20663 (N_20663,N_20304,N_20019);
and U20664 (N_20664,N_20083,N_20023);
xnor U20665 (N_20665,N_20401,N_20016);
or U20666 (N_20666,N_20445,N_20130);
and U20667 (N_20667,N_20010,N_20323);
and U20668 (N_20668,N_20459,N_20178);
xor U20669 (N_20669,N_20321,N_20205);
nor U20670 (N_20670,N_20166,N_20480);
xnor U20671 (N_20671,N_20075,N_20264);
and U20672 (N_20672,N_20159,N_20040);
and U20673 (N_20673,N_20302,N_20271);
and U20674 (N_20674,N_20058,N_20096);
nor U20675 (N_20675,N_20029,N_20208);
nor U20676 (N_20676,N_20492,N_20454);
nand U20677 (N_20677,N_20170,N_20160);
or U20678 (N_20678,N_20105,N_20000);
xnor U20679 (N_20679,N_20145,N_20003);
or U20680 (N_20680,N_20032,N_20318);
xor U20681 (N_20681,N_20289,N_20477);
nor U20682 (N_20682,N_20490,N_20356);
nand U20683 (N_20683,N_20312,N_20037);
or U20684 (N_20684,N_20171,N_20050);
nand U20685 (N_20685,N_20146,N_20483);
or U20686 (N_20686,N_20209,N_20253);
nand U20687 (N_20687,N_20174,N_20024);
xnor U20688 (N_20688,N_20395,N_20498);
nor U20689 (N_20689,N_20250,N_20382);
xor U20690 (N_20690,N_20163,N_20475);
nand U20691 (N_20691,N_20462,N_20142);
or U20692 (N_20692,N_20473,N_20081);
nand U20693 (N_20693,N_20070,N_20158);
nor U20694 (N_20694,N_20049,N_20425);
xnor U20695 (N_20695,N_20057,N_20360);
xnor U20696 (N_20696,N_20194,N_20252);
or U20697 (N_20697,N_20001,N_20424);
or U20698 (N_20698,N_20358,N_20439);
or U20699 (N_20699,N_20061,N_20053);
xor U20700 (N_20700,N_20115,N_20149);
and U20701 (N_20701,N_20421,N_20399);
xor U20702 (N_20702,N_20233,N_20438);
and U20703 (N_20703,N_20018,N_20085);
and U20704 (N_20704,N_20307,N_20151);
nor U20705 (N_20705,N_20193,N_20097);
and U20706 (N_20706,N_20243,N_20155);
or U20707 (N_20707,N_20152,N_20431);
nand U20708 (N_20708,N_20359,N_20489);
xnor U20709 (N_20709,N_20491,N_20406);
nor U20710 (N_20710,N_20333,N_20353);
and U20711 (N_20711,N_20190,N_20136);
nand U20712 (N_20712,N_20030,N_20044);
and U20713 (N_20713,N_20365,N_20474);
nor U20714 (N_20714,N_20207,N_20248);
nor U20715 (N_20715,N_20292,N_20324);
and U20716 (N_20716,N_20184,N_20288);
and U20717 (N_20717,N_20228,N_20249);
or U20718 (N_20718,N_20470,N_20245);
or U20719 (N_20719,N_20266,N_20263);
or U20720 (N_20720,N_20448,N_20457);
or U20721 (N_20721,N_20396,N_20332);
nor U20722 (N_20722,N_20165,N_20415);
nor U20723 (N_20723,N_20133,N_20309);
or U20724 (N_20724,N_20311,N_20051);
nand U20725 (N_20725,N_20404,N_20293);
nand U20726 (N_20726,N_20427,N_20244);
and U20727 (N_20727,N_20092,N_20124);
xnor U20728 (N_20728,N_20432,N_20192);
nand U20729 (N_20729,N_20257,N_20196);
xor U20730 (N_20730,N_20313,N_20035);
xor U20731 (N_20731,N_20179,N_20449);
nand U20732 (N_20732,N_20120,N_20456);
and U20733 (N_20733,N_20066,N_20284);
nor U20734 (N_20734,N_20239,N_20113);
nand U20735 (N_20735,N_20078,N_20322);
or U20736 (N_20736,N_20004,N_20076);
nor U20737 (N_20737,N_20202,N_20011);
nand U20738 (N_20738,N_20398,N_20327);
and U20739 (N_20739,N_20378,N_20175);
or U20740 (N_20740,N_20221,N_20330);
xnor U20741 (N_20741,N_20362,N_20009);
and U20742 (N_20742,N_20144,N_20173);
nand U20743 (N_20743,N_20455,N_20305);
and U20744 (N_20744,N_20346,N_20496);
xnor U20745 (N_20745,N_20048,N_20135);
or U20746 (N_20746,N_20227,N_20363);
and U20747 (N_20747,N_20063,N_20464);
or U20748 (N_20748,N_20325,N_20499);
and U20749 (N_20749,N_20287,N_20275);
nor U20750 (N_20750,N_20093,N_20138);
and U20751 (N_20751,N_20475,N_20073);
and U20752 (N_20752,N_20073,N_20281);
xnor U20753 (N_20753,N_20095,N_20222);
nand U20754 (N_20754,N_20251,N_20227);
nand U20755 (N_20755,N_20421,N_20019);
or U20756 (N_20756,N_20068,N_20387);
xor U20757 (N_20757,N_20342,N_20306);
xor U20758 (N_20758,N_20475,N_20318);
or U20759 (N_20759,N_20459,N_20010);
and U20760 (N_20760,N_20228,N_20197);
nor U20761 (N_20761,N_20075,N_20379);
or U20762 (N_20762,N_20155,N_20138);
or U20763 (N_20763,N_20185,N_20103);
nand U20764 (N_20764,N_20247,N_20128);
nor U20765 (N_20765,N_20204,N_20032);
and U20766 (N_20766,N_20440,N_20065);
xnor U20767 (N_20767,N_20483,N_20222);
nand U20768 (N_20768,N_20051,N_20108);
and U20769 (N_20769,N_20391,N_20261);
xnor U20770 (N_20770,N_20199,N_20295);
or U20771 (N_20771,N_20206,N_20343);
nor U20772 (N_20772,N_20387,N_20090);
xor U20773 (N_20773,N_20105,N_20251);
or U20774 (N_20774,N_20340,N_20184);
and U20775 (N_20775,N_20129,N_20015);
xor U20776 (N_20776,N_20492,N_20399);
and U20777 (N_20777,N_20349,N_20187);
nand U20778 (N_20778,N_20266,N_20029);
nor U20779 (N_20779,N_20052,N_20290);
nand U20780 (N_20780,N_20143,N_20360);
and U20781 (N_20781,N_20295,N_20270);
xor U20782 (N_20782,N_20013,N_20452);
nor U20783 (N_20783,N_20190,N_20431);
xor U20784 (N_20784,N_20134,N_20110);
nand U20785 (N_20785,N_20271,N_20180);
nor U20786 (N_20786,N_20406,N_20192);
xnor U20787 (N_20787,N_20071,N_20353);
or U20788 (N_20788,N_20193,N_20419);
nor U20789 (N_20789,N_20268,N_20329);
nor U20790 (N_20790,N_20102,N_20096);
xnor U20791 (N_20791,N_20242,N_20089);
nor U20792 (N_20792,N_20079,N_20045);
or U20793 (N_20793,N_20214,N_20293);
xnor U20794 (N_20794,N_20029,N_20000);
or U20795 (N_20795,N_20453,N_20215);
nand U20796 (N_20796,N_20025,N_20120);
or U20797 (N_20797,N_20438,N_20121);
or U20798 (N_20798,N_20267,N_20371);
or U20799 (N_20799,N_20192,N_20357);
or U20800 (N_20800,N_20214,N_20374);
nand U20801 (N_20801,N_20463,N_20074);
or U20802 (N_20802,N_20306,N_20457);
nor U20803 (N_20803,N_20479,N_20025);
and U20804 (N_20804,N_20044,N_20452);
xnor U20805 (N_20805,N_20483,N_20105);
or U20806 (N_20806,N_20294,N_20466);
nand U20807 (N_20807,N_20400,N_20345);
nor U20808 (N_20808,N_20395,N_20222);
nor U20809 (N_20809,N_20142,N_20112);
or U20810 (N_20810,N_20235,N_20309);
xor U20811 (N_20811,N_20408,N_20210);
or U20812 (N_20812,N_20255,N_20297);
xor U20813 (N_20813,N_20025,N_20317);
nand U20814 (N_20814,N_20478,N_20228);
nor U20815 (N_20815,N_20126,N_20207);
or U20816 (N_20816,N_20155,N_20199);
xnor U20817 (N_20817,N_20174,N_20007);
nand U20818 (N_20818,N_20277,N_20304);
nor U20819 (N_20819,N_20136,N_20401);
nand U20820 (N_20820,N_20064,N_20008);
nor U20821 (N_20821,N_20015,N_20226);
and U20822 (N_20822,N_20183,N_20248);
or U20823 (N_20823,N_20384,N_20297);
nand U20824 (N_20824,N_20285,N_20291);
and U20825 (N_20825,N_20142,N_20359);
nand U20826 (N_20826,N_20247,N_20180);
nor U20827 (N_20827,N_20169,N_20296);
and U20828 (N_20828,N_20150,N_20067);
nor U20829 (N_20829,N_20391,N_20040);
nor U20830 (N_20830,N_20384,N_20483);
nand U20831 (N_20831,N_20049,N_20371);
nor U20832 (N_20832,N_20026,N_20219);
and U20833 (N_20833,N_20341,N_20328);
xor U20834 (N_20834,N_20156,N_20444);
nand U20835 (N_20835,N_20449,N_20197);
and U20836 (N_20836,N_20443,N_20342);
nand U20837 (N_20837,N_20195,N_20063);
xor U20838 (N_20838,N_20022,N_20303);
xnor U20839 (N_20839,N_20185,N_20260);
xnor U20840 (N_20840,N_20178,N_20187);
xor U20841 (N_20841,N_20477,N_20347);
xor U20842 (N_20842,N_20152,N_20048);
and U20843 (N_20843,N_20148,N_20029);
and U20844 (N_20844,N_20280,N_20376);
and U20845 (N_20845,N_20128,N_20013);
nand U20846 (N_20846,N_20446,N_20458);
and U20847 (N_20847,N_20279,N_20451);
nor U20848 (N_20848,N_20453,N_20479);
or U20849 (N_20849,N_20162,N_20333);
nand U20850 (N_20850,N_20076,N_20200);
nand U20851 (N_20851,N_20002,N_20062);
or U20852 (N_20852,N_20400,N_20192);
nor U20853 (N_20853,N_20114,N_20165);
nor U20854 (N_20854,N_20301,N_20115);
nand U20855 (N_20855,N_20277,N_20166);
nor U20856 (N_20856,N_20060,N_20083);
or U20857 (N_20857,N_20482,N_20361);
nor U20858 (N_20858,N_20446,N_20153);
or U20859 (N_20859,N_20184,N_20420);
and U20860 (N_20860,N_20431,N_20115);
or U20861 (N_20861,N_20462,N_20157);
nor U20862 (N_20862,N_20345,N_20465);
or U20863 (N_20863,N_20362,N_20497);
and U20864 (N_20864,N_20178,N_20392);
and U20865 (N_20865,N_20346,N_20041);
nor U20866 (N_20866,N_20190,N_20407);
or U20867 (N_20867,N_20323,N_20486);
nor U20868 (N_20868,N_20447,N_20199);
nand U20869 (N_20869,N_20237,N_20206);
and U20870 (N_20870,N_20219,N_20173);
and U20871 (N_20871,N_20080,N_20393);
nor U20872 (N_20872,N_20483,N_20283);
and U20873 (N_20873,N_20355,N_20378);
and U20874 (N_20874,N_20413,N_20043);
and U20875 (N_20875,N_20419,N_20238);
or U20876 (N_20876,N_20122,N_20016);
and U20877 (N_20877,N_20329,N_20113);
and U20878 (N_20878,N_20140,N_20288);
nand U20879 (N_20879,N_20498,N_20323);
xnor U20880 (N_20880,N_20253,N_20479);
or U20881 (N_20881,N_20051,N_20197);
nor U20882 (N_20882,N_20408,N_20498);
and U20883 (N_20883,N_20300,N_20440);
nor U20884 (N_20884,N_20212,N_20404);
nor U20885 (N_20885,N_20199,N_20367);
nor U20886 (N_20886,N_20172,N_20112);
or U20887 (N_20887,N_20297,N_20241);
and U20888 (N_20888,N_20263,N_20370);
or U20889 (N_20889,N_20321,N_20323);
xnor U20890 (N_20890,N_20188,N_20202);
and U20891 (N_20891,N_20316,N_20449);
nand U20892 (N_20892,N_20370,N_20120);
or U20893 (N_20893,N_20410,N_20422);
xnor U20894 (N_20894,N_20225,N_20001);
or U20895 (N_20895,N_20316,N_20217);
or U20896 (N_20896,N_20470,N_20209);
xnor U20897 (N_20897,N_20254,N_20204);
nor U20898 (N_20898,N_20381,N_20252);
xor U20899 (N_20899,N_20300,N_20335);
xor U20900 (N_20900,N_20217,N_20490);
or U20901 (N_20901,N_20223,N_20159);
or U20902 (N_20902,N_20204,N_20329);
or U20903 (N_20903,N_20280,N_20467);
and U20904 (N_20904,N_20280,N_20150);
nand U20905 (N_20905,N_20138,N_20390);
xor U20906 (N_20906,N_20212,N_20070);
xor U20907 (N_20907,N_20463,N_20407);
and U20908 (N_20908,N_20046,N_20238);
or U20909 (N_20909,N_20264,N_20427);
nand U20910 (N_20910,N_20010,N_20220);
nor U20911 (N_20911,N_20099,N_20083);
nand U20912 (N_20912,N_20442,N_20170);
or U20913 (N_20913,N_20148,N_20108);
nand U20914 (N_20914,N_20107,N_20131);
xnor U20915 (N_20915,N_20247,N_20093);
nand U20916 (N_20916,N_20220,N_20163);
xor U20917 (N_20917,N_20101,N_20034);
nand U20918 (N_20918,N_20198,N_20437);
and U20919 (N_20919,N_20418,N_20053);
and U20920 (N_20920,N_20460,N_20335);
nor U20921 (N_20921,N_20294,N_20328);
or U20922 (N_20922,N_20243,N_20453);
and U20923 (N_20923,N_20192,N_20465);
xnor U20924 (N_20924,N_20210,N_20469);
and U20925 (N_20925,N_20259,N_20027);
and U20926 (N_20926,N_20057,N_20215);
and U20927 (N_20927,N_20445,N_20428);
xnor U20928 (N_20928,N_20142,N_20258);
and U20929 (N_20929,N_20335,N_20154);
nand U20930 (N_20930,N_20035,N_20270);
nand U20931 (N_20931,N_20035,N_20232);
or U20932 (N_20932,N_20126,N_20427);
and U20933 (N_20933,N_20068,N_20470);
nand U20934 (N_20934,N_20467,N_20087);
nand U20935 (N_20935,N_20099,N_20478);
nand U20936 (N_20936,N_20231,N_20103);
nor U20937 (N_20937,N_20464,N_20111);
nand U20938 (N_20938,N_20369,N_20148);
and U20939 (N_20939,N_20276,N_20190);
and U20940 (N_20940,N_20046,N_20324);
xnor U20941 (N_20941,N_20291,N_20267);
xnor U20942 (N_20942,N_20209,N_20367);
xnor U20943 (N_20943,N_20190,N_20279);
and U20944 (N_20944,N_20430,N_20173);
and U20945 (N_20945,N_20169,N_20205);
and U20946 (N_20946,N_20120,N_20069);
xor U20947 (N_20947,N_20141,N_20454);
or U20948 (N_20948,N_20432,N_20072);
nand U20949 (N_20949,N_20455,N_20327);
nand U20950 (N_20950,N_20101,N_20189);
or U20951 (N_20951,N_20028,N_20109);
xnor U20952 (N_20952,N_20187,N_20097);
nor U20953 (N_20953,N_20109,N_20366);
xor U20954 (N_20954,N_20064,N_20300);
xnor U20955 (N_20955,N_20229,N_20499);
nand U20956 (N_20956,N_20375,N_20162);
nor U20957 (N_20957,N_20210,N_20092);
and U20958 (N_20958,N_20096,N_20283);
and U20959 (N_20959,N_20018,N_20113);
and U20960 (N_20960,N_20266,N_20302);
nand U20961 (N_20961,N_20391,N_20023);
or U20962 (N_20962,N_20029,N_20272);
or U20963 (N_20963,N_20018,N_20409);
or U20964 (N_20964,N_20359,N_20111);
xnor U20965 (N_20965,N_20005,N_20397);
or U20966 (N_20966,N_20462,N_20228);
and U20967 (N_20967,N_20087,N_20459);
nor U20968 (N_20968,N_20271,N_20140);
xor U20969 (N_20969,N_20474,N_20243);
or U20970 (N_20970,N_20279,N_20499);
nand U20971 (N_20971,N_20120,N_20104);
and U20972 (N_20972,N_20168,N_20132);
nand U20973 (N_20973,N_20111,N_20477);
and U20974 (N_20974,N_20183,N_20497);
nor U20975 (N_20975,N_20186,N_20226);
or U20976 (N_20976,N_20025,N_20128);
or U20977 (N_20977,N_20137,N_20269);
xnor U20978 (N_20978,N_20405,N_20452);
nor U20979 (N_20979,N_20223,N_20262);
xor U20980 (N_20980,N_20352,N_20385);
nor U20981 (N_20981,N_20399,N_20176);
nand U20982 (N_20982,N_20326,N_20432);
nand U20983 (N_20983,N_20033,N_20357);
xor U20984 (N_20984,N_20462,N_20294);
or U20985 (N_20985,N_20248,N_20134);
or U20986 (N_20986,N_20215,N_20049);
nor U20987 (N_20987,N_20323,N_20424);
nor U20988 (N_20988,N_20496,N_20477);
xnor U20989 (N_20989,N_20092,N_20091);
nor U20990 (N_20990,N_20259,N_20269);
nor U20991 (N_20991,N_20216,N_20253);
xor U20992 (N_20992,N_20379,N_20355);
nor U20993 (N_20993,N_20329,N_20017);
xnor U20994 (N_20994,N_20423,N_20244);
nor U20995 (N_20995,N_20159,N_20231);
or U20996 (N_20996,N_20224,N_20064);
xor U20997 (N_20997,N_20039,N_20455);
and U20998 (N_20998,N_20466,N_20434);
nor U20999 (N_20999,N_20422,N_20322);
nor U21000 (N_21000,N_20530,N_20635);
nand U21001 (N_21001,N_20902,N_20613);
nor U21002 (N_21002,N_20550,N_20839);
and U21003 (N_21003,N_20802,N_20698);
or U21004 (N_21004,N_20812,N_20503);
or U21005 (N_21005,N_20685,N_20844);
and U21006 (N_21006,N_20549,N_20720);
nand U21007 (N_21007,N_20790,N_20900);
nor U21008 (N_21008,N_20825,N_20568);
nor U21009 (N_21009,N_20892,N_20907);
xor U21010 (N_21010,N_20584,N_20727);
nor U21011 (N_21011,N_20578,N_20796);
nor U21012 (N_21012,N_20774,N_20716);
nand U21013 (N_21013,N_20800,N_20606);
nand U21014 (N_21014,N_20940,N_20598);
nor U21015 (N_21015,N_20577,N_20687);
xor U21016 (N_21016,N_20586,N_20982);
nand U21017 (N_21017,N_20762,N_20511);
or U21018 (N_21018,N_20832,N_20706);
nor U21019 (N_21019,N_20817,N_20527);
and U21020 (N_21020,N_20905,N_20763);
xor U21021 (N_21021,N_20792,N_20740);
nand U21022 (N_21022,N_20996,N_20827);
or U21023 (N_21023,N_20820,N_20971);
xor U21024 (N_21024,N_20741,N_20618);
or U21025 (N_21025,N_20871,N_20912);
nand U21026 (N_21026,N_20582,N_20933);
nand U21027 (N_21027,N_20724,N_20835);
nor U21028 (N_21028,N_20742,N_20688);
nand U21029 (N_21029,N_20773,N_20850);
xor U21030 (N_21030,N_20917,N_20677);
and U21031 (N_21031,N_20903,N_20631);
and U21032 (N_21032,N_20608,N_20623);
xnor U21033 (N_21033,N_20587,N_20806);
xor U21034 (N_21034,N_20506,N_20733);
nand U21035 (N_21035,N_20918,N_20634);
xnor U21036 (N_21036,N_20599,N_20620);
or U21037 (N_21037,N_20514,N_20602);
or U21038 (N_21038,N_20952,N_20922);
nor U21039 (N_21039,N_20969,N_20597);
nor U21040 (N_21040,N_20821,N_20546);
nor U21041 (N_21041,N_20668,N_20566);
and U21042 (N_21042,N_20833,N_20767);
nand U21043 (N_21043,N_20761,N_20968);
nor U21044 (N_21044,N_20998,N_20950);
xor U21045 (N_21045,N_20769,N_20883);
or U21046 (N_21046,N_20652,N_20713);
nor U21047 (N_21047,N_20845,N_20964);
and U21048 (N_21048,N_20801,N_20736);
or U21049 (N_21049,N_20849,N_20941);
xor U21050 (N_21050,N_20818,N_20703);
or U21051 (N_21051,N_20533,N_20548);
nand U21052 (N_21052,N_20787,N_20663);
and U21053 (N_21053,N_20671,N_20714);
nand U21054 (N_21054,N_20877,N_20939);
xnor U21055 (N_21055,N_20689,N_20955);
nor U21056 (N_21056,N_20643,N_20837);
and U21057 (N_21057,N_20965,N_20794);
nand U21058 (N_21058,N_20650,N_20782);
nand U21059 (N_21059,N_20680,N_20945);
xnor U21060 (N_21060,N_20557,N_20861);
nand U21061 (N_21061,N_20811,N_20691);
xor U21062 (N_21062,N_20766,N_20658);
nand U21063 (N_21063,N_20531,N_20977);
nand U21064 (N_21064,N_20534,N_20615);
xnor U21065 (N_21065,N_20633,N_20528);
xnor U21066 (N_21066,N_20522,N_20904);
nand U21067 (N_21067,N_20610,N_20656);
and U21068 (N_21068,N_20639,N_20932);
nor U21069 (N_21069,N_20651,N_20626);
nor U21070 (N_21070,N_20661,N_20931);
or U21071 (N_21071,N_20573,N_20664);
or U21072 (N_21072,N_20753,N_20757);
nand U21073 (N_21073,N_20799,N_20659);
and U21074 (N_21074,N_20579,N_20665);
and U21075 (N_21075,N_20637,N_20981);
and U21076 (N_21076,N_20589,N_20684);
xor U21077 (N_21077,N_20654,N_20819);
nor U21078 (N_21078,N_20937,N_20916);
nor U21079 (N_21079,N_20576,N_20921);
and U21080 (N_21080,N_20824,N_20695);
xnor U21081 (N_21081,N_20810,N_20959);
and U21082 (N_21082,N_20788,N_20508);
and U21083 (N_21083,N_20580,N_20644);
and U21084 (N_21084,N_20726,N_20739);
xor U21085 (N_21085,N_20700,N_20744);
or U21086 (N_21086,N_20667,N_20673);
xor U21087 (N_21087,N_20641,N_20983);
or U21088 (N_21088,N_20847,N_20961);
nand U21089 (N_21089,N_20552,N_20997);
and U21090 (N_21090,N_20660,N_20722);
nor U21091 (N_21091,N_20963,N_20554);
nand U21092 (N_21092,N_20875,N_20509);
nor U21093 (N_21093,N_20710,N_20947);
or U21094 (N_21094,N_20897,N_20666);
nand U21095 (N_21095,N_20856,N_20798);
xnor U21096 (N_21096,N_20860,N_20809);
or U21097 (N_21097,N_20542,N_20866);
nor U21098 (N_21098,N_20976,N_20814);
or U21099 (N_21099,N_20913,N_20719);
or U21100 (N_21100,N_20953,N_20693);
and U21101 (N_21101,N_20775,N_20884);
xnor U21102 (N_21102,N_20681,N_20789);
nand U21103 (N_21103,N_20797,N_20914);
and U21104 (N_21104,N_20994,N_20887);
or U21105 (N_21105,N_20778,N_20867);
and U21106 (N_21106,N_20760,N_20600);
and U21107 (N_21107,N_20901,N_20747);
nand U21108 (N_21108,N_20536,N_20885);
and U21109 (N_21109,N_20628,N_20540);
xor U21110 (N_21110,N_20516,N_20771);
nand U21111 (N_21111,N_20838,N_20951);
nand U21112 (N_21112,N_20865,N_20559);
xor U21113 (N_21113,N_20975,N_20642);
or U21114 (N_21114,N_20785,N_20957);
and U21115 (N_21115,N_20803,N_20614);
xnor U21116 (N_21116,N_20715,N_20978);
xor U21117 (N_21117,N_20864,N_20970);
xnor U21118 (N_21118,N_20855,N_20672);
or U21119 (N_21119,N_20670,N_20807);
nor U21120 (N_21120,N_20570,N_20906);
nand U21121 (N_21121,N_20991,N_20946);
or U21122 (N_21122,N_20928,N_20718);
or U21123 (N_21123,N_20513,N_20510);
nor U21124 (N_21124,N_20836,N_20874);
nor U21125 (N_21125,N_20565,N_20966);
nor U21126 (N_21126,N_20571,N_20752);
xor U21127 (N_21127,N_20842,N_20754);
nor U21128 (N_21128,N_20823,N_20558);
and U21129 (N_21129,N_20888,N_20621);
nor U21130 (N_21130,N_20869,N_20980);
nand U21131 (N_21131,N_20609,N_20686);
and U21132 (N_21132,N_20699,N_20882);
and U21133 (N_21133,N_20611,N_20772);
or U21134 (N_21134,N_20958,N_20910);
and U21135 (N_21135,N_20786,N_20784);
nor U21136 (N_21136,N_20935,N_20783);
and U21137 (N_21137,N_20507,N_20622);
and U21138 (N_21138,N_20841,N_20857);
and U21139 (N_21139,N_20944,N_20828);
and U21140 (N_21140,N_20898,N_20676);
nor U21141 (N_21141,N_20596,N_20702);
nand U21142 (N_21142,N_20630,N_20529);
or U21143 (N_21143,N_20505,N_20585);
nand U21144 (N_21144,N_20831,N_20759);
nor U21145 (N_21145,N_20541,N_20690);
nand U21146 (N_21146,N_20646,N_20524);
nand U21147 (N_21147,N_20737,N_20924);
or U21148 (N_21148,N_20822,N_20696);
and U21149 (N_21149,N_20590,N_20776);
xnor U21150 (N_21150,N_20601,N_20848);
or U21151 (N_21151,N_20567,N_20657);
nor U21152 (N_21152,N_20562,N_20834);
nor U21153 (N_21153,N_20735,N_20758);
xnor U21154 (N_21154,N_20525,N_20595);
or U21155 (N_21155,N_20972,N_20777);
nand U21156 (N_21156,N_20556,N_20632);
nand U21157 (N_21157,N_20537,N_20645);
nor U21158 (N_21158,N_20925,N_20619);
xor U21159 (N_21159,N_20605,N_20746);
nor U21160 (N_21160,N_20563,N_20880);
nor U21161 (N_21161,N_20697,N_20692);
xor U21162 (N_21162,N_20535,N_20738);
and U21163 (N_21163,N_20942,N_20526);
nand U21164 (N_21164,N_20625,N_20588);
or U21165 (N_21165,N_20551,N_20675);
or U21166 (N_21166,N_20518,N_20859);
or U21167 (N_21167,N_20593,N_20929);
nand U21168 (N_21168,N_20749,N_20872);
nand U21169 (N_21169,N_20545,N_20729);
nor U21170 (N_21170,N_20581,N_20674);
nand U21171 (N_21171,N_20755,N_20889);
and U21172 (N_21172,N_20725,N_20934);
xor U21173 (N_21173,N_20868,N_20895);
and U21174 (N_21174,N_20854,N_20879);
or U21175 (N_21175,N_20574,N_20992);
and U21176 (N_21176,N_20985,N_20682);
nand U21177 (N_21177,N_20617,N_20960);
xor U21178 (N_21178,N_20500,N_20543);
nor U21179 (N_21179,N_20701,N_20962);
or U21180 (N_21180,N_20569,N_20795);
nand U21181 (N_21181,N_20829,N_20683);
and U21182 (N_21182,N_20748,N_20560);
nor U21183 (N_21183,N_20919,N_20804);
and U21184 (N_21184,N_20911,N_20561);
and U21185 (N_21185,N_20915,N_20878);
or U21186 (N_21186,N_20908,N_20764);
xor U21187 (N_21187,N_20539,N_20979);
and U21188 (N_21188,N_20708,N_20765);
and U21189 (N_21189,N_20927,N_20876);
and U21190 (N_21190,N_20743,N_20793);
xor U21191 (N_21191,N_20949,N_20986);
and U21192 (N_21192,N_20555,N_20502);
or U21193 (N_21193,N_20731,N_20893);
xor U21194 (N_21194,N_20943,N_20732);
xor U21195 (N_21195,N_20781,N_20583);
nor U21196 (N_21196,N_20638,N_20873);
or U21197 (N_21197,N_20974,N_20948);
nor U21198 (N_21198,N_20896,N_20538);
xnor U21199 (N_21199,N_20840,N_20851);
and U21200 (N_21200,N_20648,N_20770);
xnor U21201 (N_21201,N_20909,N_20808);
or U21202 (N_21202,N_20603,N_20575);
nand U21203 (N_21203,N_20512,N_20515);
xor U21204 (N_21204,N_20993,N_20858);
nor U21205 (N_21205,N_20779,N_20519);
nand U21206 (N_21206,N_20709,N_20521);
nor U21207 (N_21207,N_20572,N_20707);
xnor U21208 (N_21208,N_20973,N_20930);
nand U21209 (N_21209,N_20830,N_20751);
and U21210 (N_21210,N_20768,N_20678);
or U21211 (N_21211,N_20846,N_20624);
and U21212 (N_21212,N_20890,N_20954);
xnor U21213 (N_21213,N_20734,N_20923);
or U21214 (N_21214,N_20501,N_20591);
xor U21215 (N_21215,N_20988,N_20629);
xor U21216 (N_21216,N_20721,N_20843);
and U21217 (N_21217,N_20564,N_20532);
nor U21218 (N_21218,N_20504,N_20612);
nand U21219 (N_21219,N_20547,N_20881);
and U21220 (N_21220,N_20640,N_20544);
and U21221 (N_21221,N_20662,N_20679);
nor U21222 (N_21222,N_20723,N_20853);
or U21223 (N_21223,N_20711,N_20712);
and U21224 (N_21224,N_20805,N_20704);
nand U21225 (N_21225,N_20627,N_20780);
nand U21226 (N_21226,N_20517,N_20938);
or U21227 (N_21227,N_20636,N_20995);
and U21228 (N_21228,N_20926,N_20594);
nand U21229 (N_21229,N_20862,N_20655);
xor U21230 (N_21230,N_20653,N_20745);
xor U21231 (N_21231,N_20863,N_20730);
nor U21232 (N_21232,N_20815,N_20891);
nand U21233 (N_21233,N_20669,N_20728);
or U21234 (N_21234,N_20870,N_20647);
and U21235 (N_21235,N_20956,N_20826);
nor U21236 (N_21236,N_20852,N_20756);
and U21237 (N_21237,N_20967,N_20592);
xnor U21238 (N_21238,N_20886,N_20604);
xnor U21239 (N_21239,N_20984,N_20750);
nor U21240 (N_21240,N_20987,N_20813);
and U21241 (N_21241,N_20894,N_20899);
or U21242 (N_21242,N_20989,N_20607);
or U21243 (N_21243,N_20649,N_20791);
or U21244 (N_21244,N_20705,N_20553);
xor U21245 (N_21245,N_20999,N_20990);
and U21246 (N_21246,N_20920,N_20936);
xnor U21247 (N_21247,N_20717,N_20520);
nand U21248 (N_21248,N_20523,N_20694);
and U21249 (N_21249,N_20816,N_20616);
nand U21250 (N_21250,N_20652,N_20922);
or U21251 (N_21251,N_20885,N_20983);
nand U21252 (N_21252,N_20793,N_20776);
and U21253 (N_21253,N_20524,N_20597);
or U21254 (N_21254,N_20960,N_20774);
and U21255 (N_21255,N_20621,N_20662);
or U21256 (N_21256,N_20626,N_20732);
nor U21257 (N_21257,N_20518,N_20534);
xnor U21258 (N_21258,N_20885,N_20725);
nor U21259 (N_21259,N_20727,N_20698);
or U21260 (N_21260,N_20989,N_20676);
nand U21261 (N_21261,N_20717,N_20858);
xor U21262 (N_21262,N_20853,N_20771);
nand U21263 (N_21263,N_20660,N_20784);
xor U21264 (N_21264,N_20891,N_20861);
nor U21265 (N_21265,N_20695,N_20745);
xor U21266 (N_21266,N_20900,N_20587);
nand U21267 (N_21267,N_20662,N_20569);
and U21268 (N_21268,N_20731,N_20641);
and U21269 (N_21269,N_20922,N_20833);
and U21270 (N_21270,N_20926,N_20837);
xor U21271 (N_21271,N_20783,N_20742);
xor U21272 (N_21272,N_20513,N_20736);
nor U21273 (N_21273,N_20784,N_20622);
and U21274 (N_21274,N_20928,N_20747);
and U21275 (N_21275,N_20878,N_20697);
xor U21276 (N_21276,N_20560,N_20760);
nor U21277 (N_21277,N_20996,N_20673);
or U21278 (N_21278,N_20938,N_20593);
nor U21279 (N_21279,N_20884,N_20967);
nor U21280 (N_21280,N_20998,N_20756);
xnor U21281 (N_21281,N_20733,N_20761);
or U21282 (N_21282,N_20818,N_20708);
nor U21283 (N_21283,N_20829,N_20846);
nor U21284 (N_21284,N_20981,N_20606);
xnor U21285 (N_21285,N_20703,N_20617);
and U21286 (N_21286,N_20946,N_20815);
nand U21287 (N_21287,N_20637,N_20825);
nor U21288 (N_21288,N_20648,N_20631);
or U21289 (N_21289,N_20945,N_20861);
nand U21290 (N_21290,N_20592,N_20516);
nor U21291 (N_21291,N_20817,N_20847);
and U21292 (N_21292,N_20767,N_20939);
nand U21293 (N_21293,N_20909,N_20628);
or U21294 (N_21294,N_20867,N_20558);
and U21295 (N_21295,N_20546,N_20993);
xnor U21296 (N_21296,N_20502,N_20764);
nor U21297 (N_21297,N_20773,N_20662);
xnor U21298 (N_21298,N_20616,N_20946);
xnor U21299 (N_21299,N_20954,N_20892);
or U21300 (N_21300,N_20724,N_20841);
nand U21301 (N_21301,N_20504,N_20643);
xnor U21302 (N_21302,N_20811,N_20696);
and U21303 (N_21303,N_20830,N_20505);
and U21304 (N_21304,N_20612,N_20702);
nand U21305 (N_21305,N_20717,N_20875);
nand U21306 (N_21306,N_20935,N_20703);
and U21307 (N_21307,N_20965,N_20838);
and U21308 (N_21308,N_20939,N_20711);
or U21309 (N_21309,N_20540,N_20583);
nand U21310 (N_21310,N_20935,N_20714);
nor U21311 (N_21311,N_20807,N_20623);
nor U21312 (N_21312,N_20761,N_20956);
nor U21313 (N_21313,N_20879,N_20621);
nand U21314 (N_21314,N_20715,N_20614);
nor U21315 (N_21315,N_20943,N_20993);
xor U21316 (N_21316,N_20671,N_20675);
xnor U21317 (N_21317,N_20715,N_20700);
or U21318 (N_21318,N_20621,N_20893);
nor U21319 (N_21319,N_20548,N_20595);
and U21320 (N_21320,N_20587,N_20887);
nand U21321 (N_21321,N_20718,N_20548);
or U21322 (N_21322,N_20942,N_20881);
xor U21323 (N_21323,N_20763,N_20715);
nand U21324 (N_21324,N_20884,N_20989);
and U21325 (N_21325,N_20611,N_20553);
nor U21326 (N_21326,N_20867,N_20818);
nor U21327 (N_21327,N_20681,N_20923);
and U21328 (N_21328,N_20975,N_20713);
nand U21329 (N_21329,N_20925,N_20962);
or U21330 (N_21330,N_20696,N_20843);
xor U21331 (N_21331,N_20913,N_20958);
nor U21332 (N_21332,N_20638,N_20623);
xnor U21333 (N_21333,N_20956,N_20633);
xor U21334 (N_21334,N_20914,N_20677);
or U21335 (N_21335,N_20947,N_20758);
nand U21336 (N_21336,N_20995,N_20625);
nor U21337 (N_21337,N_20755,N_20912);
and U21338 (N_21338,N_20648,N_20536);
xor U21339 (N_21339,N_20756,N_20655);
or U21340 (N_21340,N_20697,N_20814);
nor U21341 (N_21341,N_20764,N_20539);
and U21342 (N_21342,N_20656,N_20646);
nor U21343 (N_21343,N_20953,N_20508);
xor U21344 (N_21344,N_20956,N_20885);
nor U21345 (N_21345,N_20541,N_20877);
nor U21346 (N_21346,N_20650,N_20918);
xnor U21347 (N_21347,N_20627,N_20611);
or U21348 (N_21348,N_20815,N_20669);
and U21349 (N_21349,N_20880,N_20966);
and U21350 (N_21350,N_20793,N_20806);
nor U21351 (N_21351,N_20555,N_20981);
and U21352 (N_21352,N_20737,N_20624);
or U21353 (N_21353,N_20625,N_20716);
and U21354 (N_21354,N_20504,N_20854);
or U21355 (N_21355,N_20819,N_20708);
xor U21356 (N_21356,N_20603,N_20725);
nand U21357 (N_21357,N_20661,N_20715);
or U21358 (N_21358,N_20601,N_20851);
nor U21359 (N_21359,N_20747,N_20706);
xor U21360 (N_21360,N_20772,N_20894);
xnor U21361 (N_21361,N_20530,N_20890);
nand U21362 (N_21362,N_20935,N_20741);
nor U21363 (N_21363,N_20638,N_20790);
nor U21364 (N_21364,N_20748,N_20645);
and U21365 (N_21365,N_20851,N_20644);
or U21366 (N_21366,N_20851,N_20579);
xnor U21367 (N_21367,N_20924,N_20895);
nor U21368 (N_21368,N_20552,N_20578);
xnor U21369 (N_21369,N_20822,N_20963);
xor U21370 (N_21370,N_20715,N_20638);
and U21371 (N_21371,N_20861,N_20635);
and U21372 (N_21372,N_20767,N_20918);
or U21373 (N_21373,N_20735,N_20759);
nand U21374 (N_21374,N_20719,N_20503);
and U21375 (N_21375,N_20637,N_20878);
nand U21376 (N_21376,N_20841,N_20888);
or U21377 (N_21377,N_20861,N_20881);
nand U21378 (N_21378,N_20927,N_20847);
and U21379 (N_21379,N_20683,N_20947);
nor U21380 (N_21380,N_20997,N_20929);
nor U21381 (N_21381,N_20578,N_20586);
nand U21382 (N_21382,N_20880,N_20784);
nand U21383 (N_21383,N_20745,N_20911);
nand U21384 (N_21384,N_20913,N_20998);
or U21385 (N_21385,N_20680,N_20875);
or U21386 (N_21386,N_20985,N_20930);
nor U21387 (N_21387,N_20548,N_20714);
xor U21388 (N_21388,N_20967,N_20851);
and U21389 (N_21389,N_20924,N_20557);
or U21390 (N_21390,N_20528,N_20554);
and U21391 (N_21391,N_20972,N_20884);
or U21392 (N_21392,N_20689,N_20663);
nand U21393 (N_21393,N_20506,N_20650);
and U21394 (N_21394,N_20503,N_20857);
nand U21395 (N_21395,N_20745,N_20690);
nand U21396 (N_21396,N_20993,N_20509);
or U21397 (N_21397,N_20946,N_20842);
nand U21398 (N_21398,N_20958,N_20578);
and U21399 (N_21399,N_20933,N_20886);
nand U21400 (N_21400,N_20804,N_20970);
xnor U21401 (N_21401,N_20943,N_20973);
nor U21402 (N_21402,N_20587,N_20879);
xor U21403 (N_21403,N_20812,N_20888);
nand U21404 (N_21404,N_20785,N_20844);
and U21405 (N_21405,N_20607,N_20804);
nand U21406 (N_21406,N_20963,N_20775);
xnor U21407 (N_21407,N_20527,N_20933);
nor U21408 (N_21408,N_20626,N_20937);
nand U21409 (N_21409,N_20889,N_20986);
or U21410 (N_21410,N_20745,N_20995);
nand U21411 (N_21411,N_20582,N_20693);
xnor U21412 (N_21412,N_20821,N_20792);
and U21413 (N_21413,N_20563,N_20908);
or U21414 (N_21414,N_20952,N_20985);
or U21415 (N_21415,N_20581,N_20736);
nor U21416 (N_21416,N_20829,N_20543);
nand U21417 (N_21417,N_20817,N_20660);
xnor U21418 (N_21418,N_20623,N_20911);
and U21419 (N_21419,N_20596,N_20914);
or U21420 (N_21420,N_20655,N_20943);
and U21421 (N_21421,N_20854,N_20776);
xor U21422 (N_21422,N_20935,N_20596);
and U21423 (N_21423,N_20621,N_20613);
or U21424 (N_21424,N_20976,N_20764);
and U21425 (N_21425,N_20576,N_20825);
nand U21426 (N_21426,N_20699,N_20556);
and U21427 (N_21427,N_20807,N_20987);
nor U21428 (N_21428,N_20888,N_20677);
or U21429 (N_21429,N_20914,N_20840);
and U21430 (N_21430,N_20578,N_20809);
xor U21431 (N_21431,N_20682,N_20923);
and U21432 (N_21432,N_20654,N_20865);
nand U21433 (N_21433,N_20816,N_20951);
nor U21434 (N_21434,N_20636,N_20739);
or U21435 (N_21435,N_20962,N_20658);
or U21436 (N_21436,N_20804,N_20615);
and U21437 (N_21437,N_20602,N_20511);
or U21438 (N_21438,N_20969,N_20847);
nor U21439 (N_21439,N_20678,N_20873);
or U21440 (N_21440,N_20815,N_20523);
or U21441 (N_21441,N_20947,N_20672);
nand U21442 (N_21442,N_20822,N_20695);
xor U21443 (N_21443,N_20868,N_20658);
nor U21444 (N_21444,N_20891,N_20821);
or U21445 (N_21445,N_20928,N_20669);
nor U21446 (N_21446,N_20597,N_20928);
or U21447 (N_21447,N_20867,N_20503);
nor U21448 (N_21448,N_20616,N_20688);
nor U21449 (N_21449,N_20749,N_20682);
or U21450 (N_21450,N_20910,N_20733);
nor U21451 (N_21451,N_20516,N_20726);
xnor U21452 (N_21452,N_20657,N_20798);
nand U21453 (N_21453,N_20512,N_20852);
xor U21454 (N_21454,N_20605,N_20525);
xnor U21455 (N_21455,N_20545,N_20987);
nor U21456 (N_21456,N_20733,N_20991);
or U21457 (N_21457,N_20740,N_20940);
nand U21458 (N_21458,N_20869,N_20935);
nor U21459 (N_21459,N_20973,N_20794);
nor U21460 (N_21460,N_20865,N_20897);
nor U21461 (N_21461,N_20794,N_20960);
nor U21462 (N_21462,N_20814,N_20960);
nand U21463 (N_21463,N_20557,N_20563);
and U21464 (N_21464,N_20744,N_20808);
or U21465 (N_21465,N_20782,N_20621);
and U21466 (N_21466,N_20959,N_20612);
nor U21467 (N_21467,N_20780,N_20935);
and U21468 (N_21468,N_20842,N_20627);
and U21469 (N_21469,N_20842,N_20707);
nand U21470 (N_21470,N_20500,N_20744);
or U21471 (N_21471,N_20620,N_20764);
nand U21472 (N_21472,N_20895,N_20548);
nand U21473 (N_21473,N_20537,N_20658);
and U21474 (N_21474,N_20815,N_20569);
nor U21475 (N_21475,N_20953,N_20983);
xor U21476 (N_21476,N_20806,N_20558);
nand U21477 (N_21477,N_20862,N_20886);
nor U21478 (N_21478,N_20584,N_20869);
or U21479 (N_21479,N_20926,N_20854);
nor U21480 (N_21480,N_20867,N_20855);
or U21481 (N_21481,N_20806,N_20789);
and U21482 (N_21482,N_20622,N_20872);
nor U21483 (N_21483,N_20696,N_20557);
or U21484 (N_21484,N_20580,N_20729);
nand U21485 (N_21485,N_20560,N_20997);
nor U21486 (N_21486,N_20602,N_20526);
xor U21487 (N_21487,N_20856,N_20610);
nor U21488 (N_21488,N_20989,N_20977);
nor U21489 (N_21489,N_20900,N_20558);
xnor U21490 (N_21490,N_20770,N_20843);
or U21491 (N_21491,N_20701,N_20583);
nand U21492 (N_21492,N_20540,N_20809);
xor U21493 (N_21493,N_20943,N_20790);
or U21494 (N_21494,N_20990,N_20629);
nor U21495 (N_21495,N_20646,N_20573);
or U21496 (N_21496,N_20505,N_20989);
nand U21497 (N_21497,N_20852,N_20763);
and U21498 (N_21498,N_20953,N_20598);
nand U21499 (N_21499,N_20634,N_20529);
nand U21500 (N_21500,N_21402,N_21493);
nor U21501 (N_21501,N_21334,N_21478);
xor U21502 (N_21502,N_21224,N_21248);
nor U21503 (N_21503,N_21260,N_21379);
nor U21504 (N_21504,N_21044,N_21229);
nor U21505 (N_21505,N_21182,N_21002);
nand U21506 (N_21506,N_21169,N_21181);
or U21507 (N_21507,N_21395,N_21098);
nand U21508 (N_21508,N_21313,N_21436);
and U21509 (N_21509,N_21107,N_21339);
nor U21510 (N_21510,N_21490,N_21352);
xnor U21511 (N_21511,N_21294,N_21285);
xor U21512 (N_21512,N_21400,N_21265);
nor U21513 (N_21513,N_21037,N_21468);
or U21514 (N_21514,N_21286,N_21299);
or U21515 (N_21515,N_21159,N_21177);
nor U21516 (N_21516,N_21201,N_21045);
and U21517 (N_21517,N_21350,N_21043);
and U21518 (N_21518,N_21443,N_21122);
nor U21519 (N_21519,N_21251,N_21087);
and U21520 (N_21520,N_21430,N_21276);
or U21521 (N_21521,N_21047,N_21228);
xor U21522 (N_21522,N_21115,N_21289);
xnor U21523 (N_21523,N_21155,N_21396);
nand U21524 (N_21524,N_21462,N_21358);
nor U21525 (N_21525,N_21267,N_21000);
xnor U21526 (N_21526,N_21009,N_21481);
or U21527 (N_21527,N_21231,N_21453);
nand U21528 (N_21528,N_21070,N_21382);
or U21529 (N_21529,N_21372,N_21046);
and U21530 (N_21530,N_21357,N_21280);
xnor U21531 (N_21531,N_21381,N_21342);
xor U21532 (N_21532,N_21494,N_21326);
or U21533 (N_21533,N_21405,N_21208);
xor U21534 (N_21534,N_21362,N_21364);
xor U21535 (N_21535,N_21300,N_21034);
or U21536 (N_21536,N_21190,N_21001);
nor U21537 (N_21537,N_21214,N_21234);
or U21538 (N_21538,N_21380,N_21288);
and U21539 (N_21539,N_21345,N_21124);
xor U21540 (N_21540,N_21466,N_21007);
nor U21541 (N_21541,N_21471,N_21066);
nor U21542 (N_21542,N_21212,N_21096);
xor U21543 (N_21543,N_21186,N_21366);
or U21544 (N_21544,N_21135,N_21061);
and U21545 (N_21545,N_21447,N_21119);
and U21546 (N_21546,N_21144,N_21051);
xor U21547 (N_21547,N_21189,N_21220);
xnor U21548 (N_21548,N_21164,N_21238);
xor U21549 (N_21549,N_21239,N_21129);
nor U21550 (N_21550,N_21069,N_21469);
nand U21551 (N_21551,N_21480,N_21010);
nand U21552 (N_21552,N_21290,N_21021);
nor U21553 (N_21553,N_21012,N_21036);
or U21554 (N_21554,N_21424,N_21148);
nand U21555 (N_21555,N_21143,N_21329);
xor U21556 (N_21556,N_21355,N_21261);
nand U21557 (N_21557,N_21196,N_21470);
xor U21558 (N_21558,N_21211,N_21052);
xnor U21559 (N_21559,N_21183,N_21132);
xnor U21560 (N_21560,N_21247,N_21095);
or U21561 (N_21561,N_21316,N_21445);
nand U21562 (N_21562,N_21412,N_21141);
nor U21563 (N_21563,N_21496,N_21423);
and U21564 (N_21564,N_21409,N_21093);
and U21565 (N_21565,N_21333,N_21439);
and U21566 (N_21566,N_21078,N_21308);
or U21567 (N_21567,N_21246,N_21040);
xor U21568 (N_21568,N_21179,N_21109);
nor U21569 (N_21569,N_21207,N_21136);
and U21570 (N_21570,N_21374,N_21121);
xor U21571 (N_21571,N_21283,N_21270);
nor U21572 (N_21572,N_21198,N_21112);
and U21573 (N_21573,N_21337,N_21172);
xor U21574 (N_21574,N_21204,N_21076);
xnor U21575 (N_21575,N_21346,N_21020);
xnor U21576 (N_21576,N_21406,N_21079);
or U21577 (N_21577,N_21319,N_21278);
nand U21578 (N_21578,N_21206,N_21476);
xor U21579 (N_21579,N_21483,N_21097);
nor U21580 (N_21580,N_21279,N_21178);
xor U21581 (N_21581,N_21318,N_21033);
nor U21582 (N_21582,N_21042,N_21477);
nand U21583 (N_21583,N_21486,N_21029);
or U21584 (N_21584,N_21213,N_21099);
nor U21585 (N_21585,N_21360,N_21056);
nand U21586 (N_21586,N_21041,N_21418);
nand U21587 (N_21587,N_21084,N_21072);
and U21588 (N_21588,N_21101,N_21293);
xor U21589 (N_21589,N_21442,N_21343);
nand U21590 (N_21590,N_21106,N_21068);
nand U21591 (N_21591,N_21088,N_21230);
or U21592 (N_21592,N_21272,N_21348);
nor U21593 (N_21593,N_21451,N_21365);
nand U21594 (N_21594,N_21315,N_21401);
nand U21595 (N_21595,N_21243,N_21487);
or U21596 (N_21596,N_21254,N_21473);
nand U21597 (N_21597,N_21377,N_21398);
nand U21598 (N_21598,N_21393,N_21140);
nor U21599 (N_21599,N_21387,N_21197);
xnor U21600 (N_21600,N_21306,N_21336);
or U21601 (N_21601,N_21128,N_21018);
or U21602 (N_21602,N_21110,N_21347);
or U21603 (N_21603,N_21323,N_21085);
nor U21604 (N_21604,N_21116,N_21497);
or U21605 (N_21605,N_21351,N_21369);
nor U21606 (N_21606,N_21062,N_21103);
nand U21607 (N_21607,N_21199,N_21367);
xor U21608 (N_21608,N_21475,N_21435);
or U21609 (N_21609,N_21269,N_21499);
nor U21610 (N_21610,N_21174,N_21138);
and U21611 (N_21611,N_21147,N_21472);
or U21612 (N_21612,N_21322,N_21263);
and U21613 (N_21613,N_21287,N_21422);
xor U21614 (N_21614,N_21053,N_21038);
and U21615 (N_21615,N_21474,N_21091);
and U21616 (N_21616,N_21222,N_21495);
nand U21617 (N_21617,N_21026,N_21166);
nand U21618 (N_21618,N_21489,N_21421);
and U21619 (N_21619,N_21003,N_21118);
or U21620 (N_21620,N_21014,N_21125);
nand U21621 (N_21621,N_21117,N_21426);
and U21622 (N_21622,N_21253,N_21139);
nor U21623 (N_21623,N_21258,N_21344);
xnor U21624 (N_21624,N_21416,N_21448);
nor U21625 (N_21625,N_21295,N_21071);
and U21626 (N_21626,N_21185,N_21356);
and U21627 (N_21627,N_21301,N_21375);
or U21628 (N_21628,N_21063,N_21249);
nor U21629 (N_21629,N_21321,N_21149);
and U21630 (N_21630,N_21310,N_21142);
nor U21631 (N_21631,N_21349,N_21391);
nand U21632 (N_21632,N_21011,N_21039);
nor U21633 (N_21633,N_21060,N_21492);
or U21634 (N_21634,N_21081,N_21153);
or U21635 (N_21635,N_21394,N_21219);
nand U21636 (N_21636,N_21378,N_21429);
or U21637 (N_21637,N_21274,N_21331);
xnor U21638 (N_21638,N_21126,N_21386);
and U21639 (N_21639,N_21027,N_21160);
and U21640 (N_21640,N_21077,N_21428);
nand U21641 (N_21641,N_21111,N_21432);
xnor U21642 (N_21642,N_21022,N_21216);
nor U21643 (N_21643,N_21427,N_21089);
nor U21644 (N_21644,N_21498,N_21371);
nor U21645 (N_21645,N_21232,N_21217);
and U21646 (N_21646,N_21059,N_21328);
nor U21647 (N_21647,N_21291,N_21008);
nand U21648 (N_21648,N_21171,N_21242);
nor U21649 (N_21649,N_21438,N_21457);
nor U21650 (N_21650,N_21067,N_21168);
nand U21651 (N_21651,N_21028,N_21163);
nor U21652 (N_21652,N_21414,N_21210);
xnor U21653 (N_21653,N_21048,N_21105);
or U21654 (N_21654,N_21170,N_21373);
or U21655 (N_21655,N_21410,N_21146);
nor U21656 (N_21656,N_21444,N_21407);
and U21657 (N_21657,N_21311,N_21463);
nand U21658 (N_21658,N_21131,N_21479);
xnor U21659 (N_21659,N_21133,N_21244);
xor U21660 (N_21660,N_21054,N_21092);
nor U21661 (N_21661,N_21123,N_21455);
nand U21662 (N_21662,N_21102,N_21433);
xor U21663 (N_21663,N_21031,N_21388);
nand U21664 (N_21664,N_21454,N_21297);
and U21665 (N_21665,N_21257,N_21441);
or U21666 (N_21666,N_21165,N_21275);
nand U21667 (N_21667,N_21024,N_21403);
xnor U21668 (N_21668,N_21237,N_21006);
xnor U21669 (N_21669,N_21245,N_21145);
nor U21670 (N_21670,N_21184,N_21465);
or U21671 (N_21671,N_21284,N_21200);
xor U21672 (N_21672,N_21137,N_21361);
xor U21673 (N_21673,N_21055,N_21440);
nand U21674 (N_21674,N_21425,N_21157);
and U21675 (N_21675,N_21241,N_21385);
nand U21676 (N_21676,N_21233,N_21307);
and U21677 (N_21677,N_21151,N_21359);
xor U21678 (N_21678,N_21057,N_21017);
nand U21679 (N_21679,N_21113,N_21223);
and U21680 (N_21680,N_21235,N_21456);
and U21681 (N_21681,N_21491,N_21152);
and U21682 (N_21682,N_21074,N_21446);
nand U21683 (N_21683,N_21005,N_21209);
nor U21684 (N_21684,N_21205,N_21281);
and U21685 (N_21685,N_21392,N_21314);
xor U21686 (N_21686,N_21127,N_21282);
nor U21687 (N_21687,N_21187,N_21277);
nor U21688 (N_21688,N_21353,N_21094);
nand U21689 (N_21689,N_21298,N_21332);
xor U21690 (N_21690,N_21108,N_21255);
or U21691 (N_21691,N_21134,N_21156);
and U21692 (N_21692,N_21459,N_21354);
nand U21693 (N_21693,N_21023,N_21188);
xor U21694 (N_21694,N_21384,N_21218);
and U21695 (N_21695,N_21399,N_21050);
xor U21696 (N_21696,N_21450,N_21065);
xnor U21697 (N_21697,N_21192,N_21317);
and U21698 (N_21698,N_21240,N_21415);
xnor U21699 (N_21699,N_21340,N_21130);
or U21700 (N_21700,N_21058,N_21485);
or U21701 (N_21701,N_21266,N_21082);
nand U21702 (N_21702,N_21452,N_21049);
and U21703 (N_21703,N_21458,N_21324);
nor U21704 (N_21704,N_21335,N_21161);
and U21705 (N_21705,N_21173,N_21404);
or U21706 (N_21706,N_21086,N_21175);
or U21707 (N_21707,N_21488,N_21252);
nor U21708 (N_21708,N_21083,N_21449);
or U21709 (N_21709,N_21104,N_21389);
or U21710 (N_21710,N_21154,N_21193);
and U21711 (N_21711,N_21019,N_21312);
or U21712 (N_21712,N_21180,N_21413);
or U21713 (N_21713,N_21194,N_21268);
and U21714 (N_21714,N_21075,N_21195);
nor U21715 (N_21715,N_21484,N_21273);
xor U21716 (N_21716,N_21202,N_21460);
nand U21717 (N_21717,N_21417,N_21176);
and U21718 (N_21718,N_21408,N_21397);
nand U21719 (N_21719,N_21383,N_21271);
or U21720 (N_21720,N_21013,N_21330);
or U21721 (N_21721,N_21437,N_21150);
and U21722 (N_21722,N_21461,N_21376);
and U21723 (N_21723,N_21225,N_21305);
nor U21724 (N_21724,N_21368,N_21226);
xor U21725 (N_21725,N_21030,N_21025);
nor U21726 (N_21726,N_21292,N_21370);
nand U21727 (N_21727,N_21325,N_21302);
nor U21728 (N_21728,N_21073,N_21304);
nor U21729 (N_21729,N_21327,N_21221);
nand U21730 (N_21730,N_21309,N_21215);
nor U21731 (N_21731,N_21250,N_21035);
xor U21732 (N_21732,N_21259,N_21004);
and U21733 (N_21733,N_21341,N_21016);
and U21734 (N_21734,N_21167,N_21467);
xnor U21735 (N_21735,N_21032,N_21064);
nor U21736 (N_21736,N_21264,N_21482);
nand U21737 (N_21737,N_21100,N_21363);
and U21738 (N_21738,N_21262,N_21419);
xnor U21739 (N_21739,N_21256,N_21411);
nor U21740 (N_21740,N_21338,N_21236);
and U21741 (N_21741,N_21080,N_21191);
nand U21742 (N_21742,N_21158,N_21303);
and U21743 (N_21743,N_21434,N_21320);
and U21744 (N_21744,N_21390,N_21464);
nor U21745 (N_21745,N_21114,N_21420);
nand U21746 (N_21746,N_21015,N_21162);
and U21747 (N_21747,N_21431,N_21203);
and U21748 (N_21748,N_21090,N_21120);
and U21749 (N_21749,N_21227,N_21296);
and U21750 (N_21750,N_21252,N_21431);
nand U21751 (N_21751,N_21469,N_21327);
xnor U21752 (N_21752,N_21409,N_21118);
nand U21753 (N_21753,N_21224,N_21119);
or U21754 (N_21754,N_21441,N_21401);
and U21755 (N_21755,N_21431,N_21273);
and U21756 (N_21756,N_21177,N_21036);
xor U21757 (N_21757,N_21239,N_21080);
nand U21758 (N_21758,N_21476,N_21345);
or U21759 (N_21759,N_21090,N_21248);
nand U21760 (N_21760,N_21025,N_21472);
xor U21761 (N_21761,N_21196,N_21323);
or U21762 (N_21762,N_21201,N_21008);
nand U21763 (N_21763,N_21292,N_21447);
nand U21764 (N_21764,N_21451,N_21216);
nand U21765 (N_21765,N_21262,N_21086);
nor U21766 (N_21766,N_21343,N_21438);
and U21767 (N_21767,N_21108,N_21190);
xor U21768 (N_21768,N_21142,N_21053);
nand U21769 (N_21769,N_21423,N_21209);
and U21770 (N_21770,N_21171,N_21177);
or U21771 (N_21771,N_21381,N_21327);
xnor U21772 (N_21772,N_21221,N_21027);
nor U21773 (N_21773,N_21249,N_21011);
xnor U21774 (N_21774,N_21393,N_21449);
nand U21775 (N_21775,N_21013,N_21450);
and U21776 (N_21776,N_21154,N_21375);
nor U21777 (N_21777,N_21232,N_21137);
nor U21778 (N_21778,N_21149,N_21052);
or U21779 (N_21779,N_21258,N_21291);
or U21780 (N_21780,N_21450,N_21347);
nand U21781 (N_21781,N_21212,N_21302);
or U21782 (N_21782,N_21204,N_21110);
nor U21783 (N_21783,N_21028,N_21365);
nor U21784 (N_21784,N_21458,N_21295);
xnor U21785 (N_21785,N_21374,N_21204);
and U21786 (N_21786,N_21172,N_21346);
or U21787 (N_21787,N_21383,N_21381);
or U21788 (N_21788,N_21093,N_21132);
xor U21789 (N_21789,N_21183,N_21121);
or U21790 (N_21790,N_21475,N_21073);
xnor U21791 (N_21791,N_21422,N_21470);
nand U21792 (N_21792,N_21454,N_21289);
and U21793 (N_21793,N_21087,N_21222);
and U21794 (N_21794,N_21155,N_21030);
nor U21795 (N_21795,N_21479,N_21219);
and U21796 (N_21796,N_21021,N_21047);
and U21797 (N_21797,N_21380,N_21395);
or U21798 (N_21798,N_21115,N_21459);
nand U21799 (N_21799,N_21070,N_21118);
and U21800 (N_21800,N_21409,N_21316);
nand U21801 (N_21801,N_21304,N_21121);
and U21802 (N_21802,N_21326,N_21437);
or U21803 (N_21803,N_21288,N_21232);
or U21804 (N_21804,N_21160,N_21111);
nor U21805 (N_21805,N_21193,N_21358);
nand U21806 (N_21806,N_21059,N_21389);
or U21807 (N_21807,N_21430,N_21306);
nand U21808 (N_21808,N_21390,N_21391);
and U21809 (N_21809,N_21052,N_21294);
nand U21810 (N_21810,N_21199,N_21090);
nor U21811 (N_21811,N_21404,N_21080);
or U21812 (N_21812,N_21352,N_21333);
or U21813 (N_21813,N_21147,N_21461);
and U21814 (N_21814,N_21443,N_21034);
nand U21815 (N_21815,N_21200,N_21410);
nor U21816 (N_21816,N_21374,N_21164);
xnor U21817 (N_21817,N_21274,N_21150);
and U21818 (N_21818,N_21344,N_21448);
and U21819 (N_21819,N_21031,N_21333);
nor U21820 (N_21820,N_21402,N_21379);
nor U21821 (N_21821,N_21314,N_21089);
nor U21822 (N_21822,N_21418,N_21119);
or U21823 (N_21823,N_21326,N_21146);
nor U21824 (N_21824,N_21054,N_21375);
or U21825 (N_21825,N_21128,N_21016);
xnor U21826 (N_21826,N_21109,N_21018);
and U21827 (N_21827,N_21296,N_21065);
and U21828 (N_21828,N_21307,N_21121);
or U21829 (N_21829,N_21018,N_21313);
and U21830 (N_21830,N_21434,N_21154);
nand U21831 (N_21831,N_21347,N_21454);
xor U21832 (N_21832,N_21468,N_21379);
or U21833 (N_21833,N_21137,N_21061);
and U21834 (N_21834,N_21231,N_21351);
nand U21835 (N_21835,N_21315,N_21233);
xor U21836 (N_21836,N_21282,N_21213);
nand U21837 (N_21837,N_21125,N_21213);
and U21838 (N_21838,N_21018,N_21335);
and U21839 (N_21839,N_21108,N_21336);
nand U21840 (N_21840,N_21253,N_21026);
xnor U21841 (N_21841,N_21311,N_21385);
xor U21842 (N_21842,N_21340,N_21006);
nand U21843 (N_21843,N_21248,N_21189);
xor U21844 (N_21844,N_21193,N_21105);
and U21845 (N_21845,N_21199,N_21052);
and U21846 (N_21846,N_21339,N_21099);
nand U21847 (N_21847,N_21255,N_21310);
or U21848 (N_21848,N_21396,N_21235);
nand U21849 (N_21849,N_21030,N_21188);
nand U21850 (N_21850,N_21095,N_21394);
and U21851 (N_21851,N_21230,N_21221);
and U21852 (N_21852,N_21441,N_21074);
nor U21853 (N_21853,N_21130,N_21071);
xor U21854 (N_21854,N_21101,N_21094);
nand U21855 (N_21855,N_21334,N_21108);
nor U21856 (N_21856,N_21330,N_21158);
xnor U21857 (N_21857,N_21339,N_21376);
or U21858 (N_21858,N_21465,N_21349);
xor U21859 (N_21859,N_21127,N_21374);
nand U21860 (N_21860,N_21363,N_21455);
nor U21861 (N_21861,N_21002,N_21439);
xnor U21862 (N_21862,N_21451,N_21271);
nor U21863 (N_21863,N_21313,N_21035);
or U21864 (N_21864,N_21408,N_21019);
or U21865 (N_21865,N_21095,N_21435);
nand U21866 (N_21866,N_21355,N_21071);
or U21867 (N_21867,N_21035,N_21339);
and U21868 (N_21868,N_21491,N_21499);
or U21869 (N_21869,N_21260,N_21440);
or U21870 (N_21870,N_21105,N_21016);
nor U21871 (N_21871,N_21231,N_21321);
and U21872 (N_21872,N_21202,N_21138);
nor U21873 (N_21873,N_21194,N_21202);
nand U21874 (N_21874,N_21412,N_21434);
xnor U21875 (N_21875,N_21287,N_21070);
nor U21876 (N_21876,N_21189,N_21212);
xnor U21877 (N_21877,N_21133,N_21220);
xnor U21878 (N_21878,N_21093,N_21320);
nor U21879 (N_21879,N_21254,N_21464);
nand U21880 (N_21880,N_21174,N_21366);
xnor U21881 (N_21881,N_21051,N_21137);
or U21882 (N_21882,N_21035,N_21410);
xnor U21883 (N_21883,N_21087,N_21080);
or U21884 (N_21884,N_21322,N_21381);
nor U21885 (N_21885,N_21493,N_21166);
nand U21886 (N_21886,N_21338,N_21212);
nor U21887 (N_21887,N_21186,N_21357);
nor U21888 (N_21888,N_21447,N_21269);
or U21889 (N_21889,N_21395,N_21471);
xnor U21890 (N_21890,N_21478,N_21482);
xnor U21891 (N_21891,N_21220,N_21419);
xor U21892 (N_21892,N_21063,N_21257);
nand U21893 (N_21893,N_21167,N_21450);
and U21894 (N_21894,N_21438,N_21252);
nand U21895 (N_21895,N_21194,N_21409);
nand U21896 (N_21896,N_21025,N_21039);
nand U21897 (N_21897,N_21464,N_21322);
nor U21898 (N_21898,N_21465,N_21162);
or U21899 (N_21899,N_21481,N_21334);
nand U21900 (N_21900,N_21302,N_21101);
or U21901 (N_21901,N_21453,N_21161);
or U21902 (N_21902,N_21471,N_21332);
and U21903 (N_21903,N_21434,N_21391);
nor U21904 (N_21904,N_21103,N_21035);
and U21905 (N_21905,N_21056,N_21209);
and U21906 (N_21906,N_21033,N_21217);
or U21907 (N_21907,N_21182,N_21383);
or U21908 (N_21908,N_21243,N_21401);
nand U21909 (N_21909,N_21335,N_21423);
nor U21910 (N_21910,N_21212,N_21129);
nand U21911 (N_21911,N_21339,N_21121);
or U21912 (N_21912,N_21027,N_21385);
and U21913 (N_21913,N_21392,N_21457);
xnor U21914 (N_21914,N_21377,N_21137);
and U21915 (N_21915,N_21280,N_21149);
and U21916 (N_21916,N_21295,N_21052);
and U21917 (N_21917,N_21152,N_21279);
nand U21918 (N_21918,N_21112,N_21038);
nor U21919 (N_21919,N_21055,N_21050);
and U21920 (N_21920,N_21189,N_21079);
nor U21921 (N_21921,N_21442,N_21041);
or U21922 (N_21922,N_21167,N_21006);
nor U21923 (N_21923,N_21357,N_21079);
or U21924 (N_21924,N_21467,N_21185);
and U21925 (N_21925,N_21121,N_21155);
xor U21926 (N_21926,N_21143,N_21252);
nor U21927 (N_21927,N_21036,N_21077);
nor U21928 (N_21928,N_21450,N_21318);
nand U21929 (N_21929,N_21261,N_21469);
and U21930 (N_21930,N_21128,N_21436);
nand U21931 (N_21931,N_21226,N_21439);
xnor U21932 (N_21932,N_21498,N_21409);
or U21933 (N_21933,N_21361,N_21132);
xor U21934 (N_21934,N_21471,N_21211);
nand U21935 (N_21935,N_21281,N_21141);
and U21936 (N_21936,N_21158,N_21370);
or U21937 (N_21937,N_21152,N_21227);
xor U21938 (N_21938,N_21131,N_21439);
xor U21939 (N_21939,N_21123,N_21478);
and U21940 (N_21940,N_21497,N_21128);
nand U21941 (N_21941,N_21077,N_21403);
and U21942 (N_21942,N_21438,N_21317);
nor U21943 (N_21943,N_21101,N_21193);
and U21944 (N_21944,N_21229,N_21047);
nand U21945 (N_21945,N_21282,N_21057);
xor U21946 (N_21946,N_21290,N_21270);
and U21947 (N_21947,N_21288,N_21075);
xor U21948 (N_21948,N_21147,N_21315);
or U21949 (N_21949,N_21230,N_21360);
nor U21950 (N_21950,N_21064,N_21410);
nor U21951 (N_21951,N_21405,N_21059);
nand U21952 (N_21952,N_21100,N_21293);
nand U21953 (N_21953,N_21037,N_21108);
xnor U21954 (N_21954,N_21048,N_21081);
nor U21955 (N_21955,N_21169,N_21221);
or U21956 (N_21956,N_21314,N_21269);
and U21957 (N_21957,N_21318,N_21087);
xnor U21958 (N_21958,N_21301,N_21383);
nand U21959 (N_21959,N_21118,N_21460);
or U21960 (N_21960,N_21427,N_21236);
and U21961 (N_21961,N_21327,N_21273);
and U21962 (N_21962,N_21400,N_21192);
or U21963 (N_21963,N_21349,N_21419);
nand U21964 (N_21964,N_21479,N_21134);
nor U21965 (N_21965,N_21185,N_21212);
nor U21966 (N_21966,N_21317,N_21231);
nand U21967 (N_21967,N_21241,N_21027);
or U21968 (N_21968,N_21488,N_21069);
or U21969 (N_21969,N_21302,N_21383);
nand U21970 (N_21970,N_21313,N_21334);
or U21971 (N_21971,N_21280,N_21199);
nand U21972 (N_21972,N_21214,N_21040);
and U21973 (N_21973,N_21125,N_21387);
xnor U21974 (N_21974,N_21067,N_21381);
nand U21975 (N_21975,N_21283,N_21441);
nor U21976 (N_21976,N_21034,N_21467);
and U21977 (N_21977,N_21108,N_21221);
nand U21978 (N_21978,N_21343,N_21336);
nand U21979 (N_21979,N_21239,N_21451);
nor U21980 (N_21980,N_21400,N_21256);
or U21981 (N_21981,N_21169,N_21019);
and U21982 (N_21982,N_21411,N_21268);
nand U21983 (N_21983,N_21053,N_21096);
nand U21984 (N_21984,N_21019,N_21176);
or U21985 (N_21985,N_21082,N_21239);
and U21986 (N_21986,N_21132,N_21079);
nor U21987 (N_21987,N_21079,N_21461);
and U21988 (N_21988,N_21119,N_21081);
xor U21989 (N_21989,N_21414,N_21386);
and U21990 (N_21990,N_21300,N_21269);
xor U21991 (N_21991,N_21292,N_21315);
nand U21992 (N_21992,N_21325,N_21497);
or U21993 (N_21993,N_21136,N_21377);
xnor U21994 (N_21994,N_21456,N_21448);
or U21995 (N_21995,N_21378,N_21192);
nand U21996 (N_21996,N_21061,N_21155);
and U21997 (N_21997,N_21212,N_21218);
and U21998 (N_21998,N_21089,N_21382);
nand U21999 (N_21999,N_21467,N_21432);
and U22000 (N_22000,N_21678,N_21930);
xnor U22001 (N_22001,N_21697,N_21557);
and U22002 (N_22002,N_21917,N_21534);
nor U22003 (N_22003,N_21919,N_21927);
and U22004 (N_22004,N_21967,N_21910);
xor U22005 (N_22005,N_21825,N_21833);
or U22006 (N_22006,N_21634,N_21716);
xor U22007 (N_22007,N_21998,N_21527);
nor U22008 (N_22008,N_21884,N_21845);
nor U22009 (N_22009,N_21658,N_21773);
xor U22010 (N_22010,N_21758,N_21511);
xnor U22011 (N_22011,N_21711,N_21821);
and U22012 (N_22012,N_21733,N_21705);
nand U22013 (N_22013,N_21620,N_21769);
xor U22014 (N_22014,N_21871,N_21581);
nor U22015 (N_22015,N_21928,N_21726);
nor U22016 (N_22016,N_21583,N_21513);
nand U22017 (N_22017,N_21706,N_21575);
nand U22018 (N_22018,N_21695,N_21935);
nand U22019 (N_22019,N_21606,N_21961);
nand U22020 (N_22020,N_21963,N_21731);
and U22021 (N_22021,N_21797,N_21756);
xor U22022 (N_22022,N_21549,N_21904);
and U22023 (N_22023,N_21937,N_21612);
and U22024 (N_22024,N_21569,N_21582);
xnor U22025 (N_22025,N_21799,N_21601);
xnor U22026 (N_22026,N_21991,N_21828);
or U22027 (N_22027,N_21692,N_21578);
or U22028 (N_22028,N_21512,N_21587);
nand U22029 (N_22029,N_21619,N_21889);
nand U22030 (N_22030,N_21616,N_21950);
or U22031 (N_22031,N_21929,N_21519);
xnor U22032 (N_22032,N_21816,N_21611);
or U22033 (N_22033,N_21891,N_21800);
or U22034 (N_22034,N_21536,N_21992);
and U22035 (N_22035,N_21514,N_21759);
nor U22036 (N_22036,N_21802,N_21547);
xnor U22037 (N_22037,N_21923,N_21528);
nand U22038 (N_22038,N_21674,N_21520);
and U22039 (N_22039,N_21651,N_21755);
nor U22040 (N_22040,N_21550,N_21903);
xnor U22041 (N_22041,N_21772,N_21783);
nor U22042 (N_22042,N_21595,N_21741);
nand U22043 (N_22043,N_21648,N_21883);
nor U22044 (N_22044,N_21691,N_21909);
nor U22045 (N_22045,N_21541,N_21771);
or U22046 (N_22046,N_21625,N_21907);
nor U22047 (N_22047,N_21842,N_21559);
nor U22048 (N_22048,N_21510,N_21949);
xor U22049 (N_22049,N_21742,N_21982);
xnor U22050 (N_22050,N_21894,N_21641);
and U22051 (N_22051,N_21867,N_21724);
or U22052 (N_22052,N_21996,N_21844);
or U22053 (N_22053,N_21934,N_21859);
xnor U22054 (N_22054,N_21675,N_21866);
and U22055 (N_22055,N_21526,N_21556);
nor U22056 (N_22056,N_21723,N_21886);
nand U22057 (N_22057,N_21503,N_21795);
xnor U22058 (N_22058,N_21926,N_21836);
or U22059 (N_22059,N_21743,N_21734);
and U22060 (N_22060,N_21668,N_21990);
and U22061 (N_22061,N_21945,N_21905);
or U22062 (N_22062,N_21857,N_21672);
xor U22063 (N_22063,N_21656,N_21822);
nor U22064 (N_22064,N_21993,N_21515);
nor U22065 (N_22065,N_21747,N_21545);
nor U22066 (N_22066,N_21679,N_21776);
nand U22067 (N_22067,N_21848,N_21570);
xnor U22068 (N_22068,N_21804,N_21732);
nand U22069 (N_22069,N_21596,N_21649);
nand U22070 (N_22070,N_21626,N_21631);
nand U22071 (N_22071,N_21636,N_21699);
nor U22072 (N_22072,N_21737,N_21818);
nor U22073 (N_22073,N_21829,N_21554);
or U22074 (N_22074,N_21947,N_21666);
xor U22075 (N_22075,N_21813,N_21968);
xnor U22076 (N_22076,N_21817,N_21688);
xnor U22077 (N_22077,N_21876,N_21878);
nor U22078 (N_22078,N_21805,N_21622);
and U22079 (N_22079,N_21718,N_21767);
nor U22080 (N_22080,N_21738,N_21750);
xnor U22081 (N_22081,N_21643,N_21975);
nand U22082 (N_22082,N_21887,N_21918);
and U22083 (N_22083,N_21940,N_21603);
nand U22084 (N_22084,N_21574,N_21739);
nor U22085 (N_22085,N_21779,N_21749);
and U22086 (N_22086,N_21555,N_21501);
xnor U22087 (N_22087,N_21689,N_21809);
nor U22088 (N_22088,N_21959,N_21915);
xnor U22089 (N_22089,N_21610,N_21702);
nor U22090 (N_22090,N_21785,N_21708);
nand U22091 (N_22091,N_21869,N_21644);
and U22092 (N_22092,N_21599,N_21953);
or U22093 (N_22093,N_21645,N_21714);
xnor U22094 (N_22094,N_21676,N_21593);
nand U22095 (N_22095,N_21812,N_21916);
nand U22096 (N_22096,N_21988,N_21647);
or U22097 (N_22097,N_21524,N_21703);
and U22098 (N_22098,N_21589,N_21529);
xnor U22099 (N_22099,N_21505,N_21815);
or U22100 (N_22100,N_21893,N_21720);
nor U22101 (N_22101,N_21725,N_21572);
xnor U22102 (N_22102,N_21908,N_21664);
nor U22103 (N_22103,N_21875,N_21814);
or U22104 (N_22104,N_21605,N_21826);
xor U22105 (N_22105,N_21850,N_21840);
or U22106 (N_22106,N_21573,N_21685);
and U22107 (N_22107,N_21538,N_21901);
and U22108 (N_22108,N_21969,N_21663);
or U22109 (N_22109,N_21775,N_21553);
nor U22110 (N_22110,N_21760,N_21540);
xor U22111 (N_22111,N_21687,N_21965);
or U22112 (N_22112,N_21820,N_21838);
nor U22113 (N_22113,N_21925,N_21964);
and U22114 (N_22114,N_21757,N_21660);
nand U22115 (N_22115,N_21696,N_21704);
nand U22116 (N_22116,N_21640,N_21786);
or U22117 (N_22117,N_21564,N_21667);
nand U22118 (N_22118,N_21933,N_21787);
xnor U22119 (N_22119,N_21966,N_21604);
nor U22120 (N_22120,N_21892,N_21618);
or U22121 (N_22121,N_21890,N_21806);
or U22122 (N_22122,N_21897,N_21985);
nand U22123 (N_22123,N_21698,N_21517);
or U22124 (N_22124,N_21584,N_21630);
nor U22125 (N_22125,N_21753,N_21751);
nand U22126 (N_22126,N_21763,N_21721);
nand U22127 (N_22127,N_21650,N_21877);
and U22128 (N_22128,N_21788,N_21989);
and U22129 (N_22129,N_21983,N_21868);
nor U22130 (N_22130,N_21843,N_21971);
and U22131 (N_22131,N_21880,N_21943);
nor U22132 (N_22132,N_21754,N_21854);
or U22133 (N_22133,N_21661,N_21782);
xor U22134 (N_22134,N_21946,N_21562);
xor U22135 (N_22135,N_21592,N_21994);
or U22136 (N_22136,N_21986,N_21936);
nor U22137 (N_22137,N_21567,N_21594);
nor U22138 (N_22138,N_21921,N_21899);
xor U22139 (N_22139,N_21521,N_21970);
nand U22140 (N_22140,N_21861,N_21712);
nand U22141 (N_22141,N_21765,N_21774);
xnor U22142 (N_22142,N_21745,N_21638);
or U22143 (N_22143,N_21849,N_21655);
xor U22144 (N_22144,N_21632,N_21987);
or U22145 (N_22145,N_21780,N_21939);
nor U22146 (N_22146,N_21748,N_21639);
xnor U22147 (N_22147,N_21671,N_21951);
xnor U22148 (N_22148,N_21944,N_21914);
nor U22149 (N_22149,N_21518,N_21700);
xnor U22150 (N_22150,N_21588,N_21981);
or U22151 (N_22151,N_21954,N_21823);
nor U22152 (N_22152,N_21542,N_21615);
xnor U22153 (N_22153,N_21853,N_21879);
xor U22154 (N_22154,N_21709,N_21865);
and U22155 (N_22155,N_21955,N_21977);
xor U22156 (N_22156,N_21938,N_21902);
or U22157 (N_22157,N_21932,N_21614);
nand U22158 (N_22158,N_21942,N_21624);
nand U22159 (N_22159,N_21803,N_21789);
xor U22160 (N_22160,N_21864,N_21607);
or U22161 (N_22161,N_21924,N_21922);
xor U22162 (N_22162,N_21681,N_21635);
and U22163 (N_22163,N_21654,N_21973);
and U22164 (N_22164,N_21997,N_21835);
xor U22165 (N_22165,N_21535,N_21621);
xnor U22166 (N_22166,N_21911,N_21531);
and U22167 (N_22167,N_21837,N_21677);
nor U22168 (N_22168,N_21960,N_21613);
and U22169 (N_22169,N_21847,N_21863);
nor U22170 (N_22170,N_21602,N_21623);
xor U22171 (N_22171,N_21686,N_21522);
nor U22172 (N_22172,N_21590,N_21752);
nor U22173 (N_22173,N_21552,N_21710);
xor U22174 (N_22174,N_21808,N_21796);
and U22175 (N_22175,N_21558,N_21834);
nand U22176 (N_22176,N_21683,N_21508);
nand U22177 (N_22177,N_21577,N_21778);
nand U22178 (N_22178,N_21713,N_21670);
xnor U22179 (N_22179,N_21931,N_21551);
xnor U22180 (N_22180,N_21860,N_21563);
nor U22181 (N_22181,N_21770,N_21855);
or U22182 (N_22182,N_21546,N_21827);
nand U22183 (N_22183,N_21662,N_21608);
or U22184 (N_22184,N_21565,N_21962);
nand U22185 (N_22185,N_21792,N_21768);
and U22186 (N_22186,N_21652,N_21539);
nor U22187 (N_22187,N_21858,N_21653);
xnor U22188 (N_22188,N_21707,N_21609);
nand U22189 (N_22189,N_21740,N_21730);
nand U22190 (N_22190,N_21715,N_21506);
nor U22191 (N_22191,N_21762,N_21585);
xnor U22192 (N_22192,N_21597,N_21735);
and U22193 (N_22193,N_21791,N_21537);
nand U22194 (N_22194,N_21995,N_21941);
nor U22195 (N_22195,N_21895,N_21717);
and U22196 (N_22196,N_21533,N_21657);
and U22197 (N_22197,N_21839,N_21500);
nand U22198 (N_22198,N_21896,N_21764);
and U22199 (N_22199,N_21972,N_21684);
or U22200 (N_22200,N_21722,N_21633);
or U22201 (N_22201,N_21790,N_21984);
and U22202 (N_22202,N_21682,N_21669);
nor U22203 (N_22203,N_21580,N_21888);
nor U22204 (N_22204,N_21976,N_21532);
xnor U22205 (N_22205,N_21956,N_21980);
and U22206 (N_22206,N_21824,N_21646);
xor U22207 (N_22207,N_21832,N_21862);
or U22208 (N_22208,N_21548,N_21637);
nor U22209 (N_22209,N_21576,N_21560);
and U22210 (N_22210,N_21665,N_21811);
nor U22211 (N_22211,N_21952,N_21507);
nor U22212 (N_22212,N_21798,N_21543);
or U22213 (N_22213,N_21974,N_21979);
nor U22214 (N_22214,N_21906,N_21680);
nand U22215 (N_22215,N_21801,N_21694);
xnor U22216 (N_22216,N_21777,N_21874);
and U22217 (N_22217,N_21746,N_21617);
or U22218 (N_22218,N_21841,N_21628);
xor U22219 (N_22219,N_21729,N_21856);
and U22220 (N_22220,N_21846,N_21807);
or U22221 (N_22221,N_21744,N_21544);
nand U22222 (N_22222,N_21852,N_21693);
and U22223 (N_22223,N_21642,N_21502);
or U22224 (N_22224,N_21579,N_21873);
and U22225 (N_22225,N_21598,N_21516);
nand U22226 (N_22226,N_21784,N_21659);
and U22227 (N_22227,N_21872,N_21999);
nand U22228 (N_22228,N_21978,N_21673);
nand U22229 (N_22229,N_21870,N_21571);
nand U22230 (N_22230,N_21882,N_21948);
xnor U22231 (N_22231,N_21881,N_21690);
nor U22232 (N_22232,N_21810,N_21600);
xor U22233 (N_22233,N_21920,N_21851);
nor U22234 (N_22234,N_21728,N_21568);
nand U22235 (N_22235,N_21561,N_21761);
nor U22236 (N_22236,N_21958,N_21900);
and U22237 (N_22237,N_21627,N_21530);
xnor U22238 (N_22238,N_21566,N_21504);
nor U22239 (N_22239,N_21727,N_21719);
xnor U22240 (N_22240,N_21830,N_21819);
and U22241 (N_22241,N_21629,N_21523);
nor U22242 (N_22242,N_21912,N_21591);
and U22243 (N_22243,N_21525,N_21898);
nand U22244 (N_22244,N_21913,N_21509);
nor U22245 (N_22245,N_21885,N_21586);
and U22246 (N_22246,N_21957,N_21701);
or U22247 (N_22247,N_21736,N_21794);
or U22248 (N_22248,N_21793,N_21831);
nand U22249 (N_22249,N_21766,N_21781);
xnor U22250 (N_22250,N_21595,N_21542);
and U22251 (N_22251,N_21622,N_21598);
or U22252 (N_22252,N_21721,N_21894);
and U22253 (N_22253,N_21851,N_21628);
and U22254 (N_22254,N_21796,N_21744);
nand U22255 (N_22255,N_21781,N_21996);
or U22256 (N_22256,N_21617,N_21920);
xor U22257 (N_22257,N_21793,N_21674);
and U22258 (N_22258,N_21526,N_21935);
nand U22259 (N_22259,N_21633,N_21571);
and U22260 (N_22260,N_21500,N_21859);
nand U22261 (N_22261,N_21674,N_21904);
or U22262 (N_22262,N_21652,N_21536);
or U22263 (N_22263,N_21878,N_21655);
and U22264 (N_22264,N_21835,N_21891);
and U22265 (N_22265,N_21610,N_21994);
or U22266 (N_22266,N_21914,N_21907);
nand U22267 (N_22267,N_21564,N_21638);
and U22268 (N_22268,N_21974,N_21661);
nand U22269 (N_22269,N_21869,N_21618);
xor U22270 (N_22270,N_21522,N_21913);
nand U22271 (N_22271,N_21552,N_21706);
or U22272 (N_22272,N_21565,N_21696);
nand U22273 (N_22273,N_21657,N_21773);
xnor U22274 (N_22274,N_21797,N_21811);
nor U22275 (N_22275,N_21806,N_21768);
or U22276 (N_22276,N_21846,N_21754);
or U22277 (N_22277,N_21557,N_21928);
nor U22278 (N_22278,N_21968,N_21865);
nor U22279 (N_22279,N_21788,N_21999);
nor U22280 (N_22280,N_21564,N_21738);
and U22281 (N_22281,N_21849,N_21621);
nor U22282 (N_22282,N_21854,N_21656);
xnor U22283 (N_22283,N_21712,N_21792);
or U22284 (N_22284,N_21930,N_21747);
nand U22285 (N_22285,N_21729,N_21772);
nand U22286 (N_22286,N_21792,N_21913);
nand U22287 (N_22287,N_21797,N_21553);
nand U22288 (N_22288,N_21875,N_21526);
nor U22289 (N_22289,N_21779,N_21581);
xnor U22290 (N_22290,N_21985,N_21705);
or U22291 (N_22291,N_21567,N_21722);
nor U22292 (N_22292,N_21707,N_21978);
or U22293 (N_22293,N_21678,N_21700);
and U22294 (N_22294,N_21724,N_21625);
nor U22295 (N_22295,N_21660,N_21652);
nor U22296 (N_22296,N_21813,N_21965);
nor U22297 (N_22297,N_21623,N_21872);
and U22298 (N_22298,N_21634,N_21602);
xnor U22299 (N_22299,N_21616,N_21778);
xor U22300 (N_22300,N_21897,N_21930);
and U22301 (N_22301,N_21974,N_21670);
nor U22302 (N_22302,N_21651,N_21745);
nor U22303 (N_22303,N_21944,N_21831);
xor U22304 (N_22304,N_21883,N_21896);
nor U22305 (N_22305,N_21857,N_21684);
nor U22306 (N_22306,N_21852,N_21689);
xor U22307 (N_22307,N_21973,N_21934);
or U22308 (N_22308,N_21770,N_21815);
and U22309 (N_22309,N_21705,N_21825);
and U22310 (N_22310,N_21507,N_21937);
xnor U22311 (N_22311,N_21892,N_21675);
nand U22312 (N_22312,N_21630,N_21635);
nor U22313 (N_22313,N_21808,N_21943);
and U22314 (N_22314,N_21915,N_21735);
or U22315 (N_22315,N_21807,N_21984);
nor U22316 (N_22316,N_21735,N_21737);
nor U22317 (N_22317,N_21963,N_21510);
xnor U22318 (N_22318,N_21826,N_21917);
and U22319 (N_22319,N_21896,N_21521);
nor U22320 (N_22320,N_21560,N_21856);
and U22321 (N_22321,N_21557,N_21519);
nand U22322 (N_22322,N_21995,N_21532);
or U22323 (N_22323,N_21693,N_21543);
nand U22324 (N_22324,N_21899,N_21564);
xor U22325 (N_22325,N_21636,N_21790);
xnor U22326 (N_22326,N_21986,N_21604);
or U22327 (N_22327,N_21664,N_21786);
or U22328 (N_22328,N_21733,N_21915);
xnor U22329 (N_22329,N_21501,N_21681);
and U22330 (N_22330,N_21834,N_21799);
xor U22331 (N_22331,N_21628,N_21860);
and U22332 (N_22332,N_21834,N_21605);
nand U22333 (N_22333,N_21791,N_21974);
nand U22334 (N_22334,N_21936,N_21539);
and U22335 (N_22335,N_21605,N_21529);
nand U22336 (N_22336,N_21947,N_21839);
or U22337 (N_22337,N_21920,N_21692);
or U22338 (N_22338,N_21502,N_21954);
nand U22339 (N_22339,N_21569,N_21810);
nor U22340 (N_22340,N_21836,N_21769);
nor U22341 (N_22341,N_21885,N_21883);
or U22342 (N_22342,N_21726,N_21580);
nand U22343 (N_22343,N_21710,N_21894);
xor U22344 (N_22344,N_21972,N_21622);
xor U22345 (N_22345,N_21536,N_21577);
nor U22346 (N_22346,N_21547,N_21897);
nor U22347 (N_22347,N_21861,N_21635);
xnor U22348 (N_22348,N_21538,N_21930);
or U22349 (N_22349,N_21937,N_21627);
nor U22350 (N_22350,N_21798,N_21762);
and U22351 (N_22351,N_21723,N_21613);
xnor U22352 (N_22352,N_21783,N_21642);
xor U22353 (N_22353,N_21762,N_21976);
nand U22354 (N_22354,N_21525,N_21686);
nand U22355 (N_22355,N_21643,N_21577);
nor U22356 (N_22356,N_21719,N_21638);
and U22357 (N_22357,N_21600,N_21593);
and U22358 (N_22358,N_21856,N_21612);
nor U22359 (N_22359,N_21590,N_21925);
nand U22360 (N_22360,N_21703,N_21613);
or U22361 (N_22361,N_21733,N_21609);
xnor U22362 (N_22362,N_21686,N_21578);
xor U22363 (N_22363,N_21545,N_21769);
and U22364 (N_22364,N_21776,N_21795);
nand U22365 (N_22365,N_21639,N_21837);
and U22366 (N_22366,N_21806,N_21609);
and U22367 (N_22367,N_21500,N_21596);
and U22368 (N_22368,N_21751,N_21546);
nor U22369 (N_22369,N_21648,N_21930);
nor U22370 (N_22370,N_21874,N_21663);
xor U22371 (N_22371,N_21577,N_21929);
nand U22372 (N_22372,N_21847,N_21666);
and U22373 (N_22373,N_21881,N_21936);
nand U22374 (N_22374,N_21662,N_21659);
and U22375 (N_22375,N_21865,N_21540);
nand U22376 (N_22376,N_21881,N_21753);
and U22377 (N_22377,N_21542,N_21892);
nand U22378 (N_22378,N_21785,N_21581);
and U22379 (N_22379,N_21528,N_21720);
xnor U22380 (N_22380,N_21664,N_21836);
xor U22381 (N_22381,N_21698,N_21952);
nand U22382 (N_22382,N_21929,N_21909);
nand U22383 (N_22383,N_21831,N_21764);
nand U22384 (N_22384,N_21970,N_21707);
xnor U22385 (N_22385,N_21844,N_21700);
xnor U22386 (N_22386,N_21975,N_21990);
nor U22387 (N_22387,N_21621,N_21660);
or U22388 (N_22388,N_21697,N_21861);
xor U22389 (N_22389,N_21554,N_21711);
and U22390 (N_22390,N_21740,N_21720);
and U22391 (N_22391,N_21948,N_21957);
nor U22392 (N_22392,N_21600,N_21823);
nor U22393 (N_22393,N_21841,N_21825);
and U22394 (N_22394,N_21673,N_21567);
xnor U22395 (N_22395,N_21918,N_21576);
nor U22396 (N_22396,N_21753,N_21937);
nand U22397 (N_22397,N_21713,N_21817);
and U22398 (N_22398,N_21909,N_21828);
nor U22399 (N_22399,N_21804,N_21780);
nand U22400 (N_22400,N_21829,N_21960);
nor U22401 (N_22401,N_21844,N_21999);
nand U22402 (N_22402,N_21541,N_21607);
and U22403 (N_22403,N_21502,N_21731);
nor U22404 (N_22404,N_21599,N_21671);
or U22405 (N_22405,N_21728,N_21986);
nand U22406 (N_22406,N_21877,N_21863);
nor U22407 (N_22407,N_21728,N_21585);
nor U22408 (N_22408,N_21713,N_21729);
or U22409 (N_22409,N_21699,N_21940);
and U22410 (N_22410,N_21865,N_21960);
and U22411 (N_22411,N_21785,N_21806);
and U22412 (N_22412,N_21666,N_21922);
or U22413 (N_22413,N_21731,N_21500);
and U22414 (N_22414,N_21712,N_21967);
nor U22415 (N_22415,N_21877,N_21866);
nand U22416 (N_22416,N_21975,N_21817);
nor U22417 (N_22417,N_21856,N_21508);
nand U22418 (N_22418,N_21940,N_21559);
nor U22419 (N_22419,N_21918,N_21899);
or U22420 (N_22420,N_21779,N_21624);
and U22421 (N_22421,N_21621,N_21834);
xnor U22422 (N_22422,N_21957,N_21527);
and U22423 (N_22423,N_21812,N_21980);
xor U22424 (N_22424,N_21731,N_21899);
xor U22425 (N_22425,N_21683,N_21722);
or U22426 (N_22426,N_21570,N_21711);
nand U22427 (N_22427,N_21532,N_21708);
nand U22428 (N_22428,N_21764,N_21870);
nand U22429 (N_22429,N_21567,N_21688);
xnor U22430 (N_22430,N_21563,N_21865);
nor U22431 (N_22431,N_21696,N_21600);
nor U22432 (N_22432,N_21890,N_21638);
and U22433 (N_22433,N_21599,N_21788);
nor U22434 (N_22434,N_21617,N_21776);
nand U22435 (N_22435,N_21699,N_21966);
or U22436 (N_22436,N_21735,N_21703);
xor U22437 (N_22437,N_21876,N_21705);
xnor U22438 (N_22438,N_21674,N_21852);
xor U22439 (N_22439,N_21597,N_21566);
nand U22440 (N_22440,N_21798,N_21981);
nor U22441 (N_22441,N_21984,N_21885);
or U22442 (N_22442,N_21818,N_21771);
xor U22443 (N_22443,N_21896,N_21990);
nor U22444 (N_22444,N_21640,N_21668);
nand U22445 (N_22445,N_21841,N_21986);
and U22446 (N_22446,N_21511,N_21990);
and U22447 (N_22447,N_21623,N_21593);
xor U22448 (N_22448,N_21578,N_21823);
xnor U22449 (N_22449,N_21547,N_21824);
and U22450 (N_22450,N_21660,N_21517);
and U22451 (N_22451,N_21949,N_21681);
and U22452 (N_22452,N_21613,N_21746);
and U22453 (N_22453,N_21649,N_21967);
nand U22454 (N_22454,N_21520,N_21779);
and U22455 (N_22455,N_21682,N_21986);
nor U22456 (N_22456,N_21894,N_21739);
and U22457 (N_22457,N_21711,N_21714);
or U22458 (N_22458,N_21737,N_21967);
or U22459 (N_22459,N_21949,N_21984);
xnor U22460 (N_22460,N_21815,N_21929);
xor U22461 (N_22461,N_21546,N_21579);
or U22462 (N_22462,N_21626,N_21720);
xor U22463 (N_22463,N_21936,N_21925);
xor U22464 (N_22464,N_21710,N_21645);
nor U22465 (N_22465,N_21765,N_21533);
or U22466 (N_22466,N_21840,N_21709);
and U22467 (N_22467,N_21903,N_21969);
and U22468 (N_22468,N_21891,N_21507);
and U22469 (N_22469,N_21885,N_21888);
nor U22470 (N_22470,N_21736,N_21774);
xor U22471 (N_22471,N_21703,N_21907);
nor U22472 (N_22472,N_21687,N_21519);
nand U22473 (N_22473,N_21805,N_21679);
xor U22474 (N_22474,N_21836,N_21569);
nor U22475 (N_22475,N_21990,N_21939);
nor U22476 (N_22476,N_21950,N_21857);
or U22477 (N_22477,N_21763,N_21869);
nand U22478 (N_22478,N_21663,N_21628);
and U22479 (N_22479,N_21983,N_21893);
and U22480 (N_22480,N_21741,N_21514);
xor U22481 (N_22481,N_21898,N_21557);
and U22482 (N_22482,N_21528,N_21547);
or U22483 (N_22483,N_21720,N_21501);
nand U22484 (N_22484,N_21662,N_21524);
xor U22485 (N_22485,N_21570,N_21935);
xor U22486 (N_22486,N_21503,N_21904);
and U22487 (N_22487,N_21903,N_21915);
nor U22488 (N_22488,N_21728,N_21904);
xnor U22489 (N_22489,N_21998,N_21819);
nor U22490 (N_22490,N_21578,N_21702);
nor U22491 (N_22491,N_21959,N_21591);
or U22492 (N_22492,N_21576,N_21586);
nand U22493 (N_22493,N_21974,N_21505);
xor U22494 (N_22494,N_21622,N_21981);
xnor U22495 (N_22495,N_21668,N_21897);
nor U22496 (N_22496,N_21554,N_21529);
nor U22497 (N_22497,N_21618,N_21627);
nor U22498 (N_22498,N_21639,N_21702);
xnor U22499 (N_22499,N_21514,N_21791);
nor U22500 (N_22500,N_22354,N_22012);
nand U22501 (N_22501,N_22101,N_22088);
xor U22502 (N_22502,N_22257,N_22138);
xor U22503 (N_22503,N_22258,N_22104);
or U22504 (N_22504,N_22166,N_22150);
nor U22505 (N_22505,N_22411,N_22145);
xor U22506 (N_22506,N_22372,N_22248);
xor U22507 (N_22507,N_22063,N_22427);
or U22508 (N_22508,N_22139,N_22426);
or U22509 (N_22509,N_22470,N_22475);
nand U22510 (N_22510,N_22234,N_22238);
and U22511 (N_22511,N_22442,N_22283);
xnor U22512 (N_22512,N_22018,N_22186);
or U22513 (N_22513,N_22105,N_22221);
or U22514 (N_22514,N_22276,N_22013);
nor U22515 (N_22515,N_22130,N_22264);
xor U22516 (N_22516,N_22022,N_22259);
and U22517 (N_22517,N_22240,N_22453);
and U22518 (N_22518,N_22297,N_22394);
or U22519 (N_22519,N_22436,N_22312);
xor U22520 (N_22520,N_22144,N_22398);
or U22521 (N_22521,N_22143,N_22383);
and U22522 (N_22522,N_22050,N_22365);
nand U22523 (N_22523,N_22195,N_22483);
nor U22524 (N_22524,N_22054,N_22302);
or U22525 (N_22525,N_22147,N_22493);
or U22526 (N_22526,N_22447,N_22111);
nor U22527 (N_22527,N_22078,N_22304);
xnor U22528 (N_22528,N_22488,N_22106);
nor U22529 (N_22529,N_22115,N_22128);
nor U22530 (N_22530,N_22017,N_22038);
or U22531 (N_22531,N_22396,N_22112);
xor U22532 (N_22532,N_22005,N_22065);
nand U22533 (N_22533,N_22167,N_22352);
nor U22534 (N_22534,N_22096,N_22321);
and U22535 (N_22535,N_22430,N_22349);
nand U22536 (N_22536,N_22410,N_22045);
and U22537 (N_22537,N_22351,N_22343);
or U22538 (N_22538,N_22233,N_22204);
or U22539 (N_22539,N_22253,N_22353);
nor U22540 (N_22540,N_22420,N_22189);
nand U22541 (N_22541,N_22319,N_22114);
or U22542 (N_22542,N_22367,N_22194);
xor U22543 (N_22543,N_22217,N_22132);
nor U22544 (N_22544,N_22187,N_22039);
xor U22545 (N_22545,N_22040,N_22268);
and U22546 (N_22546,N_22279,N_22043);
and U22547 (N_22547,N_22051,N_22382);
nand U22548 (N_22548,N_22228,N_22177);
xnor U22549 (N_22549,N_22429,N_22026);
or U22550 (N_22550,N_22237,N_22301);
nand U22551 (N_22551,N_22211,N_22361);
nand U22552 (N_22552,N_22317,N_22363);
nand U22553 (N_22553,N_22030,N_22216);
and U22554 (N_22554,N_22338,N_22417);
nor U22555 (N_22555,N_22327,N_22048);
and U22556 (N_22556,N_22289,N_22094);
xnor U22557 (N_22557,N_22056,N_22295);
and U22558 (N_22558,N_22294,N_22015);
xnor U22559 (N_22559,N_22061,N_22073);
nand U22560 (N_22560,N_22440,N_22368);
nor U22561 (N_22561,N_22346,N_22097);
or U22562 (N_22562,N_22154,N_22247);
or U22563 (N_22563,N_22270,N_22116);
and U22564 (N_22564,N_22122,N_22308);
xnor U22565 (N_22565,N_22403,N_22454);
nor U22566 (N_22566,N_22291,N_22451);
xor U22567 (N_22567,N_22163,N_22311);
or U22568 (N_22568,N_22318,N_22445);
xnor U22569 (N_22569,N_22497,N_22266);
and U22570 (N_22570,N_22439,N_22472);
nand U22571 (N_22571,N_22332,N_22347);
xnor U22572 (N_22572,N_22405,N_22255);
and U22573 (N_22573,N_22009,N_22498);
or U22574 (N_22574,N_22156,N_22466);
or U22575 (N_22575,N_22029,N_22322);
and U22576 (N_22576,N_22070,N_22408);
nand U22577 (N_22577,N_22016,N_22386);
nand U22578 (N_22578,N_22371,N_22159);
nor U22579 (N_22579,N_22397,N_22236);
or U22580 (N_22580,N_22437,N_22335);
and U22581 (N_22581,N_22305,N_22377);
nand U22582 (N_22582,N_22188,N_22066);
and U22583 (N_22583,N_22339,N_22269);
and U22584 (N_22584,N_22084,N_22197);
nor U22585 (N_22585,N_22409,N_22249);
or U22586 (N_22586,N_22239,N_22362);
xor U22587 (N_22587,N_22041,N_22370);
or U22588 (N_22588,N_22281,N_22406);
xor U22589 (N_22589,N_22285,N_22243);
or U22590 (N_22590,N_22441,N_22288);
nor U22591 (N_22591,N_22213,N_22328);
or U22592 (N_22592,N_22345,N_22395);
or U22593 (N_22593,N_22284,N_22256);
or U22594 (N_22594,N_22496,N_22200);
xnor U22595 (N_22595,N_22059,N_22171);
or U22596 (N_22596,N_22082,N_22032);
nor U22597 (N_22597,N_22080,N_22024);
and U22598 (N_22598,N_22309,N_22303);
xnor U22599 (N_22599,N_22344,N_22476);
nor U22600 (N_22600,N_22485,N_22174);
nor U22601 (N_22601,N_22047,N_22385);
xnor U22602 (N_22602,N_22314,N_22090);
and U22603 (N_22603,N_22412,N_22337);
nand U22604 (N_22604,N_22086,N_22422);
nor U22605 (N_22605,N_22468,N_22350);
or U22606 (N_22606,N_22108,N_22356);
or U22607 (N_22607,N_22117,N_22263);
and U22608 (N_22608,N_22444,N_22275);
nor U22609 (N_22609,N_22452,N_22103);
nor U22610 (N_22610,N_22359,N_22494);
xor U22611 (N_22611,N_22495,N_22191);
xor U22612 (N_22612,N_22374,N_22089);
nand U22613 (N_22613,N_22230,N_22486);
nor U22614 (N_22614,N_22260,N_22055);
and U22615 (N_22615,N_22164,N_22298);
or U22616 (N_22616,N_22180,N_22028);
or U22617 (N_22617,N_22225,N_22379);
or U22618 (N_22618,N_22340,N_22250);
and U22619 (N_22619,N_22146,N_22124);
nor U22620 (N_22620,N_22182,N_22058);
xnor U22621 (N_22621,N_22300,N_22099);
nand U22622 (N_22622,N_22196,N_22052);
nor U22623 (N_22623,N_22469,N_22183);
xnor U22624 (N_22624,N_22241,N_22219);
and U22625 (N_22625,N_22387,N_22252);
and U22626 (N_22626,N_22490,N_22169);
xnor U22627 (N_22627,N_22160,N_22118);
xor U22628 (N_22628,N_22181,N_22480);
and U22629 (N_22629,N_22210,N_22165);
nor U22630 (N_22630,N_22399,N_22325);
nand U22631 (N_22631,N_22273,N_22330);
xnor U22632 (N_22632,N_22098,N_22198);
or U22633 (N_22633,N_22113,N_22320);
xnor U22634 (N_22634,N_22334,N_22120);
xor U22635 (N_22635,N_22119,N_22037);
and U22636 (N_22636,N_22244,N_22381);
nor U22637 (N_22637,N_22172,N_22267);
nor U22638 (N_22638,N_22432,N_22060);
nand U22639 (N_22639,N_22404,N_22036);
xnor U22640 (N_22640,N_22373,N_22499);
xnor U22641 (N_22641,N_22460,N_22072);
nand U22642 (N_22642,N_22401,N_22313);
or U22643 (N_22643,N_22185,N_22175);
or U22644 (N_22644,N_22232,N_22014);
and U22645 (N_22645,N_22455,N_22315);
nor U22646 (N_22646,N_22134,N_22202);
xnor U22647 (N_22647,N_22133,N_22464);
and U22648 (N_22648,N_22007,N_22482);
xor U22649 (N_22649,N_22075,N_22087);
xor U22650 (N_22650,N_22481,N_22074);
xor U22651 (N_22651,N_22076,N_22042);
xor U22652 (N_22652,N_22023,N_22388);
or U22653 (N_22653,N_22158,N_22215);
and U22654 (N_22654,N_22004,N_22380);
and U22655 (N_22655,N_22431,N_22272);
nor U22656 (N_22656,N_22246,N_22254);
xor U22657 (N_22657,N_22278,N_22077);
or U22658 (N_22658,N_22110,N_22364);
nor U22659 (N_22659,N_22418,N_22001);
nand U22660 (N_22660,N_22173,N_22020);
nor U22661 (N_22661,N_22433,N_22391);
nand U22662 (N_22662,N_22282,N_22235);
and U22663 (N_22663,N_22067,N_22292);
xnor U22664 (N_22664,N_22324,N_22000);
and U22665 (N_22665,N_22136,N_22127);
nor U22666 (N_22666,N_22025,N_22473);
and U22667 (N_22667,N_22223,N_22226);
or U22668 (N_22668,N_22207,N_22416);
and U22669 (N_22669,N_22425,N_22393);
nor U22670 (N_22670,N_22389,N_22019);
nand U22671 (N_22671,N_22456,N_22192);
nor U22672 (N_22672,N_22044,N_22378);
or U22673 (N_22673,N_22449,N_22142);
and U22674 (N_22674,N_22224,N_22205);
or U22675 (N_22675,N_22179,N_22137);
nor U22676 (N_22676,N_22438,N_22290);
nor U22677 (N_22677,N_22277,N_22203);
xor U22678 (N_22678,N_22027,N_22492);
and U22679 (N_22679,N_22125,N_22326);
nand U22680 (N_22680,N_22414,N_22222);
or U22681 (N_22681,N_22390,N_22446);
or U22682 (N_22682,N_22419,N_22458);
and U22683 (N_22683,N_22126,N_22218);
xnor U22684 (N_22684,N_22467,N_22161);
xor U22685 (N_22685,N_22057,N_22450);
xor U22686 (N_22686,N_22231,N_22095);
and U22687 (N_22687,N_22428,N_22474);
or U22688 (N_22688,N_22357,N_22049);
nand U22689 (N_22689,N_22184,N_22129);
or U22690 (N_22690,N_22011,N_22068);
xor U22691 (N_22691,N_22162,N_22034);
or U22692 (N_22692,N_22245,N_22471);
nor U22693 (N_22693,N_22081,N_22155);
and U22694 (N_22694,N_22376,N_22369);
xnor U22695 (N_22695,N_22168,N_22107);
and U22696 (N_22696,N_22287,N_22021);
xor U22697 (N_22697,N_22153,N_22033);
and U22698 (N_22698,N_22157,N_22421);
nand U22699 (N_22699,N_22131,N_22358);
xor U22700 (N_22700,N_22448,N_22190);
and U22701 (N_22701,N_22491,N_22229);
or U22702 (N_22702,N_22206,N_22375);
and U22703 (N_22703,N_22400,N_22331);
and U22704 (N_22704,N_22461,N_22342);
xnor U22705 (N_22705,N_22053,N_22462);
nor U22706 (N_22706,N_22274,N_22227);
and U22707 (N_22707,N_22434,N_22193);
and U22708 (N_22708,N_22092,N_22392);
or U22709 (N_22709,N_22293,N_22280);
xor U22710 (N_22710,N_22307,N_22006);
or U22711 (N_22711,N_22008,N_22083);
and U22712 (N_22712,N_22316,N_22271);
nor U22713 (N_22713,N_22010,N_22069);
or U22714 (N_22714,N_22151,N_22178);
and U22715 (N_22715,N_22152,N_22085);
and U22716 (N_22716,N_22208,N_22212);
xnor U22717 (N_22717,N_22123,N_22402);
or U22718 (N_22718,N_22384,N_22170);
or U22719 (N_22719,N_22413,N_22306);
and U22720 (N_22720,N_22484,N_22435);
nand U22721 (N_22721,N_22140,N_22199);
nand U22722 (N_22722,N_22220,N_22093);
nand U22723 (N_22723,N_22487,N_22415);
nand U22724 (N_22724,N_22176,N_22355);
nor U22725 (N_22725,N_22002,N_22242);
and U22726 (N_22726,N_22477,N_22333);
and U22727 (N_22727,N_22102,N_22214);
nand U22728 (N_22728,N_22360,N_22031);
or U22729 (N_22729,N_22091,N_22296);
or U22730 (N_22730,N_22003,N_22341);
xnor U22731 (N_22731,N_22035,N_22457);
nor U22732 (N_22732,N_22423,N_22463);
nor U22733 (N_22733,N_22148,N_22329);
xnor U22734 (N_22734,N_22109,N_22201);
or U22735 (N_22735,N_22121,N_22265);
nor U22736 (N_22736,N_22443,N_22407);
nor U22737 (N_22737,N_22459,N_22062);
and U22738 (N_22738,N_22479,N_22336);
and U22739 (N_22739,N_22251,N_22310);
and U22740 (N_22740,N_22348,N_22262);
and U22741 (N_22741,N_22141,N_22424);
xor U22742 (N_22742,N_22135,N_22064);
and U22743 (N_22743,N_22323,N_22149);
nor U22744 (N_22744,N_22366,N_22489);
and U22745 (N_22745,N_22046,N_22100);
xor U22746 (N_22746,N_22079,N_22286);
nor U22747 (N_22747,N_22465,N_22261);
nand U22748 (N_22748,N_22299,N_22209);
xnor U22749 (N_22749,N_22071,N_22478);
xnor U22750 (N_22750,N_22441,N_22403);
xnor U22751 (N_22751,N_22182,N_22398);
and U22752 (N_22752,N_22145,N_22455);
xor U22753 (N_22753,N_22396,N_22441);
xor U22754 (N_22754,N_22413,N_22439);
or U22755 (N_22755,N_22033,N_22223);
or U22756 (N_22756,N_22279,N_22263);
or U22757 (N_22757,N_22367,N_22112);
nor U22758 (N_22758,N_22401,N_22464);
nand U22759 (N_22759,N_22374,N_22323);
or U22760 (N_22760,N_22212,N_22102);
nand U22761 (N_22761,N_22000,N_22342);
xor U22762 (N_22762,N_22427,N_22320);
or U22763 (N_22763,N_22205,N_22447);
xor U22764 (N_22764,N_22106,N_22334);
nand U22765 (N_22765,N_22092,N_22008);
xor U22766 (N_22766,N_22091,N_22276);
xnor U22767 (N_22767,N_22362,N_22184);
and U22768 (N_22768,N_22176,N_22348);
nand U22769 (N_22769,N_22337,N_22371);
and U22770 (N_22770,N_22029,N_22479);
nor U22771 (N_22771,N_22292,N_22430);
nand U22772 (N_22772,N_22426,N_22480);
or U22773 (N_22773,N_22411,N_22353);
or U22774 (N_22774,N_22372,N_22034);
and U22775 (N_22775,N_22362,N_22477);
and U22776 (N_22776,N_22054,N_22261);
or U22777 (N_22777,N_22222,N_22252);
xnor U22778 (N_22778,N_22499,N_22475);
and U22779 (N_22779,N_22184,N_22156);
or U22780 (N_22780,N_22037,N_22173);
and U22781 (N_22781,N_22098,N_22173);
nand U22782 (N_22782,N_22233,N_22155);
and U22783 (N_22783,N_22188,N_22236);
nand U22784 (N_22784,N_22101,N_22290);
nand U22785 (N_22785,N_22485,N_22098);
nor U22786 (N_22786,N_22391,N_22296);
xor U22787 (N_22787,N_22174,N_22152);
or U22788 (N_22788,N_22452,N_22400);
or U22789 (N_22789,N_22348,N_22300);
nor U22790 (N_22790,N_22008,N_22005);
or U22791 (N_22791,N_22200,N_22474);
nand U22792 (N_22792,N_22369,N_22186);
and U22793 (N_22793,N_22276,N_22099);
xor U22794 (N_22794,N_22075,N_22497);
xnor U22795 (N_22795,N_22489,N_22245);
nand U22796 (N_22796,N_22191,N_22249);
or U22797 (N_22797,N_22091,N_22180);
or U22798 (N_22798,N_22266,N_22118);
xor U22799 (N_22799,N_22334,N_22263);
or U22800 (N_22800,N_22390,N_22434);
nand U22801 (N_22801,N_22309,N_22328);
xnor U22802 (N_22802,N_22035,N_22484);
and U22803 (N_22803,N_22246,N_22495);
and U22804 (N_22804,N_22021,N_22357);
nor U22805 (N_22805,N_22410,N_22047);
nor U22806 (N_22806,N_22324,N_22471);
and U22807 (N_22807,N_22408,N_22245);
nor U22808 (N_22808,N_22484,N_22342);
nor U22809 (N_22809,N_22305,N_22460);
nand U22810 (N_22810,N_22347,N_22417);
nand U22811 (N_22811,N_22321,N_22059);
and U22812 (N_22812,N_22398,N_22049);
and U22813 (N_22813,N_22445,N_22410);
nand U22814 (N_22814,N_22328,N_22240);
nand U22815 (N_22815,N_22057,N_22288);
xnor U22816 (N_22816,N_22214,N_22314);
or U22817 (N_22817,N_22204,N_22247);
or U22818 (N_22818,N_22055,N_22402);
nand U22819 (N_22819,N_22278,N_22432);
xnor U22820 (N_22820,N_22208,N_22363);
or U22821 (N_22821,N_22458,N_22474);
and U22822 (N_22822,N_22216,N_22290);
or U22823 (N_22823,N_22448,N_22340);
nand U22824 (N_22824,N_22360,N_22424);
xor U22825 (N_22825,N_22059,N_22264);
xnor U22826 (N_22826,N_22110,N_22398);
and U22827 (N_22827,N_22175,N_22340);
and U22828 (N_22828,N_22302,N_22361);
nor U22829 (N_22829,N_22076,N_22093);
or U22830 (N_22830,N_22198,N_22046);
or U22831 (N_22831,N_22105,N_22381);
xnor U22832 (N_22832,N_22174,N_22040);
xnor U22833 (N_22833,N_22278,N_22152);
xor U22834 (N_22834,N_22283,N_22219);
nand U22835 (N_22835,N_22252,N_22010);
and U22836 (N_22836,N_22055,N_22090);
nand U22837 (N_22837,N_22148,N_22106);
nand U22838 (N_22838,N_22483,N_22257);
nor U22839 (N_22839,N_22023,N_22292);
nand U22840 (N_22840,N_22016,N_22191);
xnor U22841 (N_22841,N_22202,N_22208);
nor U22842 (N_22842,N_22211,N_22263);
xor U22843 (N_22843,N_22195,N_22106);
and U22844 (N_22844,N_22344,N_22152);
or U22845 (N_22845,N_22407,N_22148);
xor U22846 (N_22846,N_22399,N_22257);
nand U22847 (N_22847,N_22251,N_22174);
nand U22848 (N_22848,N_22174,N_22460);
and U22849 (N_22849,N_22039,N_22248);
and U22850 (N_22850,N_22351,N_22472);
nor U22851 (N_22851,N_22067,N_22234);
xor U22852 (N_22852,N_22117,N_22186);
nor U22853 (N_22853,N_22265,N_22295);
xor U22854 (N_22854,N_22334,N_22294);
and U22855 (N_22855,N_22497,N_22240);
and U22856 (N_22856,N_22269,N_22305);
nor U22857 (N_22857,N_22085,N_22126);
nor U22858 (N_22858,N_22184,N_22343);
or U22859 (N_22859,N_22482,N_22147);
xor U22860 (N_22860,N_22312,N_22332);
and U22861 (N_22861,N_22344,N_22133);
and U22862 (N_22862,N_22394,N_22207);
nand U22863 (N_22863,N_22364,N_22465);
nor U22864 (N_22864,N_22305,N_22412);
nor U22865 (N_22865,N_22186,N_22260);
or U22866 (N_22866,N_22170,N_22053);
or U22867 (N_22867,N_22243,N_22269);
nor U22868 (N_22868,N_22484,N_22221);
nand U22869 (N_22869,N_22334,N_22340);
or U22870 (N_22870,N_22376,N_22190);
or U22871 (N_22871,N_22351,N_22378);
or U22872 (N_22872,N_22308,N_22427);
nor U22873 (N_22873,N_22139,N_22363);
xor U22874 (N_22874,N_22135,N_22050);
or U22875 (N_22875,N_22489,N_22428);
nand U22876 (N_22876,N_22447,N_22251);
or U22877 (N_22877,N_22097,N_22210);
or U22878 (N_22878,N_22038,N_22258);
nor U22879 (N_22879,N_22059,N_22229);
or U22880 (N_22880,N_22172,N_22437);
or U22881 (N_22881,N_22105,N_22223);
and U22882 (N_22882,N_22145,N_22282);
and U22883 (N_22883,N_22017,N_22193);
xnor U22884 (N_22884,N_22098,N_22342);
or U22885 (N_22885,N_22386,N_22495);
nor U22886 (N_22886,N_22285,N_22363);
xor U22887 (N_22887,N_22477,N_22290);
and U22888 (N_22888,N_22121,N_22021);
xor U22889 (N_22889,N_22199,N_22269);
or U22890 (N_22890,N_22118,N_22269);
nor U22891 (N_22891,N_22048,N_22018);
nor U22892 (N_22892,N_22107,N_22014);
nor U22893 (N_22893,N_22457,N_22007);
nor U22894 (N_22894,N_22133,N_22242);
or U22895 (N_22895,N_22404,N_22189);
nand U22896 (N_22896,N_22033,N_22339);
xor U22897 (N_22897,N_22036,N_22453);
and U22898 (N_22898,N_22198,N_22169);
nor U22899 (N_22899,N_22364,N_22149);
and U22900 (N_22900,N_22009,N_22314);
nand U22901 (N_22901,N_22230,N_22424);
or U22902 (N_22902,N_22088,N_22285);
nor U22903 (N_22903,N_22339,N_22352);
nor U22904 (N_22904,N_22118,N_22493);
nor U22905 (N_22905,N_22424,N_22051);
nor U22906 (N_22906,N_22109,N_22440);
or U22907 (N_22907,N_22316,N_22435);
nand U22908 (N_22908,N_22105,N_22279);
nand U22909 (N_22909,N_22068,N_22305);
xnor U22910 (N_22910,N_22133,N_22478);
or U22911 (N_22911,N_22424,N_22280);
nor U22912 (N_22912,N_22057,N_22426);
nor U22913 (N_22913,N_22391,N_22121);
xor U22914 (N_22914,N_22205,N_22323);
nand U22915 (N_22915,N_22029,N_22155);
nand U22916 (N_22916,N_22121,N_22046);
or U22917 (N_22917,N_22034,N_22102);
xor U22918 (N_22918,N_22060,N_22087);
nand U22919 (N_22919,N_22228,N_22199);
and U22920 (N_22920,N_22049,N_22389);
xnor U22921 (N_22921,N_22385,N_22017);
nand U22922 (N_22922,N_22457,N_22104);
and U22923 (N_22923,N_22011,N_22414);
nand U22924 (N_22924,N_22116,N_22291);
and U22925 (N_22925,N_22092,N_22044);
nor U22926 (N_22926,N_22424,N_22090);
nor U22927 (N_22927,N_22324,N_22344);
or U22928 (N_22928,N_22157,N_22427);
or U22929 (N_22929,N_22332,N_22325);
nor U22930 (N_22930,N_22132,N_22498);
xor U22931 (N_22931,N_22371,N_22380);
or U22932 (N_22932,N_22295,N_22070);
or U22933 (N_22933,N_22363,N_22147);
and U22934 (N_22934,N_22224,N_22119);
xor U22935 (N_22935,N_22382,N_22001);
nor U22936 (N_22936,N_22199,N_22224);
nand U22937 (N_22937,N_22400,N_22265);
nor U22938 (N_22938,N_22030,N_22475);
nand U22939 (N_22939,N_22343,N_22357);
and U22940 (N_22940,N_22177,N_22237);
nand U22941 (N_22941,N_22419,N_22250);
nand U22942 (N_22942,N_22323,N_22139);
or U22943 (N_22943,N_22103,N_22164);
or U22944 (N_22944,N_22466,N_22222);
or U22945 (N_22945,N_22334,N_22293);
xnor U22946 (N_22946,N_22450,N_22213);
xnor U22947 (N_22947,N_22032,N_22357);
nor U22948 (N_22948,N_22101,N_22189);
nand U22949 (N_22949,N_22323,N_22121);
nand U22950 (N_22950,N_22488,N_22107);
or U22951 (N_22951,N_22142,N_22487);
nor U22952 (N_22952,N_22488,N_22497);
or U22953 (N_22953,N_22028,N_22086);
or U22954 (N_22954,N_22119,N_22436);
xor U22955 (N_22955,N_22300,N_22070);
nand U22956 (N_22956,N_22343,N_22308);
nor U22957 (N_22957,N_22039,N_22478);
xnor U22958 (N_22958,N_22387,N_22388);
or U22959 (N_22959,N_22457,N_22061);
and U22960 (N_22960,N_22277,N_22345);
or U22961 (N_22961,N_22066,N_22323);
and U22962 (N_22962,N_22224,N_22138);
nand U22963 (N_22963,N_22008,N_22376);
nand U22964 (N_22964,N_22024,N_22400);
nand U22965 (N_22965,N_22217,N_22457);
xor U22966 (N_22966,N_22208,N_22440);
nor U22967 (N_22967,N_22374,N_22383);
xor U22968 (N_22968,N_22023,N_22117);
nand U22969 (N_22969,N_22354,N_22126);
or U22970 (N_22970,N_22493,N_22186);
xnor U22971 (N_22971,N_22211,N_22453);
xor U22972 (N_22972,N_22120,N_22177);
xor U22973 (N_22973,N_22321,N_22313);
and U22974 (N_22974,N_22346,N_22451);
nor U22975 (N_22975,N_22245,N_22487);
and U22976 (N_22976,N_22130,N_22243);
or U22977 (N_22977,N_22075,N_22273);
or U22978 (N_22978,N_22203,N_22368);
xor U22979 (N_22979,N_22057,N_22479);
nor U22980 (N_22980,N_22413,N_22363);
nor U22981 (N_22981,N_22283,N_22012);
or U22982 (N_22982,N_22279,N_22435);
nor U22983 (N_22983,N_22290,N_22175);
nor U22984 (N_22984,N_22205,N_22277);
or U22985 (N_22985,N_22151,N_22046);
and U22986 (N_22986,N_22187,N_22449);
nand U22987 (N_22987,N_22164,N_22193);
and U22988 (N_22988,N_22427,N_22317);
xor U22989 (N_22989,N_22077,N_22083);
and U22990 (N_22990,N_22478,N_22408);
or U22991 (N_22991,N_22007,N_22470);
and U22992 (N_22992,N_22477,N_22298);
and U22993 (N_22993,N_22328,N_22162);
xor U22994 (N_22994,N_22278,N_22414);
and U22995 (N_22995,N_22362,N_22085);
xor U22996 (N_22996,N_22233,N_22183);
or U22997 (N_22997,N_22415,N_22185);
nor U22998 (N_22998,N_22109,N_22388);
xnor U22999 (N_22999,N_22338,N_22035);
nand U23000 (N_23000,N_22833,N_22881);
xnor U23001 (N_23001,N_22559,N_22836);
and U23002 (N_23002,N_22651,N_22727);
and U23003 (N_23003,N_22840,N_22521);
xnor U23004 (N_23004,N_22854,N_22972);
and U23005 (N_23005,N_22815,N_22907);
nand U23006 (N_23006,N_22762,N_22797);
or U23007 (N_23007,N_22548,N_22844);
or U23008 (N_23008,N_22691,N_22582);
nand U23009 (N_23009,N_22565,N_22978);
nor U23010 (N_23010,N_22624,N_22864);
or U23011 (N_23011,N_22925,N_22641);
and U23012 (N_23012,N_22566,N_22976);
or U23013 (N_23013,N_22540,N_22979);
or U23014 (N_23014,N_22583,N_22749);
nand U23015 (N_23015,N_22576,N_22769);
xnor U23016 (N_23016,N_22534,N_22975);
or U23017 (N_23017,N_22822,N_22658);
nor U23018 (N_23018,N_22577,N_22929);
and U23019 (N_23019,N_22814,N_22660);
or U23020 (N_23020,N_22984,N_22717);
and U23021 (N_23021,N_22832,N_22595);
and U23022 (N_23022,N_22747,N_22688);
or U23023 (N_23023,N_22613,N_22952);
and U23024 (N_23024,N_22838,N_22849);
nand U23025 (N_23025,N_22689,N_22648);
nor U23026 (N_23026,N_22945,N_22914);
or U23027 (N_23027,N_22805,N_22752);
or U23028 (N_23028,N_22897,N_22650);
or U23029 (N_23029,N_22842,N_22807);
or U23030 (N_23030,N_22821,N_22639);
and U23031 (N_23031,N_22537,N_22712);
nor U23032 (N_23032,N_22923,N_22708);
nor U23033 (N_23033,N_22709,N_22685);
or U23034 (N_23034,N_22529,N_22845);
nand U23035 (N_23035,N_22726,N_22678);
and U23036 (N_23036,N_22516,N_22578);
nor U23037 (N_23037,N_22900,N_22987);
nand U23038 (N_23038,N_22974,N_22718);
nand U23039 (N_23039,N_22948,N_22526);
xor U23040 (N_23040,N_22629,N_22930);
xnor U23041 (N_23041,N_22954,N_22783);
xor U23042 (N_23042,N_22596,N_22612);
and U23043 (N_23043,N_22883,N_22561);
nor U23044 (N_23044,N_22563,N_22922);
or U23045 (N_23045,N_22674,N_22887);
and U23046 (N_23046,N_22643,N_22620);
nand U23047 (N_23047,N_22818,N_22743);
and U23048 (N_23048,N_22611,N_22502);
nor U23049 (N_23049,N_22697,N_22757);
and U23050 (N_23050,N_22763,N_22637);
nor U23051 (N_23051,N_22847,N_22985);
nand U23052 (N_23052,N_22915,N_22720);
xnor U23053 (N_23053,N_22823,N_22667);
nand U23054 (N_23054,N_22879,N_22765);
and U23055 (N_23055,N_22852,N_22776);
nand U23056 (N_23056,N_22575,N_22947);
xnor U23057 (N_23057,N_22848,N_22995);
xor U23058 (N_23058,N_22969,N_22895);
and U23059 (N_23059,N_22638,N_22524);
nor U23060 (N_23060,N_22920,N_22971);
or U23061 (N_23061,N_22535,N_22692);
or U23062 (N_23062,N_22801,N_22562);
nor U23063 (N_23063,N_22991,N_22675);
xnor U23064 (N_23064,N_22507,N_22905);
nand U23065 (N_23065,N_22817,N_22919);
xnor U23066 (N_23066,N_22508,N_22775);
xor U23067 (N_23067,N_22878,N_22835);
xor U23068 (N_23068,N_22735,N_22795);
nor U23069 (N_23069,N_22820,N_22789);
or U23070 (N_23070,N_22786,N_22874);
xnor U23071 (N_23071,N_22531,N_22656);
nor U23072 (N_23072,N_22500,N_22800);
or U23073 (N_23073,N_22545,N_22996);
nor U23074 (N_23074,N_22664,N_22606);
xor U23075 (N_23075,N_22501,N_22690);
nand U23076 (N_23076,N_22777,N_22773);
nor U23077 (N_23077,N_22544,N_22604);
and U23078 (N_23078,N_22716,N_22600);
or U23079 (N_23079,N_22748,N_22630);
and U23080 (N_23080,N_22659,N_22702);
and U23081 (N_23081,N_22610,N_22779);
or U23082 (N_23082,N_22937,N_22888);
or U23083 (N_23083,N_22810,N_22877);
nor U23084 (N_23084,N_22599,N_22868);
and U23085 (N_23085,N_22580,N_22568);
or U23086 (N_23086,N_22686,N_22645);
nand U23087 (N_23087,N_22569,N_22994);
nand U23088 (N_23088,N_22703,N_22760);
nor U23089 (N_23089,N_22839,N_22533);
or U23090 (N_23090,N_22867,N_22944);
or U23091 (N_23091,N_22661,N_22764);
xor U23092 (N_23092,N_22593,N_22999);
or U23093 (N_23093,N_22572,N_22943);
or U23094 (N_23094,N_22668,N_22767);
and U23095 (N_23095,N_22632,N_22935);
nor U23096 (N_23096,N_22819,N_22701);
nor U23097 (N_23097,N_22858,N_22706);
or U23098 (N_23098,N_22546,N_22998);
xor U23099 (N_23099,N_22594,N_22636);
xnor U23100 (N_23100,N_22557,N_22970);
and U23101 (N_23101,N_22621,N_22758);
nand U23102 (N_23102,N_22704,N_22790);
nand U23103 (N_23103,N_22737,N_22680);
or U23104 (N_23104,N_22555,N_22542);
or U23105 (N_23105,N_22591,N_22654);
nand U23106 (N_23106,N_22761,N_22850);
xor U23107 (N_23107,N_22513,N_22913);
nor U23108 (N_23108,N_22855,N_22541);
nand U23109 (N_23109,N_22928,N_22870);
xnor U23110 (N_23110,N_22901,N_22753);
xnor U23111 (N_23111,N_22579,N_22552);
and U23112 (N_23112,N_22927,N_22687);
nand U23113 (N_23113,N_22707,N_22585);
xnor U23114 (N_23114,N_22738,N_22791);
nor U23115 (N_23115,N_22977,N_22967);
nor U23116 (N_23116,N_22917,N_22682);
nor U23117 (N_23117,N_22861,N_22644);
nand U23118 (N_23118,N_22571,N_22902);
nor U23119 (N_23119,N_22560,N_22556);
nor U23120 (N_23120,N_22955,N_22856);
xnor U23121 (N_23121,N_22742,N_22505);
xnor U23122 (N_23122,N_22514,N_22581);
nor U23123 (N_23123,N_22906,N_22730);
nor U23124 (N_23124,N_22898,N_22676);
xnor U23125 (N_23125,N_22677,N_22517);
and U23126 (N_23126,N_22802,N_22695);
and U23127 (N_23127,N_22951,N_22640);
and U23128 (N_23128,N_22882,N_22592);
nor U23129 (N_23129,N_22587,N_22550);
nand U23130 (N_23130,N_22586,N_22705);
and U23131 (N_23131,N_22798,N_22916);
or U23132 (N_23132,N_22744,N_22780);
xnor U23133 (N_23133,N_22741,N_22506);
or U23134 (N_23134,N_22736,N_22788);
nand U23135 (N_23135,N_22518,N_22733);
xor U23136 (N_23136,N_22627,N_22869);
xnor U23137 (N_23137,N_22792,N_22921);
nor U23138 (N_23138,N_22710,N_22723);
or U23139 (N_23139,N_22511,N_22778);
nand U23140 (N_23140,N_22931,N_22891);
and U23141 (N_23141,N_22831,N_22631);
and U23142 (N_23142,N_22816,N_22665);
xor U23143 (N_23143,N_22597,N_22886);
nor U23144 (N_23144,N_22826,N_22957);
or U23145 (N_23145,N_22616,N_22766);
or U23146 (N_23146,N_22655,N_22993);
and U23147 (N_23147,N_22598,N_22809);
and U23148 (N_23148,N_22522,N_22918);
nor U23149 (N_23149,N_22670,N_22950);
nor U23150 (N_23150,N_22772,N_22669);
nor U23151 (N_23151,N_22890,N_22997);
and U23152 (N_23152,N_22862,N_22963);
xnor U23153 (N_23153,N_22846,N_22553);
and U23154 (N_23154,N_22527,N_22990);
nand U23155 (N_23155,N_22756,N_22543);
or U23156 (N_23156,N_22635,N_22625);
xnor U23157 (N_23157,N_22924,N_22731);
xnor U23158 (N_23158,N_22770,N_22681);
nor U23159 (N_23159,N_22796,N_22829);
xor U23160 (N_23160,N_22892,N_22893);
nand U23161 (N_23161,N_22649,N_22983);
and U23162 (N_23162,N_22503,N_22806);
xor U23163 (N_23163,N_22872,N_22768);
nor U23164 (N_23164,N_22729,N_22671);
xnor U23165 (N_23165,N_22605,N_22549);
and U23166 (N_23166,N_22837,N_22713);
xor U23167 (N_23167,N_22590,N_22618);
nand U23168 (N_23168,N_22968,N_22841);
or U23169 (N_23169,N_22700,N_22693);
and U23170 (N_23170,N_22714,N_22628);
and U23171 (N_23171,N_22719,N_22982);
and U23172 (N_23172,N_22732,N_22721);
nand U23173 (N_23173,N_22759,N_22853);
xnor U23174 (N_23174,N_22932,N_22804);
nand U23175 (N_23175,N_22986,N_22940);
nor U23176 (N_23176,N_22647,N_22679);
xor U23177 (N_23177,N_22751,N_22958);
xnor U23178 (N_23178,N_22603,N_22964);
and U23179 (N_23179,N_22953,N_22532);
nand U23180 (N_23180,N_22812,N_22966);
or U23181 (N_23181,N_22782,N_22828);
nand U23182 (N_23182,N_22910,N_22754);
and U23183 (N_23183,N_22683,N_22699);
or U23184 (N_23184,N_22904,N_22539);
nand U23185 (N_23185,N_22811,N_22623);
or U23186 (N_23186,N_22684,N_22504);
nor U23187 (N_23187,N_22573,N_22851);
nand U23188 (N_23188,N_22739,N_22755);
or U23189 (N_23189,N_22673,N_22885);
xnor U23190 (N_23190,N_22512,N_22908);
xnor U23191 (N_23191,N_22525,N_22871);
nand U23192 (N_23192,N_22934,N_22634);
nand U23193 (N_23193,N_22528,N_22936);
xor U23194 (N_23194,N_22750,N_22989);
nor U23195 (N_23195,N_22551,N_22912);
and U23196 (N_23196,N_22567,N_22992);
nand U23197 (N_23197,N_22911,N_22946);
nor U23198 (N_23198,N_22961,N_22515);
xnor U23199 (N_23199,N_22574,N_22509);
and U23200 (N_23200,N_22745,N_22857);
and U23201 (N_23201,N_22715,N_22698);
or U23202 (N_23202,N_22523,N_22781);
nor U23203 (N_23203,N_22926,N_22909);
or U23204 (N_23204,N_22564,N_22949);
or U23205 (N_23205,N_22799,N_22663);
nor U23206 (N_23206,N_22941,N_22547);
or U23207 (N_23207,N_22884,N_22962);
nand U23208 (N_23208,N_22602,N_22642);
and U23209 (N_23209,N_22558,N_22834);
nor U23210 (N_23210,N_22740,N_22771);
xor U23211 (N_23211,N_22813,N_22875);
and U23212 (N_23212,N_22725,N_22903);
xor U23213 (N_23213,N_22666,N_22960);
and U23214 (N_23214,N_22633,N_22601);
and U23215 (N_23215,N_22942,N_22859);
nor U23216 (N_23216,N_22711,N_22787);
nand U23217 (N_23217,N_22728,N_22785);
xor U23218 (N_23218,N_22825,N_22863);
and U23219 (N_23219,N_22734,N_22824);
xor U23220 (N_23220,N_22784,N_22959);
xor U23221 (N_23221,N_22866,N_22510);
xnor U23222 (N_23222,N_22696,N_22617);
nand U23223 (N_23223,N_22589,N_22774);
and U23224 (N_23224,N_22880,N_22536);
and U23225 (N_23225,N_22746,N_22722);
nand U23226 (N_23226,N_22619,N_22981);
nand U23227 (N_23227,N_22793,N_22894);
nor U23228 (N_23228,N_22808,N_22873);
and U23229 (N_23229,N_22843,N_22584);
nor U23230 (N_23230,N_22554,N_22652);
nor U23231 (N_23231,N_22794,N_22520);
and U23232 (N_23232,N_22876,N_22988);
and U23233 (N_23233,N_22939,N_22538);
and U23234 (N_23234,N_22646,N_22607);
xor U23235 (N_23235,N_22896,N_22662);
xor U23236 (N_23236,N_22827,N_22519);
and U23237 (N_23237,N_22889,N_22803);
and U23238 (N_23238,N_22626,N_22614);
or U23239 (N_23239,N_22588,N_22653);
or U23240 (N_23240,N_22980,N_22830);
and U23241 (N_23241,N_22933,N_22965);
nor U23242 (N_23242,N_22609,N_22608);
xor U23243 (N_23243,N_22657,N_22860);
and U23244 (N_23244,N_22622,N_22938);
xor U23245 (N_23245,N_22899,N_22973);
or U23246 (N_23246,N_22956,N_22615);
or U23247 (N_23247,N_22570,N_22724);
or U23248 (N_23248,N_22672,N_22530);
nand U23249 (N_23249,N_22694,N_22865);
nand U23250 (N_23250,N_22592,N_22775);
and U23251 (N_23251,N_22702,N_22716);
or U23252 (N_23252,N_22745,N_22889);
and U23253 (N_23253,N_22670,N_22857);
nand U23254 (N_23254,N_22998,N_22502);
nand U23255 (N_23255,N_22947,N_22527);
nand U23256 (N_23256,N_22536,N_22963);
xor U23257 (N_23257,N_22886,N_22838);
nor U23258 (N_23258,N_22751,N_22703);
nor U23259 (N_23259,N_22724,N_22667);
xnor U23260 (N_23260,N_22943,N_22533);
nor U23261 (N_23261,N_22628,N_22655);
nor U23262 (N_23262,N_22687,N_22813);
or U23263 (N_23263,N_22791,N_22804);
or U23264 (N_23264,N_22800,N_22614);
nor U23265 (N_23265,N_22581,N_22529);
nand U23266 (N_23266,N_22625,N_22505);
nor U23267 (N_23267,N_22862,N_22911);
and U23268 (N_23268,N_22645,N_22921);
nand U23269 (N_23269,N_22540,N_22869);
or U23270 (N_23270,N_22564,N_22542);
or U23271 (N_23271,N_22639,N_22609);
xor U23272 (N_23272,N_22953,N_22607);
xnor U23273 (N_23273,N_22898,N_22572);
xnor U23274 (N_23274,N_22585,N_22850);
or U23275 (N_23275,N_22617,N_22597);
nand U23276 (N_23276,N_22665,N_22906);
nand U23277 (N_23277,N_22917,N_22753);
and U23278 (N_23278,N_22932,N_22808);
nor U23279 (N_23279,N_22947,N_22584);
and U23280 (N_23280,N_22566,N_22798);
xnor U23281 (N_23281,N_22937,N_22981);
or U23282 (N_23282,N_22826,N_22945);
nor U23283 (N_23283,N_22833,N_22669);
nand U23284 (N_23284,N_22607,N_22832);
nor U23285 (N_23285,N_22730,N_22779);
nor U23286 (N_23286,N_22983,N_22640);
or U23287 (N_23287,N_22987,N_22723);
nor U23288 (N_23288,N_22620,N_22813);
or U23289 (N_23289,N_22886,N_22981);
and U23290 (N_23290,N_22728,N_22717);
xnor U23291 (N_23291,N_22704,N_22878);
and U23292 (N_23292,N_22790,N_22871);
xor U23293 (N_23293,N_22851,N_22613);
xor U23294 (N_23294,N_22683,N_22701);
nand U23295 (N_23295,N_22555,N_22651);
xor U23296 (N_23296,N_22693,N_22788);
and U23297 (N_23297,N_22953,N_22741);
and U23298 (N_23298,N_22545,N_22515);
and U23299 (N_23299,N_22926,N_22907);
nand U23300 (N_23300,N_22521,N_22559);
nand U23301 (N_23301,N_22901,N_22953);
xnor U23302 (N_23302,N_22850,N_22994);
and U23303 (N_23303,N_22804,N_22969);
or U23304 (N_23304,N_22625,N_22797);
and U23305 (N_23305,N_22669,N_22797);
and U23306 (N_23306,N_22963,N_22864);
nor U23307 (N_23307,N_22600,N_22804);
or U23308 (N_23308,N_22569,N_22508);
nand U23309 (N_23309,N_22918,N_22779);
nand U23310 (N_23310,N_22845,N_22824);
and U23311 (N_23311,N_22665,N_22799);
xor U23312 (N_23312,N_22524,N_22751);
and U23313 (N_23313,N_22954,N_22626);
xnor U23314 (N_23314,N_22731,N_22551);
xnor U23315 (N_23315,N_22950,N_22873);
and U23316 (N_23316,N_22604,N_22805);
or U23317 (N_23317,N_22730,N_22733);
and U23318 (N_23318,N_22679,N_22916);
nand U23319 (N_23319,N_22992,N_22674);
or U23320 (N_23320,N_22543,N_22571);
nand U23321 (N_23321,N_22815,N_22995);
and U23322 (N_23322,N_22590,N_22935);
nor U23323 (N_23323,N_22561,N_22623);
nand U23324 (N_23324,N_22973,N_22965);
xor U23325 (N_23325,N_22623,N_22711);
or U23326 (N_23326,N_22807,N_22865);
nand U23327 (N_23327,N_22897,N_22560);
or U23328 (N_23328,N_22803,N_22983);
xor U23329 (N_23329,N_22989,N_22909);
nand U23330 (N_23330,N_22847,N_22575);
and U23331 (N_23331,N_22508,N_22825);
and U23332 (N_23332,N_22585,N_22794);
nor U23333 (N_23333,N_22990,N_22515);
or U23334 (N_23334,N_22605,N_22983);
nand U23335 (N_23335,N_22619,N_22860);
nand U23336 (N_23336,N_22894,N_22788);
nor U23337 (N_23337,N_22731,N_22623);
nor U23338 (N_23338,N_22679,N_22817);
nor U23339 (N_23339,N_22528,N_22586);
and U23340 (N_23340,N_22739,N_22848);
nor U23341 (N_23341,N_22800,N_22978);
and U23342 (N_23342,N_22730,N_22670);
nor U23343 (N_23343,N_22758,N_22662);
and U23344 (N_23344,N_22997,N_22967);
or U23345 (N_23345,N_22753,N_22996);
nand U23346 (N_23346,N_22658,N_22881);
or U23347 (N_23347,N_22961,N_22687);
xnor U23348 (N_23348,N_22848,N_22558);
nand U23349 (N_23349,N_22662,N_22716);
and U23350 (N_23350,N_22713,N_22527);
xnor U23351 (N_23351,N_22844,N_22713);
or U23352 (N_23352,N_22594,N_22886);
xnor U23353 (N_23353,N_22513,N_22757);
and U23354 (N_23354,N_22850,N_22931);
nor U23355 (N_23355,N_22533,N_22671);
nor U23356 (N_23356,N_22988,N_22804);
and U23357 (N_23357,N_22684,N_22669);
nor U23358 (N_23358,N_22913,N_22848);
and U23359 (N_23359,N_22802,N_22883);
nor U23360 (N_23360,N_22653,N_22570);
and U23361 (N_23361,N_22932,N_22906);
nor U23362 (N_23362,N_22555,N_22863);
nand U23363 (N_23363,N_22999,N_22939);
nor U23364 (N_23364,N_22963,N_22717);
and U23365 (N_23365,N_22797,N_22664);
nor U23366 (N_23366,N_22863,N_22923);
nor U23367 (N_23367,N_22566,N_22504);
nand U23368 (N_23368,N_22567,N_22727);
or U23369 (N_23369,N_22512,N_22547);
nand U23370 (N_23370,N_22517,N_22973);
nor U23371 (N_23371,N_22642,N_22693);
nand U23372 (N_23372,N_22567,N_22833);
nand U23373 (N_23373,N_22733,N_22909);
xor U23374 (N_23374,N_22885,N_22911);
nor U23375 (N_23375,N_22576,N_22808);
nand U23376 (N_23376,N_22633,N_22550);
xnor U23377 (N_23377,N_22831,N_22774);
and U23378 (N_23378,N_22612,N_22923);
nand U23379 (N_23379,N_22672,N_22876);
nand U23380 (N_23380,N_22511,N_22580);
xnor U23381 (N_23381,N_22737,N_22793);
nand U23382 (N_23382,N_22871,N_22589);
nand U23383 (N_23383,N_22657,N_22786);
or U23384 (N_23384,N_22641,N_22718);
xor U23385 (N_23385,N_22833,N_22999);
xnor U23386 (N_23386,N_22890,N_22751);
nand U23387 (N_23387,N_22892,N_22939);
and U23388 (N_23388,N_22518,N_22756);
nand U23389 (N_23389,N_22559,N_22872);
xnor U23390 (N_23390,N_22584,N_22769);
nor U23391 (N_23391,N_22784,N_22700);
nand U23392 (N_23392,N_22910,N_22840);
or U23393 (N_23393,N_22922,N_22501);
or U23394 (N_23394,N_22873,N_22944);
xnor U23395 (N_23395,N_22724,N_22980);
nor U23396 (N_23396,N_22959,N_22797);
and U23397 (N_23397,N_22784,N_22738);
nand U23398 (N_23398,N_22614,N_22633);
nor U23399 (N_23399,N_22960,N_22829);
nor U23400 (N_23400,N_22862,N_22723);
nor U23401 (N_23401,N_22698,N_22610);
and U23402 (N_23402,N_22866,N_22938);
xor U23403 (N_23403,N_22702,N_22867);
and U23404 (N_23404,N_22862,N_22733);
and U23405 (N_23405,N_22983,N_22912);
nor U23406 (N_23406,N_22915,N_22775);
or U23407 (N_23407,N_22586,N_22745);
xnor U23408 (N_23408,N_22797,N_22910);
nand U23409 (N_23409,N_22782,N_22643);
nand U23410 (N_23410,N_22554,N_22847);
nor U23411 (N_23411,N_22834,N_22827);
nor U23412 (N_23412,N_22761,N_22806);
and U23413 (N_23413,N_22824,N_22922);
nor U23414 (N_23414,N_22845,N_22770);
nor U23415 (N_23415,N_22628,N_22807);
xnor U23416 (N_23416,N_22996,N_22540);
and U23417 (N_23417,N_22791,N_22616);
and U23418 (N_23418,N_22983,N_22886);
or U23419 (N_23419,N_22512,N_22979);
or U23420 (N_23420,N_22563,N_22577);
nor U23421 (N_23421,N_22544,N_22657);
nand U23422 (N_23422,N_22935,N_22682);
nor U23423 (N_23423,N_22988,N_22894);
and U23424 (N_23424,N_22590,N_22811);
nand U23425 (N_23425,N_22956,N_22716);
or U23426 (N_23426,N_22617,N_22549);
nand U23427 (N_23427,N_22736,N_22608);
and U23428 (N_23428,N_22525,N_22588);
or U23429 (N_23429,N_22528,N_22631);
xnor U23430 (N_23430,N_22619,N_22844);
xor U23431 (N_23431,N_22855,N_22934);
or U23432 (N_23432,N_22720,N_22711);
or U23433 (N_23433,N_22739,N_22808);
and U23434 (N_23434,N_22589,N_22916);
or U23435 (N_23435,N_22809,N_22652);
or U23436 (N_23436,N_22912,N_22659);
and U23437 (N_23437,N_22788,N_22782);
or U23438 (N_23438,N_22616,N_22500);
nor U23439 (N_23439,N_22663,N_22766);
nand U23440 (N_23440,N_22577,N_22777);
xnor U23441 (N_23441,N_22688,N_22810);
xnor U23442 (N_23442,N_22536,N_22528);
xor U23443 (N_23443,N_22905,N_22720);
xor U23444 (N_23444,N_22891,N_22790);
or U23445 (N_23445,N_22502,N_22883);
nor U23446 (N_23446,N_22692,N_22931);
xnor U23447 (N_23447,N_22797,N_22761);
nor U23448 (N_23448,N_22681,N_22902);
nor U23449 (N_23449,N_22647,N_22859);
xor U23450 (N_23450,N_22596,N_22892);
and U23451 (N_23451,N_22826,N_22886);
nand U23452 (N_23452,N_22782,N_22762);
or U23453 (N_23453,N_22976,N_22860);
xnor U23454 (N_23454,N_22543,N_22819);
and U23455 (N_23455,N_22885,N_22901);
nand U23456 (N_23456,N_22655,N_22566);
xnor U23457 (N_23457,N_22618,N_22611);
xor U23458 (N_23458,N_22557,N_22502);
and U23459 (N_23459,N_22872,N_22814);
nor U23460 (N_23460,N_22579,N_22632);
and U23461 (N_23461,N_22826,N_22879);
nor U23462 (N_23462,N_22671,N_22844);
and U23463 (N_23463,N_22878,N_22913);
xor U23464 (N_23464,N_22682,N_22817);
or U23465 (N_23465,N_22998,N_22723);
nand U23466 (N_23466,N_22639,N_22587);
nor U23467 (N_23467,N_22730,N_22942);
and U23468 (N_23468,N_22811,N_22537);
xnor U23469 (N_23469,N_22836,N_22992);
nor U23470 (N_23470,N_22782,N_22723);
nand U23471 (N_23471,N_22989,N_22937);
or U23472 (N_23472,N_22877,N_22558);
or U23473 (N_23473,N_22787,N_22608);
or U23474 (N_23474,N_22683,N_22573);
nor U23475 (N_23475,N_22828,N_22661);
xor U23476 (N_23476,N_22784,N_22561);
or U23477 (N_23477,N_22640,N_22879);
nand U23478 (N_23478,N_22582,N_22696);
xnor U23479 (N_23479,N_22506,N_22929);
nor U23480 (N_23480,N_22966,N_22768);
and U23481 (N_23481,N_22510,N_22541);
and U23482 (N_23482,N_22709,N_22554);
xor U23483 (N_23483,N_22779,N_22543);
nand U23484 (N_23484,N_22628,N_22506);
or U23485 (N_23485,N_22940,N_22893);
nand U23486 (N_23486,N_22966,N_22561);
xnor U23487 (N_23487,N_22602,N_22575);
and U23488 (N_23488,N_22755,N_22798);
and U23489 (N_23489,N_22929,N_22999);
nand U23490 (N_23490,N_22616,N_22765);
or U23491 (N_23491,N_22938,N_22503);
xor U23492 (N_23492,N_22972,N_22524);
nor U23493 (N_23493,N_22900,N_22849);
nor U23494 (N_23494,N_22994,N_22966);
xnor U23495 (N_23495,N_22784,N_22590);
nor U23496 (N_23496,N_22894,N_22720);
nand U23497 (N_23497,N_22797,N_22702);
nand U23498 (N_23498,N_22590,N_22658);
nand U23499 (N_23499,N_22840,N_22659);
or U23500 (N_23500,N_23272,N_23279);
nand U23501 (N_23501,N_23163,N_23074);
or U23502 (N_23502,N_23248,N_23099);
and U23503 (N_23503,N_23239,N_23066);
nor U23504 (N_23504,N_23393,N_23377);
or U23505 (N_23505,N_23112,N_23422);
xnor U23506 (N_23506,N_23498,N_23294);
xor U23507 (N_23507,N_23165,N_23494);
nor U23508 (N_23508,N_23076,N_23020);
and U23509 (N_23509,N_23042,N_23173);
xor U23510 (N_23510,N_23113,N_23499);
xor U23511 (N_23511,N_23282,N_23087);
xnor U23512 (N_23512,N_23206,N_23417);
or U23513 (N_23513,N_23055,N_23432);
nand U23514 (N_23514,N_23465,N_23453);
nor U23515 (N_23515,N_23410,N_23375);
or U23516 (N_23516,N_23396,N_23149);
or U23517 (N_23517,N_23265,N_23164);
nor U23518 (N_23518,N_23230,N_23110);
xor U23519 (N_23519,N_23335,N_23053);
nor U23520 (N_23520,N_23235,N_23362);
or U23521 (N_23521,N_23078,N_23211);
and U23522 (N_23522,N_23072,N_23109);
nand U23523 (N_23523,N_23260,N_23405);
nand U23524 (N_23524,N_23415,N_23243);
or U23525 (N_23525,N_23141,N_23142);
and U23526 (N_23526,N_23025,N_23010);
or U23527 (N_23527,N_23478,N_23322);
nor U23528 (N_23528,N_23296,N_23463);
nand U23529 (N_23529,N_23314,N_23472);
and U23530 (N_23530,N_23287,N_23372);
nand U23531 (N_23531,N_23263,N_23481);
xor U23532 (N_23532,N_23218,N_23430);
nand U23533 (N_23533,N_23217,N_23283);
xnor U23534 (N_23534,N_23166,N_23345);
nor U23535 (N_23535,N_23212,N_23070);
nand U23536 (N_23536,N_23075,N_23379);
nand U23537 (N_23537,N_23444,N_23101);
xor U23538 (N_23538,N_23416,N_23147);
nor U23539 (N_23539,N_23355,N_23056);
nand U23540 (N_23540,N_23023,N_23100);
xnor U23541 (N_23541,N_23452,N_23464);
xnor U23542 (N_23542,N_23445,N_23057);
nand U23543 (N_23543,N_23306,N_23016);
nor U23544 (N_23544,N_23352,N_23387);
nand U23545 (N_23545,N_23493,N_23441);
or U23546 (N_23546,N_23238,N_23450);
and U23547 (N_23547,N_23143,N_23374);
nand U23548 (N_23548,N_23304,N_23367);
nor U23549 (N_23549,N_23346,N_23083);
or U23550 (N_23550,N_23333,N_23246);
and U23551 (N_23551,N_23161,N_23037);
and U23552 (N_23552,N_23199,N_23407);
nor U23553 (N_23553,N_23006,N_23220);
nand U23554 (N_23554,N_23122,N_23266);
xnor U23555 (N_23555,N_23026,N_23431);
or U23556 (N_23556,N_23135,N_23390);
xnor U23557 (N_23557,N_23124,N_23286);
nor U23558 (N_23558,N_23492,N_23085);
nand U23559 (N_23559,N_23082,N_23244);
nor U23560 (N_23560,N_23240,N_23301);
or U23561 (N_23561,N_23414,N_23205);
or U23562 (N_23562,N_23348,N_23029);
xnor U23563 (N_23563,N_23257,N_23326);
nor U23564 (N_23564,N_23136,N_23221);
and U23565 (N_23565,N_23412,N_23419);
and U23566 (N_23566,N_23245,N_23151);
and U23567 (N_23567,N_23247,N_23292);
nand U23568 (N_23568,N_23406,N_23285);
or U23569 (N_23569,N_23328,N_23090);
nor U23570 (N_23570,N_23378,N_23293);
or U23571 (N_23571,N_23490,N_23486);
nor U23572 (N_23572,N_23137,N_23261);
nor U23573 (N_23573,N_23232,N_23035);
nand U23574 (N_23574,N_23096,N_23125);
nand U23575 (N_23575,N_23024,N_23021);
and U23576 (N_23576,N_23373,N_23106);
or U23577 (N_23577,N_23357,N_23114);
or U23578 (N_23578,N_23187,N_23005);
xor U23579 (N_23579,N_23309,N_23330);
nor U23580 (N_23580,N_23116,N_23288);
nand U23581 (N_23581,N_23302,N_23281);
nand U23582 (N_23582,N_23267,N_23289);
and U23583 (N_23583,N_23475,N_23466);
nor U23584 (N_23584,N_23229,N_23204);
or U23585 (N_23585,N_23256,N_23000);
xor U23586 (N_23586,N_23155,N_23157);
or U23587 (N_23587,N_23371,N_23473);
nor U23588 (N_23588,N_23086,N_23191);
xor U23589 (N_23589,N_23284,N_23300);
and U23590 (N_23590,N_23434,N_23435);
or U23591 (N_23591,N_23456,N_23255);
nand U23592 (N_23592,N_23403,N_23159);
xor U23593 (N_23593,N_23258,N_23144);
nor U23594 (N_23594,N_23047,N_23438);
nand U23595 (N_23595,N_23389,N_23369);
or U23596 (N_23596,N_23059,N_23012);
xnor U23597 (N_23597,N_23420,N_23226);
nand U23598 (N_23598,N_23034,N_23234);
xnor U23599 (N_23599,N_23172,N_23017);
nand U23600 (N_23600,N_23152,N_23111);
xor U23601 (N_23601,N_23118,N_23095);
or U23602 (N_23602,N_23311,N_23168);
and U23603 (N_23603,N_23084,N_23320);
xor U23604 (N_23604,N_23052,N_23158);
nand U23605 (N_23605,N_23477,N_23397);
xor U23606 (N_23606,N_23426,N_23337);
and U23607 (N_23607,N_23359,N_23327);
xnor U23608 (N_23608,N_23252,N_23041);
nand U23609 (N_23609,N_23196,N_23303);
nand U23610 (N_23610,N_23033,N_23081);
nand U23611 (N_23611,N_23358,N_23398);
and U23612 (N_23612,N_23364,N_23439);
or U23613 (N_23613,N_23079,N_23065);
nor U23614 (N_23614,N_23479,N_23262);
nand U23615 (N_23615,N_23154,N_23175);
or U23616 (N_23616,N_23485,N_23411);
and U23617 (N_23617,N_23132,N_23380);
xnor U23618 (N_23618,N_23331,N_23278);
nand U23619 (N_23619,N_23323,N_23190);
and U23620 (N_23620,N_23071,N_23058);
xor U23621 (N_23621,N_23421,N_23496);
and U23622 (N_23622,N_23186,N_23051);
nor U23623 (N_23623,N_23324,N_23436);
nor U23624 (N_23624,N_23241,N_23148);
or U23625 (N_23625,N_23145,N_23370);
and U23626 (N_23626,N_23134,N_23340);
or U23627 (N_23627,N_23044,N_23332);
nor U23628 (N_23628,N_23117,N_23404);
nand U23629 (N_23629,N_23031,N_23097);
nand U23630 (N_23630,N_23063,N_23138);
nor U23631 (N_23631,N_23350,N_23068);
or U23632 (N_23632,N_23150,N_23022);
and U23633 (N_23633,N_23461,N_23185);
and U23634 (N_23634,N_23448,N_23394);
and U23635 (N_23635,N_23233,N_23127);
or U23636 (N_23636,N_23131,N_23197);
and U23637 (N_23637,N_23179,N_23305);
xnor U23638 (N_23638,N_23356,N_23128);
nand U23639 (N_23639,N_23093,N_23313);
nand U23640 (N_23640,N_23440,N_23334);
and U23641 (N_23641,N_23170,N_23178);
nor U23642 (N_23642,N_23013,N_23329);
xnor U23643 (N_23643,N_23360,N_23318);
xor U23644 (N_23644,N_23400,N_23443);
nand U23645 (N_23645,N_23019,N_23146);
nand U23646 (N_23646,N_23181,N_23160);
nand U23647 (N_23647,N_23073,N_23468);
nor U23648 (N_23648,N_23015,N_23429);
or U23649 (N_23649,N_23080,N_23209);
and U23650 (N_23650,N_23126,N_23325);
xor U23651 (N_23651,N_23480,N_23408);
nor U23652 (N_23652,N_23169,N_23195);
or U23653 (N_23653,N_23268,N_23129);
nor U23654 (N_23654,N_23295,N_23269);
or U23655 (N_23655,N_23385,N_23460);
nor U23656 (N_23656,N_23089,N_23028);
and U23657 (N_23657,N_23382,N_23094);
or U23658 (N_23658,N_23036,N_23476);
and U23659 (N_23659,N_23183,N_23353);
or U23660 (N_23660,N_23088,N_23105);
xnor U23661 (N_23661,N_23216,N_23457);
and U23662 (N_23662,N_23280,N_23275);
or U23663 (N_23663,N_23001,N_23140);
nand U23664 (N_23664,N_23446,N_23038);
or U23665 (N_23665,N_23402,N_23366);
or U23666 (N_23666,N_23315,N_23391);
nand U23667 (N_23667,N_23351,N_23208);
nor U23668 (N_23668,N_23049,N_23227);
or U23669 (N_23669,N_23484,N_23054);
xnor U23670 (N_23670,N_23188,N_23067);
nor U23671 (N_23671,N_23491,N_23384);
nand U23672 (N_23672,N_23317,N_23123);
nand U23673 (N_23673,N_23427,N_23338);
nand U23674 (N_23674,N_23392,N_23399);
and U23675 (N_23675,N_23433,N_23046);
xnor U23676 (N_23676,N_23413,N_23139);
or U23677 (N_23677,N_23189,N_23250);
xor U23678 (N_23678,N_23277,N_23459);
and U23679 (N_23679,N_23039,N_23349);
xor U23680 (N_23680,N_23177,N_23098);
nor U23681 (N_23681,N_23249,N_23455);
xnor U23682 (N_23682,N_23062,N_23254);
xor U23683 (N_23683,N_23027,N_23401);
and U23684 (N_23684,N_23102,N_23447);
or U23685 (N_23685,N_23184,N_23045);
nand U23686 (N_23686,N_23471,N_23061);
or U23687 (N_23687,N_23470,N_23291);
xor U23688 (N_23688,N_23032,N_23210);
nand U23689 (N_23689,N_23043,N_23174);
xor U23690 (N_23690,N_23454,N_23451);
or U23691 (N_23691,N_23307,N_23270);
and U23692 (N_23692,N_23009,N_23368);
nand U23693 (N_23693,N_23194,N_23004);
nor U23694 (N_23694,N_23495,N_23092);
nor U23695 (N_23695,N_23365,N_23231);
and U23696 (N_23696,N_23201,N_23363);
nor U23697 (N_23697,N_23299,N_23060);
or U23698 (N_23698,N_23409,N_23316);
xnor U23699 (N_23699,N_23395,N_23488);
nand U23700 (N_23700,N_23424,N_23215);
nor U23701 (N_23701,N_23467,N_23388);
nand U23702 (N_23702,N_23386,N_23347);
or U23703 (N_23703,N_23180,N_23003);
nor U23704 (N_23704,N_23298,N_23202);
nor U23705 (N_23705,N_23271,N_23156);
xnor U23706 (N_23706,N_23253,N_23171);
and U23707 (N_23707,N_23251,N_23489);
xnor U23708 (N_23708,N_23091,N_23469);
nand U23709 (N_23709,N_23276,N_23119);
nand U23710 (N_23710,N_23236,N_23319);
or U23711 (N_23711,N_23458,N_23418);
and U23712 (N_23712,N_23361,N_23064);
nand U23713 (N_23713,N_23050,N_23048);
and U23714 (N_23714,N_23310,N_23008);
nor U23715 (N_23715,N_23107,N_23462);
nor U23716 (N_23716,N_23040,N_23030);
nor U23717 (N_23717,N_23381,N_23176);
nand U23718 (N_23718,N_23069,N_23222);
xnor U23719 (N_23719,N_23115,N_23290);
xnor U23720 (N_23720,N_23336,N_23297);
xor U23721 (N_23721,N_23214,N_23120);
xnor U23722 (N_23722,N_23449,N_23274);
or U23723 (N_23723,N_23193,N_23228);
or U23724 (N_23724,N_23259,N_23121);
nand U23725 (N_23725,N_23341,N_23482);
and U23726 (N_23726,N_23312,N_23167);
and U23727 (N_23727,N_23014,N_23153);
nand U23728 (N_23728,N_23423,N_23383);
xor U23729 (N_23729,N_23207,N_23497);
or U23730 (N_23730,N_23442,N_23133);
and U23731 (N_23731,N_23225,N_23002);
nand U23732 (N_23732,N_23182,N_23203);
or U23733 (N_23733,N_23428,N_23343);
or U23734 (N_23734,N_23344,N_23339);
xnor U23735 (N_23735,N_23242,N_23103);
nor U23736 (N_23736,N_23223,N_23104);
or U23737 (N_23737,N_23483,N_23273);
or U23738 (N_23738,N_23264,N_23425);
nor U23739 (N_23739,N_23077,N_23200);
nor U23740 (N_23740,N_23487,N_23198);
nor U23741 (N_23741,N_23376,N_23219);
and U23742 (N_23742,N_23018,N_23308);
nand U23743 (N_23743,N_23342,N_23224);
or U23744 (N_23744,N_23007,N_23192);
nand U23745 (N_23745,N_23354,N_23237);
nand U23746 (N_23746,N_23108,N_23437);
xor U23747 (N_23747,N_23213,N_23011);
nand U23748 (N_23748,N_23162,N_23321);
and U23749 (N_23749,N_23130,N_23474);
and U23750 (N_23750,N_23184,N_23180);
xor U23751 (N_23751,N_23036,N_23351);
or U23752 (N_23752,N_23224,N_23474);
or U23753 (N_23753,N_23125,N_23034);
nor U23754 (N_23754,N_23388,N_23271);
or U23755 (N_23755,N_23352,N_23128);
or U23756 (N_23756,N_23309,N_23233);
or U23757 (N_23757,N_23228,N_23024);
and U23758 (N_23758,N_23136,N_23030);
or U23759 (N_23759,N_23234,N_23054);
nor U23760 (N_23760,N_23400,N_23076);
or U23761 (N_23761,N_23174,N_23064);
or U23762 (N_23762,N_23052,N_23480);
or U23763 (N_23763,N_23327,N_23481);
xnor U23764 (N_23764,N_23182,N_23395);
nand U23765 (N_23765,N_23223,N_23116);
nor U23766 (N_23766,N_23428,N_23383);
and U23767 (N_23767,N_23476,N_23322);
or U23768 (N_23768,N_23108,N_23265);
or U23769 (N_23769,N_23040,N_23087);
or U23770 (N_23770,N_23425,N_23105);
or U23771 (N_23771,N_23437,N_23059);
xor U23772 (N_23772,N_23085,N_23213);
and U23773 (N_23773,N_23453,N_23226);
or U23774 (N_23774,N_23058,N_23014);
nand U23775 (N_23775,N_23446,N_23088);
or U23776 (N_23776,N_23373,N_23462);
xor U23777 (N_23777,N_23341,N_23056);
nand U23778 (N_23778,N_23377,N_23000);
xnor U23779 (N_23779,N_23395,N_23154);
or U23780 (N_23780,N_23286,N_23313);
nand U23781 (N_23781,N_23312,N_23223);
or U23782 (N_23782,N_23381,N_23213);
xor U23783 (N_23783,N_23165,N_23403);
and U23784 (N_23784,N_23136,N_23169);
or U23785 (N_23785,N_23230,N_23415);
xor U23786 (N_23786,N_23367,N_23196);
xnor U23787 (N_23787,N_23415,N_23041);
or U23788 (N_23788,N_23168,N_23171);
or U23789 (N_23789,N_23209,N_23231);
nor U23790 (N_23790,N_23001,N_23397);
nor U23791 (N_23791,N_23166,N_23098);
xor U23792 (N_23792,N_23230,N_23085);
and U23793 (N_23793,N_23003,N_23134);
or U23794 (N_23794,N_23101,N_23386);
or U23795 (N_23795,N_23277,N_23410);
or U23796 (N_23796,N_23004,N_23274);
and U23797 (N_23797,N_23203,N_23332);
nor U23798 (N_23798,N_23384,N_23051);
and U23799 (N_23799,N_23027,N_23257);
nand U23800 (N_23800,N_23361,N_23229);
xor U23801 (N_23801,N_23384,N_23143);
nand U23802 (N_23802,N_23061,N_23292);
nor U23803 (N_23803,N_23138,N_23416);
nor U23804 (N_23804,N_23188,N_23109);
nor U23805 (N_23805,N_23092,N_23441);
xor U23806 (N_23806,N_23129,N_23490);
and U23807 (N_23807,N_23154,N_23000);
xor U23808 (N_23808,N_23297,N_23036);
and U23809 (N_23809,N_23487,N_23438);
nor U23810 (N_23810,N_23302,N_23190);
or U23811 (N_23811,N_23329,N_23491);
nand U23812 (N_23812,N_23335,N_23257);
or U23813 (N_23813,N_23345,N_23183);
nand U23814 (N_23814,N_23201,N_23319);
nor U23815 (N_23815,N_23245,N_23370);
nor U23816 (N_23816,N_23267,N_23183);
nor U23817 (N_23817,N_23087,N_23255);
xor U23818 (N_23818,N_23473,N_23082);
or U23819 (N_23819,N_23054,N_23037);
or U23820 (N_23820,N_23092,N_23361);
nor U23821 (N_23821,N_23415,N_23190);
nor U23822 (N_23822,N_23048,N_23056);
nor U23823 (N_23823,N_23360,N_23188);
nand U23824 (N_23824,N_23298,N_23077);
nand U23825 (N_23825,N_23145,N_23374);
xnor U23826 (N_23826,N_23360,N_23114);
xor U23827 (N_23827,N_23437,N_23114);
nand U23828 (N_23828,N_23331,N_23083);
nand U23829 (N_23829,N_23322,N_23400);
nand U23830 (N_23830,N_23422,N_23347);
or U23831 (N_23831,N_23035,N_23135);
nor U23832 (N_23832,N_23162,N_23085);
xor U23833 (N_23833,N_23416,N_23299);
and U23834 (N_23834,N_23351,N_23030);
nor U23835 (N_23835,N_23018,N_23274);
nor U23836 (N_23836,N_23197,N_23449);
or U23837 (N_23837,N_23182,N_23141);
xor U23838 (N_23838,N_23028,N_23027);
nor U23839 (N_23839,N_23467,N_23074);
and U23840 (N_23840,N_23285,N_23261);
and U23841 (N_23841,N_23474,N_23146);
or U23842 (N_23842,N_23380,N_23360);
xnor U23843 (N_23843,N_23321,N_23441);
xnor U23844 (N_23844,N_23235,N_23390);
or U23845 (N_23845,N_23217,N_23056);
and U23846 (N_23846,N_23382,N_23195);
nor U23847 (N_23847,N_23260,N_23287);
nor U23848 (N_23848,N_23253,N_23287);
and U23849 (N_23849,N_23445,N_23211);
nand U23850 (N_23850,N_23473,N_23378);
nor U23851 (N_23851,N_23106,N_23296);
or U23852 (N_23852,N_23124,N_23122);
and U23853 (N_23853,N_23099,N_23340);
or U23854 (N_23854,N_23334,N_23097);
nor U23855 (N_23855,N_23326,N_23216);
nor U23856 (N_23856,N_23096,N_23121);
nor U23857 (N_23857,N_23492,N_23459);
nand U23858 (N_23858,N_23409,N_23098);
and U23859 (N_23859,N_23004,N_23454);
nor U23860 (N_23860,N_23233,N_23199);
xnor U23861 (N_23861,N_23233,N_23387);
or U23862 (N_23862,N_23271,N_23362);
xor U23863 (N_23863,N_23336,N_23076);
xor U23864 (N_23864,N_23251,N_23116);
nor U23865 (N_23865,N_23404,N_23027);
xor U23866 (N_23866,N_23488,N_23196);
nand U23867 (N_23867,N_23302,N_23425);
nand U23868 (N_23868,N_23096,N_23430);
nand U23869 (N_23869,N_23328,N_23409);
and U23870 (N_23870,N_23412,N_23212);
nor U23871 (N_23871,N_23409,N_23321);
or U23872 (N_23872,N_23159,N_23308);
or U23873 (N_23873,N_23272,N_23008);
nor U23874 (N_23874,N_23488,N_23124);
xor U23875 (N_23875,N_23436,N_23263);
xor U23876 (N_23876,N_23387,N_23289);
nor U23877 (N_23877,N_23213,N_23251);
nand U23878 (N_23878,N_23191,N_23139);
nor U23879 (N_23879,N_23235,N_23210);
or U23880 (N_23880,N_23374,N_23424);
xnor U23881 (N_23881,N_23203,N_23028);
nor U23882 (N_23882,N_23042,N_23430);
and U23883 (N_23883,N_23331,N_23089);
xor U23884 (N_23884,N_23115,N_23318);
nand U23885 (N_23885,N_23200,N_23029);
or U23886 (N_23886,N_23210,N_23263);
or U23887 (N_23887,N_23296,N_23437);
xnor U23888 (N_23888,N_23487,N_23172);
nand U23889 (N_23889,N_23222,N_23235);
xnor U23890 (N_23890,N_23447,N_23011);
and U23891 (N_23891,N_23038,N_23385);
or U23892 (N_23892,N_23155,N_23061);
or U23893 (N_23893,N_23079,N_23244);
nor U23894 (N_23894,N_23130,N_23196);
or U23895 (N_23895,N_23057,N_23015);
nand U23896 (N_23896,N_23352,N_23284);
and U23897 (N_23897,N_23122,N_23013);
nor U23898 (N_23898,N_23147,N_23140);
or U23899 (N_23899,N_23150,N_23112);
nor U23900 (N_23900,N_23152,N_23042);
and U23901 (N_23901,N_23049,N_23116);
nor U23902 (N_23902,N_23268,N_23183);
nand U23903 (N_23903,N_23178,N_23204);
nand U23904 (N_23904,N_23067,N_23237);
or U23905 (N_23905,N_23004,N_23078);
nand U23906 (N_23906,N_23109,N_23302);
nor U23907 (N_23907,N_23214,N_23303);
or U23908 (N_23908,N_23418,N_23140);
xnor U23909 (N_23909,N_23426,N_23388);
or U23910 (N_23910,N_23288,N_23290);
nand U23911 (N_23911,N_23342,N_23185);
nand U23912 (N_23912,N_23483,N_23257);
xnor U23913 (N_23913,N_23471,N_23109);
nand U23914 (N_23914,N_23313,N_23118);
and U23915 (N_23915,N_23302,N_23025);
and U23916 (N_23916,N_23330,N_23305);
and U23917 (N_23917,N_23161,N_23173);
and U23918 (N_23918,N_23433,N_23032);
and U23919 (N_23919,N_23093,N_23228);
and U23920 (N_23920,N_23296,N_23013);
xnor U23921 (N_23921,N_23321,N_23043);
or U23922 (N_23922,N_23332,N_23093);
nor U23923 (N_23923,N_23120,N_23464);
xor U23924 (N_23924,N_23293,N_23130);
and U23925 (N_23925,N_23499,N_23485);
xnor U23926 (N_23926,N_23048,N_23210);
nor U23927 (N_23927,N_23102,N_23082);
nand U23928 (N_23928,N_23374,N_23084);
nand U23929 (N_23929,N_23407,N_23089);
xnor U23930 (N_23930,N_23247,N_23353);
xnor U23931 (N_23931,N_23019,N_23389);
xnor U23932 (N_23932,N_23453,N_23156);
xor U23933 (N_23933,N_23422,N_23229);
and U23934 (N_23934,N_23478,N_23259);
nor U23935 (N_23935,N_23408,N_23308);
or U23936 (N_23936,N_23152,N_23255);
nor U23937 (N_23937,N_23497,N_23407);
xnor U23938 (N_23938,N_23138,N_23219);
nor U23939 (N_23939,N_23165,N_23119);
and U23940 (N_23940,N_23112,N_23147);
or U23941 (N_23941,N_23351,N_23059);
nor U23942 (N_23942,N_23156,N_23384);
nand U23943 (N_23943,N_23456,N_23395);
nand U23944 (N_23944,N_23029,N_23138);
xor U23945 (N_23945,N_23074,N_23095);
and U23946 (N_23946,N_23163,N_23361);
nand U23947 (N_23947,N_23328,N_23248);
and U23948 (N_23948,N_23306,N_23436);
nor U23949 (N_23949,N_23242,N_23317);
xor U23950 (N_23950,N_23269,N_23112);
and U23951 (N_23951,N_23176,N_23443);
nand U23952 (N_23952,N_23357,N_23468);
or U23953 (N_23953,N_23199,N_23113);
xor U23954 (N_23954,N_23348,N_23162);
nand U23955 (N_23955,N_23289,N_23321);
nor U23956 (N_23956,N_23059,N_23492);
nand U23957 (N_23957,N_23359,N_23060);
xnor U23958 (N_23958,N_23037,N_23367);
nor U23959 (N_23959,N_23119,N_23167);
nor U23960 (N_23960,N_23259,N_23280);
xnor U23961 (N_23961,N_23285,N_23134);
and U23962 (N_23962,N_23332,N_23420);
or U23963 (N_23963,N_23308,N_23492);
xor U23964 (N_23964,N_23310,N_23222);
nor U23965 (N_23965,N_23339,N_23372);
or U23966 (N_23966,N_23469,N_23425);
and U23967 (N_23967,N_23437,N_23233);
nand U23968 (N_23968,N_23319,N_23416);
and U23969 (N_23969,N_23235,N_23051);
and U23970 (N_23970,N_23219,N_23006);
and U23971 (N_23971,N_23302,N_23121);
and U23972 (N_23972,N_23174,N_23186);
xnor U23973 (N_23973,N_23234,N_23433);
or U23974 (N_23974,N_23392,N_23126);
and U23975 (N_23975,N_23146,N_23459);
nand U23976 (N_23976,N_23055,N_23018);
and U23977 (N_23977,N_23384,N_23110);
nor U23978 (N_23978,N_23062,N_23381);
or U23979 (N_23979,N_23041,N_23007);
nor U23980 (N_23980,N_23255,N_23212);
xor U23981 (N_23981,N_23403,N_23284);
nand U23982 (N_23982,N_23495,N_23127);
xor U23983 (N_23983,N_23170,N_23246);
and U23984 (N_23984,N_23103,N_23144);
or U23985 (N_23985,N_23098,N_23193);
xor U23986 (N_23986,N_23482,N_23075);
and U23987 (N_23987,N_23202,N_23113);
xor U23988 (N_23988,N_23283,N_23187);
or U23989 (N_23989,N_23372,N_23008);
xnor U23990 (N_23990,N_23163,N_23474);
nand U23991 (N_23991,N_23116,N_23169);
xnor U23992 (N_23992,N_23144,N_23467);
and U23993 (N_23993,N_23055,N_23118);
and U23994 (N_23994,N_23050,N_23409);
xor U23995 (N_23995,N_23236,N_23018);
or U23996 (N_23996,N_23390,N_23175);
xnor U23997 (N_23997,N_23329,N_23169);
or U23998 (N_23998,N_23297,N_23477);
and U23999 (N_23999,N_23208,N_23030);
xnor U24000 (N_24000,N_23535,N_23575);
nand U24001 (N_24001,N_23579,N_23619);
xor U24002 (N_24002,N_23545,N_23692);
nor U24003 (N_24003,N_23682,N_23863);
and U24004 (N_24004,N_23639,N_23968);
and U24005 (N_24005,N_23955,N_23733);
nor U24006 (N_24006,N_23807,N_23608);
and U24007 (N_24007,N_23844,N_23614);
or U24008 (N_24008,N_23696,N_23727);
and U24009 (N_24009,N_23930,N_23793);
and U24010 (N_24010,N_23675,N_23525);
nor U24011 (N_24011,N_23710,N_23849);
nor U24012 (N_24012,N_23636,N_23905);
or U24013 (N_24013,N_23702,N_23683);
and U24014 (N_24014,N_23739,N_23780);
xor U24015 (N_24015,N_23981,N_23559);
nand U24016 (N_24016,N_23956,N_23630);
and U24017 (N_24017,N_23954,N_23519);
or U24018 (N_24018,N_23982,N_23843);
and U24019 (N_24019,N_23764,N_23516);
xor U24020 (N_24020,N_23848,N_23761);
nand U24021 (N_24021,N_23914,N_23911);
or U24022 (N_24022,N_23817,N_23753);
or U24023 (N_24023,N_23534,N_23985);
xor U24024 (N_24024,N_23653,N_23869);
or U24025 (N_24025,N_23508,N_23890);
or U24026 (N_24026,N_23862,N_23677);
xnor U24027 (N_24027,N_23812,N_23760);
and U24028 (N_24028,N_23897,N_23808);
or U24029 (N_24029,N_23586,N_23705);
nor U24030 (N_24030,N_23703,N_23504);
nand U24031 (N_24031,N_23917,N_23767);
nand U24032 (N_24032,N_23782,N_23510);
or U24033 (N_24033,N_23688,N_23878);
nor U24034 (N_24034,N_23741,N_23737);
nor U24035 (N_24035,N_23648,N_23864);
or U24036 (N_24036,N_23563,N_23666);
nand U24037 (N_24037,N_23515,N_23526);
nand U24038 (N_24038,N_23555,N_23691);
nor U24039 (N_24039,N_23997,N_23953);
nor U24040 (N_24040,N_23960,N_23934);
nor U24041 (N_24041,N_23607,N_23791);
xor U24042 (N_24042,N_23789,N_23859);
xor U24043 (N_24043,N_23771,N_23970);
or U24044 (N_24044,N_23899,N_23883);
and U24045 (N_24045,N_23920,N_23731);
xnor U24046 (N_24046,N_23669,N_23501);
xor U24047 (N_24047,N_23873,N_23673);
nor U24048 (N_24048,N_23720,N_23948);
or U24049 (N_24049,N_23821,N_23540);
nand U24050 (N_24050,N_23832,N_23689);
or U24051 (N_24051,N_23854,N_23625);
and U24052 (N_24052,N_23851,N_23907);
and U24053 (N_24053,N_23750,N_23941);
nand U24054 (N_24054,N_23949,N_23599);
xor U24055 (N_24055,N_23923,N_23749);
and U24056 (N_24056,N_23711,N_23822);
or U24057 (N_24057,N_23751,N_23712);
xor U24058 (N_24058,N_23814,N_23652);
xnor U24059 (N_24059,N_23824,N_23600);
nor U24060 (N_24060,N_23745,N_23725);
and U24061 (N_24061,N_23581,N_23552);
xnor U24062 (N_24062,N_23604,N_23665);
xor U24063 (N_24063,N_23913,N_23734);
xnor U24064 (N_24064,N_23798,N_23646);
xor U24065 (N_24065,N_23518,N_23826);
or U24066 (N_24066,N_23717,N_23879);
or U24067 (N_24067,N_23908,N_23966);
xnor U24068 (N_24068,N_23950,N_23632);
xnor U24069 (N_24069,N_23794,N_23549);
or U24070 (N_24070,N_23983,N_23592);
and U24071 (N_24071,N_23947,N_23989);
and U24072 (N_24072,N_23620,N_23724);
nor U24073 (N_24073,N_23991,N_23583);
nand U24074 (N_24074,N_23503,N_23827);
and U24075 (N_24075,N_23758,N_23774);
xnor U24076 (N_24076,N_23886,N_23611);
nor U24077 (N_24077,N_23538,N_23634);
nor U24078 (N_24078,N_23776,N_23609);
nor U24079 (N_24079,N_23781,N_23603);
or U24080 (N_24080,N_23881,N_23612);
xor U24081 (N_24081,N_23649,N_23802);
nor U24082 (N_24082,N_23972,N_23938);
and U24083 (N_24083,N_23887,N_23530);
and U24084 (N_24084,N_23999,N_23514);
and U24085 (N_24085,N_23748,N_23763);
and U24086 (N_24086,N_23628,N_23617);
and U24087 (N_24087,N_23871,N_23951);
and U24088 (N_24088,N_23664,N_23942);
and U24089 (N_24089,N_23925,N_23594);
nor U24090 (N_24090,N_23513,N_23945);
nor U24091 (N_24091,N_23805,N_23896);
xnor U24092 (N_24092,N_23690,N_23796);
nor U24093 (N_24093,N_23775,N_23736);
nand U24094 (N_24094,N_23523,N_23909);
xnor U24095 (N_24095,N_23837,N_23527);
and U24096 (N_24096,N_23671,N_23921);
nand U24097 (N_24097,N_23601,N_23860);
nand U24098 (N_24098,N_23961,N_23517);
or U24099 (N_24099,N_23557,N_23658);
and U24100 (N_24100,N_23766,N_23926);
nor U24101 (N_24101,N_23792,N_23865);
xor U24102 (N_24102,N_23719,N_23629);
xor U24103 (N_24103,N_23606,N_23644);
nand U24104 (N_24104,N_23651,N_23694);
and U24105 (N_24105,N_23810,N_23785);
nor U24106 (N_24106,N_23853,N_23996);
nand U24107 (N_24107,N_23901,N_23551);
or U24108 (N_24108,N_23744,N_23521);
and U24109 (N_24109,N_23550,N_23693);
or U24110 (N_24110,N_23795,N_23978);
nor U24111 (N_24111,N_23566,N_23536);
and U24112 (N_24112,N_23587,N_23732);
and U24113 (N_24113,N_23828,N_23969);
nand U24114 (N_24114,N_23624,N_23957);
and U24115 (N_24115,N_23927,N_23561);
and U24116 (N_24116,N_23809,N_23786);
nor U24117 (N_24117,N_23856,N_23556);
nor U24118 (N_24118,N_23709,N_23505);
nand U24119 (N_24119,N_23582,N_23784);
nand U24120 (N_24120,N_23943,N_23571);
and U24121 (N_24121,N_23621,N_23993);
nand U24122 (N_24122,N_23546,N_23919);
or U24123 (N_24123,N_23880,N_23799);
nor U24124 (N_24124,N_23980,N_23532);
xnor U24125 (N_24125,N_23623,N_23512);
or U24126 (N_24126,N_23971,N_23678);
and U24127 (N_24127,N_23576,N_23506);
xor U24128 (N_24128,N_23681,N_23788);
xnor U24129 (N_24129,N_23698,N_23715);
and U24130 (N_24130,N_23700,N_23577);
nor U24131 (N_24131,N_23975,N_23801);
and U24132 (N_24132,N_23833,N_23752);
nand U24133 (N_24133,N_23936,N_23699);
xor U24134 (N_24134,N_23631,N_23830);
xnor U24135 (N_24135,N_23906,N_23659);
nor U24136 (N_24136,N_23730,N_23595);
or U24137 (N_24137,N_23959,N_23772);
and U24138 (N_24138,N_23935,N_23618);
or U24139 (N_24139,N_23918,N_23662);
or U24140 (N_24140,N_23637,N_23965);
nand U24141 (N_24141,N_23858,N_23522);
xnor U24142 (N_24142,N_23850,N_23584);
and U24143 (N_24143,N_23687,N_23861);
nand U24144 (N_24144,N_23562,N_23531);
xnor U24145 (N_24145,N_23539,N_23667);
nor U24146 (N_24146,N_23759,N_23819);
nand U24147 (N_24147,N_23708,N_23726);
nand U24148 (N_24148,N_23568,N_23963);
xnor U24149 (N_24149,N_23613,N_23704);
nor U24150 (N_24150,N_23580,N_23656);
nand U24151 (N_24151,N_23891,N_23500);
xor U24152 (N_24152,N_23533,N_23615);
nor U24153 (N_24153,N_23770,N_23790);
and U24154 (N_24154,N_23610,N_23962);
or U24155 (N_24155,N_23952,N_23984);
xnor U24156 (N_24156,N_23643,N_23815);
or U24157 (N_24157,N_23787,N_23835);
nand U24158 (N_24158,N_23569,N_23976);
and U24159 (N_24159,N_23560,N_23912);
or U24160 (N_24160,N_23820,N_23910);
xnor U24161 (N_24161,N_23857,N_23695);
nor U24162 (N_24162,N_23627,N_23834);
and U24163 (N_24163,N_23803,N_23944);
xor U24164 (N_24164,N_23616,N_23721);
and U24165 (N_24165,N_23564,N_23924);
nor U24166 (N_24166,N_23641,N_23977);
and U24167 (N_24167,N_23742,N_23738);
and U24168 (N_24168,N_23757,N_23988);
xnor U24169 (N_24169,N_23929,N_23686);
and U24170 (N_24170,N_23747,N_23816);
xor U24171 (N_24171,N_23697,N_23889);
nor U24172 (N_24172,N_23893,N_23746);
nand U24173 (N_24173,N_23855,N_23638);
nand U24174 (N_24174,N_23846,N_23743);
xnor U24175 (N_24175,N_23544,N_23847);
nor U24176 (N_24176,N_23633,N_23818);
or U24177 (N_24177,N_23714,N_23645);
or U24178 (N_24178,N_23868,N_23663);
and U24179 (N_24179,N_23845,N_23797);
or U24180 (N_24180,N_23565,N_23773);
nand U24181 (N_24181,N_23900,N_23590);
and U24182 (N_24182,N_23933,N_23554);
or U24183 (N_24183,N_23779,N_23931);
nor U24184 (N_24184,N_23578,N_23529);
nor U24185 (N_24185,N_23718,N_23974);
xnor U24186 (N_24186,N_23660,N_23867);
xnor U24187 (N_24187,N_23994,N_23622);
nand U24188 (N_24188,N_23987,N_23602);
or U24189 (N_24189,N_23588,N_23574);
and U24190 (N_24190,N_23528,N_23716);
and U24191 (N_24191,N_23915,N_23876);
and U24192 (N_24192,N_23916,N_23995);
xnor U24193 (N_24193,N_23713,N_23740);
nand U24194 (N_24194,N_23542,N_23946);
xnor U24195 (N_24195,N_23940,N_23875);
or U24196 (N_24196,N_23813,N_23723);
and U24197 (N_24197,N_23657,N_23573);
and U24198 (N_24198,N_23898,N_23722);
xor U24199 (N_24199,N_23676,N_23904);
nand U24200 (N_24200,N_23967,N_23836);
nor U24201 (N_24201,N_23992,N_23838);
nor U24202 (N_24202,N_23585,N_23541);
or U24203 (N_24203,N_23754,N_23706);
nand U24204 (N_24204,N_23597,N_23509);
or U24205 (N_24205,N_23511,N_23670);
and U24206 (N_24206,N_23762,N_23635);
and U24207 (N_24207,N_23894,N_23668);
xnor U24208 (N_24208,N_23884,N_23558);
or U24209 (N_24209,N_23839,N_23800);
xnor U24210 (N_24210,N_23735,N_23902);
nand U24211 (N_24211,N_23567,N_23877);
and U24212 (N_24212,N_23928,N_23769);
or U24213 (N_24213,N_23507,N_23661);
and U24214 (N_24214,N_23804,N_23707);
or U24215 (N_24215,N_23885,N_23841);
xnor U24216 (N_24216,N_23755,N_23605);
xnor U24217 (N_24217,N_23502,N_23840);
nor U24218 (N_24218,N_23593,N_23680);
nor U24219 (N_24219,N_23852,N_23831);
or U24220 (N_24220,N_23765,N_23537);
nand U24221 (N_24221,N_23986,N_23958);
and U24222 (N_24222,N_23672,N_23874);
and U24223 (N_24223,N_23596,N_23778);
or U24224 (N_24224,N_23570,N_23685);
and U24225 (N_24225,N_23728,N_23655);
xor U24226 (N_24226,N_23870,N_23756);
and U24227 (N_24227,N_23811,N_23640);
nor U24228 (N_24228,N_23524,N_23679);
and U24229 (N_24229,N_23547,N_23973);
nor U24230 (N_24230,N_23990,N_23591);
and U24231 (N_24231,N_23895,N_23939);
and U24232 (N_24232,N_23642,N_23674);
nor U24233 (N_24233,N_23892,N_23598);
and U24234 (N_24234,N_23806,N_23866);
and U24235 (N_24235,N_23882,N_23553);
or U24236 (N_24236,N_23729,N_23872);
xor U24237 (N_24237,N_23903,N_23829);
and U24238 (N_24238,N_23589,N_23932);
and U24239 (N_24239,N_23998,N_23701);
nor U24240 (N_24240,N_23654,N_23572);
nor U24241 (N_24241,N_23842,N_23543);
or U24242 (N_24242,N_23647,N_23979);
xnor U24243 (N_24243,N_23684,N_23823);
nor U24244 (N_24244,N_23626,N_23964);
and U24245 (N_24245,N_23777,N_23922);
and U24246 (N_24246,N_23768,N_23783);
and U24247 (N_24247,N_23888,N_23825);
and U24248 (N_24248,N_23937,N_23520);
nor U24249 (N_24249,N_23548,N_23650);
or U24250 (N_24250,N_23949,N_23989);
nand U24251 (N_24251,N_23880,N_23541);
xnor U24252 (N_24252,N_23523,N_23582);
xor U24253 (N_24253,N_23521,N_23904);
xnor U24254 (N_24254,N_23642,N_23949);
nor U24255 (N_24255,N_23796,N_23738);
or U24256 (N_24256,N_23604,N_23775);
nor U24257 (N_24257,N_23890,N_23800);
xnor U24258 (N_24258,N_23716,N_23824);
or U24259 (N_24259,N_23574,N_23870);
nand U24260 (N_24260,N_23840,N_23620);
or U24261 (N_24261,N_23850,N_23981);
and U24262 (N_24262,N_23961,N_23860);
nor U24263 (N_24263,N_23967,N_23527);
nor U24264 (N_24264,N_23951,N_23916);
and U24265 (N_24265,N_23730,N_23502);
and U24266 (N_24266,N_23609,N_23554);
and U24267 (N_24267,N_23928,N_23604);
xnor U24268 (N_24268,N_23506,N_23765);
and U24269 (N_24269,N_23566,N_23879);
nor U24270 (N_24270,N_23507,N_23994);
or U24271 (N_24271,N_23963,N_23818);
nor U24272 (N_24272,N_23809,N_23968);
and U24273 (N_24273,N_23583,N_23773);
nand U24274 (N_24274,N_23538,N_23777);
or U24275 (N_24275,N_23702,N_23892);
xnor U24276 (N_24276,N_23938,N_23704);
nor U24277 (N_24277,N_23570,N_23529);
or U24278 (N_24278,N_23999,N_23552);
xor U24279 (N_24279,N_23835,N_23834);
nor U24280 (N_24280,N_23709,N_23537);
or U24281 (N_24281,N_23635,N_23843);
nor U24282 (N_24282,N_23622,N_23626);
and U24283 (N_24283,N_23663,N_23693);
nor U24284 (N_24284,N_23809,N_23623);
or U24285 (N_24285,N_23954,N_23552);
xnor U24286 (N_24286,N_23554,N_23514);
or U24287 (N_24287,N_23837,N_23918);
and U24288 (N_24288,N_23707,N_23934);
nor U24289 (N_24289,N_23829,N_23966);
nand U24290 (N_24290,N_23550,N_23974);
and U24291 (N_24291,N_23546,N_23511);
xor U24292 (N_24292,N_23819,N_23908);
or U24293 (N_24293,N_23770,N_23776);
nand U24294 (N_24294,N_23724,N_23817);
or U24295 (N_24295,N_23751,N_23851);
nor U24296 (N_24296,N_23726,N_23730);
and U24297 (N_24297,N_23785,N_23560);
or U24298 (N_24298,N_23697,N_23835);
or U24299 (N_24299,N_23536,N_23859);
or U24300 (N_24300,N_23736,N_23529);
nor U24301 (N_24301,N_23966,N_23888);
and U24302 (N_24302,N_23705,N_23635);
nand U24303 (N_24303,N_23746,N_23691);
xnor U24304 (N_24304,N_23738,N_23828);
nor U24305 (N_24305,N_23632,N_23649);
xor U24306 (N_24306,N_23945,N_23984);
nand U24307 (N_24307,N_23533,N_23690);
nor U24308 (N_24308,N_23670,N_23604);
or U24309 (N_24309,N_23540,N_23786);
or U24310 (N_24310,N_23695,N_23963);
nor U24311 (N_24311,N_23817,N_23592);
and U24312 (N_24312,N_23609,N_23685);
nor U24313 (N_24313,N_23703,N_23981);
nand U24314 (N_24314,N_23517,N_23827);
xnor U24315 (N_24315,N_23995,N_23509);
xor U24316 (N_24316,N_23644,N_23773);
nor U24317 (N_24317,N_23699,N_23889);
or U24318 (N_24318,N_23701,N_23987);
and U24319 (N_24319,N_23695,N_23527);
or U24320 (N_24320,N_23788,N_23957);
nor U24321 (N_24321,N_23916,N_23810);
and U24322 (N_24322,N_23792,N_23535);
nand U24323 (N_24323,N_23665,N_23519);
xor U24324 (N_24324,N_23535,N_23801);
or U24325 (N_24325,N_23793,N_23605);
xor U24326 (N_24326,N_23931,N_23816);
and U24327 (N_24327,N_23730,N_23917);
and U24328 (N_24328,N_23548,N_23882);
and U24329 (N_24329,N_23802,N_23579);
nand U24330 (N_24330,N_23848,N_23770);
nor U24331 (N_24331,N_23845,N_23787);
xnor U24332 (N_24332,N_23515,N_23736);
nand U24333 (N_24333,N_23534,N_23535);
and U24334 (N_24334,N_23844,N_23796);
xor U24335 (N_24335,N_23999,N_23804);
nand U24336 (N_24336,N_23575,N_23697);
and U24337 (N_24337,N_23872,N_23632);
or U24338 (N_24338,N_23905,N_23903);
nor U24339 (N_24339,N_23558,N_23517);
nand U24340 (N_24340,N_23760,N_23687);
nand U24341 (N_24341,N_23921,N_23576);
nor U24342 (N_24342,N_23548,N_23962);
nor U24343 (N_24343,N_23602,N_23940);
xnor U24344 (N_24344,N_23888,N_23943);
nand U24345 (N_24345,N_23710,N_23574);
and U24346 (N_24346,N_23553,N_23579);
or U24347 (N_24347,N_23524,N_23836);
xnor U24348 (N_24348,N_23839,N_23684);
and U24349 (N_24349,N_23946,N_23947);
xnor U24350 (N_24350,N_23854,N_23601);
or U24351 (N_24351,N_23789,N_23722);
and U24352 (N_24352,N_23833,N_23747);
xor U24353 (N_24353,N_23982,N_23999);
nor U24354 (N_24354,N_23546,N_23660);
nand U24355 (N_24355,N_23549,N_23577);
nand U24356 (N_24356,N_23592,N_23978);
xor U24357 (N_24357,N_23667,N_23850);
xor U24358 (N_24358,N_23853,N_23713);
xor U24359 (N_24359,N_23721,N_23888);
and U24360 (N_24360,N_23528,N_23920);
xnor U24361 (N_24361,N_23847,N_23970);
and U24362 (N_24362,N_23502,N_23718);
xor U24363 (N_24363,N_23544,N_23659);
and U24364 (N_24364,N_23742,N_23897);
and U24365 (N_24365,N_23859,N_23745);
nor U24366 (N_24366,N_23798,N_23700);
or U24367 (N_24367,N_23887,N_23863);
xor U24368 (N_24368,N_23522,N_23620);
and U24369 (N_24369,N_23650,N_23565);
and U24370 (N_24370,N_23995,N_23752);
nor U24371 (N_24371,N_23877,N_23722);
or U24372 (N_24372,N_23925,N_23949);
nor U24373 (N_24373,N_23629,N_23976);
nand U24374 (N_24374,N_23690,N_23640);
and U24375 (N_24375,N_23772,N_23588);
nor U24376 (N_24376,N_23751,N_23721);
or U24377 (N_24377,N_23602,N_23855);
or U24378 (N_24378,N_23616,N_23760);
and U24379 (N_24379,N_23710,N_23627);
xnor U24380 (N_24380,N_23811,N_23520);
or U24381 (N_24381,N_23980,N_23865);
and U24382 (N_24382,N_23950,N_23552);
nor U24383 (N_24383,N_23643,N_23562);
or U24384 (N_24384,N_23786,N_23615);
nand U24385 (N_24385,N_23816,N_23518);
nand U24386 (N_24386,N_23591,N_23576);
nor U24387 (N_24387,N_23994,N_23517);
xor U24388 (N_24388,N_23964,N_23829);
nor U24389 (N_24389,N_23674,N_23916);
nor U24390 (N_24390,N_23911,N_23743);
and U24391 (N_24391,N_23914,N_23832);
nor U24392 (N_24392,N_23598,N_23796);
and U24393 (N_24393,N_23769,N_23654);
nor U24394 (N_24394,N_23501,N_23582);
xor U24395 (N_24395,N_23779,N_23751);
or U24396 (N_24396,N_23753,N_23762);
nor U24397 (N_24397,N_23859,N_23874);
xor U24398 (N_24398,N_23888,N_23983);
and U24399 (N_24399,N_23827,N_23572);
nor U24400 (N_24400,N_23955,N_23985);
nor U24401 (N_24401,N_23624,N_23688);
xor U24402 (N_24402,N_23932,N_23906);
xor U24403 (N_24403,N_23680,N_23717);
or U24404 (N_24404,N_23951,N_23600);
and U24405 (N_24405,N_23999,N_23596);
and U24406 (N_24406,N_23502,N_23702);
nor U24407 (N_24407,N_23597,N_23691);
or U24408 (N_24408,N_23585,N_23829);
or U24409 (N_24409,N_23982,N_23896);
nand U24410 (N_24410,N_23774,N_23869);
nor U24411 (N_24411,N_23861,N_23926);
nand U24412 (N_24412,N_23844,N_23574);
or U24413 (N_24413,N_23545,N_23591);
nand U24414 (N_24414,N_23841,N_23592);
nand U24415 (N_24415,N_23830,N_23717);
nand U24416 (N_24416,N_23780,N_23741);
nor U24417 (N_24417,N_23830,N_23998);
nand U24418 (N_24418,N_23643,N_23904);
and U24419 (N_24419,N_23871,N_23558);
nor U24420 (N_24420,N_23795,N_23555);
and U24421 (N_24421,N_23639,N_23652);
nand U24422 (N_24422,N_23984,N_23961);
xor U24423 (N_24423,N_23570,N_23621);
and U24424 (N_24424,N_23591,N_23750);
nor U24425 (N_24425,N_23675,N_23897);
and U24426 (N_24426,N_23907,N_23692);
or U24427 (N_24427,N_23748,N_23894);
and U24428 (N_24428,N_23976,N_23827);
xor U24429 (N_24429,N_23850,N_23505);
nor U24430 (N_24430,N_23675,N_23917);
xor U24431 (N_24431,N_23827,N_23874);
nor U24432 (N_24432,N_23541,N_23540);
or U24433 (N_24433,N_23817,N_23751);
and U24434 (N_24434,N_23654,N_23971);
and U24435 (N_24435,N_23605,N_23981);
and U24436 (N_24436,N_23674,N_23502);
nor U24437 (N_24437,N_23700,N_23790);
xor U24438 (N_24438,N_23879,N_23900);
or U24439 (N_24439,N_23728,N_23886);
nand U24440 (N_24440,N_23589,N_23882);
or U24441 (N_24441,N_23931,N_23608);
xnor U24442 (N_24442,N_23871,N_23959);
and U24443 (N_24443,N_23701,N_23883);
or U24444 (N_24444,N_23543,N_23692);
or U24445 (N_24445,N_23945,N_23542);
nand U24446 (N_24446,N_23630,N_23544);
or U24447 (N_24447,N_23983,N_23576);
nor U24448 (N_24448,N_23991,N_23901);
nor U24449 (N_24449,N_23834,N_23761);
xnor U24450 (N_24450,N_23744,N_23570);
xor U24451 (N_24451,N_23869,N_23977);
xor U24452 (N_24452,N_23615,N_23593);
and U24453 (N_24453,N_23731,N_23647);
xnor U24454 (N_24454,N_23601,N_23924);
nor U24455 (N_24455,N_23512,N_23884);
nor U24456 (N_24456,N_23892,N_23813);
nor U24457 (N_24457,N_23523,N_23861);
nor U24458 (N_24458,N_23708,N_23721);
and U24459 (N_24459,N_23822,N_23717);
xor U24460 (N_24460,N_23966,N_23601);
xnor U24461 (N_24461,N_23504,N_23840);
nor U24462 (N_24462,N_23897,N_23946);
or U24463 (N_24463,N_23715,N_23605);
xor U24464 (N_24464,N_23639,N_23630);
and U24465 (N_24465,N_23654,N_23506);
or U24466 (N_24466,N_23662,N_23863);
or U24467 (N_24467,N_23627,N_23823);
nor U24468 (N_24468,N_23585,N_23758);
and U24469 (N_24469,N_23617,N_23696);
nor U24470 (N_24470,N_23948,N_23696);
and U24471 (N_24471,N_23851,N_23512);
nand U24472 (N_24472,N_23889,N_23547);
nand U24473 (N_24473,N_23843,N_23868);
nand U24474 (N_24474,N_23628,N_23816);
nand U24475 (N_24475,N_23546,N_23996);
xnor U24476 (N_24476,N_23765,N_23606);
nor U24477 (N_24477,N_23576,N_23773);
nor U24478 (N_24478,N_23509,N_23810);
or U24479 (N_24479,N_23743,N_23598);
nand U24480 (N_24480,N_23906,N_23646);
and U24481 (N_24481,N_23843,N_23634);
nor U24482 (N_24482,N_23580,N_23617);
nand U24483 (N_24483,N_23707,N_23596);
nor U24484 (N_24484,N_23707,N_23915);
and U24485 (N_24485,N_23683,N_23728);
nor U24486 (N_24486,N_23562,N_23558);
nand U24487 (N_24487,N_23534,N_23577);
and U24488 (N_24488,N_23528,N_23805);
and U24489 (N_24489,N_23577,N_23690);
xor U24490 (N_24490,N_23659,N_23986);
xnor U24491 (N_24491,N_23774,N_23608);
xor U24492 (N_24492,N_23625,N_23987);
xor U24493 (N_24493,N_23669,N_23585);
nor U24494 (N_24494,N_23610,N_23906);
nand U24495 (N_24495,N_23846,N_23702);
or U24496 (N_24496,N_23536,N_23540);
nor U24497 (N_24497,N_23606,N_23907);
nand U24498 (N_24498,N_23588,N_23963);
nand U24499 (N_24499,N_23569,N_23854);
nor U24500 (N_24500,N_24394,N_24267);
nor U24501 (N_24501,N_24068,N_24283);
or U24502 (N_24502,N_24027,N_24390);
nor U24503 (N_24503,N_24452,N_24365);
nand U24504 (N_24504,N_24228,N_24181);
and U24505 (N_24505,N_24387,N_24045);
nor U24506 (N_24506,N_24429,N_24257);
or U24507 (N_24507,N_24233,N_24080);
and U24508 (N_24508,N_24310,N_24294);
or U24509 (N_24509,N_24292,N_24477);
nand U24510 (N_24510,N_24434,N_24130);
and U24511 (N_24511,N_24026,N_24082);
xor U24512 (N_24512,N_24201,N_24030);
and U24513 (N_24513,N_24316,N_24115);
or U24514 (N_24514,N_24392,N_24352);
nand U24515 (N_24515,N_24448,N_24170);
nand U24516 (N_24516,N_24290,N_24463);
or U24517 (N_24517,N_24091,N_24043);
nand U24518 (N_24518,N_24395,N_24203);
or U24519 (N_24519,N_24286,N_24415);
or U24520 (N_24520,N_24156,N_24111);
nor U24521 (N_24521,N_24260,N_24422);
or U24522 (N_24522,N_24213,N_24424);
or U24523 (N_24523,N_24188,N_24447);
or U24524 (N_24524,N_24299,N_24140);
or U24525 (N_24525,N_24276,N_24350);
nor U24526 (N_24526,N_24024,N_24278);
and U24527 (N_24527,N_24444,N_24218);
or U24528 (N_24528,N_24410,N_24133);
nor U24529 (N_24529,N_24139,N_24351);
or U24530 (N_24530,N_24408,N_24012);
nor U24531 (N_24531,N_24479,N_24000);
and U24532 (N_24532,N_24413,N_24281);
nand U24533 (N_24533,N_24186,N_24033);
or U24534 (N_24534,N_24246,N_24102);
nor U24535 (N_24535,N_24377,N_24226);
nand U24536 (N_24536,N_24180,N_24343);
nor U24537 (N_24537,N_24255,N_24028);
xor U24538 (N_24538,N_24245,N_24217);
and U24539 (N_24539,N_24264,N_24402);
xor U24540 (N_24540,N_24490,N_24083);
nor U24541 (N_24541,N_24442,N_24318);
and U24542 (N_24542,N_24456,N_24306);
xnor U24543 (N_24543,N_24090,N_24057);
and U24544 (N_24544,N_24066,N_24248);
or U24545 (N_24545,N_24164,N_24025);
xnor U24546 (N_24546,N_24104,N_24037);
and U24547 (N_24547,N_24337,N_24240);
xor U24548 (N_24548,N_24405,N_24055);
xor U24549 (N_24549,N_24342,N_24443);
xnor U24550 (N_24550,N_24189,N_24330);
and U24551 (N_24551,N_24433,N_24389);
or U24552 (N_24552,N_24348,N_24372);
nor U24553 (N_24553,N_24417,N_24259);
xor U24554 (N_24554,N_24344,N_24438);
xnor U24555 (N_24555,N_24145,N_24089);
nor U24556 (N_24556,N_24243,N_24385);
xor U24557 (N_24557,N_24063,N_24303);
xnor U24558 (N_24558,N_24093,N_24378);
or U24559 (N_24559,N_24108,N_24038);
or U24560 (N_24560,N_24478,N_24244);
nor U24561 (N_24561,N_24101,N_24483);
xor U24562 (N_24562,N_24430,N_24197);
or U24563 (N_24563,N_24056,N_24327);
nand U24564 (N_24564,N_24380,N_24224);
and U24565 (N_24565,N_24031,N_24412);
nand U24566 (N_24566,N_24127,N_24174);
and U24567 (N_24567,N_24455,N_24453);
nor U24568 (N_24568,N_24166,N_24185);
nand U24569 (N_24569,N_24150,N_24153);
or U24570 (N_24570,N_24268,N_24262);
nor U24571 (N_24571,N_24288,N_24274);
nor U24572 (N_24572,N_24225,N_24400);
nor U24573 (N_24573,N_24032,N_24103);
or U24574 (N_24574,N_24016,N_24003);
and U24575 (N_24575,N_24357,N_24207);
nor U24576 (N_24576,N_24148,N_24009);
or U24577 (N_24577,N_24384,N_24237);
xnor U24578 (N_24578,N_24250,N_24152);
nand U24579 (N_24579,N_24311,N_24285);
xnor U24580 (N_24580,N_24323,N_24060);
nand U24581 (N_24581,N_24113,N_24086);
nand U24582 (N_24582,N_24373,N_24094);
and U24583 (N_24583,N_24110,N_24044);
or U24584 (N_24584,N_24041,N_24142);
nor U24585 (N_24585,N_24172,N_24469);
nand U24586 (N_24586,N_24013,N_24079);
nand U24587 (N_24587,N_24336,N_24229);
nand U24588 (N_24588,N_24121,N_24124);
and U24589 (N_24589,N_24070,N_24112);
or U24590 (N_24590,N_24282,N_24129);
and U24591 (N_24591,N_24100,N_24474);
xor U24592 (N_24592,N_24499,N_24252);
nand U24593 (N_24593,N_24401,N_24017);
and U24594 (N_24594,N_24418,N_24349);
nor U24595 (N_24595,N_24374,N_24048);
and U24596 (N_24596,N_24460,N_24138);
and U24597 (N_24597,N_24347,N_24194);
nand U24598 (N_24598,N_24409,N_24004);
and U24599 (N_24599,N_24445,N_24471);
and U24600 (N_24600,N_24404,N_24457);
xnor U24601 (N_24601,N_24298,N_24010);
and U24602 (N_24602,N_24488,N_24297);
xor U24603 (N_24603,N_24398,N_24362);
xor U24604 (N_24604,N_24493,N_24421);
and U24605 (N_24605,N_24314,N_24432);
nand U24606 (N_24606,N_24122,N_24458);
nor U24607 (N_24607,N_24466,N_24162);
or U24608 (N_24608,N_24269,N_24085);
xnor U24609 (N_24609,N_24075,N_24007);
nor U24610 (N_24610,N_24489,N_24454);
or U24611 (N_24611,N_24420,N_24199);
nor U24612 (N_24612,N_24114,N_24258);
xnor U24613 (N_24613,N_24099,N_24064);
nor U24614 (N_24614,N_24161,N_24339);
nor U24615 (N_24615,N_24325,N_24036);
and U24616 (N_24616,N_24497,N_24359);
and U24617 (N_24617,N_24241,N_24220);
or U24618 (N_24618,N_24173,N_24167);
nor U24619 (N_24619,N_24144,N_24334);
xnor U24620 (N_24620,N_24169,N_24480);
nor U24621 (N_24621,N_24072,N_24295);
and U24622 (N_24622,N_24071,N_24467);
xor U24623 (N_24623,N_24475,N_24096);
xor U24624 (N_24624,N_24222,N_24053);
and U24625 (N_24625,N_24427,N_24481);
xor U24626 (N_24626,N_24216,N_24494);
xnor U24627 (N_24627,N_24131,N_24040);
or U24628 (N_24628,N_24440,N_24046);
or U24629 (N_24629,N_24491,N_24206);
or U24630 (N_24630,N_24451,N_24322);
and U24631 (N_24631,N_24340,N_24472);
xnor U24632 (N_24632,N_24204,N_24035);
and U24633 (N_24633,N_24230,N_24338);
nand U24634 (N_24634,N_24446,N_24183);
xnor U24635 (N_24635,N_24239,N_24158);
nand U24636 (N_24636,N_24175,N_24399);
nand U24637 (N_24637,N_24134,N_24386);
xor U24638 (N_24638,N_24067,N_24461);
nor U24639 (N_24639,N_24118,N_24223);
xnor U24640 (N_24640,N_24371,N_24363);
nand U24641 (N_24641,N_24383,N_24059);
nor U24642 (N_24642,N_24492,N_24021);
nor U24643 (N_24643,N_24346,N_24023);
xor U24644 (N_24644,N_24496,N_24088);
xor U24645 (N_24645,N_24095,N_24279);
and U24646 (N_24646,N_24272,N_24428);
or U24647 (N_24647,N_24084,N_24092);
and U24648 (N_24648,N_24050,N_24355);
nor U24649 (N_24649,N_24304,N_24202);
xor U24650 (N_24650,N_24317,N_24368);
and U24651 (N_24651,N_24253,N_24136);
nand U24652 (N_24652,N_24198,N_24366);
and U24653 (N_24653,N_24364,N_24081);
nor U24654 (N_24654,N_24116,N_24414);
xor U24655 (N_24655,N_24179,N_24293);
or U24656 (N_24656,N_24097,N_24157);
and U24657 (N_24657,N_24376,N_24196);
nor U24658 (N_24658,N_24423,N_24263);
and U24659 (N_24659,N_24192,N_24087);
nor U24660 (N_24660,N_24375,N_24411);
nor U24661 (N_24661,N_24464,N_24242);
xnor U24662 (N_24662,N_24042,N_24333);
xnor U24663 (N_24663,N_24345,N_24277);
xor U24664 (N_24664,N_24117,N_24001);
nand U24665 (N_24665,N_24227,N_24331);
nor U24666 (N_24666,N_24234,N_24212);
nor U24667 (N_24667,N_24495,N_24238);
nor U24668 (N_24668,N_24107,N_24356);
nor U24669 (N_24669,N_24190,N_24321);
xor U24670 (N_24670,N_24221,N_24052);
and U24671 (N_24671,N_24369,N_24120);
or U24672 (N_24672,N_24441,N_24029);
nor U24673 (N_24673,N_24098,N_24315);
and U24674 (N_24674,N_24137,N_24284);
xor U24675 (N_24675,N_24425,N_24486);
nand U24676 (N_24676,N_24435,N_24119);
or U24677 (N_24677,N_24125,N_24065);
nand U24678 (N_24678,N_24312,N_24436);
nor U24679 (N_24679,N_24014,N_24476);
and U24680 (N_24680,N_24002,N_24324);
xnor U24681 (N_24681,N_24379,N_24426);
or U24682 (N_24682,N_24210,N_24354);
or U24683 (N_24683,N_24008,N_24132);
nor U24684 (N_24684,N_24465,N_24361);
nand U24685 (N_24685,N_24236,N_24209);
and U24686 (N_24686,N_24177,N_24047);
nand U24687 (N_24687,N_24232,N_24215);
nand U24688 (N_24688,N_24431,N_24061);
xor U24689 (N_24689,N_24256,N_24069);
and U24690 (N_24690,N_24214,N_24468);
nand U24691 (N_24691,N_24109,N_24291);
and U24692 (N_24692,N_24018,N_24039);
and U24693 (N_24693,N_24473,N_24074);
and U24694 (N_24694,N_24105,N_24106);
or U24695 (N_24695,N_24126,N_24205);
or U24696 (N_24696,N_24459,N_24320);
nor U24697 (N_24697,N_24020,N_24381);
nand U24698 (N_24698,N_24128,N_24187);
nand U24699 (N_24699,N_24271,N_24329);
xor U24700 (N_24700,N_24151,N_24358);
xor U24701 (N_24701,N_24309,N_24034);
xor U24702 (N_24702,N_24165,N_24168);
or U24703 (N_24703,N_24022,N_24076);
nor U24704 (N_24704,N_24270,N_24154);
and U24705 (N_24705,N_24184,N_24077);
and U24706 (N_24706,N_24247,N_24135);
nand U24707 (N_24707,N_24307,N_24388);
and U24708 (N_24708,N_24178,N_24147);
nor U24709 (N_24709,N_24054,N_24470);
nand U24710 (N_24710,N_24498,N_24300);
nor U24711 (N_24711,N_24419,N_24397);
xnor U24712 (N_24712,N_24462,N_24005);
nor U24713 (N_24713,N_24332,N_24328);
nor U24714 (N_24714,N_24249,N_24143);
xor U24715 (N_24715,N_24275,N_24261);
xor U24716 (N_24716,N_24266,N_24406);
nand U24717 (N_24717,N_24211,N_24171);
or U24718 (N_24718,N_24407,N_24254);
or U24719 (N_24719,N_24450,N_24319);
nor U24720 (N_24720,N_24302,N_24195);
and U24721 (N_24721,N_24487,N_24200);
xnor U24722 (N_24722,N_24123,N_24287);
nand U24723 (N_24723,N_24208,N_24073);
nor U24724 (N_24724,N_24437,N_24149);
nor U24725 (N_24725,N_24191,N_24391);
nand U24726 (N_24726,N_24360,N_24019);
nor U24727 (N_24727,N_24155,N_24078);
and U24728 (N_24728,N_24062,N_24051);
nand U24729 (N_24729,N_24289,N_24382);
nor U24730 (N_24730,N_24308,N_24058);
or U24731 (N_24731,N_24403,N_24439);
nand U24732 (N_24732,N_24273,N_24393);
nor U24733 (N_24733,N_24301,N_24163);
or U24734 (N_24734,N_24416,N_24231);
xor U24735 (N_24735,N_24193,N_24296);
nor U24736 (N_24736,N_24341,N_24305);
nand U24737 (N_24737,N_24141,N_24011);
nor U24738 (N_24738,N_24265,N_24335);
xnor U24739 (N_24739,N_24251,N_24449);
or U24740 (N_24740,N_24049,N_24485);
nand U24741 (N_24741,N_24313,N_24367);
or U24742 (N_24742,N_24482,N_24160);
nor U24743 (N_24743,N_24219,N_24396);
nand U24744 (N_24744,N_24176,N_24146);
nand U24745 (N_24745,N_24353,N_24159);
or U24746 (N_24746,N_24015,N_24006);
nand U24747 (N_24747,N_24484,N_24182);
nor U24748 (N_24748,N_24326,N_24370);
nand U24749 (N_24749,N_24235,N_24280);
and U24750 (N_24750,N_24074,N_24398);
xor U24751 (N_24751,N_24089,N_24020);
xnor U24752 (N_24752,N_24190,N_24128);
and U24753 (N_24753,N_24068,N_24461);
or U24754 (N_24754,N_24272,N_24233);
and U24755 (N_24755,N_24138,N_24335);
and U24756 (N_24756,N_24094,N_24231);
xor U24757 (N_24757,N_24076,N_24289);
nor U24758 (N_24758,N_24163,N_24091);
xor U24759 (N_24759,N_24387,N_24193);
and U24760 (N_24760,N_24094,N_24392);
nand U24761 (N_24761,N_24405,N_24251);
nand U24762 (N_24762,N_24068,N_24491);
nor U24763 (N_24763,N_24111,N_24140);
nand U24764 (N_24764,N_24289,N_24332);
xnor U24765 (N_24765,N_24231,N_24469);
nand U24766 (N_24766,N_24330,N_24115);
and U24767 (N_24767,N_24310,N_24311);
or U24768 (N_24768,N_24358,N_24338);
and U24769 (N_24769,N_24276,N_24294);
or U24770 (N_24770,N_24035,N_24278);
xnor U24771 (N_24771,N_24118,N_24421);
xor U24772 (N_24772,N_24302,N_24270);
xor U24773 (N_24773,N_24363,N_24031);
or U24774 (N_24774,N_24421,N_24161);
or U24775 (N_24775,N_24146,N_24413);
or U24776 (N_24776,N_24410,N_24283);
nand U24777 (N_24777,N_24361,N_24379);
and U24778 (N_24778,N_24367,N_24086);
and U24779 (N_24779,N_24270,N_24304);
nor U24780 (N_24780,N_24118,N_24462);
nand U24781 (N_24781,N_24454,N_24194);
xnor U24782 (N_24782,N_24077,N_24297);
or U24783 (N_24783,N_24434,N_24479);
xor U24784 (N_24784,N_24270,N_24228);
nand U24785 (N_24785,N_24097,N_24234);
xnor U24786 (N_24786,N_24378,N_24236);
nand U24787 (N_24787,N_24139,N_24227);
nand U24788 (N_24788,N_24452,N_24021);
nor U24789 (N_24789,N_24488,N_24150);
nor U24790 (N_24790,N_24071,N_24216);
nor U24791 (N_24791,N_24109,N_24459);
nor U24792 (N_24792,N_24352,N_24434);
nor U24793 (N_24793,N_24356,N_24265);
or U24794 (N_24794,N_24498,N_24383);
or U24795 (N_24795,N_24087,N_24404);
or U24796 (N_24796,N_24095,N_24478);
and U24797 (N_24797,N_24214,N_24057);
and U24798 (N_24798,N_24045,N_24053);
or U24799 (N_24799,N_24280,N_24313);
nor U24800 (N_24800,N_24043,N_24491);
nor U24801 (N_24801,N_24238,N_24200);
nand U24802 (N_24802,N_24374,N_24226);
nand U24803 (N_24803,N_24319,N_24122);
and U24804 (N_24804,N_24240,N_24333);
and U24805 (N_24805,N_24365,N_24062);
or U24806 (N_24806,N_24280,N_24037);
or U24807 (N_24807,N_24464,N_24357);
xor U24808 (N_24808,N_24466,N_24195);
xor U24809 (N_24809,N_24200,N_24256);
or U24810 (N_24810,N_24473,N_24152);
and U24811 (N_24811,N_24128,N_24478);
or U24812 (N_24812,N_24040,N_24258);
and U24813 (N_24813,N_24120,N_24071);
or U24814 (N_24814,N_24307,N_24135);
xnor U24815 (N_24815,N_24065,N_24239);
nor U24816 (N_24816,N_24385,N_24349);
or U24817 (N_24817,N_24369,N_24065);
nand U24818 (N_24818,N_24236,N_24456);
xnor U24819 (N_24819,N_24077,N_24390);
xor U24820 (N_24820,N_24309,N_24445);
nor U24821 (N_24821,N_24111,N_24339);
nor U24822 (N_24822,N_24152,N_24347);
nand U24823 (N_24823,N_24195,N_24277);
or U24824 (N_24824,N_24119,N_24413);
and U24825 (N_24825,N_24018,N_24315);
nor U24826 (N_24826,N_24472,N_24218);
nor U24827 (N_24827,N_24016,N_24238);
xnor U24828 (N_24828,N_24312,N_24335);
nand U24829 (N_24829,N_24268,N_24293);
nand U24830 (N_24830,N_24386,N_24317);
and U24831 (N_24831,N_24490,N_24184);
or U24832 (N_24832,N_24497,N_24187);
nor U24833 (N_24833,N_24423,N_24122);
and U24834 (N_24834,N_24304,N_24204);
nor U24835 (N_24835,N_24336,N_24152);
or U24836 (N_24836,N_24332,N_24337);
nor U24837 (N_24837,N_24098,N_24474);
xnor U24838 (N_24838,N_24292,N_24448);
xnor U24839 (N_24839,N_24244,N_24222);
nor U24840 (N_24840,N_24479,N_24273);
nor U24841 (N_24841,N_24085,N_24048);
nor U24842 (N_24842,N_24011,N_24026);
and U24843 (N_24843,N_24456,N_24080);
nor U24844 (N_24844,N_24324,N_24087);
or U24845 (N_24845,N_24213,N_24053);
nor U24846 (N_24846,N_24092,N_24200);
and U24847 (N_24847,N_24184,N_24222);
and U24848 (N_24848,N_24021,N_24211);
and U24849 (N_24849,N_24015,N_24132);
xor U24850 (N_24850,N_24364,N_24052);
nor U24851 (N_24851,N_24279,N_24420);
xnor U24852 (N_24852,N_24192,N_24387);
xor U24853 (N_24853,N_24016,N_24082);
nor U24854 (N_24854,N_24069,N_24417);
nand U24855 (N_24855,N_24232,N_24090);
and U24856 (N_24856,N_24435,N_24149);
xnor U24857 (N_24857,N_24235,N_24291);
nand U24858 (N_24858,N_24421,N_24196);
nand U24859 (N_24859,N_24026,N_24303);
and U24860 (N_24860,N_24282,N_24367);
and U24861 (N_24861,N_24365,N_24481);
nand U24862 (N_24862,N_24284,N_24214);
xor U24863 (N_24863,N_24409,N_24372);
nor U24864 (N_24864,N_24019,N_24009);
or U24865 (N_24865,N_24119,N_24016);
or U24866 (N_24866,N_24117,N_24101);
and U24867 (N_24867,N_24344,N_24119);
or U24868 (N_24868,N_24330,N_24080);
nand U24869 (N_24869,N_24354,N_24338);
nand U24870 (N_24870,N_24089,N_24099);
or U24871 (N_24871,N_24073,N_24415);
nor U24872 (N_24872,N_24148,N_24256);
and U24873 (N_24873,N_24464,N_24143);
or U24874 (N_24874,N_24049,N_24140);
and U24875 (N_24875,N_24266,N_24150);
xor U24876 (N_24876,N_24256,N_24232);
nor U24877 (N_24877,N_24385,N_24205);
xnor U24878 (N_24878,N_24448,N_24101);
and U24879 (N_24879,N_24451,N_24376);
xor U24880 (N_24880,N_24205,N_24115);
xor U24881 (N_24881,N_24081,N_24137);
nand U24882 (N_24882,N_24048,N_24416);
and U24883 (N_24883,N_24024,N_24321);
or U24884 (N_24884,N_24436,N_24069);
nor U24885 (N_24885,N_24075,N_24185);
nor U24886 (N_24886,N_24445,N_24257);
or U24887 (N_24887,N_24141,N_24496);
nor U24888 (N_24888,N_24449,N_24415);
nand U24889 (N_24889,N_24114,N_24023);
xnor U24890 (N_24890,N_24170,N_24272);
nor U24891 (N_24891,N_24075,N_24488);
and U24892 (N_24892,N_24313,N_24306);
xnor U24893 (N_24893,N_24358,N_24197);
xnor U24894 (N_24894,N_24390,N_24324);
nor U24895 (N_24895,N_24175,N_24212);
or U24896 (N_24896,N_24467,N_24464);
xnor U24897 (N_24897,N_24143,N_24172);
and U24898 (N_24898,N_24053,N_24362);
or U24899 (N_24899,N_24028,N_24333);
or U24900 (N_24900,N_24458,N_24292);
and U24901 (N_24901,N_24340,N_24353);
xor U24902 (N_24902,N_24280,N_24103);
nand U24903 (N_24903,N_24437,N_24014);
nor U24904 (N_24904,N_24320,N_24340);
xnor U24905 (N_24905,N_24289,N_24050);
nand U24906 (N_24906,N_24115,N_24271);
nor U24907 (N_24907,N_24131,N_24322);
and U24908 (N_24908,N_24353,N_24396);
nand U24909 (N_24909,N_24461,N_24037);
nor U24910 (N_24910,N_24118,N_24228);
and U24911 (N_24911,N_24262,N_24125);
nand U24912 (N_24912,N_24115,N_24112);
nand U24913 (N_24913,N_24257,N_24181);
or U24914 (N_24914,N_24106,N_24441);
nand U24915 (N_24915,N_24441,N_24185);
nor U24916 (N_24916,N_24262,N_24283);
xor U24917 (N_24917,N_24490,N_24100);
and U24918 (N_24918,N_24288,N_24120);
or U24919 (N_24919,N_24064,N_24302);
xor U24920 (N_24920,N_24165,N_24414);
and U24921 (N_24921,N_24281,N_24439);
or U24922 (N_24922,N_24176,N_24257);
nor U24923 (N_24923,N_24100,N_24411);
xor U24924 (N_24924,N_24284,N_24317);
or U24925 (N_24925,N_24255,N_24359);
nor U24926 (N_24926,N_24318,N_24026);
or U24927 (N_24927,N_24417,N_24135);
xnor U24928 (N_24928,N_24451,N_24041);
nand U24929 (N_24929,N_24275,N_24151);
and U24930 (N_24930,N_24499,N_24481);
nor U24931 (N_24931,N_24369,N_24477);
and U24932 (N_24932,N_24411,N_24418);
or U24933 (N_24933,N_24220,N_24261);
xor U24934 (N_24934,N_24447,N_24255);
xnor U24935 (N_24935,N_24041,N_24220);
nand U24936 (N_24936,N_24278,N_24490);
nand U24937 (N_24937,N_24415,N_24135);
xnor U24938 (N_24938,N_24383,N_24487);
and U24939 (N_24939,N_24359,N_24061);
nand U24940 (N_24940,N_24309,N_24454);
nand U24941 (N_24941,N_24099,N_24117);
nor U24942 (N_24942,N_24201,N_24094);
xor U24943 (N_24943,N_24401,N_24423);
and U24944 (N_24944,N_24121,N_24091);
xor U24945 (N_24945,N_24176,N_24134);
and U24946 (N_24946,N_24320,N_24087);
or U24947 (N_24947,N_24391,N_24246);
nand U24948 (N_24948,N_24150,N_24121);
xor U24949 (N_24949,N_24305,N_24071);
xor U24950 (N_24950,N_24313,N_24344);
nor U24951 (N_24951,N_24473,N_24392);
and U24952 (N_24952,N_24114,N_24480);
or U24953 (N_24953,N_24102,N_24041);
or U24954 (N_24954,N_24401,N_24163);
and U24955 (N_24955,N_24186,N_24465);
or U24956 (N_24956,N_24447,N_24495);
xnor U24957 (N_24957,N_24116,N_24183);
nor U24958 (N_24958,N_24172,N_24373);
xor U24959 (N_24959,N_24003,N_24437);
nor U24960 (N_24960,N_24378,N_24064);
xnor U24961 (N_24961,N_24372,N_24319);
and U24962 (N_24962,N_24043,N_24180);
nor U24963 (N_24963,N_24092,N_24426);
xor U24964 (N_24964,N_24324,N_24350);
xor U24965 (N_24965,N_24304,N_24252);
or U24966 (N_24966,N_24254,N_24401);
nor U24967 (N_24967,N_24368,N_24144);
nand U24968 (N_24968,N_24117,N_24351);
nor U24969 (N_24969,N_24168,N_24041);
xor U24970 (N_24970,N_24389,N_24215);
and U24971 (N_24971,N_24233,N_24070);
or U24972 (N_24972,N_24399,N_24436);
nor U24973 (N_24973,N_24262,N_24373);
and U24974 (N_24974,N_24252,N_24163);
nand U24975 (N_24975,N_24379,N_24013);
and U24976 (N_24976,N_24247,N_24161);
or U24977 (N_24977,N_24421,N_24460);
nor U24978 (N_24978,N_24441,N_24065);
xnor U24979 (N_24979,N_24199,N_24246);
xor U24980 (N_24980,N_24413,N_24164);
nor U24981 (N_24981,N_24423,N_24381);
nor U24982 (N_24982,N_24261,N_24262);
nand U24983 (N_24983,N_24068,N_24008);
nor U24984 (N_24984,N_24065,N_24006);
xor U24985 (N_24985,N_24281,N_24054);
xor U24986 (N_24986,N_24341,N_24285);
nor U24987 (N_24987,N_24393,N_24187);
or U24988 (N_24988,N_24179,N_24386);
or U24989 (N_24989,N_24472,N_24005);
xnor U24990 (N_24990,N_24182,N_24195);
xnor U24991 (N_24991,N_24157,N_24175);
nor U24992 (N_24992,N_24037,N_24161);
nor U24993 (N_24993,N_24231,N_24312);
or U24994 (N_24994,N_24262,N_24485);
xnor U24995 (N_24995,N_24199,N_24498);
xnor U24996 (N_24996,N_24230,N_24043);
or U24997 (N_24997,N_24177,N_24381);
nor U24998 (N_24998,N_24239,N_24396);
xor U24999 (N_24999,N_24099,N_24438);
nand U25000 (N_25000,N_24703,N_24524);
and U25001 (N_25001,N_24827,N_24509);
xor U25002 (N_25002,N_24905,N_24987);
xnor U25003 (N_25003,N_24923,N_24896);
and U25004 (N_25004,N_24815,N_24969);
nor U25005 (N_25005,N_24714,N_24706);
nor U25006 (N_25006,N_24806,N_24548);
nor U25007 (N_25007,N_24661,N_24856);
or U25008 (N_25008,N_24971,N_24842);
and U25009 (N_25009,N_24704,N_24841);
xor U25010 (N_25010,N_24768,N_24824);
xor U25011 (N_25011,N_24745,N_24920);
and U25012 (N_25012,N_24958,N_24710);
nor U25013 (N_25013,N_24525,N_24775);
nor U25014 (N_25014,N_24630,N_24544);
nand U25015 (N_25015,N_24577,N_24879);
nand U25016 (N_25016,N_24594,N_24847);
or U25017 (N_25017,N_24926,N_24774);
xnor U25018 (N_25018,N_24501,N_24742);
nand U25019 (N_25019,N_24554,N_24688);
nor U25020 (N_25020,N_24946,N_24616);
xnor U25021 (N_25021,N_24904,N_24875);
and U25022 (N_25022,N_24508,N_24782);
xnor U25023 (N_25023,N_24981,N_24695);
and U25024 (N_25024,N_24826,N_24895);
or U25025 (N_25025,N_24683,N_24939);
or U25026 (N_25026,N_24729,N_24892);
nand U25027 (N_25027,N_24680,N_24913);
or U25028 (N_25028,N_24656,N_24897);
or U25029 (N_25029,N_24592,N_24919);
nand U25030 (N_25030,N_24511,N_24619);
and U25031 (N_25031,N_24655,N_24686);
xnor U25032 (N_25032,N_24870,N_24909);
nor U25033 (N_25033,N_24541,N_24528);
nor U25034 (N_25034,N_24907,N_24948);
nand U25035 (N_25035,N_24889,N_24522);
xnor U25036 (N_25036,N_24766,N_24860);
nand U25037 (N_25037,N_24823,N_24613);
and U25038 (N_25038,N_24581,N_24990);
nor U25039 (N_25039,N_24708,N_24821);
and U25040 (N_25040,N_24899,N_24657);
xnor U25041 (N_25041,N_24622,N_24790);
nor U25042 (N_25042,N_24550,N_24719);
nand U25043 (N_25043,N_24608,N_24781);
nor U25044 (N_25044,N_24574,N_24993);
or U25045 (N_25045,N_24685,N_24831);
xnor U25046 (N_25046,N_24615,N_24961);
nor U25047 (N_25047,N_24644,N_24885);
and U25048 (N_25048,N_24694,N_24911);
or U25049 (N_25049,N_24994,N_24716);
nor U25050 (N_25050,N_24857,N_24957);
nand U25051 (N_25051,N_24829,N_24910);
nand U25052 (N_25052,N_24677,N_24898);
or U25053 (N_25053,N_24789,N_24506);
or U25054 (N_25054,N_24747,N_24967);
nor U25055 (N_25055,N_24908,N_24586);
or U25056 (N_25056,N_24974,N_24848);
and U25057 (N_25057,N_24549,N_24606);
nand U25058 (N_25058,N_24794,N_24835);
and U25059 (N_25059,N_24503,N_24759);
xnor U25060 (N_25060,N_24949,N_24873);
xnor U25061 (N_25061,N_24854,N_24855);
or U25062 (N_25062,N_24748,N_24998);
or U25063 (N_25063,N_24517,N_24669);
nor U25064 (N_25064,N_24725,N_24927);
nor U25065 (N_25065,N_24651,N_24798);
nor U25066 (N_25066,N_24846,N_24523);
nand U25067 (N_25067,N_24930,N_24746);
xor U25068 (N_25068,N_24894,N_24795);
nor U25069 (N_25069,N_24696,N_24991);
nor U25070 (N_25070,N_24880,N_24738);
and U25071 (N_25071,N_24652,N_24721);
xnor U25072 (N_25072,N_24833,N_24972);
and U25073 (N_25073,N_24727,N_24646);
nor U25074 (N_25074,N_24955,N_24785);
or U25075 (N_25075,N_24647,N_24830);
nand U25076 (N_25076,N_24840,N_24876);
nor U25077 (N_25077,N_24807,N_24763);
nand U25078 (N_25078,N_24960,N_24845);
or U25079 (N_25079,N_24802,N_24893);
xor U25080 (N_25080,N_24772,N_24773);
and U25081 (N_25081,N_24822,N_24660);
or U25082 (N_25082,N_24954,N_24771);
nand U25083 (N_25083,N_24530,N_24617);
xnor U25084 (N_25084,N_24576,N_24862);
xnor U25085 (N_25085,N_24739,N_24610);
xor U25086 (N_25086,N_24874,N_24539);
xnor U25087 (N_25087,N_24755,N_24609);
nor U25088 (N_25088,N_24780,N_24736);
and U25089 (N_25089,N_24940,N_24596);
nor U25090 (N_25090,N_24836,N_24654);
nand U25091 (N_25091,N_24865,N_24565);
and U25092 (N_25092,N_24663,N_24935);
nor U25093 (N_25093,N_24881,N_24621);
or U25094 (N_25094,N_24784,N_24653);
xnor U25095 (N_25095,N_24963,N_24582);
nand U25096 (N_25096,N_24546,N_24984);
nand U25097 (N_25097,N_24666,N_24510);
xnor U25098 (N_25098,N_24545,N_24563);
nor U25099 (N_25099,N_24558,N_24850);
xnor U25100 (N_25100,N_24968,N_24891);
nand U25101 (N_25101,N_24741,N_24593);
nand U25102 (N_25102,N_24912,N_24816);
nor U25103 (N_25103,N_24752,N_24733);
nor U25104 (N_25104,N_24579,N_24867);
xor U25105 (N_25105,N_24534,N_24635);
xnor U25106 (N_25106,N_24602,N_24995);
or U25107 (N_25107,N_24561,N_24702);
nor U25108 (N_25108,N_24849,N_24753);
nand U25109 (N_25109,N_24637,N_24571);
xor U25110 (N_25110,N_24864,N_24756);
or U25111 (N_25111,N_24884,N_24769);
xnor U25112 (N_25112,N_24735,N_24730);
nand U25113 (N_25113,N_24888,N_24671);
nor U25114 (N_25114,N_24591,N_24814);
nand U25115 (N_25115,N_24679,N_24731);
or U25116 (N_25116,N_24760,N_24743);
nand U25117 (N_25117,N_24925,N_24595);
nand U25118 (N_25118,N_24690,N_24882);
or U25119 (N_25119,N_24504,N_24744);
or U25120 (N_25120,N_24783,N_24623);
nor U25121 (N_25121,N_24877,N_24985);
xor U25122 (N_25122,N_24953,N_24700);
nand U25123 (N_25123,N_24667,N_24723);
and U25124 (N_25124,N_24754,N_24917);
and U25125 (N_25125,N_24650,N_24749);
and U25126 (N_25126,N_24761,N_24553);
nor U25127 (N_25127,N_24936,N_24997);
and U25128 (N_25128,N_24639,N_24628);
and U25129 (N_25129,N_24793,N_24536);
nand U25130 (N_25130,N_24964,N_24674);
nor U25131 (N_25131,N_24612,N_24705);
and U25132 (N_25132,N_24989,N_24810);
nand U25133 (N_25133,N_24914,N_24799);
xnor U25134 (N_25134,N_24776,N_24934);
or U25135 (N_25135,N_24600,N_24531);
nand U25136 (N_25136,N_24871,N_24668);
nor U25137 (N_25137,N_24691,N_24859);
nand U25138 (N_25138,N_24529,N_24804);
xnor U25139 (N_25139,N_24812,N_24540);
xor U25140 (N_25140,N_24980,N_24979);
or U25141 (N_25141,N_24779,N_24931);
xor U25142 (N_25142,N_24502,N_24765);
or U25143 (N_25143,N_24662,N_24924);
or U25144 (N_25144,N_24570,N_24797);
nand U25145 (N_25145,N_24603,N_24901);
nand U25146 (N_25146,N_24518,N_24777);
nor U25147 (N_25147,N_24868,N_24869);
nand U25148 (N_25148,N_24689,N_24599);
nor U25149 (N_25149,N_24838,N_24672);
nor U25150 (N_25150,N_24767,N_24751);
nand U25151 (N_25151,N_24809,N_24638);
xnor U25152 (N_25152,N_24837,N_24538);
nor U25153 (N_25153,N_24801,N_24986);
nand U25154 (N_25154,N_24658,N_24861);
nand U25155 (N_25155,N_24813,N_24915);
or U25156 (N_25156,N_24645,N_24734);
and U25157 (N_25157,N_24872,N_24665);
and U25158 (N_25158,N_24852,N_24629);
xor U25159 (N_25159,N_24684,N_24559);
xnor U25160 (N_25160,N_24693,N_24516);
and U25161 (N_25161,N_24718,N_24520);
nor U25162 (N_25162,N_24641,N_24555);
xor U25163 (N_25163,N_24547,N_24726);
or U25164 (N_25164,N_24999,N_24944);
nor U25165 (N_25165,N_24604,N_24560);
xor U25166 (N_25166,N_24977,N_24933);
nand U25167 (N_25167,N_24687,N_24699);
nor U25168 (N_25168,N_24675,N_24803);
nand U25169 (N_25169,N_24648,N_24631);
or U25170 (N_25170,N_24601,N_24973);
nand U25171 (N_25171,N_24519,N_24620);
xnor U25172 (N_25172,N_24614,N_24659);
xor U25173 (N_25173,N_24942,N_24758);
xor U25174 (N_25174,N_24634,N_24642);
and U25175 (N_25175,N_24791,N_24922);
and U25176 (N_25176,N_24740,N_24982);
xor U25177 (N_25177,N_24632,N_24858);
nand U25178 (N_25178,N_24737,N_24527);
xor U25179 (N_25179,N_24952,N_24564);
nor U25180 (N_25180,N_24692,N_24572);
and U25181 (N_25181,N_24588,N_24866);
nand U25182 (N_25182,N_24786,N_24578);
and U25183 (N_25183,N_24978,N_24764);
and U25184 (N_25184,N_24788,N_24724);
nand U25185 (N_25185,N_24863,N_24720);
and U25186 (N_25186,N_24607,N_24844);
and U25187 (N_25187,N_24521,N_24945);
nand U25188 (N_25188,N_24513,N_24711);
xor U25189 (N_25189,N_24573,N_24543);
nor U25190 (N_25190,N_24805,N_24636);
nor U25191 (N_25191,N_24757,N_24698);
nand U25192 (N_25192,N_24817,N_24825);
xnor U25193 (N_25193,N_24562,N_24713);
nand U25194 (N_25194,N_24992,N_24681);
nor U25195 (N_25195,N_24903,N_24682);
and U25196 (N_25196,N_24937,N_24928);
nor U25197 (N_25197,N_24709,N_24983);
xor U25198 (N_25198,N_24505,N_24787);
nand U25199 (N_25199,N_24770,N_24959);
and U25200 (N_25200,N_24728,N_24938);
nor U25201 (N_25201,N_24537,N_24878);
or U25202 (N_25202,N_24717,N_24569);
nor U25203 (N_25203,N_24587,N_24929);
xnor U25204 (N_25204,N_24673,N_24951);
and U25205 (N_25205,N_24811,N_24932);
nor U25206 (N_25206,N_24918,N_24828);
and U25207 (N_25207,N_24512,N_24567);
and U25208 (N_25208,N_24584,N_24839);
and U25209 (N_25209,N_24568,N_24526);
nand U25210 (N_25210,N_24970,N_24598);
or U25211 (N_25211,N_24800,N_24843);
nand U25212 (N_25212,N_24966,N_24834);
xnor U25213 (N_25213,N_24883,N_24916);
nor U25214 (N_25214,N_24965,N_24627);
xor U25215 (N_25215,N_24900,N_24590);
and U25216 (N_25216,N_24625,N_24583);
xnor U25217 (N_25217,N_24976,N_24808);
or U25218 (N_25218,N_24626,N_24886);
or U25219 (N_25219,N_24853,N_24796);
and U25220 (N_25220,N_24988,N_24676);
nor U25221 (N_25221,N_24832,N_24552);
or U25222 (N_25222,N_24542,N_24697);
or U25223 (N_25223,N_24575,N_24611);
and U25224 (N_25224,N_24678,N_24643);
or U25225 (N_25225,N_24566,N_24722);
xor U25226 (N_25226,N_24640,N_24941);
xnor U25227 (N_25227,N_24996,N_24818);
nand U25228 (N_25228,N_24921,N_24515);
xnor U25229 (N_25229,N_24580,N_24902);
or U25230 (N_25230,N_24605,N_24649);
xnor U25231 (N_25231,N_24732,N_24819);
nor U25232 (N_25232,N_24633,N_24585);
nand U25233 (N_25233,N_24950,N_24624);
or U25234 (N_25234,N_24551,N_24906);
nand U25235 (N_25235,N_24589,N_24507);
and U25236 (N_25236,N_24500,N_24947);
xor U25237 (N_25237,N_24943,N_24851);
or U25238 (N_25238,N_24701,N_24887);
and U25239 (N_25239,N_24715,N_24750);
and U25240 (N_25240,N_24956,N_24778);
and U25241 (N_25241,N_24532,N_24762);
nand U25242 (N_25242,N_24962,N_24535);
xor U25243 (N_25243,N_24597,N_24556);
nor U25244 (N_25244,N_24664,N_24670);
xnor U25245 (N_25245,N_24975,N_24533);
nand U25246 (N_25246,N_24514,N_24707);
or U25247 (N_25247,N_24712,N_24792);
and U25248 (N_25248,N_24557,N_24890);
xnor U25249 (N_25249,N_24820,N_24618);
nor U25250 (N_25250,N_24846,N_24698);
nor U25251 (N_25251,N_24503,N_24858);
nand U25252 (N_25252,N_24557,N_24727);
or U25253 (N_25253,N_24852,N_24536);
xnor U25254 (N_25254,N_24965,N_24863);
nor U25255 (N_25255,N_24685,N_24706);
xor U25256 (N_25256,N_24953,N_24558);
xor U25257 (N_25257,N_24715,N_24646);
and U25258 (N_25258,N_24834,N_24901);
or U25259 (N_25259,N_24876,N_24529);
nor U25260 (N_25260,N_24998,N_24941);
nand U25261 (N_25261,N_24865,N_24801);
xor U25262 (N_25262,N_24847,N_24581);
nand U25263 (N_25263,N_24546,N_24774);
and U25264 (N_25264,N_24680,N_24651);
and U25265 (N_25265,N_24886,N_24901);
nor U25266 (N_25266,N_24505,N_24617);
or U25267 (N_25267,N_24691,N_24897);
and U25268 (N_25268,N_24709,N_24792);
nor U25269 (N_25269,N_24588,N_24582);
xnor U25270 (N_25270,N_24558,N_24845);
nor U25271 (N_25271,N_24805,N_24810);
and U25272 (N_25272,N_24622,N_24772);
nand U25273 (N_25273,N_24609,N_24954);
and U25274 (N_25274,N_24954,N_24910);
xor U25275 (N_25275,N_24606,N_24582);
nor U25276 (N_25276,N_24793,N_24646);
nand U25277 (N_25277,N_24962,N_24631);
nor U25278 (N_25278,N_24525,N_24633);
and U25279 (N_25279,N_24502,N_24947);
or U25280 (N_25280,N_24978,N_24866);
nand U25281 (N_25281,N_24595,N_24618);
xnor U25282 (N_25282,N_24678,N_24659);
nand U25283 (N_25283,N_24900,N_24774);
or U25284 (N_25284,N_24794,N_24613);
nand U25285 (N_25285,N_24635,N_24554);
xor U25286 (N_25286,N_24634,N_24553);
nand U25287 (N_25287,N_24912,N_24594);
and U25288 (N_25288,N_24869,N_24561);
nor U25289 (N_25289,N_24699,N_24993);
or U25290 (N_25290,N_24824,N_24668);
and U25291 (N_25291,N_24740,N_24630);
nor U25292 (N_25292,N_24909,N_24723);
and U25293 (N_25293,N_24948,N_24974);
nor U25294 (N_25294,N_24641,N_24800);
and U25295 (N_25295,N_24748,N_24882);
and U25296 (N_25296,N_24603,N_24753);
nand U25297 (N_25297,N_24949,N_24975);
nand U25298 (N_25298,N_24602,N_24700);
nor U25299 (N_25299,N_24644,N_24910);
nand U25300 (N_25300,N_24940,N_24642);
nor U25301 (N_25301,N_24927,N_24578);
and U25302 (N_25302,N_24555,N_24926);
nand U25303 (N_25303,N_24598,N_24787);
and U25304 (N_25304,N_24752,N_24518);
nand U25305 (N_25305,N_24597,N_24922);
nor U25306 (N_25306,N_24912,N_24715);
and U25307 (N_25307,N_24535,N_24903);
or U25308 (N_25308,N_24928,N_24517);
or U25309 (N_25309,N_24773,N_24903);
or U25310 (N_25310,N_24704,N_24648);
xnor U25311 (N_25311,N_24509,N_24693);
nor U25312 (N_25312,N_24990,N_24864);
and U25313 (N_25313,N_24822,N_24610);
nand U25314 (N_25314,N_24844,N_24553);
and U25315 (N_25315,N_24873,N_24846);
nor U25316 (N_25316,N_24574,N_24716);
and U25317 (N_25317,N_24568,N_24929);
nor U25318 (N_25318,N_24658,N_24617);
and U25319 (N_25319,N_24632,N_24631);
xor U25320 (N_25320,N_24501,N_24666);
xnor U25321 (N_25321,N_24783,N_24603);
or U25322 (N_25322,N_24755,N_24915);
and U25323 (N_25323,N_24964,N_24514);
xor U25324 (N_25324,N_24606,N_24862);
and U25325 (N_25325,N_24869,N_24989);
xnor U25326 (N_25326,N_24522,N_24891);
xnor U25327 (N_25327,N_24824,N_24877);
nand U25328 (N_25328,N_24687,N_24751);
and U25329 (N_25329,N_24899,N_24913);
xor U25330 (N_25330,N_24571,N_24972);
or U25331 (N_25331,N_24611,N_24641);
or U25332 (N_25332,N_24653,N_24534);
nand U25333 (N_25333,N_24820,N_24692);
nor U25334 (N_25334,N_24647,N_24664);
or U25335 (N_25335,N_24943,N_24890);
nor U25336 (N_25336,N_24719,N_24906);
or U25337 (N_25337,N_24692,N_24906);
xnor U25338 (N_25338,N_24687,N_24863);
or U25339 (N_25339,N_24676,N_24510);
xor U25340 (N_25340,N_24512,N_24824);
nor U25341 (N_25341,N_24844,N_24953);
or U25342 (N_25342,N_24980,N_24562);
and U25343 (N_25343,N_24568,N_24914);
xor U25344 (N_25344,N_24933,N_24930);
and U25345 (N_25345,N_24759,N_24858);
xnor U25346 (N_25346,N_24794,N_24649);
nand U25347 (N_25347,N_24783,N_24957);
and U25348 (N_25348,N_24915,N_24789);
or U25349 (N_25349,N_24917,N_24727);
nand U25350 (N_25350,N_24781,N_24558);
nor U25351 (N_25351,N_24550,N_24897);
and U25352 (N_25352,N_24622,N_24799);
xnor U25353 (N_25353,N_24578,N_24652);
xnor U25354 (N_25354,N_24594,N_24918);
and U25355 (N_25355,N_24825,N_24930);
xnor U25356 (N_25356,N_24561,N_24537);
and U25357 (N_25357,N_24672,N_24633);
or U25358 (N_25358,N_24617,N_24908);
nor U25359 (N_25359,N_24995,N_24714);
and U25360 (N_25360,N_24680,N_24995);
or U25361 (N_25361,N_24603,N_24830);
and U25362 (N_25362,N_24964,N_24967);
and U25363 (N_25363,N_24938,N_24794);
nand U25364 (N_25364,N_24898,N_24581);
or U25365 (N_25365,N_24924,N_24690);
nand U25366 (N_25366,N_24611,N_24910);
and U25367 (N_25367,N_24810,N_24839);
and U25368 (N_25368,N_24543,N_24764);
nand U25369 (N_25369,N_24650,N_24824);
nand U25370 (N_25370,N_24517,N_24575);
nor U25371 (N_25371,N_24952,N_24779);
nand U25372 (N_25372,N_24957,N_24688);
nor U25373 (N_25373,N_24888,N_24768);
and U25374 (N_25374,N_24670,N_24762);
nand U25375 (N_25375,N_24924,N_24951);
and U25376 (N_25376,N_24583,N_24669);
nor U25377 (N_25377,N_24799,N_24944);
and U25378 (N_25378,N_24869,N_24670);
or U25379 (N_25379,N_24656,N_24678);
and U25380 (N_25380,N_24980,N_24913);
nand U25381 (N_25381,N_24682,N_24920);
nor U25382 (N_25382,N_24792,N_24904);
xor U25383 (N_25383,N_24640,N_24835);
and U25384 (N_25384,N_24934,N_24858);
nand U25385 (N_25385,N_24615,N_24635);
nor U25386 (N_25386,N_24731,N_24718);
xnor U25387 (N_25387,N_24867,N_24950);
nor U25388 (N_25388,N_24796,N_24870);
nor U25389 (N_25389,N_24503,N_24830);
nor U25390 (N_25390,N_24998,N_24608);
nand U25391 (N_25391,N_24519,N_24710);
nor U25392 (N_25392,N_24768,N_24872);
nand U25393 (N_25393,N_24727,N_24608);
or U25394 (N_25394,N_24862,N_24802);
nor U25395 (N_25395,N_24876,N_24992);
nand U25396 (N_25396,N_24925,N_24789);
nand U25397 (N_25397,N_24770,N_24733);
nor U25398 (N_25398,N_24688,N_24840);
xnor U25399 (N_25399,N_24892,N_24513);
nand U25400 (N_25400,N_24542,N_24536);
nor U25401 (N_25401,N_24906,N_24954);
xor U25402 (N_25402,N_24620,N_24962);
nor U25403 (N_25403,N_24711,N_24818);
nand U25404 (N_25404,N_24867,N_24832);
and U25405 (N_25405,N_24831,N_24543);
nor U25406 (N_25406,N_24795,N_24578);
nor U25407 (N_25407,N_24620,N_24740);
or U25408 (N_25408,N_24965,N_24761);
and U25409 (N_25409,N_24753,N_24766);
and U25410 (N_25410,N_24927,N_24712);
nor U25411 (N_25411,N_24618,N_24715);
or U25412 (N_25412,N_24647,N_24766);
nor U25413 (N_25413,N_24595,N_24940);
nor U25414 (N_25414,N_24898,N_24538);
nand U25415 (N_25415,N_24645,N_24819);
xor U25416 (N_25416,N_24623,N_24515);
nor U25417 (N_25417,N_24731,N_24751);
and U25418 (N_25418,N_24615,N_24654);
or U25419 (N_25419,N_24684,N_24653);
or U25420 (N_25420,N_24972,N_24876);
or U25421 (N_25421,N_24765,N_24573);
xnor U25422 (N_25422,N_24577,N_24828);
or U25423 (N_25423,N_24794,N_24973);
or U25424 (N_25424,N_24508,N_24968);
or U25425 (N_25425,N_24575,N_24727);
nor U25426 (N_25426,N_24796,N_24530);
nand U25427 (N_25427,N_24873,N_24996);
nor U25428 (N_25428,N_24906,N_24912);
and U25429 (N_25429,N_24654,N_24552);
or U25430 (N_25430,N_24519,N_24704);
or U25431 (N_25431,N_24854,N_24686);
nor U25432 (N_25432,N_24663,N_24636);
xnor U25433 (N_25433,N_24894,N_24917);
or U25434 (N_25434,N_24845,N_24641);
nand U25435 (N_25435,N_24697,N_24983);
nand U25436 (N_25436,N_24610,N_24595);
and U25437 (N_25437,N_24927,N_24813);
xor U25438 (N_25438,N_24699,N_24579);
xor U25439 (N_25439,N_24803,N_24865);
xor U25440 (N_25440,N_24940,N_24593);
nand U25441 (N_25441,N_24538,N_24993);
nor U25442 (N_25442,N_24677,N_24819);
xor U25443 (N_25443,N_24618,N_24869);
nand U25444 (N_25444,N_24576,N_24801);
nor U25445 (N_25445,N_24853,N_24700);
nor U25446 (N_25446,N_24911,N_24981);
xor U25447 (N_25447,N_24531,N_24666);
or U25448 (N_25448,N_24610,N_24527);
nand U25449 (N_25449,N_24547,N_24687);
nand U25450 (N_25450,N_24924,N_24767);
nand U25451 (N_25451,N_24715,N_24526);
nand U25452 (N_25452,N_24614,N_24600);
nand U25453 (N_25453,N_24810,N_24737);
and U25454 (N_25454,N_24846,N_24983);
xnor U25455 (N_25455,N_24840,N_24998);
and U25456 (N_25456,N_24767,N_24987);
nor U25457 (N_25457,N_24860,N_24981);
nand U25458 (N_25458,N_24530,N_24585);
nor U25459 (N_25459,N_24791,N_24746);
or U25460 (N_25460,N_24907,N_24872);
nor U25461 (N_25461,N_24756,N_24663);
nand U25462 (N_25462,N_24837,N_24918);
xor U25463 (N_25463,N_24682,N_24566);
nor U25464 (N_25464,N_24527,N_24758);
nand U25465 (N_25465,N_24918,N_24576);
or U25466 (N_25466,N_24856,N_24857);
or U25467 (N_25467,N_24806,N_24553);
nand U25468 (N_25468,N_24705,N_24992);
and U25469 (N_25469,N_24672,N_24688);
nor U25470 (N_25470,N_24612,N_24901);
or U25471 (N_25471,N_24790,N_24555);
xnor U25472 (N_25472,N_24850,N_24653);
nor U25473 (N_25473,N_24790,N_24854);
nor U25474 (N_25474,N_24948,N_24831);
nor U25475 (N_25475,N_24656,N_24571);
nor U25476 (N_25476,N_24605,N_24930);
xor U25477 (N_25477,N_24749,N_24561);
xor U25478 (N_25478,N_24931,N_24557);
xor U25479 (N_25479,N_24853,N_24530);
xor U25480 (N_25480,N_24809,N_24745);
nor U25481 (N_25481,N_24515,N_24697);
nand U25482 (N_25482,N_24668,N_24607);
and U25483 (N_25483,N_24571,N_24699);
and U25484 (N_25484,N_24784,N_24932);
nor U25485 (N_25485,N_24959,N_24843);
nor U25486 (N_25486,N_24899,N_24682);
nand U25487 (N_25487,N_24562,N_24778);
xnor U25488 (N_25488,N_24720,N_24612);
and U25489 (N_25489,N_24857,N_24815);
xor U25490 (N_25490,N_24637,N_24511);
or U25491 (N_25491,N_24682,N_24660);
nand U25492 (N_25492,N_24968,N_24788);
nand U25493 (N_25493,N_24596,N_24706);
xor U25494 (N_25494,N_24826,N_24974);
and U25495 (N_25495,N_24667,N_24814);
nand U25496 (N_25496,N_24558,N_24924);
and U25497 (N_25497,N_24644,N_24673);
nor U25498 (N_25498,N_24900,N_24794);
xnor U25499 (N_25499,N_24581,N_24530);
nand U25500 (N_25500,N_25405,N_25462);
xor U25501 (N_25501,N_25351,N_25224);
and U25502 (N_25502,N_25311,N_25061);
xnor U25503 (N_25503,N_25295,N_25360);
and U25504 (N_25504,N_25208,N_25085);
nor U25505 (N_25505,N_25017,N_25095);
nor U25506 (N_25506,N_25452,N_25410);
or U25507 (N_25507,N_25358,N_25094);
xnor U25508 (N_25508,N_25156,N_25484);
or U25509 (N_25509,N_25449,N_25428);
and U25510 (N_25510,N_25315,N_25498);
nand U25511 (N_25511,N_25236,N_25263);
xnor U25512 (N_25512,N_25005,N_25468);
nand U25513 (N_25513,N_25268,N_25004);
or U25514 (N_25514,N_25496,N_25341);
and U25515 (N_25515,N_25161,N_25321);
nand U25516 (N_25516,N_25026,N_25016);
nor U25517 (N_25517,N_25381,N_25011);
nor U25518 (N_25518,N_25261,N_25255);
and U25519 (N_25519,N_25160,N_25007);
or U25520 (N_25520,N_25336,N_25273);
xnor U25521 (N_25521,N_25097,N_25038);
or U25522 (N_25522,N_25416,N_25418);
nand U25523 (N_25523,N_25213,N_25349);
or U25524 (N_25524,N_25362,N_25251);
xnor U25525 (N_25525,N_25066,N_25126);
nor U25526 (N_25526,N_25434,N_25404);
or U25527 (N_25527,N_25361,N_25426);
nand U25528 (N_25528,N_25194,N_25390);
nand U25529 (N_25529,N_25317,N_25271);
nand U25530 (N_25530,N_25267,N_25045);
and U25531 (N_25531,N_25483,N_25327);
nand U25532 (N_25532,N_25056,N_25240);
or U25533 (N_25533,N_25074,N_25403);
xor U25534 (N_25534,N_25128,N_25103);
or U25535 (N_25535,N_25367,N_25154);
xnor U25536 (N_25536,N_25386,N_25046);
and U25537 (N_25537,N_25306,N_25117);
xnor U25538 (N_25538,N_25125,N_25116);
nand U25539 (N_25539,N_25150,N_25185);
nor U25540 (N_25540,N_25423,N_25174);
and U25541 (N_25541,N_25137,N_25466);
or U25542 (N_25542,N_25412,N_25018);
or U25543 (N_25543,N_25356,N_25009);
and U25544 (N_25544,N_25297,N_25371);
nand U25545 (N_25545,N_25107,N_25312);
nand U25546 (N_25546,N_25051,N_25221);
xnor U25547 (N_25547,N_25425,N_25023);
xor U25548 (N_25548,N_25069,N_25435);
or U25549 (N_25549,N_25063,N_25122);
xor U25550 (N_25550,N_25298,N_25451);
nand U25551 (N_25551,N_25021,N_25269);
xor U25552 (N_25552,N_25422,N_25303);
and U25553 (N_25553,N_25214,N_25012);
xnor U25554 (N_25554,N_25165,N_25256);
and U25555 (N_25555,N_25391,N_25470);
and U25556 (N_25556,N_25060,N_25393);
nor U25557 (N_25557,N_25233,N_25415);
and U25558 (N_25558,N_25022,N_25105);
or U25559 (N_25559,N_25257,N_25417);
nor U25560 (N_25560,N_25474,N_25025);
or U25561 (N_25561,N_25197,N_25278);
or U25562 (N_25562,N_25379,N_25402);
xor U25563 (N_25563,N_25162,N_25326);
and U25564 (N_25564,N_25033,N_25102);
xor U25565 (N_25565,N_25175,N_25438);
or U25566 (N_25566,N_25072,N_25200);
nand U25567 (N_25567,N_25433,N_25274);
nor U25568 (N_25568,N_25293,N_25113);
nand U25569 (N_25569,N_25247,N_25226);
xor U25570 (N_25570,N_25409,N_25280);
nor U25571 (N_25571,N_25186,N_25169);
nor U25572 (N_25572,N_25461,N_25210);
xor U25573 (N_25573,N_25333,N_25147);
xor U25574 (N_25574,N_25318,N_25028);
or U25575 (N_25575,N_25444,N_25395);
nor U25576 (N_25576,N_25291,N_25345);
and U25577 (N_25577,N_25244,N_25387);
nand U25578 (N_25578,N_25181,N_25075);
or U25579 (N_25579,N_25058,N_25490);
xor U25580 (N_25580,N_25144,N_25164);
nand U25581 (N_25581,N_25302,N_25220);
or U25582 (N_25582,N_25299,N_25335);
nand U25583 (N_25583,N_25237,N_25043);
nand U25584 (N_25584,N_25231,N_25006);
and U25585 (N_25585,N_25266,N_25467);
xnor U25586 (N_25586,N_25471,N_25301);
nand U25587 (N_25587,N_25348,N_25152);
xor U25588 (N_25588,N_25448,N_25472);
nor U25589 (N_25589,N_25114,N_25119);
or U25590 (N_25590,N_25290,N_25440);
or U25591 (N_25591,N_25173,N_25049);
xnor U25592 (N_25592,N_25133,N_25222);
nor U25593 (N_25593,N_25101,N_25129);
nand U25594 (N_25594,N_25457,N_25041);
xor U25595 (N_25595,N_25488,N_25053);
or U25596 (N_25596,N_25157,N_25242);
and U25597 (N_25597,N_25482,N_25453);
or U25598 (N_25598,N_25248,N_25149);
nand U25599 (N_25599,N_25316,N_25190);
xor U25600 (N_25600,N_25218,N_25464);
or U25601 (N_25601,N_25239,N_25437);
xor U25602 (N_25602,N_25040,N_25037);
and U25603 (N_25603,N_25146,N_25365);
xor U25604 (N_25604,N_25459,N_25332);
xnor U25605 (N_25605,N_25188,N_25115);
or U25606 (N_25606,N_25153,N_25491);
or U25607 (N_25607,N_25486,N_25091);
or U25608 (N_25608,N_25187,N_25065);
or U25609 (N_25609,N_25118,N_25143);
nor U25610 (N_25610,N_25087,N_25343);
xnor U25611 (N_25611,N_25401,N_25176);
nand U25612 (N_25612,N_25195,N_25347);
xor U25613 (N_25613,N_25110,N_25155);
nand U25614 (N_25614,N_25008,N_25178);
and U25615 (N_25615,N_25229,N_25480);
nor U25616 (N_25616,N_25396,N_25377);
xnor U25617 (N_25617,N_25414,N_25394);
xor U25618 (N_25618,N_25071,N_25436);
nand U25619 (N_25619,N_25177,N_25346);
or U25620 (N_25620,N_25015,N_25034);
and U25621 (N_25621,N_25003,N_25127);
and U25622 (N_25622,N_25215,N_25310);
nor U25623 (N_25623,N_25232,N_25262);
and U25624 (N_25624,N_25443,N_25424);
or U25625 (N_25625,N_25389,N_25198);
xnor U25626 (N_25626,N_25171,N_25324);
and U25627 (N_25627,N_25392,N_25182);
or U25628 (N_25628,N_25441,N_25052);
xor U25629 (N_25629,N_25294,N_25193);
nor U25630 (N_25630,N_25047,N_25132);
nand U25631 (N_25631,N_25179,N_25206);
nand U25632 (N_25632,N_25407,N_25477);
and U25633 (N_25633,N_25366,N_25265);
nand U25634 (N_25634,N_25427,N_25330);
or U25635 (N_25635,N_25319,N_25357);
or U25636 (N_25636,N_25442,N_25282);
and U25637 (N_25637,N_25070,N_25138);
nor U25638 (N_25638,N_25172,N_25429);
nor U25639 (N_25639,N_25339,N_25322);
and U25640 (N_25640,N_25277,N_25082);
nand U25641 (N_25641,N_25369,N_25399);
and U25642 (N_25642,N_25374,N_25002);
nand U25643 (N_25643,N_25245,N_25260);
xnor U25644 (N_25644,N_25227,N_25170);
or U25645 (N_25645,N_25090,N_25376);
nand U25646 (N_25646,N_25281,N_25373);
and U25647 (N_25647,N_25338,N_25064);
nand U25648 (N_25648,N_25201,N_25334);
nor U25649 (N_25649,N_25135,N_25305);
nand U25650 (N_25650,N_25100,N_25035);
or U25651 (N_25651,N_25272,N_25159);
xor U25652 (N_25652,N_25384,N_25406);
or U25653 (N_25653,N_25493,N_25411);
nand U25654 (N_25654,N_25039,N_25109);
and U25655 (N_25655,N_25032,N_25340);
and U25656 (N_25656,N_25130,N_25168);
xor U25657 (N_25657,N_25350,N_25455);
or U25658 (N_25658,N_25314,N_25142);
or U25659 (N_25659,N_25353,N_25495);
or U25660 (N_25660,N_25010,N_25059);
xnor U25661 (N_25661,N_25445,N_25104);
and U25662 (N_25662,N_25136,N_25275);
xor U25663 (N_25663,N_25238,N_25092);
nor U25664 (N_25664,N_25014,N_25355);
and U25665 (N_25665,N_25131,N_25029);
and U25666 (N_25666,N_25292,N_25096);
and U25667 (N_25667,N_25243,N_25079);
and U25668 (N_25668,N_25123,N_25383);
or U25669 (N_25669,N_25372,N_25432);
or U25670 (N_25670,N_25308,N_25254);
nand U25671 (N_25671,N_25469,N_25189);
nor U25672 (N_25672,N_25456,N_25027);
and U25673 (N_25673,N_25252,N_25344);
xnor U25674 (N_25674,N_25478,N_25329);
or U25675 (N_25675,N_25489,N_25458);
nand U25676 (N_25676,N_25228,N_25241);
nand U25677 (N_25677,N_25086,N_25283);
nand U25678 (N_25678,N_25364,N_25378);
nor U25679 (N_25679,N_25076,N_25108);
or U25680 (N_25680,N_25199,N_25419);
or U25681 (N_25681,N_25088,N_25259);
xnor U25682 (N_25682,N_25430,N_25068);
and U25683 (N_25683,N_25099,N_25209);
nor U25684 (N_25684,N_25447,N_25120);
xor U25685 (N_25685,N_25207,N_25098);
xor U25686 (N_25686,N_25180,N_25439);
xnor U25687 (N_25687,N_25288,N_25380);
nand U25688 (N_25688,N_25475,N_25300);
or U25689 (N_25689,N_25036,N_25368);
xor U25690 (N_25690,N_25212,N_25184);
or U25691 (N_25691,N_25078,N_25270);
and U25692 (N_25692,N_25205,N_25485);
nand U25693 (N_25693,N_25048,N_25492);
and U25694 (N_25694,N_25084,N_25320);
nand U25695 (N_25695,N_25134,N_25313);
or U25696 (N_25696,N_25001,N_25285);
nor U25697 (N_25697,N_25473,N_25323);
nand U25698 (N_25698,N_25494,N_25354);
nand U25699 (N_25699,N_25276,N_25225);
or U25700 (N_25700,N_25375,N_25158);
nor U25701 (N_25701,N_25309,N_25450);
nand U25702 (N_25702,N_25000,N_25287);
xor U25703 (N_25703,N_25141,N_25400);
xor U25704 (N_25704,N_25479,N_25286);
nor U25705 (N_25705,N_25055,N_25083);
or U25706 (N_25706,N_25081,N_25246);
and U25707 (N_25707,N_25408,N_25013);
and U25708 (N_25708,N_25499,N_25385);
nand U25709 (N_25709,N_25421,N_25235);
and U25710 (N_25710,N_25465,N_25454);
or U25711 (N_25711,N_25050,N_25163);
or U25712 (N_25712,N_25112,N_25121);
or U25713 (N_25713,N_25398,N_25420);
nor U25714 (N_25714,N_25019,N_25223);
xnor U25715 (N_25715,N_25284,N_25093);
nor U25716 (N_25716,N_25151,N_25382);
nor U25717 (N_25717,N_25089,N_25031);
and U25718 (N_25718,N_25148,N_25183);
and U25719 (N_25719,N_25062,N_25497);
xnor U25720 (N_25720,N_25397,N_25359);
nor U25721 (N_25721,N_25307,N_25073);
xnor U25722 (N_25722,N_25258,N_25044);
nor U25723 (N_25723,N_25211,N_25124);
xor U25724 (N_25724,N_25219,N_25325);
xor U25725 (N_25725,N_25352,N_25145);
xor U25726 (N_25726,N_25111,N_25140);
nand U25727 (N_25727,N_25413,N_25234);
and U25728 (N_25728,N_25264,N_25020);
xor U25729 (N_25729,N_25487,N_25106);
xor U25730 (N_25730,N_25388,N_25370);
nand U25731 (N_25731,N_25077,N_25030);
xor U25732 (N_25732,N_25217,N_25067);
nor U25733 (N_25733,N_25296,N_25139);
xnor U25734 (N_25734,N_25249,N_25481);
nor U25735 (N_25735,N_25331,N_25192);
or U25736 (N_25736,N_25080,N_25216);
or U25737 (N_25737,N_25253,N_25289);
nand U25738 (N_25738,N_25328,N_25204);
nand U25739 (N_25739,N_25054,N_25202);
or U25740 (N_25740,N_25250,N_25337);
nand U25741 (N_25741,N_25476,N_25431);
nand U25742 (N_25742,N_25446,N_25191);
or U25743 (N_25743,N_25024,N_25463);
nand U25744 (N_25744,N_25304,N_25203);
xnor U25745 (N_25745,N_25279,N_25167);
nand U25746 (N_25746,N_25460,N_25230);
or U25747 (N_25747,N_25057,N_25342);
nor U25748 (N_25748,N_25196,N_25166);
nor U25749 (N_25749,N_25042,N_25363);
xnor U25750 (N_25750,N_25440,N_25299);
or U25751 (N_25751,N_25314,N_25430);
nor U25752 (N_25752,N_25393,N_25225);
and U25753 (N_25753,N_25272,N_25449);
nor U25754 (N_25754,N_25436,N_25182);
xor U25755 (N_25755,N_25332,N_25116);
nand U25756 (N_25756,N_25151,N_25399);
nand U25757 (N_25757,N_25352,N_25182);
xnor U25758 (N_25758,N_25056,N_25434);
or U25759 (N_25759,N_25395,N_25138);
xor U25760 (N_25760,N_25375,N_25246);
or U25761 (N_25761,N_25146,N_25055);
nand U25762 (N_25762,N_25305,N_25023);
nor U25763 (N_25763,N_25405,N_25363);
or U25764 (N_25764,N_25022,N_25379);
and U25765 (N_25765,N_25053,N_25245);
or U25766 (N_25766,N_25322,N_25164);
nor U25767 (N_25767,N_25399,N_25164);
nor U25768 (N_25768,N_25193,N_25369);
and U25769 (N_25769,N_25279,N_25265);
and U25770 (N_25770,N_25478,N_25000);
and U25771 (N_25771,N_25428,N_25077);
and U25772 (N_25772,N_25187,N_25411);
xor U25773 (N_25773,N_25408,N_25360);
nand U25774 (N_25774,N_25467,N_25376);
xnor U25775 (N_25775,N_25349,N_25208);
xor U25776 (N_25776,N_25337,N_25207);
and U25777 (N_25777,N_25372,N_25391);
and U25778 (N_25778,N_25421,N_25124);
xor U25779 (N_25779,N_25028,N_25154);
nand U25780 (N_25780,N_25349,N_25378);
nor U25781 (N_25781,N_25160,N_25335);
xor U25782 (N_25782,N_25173,N_25455);
nor U25783 (N_25783,N_25308,N_25147);
nand U25784 (N_25784,N_25175,N_25402);
xor U25785 (N_25785,N_25142,N_25414);
nand U25786 (N_25786,N_25340,N_25424);
xnor U25787 (N_25787,N_25475,N_25046);
nand U25788 (N_25788,N_25471,N_25142);
or U25789 (N_25789,N_25175,N_25397);
and U25790 (N_25790,N_25434,N_25409);
nand U25791 (N_25791,N_25063,N_25218);
and U25792 (N_25792,N_25028,N_25450);
and U25793 (N_25793,N_25060,N_25053);
nand U25794 (N_25794,N_25447,N_25253);
or U25795 (N_25795,N_25177,N_25498);
nand U25796 (N_25796,N_25417,N_25180);
and U25797 (N_25797,N_25231,N_25299);
xnor U25798 (N_25798,N_25151,N_25437);
and U25799 (N_25799,N_25294,N_25464);
nor U25800 (N_25800,N_25355,N_25457);
and U25801 (N_25801,N_25117,N_25327);
xnor U25802 (N_25802,N_25178,N_25012);
or U25803 (N_25803,N_25039,N_25402);
xnor U25804 (N_25804,N_25339,N_25179);
xor U25805 (N_25805,N_25210,N_25135);
and U25806 (N_25806,N_25493,N_25220);
and U25807 (N_25807,N_25130,N_25266);
nand U25808 (N_25808,N_25186,N_25215);
nor U25809 (N_25809,N_25323,N_25053);
nand U25810 (N_25810,N_25440,N_25377);
nand U25811 (N_25811,N_25048,N_25092);
nor U25812 (N_25812,N_25103,N_25132);
nand U25813 (N_25813,N_25379,N_25481);
nand U25814 (N_25814,N_25233,N_25301);
nor U25815 (N_25815,N_25164,N_25077);
nand U25816 (N_25816,N_25251,N_25357);
and U25817 (N_25817,N_25285,N_25007);
nand U25818 (N_25818,N_25360,N_25057);
or U25819 (N_25819,N_25141,N_25486);
xor U25820 (N_25820,N_25436,N_25032);
and U25821 (N_25821,N_25111,N_25487);
or U25822 (N_25822,N_25367,N_25488);
xor U25823 (N_25823,N_25061,N_25342);
and U25824 (N_25824,N_25264,N_25324);
and U25825 (N_25825,N_25170,N_25361);
nor U25826 (N_25826,N_25360,N_25260);
nor U25827 (N_25827,N_25312,N_25273);
xor U25828 (N_25828,N_25356,N_25360);
xor U25829 (N_25829,N_25193,N_25018);
nor U25830 (N_25830,N_25282,N_25024);
xor U25831 (N_25831,N_25317,N_25395);
nand U25832 (N_25832,N_25057,N_25440);
nand U25833 (N_25833,N_25241,N_25433);
or U25834 (N_25834,N_25238,N_25173);
or U25835 (N_25835,N_25491,N_25039);
nand U25836 (N_25836,N_25171,N_25326);
or U25837 (N_25837,N_25440,N_25162);
or U25838 (N_25838,N_25383,N_25003);
nor U25839 (N_25839,N_25186,N_25489);
nor U25840 (N_25840,N_25087,N_25028);
or U25841 (N_25841,N_25006,N_25288);
xnor U25842 (N_25842,N_25170,N_25366);
nor U25843 (N_25843,N_25300,N_25019);
nand U25844 (N_25844,N_25063,N_25073);
nor U25845 (N_25845,N_25433,N_25109);
or U25846 (N_25846,N_25116,N_25193);
nor U25847 (N_25847,N_25034,N_25215);
xor U25848 (N_25848,N_25228,N_25206);
nand U25849 (N_25849,N_25140,N_25036);
and U25850 (N_25850,N_25465,N_25307);
and U25851 (N_25851,N_25031,N_25218);
nand U25852 (N_25852,N_25102,N_25198);
nor U25853 (N_25853,N_25497,N_25132);
nor U25854 (N_25854,N_25096,N_25257);
and U25855 (N_25855,N_25368,N_25093);
nor U25856 (N_25856,N_25115,N_25194);
nand U25857 (N_25857,N_25317,N_25218);
or U25858 (N_25858,N_25172,N_25173);
nand U25859 (N_25859,N_25474,N_25373);
or U25860 (N_25860,N_25409,N_25183);
and U25861 (N_25861,N_25192,N_25354);
and U25862 (N_25862,N_25286,N_25186);
xnor U25863 (N_25863,N_25234,N_25313);
nand U25864 (N_25864,N_25326,N_25319);
or U25865 (N_25865,N_25393,N_25249);
nand U25866 (N_25866,N_25249,N_25470);
and U25867 (N_25867,N_25057,N_25495);
nor U25868 (N_25868,N_25431,N_25076);
xnor U25869 (N_25869,N_25359,N_25470);
and U25870 (N_25870,N_25443,N_25447);
xnor U25871 (N_25871,N_25451,N_25159);
nand U25872 (N_25872,N_25243,N_25019);
and U25873 (N_25873,N_25225,N_25019);
xnor U25874 (N_25874,N_25043,N_25415);
xnor U25875 (N_25875,N_25216,N_25044);
nor U25876 (N_25876,N_25040,N_25374);
and U25877 (N_25877,N_25040,N_25117);
nand U25878 (N_25878,N_25265,N_25227);
or U25879 (N_25879,N_25279,N_25082);
or U25880 (N_25880,N_25371,N_25173);
xor U25881 (N_25881,N_25418,N_25077);
nand U25882 (N_25882,N_25309,N_25120);
xnor U25883 (N_25883,N_25021,N_25126);
nand U25884 (N_25884,N_25276,N_25041);
nor U25885 (N_25885,N_25310,N_25354);
xor U25886 (N_25886,N_25440,N_25247);
xnor U25887 (N_25887,N_25329,N_25455);
nor U25888 (N_25888,N_25154,N_25076);
nand U25889 (N_25889,N_25404,N_25092);
or U25890 (N_25890,N_25054,N_25445);
nor U25891 (N_25891,N_25318,N_25092);
and U25892 (N_25892,N_25047,N_25006);
nand U25893 (N_25893,N_25328,N_25172);
nor U25894 (N_25894,N_25079,N_25044);
or U25895 (N_25895,N_25422,N_25250);
or U25896 (N_25896,N_25451,N_25214);
xnor U25897 (N_25897,N_25016,N_25272);
xor U25898 (N_25898,N_25248,N_25169);
or U25899 (N_25899,N_25313,N_25367);
nand U25900 (N_25900,N_25087,N_25341);
nand U25901 (N_25901,N_25370,N_25166);
nor U25902 (N_25902,N_25295,N_25228);
nand U25903 (N_25903,N_25453,N_25392);
nand U25904 (N_25904,N_25166,N_25186);
and U25905 (N_25905,N_25274,N_25340);
xnor U25906 (N_25906,N_25273,N_25436);
or U25907 (N_25907,N_25019,N_25323);
and U25908 (N_25908,N_25054,N_25225);
and U25909 (N_25909,N_25231,N_25076);
xnor U25910 (N_25910,N_25450,N_25346);
and U25911 (N_25911,N_25213,N_25152);
or U25912 (N_25912,N_25216,N_25145);
or U25913 (N_25913,N_25323,N_25171);
or U25914 (N_25914,N_25004,N_25139);
or U25915 (N_25915,N_25413,N_25435);
nor U25916 (N_25916,N_25275,N_25354);
and U25917 (N_25917,N_25158,N_25311);
nor U25918 (N_25918,N_25056,N_25372);
nand U25919 (N_25919,N_25367,N_25077);
or U25920 (N_25920,N_25027,N_25134);
nand U25921 (N_25921,N_25144,N_25155);
nand U25922 (N_25922,N_25018,N_25192);
xor U25923 (N_25923,N_25028,N_25124);
nor U25924 (N_25924,N_25272,N_25181);
and U25925 (N_25925,N_25397,N_25268);
or U25926 (N_25926,N_25082,N_25151);
nand U25927 (N_25927,N_25312,N_25392);
and U25928 (N_25928,N_25285,N_25440);
nor U25929 (N_25929,N_25015,N_25243);
nor U25930 (N_25930,N_25393,N_25288);
nand U25931 (N_25931,N_25258,N_25249);
nor U25932 (N_25932,N_25085,N_25116);
nor U25933 (N_25933,N_25290,N_25135);
xnor U25934 (N_25934,N_25204,N_25232);
or U25935 (N_25935,N_25383,N_25312);
xnor U25936 (N_25936,N_25098,N_25283);
or U25937 (N_25937,N_25374,N_25209);
nand U25938 (N_25938,N_25381,N_25400);
and U25939 (N_25939,N_25192,N_25426);
or U25940 (N_25940,N_25463,N_25180);
nor U25941 (N_25941,N_25461,N_25320);
nor U25942 (N_25942,N_25482,N_25497);
xnor U25943 (N_25943,N_25245,N_25217);
xor U25944 (N_25944,N_25458,N_25012);
or U25945 (N_25945,N_25218,N_25324);
and U25946 (N_25946,N_25317,N_25143);
nor U25947 (N_25947,N_25426,N_25106);
nand U25948 (N_25948,N_25488,N_25034);
and U25949 (N_25949,N_25281,N_25328);
or U25950 (N_25950,N_25280,N_25375);
and U25951 (N_25951,N_25464,N_25444);
or U25952 (N_25952,N_25233,N_25010);
nand U25953 (N_25953,N_25097,N_25403);
and U25954 (N_25954,N_25269,N_25052);
nand U25955 (N_25955,N_25493,N_25430);
nand U25956 (N_25956,N_25331,N_25413);
xor U25957 (N_25957,N_25154,N_25062);
nand U25958 (N_25958,N_25100,N_25321);
nor U25959 (N_25959,N_25415,N_25050);
nor U25960 (N_25960,N_25023,N_25021);
xor U25961 (N_25961,N_25214,N_25061);
and U25962 (N_25962,N_25426,N_25451);
and U25963 (N_25963,N_25252,N_25074);
nand U25964 (N_25964,N_25325,N_25054);
xor U25965 (N_25965,N_25229,N_25471);
or U25966 (N_25966,N_25408,N_25071);
and U25967 (N_25967,N_25348,N_25496);
and U25968 (N_25968,N_25319,N_25455);
nand U25969 (N_25969,N_25158,N_25232);
xor U25970 (N_25970,N_25369,N_25123);
nor U25971 (N_25971,N_25259,N_25348);
nor U25972 (N_25972,N_25474,N_25141);
nand U25973 (N_25973,N_25008,N_25160);
nor U25974 (N_25974,N_25323,N_25400);
nand U25975 (N_25975,N_25004,N_25096);
or U25976 (N_25976,N_25460,N_25118);
nand U25977 (N_25977,N_25367,N_25358);
or U25978 (N_25978,N_25285,N_25059);
or U25979 (N_25979,N_25125,N_25146);
nand U25980 (N_25980,N_25168,N_25271);
nand U25981 (N_25981,N_25149,N_25217);
or U25982 (N_25982,N_25098,N_25051);
or U25983 (N_25983,N_25322,N_25155);
nor U25984 (N_25984,N_25140,N_25112);
nand U25985 (N_25985,N_25273,N_25478);
or U25986 (N_25986,N_25030,N_25061);
or U25987 (N_25987,N_25219,N_25320);
and U25988 (N_25988,N_25425,N_25191);
xnor U25989 (N_25989,N_25460,N_25486);
or U25990 (N_25990,N_25297,N_25004);
or U25991 (N_25991,N_25419,N_25415);
nor U25992 (N_25992,N_25105,N_25409);
xor U25993 (N_25993,N_25087,N_25330);
xor U25994 (N_25994,N_25223,N_25289);
nand U25995 (N_25995,N_25424,N_25136);
nor U25996 (N_25996,N_25384,N_25298);
or U25997 (N_25997,N_25422,N_25185);
nand U25998 (N_25998,N_25094,N_25356);
xor U25999 (N_25999,N_25271,N_25345);
nor U26000 (N_26000,N_25775,N_25862);
nor U26001 (N_26001,N_25705,N_25829);
or U26002 (N_26002,N_25575,N_25815);
or U26003 (N_26003,N_25939,N_25752);
nor U26004 (N_26004,N_25649,N_25986);
and U26005 (N_26005,N_25851,N_25956);
nand U26006 (N_26006,N_25620,N_25901);
and U26007 (N_26007,N_25626,N_25698);
xnor U26008 (N_26008,N_25671,N_25670);
or U26009 (N_26009,N_25544,N_25807);
nor U26010 (N_26010,N_25703,N_25571);
or U26011 (N_26011,N_25738,N_25716);
or U26012 (N_26012,N_25542,N_25714);
and U26013 (N_26013,N_25647,N_25658);
nand U26014 (N_26014,N_25609,N_25779);
nor U26015 (N_26015,N_25751,N_25713);
xor U26016 (N_26016,N_25577,N_25761);
nand U26017 (N_26017,N_25677,N_25992);
nor U26018 (N_26018,N_25699,N_25969);
or U26019 (N_26019,N_25744,N_25719);
nand U26020 (N_26020,N_25888,N_25919);
nor U26021 (N_26021,N_25799,N_25644);
nand U26022 (N_26022,N_25927,N_25616);
or U26023 (N_26023,N_25772,N_25790);
xnor U26024 (N_26024,N_25736,N_25514);
or U26025 (N_26025,N_25859,N_25911);
nor U26026 (N_26026,N_25686,N_25688);
or U26027 (N_26027,N_25740,N_25602);
nor U26028 (N_26028,N_25648,N_25586);
nor U26029 (N_26029,N_25906,N_25619);
nand U26030 (N_26030,N_25528,N_25836);
or U26031 (N_26031,N_25650,N_25569);
xnor U26032 (N_26032,N_25959,N_25946);
and U26033 (N_26033,N_25524,N_25666);
or U26034 (N_26034,N_25513,N_25603);
nor U26035 (N_26035,N_25595,N_25725);
or U26036 (N_26036,N_25947,N_25818);
nor U26037 (N_26037,N_25503,N_25838);
nand U26038 (N_26038,N_25983,N_25715);
and U26039 (N_26039,N_25564,N_25975);
nand U26040 (N_26040,N_25668,N_25885);
or U26041 (N_26041,N_25809,N_25876);
nand U26042 (N_26042,N_25904,N_25924);
xnor U26043 (N_26043,N_25872,N_25518);
xor U26044 (N_26044,N_25664,N_25590);
nor U26045 (N_26045,N_25676,N_25501);
nand U26046 (N_26046,N_25989,N_25627);
and U26047 (N_26047,N_25723,N_25731);
nand U26048 (N_26048,N_25584,N_25921);
or U26049 (N_26049,N_25696,N_25633);
nand U26050 (N_26050,N_25635,N_25573);
nand U26051 (N_26051,N_25733,N_25870);
xor U26052 (N_26052,N_25512,N_25599);
nand U26053 (N_26053,N_25553,N_25538);
nor U26054 (N_26054,N_25808,N_25614);
and U26055 (N_26055,N_25722,N_25707);
and U26056 (N_26056,N_25995,N_25690);
nor U26057 (N_26057,N_25708,N_25710);
and U26058 (N_26058,N_25773,N_25534);
nor U26059 (N_26059,N_25873,N_25550);
xor U26060 (N_26060,N_25653,N_25706);
nand U26061 (N_26061,N_25661,N_25629);
nand U26062 (N_26062,N_25516,N_25685);
nor U26063 (N_26063,N_25502,N_25759);
or U26064 (N_26064,N_25892,N_25895);
nor U26065 (N_26065,N_25780,N_25926);
xor U26066 (N_26066,N_25566,N_25925);
nor U26067 (N_26067,N_25543,N_25929);
or U26068 (N_26068,N_25540,N_25942);
and U26069 (N_26069,N_25672,N_25581);
nand U26070 (N_26070,N_25817,N_25900);
or U26071 (N_26071,N_25789,N_25585);
or U26072 (N_26072,N_25638,N_25621);
xor U26073 (N_26073,N_25902,N_25735);
nand U26074 (N_26074,N_25548,N_25941);
nor U26075 (N_26075,N_25847,N_25530);
nand U26076 (N_26076,N_25505,N_25898);
or U26077 (N_26077,N_25631,N_25563);
nand U26078 (N_26078,N_25674,N_25804);
and U26079 (N_26079,N_25966,N_25792);
and U26080 (N_26080,N_25718,N_25742);
nor U26081 (N_26081,N_25978,N_25541);
or U26082 (N_26082,N_25506,N_25565);
nor U26083 (N_26083,N_25755,N_25915);
xor U26084 (N_26084,N_25580,N_25729);
nor U26085 (N_26085,N_25673,N_25916);
nor U26086 (N_26086,N_25618,N_25850);
nand U26087 (N_26087,N_25861,N_25857);
or U26088 (N_26088,N_25652,N_25574);
nor U26089 (N_26089,N_25637,N_25726);
or U26090 (N_26090,N_25757,N_25810);
and U26091 (N_26091,N_25932,N_25520);
nor U26092 (N_26092,N_25656,N_25796);
or U26093 (N_26093,N_25979,N_25794);
xor U26094 (N_26094,N_25788,N_25568);
or U26095 (N_26095,N_25720,N_25903);
nor U26096 (N_26096,N_25785,N_25988);
or U26097 (N_26097,N_25824,N_25877);
nor U26098 (N_26098,N_25508,N_25546);
nor U26099 (N_26099,N_25665,N_25875);
or U26100 (N_26100,N_25519,N_25953);
and U26101 (N_26101,N_25869,N_25554);
xor U26102 (N_26102,N_25991,N_25591);
or U26103 (N_26103,N_25535,N_25611);
nor U26104 (N_26104,N_25774,N_25853);
xnor U26105 (N_26105,N_25545,N_25560);
nand U26106 (N_26106,N_25860,N_25766);
nand U26107 (N_26107,N_25971,N_25990);
or U26108 (N_26108,N_25555,N_25746);
or U26109 (N_26109,N_25593,N_25823);
xor U26110 (N_26110,N_25754,N_25643);
and U26111 (N_26111,N_25570,N_25782);
xor U26112 (N_26112,N_25878,N_25525);
nand U26113 (N_26113,N_25646,N_25852);
and U26114 (N_26114,N_25510,N_25727);
nor U26115 (N_26115,N_25747,N_25511);
nor U26116 (N_26116,N_25559,N_25930);
nand U26117 (N_26117,N_25753,N_25579);
or U26118 (N_26118,N_25880,N_25693);
nor U26119 (N_26119,N_25763,N_25748);
and U26120 (N_26120,N_25890,N_25689);
nor U26121 (N_26121,N_25702,N_25684);
or U26122 (N_26122,N_25899,N_25977);
or U26123 (N_26123,N_25613,N_25737);
nor U26124 (N_26124,N_25504,N_25783);
and U26125 (N_26125,N_25944,N_25871);
nand U26126 (N_26126,N_25604,N_25743);
nor U26127 (N_26127,N_25529,N_25515);
nand U26128 (N_26128,N_25660,N_25598);
or U26129 (N_26129,N_25655,N_25980);
and U26130 (N_26130,N_25937,N_25839);
or U26131 (N_26131,N_25695,N_25928);
and U26132 (N_26132,N_25549,N_25606);
nand U26133 (N_26133,N_25771,N_25517);
or U26134 (N_26134,N_25868,N_25526);
nand U26135 (N_26135,N_25617,N_25842);
xnor U26136 (N_26136,N_25965,N_25781);
nand U26137 (N_26137,N_25663,N_25894);
nand U26138 (N_26138,N_25678,N_25594);
nand U26139 (N_26139,N_25935,N_25667);
nand U26140 (N_26140,N_25547,N_25884);
nand U26141 (N_26141,N_25951,N_25657);
xor U26142 (N_26142,N_25500,N_25948);
nor U26143 (N_26143,N_25825,N_25957);
nand U26144 (N_26144,N_25578,N_25982);
nor U26145 (N_26145,N_25955,N_25837);
and U26146 (N_26146,N_25864,N_25700);
and U26147 (N_26147,N_25642,N_25634);
xor U26148 (N_26148,N_25840,N_25600);
xor U26149 (N_26149,N_25863,N_25879);
xnor U26150 (N_26150,N_25827,N_25784);
or U26151 (N_26151,N_25994,N_25572);
nor U26152 (N_26152,N_25622,N_25592);
nand U26153 (N_26153,N_25800,N_25522);
or U26154 (N_26154,N_25610,N_25596);
xor U26155 (N_26155,N_25931,N_25917);
nand U26156 (N_26156,N_25905,N_25625);
or U26157 (N_26157,N_25636,N_25694);
or U26158 (N_26158,N_25968,N_25812);
nand U26159 (N_26159,N_25587,N_25551);
or U26160 (N_26160,N_25765,N_25999);
xor U26161 (N_26161,N_25816,N_25583);
nor U26162 (N_26162,N_25552,N_25943);
or U26163 (N_26163,N_25639,N_25760);
xor U26164 (N_26164,N_25680,N_25820);
and U26165 (N_26165,N_25833,N_25527);
and U26166 (N_26166,N_25557,N_25628);
xor U26167 (N_26167,N_25612,N_25802);
nand U26168 (N_26168,N_25866,N_25770);
xor U26169 (N_26169,N_25981,N_25728);
and U26170 (N_26170,N_25669,N_25867);
xnor U26171 (N_26171,N_25974,N_25910);
and U26172 (N_26172,N_25961,N_25923);
nor U26173 (N_26173,N_25938,N_25821);
xnor U26174 (N_26174,N_25692,N_25972);
nor U26175 (N_26175,N_25848,N_25509);
or U26176 (N_26176,N_25806,N_25683);
or U26177 (N_26177,N_25576,N_25777);
or U26178 (N_26178,N_25960,N_25913);
nand U26179 (N_26179,N_25954,N_25828);
or U26180 (N_26180,N_25623,N_25768);
and U26181 (N_26181,N_25936,N_25856);
xnor U26182 (N_26182,N_25996,N_25918);
nor U26183 (N_26183,N_25608,N_25749);
xnor U26184 (N_26184,N_25797,N_25945);
nand U26185 (N_26185,N_25822,N_25963);
nor U26186 (N_26186,N_25597,N_25865);
xor U26187 (N_26187,N_25934,N_25819);
nand U26188 (N_26188,N_25734,N_25787);
or U26189 (N_26189,N_25745,N_25632);
and U26190 (N_26190,N_25897,N_25605);
nor U26191 (N_26191,N_25507,N_25843);
and U26192 (N_26192,N_25624,N_25691);
or U26193 (N_26193,N_25532,N_25835);
xnor U26194 (N_26194,N_25589,N_25793);
xnor U26195 (N_26195,N_25687,N_25970);
or U26196 (N_26196,N_25803,N_25531);
xnor U26197 (N_26197,N_25651,N_25539);
nor U26198 (N_26198,N_25854,N_25889);
or U26199 (N_26199,N_25940,N_25834);
nand U26200 (N_26200,N_25993,N_25830);
nand U26201 (N_26201,N_25952,N_25855);
nand U26202 (N_26202,N_25769,N_25778);
or U26203 (N_26203,N_25562,N_25813);
nor U26204 (N_26204,N_25607,N_25681);
nor U26205 (N_26205,N_25891,N_25641);
nand U26206 (N_26206,N_25582,N_25984);
xnor U26207 (N_26207,N_25558,N_25561);
xor U26208 (N_26208,N_25739,N_25767);
and U26209 (N_26209,N_25724,N_25887);
and U26210 (N_26210,N_25908,N_25764);
and U26211 (N_26211,N_25893,N_25533);
and U26212 (N_26212,N_25536,N_25758);
nand U26213 (N_26213,N_25909,N_25776);
or U26214 (N_26214,N_25985,N_25659);
or U26215 (N_26215,N_25615,N_25814);
xnor U26216 (N_26216,N_25973,N_25730);
xnor U26217 (N_26217,N_25523,N_25997);
and U26218 (N_26218,N_25949,N_25711);
nand U26219 (N_26219,N_25679,N_25630);
nor U26220 (N_26220,N_25922,N_25881);
or U26221 (N_26221,N_25964,N_25967);
xor U26222 (N_26222,N_25882,N_25920);
or U26223 (N_26223,N_25762,N_25732);
nand U26224 (N_26224,N_25795,N_25709);
nor U26225 (N_26225,N_25750,N_25675);
nor U26226 (N_26226,N_25640,N_25841);
xor U26227 (N_26227,N_25654,N_25556);
and U26228 (N_26228,N_25912,N_25914);
nor U26229 (N_26229,N_25704,N_25933);
nor U26230 (N_26230,N_25907,N_25682);
xnor U26231 (N_26231,N_25831,N_25645);
nor U26232 (N_26232,N_25662,N_25811);
nand U26233 (N_26233,N_25741,N_25805);
and U26234 (N_26234,N_25756,N_25998);
nand U26235 (N_26235,N_25826,N_25717);
nand U26236 (N_26236,N_25567,N_25832);
and U26237 (N_26237,N_25845,N_25537);
and U26238 (N_26238,N_25521,N_25712);
nor U26239 (N_26239,N_25791,N_25601);
nor U26240 (N_26240,N_25588,N_25976);
and U26241 (N_26241,N_25844,N_25987);
nor U26242 (N_26242,N_25798,N_25883);
nor U26243 (N_26243,N_25962,N_25697);
xnor U26244 (N_26244,N_25721,N_25896);
nand U26245 (N_26245,N_25950,N_25846);
nand U26246 (N_26246,N_25958,N_25786);
xnor U26247 (N_26247,N_25858,N_25874);
nor U26248 (N_26248,N_25886,N_25701);
or U26249 (N_26249,N_25849,N_25801);
xor U26250 (N_26250,N_25767,N_25861);
and U26251 (N_26251,N_25770,N_25880);
nor U26252 (N_26252,N_25883,N_25619);
nor U26253 (N_26253,N_25991,N_25879);
or U26254 (N_26254,N_25649,N_25876);
nor U26255 (N_26255,N_25542,N_25626);
or U26256 (N_26256,N_25576,N_25581);
nor U26257 (N_26257,N_25953,N_25586);
xor U26258 (N_26258,N_25972,N_25584);
xnor U26259 (N_26259,N_25869,N_25888);
nand U26260 (N_26260,N_25568,N_25962);
or U26261 (N_26261,N_25801,N_25919);
and U26262 (N_26262,N_25618,N_25537);
xnor U26263 (N_26263,N_25747,N_25669);
and U26264 (N_26264,N_25631,N_25590);
nor U26265 (N_26265,N_25976,N_25711);
or U26266 (N_26266,N_25620,N_25992);
and U26267 (N_26267,N_25902,N_25625);
and U26268 (N_26268,N_25958,N_25963);
nor U26269 (N_26269,N_25918,N_25519);
xnor U26270 (N_26270,N_25983,N_25526);
and U26271 (N_26271,N_25505,N_25607);
nor U26272 (N_26272,N_25996,N_25580);
and U26273 (N_26273,N_25914,N_25670);
nor U26274 (N_26274,N_25968,N_25615);
or U26275 (N_26275,N_25890,N_25735);
and U26276 (N_26276,N_25838,N_25513);
or U26277 (N_26277,N_25506,N_25975);
nor U26278 (N_26278,N_25788,N_25767);
xnor U26279 (N_26279,N_25712,N_25564);
xor U26280 (N_26280,N_25771,N_25750);
or U26281 (N_26281,N_25570,N_25785);
nor U26282 (N_26282,N_25707,N_25758);
and U26283 (N_26283,N_25625,N_25761);
nand U26284 (N_26284,N_25812,N_25680);
nor U26285 (N_26285,N_25737,N_25800);
or U26286 (N_26286,N_25883,N_25926);
xor U26287 (N_26287,N_25977,N_25654);
nor U26288 (N_26288,N_25635,N_25653);
xor U26289 (N_26289,N_25576,N_25825);
xnor U26290 (N_26290,N_25948,N_25673);
xor U26291 (N_26291,N_25504,N_25898);
or U26292 (N_26292,N_25718,N_25644);
nor U26293 (N_26293,N_25574,N_25977);
xnor U26294 (N_26294,N_25822,N_25752);
nor U26295 (N_26295,N_25908,N_25594);
nand U26296 (N_26296,N_25553,N_25978);
and U26297 (N_26297,N_25636,N_25770);
nor U26298 (N_26298,N_25585,N_25776);
nand U26299 (N_26299,N_25998,N_25559);
or U26300 (N_26300,N_25740,N_25948);
and U26301 (N_26301,N_25694,N_25668);
nand U26302 (N_26302,N_25557,N_25523);
nand U26303 (N_26303,N_25753,N_25918);
and U26304 (N_26304,N_25568,N_25645);
or U26305 (N_26305,N_25890,N_25958);
or U26306 (N_26306,N_25578,N_25842);
or U26307 (N_26307,N_25883,N_25550);
nor U26308 (N_26308,N_25831,N_25784);
xnor U26309 (N_26309,N_25739,N_25685);
and U26310 (N_26310,N_25649,N_25554);
nor U26311 (N_26311,N_25607,N_25772);
or U26312 (N_26312,N_25933,N_25926);
or U26313 (N_26313,N_25526,N_25593);
and U26314 (N_26314,N_25529,N_25593);
and U26315 (N_26315,N_25880,N_25563);
nand U26316 (N_26316,N_25603,N_25834);
and U26317 (N_26317,N_25682,N_25630);
and U26318 (N_26318,N_25678,N_25939);
and U26319 (N_26319,N_25705,N_25894);
nor U26320 (N_26320,N_25954,N_25810);
and U26321 (N_26321,N_25796,N_25696);
and U26322 (N_26322,N_25630,N_25838);
nor U26323 (N_26323,N_25554,N_25910);
nand U26324 (N_26324,N_25665,N_25652);
xor U26325 (N_26325,N_25970,N_25675);
and U26326 (N_26326,N_25614,N_25521);
or U26327 (N_26327,N_25627,N_25572);
nor U26328 (N_26328,N_25741,N_25792);
nor U26329 (N_26329,N_25563,N_25695);
xnor U26330 (N_26330,N_25759,N_25643);
and U26331 (N_26331,N_25642,N_25756);
and U26332 (N_26332,N_25643,N_25723);
and U26333 (N_26333,N_25574,N_25952);
nor U26334 (N_26334,N_25724,N_25900);
nand U26335 (N_26335,N_25509,N_25639);
xnor U26336 (N_26336,N_25773,N_25831);
nor U26337 (N_26337,N_25751,N_25861);
and U26338 (N_26338,N_25855,N_25776);
or U26339 (N_26339,N_25759,N_25985);
nand U26340 (N_26340,N_25887,N_25643);
xor U26341 (N_26341,N_25775,N_25696);
nand U26342 (N_26342,N_25702,N_25908);
and U26343 (N_26343,N_25669,N_25529);
nand U26344 (N_26344,N_25555,N_25668);
xnor U26345 (N_26345,N_25503,N_25756);
and U26346 (N_26346,N_25607,N_25844);
nor U26347 (N_26347,N_25591,N_25662);
nand U26348 (N_26348,N_25859,N_25651);
nand U26349 (N_26349,N_25661,N_25637);
and U26350 (N_26350,N_25690,N_25755);
xnor U26351 (N_26351,N_25858,N_25656);
nor U26352 (N_26352,N_25918,N_25840);
xor U26353 (N_26353,N_25804,N_25960);
nand U26354 (N_26354,N_25658,N_25657);
or U26355 (N_26355,N_25954,N_25609);
nor U26356 (N_26356,N_25975,N_25970);
nor U26357 (N_26357,N_25622,N_25889);
or U26358 (N_26358,N_25603,N_25712);
nor U26359 (N_26359,N_25745,N_25982);
nand U26360 (N_26360,N_25894,N_25902);
nand U26361 (N_26361,N_25528,N_25786);
nand U26362 (N_26362,N_25636,N_25732);
xor U26363 (N_26363,N_25836,N_25899);
xnor U26364 (N_26364,N_25785,N_25814);
and U26365 (N_26365,N_25814,N_25523);
xor U26366 (N_26366,N_25890,N_25654);
and U26367 (N_26367,N_25673,N_25681);
nand U26368 (N_26368,N_25756,N_25910);
or U26369 (N_26369,N_25837,N_25812);
nand U26370 (N_26370,N_25963,N_25947);
nor U26371 (N_26371,N_25976,N_25962);
nor U26372 (N_26372,N_25924,N_25616);
nor U26373 (N_26373,N_25661,N_25561);
and U26374 (N_26374,N_25864,N_25836);
xnor U26375 (N_26375,N_25522,N_25638);
nand U26376 (N_26376,N_25509,N_25830);
and U26377 (N_26377,N_25576,N_25854);
nor U26378 (N_26378,N_25834,N_25898);
or U26379 (N_26379,N_25683,N_25554);
and U26380 (N_26380,N_25932,N_25954);
nand U26381 (N_26381,N_25591,N_25896);
nor U26382 (N_26382,N_25613,N_25798);
nor U26383 (N_26383,N_25729,N_25962);
and U26384 (N_26384,N_25943,N_25725);
or U26385 (N_26385,N_25750,N_25616);
or U26386 (N_26386,N_25558,N_25520);
nor U26387 (N_26387,N_25657,N_25704);
nand U26388 (N_26388,N_25918,N_25740);
and U26389 (N_26389,N_25936,N_25540);
xnor U26390 (N_26390,N_25905,N_25902);
nand U26391 (N_26391,N_25591,N_25836);
nor U26392 (N_26392,N_25906,N_25579);
and U26393 (N_26393,N_25652,N_25800);
nor U26394 (N_26394,N_25594,N_25632);
or U26395 (N_26395,N_25555,N_25939);
or U26396 (N_26396,N_25848,N_25764);
nor U26397 (N_26397,N_25768,N_25707);
nand U26398 (N_26398,N_25769,N_25910);
nand U26399 (N_26399,N_25631,N_25853);
xor U26400 (N_26400,N_25761,N_25718);
and U26401 (N_26401,N_25887,N_25796);
and U26402 (N_26402,N_25573,N_25801);
nand U26403 (N_26403,N_25552,N_25542);
xor U26404 (N_26404,N_25847,N_25728);
nand U26405 (N_26405,N_25654,N_25656);
nor U26406 (N_26406,N_25784,N_25853);
xor U26407 (N_26407,N_25685,N_25863);
and U26408 (N_26408,N_25874,N_25570);
xnor U26409 (N_26409,N_25531,N_25843);
nand U26410 (N_26410,N_25553,N_25982);
or U26411 (N_26411,N_25714,N_25734);
or U26412 (N_26412,N_25656,N_25969);
or U26413 (N_26413,N_25527,N_25669);
nand U26414 (N_26414,N_25902,N_25788);
xnor U26415 (N_26415,N_25514,N_25953);
nor U26416 (N_26416,N_25769,N_25578);
nor U26417 (N_26417,N_25559,N_25616);
xor U26418 (N_26418,N_25822,N_25958);
and U26419 (N_26419,N_25984,N_25674);
nor U26420 (N_26420,N_25912,N_25739);
and U26421 (N_26421,N_25849,N_25697);
or U26422 (N_26422,N_25905,N_25762);
nor U26423 (N_26423,N_25693,N_25658);
or U26424 (N_26424,N_25928,N_25917);
nor U26425 (N_26425,N_25802,N_25781);
and U26426 (N_26426,N_25893,N_25968);
nor U26427 (N_26427,N_25584,N_25918);
and U26428 (N_26428,N_25504,N_25532);
nand U26429 (N_26429,N_25570,N_25607);
xor U26430 (N_26430,N_25987,N_25528);
nor U26431 (N_26431,N_25544,N_25532);
and U26432 (N_26432,N_25614,N_25621);
xnor U26433 (N_26433,N_25835,N_25883);
nand U26434 (N_26434,N_25754,N_25526);
and U26435 (N_26435,N_25818,N_25802);
and U26436 (N_26436,N_25904,N_25502);
and U26437 (N_26437,N_25568,N_25658);
nand U26438 (N_26438,N_25945,N_25758);
nand U26439 (N_26439,N_25629,N_25557);
or U26440 (N_26440,N_25810,N_25621);
xor U26441 (N_26441,N_25906,N_25742);
or U26442 (N_26442,N_25743,N_25900);
nand U26443 (N_26443,N_25859,N_25714);
nor U26444 (N_26444,N_25883,N_25755);
or U26445 (N_26445,N_25538,N_25643);
nand U26446 (N_26446,N_25954,N_25802);
nand U26447 (N_26447,N_25742,N_25590);
and U26448 (N_26448,N_25787,N_25559);
or U26449 (N_26449,N_25543,N_25745);
xnor U26450 (N_26450,N_25837,N_25965);
nor U26451 (N_26451,N_25861,N_25870);
xnor U26452 (N_26452,N_25778,N_25550);
nor U26453 (N_26453,N_25677,N_25509);
nand U26454 (N_26454,N_25991,N_25677);
or U26455 (N_26455,N_25861,N_25931);
nand U26456 (N_26456,N_25674,N_25572);
nor U26457 (N_26457,N_25803,N_25908);
nor U26458 (N_26458,N_25506,N_25567);
nand U26459 (N_26459,N_25781,N_25983);
and U26460 (N_26460,N_25839,N_25805);
and U26461 (N_26461,N_25878,N_25514);
nand U26462 (N_26462,N_25524,N_25537);
or U26463 (N_26463,N_25874,N_25992);
nand U26464 (N_26464,N_25558,N_25762);
nand U26465 (N_26465,N_25967,N_25965);
xor U26466 (N_26466,N_25853,N_25587);
nand U26467 (N_26467,N_25616,N_25696);
nand U26468 (N_26468,N_25861,N_25691);
nor U26469 (N_26469,N_25636,N_25544);
or U26470 (N_26470,N_25651,N_25952);
or U26471 (N_26471,N_25629,N_25762);
nor U26472 (N_26472,N_25924,N_25653);
and U26473 (N_26473,N_25984,N_25786);
nor U26474 (N_26474,N_25906,N_25985);
and U26475 (N_26475,N_25641,N_25816);
xnor U26476 (N_26476,N_25522,N_25956);
nor U26477 (N_26477,N_25531,N_25967);
or U26478 (N_26478,N_25924,N_25948);
xor U26479 (N_26479,N_25899,N_25873);
or U26480 (N_26480,N_25517,N_25746);
nor U26481 (N_26481,N_25502,N_25741);
nor U26482 (N_26482,N_25800,N_25858);
and U26483 (N_26483,N_25976,N_25801);
nor U26484 (N_26484,N_25709,N_25802);
or U26485 (N_26485,N_25677,N_25553);
nand U26486 (N_26486,N_25864,N_25947);
and U26487 (N_26487,N_25991,N_25558);
nor U26488 (N_26488,N_25842,N_25530);
nor U26489 (N_26489,N_25577,N_25912);
nand U26490 (N_26490,N_25816,N_25914);
xnor U26491 (N_26491,N_25749,N_25732);
nand U26492 (N_26492,N_25690,N_25724);
and U26493 (N_26493,N_25560,N_25690);
nand U26494 (N_26494,N_25532,N_25864);
nand U26495 (N_26495,N_25994,N_25891);
nand U26496 (N_26496,N_25928,N_25950);
nor U26497 (N_26497,N_25812,N_25661);
or U26498 (N_26498,N_25511,N_25976);
or U26499 (N_26499,N_25950,N_25595);
and U26500 (N_26500,N_26471,N_26324);
nor U26501 (N_26501,N_26146,N_26087);
xor U26502 (N_26502,N_26103,N_26349);
and U26503 (N_26503,N_26305,N_26325);
nand U26504 (N_26504,N_26088,N_26100);
and U26505 (N_26505,N_26013,N_26322);
nand U26506 (N_26506,N_26312,N_26356);
nor U26507 (N_26507,N_26173,N_26237);
or U26508 (N_26508,N_26451,N_26002);
xnor U26509 (N_26509,N_26338,N_26093);
nor U26510 (N_26510,N_26086,N_26423);
xnor U26511 (N_26511,N_26004,N_26449);
nor U26512 (N_26512,N_26080,N_26355);
xor U26513 (N_26513,N_26094,N_26211);
xor U26514 (N_26514,N_26328,N_26192);
and U26515 (N_26515,N_26224,N_26274);
nor U26516 (N_26516,N_26134,N_26031);
nor U26517 (N_26517,N_26076,N_26268);
and U26518 (N_26518,N_26141,N_26046);
nand U26519 (N_26519,N_26118,N_26409);
and U26520 (N_26520,N_26036,N_26179);
and U26521 (N_26521,N_26114,N_26170);
xor U26522 (N_26522,N_26015,N_26207);
and U26523 (N_26523,N_26360,N_26233);
nor U26524 (N_26524,N_26099,N_26083);
and U26525 (N_26525,N_26318,N_26313);
nand U26526 (N_26526,N_26033,N_26180);
or U26527 (N_26527,N_26441,N_26149);
nand U26528 (N_26528,N_26491,N_26011);
or U26529 (N_26529,N_26055,N_26417);
and U26530 (N_26530,N_26035,N_26085);
or U26531 (N_26531,N_26369,N_26054);
nor U26532 (N_26532,N_26473,N_26479);
nor U26533 (N_26533,N_26460,N_26320);
and U26534 (N_26534,N_26095,N_26019);
or U26535 (N_26535,N_26182,N_26056);
nor U26536 (N_26536,N_26257,N_26465);
and U26537 (N_26537,N_26499,N_26112);
xnor U26538 (N_26538,N_26484,N_26452);
nor U26539 (N_26539,N_26345,N_26472);
nand U26540 (N_26540,N_26153,N_26288);
nor U26541 (N_26541,N_26271,N_26436);
nor U26542 (N_26542,N_26474,N_26202);
and U26543 (N_26543,N_26132,N_26186);
nand U26544 (N_26544,N_26163,N_26295);
or U26545 (N_26545,N_26275,N_26077);
nand U26546 (N_26546,N_26158,N_26034);
xnor U26547 (N_26547,N_26453,N_26497);
and U26548 (N_26548,N_26361,N_26287);
and U26549 (N_26549,N_26063,N_26315);
or U26550 (N_26550,N_26045,N_26062);
nor U26551 (N_26551,N_26074,N_26205);
and U26552 (N_26552,N_26379,N_26363);
nand U26553 (N_26553,N_26350,N_26286);
and U26554 (N_26554,N_26343,N_26210);
or U26555 (N_26555,N_26248,N_26492);
nor U26556 (N_26556,N_26483,N_26160);
or U26557 (N_26557,N_26388,N_26424);
and U26558 (N_26558,N_26282,N_26265);
nor U26559 (N_26559,N_26053,N_26162);
or U26560 (N_26560,N_26391,N_26220);
xor U26561 (N_26561,N_26309,N_26323);
nand U26562 (N_26562,N_26110,N_26001);
xor U26563 (N_26563,N_26425,N_26346);
or U26564 (N_26564,N_26098,N_26404);
nand U26565 (N_26565,N_26384,N_26301);
nor U26566 (N_26566,N_26129,N_26392);
nand U26567 (N_26567,N_26333,N_26281);
xor U26568 (N_26568,N_26276,N_26334);
and U26569 (N_26569,N_26406,N_26157);
xor U26570 (N_26570,N_26487,N_26000);
nor U26571 (N_26571,N_26169,N_26232);
or U26572 (N_26572,N_26168,N_26340);
nand U26573 (N_26573,N_26241,N_26475);
nand U26574 (N_26574,N_26066,N_26413);
or U26575 (N_26575,N_26300,N_26222);
xor U26576 (N_26576,N_26040,N_26032);
and U26577 (N_26577,N_26403,N_26249);
or U26578 (N_26578,N_26029,N_26234);
nor U26579 (N_26579,N_26373,N_26092);
nor U26580 (N_26580,N_26358,N_26496);
nor U26581 (N_26581,N_26044,N_26398);
and U26582 (N_26582,N_26331,N_26187);
nand U26583 (N_26583,N_26057,N_26304);
nand U26584 (N_26584,N_26172,N_26293);
nor U26585 (N_26585,N_26476,N_26364);
nand U26586 (N_26586,N_26468,N_26126);
xnor U26587 (N_26587,N_26432,N_26143);
nand U26588 (N_26588,N_26302,N_26067);
or U26589 (N_26589,N_26006,N_26127);
nor U26590 (N_26590,N_26329,N_26140);
or U26591 (N_26591,N_26101,N_26121);
or U26592 (N_26592,N_26003,N_26117);
nor U26593 (N_26593,N_26039,N_26022);
nand U26594 (N_26594,N_26156,N_26297);
and U26595 (N_26595,N_26089,N_26050);
nor U26596 (N_26596,N_26016,N_26250);
or U26597 (N_26597,N_26108,N_26240);
or U26598 (N_26598,N_26014,N_26367);
nor U26599 (N_26599,N_26113,N_26348);
xnor U26600 (N_26600,N_26339,N_26267);
or U26601 (N_26601,N_26310,N_26467);
and U26602 (N_26602,N_26221,N_26058);
nor U26603 (N_26603,N_26494,N_26381);
and U26604 (N_26604,N_26125,N_26133);
and U26605 (N_26605,N_26079,N_26081);
or U26606 (N_26606,N_26437,N_26458);
xnor U26607 (N_26607,N_26266,N_26090);
xor U26608 (N_26608,N_26445,N_26420);
nand U26609 (N_26609,N_26256,N_26226);
or U26610 (N_26610,N_26122,N_26138);
nor U26611 (N_26611,N_26236,N_26185);
and U26612 (N_26612,N_26383,N_26049);
or U26613 (N_26613,N_26390,N_26136);
or U26614 (N_26614,N_26463,N_26213);
xor U26615 (N_26615,N_26455,N_26230);
xnor U26616 (N_26616,N_26128,N_26204);
or U26617 (N_26617,N_26037,N_26135);
or U26618 (N_26618,N_26190,N_26247);
and U26619 (N_26619,N_26264,N_26308);
and U26620 (N_26620,N_26374,N_26262);
xor U26621 (N_26621,N_26464,N_26047);
or U26622 (N_26622,N_26400,N_26238);
nand U26623 (N_26623,N_26109,N_26191);
nand U26624 (N_26624,N_26407,N_26311);
nand U26625 (N_26625,N_26025,N_26270);
xnor U26626 (N_26626,N_26326,N_26450);
xnor U26627 (N_26627,N_26498,N_26064);
xor U26628 (N_26628,N_26184,N_26052);
and U26629 (N_26629,N_26106,N_26393);
nor U26630 (N_26630,N_26380,N_26427);
xnor U26631 (N_26631,N_26068,N_26072);
nand U26632 (N_26632,N_26462,N_26371);
xnor U26633 (N_26633,N_26151,N_26231);
or U26634 (N_26634,N_26102,N_26154);
xor U26635 (N_26635,N_26228,N_26477);
or U26636 (N_26636,N_26028,N_26199);
nand U26637 (N_26637,N_26330,N_26335);
nor U26638 (N_26638,N_26411,N_26147);
or U26639 (N_26639,N_26137,N_26486);
and U26640 (N_26640,N_26005,N_26303);
nor U26641 (N_26641,N_26319,N_26148);
or U26642 (N_26642,N_26219,N_26254);
nor U26643 (N_26643,N_26481,N_26489);
nand U26644 (N_26644,N_26194,N_26107);
or U26645 (N_26645,N_26278,N_26306);
nand U26646 (N_26646,N_26347,N_26239);
xnor U26647 (N_26647,N_26131,N_26024);
or U26648 (N_26648,N_26203,N_26353);
nand U26649 (N_26649,N_26327,N_26084);
and U26650 (N_26650,N_26375,N_26030);
or U26651 (N_26651,N_26442,N_26457);
nand U26652 (N_26652,N_26272,N_26292);
or U26653 (N_26653,N_26317,N_26405);
and U26654 (N_26654,N_26217,N_26454);
and U26655 (N_26655,N_26111,N_26116);
or U26656 (N_26656,N_26421,N_26161);
nor U26657 (N_26657,N_26439,N_26480);
nand U26658 (N_26658,N_26433,N_26201);
and U26659 (N_26659,N_26352,N_26428);
and U26660 (N_26660,N_26419,N_26259);
nand U26661 (N_26661,N_26060,N_26438);
xor U26662 (N_26662,N_26104,N_26115);
and U26663 (N_26663,N_26321,N_26008);
xor U26664 (N_26664,N_26478,N_26142);
nor U26665 (N_26665,N_26208,N_26470);
nor U26666 (N_26666,N_26119,N_26279);
xor U26667 (N_26667,N_26183,N_26255);
xor U26668 (N_26668,N_26395,N_26431);
xor U26669 (N_26669,N_26298,N_26469);
or U26670 (N_26670,N_26252,N_26216);
and U26671 (N_26671,N_26263,N_26408);
xor U26672 (N_26672,N_26482,N_26144);
nor U26673 (N_26673,N_26166,N_26150);
xnor U26674 (N_26674,N_26177,N_26145);
or U26675 (N_26675,N_26399,N_26466);
nand U26676 (N_26676,N_26073,N_26176);
nor U26677 (N_26677,N_26485,N_26294);
and U26678 (N_26678,N_26246,N_26260);
xnor U26679 (N_26679,N_26316,N_26357);
nor U26680 (N_26680,N_26065,N_26459);
or U26681 (N_26681,N_26043,N_26443);
xor U26682 (N_26682,N_26426,N_26382);
and U26683 (N_26683,N_26130,N_26307);
or U26684 (N_26684,N_26193,N_26446);
nand U26685 (N_26685,N_26139,N_26299);
or U26686 (N_26686,N_26447,N_26314);
xnor U26687 (N_26687,N_26189,N_26209);
xnor U26688 (N_26688,N_26261,N_26415);
or U26689 (N_26689,N_26402,N_26337);
nor U26690 (N_26690,N_26026,N_26258);
nand U26691 (N_26691,N_26244,N_26370);
nor U26692 (N_26692,N_26051,N_26386);
or U26693 (N_26693,N_26289,N_26164);
nor U26694 (N_26694,N_26215,N_26283);
and U26695 (N_26695,N_26225,N_26071);
nor U26696 (N_26696,N_26023,N_26490);
xor U26697 (N_26697,N_26253,N_26198);
or U26698 (N_26698,N_26243,N_26048);
or U26699 (N_26699,N_26200,N_26075);
nand U26700 (N_26700,N_26242,N_26082);
and U26701 (N_26701,N_26269,N_26351);
or U26702 (N_26702,N_26376,N_26285);
nand U26703 (N_26703,N_26175,N_26165);
nand U26704 (N_26704,N_26378,N_26096);
nor U26705 (N_26705,N_26010,N_26017);
nand U26706 (N_26706,N_26007,N_26493);
nand U26707 (N_26707,N_26429,N_26078);
or U26708 (N_26708,N_26488,N_26397);
and U26709 (N_26709,N_26124,N_26332);
nand U26710 (N_26710,N_26277,N_26434);
and U26711 (N_26711,N_26159,N_26495);
nor U26712 (N_26712,N_26188,N_26394);
or U26713 (N_26713,N_26422,N_26195);
or U26714 (N_26714,N_26354,N_26389);
and U26715 (N_26715,N_26021,N_26273);
nor U26716 (N_26716,N_26359,N_26181);
nor U26717 (N_26717,N_26385,N_26448);
and U26718 (N_26718,N_26218,N_26227);
or U26719 (N_26719,N_26214,N_26120);
xnor U26720 (N_26720,N_26396,N_26097);
or U26721 (N_26721,N_26196,N_26461);
or U26722 (N_26722,N_26059,N_26362);
nand U26723 (N_26723,N_26291,N_26366);
xnor U26724 (N_26724,N_26235,N_26020);
and U26725 (N_26725,N_26018,N_26412);
nor U26726 (N_26726,N_26387,N_26401);
xnor U26727 (N_26727,N_26229,N_26456);
nand U26728 (N_26728,N_26368,N_26410);
and U26729 (N_26729,N_26280,N_26105);
xnor U26730 (N_26730,N_26070,N_26344);
xor U26731 (N_26731,N_26290,N_26212);
and U26732 (N_26732,N_26206,N_26365);
xnor U26733 (N_26733,N_26223,N_26038);
or U26734 (N_26734,N_26167,N_26414);
nand U26735 (N_26735,N_26444,N_26152);
and U26736 (N_26736,N_26296,N_26178);
xor U26737 (N_26737,N_26416,N_26012);
nor U26738 (N_26738,N_26174,N_26430);
nor U26739 (N_26739,N_26061,N_26123);
nand U26740 (N_26740,N_26435,N_26155);
nand U26741 (N_26741,N_26027,N_26440);
or U26742 (N_26742,N_26009,N_26336);
or U26743 (N_26743,N_26171,N_26284);
and U26744 (N_26744,N_26418,N_26245);
nor U26745 (N_26745,N_26069,N_26342);
nor U26746 (N_26746,N_26251,N_26341);
nor U26747 (N_26747,N_26377,N_26042);
nor U26748 (N_26748,N_26091,N_26041);
nor U26749 (N_26749,N_26197,N_26372);
or U26750 (N_26750,N_26187,N_26372);
nand U26751 (N_26751,N_26067,N_26023);
nor U26752 (N_26752,N_26490,N_26487);
or U26753 (N_26753,N_26340,N_26379);
nand U26754 (N_26754,N_26433,N_26093);
or U26755 (N_26755,N_26498,N_26180);
or U26756 (N_26756,N_26052,N_26497);
or U26757 (N_26757,N_26411,N_26445);
xnor U26758 (N_26758,N_26110,N_26469);
xnor U26759 (N_26759,N_26145,N_26162);
or U26760 (N_26760,N_26425,N_26212);
xor U26761 (N_26761,N_26011,N_26303);
nor U26762 (N_26762,N_26401,N_26294);
nand U26763 (N_26763,N_26080,N_26251);
xnor U26764 (N_26764,N_26348,N_26442);
and U26765 (N_26765,N_26483,N_26046);
nor U26766 (N_26766,N_26219,N_26470);
and U26767 (N_26767,N_26359,N_26230);
or U26768 (N_26768,N_26132,N_26283);
xor U26769 (N_26769,N_26131,N_26296);
nor U26770 (N_26770,N_26021,N_26033);
nor U26771 (N_26771,N_26139,N_26145);
nor U26772 (N_26772,N_26454,N_26404);
nand U26773 (N_26773,N_26443,N_26029);
nand U26774 (N_26774,N_26272,N_26082);
and U26775 (N_26775,N_26270,N_26039);
and U26776 (N_26776,N_26191,N_26111);
xnor U26777 (N_26777,N_26099,N_26329);
nor U26778 (N_26778,N_26356,N_26372);
and U26779 (N_26779,N_26032,N_26397);
and U26780 (N_26780,N_26311,N_26184);
and U26781 (N_26781,N_26032,N_26114);
nand U26782 (N_26782,N_26064,N_26041);
xor U26783 (N_26783,N_26109,N_26265);
xnor U26784 (N_26784,N_26276,N_26467);
nand U26785 (N_26785,N_26097,N_26484);
and U26786 (N_26786,N_26195,N_26304);
nor U26787 (N_26787,N_26364,N_26191);
nor U26788 (N_26788,N_26468,N_26235);
and U26789 (N_26789,N_26178,N_26394);
nor U26790 (N_26790,N_26343,N_26143);
nand U26791 (N_26791,N_26012,N_26082);
nor U26792 (N_26792,N_26230,N_26224);
xnor U26793 (N_26793,N_26082,N_26071);
nand U26794 (N_26794,N_26444,N_26390);
nor U26795 (N_26795,N_26440,N_26290);
nor U26796 (N_26796,N_26006,N_26008);
nor U26797 (N_26797,N_26280,N_26003);
and U26798 (N_26798,N_26144,N_26463);
nand U26799 (N_26799,N_26077,N_26215);
nor U26800 (N_26800,N_26246,N_26393);
nand U26801 (N_26801,N_26308,N_26200);
or U26802 (N_26802,N_26092,N_26386);
nand U26803 (N_26803,N_26264,N_26407);
nand U26804 (N_26804,N_26289,N_26442);
nor U26805 (N_26805,N_26259,N_26196);
xnor U26806 (N_26806,N_26369,N_26235);
xor U26807 (N_26807,N_26268,N_26335);
or U26808 (N_26808,N_26055,N_26445);
and U26809 (N_26809,N_26323,N_26332);
nand U26810 (N_26810,N_26392,N_26260);
nor U26811 (N_26811,N_26487,N_26126);
and U26812 (N_26812,N_26221,N_26333);
nor U26813 (N_26813,N_26436,N_26321);
nor U26814 (N_26814,N_26056,N_26012);
or U26815 (N_26815,N_26071,N_26205);
xnor U26816 (N_26816,N_26463,N_26299);
and U26817 (N_26817,N_26206,N_26307);
or U26818 (N_26818,N_26327,N_26063);
nand U26819 (N_26819,N_26418,N_26469);
nand U26820 (N_26820,N_26193,N_26040);
nor U26821 (N_26821,N_26452,N_26373);
nor U26822 (N_26822,N_26150,N_26066);
nor U26823 (N_26823,N_26495,N_26204);
and U26824 (N_26824,N_26346,N_26208);
xor U26825 (N_26825,N_26060,N_26328);
xnor U26826 (N_26826,N_26103,N_26476);
xnor U26827 (N_26827,N_26345,N_26425);
nand U26828 (N_26828,N_26481,N_26127);
or U26829 (N_26829,N_26072,N_26199);
nor U26830 (N_26830,N_26154,N_26031);
nor U26831 (N_26831,N_26146,N_26232);
nand U26832 (N_26832,N_26069,N_26213);
nor U26833 (N_26833,N_26422,N_26173);
and U26834 (N_26834,N_26379,N_26487);
nand U26835 (N_26835,N_26468,N_26041);
or U26836 (N_26836,N_26414,N_26381);
nor U26837 (N_26837,N_26252,N_26255);
xnor U26838 (N_26838,N_26191,N_26384);
or U26839 (N_26839,N_26416,N_26017);
nand U26840 (N_26840,N_26321,N_26275);
xnor U26841 (N_26841,N_26294,N_26453);
nand U26842 (N_26842,N_26057,N_26064);
nor U26843 (N_26843,N_26462,N_26408);
nor U26844 (N_26844,N_26095,N_26147);
xnor U26845 (N_26845,N_26309,N_26003);
or U26846 (N_26846,N_26370,N_26303);
xnor U26847 (N_26847,N_26218,N_26044);
nand U26848 (N_26848,N_26017,N_26067);
nand U26849 (N_26849,N_26154,N_26244);
xnor U26850 (N_26850,N_26348,N_26301);
xnor U26851 (N_26851,N_26370,N_26327);
nand U26852 (N_26852,N_26423,N_26283);
or U26853 (N_26853,N_26011,N_26172);
or U26854 (N_26854,N_26086,N_26081);
nand U26855 (N_26855,N_26131,N_26462);
nor U26856 (N_26856,N_26274,N_26356);
nor U26857 (N_26857,N_26279,N_26068);
or U26858 (N_26858,N_26234,N_26360);
nor U26859 (N_26859,N_26463,N_26402);
nor U26860 (N_26860,N_26332,N_26139);
nand U26861 (N_26861,N_26115,N_26259);
xor U26862 (N_26862,N_26076,N_26277);
nand U26863 (N_26863,N_26096,N_26270);
or U26864 (N_26864,N_26352,N_26366);
nand U26865 (N_26865,N_26024,N_26389);
and U26866 (N_26866,N_26055,N_26312);
nor U26867 (N_26867,N_26452,N_26210);
xor U26868 (N_26868,N_26443,N_26136);
or U26869 (N_26869,N_26194,N_26345);
or U26870 (N_26870,N_26125,N_26365);
nand U26871 (N_26871,N_26089,N_26196);
and U26872 (N_26872,N_26012,N_26038);
nand U26873 (N_26873,N_26154,N_26239);
nor U26874 (N_26874,N_26293,N_26379);
or U26875 (N_26875,N_26271,N_26326);
or U26876 (N_26876,N_26348,N_26330);
and U26877 (N_26877,N_26063,N_26403);
and U26878 (N_26878,N_26272,N_26187);
xor U26879 (N_26879,N_26024,N_26393);
nor U26880 (N_26880,N_26075,N_26210);
xor U26881 (N_26881,N_26056,N_26215);
and U26882 (N_26882,N_26057,N_26373);
or U26883 (N_26883,N_26216,N_26022);
and U26884 (N_26884,N_26089,N_26139);
xor U26885 (N_26885,N_26206,N_26288);
nand U26886 (N_26886,N_26202,N_26328);
xor U26887 (N_26887,N_26240,N_26216);
xnor U26888 (N_26888,N_26343,N_26268);
nor U26889 (N_26889,N_26063,N_26310);
and U26890 (N_26890,N_26496,N_26033);
nor U26891 (N_26891,N_26429,N_26453);
nor U26892 (N_26892,N_26434,N_26423);
xor U26893 (N_26893,N_26201,N_26265);
nand U26894 (N_26894,N_26088,N_26404);
or U26895 (N_26895,N_26098,N_26106);
nor U26896 (N_26896,N_26098,N_26030);
xnor U26897 (N_26897,N_26424,N_26224);
nor U26898 (N_26898,N_26450,N_26350);
or U26899 (N_26899,N_26384,N_26151);
and U26900 (N_26900,N_26199,N_26494);
or U26901 (N_26901,N_26445,N_26240);
xnor U26902 (N_26902,N_26062,N_26230);
xnor U26903 (N_26903,N_26400,N_26367);
nand U26904 (N_26904,N_26005,N_26410);
or U26905 (N_26905,N_26120,N_26468);
nor U26906 (N_26906,N_26164,N_26378);
nand U26907 (N_26907,N_26307,N_26170);
and U26908 (N_26908,N_26230,N_26231);
nor U26909 (N_26909,N_26365,N_26065);
and U26910 (N_26910,N_26496,N_26469);
nand U26911 (N_26911,N_26155,N_26139);
xnor U26912 (N_26912,N_26401,N_26149);
and U26913 (N_26913,N_26462,N_26091);
nand U26914 (N_26914,N_26251,N_26336);
or U26915 (N_26915,N_26307,N_26123);
xnor U26916 (N_26916,N_26342,N_26437);
or U26917 (N_26917,N_26059,N_26251);
xor U26918 (N_26918,N_26310,N_26129);
and U26919 (N_26919,N_26159,N_26034);
or U26920 (N_26920,N_26172,N_26179);
nand U26921 (N_26921,N_26294,N_26227);
and U26922 (N_26922,N_26143,N_26315);
xor U26923 (N_26923,N_26106,N_26207);
nor U26924 (N_26924,N_26170,N_26149);
xnor U26925 (N_26925,N_26262,N_26438);
or U26926 (N_26926,N_26384,N_26017);
nor U26927 (N_26927,N_26318,N_26152);
or U26928 (N_26928,N_26093,N_26350);
xor U26929 (N_26929,N_26337,N_26249);
xnor U26930 (N_26930,N_26113,N_26080);
or U26931 (N_26931,N_26121,N_26037);
nand U26932 (N_26932,N_26231,N_26250);
nand U26933 (N_26933,N_26004,N_26472);
xor U26934 (N_26934,N_26454,N_26102);
or U26935 (N_26935,N_26022,N_26296);
nor U26936 (N_26936,N_26391,N_26444);
nor U26937 (N_26937,N_26364,N_26468);
xor U26938 (N_26938,N_26368,N_26219);
xnor U26939 (N_26939,N_26490,N_26070);
or U26940 (N_26940,N_26162,N_26407);
xnor U26941 (N_26941,N_26003,N_26001);
xnor U26942 (N_26942,N_26318,N_26033);
or U26943 (N_26943,N_26128,N_26284);
or U26944 (N_26944,N_26205,N_26364);
xor U26945 (N_26945,N_26172,N_26311);
or U26946 (N_26946,N_26418,N_26307);
and U26947 (N_26947,N_26311,N_26265);
xnor U26948 (N_26948,N_26125,N_26359);
nor U26949 (N_26949,N_26298,N_26369);
or U26950 (N_26950,N_26429,N_26242);
or U26951 (N_26951,N_26389,N_26431);
nor U26952 (N_26952,N_26107,N_26080);
or U26953 (N_26953,N_26207,N_26496);
and U26954 (N_26954,N_26401,N_26250);
and U26955 (N_26955,N_26293,N_26070);
and U26956 (N_26956,N_26093,N_26158);
and U26957 (N_26957,N_26311,N_26180);
xnor U26958 (N_26958,N_26432,N_26191);
nor U26959 (N_26959,N_26053,N_26201);
and U26960 (N_26960,N_26293,N_26303);
nor U26961 (N_26961,N_26259,N_26334);
nand U26962 (N_26962,N_26328,N_26013);
or U26963 (N_26963,N_26222,N_26029);
nor U26964 (N_26964,N_26441,N_26117);
nand U26965 (N_26965,N_26289,N_26084);
and U26966 (N_26966,N_26363,N_26025);
nand U26967 (N_26967,N_26435,N_26490);
and U26968 (N_26968,N_26103,N_26145);
nand U26969 (N_26969,N_26460,N_26424);
nand U26970 (N_26970,N_26084,N_26423);
or U26971 (N_26971,N_26221,N_26279);
and U26972 (N_26972,N_26240,N_26185);
xnor U26973 (N_26973,N_26296,N_26340);
or U26974 (N_26974,N_26001,N_26307);
nand U26975 (N_26975,N_26319,N_26472);
and U26976 (N_26976,N_26220,N_26138);
nand U26977 (N_26977,N_26006,N_26272);
nor U26978 (N_26978,N_26436,N_26470);
and U26979 (N_26979,N_26277,N_26219);
xor U26980 (N_26980,N_26193,N_26205);
and U26981 (N_26981,N_26036,N_26318);
or U26982 (N_26982,N_26262,N_26345);
xor U26983 (N_26983,N_26362,N_26237);
nor U26984 (N_26984,N_26346,N_26344);
or U26985 (N_26985,N_26216,N_26373);
nand U26986 (N_26986,N_26123,N_26012);
nand U26987 (N_26987,N_26321,N_26317);
nand U26988 (N_26988,N_26272,N_26308);
xnor U26989 (N_26989,N_26127,N_26490);
xor U26990 (N_26990,N_26217,N_26372);
nand U26991 (N_26991,N_26185,N_26198);
xnor U26992 (N_26992,N_26174,N_26403);
xor U26993 (N_26993,N_26020,N_26439);
nand U26994 (N_26994,N_26204,N_26355);
or U26995 (N_26995,N_26316,N_26135);
and U26996 (N_26996,N_26331,N_26285);
nand U26997 (N_26997,N_26032,N_26369);
nor U26998 (N_26998,N_26105,N_26468);
and U26999 (N_26999,N_26207,N_26369);
nor U27000 (N_27000,N_26848,N_26658);
nand U27001 (N_27001,N_26645,N_26800);
nand U27002 (N_27002,N_26503,N_26761);
or U27003 (N_27003,N_26775,N_26846);
and U27004 (N_27004,N_26587,N_26615);
xnor U27005 (N_27005,N_26888,N_26746);
and U27006 (N_27006,N_26737,N_26769);
nand U27007 (N_27007,N_26627,N_26900);
xnor U27008 (N_27008,N_26940,N_26817);
nor U27009 (N_27009,N_26763,N_26949);
nor U27010 (N_27010,N_26506,N_26918);
xnor U27011 (N_27011,N_26558,N_26859);
nor U27012 (N_27012,N_26885,N_26708);
nor U27013 (N_27013,N_26982,N_26955);
and U27014 (N_27014,N_26588,N_26738);
nand U27015 (N_27015,N_26633,N_26921);
xor U27016 (N_27016,N_26785,N_26944);
nand U27017 (N_27017,N_26592,N_26546);
nand U27018 (N_27018,N_26953,N_26826);
and U27019 (N_27019,N_26618,N_26750);
or U27020 (N_27020,N_26860,N_26976);
and U27021 (N_27021,N_26518,N_26676);
or U27022 (N_27022,N_26724,N_26901);
nand U27023 (N_27023,N_26603,N_26666);
nand U27024 (N_27024,N_26688,N_26547);
xnor U27025 (N_27025,N_26881,N_26648);
nand U27026 (N_27026,N_26698,N_26774);
nor U27027 (N_27027,N_26864,N_26757);
nand U27028 (N_27028,N_26744,N_26910);
and U27029 (N_27029,N_26788,N_26849);
nand U27030 (N_27030,N_26613,N_26543);
or U27031 (N_27031,N_26793,N_26649);
nand U27032 (N_27032,N_26689,N_26960);
or U27033 (N_27033,N_26534,N_26784);
or U27034 (N_27034,N_26959,N_26541);
and U27035 (N_27035,N_26987,N_26681);
or U27036 (N_27036,N_26725,N_26782);
nor U27037 (N_27037,N_26745,N_26805);
nor U27038 (N_27038,N_26553,N_26651);
or U27039 (N_27039,N_26971,N_26523);
xnor U27040 (N_27040,N_26994,N_26566);
nand U27041 (N_27041,N_26624,N_26515);
nand U27042 (N_27042,N_26605,N_26767);
xor U27043 (N_27043,N_26673,N_26762);
nor U27044 (N_27044,N_26884,N_26749);
or U27045 (N_27045,N_26617,N_26836);
and U27046 (N_27046,N_26781,N_26526);
or U27047 (N_27047,N_26520,N_26913);
nor U27048 (N_27048,N_26926,N_26650);
xnor U27049 (N_27049,N_26716,N_26586);
nand U27050 (N_27050,N_26896,N_26943);
nor U27051 (N_27051,N_26683,N_26659);
nand U27052 (N_27052,N_26766,N_26593);
nor U27053 (N_27053,N_26642,N_26908);
nand U27054 (N_27054,N_26614,N_26606);
or U27055 (N_27055,N_26760,N_26705);
nand U27056 (N_27056,N_26721,N_26616);
nand U27057 (N_27057,N_26679,N_26641);
nor U27058 (N_27058,N_26646,N_26776);
nand U27059 (N_27059,N_26741,N_26902);
nor U27060 (N_27060,N_26999,N_26570);
xnor U27061 (N_27061,N_26956,N_26667);
nand U27062 (N_27062,N_26561,N_26858);
nor U27063 (N_27063,N_26704,N_26925);
nand U27064 (N_27064,N_26713,N_26535);
xnor U27065 (N_27065,N_26540,N_26796);
or U27066 (N_27066,N_26829,N_26664);
nor U27067 (N_27067,N_26780,N_26807);
nand U27068 (N_27068,N_26564,N_26604);
and U27069 (N_27069,N_26810,N_26983);
nor U27070 (N_27070,N_26854,N_26549);
or U27071 (N_27071,N_26717,N_26815);
xnor U27072 (N_27072,N_26873,N_26772);
or U27073 (N_27073,N_26692,N_26516);
xor U27074 (N_27074,N_26719,N_26919);
and U27075 (N_27075,N_26878,N_26813);
and U27076 (N_27076,N_26928,N_26690);
nand U27077 (N_27077,N_26590,N_26920);
xnor U27078 (N_27078,N_26947,N_26609);
and U27079 (N_27079,N_26801,N_26711);
xnor U27080 (N_27080,N_26795,N_26970);
and U27081 (N_27081,N_26509,N_26968);
nand U27082 (N_27082,N_26922,N_26589);
xnor U27083 (N_27083,N_26519,N_26841);
xnor U27084 (N_27084,N_26967,N_26798);
nor U27085 (N_27085,N_26504,N_26988);
nor U27086 (N_27086,N_26906,N_26661);
nor U27087 (N_27087,N_26731,N_26771);
and U27088 (N_27088,N_26961,N_26612);
xnor U27089 (N_27089,N_26662,N_26954);
xor U27090 (N_27090,N_26891,N_26998);
nand U27091 (N_27091,N_26533,N_26685);
xor U27092 (N_27092,N_26638,N_26691);
and U27093 (N_27093,N_26554,N_26652);
nor U27094 (N_27094,N_26879,N_26522);
or U27095 (N_27095,N_26669,N_26863);
nand U27096 (N_27096,N_26977,N_26728);
xor U27097 (N_27097,N_26733,N_26814);
or U27098 (N_27098,N_26581,N_26753);
or U27099 (N_27099,N_26927,N_26735);
xor U27100 (N_27100,N_26628,N_26915);
or U27101 (N_27101,N_26840,N_26824);
xnor U27102 (N_27102,N_26935,N_26694);
nand U27103 (N_27103,N_26630,N_26585);
nand U27104 (N_27104,N_26990,N_26821);
or U27105 (N_27105,N_26752,N_26791);
nor U27106 (N_27106,N_26980,N_26839);
and U27107 (N_27107,N_26611,N_26582);
and U27108 (N_27108,N_26904,N_26660);
nor U27109 (N_27109,N_26786,N_26803);
or U27110 (N_27110,N_26828,N_26768);
and U27111 (N_27111,N_26825,N_26739);
xnor U27112 (N_27112,N_26552,N_26911);
or U27113 (N_27113,N_26555,N_26583);
xor U27114 (N_27114,N_26929,N_26591);
and U27115 (N_27115,N_26975,N_26806);
xor U27116 (N_27116,N_26778,N_26845);
nor U27117 (N_27117,N_26742,N_26684);
nor U27118 (N_27118,N_26889,N_26783);
nand U27119 (N_27119,N_26811,N_26963);
or U27120 (N_27120,N_26872,N_26899);
and U27121 (N_27121,N_26748,N_26507);
nand U27122 (N_27122,N_26972,N_26951);
nor U27123 (N_27123,N_26945,N_26703);
xnor U27124 (N_27124,N_26957,N_26527);
nor U27125 (N_27125,N_26644,N_26632);
nand U27126 (N_27126,N_26563,N_26898);
xnor U27127 (N_27127,N_26635,N_26702);
xnor U27128 (N_27128,N_26625,N_26812);
xor U27129 (N_27129,N_26973,N_26835);
nor U27130 (N_27130,N_26675,N_26559);
or U27131 (N_27131,N_26505,N_26777);
nor U27132 (N_27132,N_26917,N_26720);
nand U27133 (N_27133,N_26529,N_26512);
nor U27134 (N_27134,N_26599,N_26671);
or U27135 (N_27135,N_26653,N_26797);
and U27136 (N_27136,N_26802,N_26707);
or U27137 (N_27137,N_26962,N_26756);
nand U27138 (N_27138,N_26779,N_26809);
and U27139 (N_27139,N_26610,N_26897);
or U27140 (N_27140,N_26799,N_26510);
and U27141 (N_27141,N_26657,N_26823);
xnor U27142 (N_27142,N_26542,N_26579);
xor U27143 (N_27143,N_26939,N_26852);
or U27144 (N_27144,N_26964,N_26548);
and U27145 (N_27145,N_26847,N_26573);
nand U27146 (N_27146,N_26537,N_26936);
xor U27147 (N_27147,N_26536,N_26508);
nor U27148 (N_27148,N_26528,N_26511);
xnor U27149 (N_27149,N_26984,N_26577);
and U27150 (N_27150,N_26706,N_26819);
nand U27151 (N_27151,N_26727,N_26709);
xor U27152 (N_27152,N_26730,N_26816);
nor U27153 (N_27153,N_26521,N_26574);
nand U27154 (N_27154,N_26710,N_26770);
or U27155 (N_27155,N_26933,N_26804);
nor U27156 (N_27156,N_26595,N_26647);
and U27157 (N_27157,N_26697,N_26726);
nor U27158 (N_27158,N_26822,N_26887);
xnor U27159 (N_27159,N_26514,N_26993);
nor U27160 (N_27160,N_26575,N_26668);
and U27161 (N_27161,N_26997,N_26890);
xor U27162 (N_27162,N_26562,N_26861);
nand U27163 (N_27163,N_26886,N_26620);
or U27164 (N_27164,N_26594,N_26789);
xnor U27165 (N_27165,N_26818,N_26576);
and U27166 (N_27166,N_26754,N_26712);
nor U27167 (N_27167,N_26865,N_26912);
nand U27168 (N_27168,N_26856,N_26545);
or U27169 (N_27169,N_26907,N_26608);
or U27170 (N_27170,N_26895,N_26996);
nand U27171 (N_27171,N_26640,N_26938);
xor U27172 (N_27172,N_26843,N_26867);
nor U27173 (N_27173,N_26714,N_26837);
and U27174 (N_27174,N_26851,N_26893);
nor U27175 (N_27175,N_26755,N_26531);
and U27176 (N_27176,N_26623,N_26868);
and U27177 (N_27177,N_26787,N_26655);
or U27178 (N_27178,N_26544,N_26621);
and U27179 (N_27179,N_26699,N_26600);
or U27180 (N_27180,N_26571,N_26924);
xor U27181 (N_27181,N_26530,N_26877);
xnor U27182 (N_27182,N_26656,N_26654);
nand U27183 (N_27183,N_26978,N_26974);
or U27184 (N_27184,N_26905,N_26958);
or U27185 (N_27185,N_26693,N_26670);
and U27186 (N_27186,N_26567,N_26869);
nor U27187 (N_27187,N_26565,N_26700);
and U27188 (N_27188,N_26517,N_26629);
xor U27189 (N_27189,N_26991,N_26820);
xnor U27190 (N_27190,N_26833,N_26870);
nor U27191 (N_27191,N_26674,N_26732);
xnor U27192 (N_27192,N_26580,N_26827);
nor U27193 (N_27193,N_26619,N_26923);
xor U27194 (N_27194,N_26903,N_26930);
nand U27195 (N_27195,N_26950,N_26857);
xnor U27196 (N_27196,N_26557,N_26916);
and U27197 (N_27197,N_26502,N_26937);
nor U27198 (N_27198,N_26538,N_26792);
nor U27199 (N_27199,N_26914,N_26695);
or U27200 (N_27200,N_26672,N_26663);
and U27201 (N_27201,N_26513,N_26539);
xor U27202 (N_27202,N_26639,N_26773);
and U27203 (N_27203,N_26995,N_26637);
nor U27204 (N_27204,N_26831,N_26550);
nor U27205 (N_27205,N_26855,N_26952);
or U27206 (N_27206,N_26686,N_26934);
or U27207 (N_27207,N_26665,N_26894);
nor U27208 (N_27208,N_26992,N_26634);
and U27209 (N_27209,N_26931,N_26524);
xnor U27210 (N_27210,N_26607,N_26834);
xnor U27211 (N_27211,N_26862,N_26985);
nand U27212 (N_27212,N_26677,N_26734);
or U27213 (N_27213,N_26596,N_26842);
and U27214 (N_27214,N_26759,N_26636);
nor U27215 (N_27215,N_26875,N_26747);
nor U27216 (N_27216,N_26942,N_26969);
nor U27217 (N_27217,N_26678,N_26965);
and U27218 (N_27218,N_26701,N_26682);
nand U27219 (N_27219,N_26853,N_26740);
nand U27220 (N_27220,N_26989,N_26764);
and U27221 (N_27221,N_26850,N_26844);
or U27222 (N_27222,N_26830,N_26743);
nand U27223 (N_27223,N_26979,N_26601);
nand U27224 (N_27224,N_26981,N_26874);
or U27225 (N_27225,N_26680,N_26883);
or U27226 (N_27226,N_26736,N_26643);
or U27227 (N_27227,N_26794,N_26751);
nand U27228 (N_27228,N_26932,N_26946);
nand U27229 (N_27229,N_26729,N_26765);
nor U27230 (N_27230,N_26696,N_26880);
or U27231 (N_27231,N_26718,N_26626);
nand U27232 (N_27232,N_26715,N_26909);
nand U27233 (N_27233,N_26948,N_26758);
or U27234 (N_27234,N_26602,N_26598);
xnor U27235 (N_27235,N_26876,N_26808);
xor U27236 (N_27236,N_26986,N_26838);
and U27237 (N_27237,N_26556,N_26790);
nor U27238 (N_27238,N_26687,N_26722);
or U27239 (N_27239,N_26551,N_26941);
nor U27240 (N_27240,N_26723,N_26584);
nand U27241 (N_27241,N_26882,N_26500);
or U27242 (N_27242,N_26560,N_26866);
and U27243 (N_27243,N_26832,N_26532);
or U27244 (N_27244,N_26568,N_26525);
and U27245 (N_27245,N_26892,N_26597);
nand U27246 (N_27246,N_26578,N_26572);
nor U27247 (N_27247,N_26569,N_26622);
nand U27248 (N_27248,N_26631,N_26501);
xnor U27249 (N_27249,N_26871,N_26966);
nor U27250 (N_27250,N_26888,N_26702);
nand U27251 (N_27251,N_26908,N_26752);
and U27252 (N_27252,N_26673,N_26589);
nand U27253 (N_27253,N_26741,N_26539);
or U27254 (N_27254,N_26688,N_26903);
and U27255 (N_27255,N_26784,N_26524);
xnor U27256 (N_27256,N_26741,N_26792);
nor U27257 (N_27257,N_26613,N_26785);
nor U27258 (N_27258,N_26523,N_26959);
and U27259 (N_27259,N_26527,N_26895);
xnor U27260 (N_27260,N_26932,N_26956);
and U27261 (N_27261,N_26820,N_26959);
nand U27262 (N_27262,N_26820,N_26586);
and U27263 (N_27263,N_26578,N_26864);
nand U27264 (N_27264,N_26792,N_26931);
xnor U27265 (N_27265,N_26851,N_26564);
nand U27266 (N_27266,N_26584,N_26920);
and U27267 (N_27267,N_26765,N_26863);
nand U27268 (N_27268,N_26626,N_26636);
nor U27269 (N_27269,N_26627,N_26584);
nor U27270 (N_27270,N_26866,N_26862);
or U27271 (N_27271,N_26957,N_26886);
and U27272 (N_27272,N_26665,N_26601);
or U27273 (N_27273,N_26639,N_26514);
and U27274 (N_27274,N_26541,N_26746);
and U27275 (N_27275,N_26830,N_26669);
nand U27276 (N_27276,N_26974,N_26893);
xnor U27277 (N_27277,N_26994,N_26591);
and U27278 (N_27278,N_26793,N_26943);
nor U27279 (N_27279,N_26871,N_26656);
and U27280 (N_27280,N_26555,N_26607);
nand U27281 (N_27281,N_26594,N_26984);
nor U27282 (N_27282,N_26805,N_26775);
nor U27283 (N_27283,N_26652,N_26690);
and U27284 (N_27284,N_26903,N_26958);
or U27285 (N_27285,N_26781,N_26577);
xor U27286 (N_27286,N_26854,N_26618);
or U27287 (N_27287,N_26507,N_26864);
and U27288 (N_27288,N_26564,N_26506);
or U27289 (N_27289,N_26938,N_26759);
nor U27290 (N_27290,N_26825,N_26943);
or U27291 (N_27291,N_26997,N_26542);
xor U27292 (N_27292,N_26689,N_26783);
xor U27293 (N_27293,N_26858,N_26546);
xnor U27294 (N_27294,N_26661,N_26737);
and U27295 (N_27295,N_26862,N_26978);
or U27296 (N_27296,N_26915,N_26506);
nor U27297 (N_27297,N_26790,N_26849);
and U27298 (N_27298,N_26942,N_26512);
and U27299 (N_27299,N_26500,N_26723);
nor U27300 (N_27300,N_26942,N_26726);
xnor U27301 (N_27301,N_26972,N_26738);
or U27302 (N_27302,N_26560,N_26952);
nand U27303 (N_27303,N_26654,N_26867);
or U27304 (N_27304,N_26783,N_26584);
and U27305 (N_27305,N_26587,N_26715);
or U27306 (N_27306,N_26596,N_26686);
and U27307 (N_27307,N_26735,N_26724);
or U27308 (N_27308,N_26863,N_26648);
xor U27309 (N_27309,N_26820,N_26861);
or U27310 (N_27310,N_26644,N_26682);
and U27311 (N_27311,N_26822,N_26738);
xor U27312 (N_27312,N_26906,N_26850);
nand U27313 (N_27313,N_26796,N_26945);
nand U27314 (N_27314,N_26747,N_26548);
or U27315 (N_27315,N_26897,N_26522);
nand U27316 (N_27316,N_26729,N_26839);
xnor U27317 (N_27317,N_26727,N_26729);
xnor U27318 (N_27318,N_26960,N_26810);
nor U27319 (N_27319,N_26707,N_26899);
and U27320 (N_27320,N_26773,N_26582);
or U27321 (N_27321,N_26509,N_26961);
nor U27322 (N_27322,N_26938,N_26517);
xnor U27323 (N_27323,N_26811,N_26629);
and U27324 (N_27324,N_26802,N_26967);
or U27325 (N_27325,N_26601,N_26692);
nand U27326 (N_27326,N_26664,N_26789);
nor U27327 (N_27327,N_26953,N_26547);
nand U27328 (N_27328,N_26827,N_26500);
or U27329 (N_27329,N_26558,N_26741);
and U27330 (N_27330,N_26998,N_26955);
nor U27331 (N_27331,N_26667,N_26665);
nand U27332 (N_27332,N_26542,N_26881);
xnor U27333 (N_27333,N_26523,N_26724);
nor U27334 (N_27334,N_26843,N_26527);
xnor U27335 (N_27335,N_26577,N_26559);
and U27336 (N_27336,N_26867,N_26655);
xnor U27337 (N_27337,N_26988,N_26680);
and U27338 (N_27338,N_26846,N_26850);
nor U27339 (N_27339,N_26661,N_26968);
and U27340 (N_27340,N_26754,N_26907);
or U27341 (N_27341,N_26863,N_26561);
or U27342 (N_27342,N_26990,N_26811);
and U27343 (N_27343,N_26927,N_26840);
nand U27344 (N_27344,N_26584,N_26830);
nor U27345 (N_27345,N_26735,N_26937);
or U27346 (N_27346,N_26505,N_26753);
nand U27347 (N_27347,N_26934,N_26707);
and U27348 (N_27348,N_26613,N_26996);
xor U27349 (N_27349,N_26925,N_26580);
and U27350 (N_27350,N_26529,N_26790);
nor U27351 (N_27351,N_26954,N_26559);
and U27352 (N_27352,N_26569,N_26968);
nor U27353 (N_27353,N_26615,N_26942);
nand U27354 (N_27354,N_26580,N_26528);
nand U27355 (N_27355,N_26878,N_26823);
nor U27356 (N_27356,N_26729,N_26906);
nor U27357 (N_27357,N_26758,N_26862);
xor U27358 (N_27358,N_26529,N_26519);
and U27359 (N_27359,N_26881,N_26546);
nand U27360 (N_27360,N_26700,N_26803);
nor U27361 (N_27361,N_26679,N_26639);
nor U27362 (N_27362,N_26924,N_26959);
nor U27363 (N_27363,N_26537,N_26779);
and U27364 (N_27364,N_26542,N_26524);
nor U27365 (N_27365,N_26610,N_26939);
nand U27366 (N_27366,N_26629,N_26877);
nand U27367 (N_27367,N_26606,N_26602);
and U27368 (N_27368,N_26862,N_26923);
nand U27369 (N_27369,N_26535,N_26572);
and U27370 (N_27370,N_26878,N_26656);
xor U27371 (N_27371,N_26791,N_26645);
and U27372 (N_27372,N_26545,N_26627);
and U27373 (N_27373,N_26572,N_26858);
nand U27374 (N_27374,N_26704,N_26561);
or U27375 (N_27375,N_26705,N_26880);
xor U27376 (N_27376,N_26917,N_26708);
and U27377 (N_27377,N_26600,N_26676);
nor U27378 (N_27378,N_26980,N_26927);
nor U27379 (N_27379,N_26987,N_26926);
xor U27380 (N_27380,N_26653,N_26901);
nand U27381 (N_27381,N_26626,N_26701);
nor U27382 (N_27382,N_26870,N_26598);
or U27383 (N_27383,N_26799,N_26798);
xor U27384 (N_27384,N_26802,N_26709);
and U27385 (N_27385,N_26944,N_26916);
xnor U27386 (N_27386,N_26875,N_26829);
and U27387 (N_27387,N_26982,N_26555);
and U27388 (N_27388,N_26949,N_26589);
nor U27389 (N_27389,N_26746,N_26873);
nand U27390 (N_27390,N_26594,N_26897);
or U27391 (N_27391,N_26829,N_26985);
nand U27392 (N_27392,N_26955,N_26846);
nor U27393 (N_27393,N_26833,N_26986);
nand U27394 (N_27394,N_26680,N_26830);
and U27395 (N_27395,N_26627,N_26676);
xnor U27396 (N_27396,N_26724,N_26727);
xnor U27397 (N_27397,N_26893,N_26731);
xor U27398 (N_27398,N_26503,N_26715);
nor U27399 (N_27399,N_26957,N_26512);
nand U27400 (N_27400,N_26640,N_26676);
nand U27401 (N_27401,N_26521,N_26621);
nand U27402 (N_27402,N_26885,N_26543);
nand U27403 (N_27403,N_26543,N_26736);
or U27404 (N_27404,N_26881,N_26591);
or U27405 (N_27405,N_26546,N_26891);
nor U27406 (N_27406,N_26688,N_26707);
nand U27407 (N_27407,N_26578,N_26662);
or U27408 (N_27408,N_26897,N_26557);
and U27409 (N_27409,N_26988,N_26534);
or U27410 (N_27410,N_26528,N_26999);
nand U27411 (N_27411,N_26612,N_26883);
xnor U27412 (N_27412,N_26798,N_26795);
or U27413 (N_27413,N_26695,N_26504);
and U27414 (N_27414,N_26969,N_26517);
and U27415 (N_27415,N_26956,N_26794);
or U27416 (N_27416,N_26647,N_26639);
or U27417 (N_27417,N_26683,N_26903);
xnor U27418 (N_27418,N_26563,N_26817);
nor U27419 (N_27419,N_26754,N_26982);
xnor U27420 (N_27420,N_26680,N_26860);
xor U27421 (N_27421,N_26910,N_26757);
nand U27422 (N_27422,N_26947,N_26522);
or U27423 (N_27423,N_26863,N_26998);
nor U27424 (N_27424,N_26544,N_26615);
nand U27425 (N_27425,N_26679,N_26501);
or U27426 (N_27426,N_26719,N_26562);
and U27427 (N_27427,N_26724,N_26620);
xnor U27428 (N_27428,N_26671,N_26911);
nor U27429 (N_27429,N_26648,N_26757);
and U27430 (N_27430,N_26861,N_26658);
or U27431 (N_27431,N_26947,N_26795);
nand U27432 (N_27432,N_26572,N_26618);
nor U27433 (N_27433,N_26641,N_26804);
nor U27434 (N_27434,N_26586,N_26525);
xnor U27435 (N_27435,N_26778,N_26592);
xnor U27436 (N_27436,N_26982,N_26953);
nand U27437 (N_27437,N_26945,N_26873);
xor U27438 (N_27438,N_26911,N_26823);
and U27439 (N_27439,N_26671,N_26718);
nand U27440 (N_27440,N_26567,N_26896);
and U27441 (N_27441,N_26636,N_26751);
nor U27442 (N_27442,N_26657,N_26780);
nor U27443 (N_27443,N_26537,N_26890);
nor U27444 (N_27444,N_26544,N_26570);
nand U27445 (N_27445,N_26571,N_26878);
nor U27446 (N_27446,N_26688,N_26997);
and U27447 (N_27447,N_26640,N_26905);
xnor U27448 (N_27448,N_26547,N_26862);
xor U27449 (N_27449,N_26760,N_26684);
or U27450 (N_27450,N_26513,N_26832);
xnor U27451 (N_27451,N_26671,N_26504);
nor U27452 (N_27452,N_26587,N_26626);
nor U27453 (N_27453,N_26823,N_26642);
xor U27454 (N_27454,N_26808,N_26972);
xor U27455 (N_27455,N_26741,N_26818);
nand U27456 (N_27456,N_26782,N_26765);
and U27457 (N_27457,N_26799,N_26906);
nand U27458 (N_27458,N_26728,N_26638);
nor U27459 (N_27459,N_26742,N_26933);
xnor U27460 (N_27460,N_26846,N_26912);
and U27461 (N_27461,N_26922,N_26762);
nand U27462 (N_27462,N_26986,N_26887);
nand U27463 (N_27463,N_26657,N_26798);
or U27464 (N_27464,N_26932,N_26582);
nor U27465 (N_27465,N_26548,N_26627);
nor U27466 (N_27466,N_26670,N_26964);
or U27467 (N_27467,N_26803,N_26730);
and U27468 (N_27468,N_26509,N_26649);
and U27469 (N_27469,N_26836,N_26597);
and U27470 (N_27470,N_26606,N_26840);
nor U27471 (N_27471,N_26743,N_26531);
or U27472 (N_27472,N_26870,N_26992);
and U27473 (N_27473,N_26791,N_26921);
and U27474 (N_27474,N_26820,N_26501);
xnor U27475 (N_27475,N_26890,N_26995);
nor U27476 (N_27476,N_26757,N_26526);
nand U27477 (N_27477,N_26586,N_26528);
and U27478 (N_27478,N_26684,N_26838);
xor U27479 (N_27479,N_26799,N_26556);
xor U27480 (N_27480,N_26753,N_26806);
or U27481 (N_27481,N_26982,N_26810);
or U27482 (N_27482,N_26744,N_26674);
xor U27483 (N_27483,N_26557,N_26600);
xor U27484 (N_27484,N_26678,N_26675);
and U27485 (N_27485,N_26557,N_26992);
nand U27486 (N_27486,N_26575,N_26999);
nor U27487 (N_27487,N_26715,N_26737);
nand U27488 (N_27488,N_26569,N_26879);
nand U27489 (N_27489,N_26735,N_26622);
xnor U27490 (N_27490,N_26978,N_26993);
nand U27491 (N_27491,N_26833,N_26937);
nor U27492 (N_27492,N_26725,N_26998);
and U27493 (N_27493,N_26558,N_26613);
and U27494 (N_27494,N_26869,N_26940);
nor U27495 (N_27495,N_26949,N_26520);
xnor U27496 (N_27496,N_26613,N_26920);
and U27497 (N_27497,N_26596,N_26640);
or U27498 (N_27498,N_26926,N_26684);
or U27499 (N_27499,N_26987,N_26784);
and U27500 (N_27500,N_27317,N_27397);
xnor U27501 (N_27501,N_27056,N_27309);
and U27502 (N_27502,N_27421,N_27346);
or U27503 (N_27503,N_27043,N_27306);
xor U27504 (N_27504,N_27032,N_27206);
xnor U27505 (N_27505,N_27130,N_27044);
nand U27506 (N_27506,N_27235,N_27188);
or U27507 (N_27507,N_27041,N_27046);
nor U27508 (N_27508,N_27377,N_27245);
or U27509 (N_27509,N_27211,N_27148);
nor U27510 (N_27510,N_27458,N_27120);
xnor U27511 (N_27511,N_27145,N_27368);
nor U27512 (N_27512,N_27493,N_27000);
or U27513 (N_27513,N_27395,N_27327);
xor U27514 (N_27514,N_27129,N_27010);
nand U27515 (N_27515,N_27385,N_27269);
nor U27516 (N_27516,N_27031,N_27356);
and U27517 (N_27517,N_27381,N_27142);
and U27518 (N_27518,N_27001,N_27020);
and U27519 (N_27519,N_27181,N_27132);
xor U27520 (N_27520,N_27049,N_27141);
nor U27521 (N_27521,N_27413,N_27326);
and U27522 (N_27522,N_27402,N_27495);
nor U27523 (N_27523,N_27399,N_27164);
nand U27524 (N_27524,N_27076,N_27005);
and U27525 (N_27525,N_27186,N_27113);
and U27526 (N_27526,N_27270,N_27171);
xnor U27527 (N_27527,N_27218,N_27446);
nor U27528 (N_27528,N_27424,N_27404);
and U27529 (N_27529,N_27344,N_27236);
xnor U27530 (N_27530,N_27203,N_27192);
xor U27531 (N_27531,N_27105,N_27065);
or U27532 (N_27532,N_27061,N_27304);
or U27533 (N_27533,N_27386,N_27284);
or U27534 (N_27534,N_27166,N_27004);
or U27535 (N_27535,N_27250,N_27018);
nand U27536 (N_27536,N_27372,N_27467);
xor U27537 (N_27537,N_27289,N_27299);
nor U27538 (N_27538,N_27360,N_27419);
nor U27539 (N_27539,N_27168,N_27311);
or U27540 (N_27540,N_27263,N_27152);
nor U27541 (N_27541,N_27157,N_27231);
or U27542 (N_27542,N_27465,N_27143);
nor U27543 (N_27543,N_27335,N_27095);
xor U27544 (N_27544,N_27430,N_27025);
nand U27545 (N_27545,N_27334,N_27225);
or U27546 (N_27546,N_27273,N_27449);
and U27547 (N_27547,N_27092,N_27472);
and U27548 (N_27548,N_27229,N_27414);
nor U27549 (N_27549,N_27153,N_27341);
nor U27550 (N_27550,N_27055,N_27349);
nor U27551 (N_27551,N_27242,N_27007);
nor U27552 (N_27552,N_27185,N_27103);
nor U27553 (N_27553,N_27451,N_27321);
or U27554 (N_27554,N_27212,N_27305);
or U27555 (N_27555,N_27358,N_27286);
nor U27556 (N_27556,N_27050,N_27114);
or U27557 (N_27557,N_27371,N_27134);
nor U27558 (N_27558,N_27183,N_27175);
and U27559 (N_27559,N_27325,N_27400);
and U27560 (N_27560,N_27080,N_27057);
or U27561 (N_27561,N_27329,N_27408);
xor U27562 (N_27562,N_27379,N_27111);
and U27563 (N_27563,N_27462,N_27337);
nor U27564 (N_27564,N_27352,N_27180);
xor U27565 (N_27565,N_27075,N_27297);
or U27566 (N_27566,N_27131,N_27435);
or U27567 (N_27567,N_27355,N_27336);
nand U27568 (N_27568,N_27087,N_27473);
xor U27569 (N_27569,N_27084,N_27301);
or U27570 (N_27570,N_27322,N_27471);
nand U27571 (N_27571,N_27416,N_27288);
nand U27572 (N_27572,N_27121,N_27478);
nor U27573 (N_27573,N_27228,N_27072);
nand U27574 (N_27574,N_27077,N_27066);
and U27575 (N_27575,N_27330,N_27173);
and U27576 (N_27576,N_27222,N_27314);
and U27577 (N_27577,N_27394,N_27426);
nand U27578 (N_27578,N_27194,N_27441);
or U27579 (N_27579,N_27088,N_27237);
and U27580 (N_27580,N_27323,N_27078);
nor U27581 (N_27581,N_27362,N_27215);
nor U27582 (N_27582,N_27124,N_27115);
xnor U27583 (N_27583,N_27223,N_27047);
and U27584 (N_27584,N_27177,N_27474);
nand U27585 (N_27585,N_27182,N_27489);
nand U27586 (N_27586,N_27476,N_27445);
nor U27587 (N_27587,N_27436,N_27195);
nand U27588 (N_27588,N_27102,N_27276);
and U27589 (N_27589,N_27285,N_27407);
nand U27590 (N_27590,N_27375,N_27331);
and U27591 (N_27591,N_27221,N_27280);
nor U27592 (N_27592,N_27296,N_27147);
nand U27593 (N_27593,N_27359,N_27108);
nor U27594 (N_27594,N_27428,N_27251);
nand U27595 (N_27595,N_27008,N_27415);
xnor U27596 (N_27596,N_27378,N_27461);
and U27597 (N_27597,N_27324,N_27468);
nand U27598 (N_27598,N_27492,N_27174);
or U27599 (N_27599,N_27275,N_27483);
nand U27600 (N_27600,N_27079,N_27442);
xor U27601 (N_27601,N_27035,N_27023);
nand U27602 (N_27602,N_27318,N_27213);
xor U27603 (N_27603,N_27156,N_27135);
or U27604 (N_27604,N_27083,N_27128);
and U27605 (N_27605,N_27034,N_27040);
nand U27606 (N_27606,N_27015,N_27464);
xnor U27607 (N_27607,N_27019,N_27205);
xor U27608 (N_27608,N_27012,N_27369);
xor U27609 (N_27609,N_27179,N_27294);
xor U27610 (N_27610,N_27351,N_27112);
nand U27611 (N_27611,N_27028,N_27137);
nand U27612 (N_27612,N_27466,N_27382);
and U27613 (N_27613,N_27456,N_27283);
nor U27614 (N_27614,N_27315,N_27051);
and U27615 (N_27615,N_27373,N_27059);
or U27616 (N_27616,N_27367,N_27486);
nor U27617 (N_27617,N_27443,N_27067);
xnor U27618 (N_27618,N_27074,N_27470);
nand U27619 (N_27619,N_27405,N_27234);
xnor U27620 (N_27620,N_27053,N_27265);
xnor U27621 (N_27621,N_27214,N_27350);
nor U27622 (N_27622,N_27406,N_27479);
xnor U27623 (N_27623,N_27126,N_27313);
and U27624 (N_27624,N_27006,N_27338);
xnor U27625 (N_27625,N_27440,N_27271);
nand U27626 (N_27626,N_27298,N_27432);
nor U27627 (N_27627,N_27480,N_27396);
or U27628 (N_27628,N_27310,N_27401);
or U27629 (N_27629,N_27009,N_27209);
nand U27630 (N_27630,N_27016,N_27160);
and U27631 (N_27631,N_27427,N_27189);
xnor U27632 (N_27632,N_27264,N_27151);
or U27633 (N_27633,N_27496,N_27398);
xor U27634 (N_27634,N_27048,N_27253);
nor U27635 (N_27635,N_27249,N_27425);
nor U27636 (N_27636,N_27109,N_27256);
xor U27637 (N_27637,N_27477,N_27469);
nand U27638 (N_27638,N_27190,N_27450);
xor U27639 (N_27639,N_27150,N_27252);
xor U27640 (N_27640,N_27353,N_27187);
nand U27641 (N_27641,N_27193,N_27411);
xnor U27642 (N_27642,N_27343,N_27376);
nand U27643 (N_27643,N_27233,N_27030);
nor U27644 (N_27644,N_27122,N_27054);
or U27645 (N_27645,N_27481,N_27340);
xor U27646 (N_27646,N_27199,N_27033);
xor U27647 (N_27647,N_27100,N_27163);
nand U27648 (N_27648,N_27014,N_27063);
and U27649 (N_27649,N_27319,N_27482);
nand U27650 (N_27650,N_27333,N_27200);
or U27651 (N_27651,N_27073,N_27403);
nand U27652 (N_27652,N_27365,N_27244);
and U27653 (N_27653,N_27216,N_27107);
and U27654 (N_27654,N_27261,N_27140);
nor U27655 (N_27655,N_27230,N_27279);
xor U27656 (N_27656,N_27312,N_27258);
nor U27657 (N_27657,N_27239,N_27259);
and U27658 (N_27658,N_27347,N_27197);
or U27659 (N_27659,N_27454,N_27292);
nand U27660 (N_27660,N_27138,N_27433);
nor U27661 (N_27661,N_27219,N_27307);
and U27662 (N_27662,N_27159,N_27452);
nor U27663 (N_27663,N_27434,N_27437);
or U27664 (N_27664,N_27184,N_27494);
nand U27665 (N_27665,N_27118,N_27220);
and U27666 (N_27666,N_27070,N_27420);
nor U27667 (N_27667,N_27243,N_27011);
xor U27668 (N_27668,N_27453,N_27257);
xor U27669 (N_27669,N_27170,N_27475);
or U27670 (N_27670,N_27086,N_27149);
and U27671 (N_27671,N_27045,N_27277);
and U27672 (N_27672,N_27062,N_27392);
and U27673 (N_27673,N_27255,N_27320);
xnor U27674 (N_27674,N_27262,N_27499);
or U27675 (N_27675,N_27422,N_27345);
xor U27676 (N_27676,N_27278,N_27357);
or U27677 (N_27677,N_27017,N_27463);
nor U27678 (N_27678,N_27207,N_27429);
or U27679 (N_27679,N_27022,N_27300);
nor U27680 (N_27680,N_27106,N_27232);
nor U27681 (N_27681,N_27196,N_27096);
nor U27682 (N_27682,N_27354,N_27390);
or U27683 (N_27683,N_27418,N_27364);
or U27684 (N_27684,N_27423,N_27052);
nor U27685 (N_27685,N_27363,N_27328);
or U27686 (N_27686,N_27457,N_27178);
nor U27687 (N_27687,N_27144,N_27487);
or U27688 (N_27688,N_27417,N_27455);
nand U27689 (N_27689,N_27302,N_27202);
and U27690 (N_27690,N_27042,N_27295);
and U27691 (N_27691,N_27036,N_27497);
nand U27692 (N_27692,N_27162,N_27094);
or U27693 (N_27693,N_27391,N_27217);
nand U27694 (N_27694,N_27133,N_27388);
nor U27695 (N_27695,N_27332,N_27389);
or U27696 (N_27696,N_27260,N_27161);
and U27697 (N_27697,N_27091,N_27082);
and U27698 (N_27698,N_27348,N_27116);
nand U27699 (N_27699,N_27387,N_27117);
or U27700 (N_27700,N_27123,N_27316);
xnor U27701 (N_27701,N_27060,N_27021);
or U27702 (N_27702,N_27029,N_27238);
nand U27703 (N_27703,N_27240,N_27058);
nor U27704 (N_27704,N_27498,N_27104);
xor U27705 (N_27705,N_27410,N_27127);
or U27706 (N_27706,N_27068,N_27383);
and U27707 (N_27707,N_27460,N_27085);
or U27708 (N_27708,N_27291,N_27393);
nor U27709 (N_27709,N_27267,N_27038);
or U27710 (N_27710,N_27201,N_27254);
nand U27711 (N_27711,N_27227,N_27125);
and U27712 (N_27712,N_27266,N_27303);
nor U27713 (N_27713,N_27158,N_27093);
xnor U27714 (N_27714,N_27241,N_27274);
xor U27715 (N_27715,N_27069,N_27169);
or U27716 (N_27716,N_27226,N_27101);
nand U27717 (N_27717,N_27064,N_27099);
nor U27718 (N_27718,N_27281,N_27380);
and U27719 (N_27719,N_27342,N_27308);
nor U27720 (N_27720,N_27272,N_27119);
nor U27721 (N_27721,N_27039,N_27037);
or U27722 (N_27722,N_27110,N_27282);
nand U27723 (N_27723,N_27439,N_27136);
and U27724 (N_27724,N_27090,N_27155);
nand U27725 (N_27725,N_27172,N_27459);
nand U27726 (N_27726,N_27210,N_27191);
nand U27727 (N_27727,N_27013,N_27208);
nand U27728 (N_27728,N_27290,N_27361);
nand U27729 (N_27729,N_27248,N_27268);
xor U27730 (N_27730,N_27293,N_27139);
xor U27731 (N_27731,N_27485,N_27490);
xnor U27732 (N_27732,N_27409,N_27438);
nand U27733 (N_27733,N_27002,N_27024);
nand U27734 (N_27734,N_27370,N_27154);
nor U27735 (N_27735,N_27491,N_27098);
xnor U27736 (N_27736,N_27412,N_27431);
or U27737 (N_27737,N_27448,N_27484);
nand U27738 (N_27738,N_27339,N_27146);
nor U27739 (N_27739,N_27198,N_27081);
xnor U27740 (N_27740,N_27176,N_27165);
xnor U27741 (N_27741,N_27097,N_27366);
xor U27742 (N_27742,N_27167,N_27026);
or U27743 (N_27743,N_27384,N_27247);
and U27744 (N_27744,N_27287,N_27444);
xnor U27745 (N_27745,N_27488,N_27224);
or U27746 (N_27746,N_27374,N_27003);
xor U27747 (N_27747,N_27447,N_27089);
or U27748 (N_27748,N_27071,N_27027);
and U27749 (N_27749,N_27246,N_27204);
xnor U27750 (N_27750,N_27222,N_27098);
nand U27751 (N_27751,N_27103,N_27049);
nand U27752 (N_27752,N_27242,N_27460);
and U27753 (N_27753,N_27461,N_27284);
xnor U27754 (N_27754,N_27081,N_27496);
and U27755 (N_27755,N_27199,N_27244);
nand U27756 (N_27756,N_27035,N_27136);
nor U27757 (N_27757,N_27311,N_27120);
xor U27758 (N_27758,N_27384,N_27131);
nor U27759 (N_27759,N_27467,N_27114);
or U27760 (N_27760,N_27437,N_27202);
nor U27761 (N_27761,N_27056,N_27223);
or U27762 (N_27762,N_27487,N_27083);
nand U27763 (N_27763,N_27134,N_27322);
nand U27764 (N_27764,N_27023,N_27449);
nand U27765 (N_27765,N_27436,N_27322);
or U27766 (N_27766,N_27193,N_27268);
nor U27767 (N_27767,N_27135,N_27309);
nor U27768 (N_27768,N_27391,N_27349);
nand U27769 (N_27769,N_27153,N_27181);
nor U27770 (N_27770,N_27070,N_27308);
nand U27771 (N_27771,N_27193,N_27267);
xnor U27772 (N_27772,N_27181,N_27419);
or U27773 (N_27773,N_27042,N_27173);
or U27774 (N_27774,N_27442,N_27227);
or U27775 (N_27775,N_27356,N_27267);
or U27776 (N_27776,N_27335,N_27313);
xor U27777 (N_27777,N_27149,N_27228);
nand U27778 (N_27778,N_27069,N_27055);
xor U27779 (N_27779,N_27461,N_27363);
nor U27780 (N_27780,N_27377,N_27200);
nand U27781 (N_27781,N_27152,N_27310);
nor U27782 (N_27782,N_27269,N_27374);
or U27783 (N_27783,N_27069,N_27091);
xnor U27784 (N_27784,N_27438,N_27167);
or U27785 (N_27785,N_27291,N_27026);
xnor U27786 (N_27786,N_27353,N_27074);
nor U27787 (N_27787,N_27182,N_27417);
nor U27788 (N_27788,N_27036,N_27139);
xnor U27789 (N_27789,N_27235,N_27244);
and U27790 (N_27790,N_27307,N_27408);
xor U27791 (N_27791,N_27085,N_27307);
and U27792 (N_27792,N_27010,N_27476);
nand U27793 (N_27793,N_27471,N_27108);
or U27794 (N_27794,N_27281,N_27172);
or U27795 (N_27795,N_27352,N_27183);
nand U27796 (N_27796,N_27032,N_27452);
xnor U27797 (N_27797,N_27087,N_27421);
or U27798 (N_27798,N_27179,N_27094);
or U27799 (N_27799,N_27085,N_27234);
and U27800 (N_27800,N_27173,N_27216);
xnor U27801 (N_27801,N_27448,N_27089);
nor U27802 (N_27802,N_27408,N_27194);
or U27803 (N_27803,N_27262,N_27059);
and U27804 (N_27804,N_27465,N_27033);
nand U27805 (N_27805,N_27113,N_27273);
or U27806 (N_27806,N_27419,N_27300);
nand U27807 (N_27807,N_27152,N_27385);
xnor U27808 (N_27808,N_27322,N_27357);
xnor U27809 (N_27809,N_27046,N_27077);
or U27810 (N_27810,N_27143,N_27397);
and U27811 (N_27811,N_27049,N_27325);
and U27812 (N_27812,N_27455,N_27121);
nand U27813 (N_27813,N_27435,N_27445);
or U27814 (N_27814,N_27077,N_27105);
and U27815 (N_27815,N_27172,N_27417);
nor U27816 (N_27816,N_27415,N_27440);
or U27817 (N_27817,N_27171,N_27341);
xnor U27818 (N_27818,N_27094,N_27309);
nand U27819 (N_27819,N_27469,N_27121);
nor U27820 (N_27820,N_27347,N_27388);
or U27821 (N_27821,N_27417,N_27286);
nor U27822 (N_27822,N_27155,N_27434);
nor U27823 (N_27823,N_27239,N_27487);
or U27824 (N_27824,N_27365,N_27043);
and U27825 (N_27825,N_27202,N_27241);
nand U27826 (N_27826,N_27455,N_27340);
and U27827 (N_27827,N_27376,N_27373);
nand U27828 (N_27828,N_27247,N_27179);
nand U27829 (N_27829,N_27067,N_27216);
and U27830 (N_27830,N_27380,N_27279);
or U27831 (N_27831,N_27435,N_27114);
and U27832 (N_27832,N_27432,N_27046);
nand U27833 (N_27833,N_27011,N_27009);
and U27834 (N_27834,N_27463,N_27226);
and U27835 (N_27835,N_27134,N_27117);
nand U27836 (N_27836,N_27032,N_27266);
nand U27837 (N_27837,N_27320,N_27191);
and U27838 (N_27838,N_27498,N_27444);
and U27839 (N_27839,N_27087,N_27207);
xnor U27840 (N_27840,N_27146,N_27162);
and U27841 (N_27841,N_27245,N_27447);
nand U27842 (N_27842,N_27470,N_27346);
nand U27843 (N_27843,N_27496,N_27277);
nand U27844 (N_27844,N_27437,N_27397);
nand U27845 (N_27845,N_27022,N_27262);
xor U27846 (N_27846,N_27348,N_27401);
nor U27847 (N_27847,N_27010,N_27265);
nand U27848 (N_27848,N_27025,N_27329);
nor U27849 (N_27849,N_27094,N_27446);
xnor U27850 (N_27850,N_27137,N_27441);
and U27851 (N_27851,N_27354,N_27200);
nor U27852 (N_27852,N_27251,N_27094);
and U27853 (N_27853,N_27171,N_27445);
and U27854 (N_27854,N_27221,N_27479);
nor U27855 (N_27855,N_27061,N_27047);
xnor U27856 (N_27856,N_27070,N_27094);
and U27857 (N_27857,N_27210,N_27308);
nor U27858 (N_27858,N_27387,N_27041);
xor U27859 (N_27859,N_27444,N_27098);
or U27860 (N_27860,N_27131,N_27109);
xor U27861 (N_27861,N_27017,N_27095);
nand U27862 (N_27862,N_27031,N_27195);
nand U27863 (N_27863,N_27293,N_27100);
xor U27864 (N_27864,N_27375,N_27397);
nand U27865 (N_27865,N_27076,N_27230);
xor U27866 (N_27866,N_27432,N_27234);
nor U27867 (N_27867,N_27036,N_27226);
nor U27868 (N_27868,N_27422,N_27061);
xnor U27869 (N_27869,N_27475,N_27470);
nand U27870 (N_27870,N_27275,N_27324);
nand U27871 (N_27871,N_27421,N_27386);
xor U27872 (N_27872,N_27435,N_27176);
nand U27873 (N_27873,N_27322,N_27426);
nor U27874 (N_27874,N_27191,N_27174);
xnor U27875 (N_27875,N_27384,N_27066);
xor U27876 (N_27876,N_27095,N_27499);
nand U27877 (N_27877,N_27305,N_27267);
and U27878 (N_27878,N_27373,N_27361);
and U27879 (N_27879,N_27132,N_27367);
nor U27880 (N_27880,N_27217,N_27477);
or U27881 (N_27881,N_27076,N_27243);
nor U27882 (N_27882,N_27229,N_27022);
xor U27883 (N_27883,N_27072,N_27306);
nand U27884 (N_27884,N_27158,N_27003);
nor U27885 (N_27885,N_27144,N_27314);
nand U27886 (N_27886,N_27339,N_27456);
xnor U27887 (N_27887,N_27460,N_27381);
or U27888 (N_27888,N_27236,N_27258);
xor U27889 (N_27889,N_27473,N_27241);
xor U27890 (N_27890,N_27405,N_27091);
and U27891 (N_27891,N_27070,N_27491);
or U27892 (N_27892,N_27104,N_27469);
nor U27893 (N_27893,N_27213,N_27046);
nor U27894 (N_27894,N_27020,N_27314);
xor U27895 (N_27895,N_27082,N_27464);
and U27896 (N_27896,N_27106,N_27040);
and U27897 (N_27897,N_27481,N_27442);
xnor U27898 (N_27898,N_27272,N_27111);
nor U27899 (N_27899,N_27020,N_27359);
xor U27900 (N_27900,N_27331,N_27124);
nor U27901 (N_27901,N_27342,N_27069);
xor U27902 (N_27902,N_27095,N_27272);
and U27903 (N_27903,N_27495,N_27020);
or U27904 (N_27904,N_27262,N_27019);
xor U27905 (N_27905,N_27453,N_27223);
or U27906 (N_27906,N_27322,N_27298);
xor U27907 (N_27907,N_27447,N_27248);
and U27908 (N_27908,N_27445,N_27193);
nand U27909 (N_27909,N_27451,N_27222);
nor U27910 (N_27910,N_27383,N_27445);
or U27911 (N_27911,N_27237,N_27058);
nand U27912 (N_27912,N_27352,N_27069);
and U27913 (N_27913,N_27408,N_27226);
and U27914 (N_27914,N_27135,N_27176);
nand U27915 (N_27915,N_27385,N_27439);
nor U27916 (N_27916,N_27415,N_27489);
nand U27917 (N_27917,N_27408,N_27366);
or U27918 (N_27918,N_27166,N_27099);
and U27919 (N_27919,N_27131,N_27345);
and U27920 (N_27920,N_27428,N_27147);
xnor U27921 (N_27921,N_27220,N_27341);
and U27922 (N_27922,N_27461,N_27140);
and U27923 (N_27923,N_27065,N_27469);
and U27924 (N_27924,N_27429,N_27039);
xnor U27925 (N_27925,N_27419,N_27227);
xnor U27926 (N_27926,N_27041,N_27410);
nand U27927 (N_27927,N_27421,N_27191);
and U27928 (N_27928,N_27190,N_27154);
or U27929 (N_27929,N_27070,N_27067);
xnor U27930 (N_27930,N_27342,N_27424);
xor U27931 (N_27931,N_27192,N_27385);
nand U27932 (N_27932,N_27229,N_27495);
or U27933 (N_27933,N_27011,N_27186);
nand U27934 (N_27934,N_27409,N_27364);
nand U27935 (N_27935,N_27255,N_27353);
or U27936 (N_27936,N_27144,N_27149);
and U27937 (N_27937,N_27429,N_27460);
xor U27938 (N_27938,N_27286,N_27204);
nor U27939 (N_27939,N_27176,N_27424);
xor U27940 (N_27940,N_27005,N_27127);
nor U27941 (N_27941,N_27195,N_27035);
or U27942 (N_27942,N_27291,N_27227);
xnor U27943 (N_27943,N_27269,N_27475);
nor U27944 (N_27944,N_27047,N_27153);
nor U27945 (N_27945,N_27419,N_27231);
or U27946 (N_27946,N_27290,N_27225);
xor U27947 (N_27947,N_27012,N_27121);
and U27948 (N_27948,N_27489,N_27198);
nand U27949 (N_27949,N_27127,N_27368);
or U27950 (N_27950,N_27249,N_27183);
or U27951 (N_27951,N_27051,N_27117);
or U27952 (N_27952,N_27269,N_27294);
nor U27953 (N_27953,N_27339,N_27190);
nor U27954 (N_27954,N_27121,N_27365);
or U27955 (N_27955,N_27371,N_27482);
and U27956 (N_27956,N_27108,N_27389);
and U27957 (N_27957,N_27361,N_27357);
nand U27958 (N_27958,N_27063,N_27086);
or U27959 (N_27959,N_27233,N_27435);
or U27960 (N_27960,N_27092,N_27382);
or U27961 (N_27961,N_27314,N_27279);
nand U27962 (N_27962,N_27476,N_27246);
and U27963 (N_27963,N_27068,N_27029);
nor U27964 (N_27964,N_27133,N_27069);
and U27965 (N_27965,N_27083,N_27007);
nand U27966 (N_27966,N_27017,N_27456);
nand U27967 (N_27967,N_27118,N_27244);
nand U27968 (N_27968,N_27468,N_27454);
nor U27969 (N_27969,N_27060,N_27367);
nor U27970 (N_27970,N_27227,N_27140);
or U27971 (N_27971,N_27042,N_27414);
or U27972 (N_27972,N_27216,N_27315);
nor U27973 (N_27973,N_27466,N_27056);
and U27974 (N_27974,N_27433,N_27372);
xor U27975 (N_27975,N_27169,N_27150);
or U27976 (N_27976,N_27139,N_27287);
and U27977 (N_27977,N_27047,N_27221);
and U27978 (N_27978,N_27022,N_27027);
or U27979 (N_27979,N_27473,N_27151);
or U27980 (N_27980,N_27290,N_27252);
or U27981 (N_27981,N_27011,N_27437);
or U27982 (N_27982,N_27441,N_27413);
nand U27983 (N_27983,N_27425,N_27299);
or U27984 (N_27984,N_27476,N_27494);
and U27985 (N_27985,N_27271,N_27126);
or U27986 (N_27986,N_27445,N_27312);
nor U27987 (N_27987,N_27251,N_27453);
or U27988 (N_27988,N_27103,N_27221);
nor U27989 (N_27989,N_27261,N_27293);
nor U27990 (N_27990,N_27478,N_27269);
nand U27991 (N_27991,N_27429,N_27067);
nand U27992 (N_27992,N_27107,N_27034);
and U27993 (N_27993,N_27356,N_27064);
nand U27994 (N_27994,N_27283,N_27288);
nand U27995 (N_27995,N_27078,N_27022);
nand U27996 (N_27996,N_27474,N_27311);
xnor U27997 (N_27997,N_27489,N_27081);
xnor U27998 (N_27998,N_27013,N_27391);
and U27999 (N_27999,N_27374,N_27207);
xnor U28000 (N_28000,N_27506,N_27648);
and U28001 (N_28001,N_27689,N_27666);
and U28002 (N_28002,N_27589,N_27528);
nor U28003 (N_28003,N_27984,N_27928);
nand U28004 (N_28004,N_27711,N_27995);
nand U28005 (N_28005,N_27594,N_27608);
or U28006 (N_28006,N_27969,N_27722);
nand U28007 (N_28007,N_27684,N_27777);
nor U28008 (N_28008,N_27664,N_27858);
or U28009 (N_28009,N_27755,N_27951);
xor U28010 (N_28010,N_27855,N_27500);
or U28011 (N_28011,N_27670,N_27844);
or U28012 (N_28012,N_27571,N_27687);
nand U28013 (N_28013,N_27636,N_27526);
nor U28014 (N_28014,N_27748,N_27902);
xor U28015 (N_28015,N_27899,N_27929);
xnor U28016 (N_28016,N_27716,N_27904);
and U28017 (N_28017,N_27602,N_27574);
and U28018 (N_28018,N_27575,N_27629);
nor U28019 (N_28019,N_27637,N_27980);
and U28020 (N_28020,N_27515,N_27861);
xor U28021 (N_28021,N_27603,N_27559);
xor U28022 (N_28022,N_27618,N_27701);
or U28023 (N_28023,N_27894,N_27531);
nor U28024 (N_28024,N_27662,N_27849);
nand U28025 (N_28025,N_27974,N_27549);
xor U28026 (N_28026,N_27674,N_27593);
or U28027 (N_28027,N_27931,N_27856);
xor U28028 (N_28028,N_27516,N_27685);
nor U28029 (N_28029,N_27600,N_27992);
nand U28030 (N_28030,N_27839,N_27537);
nand U28031 (N_28031,N_27966,N_27923);
nor U28032 (N_28032,N_27671,N_27634);
xor U28033 (N_28033,N_27681,N_27833);
nand U28034 (N_28034,N_27805,N_27884);
xor U28035 (N_28035,N_27955,N_27783);
and U28036 (N_28036,N_27732,N_27617);
nor U28037 (N_28037,N_27622,N_27672);
and U28038 (N_28038,N_27819,N_27991);
nor U28039 (N_28039,N_27640,N_27870);
or U28040 (N_28040,N_27556,N_27609);
nand U28041 (N_28041,N_27652,N_27815);
nand U28042 (N_28042,N_27802,N_27898);
nor U28043 (N_28043,N_27772,N_27958);
and U28044 (N_28044,N_27832,N_27744);
and U28045 (N_28045,N_27621,N_27710);
xor U28046 (N_28046,N_27859,N_27520);
and U28047 (N_28047,N_27665,N_27869);
nor U28048 (N_28048,N_27768,N_27653);
xnor U28049 (N_28049,N_27718,N_27809);
or U28050 (N_28050,N_27543,N_27713);
and U28051 (N_28051,N_27623,N_27517);
xor U28052 (N_28052,N_27646,N_27763);
nand U28053 (N_28053,N_27838,N_27889);
or U28054 (N_28054,N_27654,N_27503);
or U28055 (N_28055,N_27780,N_27935);
and U28056 (N_28056,N_27836,N_27944);
and U28057 (N_28057,N_27605,N_27961);
xnor U28058 (N_28058,N_27900,N_27530);
and U28059 (N_28059,N_27746,N_27803);
and U28060 (N_28060,N_27667,N_27552);
and U28061 (N_28061,N_27604,N_27632);
nor U28062 (N_28062,N_27697,N_27729);
nand U28063 (N_28063,N_27592,N_27700);
nor U28064 (N_28064,N_27705,N_27841);
xnor U28065 (N_28065,N_27797,N_27511);
nand U28066 (N_28066,N_27808,N_27734);
xor U28067 (N_28067,N_27804,N_27596);
or U28068 (N_28068,N_27913,N_27626);
xor U28069 (N_28069,N_27865,N_27998);
and U28070 (N_28070,N_27882,N_27874);
nand U28071 (N_28071,N_27577,N_27925);
nand U28072 (N_28072,N_27739,N_27989);
or U28073 (N_28073,N_27712,N_27536);
nand U28074 (N_28074,N_27581,N_27845);
or U28075 (N_28075,N_27801,N_27798);
nand U28076 (N_28076,N_27770,N_27579);
xnor U28077 (N_28077,N_27523,N_27810);
or U28078 (N_28078,N_27727,N_27541);
xor U28079 (N_28079,N_27850,N_27677);
xnor U28080 (N_28080,N_27633,N_27964);
xnor U28081 (N_28081,N_27782,N_27946);
nand U28082 (N_28082,N_27659,N_27613);
nand U28083 (N_28083,N_27878,N_27811);
or U28084 (N_28084,N_27908,N_27921);
and U28085 (N_28085,N_27828,N_27566);
xor U28086 (N_28086,N_27985,N_27578);
xor U28087 (N_28087,N_27813,N_27627);
nor U28088 (N_28088,N_27786,N_27699);
nor U28089 (N_28089,N_27942,N_27963);
and U28090 (N_28090,N_27601,N_27827);
nor U28091 (N_28091,N_27525,N_27624);
xor U28092 (N_28092,N_27831,N_27852);
and U28093 (N_28093,N_27824,N_27936);
nor U28094 (N_28094,N_27540,N_27757);
or U28095 (N_28095,N_27686,N_27821);
xor U28096 (N_28096,N_27888,N_27635);
and U28097 (N_28097,N_27726,N_27649);
and U28098 (N_28098,N_27934,N_27599);
or U28099 (N_28099,N_27708,N_27872);
nor U28100 (N_28100,N_27982,N_27837);
or U28101 (N_28101,N_27990,N_27720);
xor U28102 (N_28102,N_27897,N_27655);
xnor U28103 (N_28103,N_27639,N_27950);
nand U28104 (N_28104,N_27539,N_27721);
xor U28105 (N_28105,N_27937,N_27749);
and U28106 (N_28106,N_27534,N_27570);
and U28107 (N_28107,N_27790,N_27843);
nor U28108 (N_28108,N_27519,N_27924);
or U28109 (N_28109,N_27887,N_27905);
xor U28110 (N_28110,N_27764,N_27669);
or U28111 (N_28111,N_27789,N_27614);
nand U28112 (N_28112,N_27694,N_27943);
nor U28113 (N_28113,N_27692,N_27826);
nor U28114 (N_28114,N_27835,N_27947);
nand U28115 (N_28115,N_27619,N_27598);
or U28116 (N_28116,N_27997,N_27567);
and U28117 (N_28117,N_27703,N_27752);
nor U28118 (N_28118,N_27645,N_27817);
nor U28119 (N_28119,N_27933,N_27538);
and U28120 (N_28120,N_27794,N_27862);
nand U28121 (N_28121,N_27513,N_27676);
xnor U28122 (N_28122,N_27688,N_27557);
nand U28123 (N_28123,N_27584,N_27890);
nand U28124 (N_28124,N_27725,N_27719);
nor U28125 (N_28125,N_27760,N_27939);
and U28126 (N_28126,N_27920,N_27917);
xor U28127 (N_28127,N_27906,N_27529);
nor U28128 (N_28128,N_27930,N_27551);
nor U28129 (N_28129,N_27959,N_27548);
and U28130 (N_28130,N_27892,N_27896);
and U28131 (N_28131,N_27818,N_27883);
xnor U28132 (N_28132,N_27758,N_27799);
nor U28133 (N_28133,N_27597,N_27546);
nor U28134 (N_28134,N_27588,N_27564);
or U28135 (N_28135,N_27663,N_27524);
and U28136 (N_28136,N_27518,N_27709);
xor U28137 (N_28137,N_27550,N_27754);
or U28138 (N_28138,N_27765,N_27916);
nand U28139 (N_28139,N_27504,N_27532);
nor U28140 (N_28140,N_27971,N_27978);
and U28141 (N_28141,N_27854,N_27761);
or U28142 (N_28142,N_27871,N_27796);
or U28143 (N_28143,N_27738,N_27731);
or U28144 (N_28144,N_27848,N_27644);
and U28145 (N_28145,N_27941,N_27753);
xor U28146 (N_28146,N_27922,N_27569);
xor U28147 (N_28147,N_27730,N_27612);
or U28148 (N_28148,N_27788,N_27535);
and U28149 (N_28149,N_27996,N_27628);
xnor U28150 (N_28150,N_27501,N_27960);
and U28151 (N_28151,N_27678,N_27762);
nor U28152 (N_28152,N_27970,N_27502);
or U28153 (N_28153,N_27656,N_27658);
nor U28154 (N_28154,N_27514,N_27728);
xor U28155 (N_28155,N_27981,N_27776);
nor U28156 (N_28156,N_27693,N_27737);
or U28157 (N_28157,N_27860,N_27999);
and U28158 (N_28158,N_27555,N_27814);
or U28159 (N_28159,N_27582,N_27580);
xnor U28160 (N_28160,N_27576,N_27522);
nor U28161 (N_28161,N_27834,N_27573);
and U28162 (N_28162,N_27544,N_27868);
xor U28163 (N_28163,N_27867,N_27976);
xnor U28164 (N_28164,N_27742,N_27968);
or U28165 (N_28165,N_27553,N_27863);
xor U28166 (N_28166,N_27866,N_27812);
nand U28167 (N_28167,N_27747,N_27915);
xnor U28168 (N_28168,N_27668,N_27775);
nand U28169 (N_28169,N_27876,N_27620);
and U28170 (N_28170,N_27965,N_27926);
or U28171 (N_28171,N_27750,N_27779);
or U28172 (N_28172,N_27507,N_27512);
xor U28173 (N_28173,N_27886,N_27651);
nor U28174 (N_28174,N_27816,N_27972);
or U28175 (N_28175,N_27615,N_27660);
nand U28176 (N_28176,N_27954,N_27682);
or U28177 (N_28177,N_27723,N_27606);
xor U28178 (N_28178,N_27643,N_27988);
nor U28179 (N_28179,N_27973,N_27568);
nand U28180 (N_28180,N_27505,N_27987);
nand U28181 (N_28181,N_27759,N_27743);
nor U28182 (N_28182,N_27957,N_27927);
or U28183 (N_28183,N_27714,N_27986);
nand U28184 (N_28184,N_27702,N_27745);
or U28185 (N_28185,N_27983,N_27690);
nand U28186 (N_28186,N_27822,N_27967);
or U28187 (N_28187,N_27956,N_27829);
nor U28188 (N_28188,N_27661,N_27704);
nand U28189 (N_28189,N_27547,N_27642);
xor U28190 (N_28190,N_27751,N_27909);
xnor U28191 (N_28191,N_27771,N_27901);
nand U28192 (N_28192,N_27698,N_27853);
nor U28193 (N_28193,N_27631,N_27558);
nor U28194 (N_28194,N_27610,N_27945);
and U28195 (N_28195,N_27586,N_27953);
nor U28196 (N_28196,N_27769,N_27864);
nand U28197 (N_28197,N_27975,N_27795);
and U28198 (N_28198,N_27707,N_27949);
nor U28199 (N_28199,N_27715,N_27820);
or U28200 (N_28200,N_27825,N_27509);
nand U28201 (N_28201,N_27781,N_27706);
xor U28202 (N_28202,N_27919,N_27792);
and U28203 (N_28203,N_27683,N_27912);
or U28204 (N_28204,N_27616,N_27508);
and U28205 (N_28205,N_27911,N_27542);
nor U28206 (N_28206,N_27563,N_27979);
xnor U28207 (N_28207,N_27717,N_27885);
and U28208 (N_28208,N_27625,N_27842);
or U28209 (N_28209,N_27891,N_27527);
or U28210 (N_28210,N_27880,N_27774);
nor U28211 (N_28211,N_27641,N_27784);
xnor U28212 (N_28212,N_27607,N_27560);
or U28213 (N_28213,N_27875,N_27800);
nand U28214 (N_28214,N_27857,N_27907);
or U28215 (N_28215,N_27948,N_27793);
or U28216 (N_28216,N_27740,N_27766);
nand U28217 (N_28217,N_27733,N_27914);
nand U28218 (N_28218,N_27545,N_27572);
nand U28219 (N_28219,N_27791,N_27940);
xnor U28220 (N_28220,N_27736,N_27903);
and U28221 (N_28221,N_27846,N_27521);
nor U28222 (N_28222,N_27680,N_27840);
or U28223 (N_28223,N_27583,N_27565);
and U28224 (N_28224,N_27938,N_27873);
nand U28225 (N_28225,N_27650,N_27994);
nor U28226 (N_28226,N_27962,N_27877);
nand U28227 (N_28227,N_27756,N_27778);
nand U28228 (N_28228,N_27595,N_27695);
nand U28229 (N_28229,N_27893,N_27741);
nor U28230 (N_28230,N_27647,N_27590);
nor U28231 (N_28231,N_27910,N_27611);
nand U28232 (N_28232,N_27585,N_27785);
and U28233 (N_28233,N_27591,N_27847);
or U28234 (N_28234,N_27561,N_27554);
and U28235 (N_28235,N_27562,N_27657);
xor U28236 (N_28236,N_27993,N_27773);
or U28237 (N_28237,N_27679,N_27673);
nand U28238 (N_28238,N_27767,N_27675);
nor U28239 (N_28239,N_27895,N_27696);
nor U28240 (N_28240,N_27879,N_27830);
xnor U28241 (N_28241,N_27806,N_27807);
and U28242 (N_28242,N_27587,N_27881);
nor U28243 (N_28243,N_27977,N_27691);
nor U28244 (N_28244,N_27918,N_27630);
or U28245 (N_28245,N_27932,N_27851);
nand U28246 (N_28246,N_27952,N_27735);
or U28247 (N_28247,N_27533,N_27823);
or U28248 (N_28248,N_27787,N_27724);
or U28249 (N_28249,N_27638,N_27510);
nand U28250 (N_28250,N_27566,N_27810);
xnor U28251 (N_28251,N_27670,N_27759);
xnor U28252 (N_28252,N_27879,N_27816);
nor U28253 (N_28253,N_27580,N_27739);
xor U28254 (N_28254,N_27922,N_27603);
nand U28255 (N_28255,N_27902,N_27697);
nand U28256 (N_28256,N_27845,N_27824);
nand U28257 (N_28257,N_27871,N_27670);
nand U28258 (N_28258,N_27746,N_27715);
nand U28259 (N_28259,N_27985,N_27956);
nand U28260 (N_28260,N_27668,N_27621);
nand U28261 (N_28261,N_27625,N_27525);
or U28262 (N_28262,N_27758,N_27511);
and U28263 (N_28263,N_27770,N_27958);
nor U28264 (N_28264,N_27815,N_27902);
xnor U28265 (N_28265,N_27756,N_27636);
or U28266 (N_28266,N_27503,N_27533);
xor U28267 (N_28267,N_27697,N_27654);
or U28268 (N_28268,N_27996,N_27913);
xnor U28269 (N_28269,N_27954,N_27980);
or U28270 (N_28270,N_27750,N_27625);
xnor U28271 (N_28271,N_27616,N_27806);
or U28272 (N_28272,N_27765,N_27728);
nor U28273 (N_28273,N_27557,N_27555);
nand U28274 (N_28274,N_27702,N_27985);
or U28275 (N_28275,N_27770,N_27843);
and U28276 (N_28276,N_27537,N_27524);
nand U28277 (N_28277,N_27939,N_27571);
or U28278 (N_28278,N_27698,N_27891);
xnor U28279 (N_28279,N_27818,N_27814);
or U28280 (N_28280,N_27660,N_27624);
nand U28281 (N_28281,N_27586,N_27641);
nand U28282 (N_28282,N_27514,N_27661);
xor U28283 (N_28283,N_27977,N_27738);
nand U28284 (N_28284,N_27964,N_27831);
and U28285 (N_28285,N_27631,N_27822);
nor U28286 (N_28286,N_27890,N_27745);
xor U28287 (N_28287,N_27616,N_27529);
nand U28288 (N_28288,N_27592,N_27670);
nor U28289 (N_28289,N_27649,N_27962);
nor U28290 (N_28290,N_27788,N_27785);
nor U28291 (N_28291,N_27558,N_27872);
and U28292 (N_28292,N_27861,N_27668);
xor U28293 (N_28293,N_27890,N_27606);
xor U28294 (N_28294,N_27958,N_27642);
and U28295 (N_28295,N_27786,N_27590);
nand U28296 (N_28296,N_27897,N_27690);
and U28297 (N_28297,N_27892,N_27768);
xnor U28298 (N_28298,N_27845,N_27571);
nand U28299 (N_28299,N_27960,N_27524);
nor U28300 (N_28300,N_27514,N_27533);
nand U28301 (N_28301,N_27797,N_27686);
or U28302 (N_28302,N_27568,N_27525);
or U28303 (N_28303,N_27860,N_27785);
nor U28304 (N_28304,N_27687,N_27894);
or U28305 (N_28305,N_27619,N_27697);
nand U28306 (N_28306,N_27921,N_27545);
or U28307 (N_28307,N_27820,N_27792);
or U28308 (N_28308,N_27607,N_27561);
or U28309 (N_28309,N_27675,N_27968);
nand U28310 (N_28310,N_27696,N_27774);
nand U28311 (N_28311,N_27995,N_27761);
xor U28312 (N_28312,N_27614,N_27869);
nor U28313 (N_28313,N_27623,N_27509);
and U28314 (N_28314,N_27620,N_27639);
nor U28315 (N_28315,N_27646,N_27654);
nand U28316 (N_28316,N_27855,N_27695);
xor U28317 (N_28317,N_27555,N_27744);
nor U28318 (N_28318,N_27774,N_27751);
nand U28319 (N_28319,N_27567,N_27939);
xnor U28320 (N_28320,N_27644,N_27638);
and U28321 (N_28321,N_27812,N_27690);
or U28322 (N_28322,N_27671,N_27903);
xor U28323 (N_28323,N_27954,N_27683);
nor U28324 (N_28324,N_27600,N_27699);
or U28325 (N_28325,N_27869,N_27733);
or U28326 (N_28326,N_27626,N_27638);
nand U28327 (N_28327,N_27853,N_27607);
nor U28328 (N_28328,N_27922,N_27759);
nand U28329 (N_28329,N_27517,N_27676);
or U28330 (N_28330,N_27738,N_27859);
xor U28331 (N_28331,N_27563,N_27746);
and U28332 (N_28332,N_27780,N_27600);
and U28333 (N_28333,N_27742,N_27964);
nor U28334 (N_28334,N_27973,N_27761);
xor U28335 (N_28335,N_27888,N_27803);
nor U28336 (N_28336,N_27877,N_27722);
xor U28337 (N_28337,N_27955,N_27563);
and U28338 (N_28338,N_27956,N_27899);
nand U28339 (N_28339,N_27874,N_27587);
xnor U28340 (N_28340,N_27683,N_27612);
and U28341 (N_28341,N_27856,N_27837);
xnor U28342 (N_28342,N_27616,N_27507);
xnor U28343 (N_28343,N_27573,N_27594);
and U28344 (N_28344,N_27526,N_27624);
and U28345 (N_28345,N_27850,N_27881);
xor U28346 (N_28346,N_27650,N_27641);
or U28347 (N_28347,N_27690,N_27628);
or U28348 (N_28348,N_27781,N_27786);
or U28349 (N_28349,N_27640,N_27539);
nand U28350 (N_28350,N_27800,N_27872);
xnor U28351 (N_28351,N_27875,N_27851);
and U28352 (N_28352,N_27664,N_27652);
nand U28353 (N_28353,N_27588,N_27835);
xor U28354 (N_28354,N_27716,N_27987);
and U28355 (N_28355,N_27853,N_27703);
and U28356 (N_28356,N_27892,N_27675);
nand U28357 (N_28357,N_27908,N_27713);
xnor U28358 (N_28358,N_27720,N_27721);
xor U28359 (N_28359,N_27701,N_27759);
nor U28360 (N_28360,N_27928,N_27860);
nand U28361 (N_28361,N_27711,N_27717);
nor U28362 (N_28362,N_27802,N_27702);
and U28363 (N_28363,N_27715,N_27947);
and U28364 (N_28364,N_27569,N_27829);
xnor U28365 (N_28365,N_27822,N_27509);
or U28366 (N_28366,N_27738,N_27526);
nor U28367 (N_28367,N_27671,N_27573);
xor U28368 (N_28368,N_27786,N_27762);
or U28369 (N_28369,N_27893,N_27680);
xor U28370 (N_28370,N_27947,N_27772);
nor U28371 (N_28371,N_27508,N_27762);
nand U28372 (N_28372,N_27527,N_27828);
nand U28373 (N_28373,N_27910,N_27573);
xor U28374 (N_28374,N_27671,N_27668);
and U28375 (N_28375,N_27783,N_27903);
xor U28376 (N_28376,N_27951,N_27564);
nor U28377 (N_28377,N_27989,N_27539);
xnor U28378 (N_28378,N_27944,N_27522);
or U28379 (N_28379,N_27957,N_27573);
xnor U28380 (N_28380,N_27581,N_27972);
nor U28381 (N_28381,N_27575,N_27577);
xnor U28382 (N_28382,N_27563,N_27977);
xnor U28383 (N_28383,N_27530,N_27520);
nand U28384 (N_28384,N_27938,N_27635);
and U28385 (N_28385,N_27634,N_27531);
nand U28386 (N_28386,N_27603,N_27719);
xnor U28387 (N_28387,N_27724,N_27758);
nand U28388 (N_28388,N_27667,N_27760);
or U28389 (N_28389,N_27540,N_27809);
xnor U28390 (N_28390,N_27512,N_27611);
nand U28391 (N_28391,N_27665,N_27874);
xnor U28392 (N_28392,N_27921,N_27852);
nand U28393 (N_28393,N_27792,N_27775);
nand U28394 (N_28394,N_27918,N_27539);
and U28395 (N_28395,N_27569,N_27697);
and U28396 (N_28396,N_27727,N_27971);
nand U28397 (N_28397,N_27882,N_27805);
nor U28398 (N_28398,N_27982,N_27838);
and U28399 (N_28399,N_27582,N_27922);
or U28400 (N_28400,N_27835,N_27707);
and U28401 (N_28401,N_27704,N_27883);
and U28402 (N_28402,N_27648,N_27568);
nand U28403 (N_28403,N_27772,N_27851);
or U28404 (N_28404,N_27594,N_27944);
xnor U28405 (N_28405,N_27926,N_27684);
xor U28406 (N_28406,N_27510,N_27551);
or U28407 (N_28407,N_27792,N_27666);
and U28408 (N_28408,N_27817,N_27960);
or U28409 (N_28409,N_27596,N_27717);
or U28410 (N_28410,N_27840,N_27844);
nor U28411 (N_28411,N_27763,N_27990);
xnor U28412 (N_28412,N_27694,N_27704);
or U28413 (N_28413,N_27830,N_27809);
or U28414 (N_28414,N_27974,N_27956);
and U28415 (N_28415,N_27803,N_27530);
nand U28416 (N_28416,N_27526,N_27651);
nand U28417 (N_28417,N_27569,N_27605);
and U28418 (N_28418,N_27585,N_27927);
nand U28419 (N_28419,N_27572,N_27793);
xnor U28420 (N_28420,N_27945,N_27541);
or U28421 (N_28421,N_27956,N_27834);
and U28422 (N_28422,N_27584,N_27515);
or U28423 (N_28423,N_27764,N_27958);
nor U28424 (N_28424,N_27823,N_27662);
or U28425 (N_28425,N_27915,N_27601);
and U28426 (N_28426,N_27857,N_27939);
nor U28427 (N_28427,N_27924,N_27651);
and U28428 (N_28428,N_27630,N_27518);
and U28429 (N_28429,N_27625,N_27686);
xnor U28430 (N_28430,N_27730,N_27630);
nand U28431 (N_28431,N_27721,N_27984);
xnor U28432 (N_28432,N_27822,N_27897);
nor U28433 (N_28433,N_27602,N_27503);
nor U28434 (N_28434,N_27593,N_27727);
and U28435 (N_28435,N_27554,N_27999);
nor U28436 (N_28436,N_27548,N_27982);
and U28437 (N_28437,N_27864,N_27890);
or U28438 (N_28438,N_27644,N_27631);
xnor U28439 (N_28439,N_27675,N_27992);
and U28440 (N_28440,N_27500,N_27568);
nand U28441 (N_28441,N_27692,N_27725);
or U28442 (N_28442,N_27604,N_27800);
or U28443 (N_28443,N_27958,N_27582);
xor U28444 (N_28444,N_27891,N_27597);
and U28445 (N_28445,N_27574,N_27637);
or U28446 (N_28446,N_27660,N_27644);
or U28447 (N_28447,N_27737,N_27555);
xor U28448 (N_28448,N_27539,N_27507);
nor U28449 (N_28449,N_27589,N_27841);
nand U28450 (N_28450,N_27886,N_27715);
xor U28451 (N_28451,N_27707,N_27824);
nand U28452 (N_28452,N_27991,N_27665);
xnor U28453 (N_28453,N_27975,N_27783);
and U28454 (N_28454,N_27688,N_27924);
and U28455 (N_28455,N_27932,N_27900);
or U28456 (N_28456,N_27796,N_27544);
nand U28457 (N_28457,N_27915,N_27596);
nand U28458 (N_28458,N_27765,N_27773);
nor U28459 (N_28459,N_27659,N_27987);
and U28460 (N_28460,N_27704,N_27884);
nand U28461 (N_28461,N_27829,N_27743);
xor U28462 (N_28462,N_27805,N_27655);
and U28463 (N_28463,N_27927,N_27654);
or U28464 (N_28464,N_27812,N_27659);
nand U28465 (N_28465,N_27561,N_27956);
and U28466 (N_28466,N_27716,N_27664);
and U28467 (N_28467,N_27637,N_27569);
and U28468 (N_28468,N_27665,N_27633);
or U28469 (N_28469,N_27949,N_27910);
and U28470 (N_28470,N_27993,N_27546);
or U28471 (N_28471,N_27517,N_27685);
nor U28472 (N_28472,N_27540,N_27771);
xor U28473 (N_28473,N_27650,N_27804);
or U28474 (N_28474,N_27749,N_27596);
nor U28475 (N_28475,N_27522,N_27530);
xor U28476 (N_28476,N_27727,N_27780);
and U28477 (N_28477,N_27694,N_27899);
nand U28478 (N_28478,N_27506,N_27640);
or U28479 (N_28479,N_27891,N_27801);
nand U28480 (N_28480,N_27679,N_27530);
and U28481 (N_28481,N_27659,N_27970);
or U28482 (N_28482,N_27528,N_27963);
nor U28483 (N_28483,N_27788,N_27971);
nor U28484 (N_28484,N_27644,N_27742);
or U28485 (N_28485,N_27680,N_27612);
xnor U28486 (N_28486,N_27514,N_27645);
or U28487 (N_28487,N_27848,N_27705);
nor U28488 (N_28488,N_27809,N_27835);
or U28489 (N_28489,N_27505,N_27790);
or U28490 (N_28490,N_27896,N_27977);
and U28491 (N_28491,N_27765,N_27810);
xnor U28492 (N_28492,N_27605,N_27792);
xnor U28493 (N_28493,N_27774,N_27811);
nor U28494 (N_28494,N_27887,N_27948);
nand U28495 (N_28495,N_27685,N_27536);
nand U28496 (N_28496,N_27631,N_27586);
xor U28497 (N_28497,N_27951,N_27847);
xnor U28498 (N_28498,N_27899,N_27622);
and U28499 (N_28499,N_27969,N_27822);
nor U28500 (N_28500,N_28113,N_28232);
xor U28501 (N_28501,N_28083,N_28447);
xor U28502 (N_28502,N_28290,N_28278);
and U28503 (N_28503,N_28398,N_28238);
xnor U28504 (N_28504,N_28120,N_28117);
nor U28505 (N_28505,N_28243,N_28163);
nor U28506 (N_28506,N_28018,N_28189);
nor U28507 (N_28507,N_28431,N_28153);
and U28508 (N_28508,N_28204,N_28383);
or U28509 (N_28509,N_28344,N_28468);
or U28510 (N_28510,N_28402,N_28212);
xnor U28511 (N_28511,N_28176,N_28020);
and U28512 (N_28512,N_28361,N_28051);
or U28513 (N_28513,N_28213,N_28003);
xor U28514 (N_28514,N_28267,N_28174);
or U28515 (N_28515,N_28100,N_28218);
xor U28516 (N_28516,N_28325,N_28224);
or U28517 (N_28517,N_28064,N_28346);
nand U28518 (N_28518,N_28006,N_28122);
nand U28519 (N_28519,N_28036,N_28138);
or U28520 (N_28520,N_28130,N_28458);
nor U28521 (N_28521,N_28126,N_28420);
nand U28522 (N_28522,N_28237,N_28317);
nor U28523 (N_28523,N_28414,N_28401);
nor U28524 (N_28524,N_28305,N_28332);
or U28525 (N_28525,N_28418,N_28114);
or U28526 (N_28526,N_28086,N_28348);
or U28527 (N_28527,N_28360,N_28050);
nand U28528 (N_28528,N_28201,N_28143);
nor U28529 (N_28529,N_28301,N_28460);
and U28530 (N_28530,N_28443,N_28221);
and U28531 (N_28531,N_28375,N_28230);
nor U28532 (N_28532,N_28257,N_28466);
xor U28533 (N_28533,N_28250,N_28014);
and U28534 (N_28534,N_28098,N_28262);
nor U28535 (N_28535,N_28068,N_28388);
and U28536 (N_28536,N_28087,N_28004);
or U28537 (N_28537,N_28002,N_28371);
xor U28538 (N_28538,N_28437,N_28469);
or U28539 (N_28539,N_28181,N_28067);
or U28540 (N_28540,N_28258,N_28376);
and U28541 (N_28541,N_28467,N_28178);
nand U28542 (N_28542,N_28052,N_28075);
and U28543 (N_28543,N_28433,N_28286);
nand U28544 (N_28544,N_28477,N_28307);
nand U28545 (N_28545,N_28152,N_28311);
xnor U28546 (N_28546,N_28266,N_28043);
nor U28547 (N_28547,N_28353,N_28352);
and U28548 (N_28548,N_28233,N_28480);
or U28549 (N_28549,N_28451,N_28473);
nor U28550 (N_28550,N_28440,N_28300);
or U28551 (N_28551,N_28277,N_28161);
xnor U28552 (N_28552,N_28154,N_28298);
xnor U28553 (N_28553,N_28369,N_28125);
nor U28554 (N_28554,N_28013,N_28039);
xor U28555 (N_28555,N_28455,N_28231);
nor U28556 (N_28556,N_28435,N_28166);
xnor U28557 (N_28557,N_28157,N_28405);
nand U28558 (N_28558,N_28139,N_28072);
or U28559 (N_28559,N_28172,N_28256);
nor U28560 (N_28560,N_28488,N_28448);
xor U28561 (N_28561,N_28141,N_28194);
and U28562 (N_28562,N_28270,N_28297);
nor U28563 (N_28563,N_28310,N_28076);
and U28564 (N_28564,N_28185,N_28494);
xnor U28565 (N_28565,N_28214,N_28073);
or U28566 (N_28566,N_28019,N_28283);
xor U28567 (N_28567,N_28032,N_28343);
nor U28568 (N_28568,N_28198,N_28093);
xnor U28569 (N_28569,N_28481,N_28220);
or U28570 (N_28570,N_28490,N_28391);
nand U28571 (N_28571,N_28400,N_28392);
nor U28572 (N_28572,N_28432,N_28292);
nor U28573 (N_28573,N_28321,N_28354);
xor U28574 (N_28574,N_28336,N_28132);
or U28575 (N_28575,N_28021,N_28428);
nor U28576 (N_28576,N_28454,N_28226);
and U28577 (N_28577,N_28062,N_28190);
and U28578 (N_28578,N_28159,N_28492);
and U28579 (N_28579,N_28063,N_28082);
and U28580 (N_28580,N_28441,N_28287);
nor U28581 (N_28581,N_28121,N_28497);
nand U28582 (N_28582,N_28341,N_28498);
or U28583 (N_28583,N_28165,N_28274);
xnor U28584 (N_28584,N_28302,N_28229);
nor U28585 (N_28585,N_28394,N_28284);
or U28586 (N_28586,N_28055,N_28412);
xor U28587 (N_28587,N_28109,N_28110);
xor U28588 (N_28588,N_28404,N_28253);
xnor U28589 (N_28589,N_28041,N_28060);
and U28590 (N_28590,N_28396,N_28099);
nand U28591 (N_28591,N_28379,N_28385);
xor U28592 (N_28592,N_28340,N_28149);
xnor U28593 (N_28593,N_28471,N_28035);
nor U28594 (N_28594,N_28276,N_28180);
or U28595 (N_28595,N_28367,N_28085);
nand U28596 (N_28596,N_28235,N_28319);
or U28597 (N_28597,N_28119,N_28495);
xor U28598 (N_28598,N_28182,N_28475);
or U28599 (N_28599,N_28254,N_28049);
nand U28600 (N_28600,N_28249,N_28217);
or U28601 (N_28601,N_28461,N_28155);
or U28602 (N_28602,N_28282,N_28069);
and U28603 (N_28603,N_28417,N_28476);
nand U28604 (N_28604,N_28273,N_28025);
nor U28605 (N_28605,N_28294,N_28046);
and U28606 (N_28606,N_28016,N_28304);
xnor U28607 (N_28607,N_28101,N_28007);
nor U28608 (N_28608,N_28413,N_28255);
nor U28609 (N_28609,N_28167,N_28309);
and U28610 (N_28610,N_28116,N_28291);
xnor U28611 (N_28611,N_28091,N_28211);
or U28612 (N_28612,N_28345,N_28065);
nor U28613 (N_28613,N_28380,N_28179);
or U28614 (N_28614,N_28088,N_28489);
or U28615 (N_28615,N_28188,N_28351);
or U28616 (N_28616,N_28429,N_28406);
xnor U28617 (N_28617,N_28295,N_28339);
or U28618 (N_28618,N_28334,N_28223);
xnor U28619 (N_28619,N_28191,N_28140);
xnor U28620 (N_28620,N_28128,N_28026);
nor U28621 (N_28621,N_28430,N_28081);
xor U28622 (N_28622,N_28245,N_28260);
xor U28623 (N_28623,N_28293,N_28370);
and U28624 (N_28624,N_28170,N_28395);
or U28625 (N_28625,N_28424,N_28355);
or U28626 (N_28626,N_28029,N_28248);
xor U28627 (N_28627,N_28022,N_28337);
xor U28628 (N_28628,N_28323,N_28023);
xor U28629 (N_28629,N_28202,N_28357);
xnor U28630 (N_28630,N_28330,N_28184);
xor U28631 (N_28631,N_28078,N_28192);
nand U28632 (N_28632,N_28387,N_28107);
and U28633 (N_28633,N_28071,N_28227);
nand U28634 (N_28634,N_28005,N_28015);
xor U28635 (N_28635,N_28197,N_28483);
and U28636 (N_28636,N_28027,N_28397);
xor U28637 (N_28637,N_28491,N_28416);
or U28638 (N_28638,N_28215,N_28133);
nand U28639 (N_28639,N_28054,N_28486);
xnor U28640 (N_28640,N_28382,N_28123);
nor U28641 (N_28641,N_28144,N_28464);
and U28642 (N_28642,N_28279,N_28421);
nor U28643 (N_28643,N_28059,N_28203);
nand U28644 (N_28644,N_28285,N_28306);
and U28645 (N_28645,N_28342,N_28038);
xor U28646 (N_28646,N_28472,N_28415);
or U28647 (N_28647,N_28028,N_28303);
xor U28648 (N_28648,N_28208,N_28164);
nand U28649 (N_28649,N_28111,N_28449);
xor U28650 (N_28650,N_28024,N_28158);
nand U28651 (N_28651,N_28427,N_28146);
xor U28652 (N_28652,N_28240,N_28496);
xor U28653 (N_28653,N_28269,N_28320);
nor U28654 (N_28654,N_28044,N_28446);
xor U28655 (N_28655,N_28268,N_28225);
nor U28656 (N_28656,N_28136,N_28324);
xor U28657 (N_28657,N_28066,N_28175);
nand U28658 (N_28658,N_28493,N_28008);
nand U28659 (N_28659,N_28077,N_28372);
nor U28660 (N_28660,N_28030,N_28009);
or U28661 (N_28661,N_28210,N_28445);
or U28662 (N_28662,N_28183,N_28090);
nor U28663 (N_28663,N_28338,N_28058);
nand U28664 (N_28664,N_28187,N_28034);
nor U28665 (N_28665,N_28012,N_28042);
and U28666 (N_28666,N_28470,N_28499);
nand U28667 (N_28667,N_28033,N_28048);
or U28668 (N_28668,N_28209,N_28299);
nand U28669 (N_28669,N_28381,N_28142);
and U28670 (N_28670,N_28131,N_28053);
nand U28671 (N_28671,N_28289,N_28263);
and U28672 (N_28672,N_28423,N_28247);
xor U28673 (N_28673,N_28364,N_28102);
and U28674 (N_28674,N_28373,N_28017);
or U28675 (N_28675,N_28127,N_28228);
xnor U28676 (N_28676,N_28104,N_28156);
and U28677 (N_28677,N_28135,N_28314);
xnor U28678 (N_28678,N_28061,N_28084);
or U28679 (N_28679,N_28322,N_28374);
or U28680 (N_28680,N_28239,N_28259);
nor U28681 (N_28681,N_28089,N_28459);
nand U28682 (N_28682,N_28074,N_28331);
nand U28683 (N_28683,N_28296,N_28108);
and U28684 (N_28684,N_28205,N_28150);
and U28685 (N_28685,N_28316,N_28200);
or U28686 (N_28686,N_28329,N_28327);
xor U28687 (N_28687,N_28236,N_28453);
nand U28688 (N_28688,N_28092,N_28080);
xnor U28689 (N_28689,N_28452,N_28097);
nor U28690 (N_28690,N_28160,N_28162);
nand U28691 (N_28691,N_28251,N_28426);
and U28692 (N_28692,N_28425,N_28112);
nor U28693 (N_28693,N_28271,N_28368);
or U28694 (N_28694,N_28487,N_28362);
xor U28695 (N_28695,N_28095,N_28407);
nand U28696 (N_28696,N_28047,N_28206);
xnor U28697 (N_28697,N_28312,N_28106);
nor U28698 (N_28698,N_28328,N_28168);
and U28699 (N_28699,N_28411,N_28403);
xnor U28700 (N_28700,N_28195,N_28103);
and U28701 (N_28701,N_28275,N_28171);
xor U28702 (N_28702,N_28386,N_28000);
and U28703 (N_28703,N_28031,N_28129);
xor U28704 (N_28704,N_28105,N_28118);
and U28705 (N_28705,N_28484,N_28390);
and U28706 (N_28706,N_28399,N_28335);
and U28707 (N_28707,N_28216,N_28315);
nand U28708 (N_28708,N_28242,N_28422);
and U28709 (N_28709,N_28186,N_28389);
nand U28710 (N_28710,N_28457,N_28442);
xor U28711 (N_28711,N_28363,N_28264);
and U28712 (N_28712,N_28465,N_28384);
or U28713 (N_28713,N_28419,N_28359);
and U28714 (N_28714,N_28261,N_28057);
or U28715 (N_28715,N_28393,N_28479);
or U28716 (N_28716,N_28350,N_28288);
nand U28717 (N_28717,N_28196,N_28151);
nor U28718 (N_28718,N_28349,N_28450);
and U28719 (N_28719,N_28265,N_28070);
nor U28720 (N_28720,N_28333,N_28079);
xor U28721 (N_28721,N_28365,N_28193);
xor U28722 (N_28722,N_28115,N_28246);
and U28723 (N_28723,N_28438,N_28439);
and U28724 (N_28724,N_28037,N_28409);
nor U28725 (N_28725,N_28096,N_28222);
nand U28726 (N_28726,N_28326,N_28147);
or U28727 (N_28727,N_28356,N_28358);
nand U28728 (N_28728,N_28408,N_28478);
nor U28729 (N_28729,N_28281,N_28347);
xnor U28730 (N_28730,N_28169,N_28482);
nor U28731 (N_28731,N_28207,N_28280);
and U28732 (N_28732,N_28199,N_28366);
nor U28733 (N_28733,N_28177,N_28134);
nand U28734 (N_28734,N_28462,N_28241);
nand U28735 (N_28735,N_28137,N_28094);
xnor U28736 (N_28736,N_28124,N_28045);
nor U28737 (N_28737,N_28377,N_28463);
nor U28738 (N_28738,N_28244,N_28308);
or U28739 (N_28739,N_28056,N_28410);
xor U28740 (N_28740,N_28485,N_28010);
and U28741 (N_28741,N_28434,N_28148);
and U28742 (N_28742,N_28272,N_28040);
xor U28743 (N_28743,N_28252,N_28011);
nor U28744 (N_28744,N_28474,N_28318);
or U28745 (N_28745,N_28219,N_28145);
nand U28746 (N_28746,N_28001,N_28456);
nor U28747 (N_28747,N_28436,N_28378);
nor U28748 (N_28748,N_28313,N_28234);
xnor U28749 (N_28749,N_28444,N_28173);
nand U28750 (N_28750,N_28320,N_28219);
or U28751 (N_28751,N_28122,N_28048);
nor U28752 (N_28752,N_28253,N_28230);
nor U28753 (N_28753,N_28428,N_28189);
nor U28754 (N_28754,N_28255,N_28481);
xnor U28755 (N_28755,N_28098,N_28182);
xnor U28756 (N_28756,N_28096,N_28074);
nand U28757 (N_28757,N_28140,N_28242);
and U28758 (N_28758,N_28465,N_28438);
nand U28759 (N_28759,N_28300,N_28261);
nor U28760 (N_28760,N_28404,N_28403);
xnor U28761 (N_28761,N_28381,N_28451);
or U28762 (N_28762,N_28490,N_28321);
and U28763 (N_28763,N_28069,N_28072);
and U28764 (N_28764,N_28427,N_28063);
and U28765 (N_28765,N_28064,N_28215);
or U28766 (N_28766,N_28132,N_28166);
nor U28767 (N_28767,N_28105,N_28363);
or U28768 (N_28768,N_28216,N_28497);
nand U28769 (N_28769,N_28310,N_28347);
nand U28770 (N_28770,N_28418,N_28400);
nand U28771 (N_28771,N_28190,N_28427);
or U28772 (N_28772,N_28302,N_28478);
and U28773 (N_28773,N_28113,N_28275);
xnor U28774 (N_28774,N_28035,N_28353);
or U28775 (N_28775,N_28480,N_28001);
nand U28776 (N_28776,N_28245,N_28486);
or U28777 (N_28777,N_28256,N_28136);
nand U28778 (N_28778,N_28117,N_28188);
or U28779 (N_28779,N_28297,N_28104);
nor U28780 (N_28780,N_28379,N_28476);
or U28781 (N_28781,N_28064,N_28046);
nand U28782 (N_28782,N_28241,N_28249);
nand U28783 (N_28783,N_28489,N_28211);
xnor U28784 (N_28784,N_28058,N_28377);
nor U28785 (N_28785,N_28305,N_28207);
xnor U28786 (N_28786,N_28101,N_28100);
nor U28787 (N_28787,N_28451,N_28354);
or U28788 (N_28788,N_28499,N_28082);
or U28789 (N_28789,N_28349,N_28044);
nor U28790 (N_28790,N_28112,N_28041);
nand U28791 (N_28791,N_28463,N_28330);
and U28792 (N_28792,N_28205,N_28211);
and U28793 (N_28793,N_28043,N_28229);
xnor U28794 (N_28794,N_28282,N_28393);
nand U28795 (N_28795,N_28412,N_28101);
nor U28796 (N_28796,N_28493,N_28044);
and U28797 (N_28797,N_28313,N_28283);
xor U28798 (N_28798,N_28459,N_28033);
xor U28799 (N_28799,N_28396,N_28389);
or U28800 (N_28800,N_28123,N_28255);
nand U28801 (N_28801,N_28341,N_28412);
nor U28802 (N_28802,N_28401,N_28266);
or U28803 (N_28803,N_28078,N_28154);
and U28804 (N_28804,N_28078,N_28406);
nand U28805 (N_28805,N_28006,N_28180);
nand U28806 (N_28806,N_28210,N_28039);
nand U28807 (N_28807,N_28424,N_28359);
nand U28808 (N_28808,N_28279,N_28484);
or U28809 (N_28809,N_28400,N_28187);
nand U28810 (N_28810,N_28350,N_28443);
and U28811 (N_28811,N_28208,N_28484);
or U28812 (N_28812,N_28436,N_28179);
nor U28813 (N_28813,N_28023,N_28178);
nand U28814 (N_28814,N_28356,N_28102);
and U28815 (N_28815,N_28073,N_28202);
or U28816 (N_28816,N_28427,N_28143);
and U28817 (N_28817,N_28329,N_28493);
or U28818 (N_28818,N_28362,N_28148);
nor U28819 (N_28819,N_28367,N_28011);
and U28820 (N_28820,N_28358,N_28414);
and U28821 (N_28821,N_28444,N_28375);
nand U28822 (N_28822,N_28156,N_28494);
nor U28823 (N_28823,N_28002,N_28171);
nor U28824 (N_28824,N_28134,N_28366);
or U28825 (N_28825,N_28255,N_28212);
nand U28826 (N_28826,N_28287,N_28325);
nand U28827 (N_28827,N_28045,N_28240);
or U28828 (N_28828,N_28300,N_28194);
nand U28829 (N_28829,N_28005,N_28207);
nand U28830 (N_28830,N_28360,N_28407);
xor U28831 (N_28831,N_28345,N_28360);
and U28832 (N_28832,N_28285,N_28288);
nor U28833 (N_28833,N_28390,N_28121);
and U28834 (N_28834,N_28219,N_28364);
and U28835 (N_28835,N_28142,N_28001);
nand U28836 (N_28836,N_28086,N_28214);
or U28837 (N_28837,N_28412,N_28267);
and U28838 (N_28838,N_28349,N_28471);
nor U28839 (N_28839,N_28486,N_28161);
nor U28840 (N_28840,N_28188,N_28029);
nand U28841 (N_28841,N_28417,N_28047);
nor U28842 (N_28842,N_28291,N_28006);
nand U28843 (N_28843,N_28366,N_28176);
xnor U28844 (N_28844,N_28329,N_28019);
or U28845 (N_28845,N_28476,N_28040);
nand U28846 (N_28846,N_28032,N_28198);
and U28847 (N_28847,N_28325,N_28467);
or U28848 (N_28848,N_28236,N_28085);
nand U28849 (N_28849,N_28452,N_28216);
and U28850 (N_28850,N_28229,N_28196);
and U28851 (N_28851,N_28324,N_28496);
nor U28852 (N_28852,N_28158,N_28377);
or U28853 (N_28853,N_28075,N_28348);
nor U28854 (N_28854,N_28045,N_28343);
or U28855 (N_28855,N_28450,N_28401);
or U28856 (N_28856,N_28136,N_28037);
and U28857 (N_28857,N_28495,N_28108);
xnor U28858 (N_28858,N_28071,N_28088);
or U28859 (N_28859,N_28148,N_28015);
nand U28860 (N_28860,N_28415,N_28393);
and U28861 (N_28861,N_28326,N_28202);
xnor U28862 (N_28862,N_28364,N_28359);
and U28863 (N_28863,N_28445,N_28487);
xor U28864 (N_28864,N_28366,N_28396);
xnor U28865 (N_28865,N_28183,N_28418);
and U28866 (N_28866,N_28357,N_28139);
or U28867 (N_28867,N_28338,N_28077);
and U28868 (N_28868,N_28317,N_28042);
nor U28869 (N_28869,N_28251,N_28405);
and U28870 (N_28870,N_28486,N_28461);
nand U28871 (N_28871,N_28447,N_28352);
or U28872 (N_28872,N_28335,N_28090);
xor U28873 (N_28873,N_28006,N_28389);
and U28874 (N_28874,N_28330,N_28070);
or U28875 (N_28875,N_28298,N_28371);
nand U28876 (N_28876,N_28247,N_28042);
or U28877 (N_28877,N_28234,N_28283);
xor U28878 (N_28878,N_28296,N_28414);
xnor U28879 (N_28879,N_28136,N_28106);
and U28880 (N_28880,N_28102,N_28128);
xor U28881 (N_28881,N_28389,N_28458);
and U28882 (N_28882,N_28131,N_28473);
or U28883 (N_28883,N_28363,N_28200);
xnor U28884 (N_28884,N_28202,N_28436);
or U28885 (N_28885,N_28494,N_28435);
nand U28886 (N_28886,N_28385,N_28357);
and U28887 (N_28887,N_28296,N_28448);
nor U28888 (N_28888,N_28399,N_28343);
xor U28889 (N_28889,N_28020,N_28446);
nor U28890 (N_28890,N_28254,N_28225);
or U28891 (N_28891,N_28443,N_28489);
nor U28892 (N_28892,N_28469,N_28410);
nor U28893 (N_28893,N_28307,N_28077);
and U28894 (N_28894,N_28274,N_28311);
nand U28895 (N_28895,N_28336,N_28153);
xnor U28896 (N_28896,N_28434,N_28211);
and U28897 (N_28897,N_28233,N_28494);
or U28898 (N_28898,N_28380,N_28498);
nand U28899 (N_28899,N_28156,N_28489);
xor U28900 (N_28900,N_28273,N_28150);
nor U28901 (N_28901,N_28122,N_28487);
or U28902 (N_28902,N_28442,N_28228);
xor U28903 (N_28903,N_28327,N_28322);
or U28904 (N_28904,N_28231,N_28480);
xnor U28905 (N_28905,N_28401,N_28018);
and U28906 (N_28906,N_28174,N_28196);
or U28907 (N_28907,N_28245,N_28216);
xnor U28908 (N_28908,N_28346,N_28176);
nor U28909 (N_28909,N_28149,N_28116);
and U28910 (N_28910,N_28239,N_28153);
and U28911 (N_28911,N_28265,N_28109);
and U28912 (N_28912,N_28212,N_28157);
nor U28913 (N_28913,N_28177,N_28213);
and U28914 (N_28914,N_28048,N_28363);
xnor U28915 (N_28915,N_28106,N_28250);
and U28916 (N_28916,N_28099,N_28344);
nand U28917 (N_28917,N_28416,N_28343);
nor U28918 (N_28918,N_28230,N_28003);
and U28919 (N_28919,N_28184,N_28050);
and U28920 (N_28920,N_28232,N_28451);
nor U28921 (N_28921,N_28319,N_28499);
nand U28922 (N_28922,N_28355,N_28305);
and U28923 (N_28923,N_28235,N_28454);
nor U28924 (N_28924,N_28026,N_28067);
or U28925 (N_28925,N_28222,N_28240);
or U28926 (N_28926,N_28304,N_28229);
and U28927 (N_28927,N_28070,N_28394);
nand U28928 (N_28928,N_28419,N_28054);
nand U28929 (N_28929,N_28055,N_28202);
nor U28930 (N_28930,N_28303,N_28266);
nor U28931 (N_28931,N_28083,N_28371);
nand U28932 (N_28932,N_28162,N_28435);
and U28933 (N_28933,N_28336,N_28297);
nor U28934 (N_28934,N_28495,N_28181);
nand U28935 (N_28935,N_28242,N_28412);
and U28936 (N_28936,N_28298,N_28384);
nor U28937 (N_28937,N_28349,N_28040);
xnor U28938 (N_28938,N_28043,N_28183);
or U28939 (N_28939,N_28080,N_28340);
nor U28940 (N_28940,N_28041,N_28308);
and U28941 (N_28941,N_28321,N_28361);
or U28942 (N_28942,N_28395,N_28461);
nand U28943 (N_28943,N_28093,N_28294);
or U28944 (N_28944,N_28360,N_28088);
xnor U28945 (N_28945,N_28339,N_28340);
and U28946 (N_28946,N_28287,N_28031);
and U28947 (N_28947,N_28046,N_28231);
nor U28948 (N_28948,N_28137,N_28392);
and U28949 (N_28949,N_28453,N_28496);
and U28950 (N_28950,N_28446,N_28248);
or U28951 (N_28951,N_28188,N_28197);
xnor U28952 (N_28952,N_28089,N_28104);
and U28953 (N_28953,N_28081,N_28366);
nor U28954 (N_28954,N_28249,N_28012);
and U28955 (N_28955,N_28074,N_28122);
or U28956 (N_28956,N_28480,N_28466);
nor U28957 (N_28957,N_28238,N_28365);
xnor U28958 (N_28958,N_28147,N_28399);
nand U28959 (N_28959,N_28387,N_28364);
nand U28960 (N_28960,N_28072,N_28244);
nor U28961 (N_28961,N_28426,N_28493);
xnor U28962 (N_28962,N_28434,N_28204);
and U28963 (N_28963,N_28161,N_28434);
and U28964 (N_28964,N_28034,N_28443);
and U28965 (N_28965,N_28285,N_28302);
nor U28966 (N_28966,N_28359,N_28220);
and U28967 (N_28967,N_28490,N_28096);
xor U28968 (N_28968,N_28419,N_28160);
nor U28969 (N_28969,N_28243,N_28069);
or U28970 (N_28970,N_28101,N_28251);
xor U28971 (N_28971,N_28436,N_28165);
and U28972 (N_28972,N_28296,N_28248);
nand U28973 (N_28973,N_28465,N_28425);
nand U28974 (N_28974,N_28453,N_28139);
xor U28975 (N_28975,N_28460,N_28075);
xnor U28976 (N_28976,N_28273,N_28158);
xor U28977 (N_28977,N_28054,N_28294);
nand U28978 (N_28978,N_28072,N_28367);
nand U28979 (N_28979,N_28334,N_28028);
or U28980 (N_28980,N_28348,N_28323);
nand U28981 (N_28981,N_28206,N_28217);
or U28982 (N_28982,N_28056,N_28161);
nor U28983 (N_28983,N_28154,N_28330);
nand U28984 (N_28984,N_28445,N_28309);
and U28985 (N_28985,N_28290,N_28263);
nor U28986 (N_28986,N_28188,N_28363);
nor U28987 (N_28987,N_28195,N_28228);
nand U28988 (N_28988,N_28291,N_28060);
and U28989 (N_28989,N_28099,N_28462);
nand U28990 (N_28990,N_28434,N_28051);
and U28991 (N_28991,N_28432,N_28339);
and U28992 (N_28992,N_28017,N_28186);
and U28993 (N_28993,N_28028,N_28332);
nor U28994 (N_28994,N_28156,N_28000);
or U28995 (N_28995,N_28251,N_28370);
and U28996 (N_28996,N_28444,N_28032);
and U28997 (N_28997,N_28279,N_28440);
and U28998 (N_28998,N_28445,N_28198);
and U28999 (N_28999,N_28496,N_28376);
nand U29000 (N_29000,N_28633,N_28698);
nor U29001 (N_29001,N_28575,N_28923);
nand U29002 (N_29002,N_28825,N_28940);
xor U29003 (N_29003,N_28689,N_28513);
xor U29004 (N_29004,N_28937,N_28659);
nand U29005 (N_29005,N_28595,N_28807);
nor U29006 (N_29006,N_28535,N_28712);
nand U29007 (N_29007,N_28819,N_28510);
nand U29008 (N_29008,N_28610,N_28768);
nand U29009 (N_29009,N_28641,N_28770);
nand U29010 (N_29010,N_28545,N_28881);
nand U29011 (N_29011,N_28994,N_28838);
or U29012 (N_29012,N_28620,N_28817);
and U29013 (N_29013,N_28773,N_28836);
nor U29014 (N_29014,N_28905,N_28721);
nor U29015 (N_29015,N_28814,N_28865);
or U29016 (N_29016,N_28656,N_28928);
nand U29017 (N_29017,N_28806,N_28621);
xnor U29018 (N_29018,N_28753,N_28625);
nor U29019 (N_29019,N_28989,N_28755);
and U29020 (N_29020,N_28781,N_28861);
nor U29021 (N_29021,N_28827,N_28922);
nand U29022 (N_29022,N_28849,N_28606);
nand U29023 (N_29023,N_28846,N_28599);
nand U29024 (N_29024,N_28576,N_28563);
xor U29025 (N_29025,N_28955,N_28952);
nor U29026 (N_29026,N_28505,N_28717);
nand U29027 (N_29027,N_28748,N_28604);
or U29028 (N_29028,N_28616,N_28638);
xnor U29029 (N_29029,N_28672,N_28930);
xnor U29030 (N_29030,N_28701,N_28774);
or U29031 (N_29031,N_28848,N_28822);
nand U29032 (N_29032,N_28757,N_28518);
or U29033 (N_29033,N_28988,N_28824);
and U29034 (N_29034,N_28630,N_28697);
or U29035 (N_29035,N_28670,N_28830);
and U29036 (N_29036,N_28650,N_28761);
nand U29037 (N_29037,N_28565,N_28601);
xnor U29038 (N_29038,N_28767,N_28996);
or U29039 (N_29039,N_28614,N_28653);
or U29040 (N_29040,N_28885,N_28911);
nand U29041 (N_29041,N_28790,N_28629);
nor U29042 (N_29042,N_28933,N_28769);
xnor U29043 (N_29043,N_28847,N_28772);
and U29044 (N_29044,N_28828,N_28809);
nand U29045 (N_29045,N_28637,N_28584);
xor U29046 (N_29046,N_28890,N_28731);
or U29047 (N_29047,N_28871,N_28939);
nor U29048 (N_29048,N_28583,N_28560);
nand U29049 (N_29049,N_28805,N_28738);
nand U29050 (N_29050,N_28547,N_28568);
or U29051 (N_29051,N_28646,N_28713);
or U29052 (N_29052,N_28623,N_28661);
xnor U29053 (N_29053,N_28894,N_28617);
nand U29054 (N_29054,N_28876,N_28808);
or U29055 (N_29055,N_28874,N_28677);
and U29056 (N_29056,N_28749,N_28634);
or U29057 (N_29057,N_28973,N_28700);
nor U29058 (N_29058,N_28826,N_28694);
or U29059 (N_29059,N_28877,N_28503);
or U29060 (N_29060,N_28938,N_28902);
and U29061 (N_29061,N_28691,N_28602);
and U29062 (N_29062,N_28746,N_28685);
and U29063 (N_29063,N_28934,N_28997);
xor U29064 (N_29064,N_28715,N_28907);
nor U29065 (N_29065,N_28744,N_28842);
xor U29066 (N_29066,N_28858,N_28974);
nand U29067 (N_29067,N_28887,N_28561);
xnor U29068 (N_29068,N_28534,N_28862);
or U29069 (N_29069,N_28631,N_28850);
and U29070 (N_29070,N_28765,N_28540);
and U29071 (N_29071,N_28792,N_28883);
nand U29072 (N_29072,N_28558,N_28794);
and U29073 (N_29073,N_28798,N_28758);
nor U29074 (N_29074,N_28981,N_28737);
nor U29075 (N_29075,N_28867,N_28780);
or U29076 (N_29076,N_28980,N_28581);
or U29077 (N_29077,N_28864,N_28705);
or U29078 (N_29078,N_28533,N_28736);
nand U29079 (N_29079,N_28951,N_28692);
nand U29080 (N_29080,N_28869,N_28756);
or U29081 (N_29081,N_28734,N_28608);
or U29082 (N_29082,N_28896,N_28801);
or U29083 (N_29083,N_28530,N_28956);
and U29084 (N_29084,N_28762,N_28802);
nor U29085 (N_29085,N_28859,N_28512);
or U29086 (N_29086,N_28524,N_28613);
nand U29087 (N_29087,N_28607,N_28949);
nor U29088 (N_29088,N_28516,N_28984);
xor U29089 (N_29089,N_28562,N_28569);
nand U29090 (N_29090,N_28912,N_28662);
and U29091 (N_29091,N_28789,N_28779);
and U29092 (N_29092,N_28622,N_28666);
nor U29093 (N_29093,N_28908,N_28525);
xnor U29094 (N_29094,N_28915,N_28796);
xnor U29095 (N_29095,N_28711,N_28910);
xor U29096 (N_29096,N_28571,N_28961);
xnor U29097 (N_29097,N_28985,N_28708);
nand U29098 (N_29098,N_28935,N_28799);
or U29099 (N_29099,N_28987,N_28777);
or U29100 (N_29100,N_28900,N_28570);
xnor U29101 (N_29101,N_28831,N_28893);
and U29102 (N_29102,N_28932,N_28722);
or U29103 (N_29103,N_28837,N_28918);
and U29104 (N_29104,N_28784,N_28751);
or U29105 (N_29105,N_28600,N_28926);
or U29106 (N_29106,N_28660,N_28793);
nor U29107 (N_29107,N_28615,N_28964);
xor U29108 (N_29108,N_28603,N_28797);
nor U29109 (N_29109,N_28742,N_28840);
xnor U29110 (N_29110,N_28959,N_28665);
and U29111 (N_29111,N_28668,N_28611);
nor U29112 (N_29112,N_28657,N_28948);
nor U29113 (N_29113,N_28716,N_28550);
nor U29114 (N_29114,N_28976,N_28536);
and U29115 (N_29115,N_28592,N_28555);
xnor U29116 (N_29116,N_28573,N_28841);
or U29117 (N_29117,N_28818,N_28892);
or U29118 (N_29118,N_28686,N_28690);
and U29119 (N_29119,N_28674,N_28795);
and U29120 (N_29120,N_28834,N_28971);
and U29121 (N_29121,N_28760,N_28995);
and U29122 (N_29122,N_28552,N_28947);
and U29123 (N_29123,N_28658,N_28855);
nand U29124 (N_29124,N_28803,N_28702);
nand U29125 (N_29125,N_28732,N_28618);
xnor U29126 (N_29126,N_28577,N_28624);
xor U29127 (N_29127,N_28587,N_28927);
nor U29128 (N_29128,N_28645,N_28632);
xnor U29129 (N_29129,N_28649,N_28517);
and U29130 (N_29130,N_28833,N_28598);
nor U29131 (N_29131,N_28925,N_28875);
xnor U29132 (N_29132,N_28519,N_28782);
nor U29133 (N_29133,N_28978,N_28763);
or U29134 (N_29134,N_28678,N_28663);
nor U29135 (N_29135,N_28709,N_28993);
nand U29136 (N_29136,N_28566,N_28655);
and U29137 (N_29137,N_28707,N_28856);
xnor U29138 (N_29138,N_28917,N_28853);
and U29139 (N_29139,N_28943,N_28870);
or U29140 (N_29140,N_28586,N_28648);
xor U29141 (N_29141,N_28886,N_28747);
or U29142 (N_29142,N_28729,N_28704);
nand U29143 (N_29143,N_28873,N_28529);
or U29144 (N_29144,N_28537,N_28639);
or U29145 (N_29145,N_28636,N_28627);
nor U29146 (N_29146,N_28843,N_28968);
or U29147 (N_29147,N_28673,N_28728);
xor U29148 (N_29148,N_28942,N_28548);
xnor U29149 (N_29149,N_28889,N_28965);
or U29150 (N_29150,N_28733,N_28844);
nor U29151 (N_29151,N_28787,N_28580);
nand U29152 (N_29152,N_28643,N_28596);
xor U29153 (N_29153,N_28970,N_28866);
and U29154 (N_29154,N_28944,N_28754);
nor U29155 (N_29155,N_28688,N_28546);
nand U29156 (N_29156,N_28967,N_28557);
nand U29157 (N_29157,N_28791,N_28872);
nand U29158 (N_29158,N_28868,N_28594);
and U29159 (N_29159,N_28878,N_28882);
nand U29160 (N_29160,N_28998,N_28879);
and U29161 (N_29161,N_28609,N_28654);
xor U29162 (N_29162,N_28936,N_28589);
and U29163 (N_29163,N_28695,N_28593);
xnor U29164 (N_29164,N_28644,N_28785);
nand U29165 (N_29165,N_28854,N_28921);
xnor U29166 (N_29166,N_28895,N_28820);
nand U29167 (N_29167,N_28945,N_28521);
nor U29168 (N_29168,N_28941,N_28914);
nor U29169 (N_29169,N_28913,N_28640);
or U29170 (N_29170,N_28696,N_28954);
and U29171 (N_29171,N_28664,N_28515);
nor U29172 (N_29172,N_28815,N_28813);
nor U29173 (N_29173,N_28986,N_28901);
nor U29174 (N_29174,N_28983,N_28832);
nor U29175 (N_29175,N_28681,N_28906);
and U29176 (N_29176,N_28582,N_28891);
nor U29177 (N_29177,N_28863,N_28591);
xnor U29178 (N_29178,N_28679,N_28554);
or U29179 (N_29179,N_28957,N_28706);
nand U29180 (N_29180,N_28740,N_28538);
and U29181 (N_29181,N_28739,N_28924);
or U29182 (N_29182,N_28542,N_28991);
nor U29183 (N_29183,N_28647,N_28680);
xor U29184 (N_29184,N_28682,N_28719);
and U29185 (N_29185,N_28528,N_28675);
or U29186 (N_29186,N_28743,N_28730);
xor U29187 (N_29187,N_28597,N_28898);
nand U29188 (N_29188,N_28975,N_28523);
or U29189 (N_29189,N_28635,N_28931);
and U29190 (N_29190,N_28553,N_28511);
or U29191 (N_29191,N_28823,N_28508);
nand U29192 (N_29192,N_28960,N_28860);
xor U29193 (N_29193,N_28816,N_28720);
nand U29194 (N_29194,N_28963,N_28990);
or U29195 (N_29195,N_28556,N_28909);
xor U29196 (N_29196,N_28771,N_28532);
and U29197 (N_29197,N_28999,N_28544);
xor U29198 (N_29198,N_28919,N_28946);
or U29199 (N_29199,N_28852,N_28526);
xor U29200 (N_29200,N_28506,N_28880);
or U29201 (N_29201,N_28651,N_28687);
xnor U29202 (N_29202,N_28966,N_28703);
nor U29203 (N_29203,N_28903,N_28543);
xor U29204 (N_29204,N_28509,N_28962);
nand U29205 (N_29205,N_28958,N_28588);
and U29206 (N_29206,N_28501,N_28851);
nand U29207 (N_29207,N_28775,N_28969);
and U29208 (N_29208,N_28590,N_28745);
or U29209 (N_29209,N_28857,N_28741);
and U29210 (N_29210,N_28725,N_28531);
nand U29211 (N_29211,N_28502,N_28992);
xnor U29212 (N_29212,N_28735,N_28829);
xor U29213 (N_29213,N_28626,N_28839);
or U29214 (N_29214,N_28888,N_28667);
nor U29215 (N_29215,N_28527,N_28953);
nor U29216 (N_29216,N_28950,N_28564);
xor U29217 (N_29217,N_28619,N_28710);
nand U29218 (N_29218,N_28551,N_28788);
or U29219 (N_29219,N_28759,N_28549);
xor U29220 (N_29220,N_28642,N_28752);
nor U29221 (N_29221,N_28628,N_28776);
xnor U29222 (N_29222,N_28579,N_28567);
nand U29223 (N_29223,N_28574,N_28714);
nor U29224 (N_29224,N_28884,N_28500);
and U29225 (N_29225,N_28764,N_28520);
and U29226 (N_29226,N_28676,N_28671);
and U29227 (N_29227,N_28904,N_28804);
xnor U29228 (N_29228,N_28559,N_28612);
or U29229 (N_29229,N_28522,N_28578);
nand U29230 (N_29230,N_28699,N_28541);
and U29231 (N_29231,N_28800,N_28605);
nor U29232 (N_29232,N_28726,N_28982);
nand U29233 (N_29233,N_28972,N_28718);
nand U29234 (N_29234,N_28979,N_28897);
or U29235 (N_29235,N_28810,N_28899);
nand U29236 (N_29236,N_28652,N_28766);
nand U29237 (N_29237,N_28835,N_28916);
and U29238 (N_29238,N_28920,N_28669);
nor U29239 (N_29239,N_28929,N_28683);
or U29240 (N_29240,N_28811,N_28572);
nor U29241 (N_29241,N_28845,N_28539);
nor U29242 (N_29242,N_28504,N_28514);
xor U29243 (N_29243,N_28727,N_28507);
and U29244 (N_29244,N_28693,N_28783);
and U29245 (N_29245,N_28812,N_28977);
or U29246 (N_29246,N_28585,N_28684);
nor U29247 (N_29247,N_28778,N_28750);
xor U29248 (N_29248,N_28821,N_28786);
xnor U29249 (N_29249,N_28724,N_28723);
nor U29250 (N_29250,N_28581,N_28954);
and U29251 (N_29251,N_28554,N_28720);
xor U29252 (N_29252,N_28564,N_28685);
or U29253 (N_29253,N_28792,N_28544);
nor U29254 (N_29254,N_28946,N_28921);
or U29255 (N_29255,N_28541,N_28533);
xor U29256 (N_29256,N_28782,N_28986);
or U29257 (N_29257,N_28821,N_28913);
and U29258 (N_29258,N_28920,N_28977);
and U29259 (N_29259,N_28778,N_28988);
or U29260 (N_29260,N_28756,N_28974);
nand U29261 (N_29261,N_28934,N_28689);
or U29262 (N_29262,N_28643,N_28825);
and U29263 (N_29263,N_28848,N_28666);
and U29264 (N_29264,N_28950,N_28760);
nand U29265 (N_29265,N_28517,N_28559);
xnor U29266 (N_29266,N_28855,N_28791);
nor U29267 (N_29267,N_28813,N_28985);
xor U29268 (N_29268,N_28851,N_28652);
and U29269 (N_29269,N_28564,N_28851);
nand U29270 (N_29270,N_28935,N_28610);
nand U29271 (N_29271,N_28952,N_28684);
and U29272 (N_29272,N_28787,N_28501);
xnor U29273 (N_29273,N_28638,N_28571);
nor U29274 (N_29274,N_28973,N_28555);
nor U29275 (N_29275,N_28567,N_28561);
or U29276 (N_29276,N_28550,N_28751);
xor U29277 (N_29277,N_28682,N_28669);
nor U29278 (N_29278,N_28907,N_28708);
nand U29279 (N_29279,N_28569,N_28593);
nor U29280 (N_29280,N_28558,N_28966);
nor U29281 (N_29281,N_28635,N_28978);
nor U29282 (N_29282,N_28917,N_28621);
or U29283 (N_29283,N_28846,N_28830);
or U29284 (N_29284,N_28709,N_28510);
nor U29285 (N_29285,N_28501,N_28740);
or U29286 (N_29286,N_28891,N_28983);
nand U29287 (N_29287,N_28925,N_28674);
or U29288 (N_29288,N_28853,N_28511);
nand U29289 (N_29289,N_28633,N_28574);
nor U29290 (N_29290,N_28770,N_28659);
nor U29291 (N_29291,N_28816,N_28808);
xnor U29292 (N_29292,N_28649,N_28647);
nor U29293 (N_29293,N_28518,N_28523);
nor U29294 (N_29294,N_28610,N_28661);
xnor U29295 (N_29295,N_28834,N_28865);
xnor U29296 (N_29296,N_28666,N_28660);
nand U29297 (N_29297,N_28724,N_28963);
nor U29298 (N_29298,N_28539,N_28820);
and U29299 (N_29299,N_28927,N_28950);
nor U29300 (N_29300,N_28644,N_28976);
nor U29301 (N_29301,N_28543,N_28817);
and U29302 (N_29302,N_28581,N_28619);
xor U29303 (N_29303,N_28514,N_28832);
and U29304 (N_29304,N_28514,N_28791);
nand U29305 (N_29305,N_28742,N_28834);
and U29306 (N_29306,N_28668,N_28738);
nor U29307 (N_29307,N_28605,N_28916);
xnor U29308 (N_29308,N_28609,N_28650);
nor U29309 (N_29309,N_28681,N_28672);
nand U29310 (N_29310,N_28887,N_28925);
nand U29311 (N_29311,N_28649,N_28543);
nand U29312 (N_29312,N_28849,N_28742);
and U29313 (N_29313,N_28847,N_28539);
nand U29314 (N_29314,N_28963,N_28702);
or U29315 (N_29315,N_28633,N_28950);
xnor U29316 (N_29316,N_28827,N_28979);
nor U29317 (N_29317,N_28814,N_28978);
nor U29318 (N_29318,N_28582,N_28649);
xnor U29319 (N_29319,N_28810,N_28511);
xor U29320 (N_29320,N_28562,N_28550);
or U29321 (N_29321,N_28631,N_28678);
or U29322 (N_29322,N_28566,N_28992);
xor U29323 (N_29323,N_28796,N_28856);
nand U29324 (N_29324,N_28556,N_28839);
or U29325 (N_29325,N_28816,N_28590);
xor U29326 (N_29326,N_28936,N_28617);
or U29327 (N_29327,N_28924,N_28880);
xnor U29328 (N_29328,N_28757,N_28789);
xnor U29329 (N_29329,N_28774,N_28509);
xor U29330 (N_29330,N_28757,N_28979);
and U29331 (N_29331,N_28931,N_28996);
nor U29332 (N_29332,N_28707,N_28623);
or U29333 (N_29333,N_28651,N_28792);
or U29334 (N_29334,N_28521,N_28557);
or U29335 (N_29335,N_28755,N_28667);
or U29336 (N_29336,N_28733,N_28910);
or U29337 (N_29337,N_28573,N_28526);
nor U29338 (N_29338,N_28767,N_28617);
xnor U29339 (N_29339,N_28850,N_28510);
or U29340 (N_29340,N_28580,N_28714);
nand U29341 (N_29341,N_28544,N_28718);
and U29342 (N_29342,N_28939,N_28544);
nand U29343 (N_29343,N_28839,N_28933);
nand U29344 (N_29344,N_28510,N_28993);
or U29345 (N_29345,N_28705,N_28613);
nor U29346 (N_29346,N_28998,N_28749);
and U29347 (N_29347,N_28749,N_28538);
nand U29348 (N_29348,N_28904,N_28824);
nand U29349 (N_29349,N_28790,N_28896);
nor U29350 (N_29350,N_28974,N_28661);
xor U29351 (N_29351,N_28722,N_28653);
nand U29352 (N_29352,N_28803,N_28816);
nand U29353 (N_29353,N_28507,N_28872);
or U29354 (N_29354,N_28704,N_28833);
or U29355 (N_29355,N_28714,N_28659);
and U29356 (N_29356,N_28598,N_28524);
and U29357 (N_29357,N_28729,N_28956);
nand U29358 (N_29358,N_28863,N_28768);
nor U29359 (N_29359,N_28572,N_28733);
xnor U29360 (N_29360,N_28623,N_28806);
xnor U29361 (N_29361,N_28910,N_28922);
nand U29362 (N_29362,N_28517,N_28634);
nand U29363 (N_29363,N_28979,N_28690);
nand U29364 (N_29364,N_28728,N_28932);
and U29365 (N_29365,N_28941,N_28549);
and U29366 (N_29366,N_28555,N_28733);
nor U29367 (N_29367,N_28703,N_28595);
xnor U29368 (N_29368,N_28533,N_28572);
nor U29369 (N_29369,N_28906,N_28575);
nor U29370 (N_29370,N_28539,N_28834);
nor U29371 (N_29371,N_28517,N_28565);
xnor U29372 (N_29372,N_28593,N_28756);
and U29373 (N_29373,N_28862,N_28782);
and U29374 (N_29374,N_28926,N_28813);
nand U29375 (N_29375,N_28883,N_28905);
and U29376 (N_29376,N_28990,N_28638);
and U29377 (N_29377,N_28975,N_28742);
or U29378 (N_29378,N_28970,N_28632);
xnor U29379 (N_29379,N_28510,N_28751);
nor U29380 (N_29380,N_28596,N_28547);
nor U29381 (N_29381,N_28741,N_28637);
xnor U29382 (N_29382,N_28966,N_28760);
and U29383 (N_29383,N_28683,N_28707);
or U29384 (N_29384,N_28660,N_28863);
nand U29385 (N_29385,N_28870,N_28511);
and U29386 (N_29386,N_28676,N_28788);
nand U29387 (N_29387,N_28644,N_28599);
nand U29388 (N_29388,N_28548,N_28881);
and U29389 (N_29389,N_28933,N_28580);
nand U29390 (N_29390,N_28703,N_28998);
nand U29391 (N_29391,N_28690,N_28584);
or U29392 (N_29392,N_28981,N_28595);
nand U29393 (N_29393,N_28700,N_28926);
xnor U29394 (N_29394,N_28797,N_28526);
and U29395 (N_29395,N_28941,N_28827);
xnor U29396 (N_29396,N_28803,N_28556);
nand U29397 (N_29397,N_28627,N_28626);
or U29398 (N_29398,N_28961,N_28611);
nor U29399 (N_29399,N_28776,N_28815);
or U29400 (N_29400,N_28719,N_28862);
nor U29401 (N_29401,N_28936,N_28735);
or U29402 (N_29402,N_28704,N_28767);
nor U29403 (N_29403,N_28863,N_28621);
nand U29404 (N_29404,N_28925,N_28543);
or U29405 (N_29405,N_28638,N_28773);
and U29406 (N_29406,N_28715,N_28905);
nor U29407 (N_29407,N_28549,N_28554);
and U29408 (N_29408,N_28927,N_28973);
or U29409 (N_29409,N_28857,N_28612);
nor U29410 (N_29410,N_28998,N_28696);
nand U29411 (N_29411,N_28571,N_28977);
or U29412 (N_29412,N_28776,N_28538);
nand U29413 (N_29413,N_28968,N_28798);
nand U29414 (N_29414,N_28820,N_28754);
nor U29415 (N_29415,N_28657,N_28793);
and U29416 (N_29416,N_28543,N_28922);
nand U29417 (N_29417,N_28534,N_28688);
or U29418 (N_29418,N_28958,N_28718);
nor U29419 (N_29419,N_28932,N_28860);
xnor U29420 (N_29420,N_28964,N_28626);
nor U29421 (N_29421,N_28707,N_28666);
nor U29422 (N_29422,N_28818,N_28857);
or U29423 (N_29423,N_28695,N_28863);
xor U29424 (N_29424,N_28910,N_28689);
and U29425 (N_29425,N_28843,N_28989);
and U29426 (N_29426,N_28769,N_28878);
nor U29427 (N_29427,N_28931,N_28756);
or U29428 (N_29428,N_28725,N_28786);
or U29429 (N_29429,N_28786,N_28713);
nand U29430 (N_29430,N_28857,N_28967);
nand U29431 (N_29431,N_28743,N_28668);
and U29432 (N_29432,N_28607,N_28968);
or U29433 (N_29433,N_28724,N_28698);
nand U29434 (N_29434,N_28541,N_28579);
or U29435 (N_29435,N_28588,N_28976);
nand U29436 (N_29436,N_28815,N_28674);
and U29437 (N_29437,N_28646,N_28539);
nand U29438 (N_29438,N_28525,N_28719);
and U29439 (N_29439,N_28708,N_28710);
nand U29440 (N_29440,N_28720,N_28810);
nand U29441 (N_29441,N_28659,N_28841);
nor U29442 (N_29442,N_28745,N_28859);
xnor U29443 (N_29443,N_28602,N_28564);
xor U29444 (N_29444,N_28669,N_28532);
nand U29445 (N_29445,N_28538,N_28565);
nand U29446 (N_29446,N_28711,N_28872);
xor U29447 (N_29447,N_28681,N_28945);
and U29448 (N_29448,N_28883,N_28610);
or U29449 (N_29449,N_28556,N_28660);
and U29450 (N_29450,N_28953,N_28662);
nor U29451 (N_29451,N_28905,N_28893);
nand U29452 (N_29452,N_28968,N_28852);
nand U29453 (N_29453,N_28805,N_28769);
nand U29454 (N_29454,N_28672,N_28923);
xor U29455 (N_29455,N_28718,N_28638);
xor U29456 (N_29456,N_28706,N_28682);
nand U29457 (N_29457,N_28532,N_28953);
xor U29458 (N_29458,N_28566,N_28932);
xor U29459 (N_29459,N_28875,N_28515);
nand U29460 (N_29460,N_28778,N_28731);
nor U29461 (N_29461,N_28942,N_28665);
nand U29462 (N_29462,N_28642,N_28896);
and U29463 (N_29463,N_28664,N_28934);
xnor U29464 (N_29464,N_28747,N_28561);
nor U29465 (N_29465,N_28919,N_28897);
nand U29466 (N_29466,N_28950,N_28586);
nor U29467 (N_29467,N_28731,N_28658);
and U29468 (N_29468,N_28967,N_28786);
xor U29469 (N_29469,N_28779,N_28833);
nor U29470 (N_29470,N_28699,N_28991);
nand U29471 (N_29471,N_28695,N_28832);
or U29472 (N_29472,N_28950,N_28977);
xnor U29473 (N_29473,N_28594,N_28654);
and U29474 (N_29474,N_28915,N_28576);
nand U29475 (N_29475,N_28758,N_28934);
xnor U29476 (N_29476,N_28657,N_28527);
nand U29477 (N_29477,N_28927,N_28550);
nor U29478 (N_29478,N_28884,N_28571);
xor U29479 (N_29479,N_28751,N_28732);
nor U29480 (N_29480,N_28943,N_28577);
and U29481 (N_29481,N_28844,N_28945);
or U29482 (N_29482,N_28510,N_28876);
and U29483 (N_29483,N_28894,N_28644);
nor U29484 (N_29484,N_28504,N_28863);
xor U29485 (N_29485,N_28787,N_28687);
and U29486 (N_29486,N_28661,N_28796);
nor U29487 (N_29487,N_28737,N_28716);
nand U29488 (N_29488,N_28603,N_28618);
or U29489 (N_29489,N_28959,N_28572);
or U29490 (N_29490,N_28761,N_28644);
xor U29491 (N_29491,N_28789,N_28629);
nand U29492 (N_29492,N_28971,N_28940);
nor U29493 (N_29493,N_28560,N_28763);
and U29494 (N_29494,N_28961,N_28806);
and U29495 (N_29495,N_28746,N_28897);
nand U29496 (N_29496,N_28734,N_28738);
or U29497 (N_29497,N_28621,N_28818);
nor U29498 (N_29498,N_28655,N_28572);
nor U29499 (N_29499,N_28592,N_28998);
nor U29500 (N_29500,N_29333,N_29270);
nor U29501 (N_29501,N_29059,N_29140);
or U29502 (N_29502,N_29108,N_29267);
xor U29503 (N_29503,N_29379,N_29339);
xor U29504 (N_29504,N_29056,N_29451);
or U29505 (N_29505,N_29168,N_29234);
and U29506 (N_29506,N_29143,N_29118);
and U29507 (N_29507,N_29452,N_29362);
or U29508 (N_29508,N_29001,N_29039);
or U29509 (N_29509,N_29232,N_29058);
nor U29510 (N_29510,N_29250,N_29368);
xor U29511 (N_29511,N_29054,N_29121);
xor U29512 (N_29512,N_29315,N_29133);
xor U29513 (N_29513,N_29354,N_29295);
xnor U29514 (N_29514,N_29312,N_29216);
xor U29515 (N_29515,N_29181,N_29390);
and U29516 (N_29516,N_29255,N_29161);
nand U29517 (N_29517,N_29005,N_29188);
nand U29518 (N_29518,N_29002,N_29423);
xor U29519 (N_29519,N_29170,N_29240);
nand U29520 (N_29520,N_29266,N_29110);
xor U29521 (N_29521,N_29171,N_29237);
and U29522 (N_29522,N_29046,N_29061);
nor U29523 (N_29523,N_29205,N_29086);
xor U29524 (N_29524,N_29319,N_29416);
and U29525 (N_29525,N_29230,N_29404);
nand U29526 (N_29526,N_29100,N_29067);
nor U29527 (N_29527,N_29342,N_29124);
nor U29528 (N_29528,N_29411,N_29218);
and U29529 (N_29529,N_29183,N_29274);
nand U29530 (N_29530,N_29474,N_29034);
nor U29531 (N_29531,N_29003,N_29441);
or U29532 (N_29532,N_29393,N_29248);
nor U29533 (N_29533,N_29469,N_29285);
xor U29534 (N_29534,N_29006,N_29211);
nor U29535 (N_29535,N_29460,N_29291);
nor U29536 (N_29536,N_29208,N_29444);
nand U29537 (N_29537,N_29485,N_29296);
and U29538 (N_29538,N_29155,N_29226);
nand U29539 (N_29539,N_29088,N_29048);
xnor U29540 (N_29540,N_29357,N_29253);
nor U29541 (N_29541,N_29350,N_29351);
nor U29542 (N_29542,N_29464,N_29343);
xnor U29543 (N_29543,N_29047,N_29182);
xnor U29544 (N_29544,N_29468,N_29269);
xnor U29545 (N_29545,N_29413,N_29305);
xnor U29546 (N_29546,N_29377,N_29224);
nor U29547 (N_29547,N_29137,N_29299);
nand U29548 (N_29548,N_29284,N_29060);
or U29549 (N_29549,N_29113,N_29134);
nor U29550 (N_29550,N_29263,N_29349);
nand U29551 (N_29551,N_29149,N_29281);
and U29552 (N_29552,N_29355,N_29432);
xnor U29553 (N_29553,N_29438,N_29217);
nand U29554 (N_29554,N_29370,N_29220);
and U29555 (N_29555,N_29273,N_29352);
and U29556 (N_29556,N_29114,N_29311);
xor U29557 (N_29557,N_29064,N_29304);
nor U29558 (N_29558,N_29051,N_29150);
and U29559 (N_29559,N_29026,N_29077);
nand U29560 (N_29560,N_29489,N_29303);
and U29561 (N_29561,N_29463,N_29309);
nor U29562 (N_29562,N_29245,N_29418);
or U29563 (N_29563,N_29102,N_29282);
and U29564 (N_29564,N_29279,N_29254);
or U29565 (N_29565,N_29195,N_29020);
nand U29566 (N_29566,N_29018,N_29019);
and U29567 (N_29567,N_29201,N_29098);
nand U29568 (N_29568,N_29175,N_29180);
or U29569 (N_29569,N_29154,N_29128);
xnor U29570 (N_29570,N_29496,N_29314);
xnor U29571 (N_29571,N_29089,N_29122);
nor U29572 (N_29572,N_29052,N_29109);
and U29573 (N_29573,N_29417,N_29112);
nor U29574 (N_29574,N_29385,N_29453);
and U29575 (N_29575,N_29041,N_29492);
and U29576 (N_29576,N_29111,N_29027);
or U29577 (N_29577,N_29142,N_29164);
or U29578 (N_29578,N_29206,N_29029);
nand U29579 (N_29579,N_29317,N_29144);
nor U29580 (N_29580,N_29210,N_29330);
xnor U29581 (N_29581,N_29448,N_29367);
nand U29582 (N_29582,N_29159,N_29425);
nor U29583 (N_29583,N_29038,N_29000);
nor U29584 (N_29584,N_29035,N_29461);
and U29585 (N_29585,N_29127,N_29410);
or U29586 (N_29586,N_29078,N_29467);
xor U29587 (N_29587,N_29225,N_29079);
or U29588 (N_29588,N_29387,N_29459);
nand U29589 (N_29589,N_29158,N_29341);
or U29590 (N_29590,N_29141,N_29251);
nor U29591 (N_29591,N_29294,N_29262);
xor U29592 (N_29592,N_29353,N_29033);
or U29593 (N_29593,N_29169,N_29439);
or U29594 (N_29594,N_29484,N_29247);
or U29595 (N_29595,N_29243,N_29381);
xnor U29596 (N_29596,N_29152,N_29493);
and U29597 (N_29597,N_29313,N_29236);
xnor U29598 (N_29598,N_29395,N_29406);
xor U29599 (N_29599,N_29443,N_29199);
and U29600 (N_29600,N_29455,N_29010);
or U29601 (N_29601,N_29322,N_29136);
or U29602 (N_29602,N_29446,N_29457);
and U29603 (N_29603,N_29196,N_29138);
and U29604 (N_29604,N_29380,N_29099);
nor U29605 (N_29605,N_29289,N_29016);
or U29606 (N_29606,N_29096,N_29332);
and U29607 (N_29607,N_29302,N_29495);
xor U29608 (N_29608,N_29065,N_29049);
and U29609 (N_29609,N_29372,N_29132);
nand U29610 (N_29610,N_29095,N_29335);
nor U29611 (N_29611,N_29326,N_29375);
and U29612 (N_29612,N_29360,N_29371);
or U29613 (N_29613,N_29456,N_29013);
nand U29614 (N_29614,N_29376,N_29229);
and U29615 (N_29615,N_29298,N_29478);
and U29616 (N_29616,N_29241,N_29084);
xor U29617 (N_29617,N_29090,N_29081);
nand U29618 (N_29618,N_29023,N_29440);
or U29619 (N_29619,N_29076,N_29431);
nand U29620 (N_29620,N_29361,N_29306);
nand U29621 (N_29621,N_29369,N_29388);
nand U29622 (N_29622,N_29153,N_29396);
nand U29623 (N_29623,N_29080,N_29024);
or U29624 (N_29624,N_29400,N_29359);
and U29625 (N_29625,N_29030,N_29454);
or U29626 (N_29626,N_29316,N_29186);
xor U29627 (N_29627,N_29437,N_29257);
nor U29628 (N_29628,N_29340,N_29363);
and U29629 (N_29629,N_29106,N_29366);
or U29630 (N_29630,N_29070,N_29045);
nand U29631 (N_29631,N_29374,N_29307);
nand U29632 (N_29632,N_29085,N_29204);
nor U29633 (N_29633,N_29043,N_29434);
and U29634 (N_29634,N_29336,N_29117);
nor U29635 (N_29635,N_29429,N_29462);
nor U29636 (N_29636,N_29198,N_29228);
nor U29637 (N_29637,N_29223,N_29233);
nand U29638 (N_29638,N_29399,N_29057);
and U29639 (N_29639,N_29156,N_29215);
nor U29640 (N_29640,N_29063,N_29116);
xor U29641 (N_29641,N_29480,N_29092);
and U29642 (N_29642,N_29483,N_29135);
nor U29643 (N_29643,N_29194,N_29346);
nor U29644 (N_29644,N_29207,N_29356);
or U29645 (N_29645,N_29288,N_29327);
nand U29646 (N_29646,N_29166,N_29412);
and U29647 (N_29647,N_29261,N_29308);
nor U29648 (N_29648,N_29197,N_29328);
nor U29649 (N_29649,N_29214,N_29075);
xor U29650 (N_29650,N_29490,N_29293);
and U29651 (N_29651,N_29465,N_29222);
or U29652 (N_29652,N_29264,N_29147);
xor U29653 (N_29653,N_29424,N_29238);
nor U29654 (N_29654,N_29012,N_29320);
xnor U29655 (N_29655,N_29348,N_29126);
nand U29656 (N_29656,N_29373,N_29394);
and U29657 (N_29657,N_29167,N_29325);
nand U29658 (N_29658,N_29402,N_29358);
nand U29659 (N_29659,N_29329,N_29097);
nor U29660 (N_29660,N_29022,N_29292);
nand U29661 (N_29661,N_29318,N_29249);
and U29662 (N_29662,N_29481,N_29179);
or U29663 (N_29663,N_29157,N_29244);
nor U29664 (N_29664,N_29259,N_29151);
nor U29665 (N_29665,N_29470,N_29119);
and U29666 (N_29666,N_29290,N_29338);
or U29667 (N_29667,N_29074,N_29212);
xor U29668 (N_29668,N_29301,N_29202);
nand U29669 (N_29669,N_29331,N_29407);
and U29670 (N_29670,N_29025,N_29203);
nor U29671 (N_29671,N_29040,N_29475);
and U29672 (N_29672,N_29105,N_29130);
and U29673 (N_29673,N_29382,N_29146);
xor U29674 (N_29674,N_29427,N_29187);
or U29675 (N_29675,N_29242,N_29428);
nand U29676 (N_29676,N_29184,N_29277);
and U29677 (N_29677,N_29386,N_29499);
xor U29678 (N_29678,N_29486,N_29466);
xnor U29679 (N_29679,N_29120,N_29445);
nor U29680 (N_29680,N_29472,N_29014);
or U29681 (N_29681,N_29174,N_29419);
or U29682 (N_29682,N_29031,N_29072);
nor U29683 (N_29683,N_29408,N_29071);
nor U29684 (N_29684,N_29433,N_29115);
and U29685 (N_29685,N_29053,N_29378);
or U29686 (N_29686,N_29011,N_29148);
or U29687 (N_29687,N_29213,N_29276);
or U29688 (N_29688,N_29017,N_29091);
xor U29689 (N_29689,N_29401,N_29477);
or U29690 (N_29690,N_29103,N_29258);
and U29691 (N_29691,N_29246,N_29347);
xnor U29692 (N_29692,N_29278,N_29287);
nor U29693 (N_29693,N_29310,N_29163);
xor U29694 (N_29694,N_29009,N_29383);
or U29695 (N_29695,N_29389,N_29272);
nor U29696 (N_29696,N_29344,N_29323);
and U29697 (N_29697,N_29435,N_29008);
and U29698 (N_29698,N_29032,N_29256);
or U29699 (N_29699,N_29283,N_29069);
xor U29700 (N_29700,N_29442,N_29028);
xor U29701 (N_29701,N_29414,N_29449);
nand U29702 (N_29702,N_29139,N_29173);
nor U29703 (N_29703,N_29055,N_29337);
xor U29704 (N_29704,N_29300,N_29007);
nor U29705 (N_29705,N_29062,N_29491);
and U29706 (N_29706,N_29365,N_29498);
nor U29707 (N_29707,N_29107,N_29403);
xnor U29708 (N_29708,N_29021,N_29044);
xnor U29709 (N_29709,N_29082,N_29398);
nand U29710 (N_29710,N_29482,N_29123);
nor U29711 (N_29711,N_29036,N_29190);
xnor U29712 (N_29712,N_29479,N_29066);
nor U29713 (N_29713,N_29176,N_29209);
or U29714 (N_29714,N_29420,N_29131);
and U29715 (N_29715,N_29042,N_29200);
nand U29716 (N_29716,N_29297,N_29487);
and U29717 (N_29717,N_29391,N_29129);
nand U29718 (N_29718,N_29145,N_29193);
nand U29719 (N_29719,N_29177,N_29260);
or U29720 (N_29720,N_29405,N_29345);
and U29721 (N_29721,N_29235,N_29037);
nand U29722 (N_29722,N_29015,N_29172);
nand U29723 (N_29723,N_29286,N_29321);
or U29724 (N_29724,N_29231,N_29068);
xnor U29725 (N_29725,N_29497,N_29004);
nand U29726 (N_29726,N_29268,N_29422);
and U29727 (N_29727,N_29471,N_29073);
and U29728 (N_29728,N_29165,N_29421);
nand U29729 (N_29729,N_29227,N_29488);
and U29730 (N_29730,N_29275,N_29280);
xnor U29731 (N_29731,N_29473,N_29185);
or U29732 (N_29732,N_29101,N_29094);
or U29733 (N_29733,N_29271,N_29426);
and U29734 (N_29734,N_29436,N_29397);
nand U29735 (N_29735,N_29409,N_29191);
xnor U29736 (N_29736,N_29050,N_29324);
nor U29737 (N_29737,N_29178,N_29392);
or U29738 (N_29738,N_29334,N_29447);
and U29739 (N_29739,N_29221,N_29415);
or U29740 (N_29740,N_29104,N_29364);
and U29741 (N_29741,N_29160,N_29162);
and U29742 (N_29742,N_29093,N_29189);
or U29743 (N_29743,N_29192,N_29265);
nand U29744 (N_29744,N_29458,N_29087);
or U29745 (N_29745,N_29476,N_29450);
nand U29746 (N_29746,N_29430,N_29239);
and U29747 (N_29747,N_29384,N_29125);
and U29748 (N_29748,N_29083,N_29219);
nor U29749 (N_29749,N_29494,N_29252);
xnor U29750 (N_29750,N_29092,N_29057);
nand U29751 (N_29751,N_29250,N_29424);
nand U29752 (N_29752,N_29083,N_29084);
or U29753 (N_29753,N_29224,N_29389);
nand U29754 (N_29754,N_29110,N_29116);
or U29755 (N_29755,N_29369,N_29136);
or U29756 (N_29756,N_29325,N_29492);
nor U29757 (N_29757,N_29172,N_29334);
xnor U29758 (N_29758,N_29127,N_29457);
nor U29759 (N_29759,N_29458,N_29109);
xor U29760 (N_29760,N_29201,N_29427);
or U29761 (N_29761,N_29034,N_29379);
nor U29762 (N_29762,N_29419,N_29266);
nand U29763 (N_29763,N_29153,N_29141);
and U29764 (N_29764,N_29355,N_29338);
nand U29765 (N_29765,N_29490,N_29392);
or U29766 (N_29766,N_29095,N_29302);
nand U29767 (N_29767,N_29356,N_29241);
or U29768 (N_29768,N_29452,N_29394);
and U29769 (N_29769,N_29438,N_29117);
or U29770 (N_29770,N_29221,N_29175);
nor U29771 (N_29771,N_29031,N_29246);
xor U29772 (N_29772,N_29165,N_29173);
xor U29773 (N_29773,N_29199,N_29105);
nor U29774 (N_29774,N_29197,N_29078);
nand U29775 (N_29775,N_29327,N_29139);
xnor U29776 (N_29776,N_29457,N_29018);
xnor U29777 (N_29777,N_29271,N_29416);
nand U29778 (N_29778,N_29395,N_29471);
xnor U29779 (N_29779,N_29236,N_29165);
nand U29780 (N_29780,N_29103,N_29408);
xnor U29781 (N_29781,N_29318,N_29043);
xor U29782 (N_29782,N_29205,N_29456);
nand U29783 (N_29783,N_29251,N_29177);
nor U29784 (N_29784,N_29131,N_29015);
nor U29785 (N_29785,N_29001,N_29234);
and U29786 (N_29786,N_29145,N_29155);
or U29787 (N_29787,N_29024,N_29448);
nor U29788 (N_29788,N_29473,N_29287);
nand U29789 (N_29789,N_29412,N_29457);
and U29790 (N_29790,N_29363,N_29075);
or U29791 (N_29791,N_29206,N_29466);
or U29792 (N_29792,N_29499,N_29065);
or U29793 (N_29793,N_29040,N_29106);
nor U29794 (N_29794,N_29129,N_29056);
and U29795 (N_29795,N_29325,N_29266);
nor U29796 (N_29796,N_29309,N_29378);
xnor U29797 (N_29797,N_29399,N_29267);
nor U29798 (N_29798,N_29050,N_29287);
xor U29799 (N_29799,N_29465,N_29389);
nor U29800 (N_29800,N_29300,N_29045);
nor U29801 (N_29801,N_29226,N_29269);
nand U29802 (N_29802,N_29124,N_29076);
nor U29803 (N_29803,N_29036,N_29032);
nor U29804 (N_29804,N_29489,N_29486);
nand U29805 (N_29805,N_29440,N_29216);
nand U29806 (N_29806,N_29409,N_29226);
nor U29807 (N_29807,N_29385,N_29389);
nand U29808 (N_29808,N_29207,N_29132);
nand U29809 (N_29809,N_29072,N_29130);
nand U29810 (N_29810,N_29128,N_29349);
nand U29811 (N_29811,N_29301,N_29440);
and U29812 (N_29812,N_29105,N_29281);
nor U29813 (N_29813,N_29052,N_29126);
xnor U29814 (N_29814,N_29099,N_29027);
nor U29815 (N_29815,N_29304,N_29417);
nor U29816 (N_29816,N_29358,N_29357);
and U29817 (N_29817,N_29104,N_29387);
and U29818 (N_29818,N_29167,N_29098);
and U29819 (N_29819,N_29188,N_29300);
xnor U29820 (N_29820,N_29400,N_29493);
or U29821 (N_29821,N_29297,N_29050);
xor U29822 (N_29822,N_29146,N_29316);
nand U29823 (N_29823,N_29170,N_29142);
nand U29824 (N_29824,N_29385,N_29008);
and U29825 (N_29825,N_29438,N_29442);
nor U29826 (N_29826,N_29082,N_29422);
nand U29827 (N_29827,N_29151,N_29000);
nor U29828 (N_29828,N_29104,N_29368);
nand U29829 (N_29829,N_29412,N_29105);
or U29830 (N_29830,N_29268,N_29288);
nor U29831 (N_29831,N_29495,N_29205);
xor U29832 (N_29832,N_29426,N_29336);
or U29833 (N_29833,N_29318,N_29017);
xor U29834 (N_29834,N_29257,N_29066);
nand U29835 (N_29835,N_29018,N_29329);
or U29836 (N_29836,N_29378,N_29359);
nand U29837 (N_29837,N_29291,N_29048);
xnor U29838 (N_29838,N_29105,N_29331);
and U29839 (N_29839,N_29339,N_29403);
and U29840 (N_29840,N_29436,N_29362);
xnor U29841 (N_29841,N_29283,N_29138);
nand U29842 (N_29842,N_29348,N_29162);
xor U29843 (N_29843,N_29430,N_29484);
xnor U29844 (N_29844,N_29489,N_29455);
nand U29845 (N_29845,N_29178,N_29157);
nand U29846 (N_29846,N_29161,N_29395);
nor U29847 (N_29847,N_29202,N_29346);
nor U29848 (N_29848,N_29063,N_29104);
nor U29849 (N_29849,N_29309,N_29282);
nor U29850 (N_29850,N_29070,N_29343);
xnor U29851 (N_29851,N_29365,N_29486);
nand U29852 (N_29852,N_29171,N_29457);
nor U29853 (N_29853,N_29091,N_29238);
and U29854 (N_29854,N_29407,N_29045);
or U29855 (N_29855,N_29181,N_29174);
xor U29856 (N_29856,N_29189,N_29257);
or U29857 (N_29857,N_29320,N_29497);
nor U29858 (N_29858,N_29038,N_29326);
and U29859 (N_29859,N_29133,N_29007);
nor U29860 (N_29860,N_29472,N_29262);
xor U29861 (N_29861,N_29371,N_29352);
or U29862 (N_29862,N_29120,N_29404);
and U29863 (N_29863,N_29049,N_29279);
xor U29864 (N_29864,N_29175,N_29343);
nand U29865 (N_29865,N_29476,N_29121);
and U29866 (N_29866,N_29223,N_29314);
and U29867 (N_29867,N_29383,N_29307);
xor U29868 (N_29868,N_29499,N_29029);
or U29869 (N_29869,N_29226,N_29481);
nand U29870 (N_29870,N_29138,N_29115);
and U29871 (N_29871,N_29236,N_29192);
or U29872 (N_29872,N_29378,N_29194);
xnor U29873 (N_29873,N_29473,N_29127);
and U29874 (N_29874,N_29280,N_29192);
xor U29875 (N_29875,N_29471,N_29393);
or U29876 (N_29876,N_29289,N_29281);
nor U29877 (N_29877,N_29013,N_29316);
or U29878 (N_29878,N_29170,N_29322);
xnor U29879 (N_29879,N_29467,N_29493);
xnor U29880 (N_29880,N_29006,N_29017);
and U29881 (N_29881,N_29026,N_29136);
and U29882 (N_29882,N_29008,N_29102);
nor U29883 (N_29883,N_29018,N_29000);
xnor U29884 (N_29884,N_29160,N_29103);
nor U29885 (N_29885,N_29497,N_29034);
or U29886 (N_29886,N_29126,N_29425);
and U29887 (N_29887,N_29014,N_29237);
nand U29888 (N_29888,N_29265,N_29099);
nor U29889 (N_29889,N_29362,N_29486);
nor U29890 (N_29890,N_29308,N_29379);
nand U29891 (N_29891,N_29150,N_29086);
xnor U29892 (N_29892,N_29026,N_29347);
nand U29893 (N_29893,N_29447,N_29429);
xnor U29894 (N_29894,N_29190,N_29345);
or U29895 (N_29895,N_29451,N_29479);
xor U29896 (N_29896,N_29129,N_29132);
nor U29897 (N_29897,N_29238,N_29389);
nor U29898 (N_29898,N_29008,N_29334);
nor U29899 (N_29899,N_29456,N_29135);
nor U29900 (N_29900,N_29189,N_29032);
and U29901 (N_29901,N_29102,N_29454);
or U29902 (N_29902,N_29310,N_29370);
nand U29903 (N_29903,N_29412,N_29156);
nor U29904 (N_29904,N_29232,N_29132);
nor U29905 (N_29905,N_29103,N_29228);
xor U29906 (N_29906,N_29367,N_29248);
nand U29907 (N_29907,N_29119,N_29152);
xnor U29908 (N_29908,N_29358,N_29448);
and U29909 (N_29909,N_29489,N_29294);
nand U29910 (N_29910,N_29324,N_29100);
nor U29911 (N_29911,N_29399,N_29350);
or U29912 (N_29912,N_29251,N_29295);
xor U29913 (N_29913,N_29030,N_29083);
nand U29914 (N_29914,N_29196,N_29015);
nand U29915 (N_29915,N_29202,N_29195);
xor U29916 (N_29916,N_29161,N_29483);
xnor U29917 (N_29917,N_29264,N_29155);
xor U29918 (N_29918,N_29384,N_29286);
and U29919 (N_29919,N_29490,N_29359);
nor U29920 (N_29920,N_29460,N_29118);
and U29921 (N_29921,N_29369,N_29287);
xnor U29922 (N_29922,N_29041,N_29491);
or U29923 (N_29923,N_29461,N_29284);
nor U29924 (N_29924,N_29074,N_29085);
and U29925 (N_29925,N_29322,N_29090);
and U29926 (N_29926,N_29449,N_29318);
nor U29927 (N_29927,N_29395,N_29080);
or U29928 (N_29928,N_29258,N_29289);
nor U29929 (N_29929,N_29404,N_29340);
and U29930 (N_29930,N_29452,N_29126);
nor U29931 (N_29931,N_29450,N_29407);
nand U29932 (N_29932,N_29455,N_29072);
xnor U29933 (N_29933,N_29338,N_29474);
nand U29934 (N_29934,N_29318,N_29490);
and U29935 (N_29935,N_29261,N_29307);
and U29936 (N_29936,N_29273,N_29205);
nor U29937 (N_29937,N_29197,N_29178);
and U29938 (N_29938,N_29135,N_29345);
nor U29939 (N_29939,N_29268,N_29241);
nand U29940 (N_29940,N_29302,N_29371);
nand U29941 (N_29941,N_29130,N_29285);
xor U29942 (N_29942,N_29053,N_29487);
nor U29943 (N_29943,N_29154,N_29015);
xor U29944 (N_29944,N_29471,N_29157);
or U29945 (N_29945,N_29088,N_29209);
xor U29946 (N_29946,N_29170,N_29000);
nand U29947 (N_29947,N_29014,N_29146);
nand U29948 (N_29948,N_29478,N_29432);
nor U29949 (N_29949,N_29174,N_29430);
or U29950 (N_29950,N_29205,N_29336);
or U29951 (N_29951,N_29122,N_29019);
nor U29952 (N_29952,N_29133,N_29161);
or U29953 (N_29953,N_29120,N_29090);
and U29954 (N_29954,N_29076,N_29357);
xor U29955 (N_29955,N_29181,N_29185);
or U29956 (N_29956,N_29161,N_29384);
nor U29957 (N_29957,N_29107,N_29430);
nor U29958 (N_29958,N_29154,N_29031);
or U29959 (N_29959,N_29189,N_29415);
nand U29960 (N_29960,N_29481,N_29228);
and U29961 (N_29961,N_29056,N_29286);
nor U29962 (N_29962,N_29255,N_29196);
nand U29963 (N_29963,N_29416,N_29033);
and U29964 (N_29964,N_29473,N_29259);
and U29965 (N_29965,N_29085,N_29280);
or U29966 (N_29966,N_29285,N_29408);
nor U29967 (N_29967,N_29230,N_29316);
nor U29968 (N_29968,N_29385,N_29250);
nor U29969 (N_29969,N_29428,N_29113);
or U29970 (N_29970,N_29300,N_29323);
nor U29971 (N_29971,N_29255,N_29034);
or U29972 (N_29972,N_29100,N_29006);
xor U29973 (N_29973,N_29461,N_29270);
and U29974 (N_29974,N_29159,N_29290);
xnor U29975 (N_29975,N_29393,N_29383);
or U29976 (N_29976,N_29081,N_29043);
xnor U29977 (N_29977,N_29195,N_29156);
nor U29978 (N_29978,N_29034,N_29386);
or U29979 (N_29979,N_29001,N_29258);
nand U29980 (N_29980,N_29428,N_29332);
or U29981 (N_29981,N_29103,N_29392);
nor U29982 (N_29982,N_29496,N_29246);
xor U29983 (N_29983,N_29238,N_29421);
or U29984 (N_29984,N_29193,N_29016);
xor U29985 (N_29985,N_29000,N_29221);
nor U29986 (N_29986,N_29361,N_29205);
and U29987 (N_29987,N_29275,N_29383);
and U29988 (N_29988,N_29034,N_29212);
nor U29989 (N_29989,N_29355,N_29031);
nand U29990 (N_29990,N_29174,N_29441);
nor U29991 (N_29991,N_29024,N_29170);
or U29992 (N_29992,N_29091,N_29214);
nand U29993 (N_29993,N_29454,N_29217);
nor U29994 (N_29994,N_29219,N_29489);
nand U29995 (N_29995,N_29024,N_29219);
or U29996 (N_29996,N_29358,N_29195);
nand U29997 (N_29997,N_29122,N_29443);
and U29998 (N_29998,N_29175,N_29113);
nand U29999 (N_29999,N_29092,N_29036);
or U30000 (N_30000,N_29934,N_29686);
and U30001 (N_30001,N_29690,N_29779);
and U30002 (N_30002,N_29562,N_29748);
nor U30003 (N_30003,N_29694,N_29764);
nand U30004 (N_30004,N_29699,N_29814);
nand U30005 (N_30005,N_29731,N_29548);
nor U30006 (N_30006,N_29884,N_29727);
nor U30007 (N_30007,N_29831,N_29857);
or U30008 (N_30008,N_29914,N_29965);
nand U30009 (N_30009,N_29938,N_29796);
nor U30010 (N_30010,N_29642,N_29526);
nor U30011 (N_30011,N_29596,N_29618);
and U30012 (N_30012,N_29652,N_29542);
nor U30013 (N_30013,N_29787,N_29926);
xor U30014 (N_30014,N_29864,N_29841);
or U30015 (N_30015,N_29545,N_29718);
or U30016 (N_30016,N_29724,N_29658);
nor U30017 (N_30017,N_29912,N_29840);
and U30018 (N_30018,N_29681,N_29608);
xnor U30019 (N_30019,N_29619,N_29615);
or U30020 (N_30020,N_29881,N_29502);
nand U30021 (N_30021,N_29626,N_29676);
or U30022 (N_30022,N_29513,N_29993);
or U30023 (N_30023,N_29971,N_29709);
or U30024 (N_30024,N_29590,N_29827);
nor U30025 (N_30025,N_29917,N_29507);
nand U30026 (N_30026,N_29552,N_29722);
or U30027 (N_30027,N_29773,N_29544);
nand U30028 (N_30028,N_29999,N_29839);
or U30029 (N_30029,N_29792,N_29696);
nand U30030 (N_30030,N_29991,N_29786);
nand U30031 (N_30031,N_29894,N_29529);
nand U30032 (N_30032,N_29655,N_29768);
xnor U30033 (N_30033,N_29735,N_29711);
and U30034 (N_30034,N_29835,N_29714);
nor U30035 (N_30035,N_29911,N_29893);
xor U30036 (N_30036,N_29514,N_29720);
xor U30037 (N_30037,N_29698,N_29967);
nand U30038 (N_30038,N_29543,N_29747);
nand U30039 (N_30039,N_29879,N_29975);
nor U30040 (N_30040,N_29903,N_29907);
xor U30041 (N_30041,N_29826,N_29927);
and U30042 (N_30042,N_29920,N_29817);
and U30043 (N_30043,N_29848,N_29579);
and U30044 (N_30044,N_29828,N_29759);
or U30045 (N_30045,N_29612,N_29684);
nand U30046 (N_30046,N_29734,N_29789);
or U30047 (N_30047,N_29812,N_29795);
nand U30048 (N_30048,N_29610,N_29756);
and U30049 (N_30049,N_29508,N_29515);
nand U30050 (N_30050,N_29784,N_29942);
or U30051 (N_30051,N_29628,N_29974);
nor U30052 (N_30052,N_29892,N_29617);
xor U30053 (N_30053,N_29992,N_29749);
or U30054 (N_30054,N_29824,N_29976);
and U30055 (N_30055,N_29936,N_29876);
nor U30056 (N_30056,N_29646,N_29685);
or U30057 (N_30057,N_29743,N_29670);
nand U30058 (N_30058,N_29667,N_29570);
xnor U30059 (N_30059,N_29921,N_29822);
nor U30060 (N_30060,N_29559,N_29943);
and U30061 (N_30061,N_29950,N_29905);
nand U30062 (N_30062,N_29660,N_29973);
nor U30063 (N_30063,N_29739,N_29994);
xor U30064 (N_30064,N_29961,N_29834);
and U30065 (N_30065,N_29932,N_29772);
nor U30066 (N_30066,N_29598,N_29878);
nor U30067 (N_30067,N_29949,N_29541);
nand U30068 (N_30068,N_29673,N_29928);
and U30069 (N_30069,N_29808,N_29807);
nand U30070 (N_30070,N_29597,N_29557);
xnor U30071 (N_30071,N_29951,N_29862);
or U30072 (N_30072,N_29532,N_29611);
nand U30073 (N_30073,N_29679,N_29924);
nor U30074 (N_30074,N_29860,N_29777);
and U30075 (N_30075,N_29584,N_29701);
nor U30076 (N_30076,N_29955,N_29650);
nor U30077 (N_30077,N_29654,N_29675);
nand U30078 (N_30078,N_29763,N_29528);
and U30079 (N_30079,N_29517,N_29648);
nor U30080 (N_30080,N_29797,N_29908);
nand U30081 (N_30081,N_29639,N_29744);
and U30082 (N_30082,N_29604,N_29737);
and U30083 (N_30083,N_29916,N_29770);
nor U30084 (N_30084,N_29705,N_29762);
or U30085 (N_30085,N_29799,N_29621);
or U30086 (N_30086,N_29823,N_29883);
or U30087 (N_30087,N_29550,N_29554);
nand U30088 (N_30088,N_29940,N_29577);
and U30089 (N_30089,N_29910,N_29663);
or U30090 (N_30090,N_29697,N_29753);
nor U30091 (N_30091,N_29981,N_29668);
nand U30092 (N_30092,N_29540,N_29760);
xnor U30093 (N_30093,N_29865,N_29750);
and U30094 (N_30094,N_29637,N_29560);
nand U30095 (N_30095,N_29553,N_29820);
and U30096 (N_30096,N_29798,N_29630);
and U30097 (N_30097,N_29614,N_29632);
nor U30098 (N_30098,N_29555,N_29556);
nor U30099 (N_30099,N_29790,N_29585);
xor U30100 (N_30100,N_29861,N_29568);
nor U30101 (N_30101,N_29781,N_29998);
and U30102 (N_30102,N_29678,N_29656);
or U30103 (N_30103,N_29966,N_29674);
nor U30104 (N_30104,N_29946,N_29576);
and U30105 (N_30105,N_29886,N_29850);
nand U30106 (N_30106,N_29746,N_29672);
xor U30107 (N_30107,N_29623,N_29537);
xor U30108 (N_30108,N_29829,N_29740);
or U30109 (N_30109,N_29984,N_29855);
or U30110 (N_30110,N_29549,N_29671);
nor U30111 (N_30111,N_29713,N_29531);
xor U30112 (N_30112,N_29647,N_29653);
and U30113 (N_30113,N_29996,N_29700);
or U30114 (N_30114,N_29509,N_29870);
nand U30115 (N_30115,N_29519,N_29964);
or U30116 (N_30116,N_29906,N_29868);
and U30117 (N_30117,N_29578,N_29631);
and U30118 (N_30118,N_29582,N_29754);
and U30119 (N_30119,N_29919,N_29853);
nor U30120 (N_30120,N_29625,N_29521);
xnor U30121 (N_30121,N_29801,N_29904);
or U30122 (N_30122,N_29662,N_29702);
nand U30123 (N_30123,N_29980,N_29859);
nor U30124 (N_30124,N_29689,N_29547);
nor U30125 (N_30125,N_29669,N_29957);
xor U30126 (N_30126,N_29956,N_29869);
nand U30127 (N_30127,N_29771,N_29922);
xor U30128 (N_30128,N_29644,N_29846);
nand U30129 (N_30129,N_29988,N_29603);
xnor U30130 (N_30130,N_29539,N_29947);
nor U30131 (N_30131,N_29574,N_29536);
nand U30132 (N_30132,N_29638,N_29970);
or U30133 (N_30133,N_29629,N_29586);
or U30134 (N_30134,N_29791,N_29620);
or U30135 (N_30135,N_29587,N_29872);
xor U30136 (N_30136,N_29664,N_29983);
and U30137 (N_30137,N_29931,N_29538);
and U30138 (N_30138,N_29887,N_29504);
or U30139 (N_30139,N_29573,N_29783);
xor U30140 (N_30140,N_29794,N_29510);
nor U30141 (N_30141,N_29962,N_29785);
or U30142 (N_30142,N_29649,N_29982);
xor U30143 (N_30143,N_29845,N_29721);
nand U30144 (N_30144,N_29863,N_29852);
nand U30145 (N_30145,N_29506,N_29706);
nand U30146 (N_30146,N_29741,N_29571);
nand U30147 (N_30147,N_29851,N_29592);
xor U30148 (N_30148,N_29566,N_29635);
or U30149 (N_30149,N_29800,N_29751);
or U30150 (N_30150,N_29572,N_29583);
and U30151 (N_30151,N_29616,N_29503);
nor U30152 (N_30152,N_29890,N_29602);
xor U30153 (N_30153,N_29716,N_29821);
and U30154 (N_30154,N_29969,N_29843);
and U30155 (N_30155,N_29683,N_29809);
or U30156 (N_30156,N_29941,N_29937);
and U30157 (N_30157,N_29707,N_29935);
xnor U30158 (N_30158,N_29888,N_29929);
xor U30159 (N_30159,N_29987,N_29793);
xor U30160 (N_30160,N_29958,N_29645);
xnor U30161 (N_30161,N_29588,N_29703);
nor U30162 (N_30162,N_29640,N_29776);
nand U30163 (N_30163,N_29874,N_29591);
xnor U30164 (N_30164,N_29765,N_29715);
or U30165 (N_30165,N_29891,N_29803);
nor U30166 (N_30166,N_29682,N_29661);
or U30167 (N_30167,N_29522,N_29622);
or U30168 (N_30168,N_29717,N_29813);
xor U30169 (N_30169,N_29710,N_29636);
nand U30170 (N_30170,N_29923,N_29968);
and U30171 (N_30171,N_29516,N_29565);
nand U30172 (N_30172,N_29551,N_29815);
nor U30173 (N_30173,N_29500,N_29806);
xnor U30174 (N_30174,N_29534,N_29819);
and U30175 (N_30175,N_29844,N_29729);
nand U30176 (N_30176,N_29990,N_29595);
nand U30177 (N_30177,N_29708,N_29723);
and U30178 (N_30178,N_29527,N_29523);
xor U30179 (N_30179,N_29581,N_29594);
nor U30180 (N_30180,N_29624,N_29895);
nor U30181 (N_30181,N_29830,N_29774);
or U30182 (N_30182,N_29832,N_29691);
nand U30183 (N_30183,N_29899,N_29761);
and U30184 (N_30184,N_29885,N_29882);
and U30185 (N_30185,N_29818,N_29977);
nand U30186 (N_30186,N_29833,N_29877);
xor U30187 (N_30187,N_29858,N_29719);
and U30188 (N_30188,N_29897,N_29758);
xnor U30189 (N_30189,N_29902,N_29780);
nor U30190 (N_30190,N_29605,N_29634);
and U30191 (N_30191,N_29561,N_29520);
xor U30192 (N_30192,N_29567,N_29875);
nand U30193 (N_30193,N_29915,N_29778);
nor U30194 (N_30194,N_29930,N_29511);
and U30195 (N_30195,N_29738,N_29849);
xor U30196 (N_30196,N_29641,N_29680);
xor U30197 (N_30197,N_29802,N_29726);
and U30198 (N_30198,N_29704,N_29627);
and U30199 (N_30199,N_29898,N_29954);
nor U30200 (N_30200,N_29866,N_29530);
or U30201 (N_30201,N_29613,N_29742);
nor U30202 (N_30202,N_29525,N_29953);
nor U30203 (N_30203,N_29767,N_29816);
xnor U30204 (N_30204,N_29687,N_29952);
and U30205 (N_30205,N_29896,N_29788);
or U30206 (N_30206,N_29909,N_29593);
or U30207 (N_30207,N_29810,N_29728);
xor U30208 (N_30208,N_29838,N_29518);
nor U30209 (N_30209,N_29854,N_29979);
and U30210 (N_30210,N_29659,N_29918);
nor U30211 (N_30211,N_29871,N_29505);
xnor U30212 (N_30212,N_29733,N_29677);
nand U30213 (N_30213,N_29900,N_29643);
xor U30214 (N_30214,N_29535,N_29873);
or U30215 (N_30215,N_29825,N_29651);
xor U30216 (N_30216,N_29766,N_29558);
nand U30217 (N_30217,N_29805,N_29589);
nor U30218 (N_30218,N_29939,N_29995);
or U30219 (N_30219,N_29692,N_29836);
nand U30220 (N_30220,N_29599,N_29569);
or U30221 (N_30221,N_29901,N_29633);
nand U30222 (N_30222,N_29889,N_29501);
nand U30223 (N_30223,N_29782,N_29775);
and U30224 (N_30224,N_29725,N_29546);
nand U30225 (N_30225,N_29769,N_29847);
and U30226 (N_30226,N_29533,N_29512);
and U30227 (N_30227,N_29948,N_29732);
and U30228 (N_30228,N_29856,N_29804);
nor U30229 (N_30229,N_29842,N_29688);
and U30230 (N_30230,N_29867,N_29609);
or U30231 (N_30231,N_29986,N_29601);
or U30232 (N_30232,N_29564,N_29600);
xor U30233 (N_30233,N_29606,N_29752);
nor U30234 (N_30234,N_29693,N_29695);
and U30235 (N_30235,N_29665,N_29945);
xnor U30236 (N_30236,N_29607,N_29755);
nor U30237 (N_30237,N_29575,N_29580);
xor U30238 (N_30238,N_29563,N_29736);
nor U30239 (N_30239,N_29972,N_29933);
or U30240 (N_30240,N_29985,N_29978);
and U30241 (N_30241,N_29963,N_29757);
xnor U30242 (N_30242,N_29712,N_29960);
nor U30243 (N_30243,N_29837,N_29959);
nand U30244 (N_30244,N_29745,N_29811);
and U30245 (N_30245,N_29880,N_29730);
nand U30246 (N_30246,N_29913,N_29666);
nand U30247 (N_30247,N_29524,N_29989);
nor U30248 (N_30248,N_29944,N_29997);
or U30249 (N_30249,N_29657,N_29925);
and U30250 (N_30250,N_29502,N_29838);
nand U30251 (N_30251,N_29980,N_29636);
nand U30252 (N_30252,N_29743,N_29931);
nor U30253 (N_30253,N_29751,N_29513);
xor U30254 (N_30254,N_29896,N_29944);
nand U30255 (N_30255,N_29832,N_29557);
nor U30256 (N_30256,N_29574,N_29533);
nand U30257 (N_30257,N_29569,N_29584);
xnor U30258 (N_30258,N_29556,N_29742);
nand U30259 (N_30259,N_29545,N_29829);
nand U30260 (N_30260,N_29655,N_29943);
xor U30261 (N_30261,N_29720,N_29977);
or U30262 (N_30262,N_29748,N_29633);
xor U30263 (N_30263,N_29805,N_29709);
or U30264 (N_30264,N_29524,N_29981);
nand U30265 (N_30265,N_29731,N_29771);
xor U30266 (N_30266,N_29652,N_29867);
xnor U30267 (N_30267,N_29992,N_29559);
xnor U30268 (N_30268,N_29901,N_29871);
and U30269 (N_30269,N_29735,N_29644);
or U30270 (N_30270,N_29526,N_29782);
and U30271 (N_30271,N_29502,N_29523);
or U30272 (N_30272,N_29633,N_29519);
nor U30273 (N_30273,N_29542,N_29645);
nor U30274 (N_30274,N_29582,N_29727);
nand U30275 (N_30275,N_29602,N_29552);
nand U30276 (N_30276,N_29640,N_29843);
xor U30277 (N_30277,N_29719,N_29613);
and U30278 (N_30278,N_29779,N_29695);
nor U30279 (N_30279,N_29683,N_29824);
nor U30280 (N_30280,N_29979,N_29697);
nor U30281 (N_30281,N_29580,N_29761);
nand U30282 (N_30282,N_29661,N_29961);
xnor U30283 (N_30283,N_29622,N_29830);
xor U30284 (N_30284,N_29986,N_29613);
and U30285 (N_30285,N_29994,N_29737);
and U30286 (N_30286,N_29647,N_29881);
nand U30287 (N_30287,N_29856,N_29727);
or U30288 (N_30288,N_29951,N_29832);
and U30289 (N_30289,N_29971,N_29757);
xnor U30290 (N_30290,N_29739,N_29619);
xor U30291 (N_30291,N_29544,N_29906);
xor U30292 (N_30292,N_29963,N_29623);
nand U30293 (N_30293,N_29812,N_29952);
nor U30294 (N_30294,N_29893,N_29737);
xor U30295 (N_30295,N_29753,N_29778);
xor U30296 (N_30296,N_29986,N_29827);
nand U30297 (N_30297,N_29943,N_29680);
or U30298 (N_30298,N_29691,N_29593);
xnor U30299 (N_30299,N_29737,N_29862);
and U30300 (N_30300,N_29810,N_29665);
or U30301 (N_30301,N_29616,N_29634);
or U30302 (N_30302,N_29675,N_29502);
or U30303 (N_30303,N_29582,N_29862);
and U30304 (N_30304,N_29717,N_29771);
and U30305 (N_30305,N_29641,N_29905);
and U30306 (N_30306,N_29922,N_29677);
or U30307 (N_30307,N_29716,N_29844);
or U30308 (N_30308,N_29889,N_29838);
xnor U30309 (N_30309,N_29707,N_29550);
and U30310 (N_30310,N_29721,N_29778);
and U30311 (N_30311,N_29617,N_29934);
nor U30312 (N_30312,N_29718,N_29579);
or U30313 (N_30313,N_29621,N_29556);
nor U30314 (N_30314,N_29904,N_29626);
nand U30315 (N_30315,N_29843,N_29524);
or U30316 (N_30316,N_29738,N_29552);
nand U30317 (N_30317,N_29874,N_29853);
nand U30318 (N_30318,N_29651,N_29807);
xor U30319 (N_30319,N_29514,N_29731);
xnor U30320 (N_30320,N_29823,N_29975);
nand U30321 (N_30321,N_29645,N_29792);
xor U30322 (N_30322,N_29845,N_29596);
nand U30323 (N_30323,N_29946,N_29555);
nand U30324 (N_30324,N_29549,N_29832);
nor U30325 (N_30325,N_29514,N_29728);
nor U30326 (N_30326,N_29938,N_29898);
or U30327 (N_30327,N_29929,N_29678);
and U30328 (N_30328,N_29893,N_29575);
or U30329 (N_30329,N_29866,N_29783);
nor U30330 (N_30330,N_29594,N_29691);
nor U30331 (N_30331,N_29604,N_29868);
nand U30332 (N_30332,N_29982,N_29784);
or U30333 (N_30333,N_29840,N_29845);
or U30334 (N_30334,N_29791,N_29790);
nor U30335 (N_30335,N_29941,N_29830);
xnor U30336 (N_30336,N_29569,N_29712);
and U30337 (N_30337,N_29604,N_29698);
xor U30338 (N_30338,N_29577,N_29715);
xor U30339 (N_30339,N_29843,N_29732);
or U30340 (N_30340,N_29712,N_29889);
and U30341 (N_30341,N_29977,N_29880);
and U30342 (N_30342,N_29869,N_29617);
or U30343 (N_30343,N_29501,N_29914);
and U30344 (N_30344,N_29956,N_29690);
and U30345 (N_30345,N_29766,N_29525);
nand U30346 (N_30346,N_29732,N_29731);
nor U30347 (N_30347,N_29731,N_29821);
or U30348 (N_30348,N_29793,N_29975);
nor U30349 (N_30349,N_29678,N_29700);
xnor U30350 (N_30350,N_29654,N_29622);
or U30351 (N_30351,N_29756,N_29792);
nand U30352 (N_30352,N_29857,N_29950);
xnor U30353 (N_30353,N_29813,N_29686);
xor U30354 (N_30354,N_29825,N_29870);
xor U30355 (N_30355,N_29843,N_29673);
nor U30356 (N_30356,N_29975,N_29857);
or U30357 (N_30357,N_29588,N_29531);
xor U30358 (N_30358,N_29685,N_29949);
xor U30359 (N_30359,N_29871,N_29845);
nand U30360 (N_30360,N_29736,N_29858);
nor U30361 (N_30361,N_29774,N_29906);
nand U30362 (N_30362,N_29909,N_29791);
and U30363 (N_30363,N_29679,N_29648);
xor U30364 (N_30364,N_29662,N_29926);
nand U30365 (N_30365,N_29986,N_29971);
xnor U30366 (N_30366,N_29550,N_29598);
nand U30367 (N_30367,N_29887,N_29967);
xor U30368 (N_30368,N_29640,N_29966);
nor U30369 (N_30369,N_29838,N_29540);
nor U30370 (N_30370,N_29508,N_29688);
and U30371 (N_30371,N_29973,N_29732);
nand U30372 (N_30372,N_29581,N_29711);
or U30373 (N_30373,N_29835,N_29615);
and U30374 (N_30374,N_29863,N_29731);
and U30375 (N_30375,N_29729,N_29822);
nand U30376 (N_30376,N_29569,N_29994);
and U30377 (N_30377,N_29832,N_29856);
or U30378 (N_30378,N_29500,N_29697);
nand U30379 (N_30379,N_29914,N_29747);
or U30380 (N_30380,N_29669,N_29752);
xor U30381 (N_30381,N_29937,N_29734);
nor U30382 (N_30382,N_29508,N_29872);
or U30383 (N_30383,N_29658,N_29868);
nor U30384 (N_30384,N_29940,N_29589);
and U30385 (N_30385,N_29619,N_29730);
or U30386 (N_30386,N_29994,N_29628);
xor U30387 (N_30387,N_29949,N_29937);
xor U30388 (N_30388,N_29571,N_29748);
xor U30389 (N_30389,N_29730,N_29749);
and U30390 (N_30390,N_29846,N_29909);
nand U30391 (N_30391,N_29757,N_29506);
and U30392 (N_30392,N_29712,N_29522);
and U30393 (N_30393,N_29926,N_29684);
and U30394 (N_30394,N_29778,N_29702);
nor U30395 (N_30395,N_29906,N_29814);
xnor U30396 (N_30396,N_29737,N_29787);
or U30397 (N_30397,N_29809,N_29651);
or U30398 (N_30398,N_29519,N_29851);
and U30399 (N_30399,N_29903,N_29975);
nand U30400 (N_30400,N_29762,N_29934);
nor U30401 (N_30401,N_29663,N_29940);
and U30402 (N_30402,N_29758,N_29707);
and U30403 (N_30403,N_29765,N_29535);
xnor U30404 (N_30404,N_29505,N_29512);
nand U30405 (N_30405,N_29618,N_29686);
and U30406 (N_30406,N_29668,N_29720);
nand U30407 (N_30407,N_29758,N_29927);
xor U30408 (N_30408,N_29995,N_29905);
or U30409 (N_30409,N_29532,N_29830);
and U30410 (N_30410,N_29876,N_29725);
nand U30411 (N_30411,N_29558,N_29701);
xnor U30412 (N_30412,N_29886,N_29985);
or U30413 (N_30413,N_29755,N_29818);
nand U30414 (N_30414,N_29813,N_29924);
nor U30415 (N_30415,N_29930,N_29862);
or U30416 (N_30416,N_29614,N_29587);
or U30417 (N_30417,N_29577,N_29731);
and U30418 (N_30418,N_29539,N_29985);
or U30419 (N_30419,N_29953,N_29526);
nor U30420 (N_30420,N_29969,N_29797);
or U30421 (N_30421,N_29667,N_29946);
or U30422 (N_30422,N_29856,N_29686);
nor U30423 (N_30423,N_29993,N_29871);
nand U30424 (N_30424,N_29983,N_29530);
or U30425 (N_30425,N_29768,N_29769);
and U30426 (N_30426,N_29768,N_29843);
xnor U30427 (N_30427,N_29789,N_29836);
nor U30428 (N_30428,N_29574,N_29964);
nand U30429 (N_30429,N_29789,N_29684);
or U30430 (N_30430,N_29623,N_29575);
or U30431 (N_30431,N_29851,N_29973);
nor U30432 (N_30432,N_29750,N_29909);
or U30433 (N_30433,N_29577,N_29820);
nor U30434 (N_30434,N_29671,N_29543);
xor U30435 (N_30435,N_29892,N_29965);
or U30436 (N_30436,N_29742,N_29894);
or U30437 (N_30437,N_29500,N_29673);
nor U30438 (N_30438,N_29673,N_29984);
xnor U30439 (N_30439,N_29892,N_29563);
and U30440 (N_30440,N_29959,N_29816);
nand U30441 (N_30441,N_29735,N_29879);
or U30442 (N_30442,N_29895,N_29609);
nand U30443 (N_30443,N_29824,N_29599);
nand U30444 (N_30444,N_29894,N_29648);
or U30445 (N_30445,N_29743,N_29731);
or U30446 (N_30446,N_29757,N_29987);
and U30447 (N_30447,N_29772,N_29664);
or U30448 (N_30448,N_29921,N_29664);
or U30449 (N_30449,N_29748,N_29614);
and U30450 (N_30450,N_29574,N_29683);
nor U30451 (N_30451,N_29563,N_29859);
nor U30452 (N_30452,N_29753,N_29973);
nor U30453 (N_30453,N_29954,N_29682);
or U30454 (N_30454,N_29656,N_29584);
and U30455 (N_30455,N_29935,N_29898);
or U30456 (N_30456,N_29584,N_29967);
nor U30457 (N_30457,N_29669,N_29845);
nand U30458 (N_30458,N_29904,N_29625);
and U30459 (N_30459,N_29915,N_29523);
nor U30460 (N_30460,N_29934,N_29837);
or U30461 (N_30461,N_29553,N_29952);
and U30462 (N_30462,N_29910,N_29879);
or U30463 (N_30463,N_29935,N_29982);
xor U30464 (N_30464,N_29843,N_29678);
xor U30465 (N_30465,N_29964,N_29730);
nor U30466 (N_30466,N_29957,N_29564);
or U30467 (N_30467,N_29792,N_29692);
or U30468 (N_30468,N_29585,N_29720);
and U30469 (N_30469,N_29804,N_29732);
nor U30470 (N_30470,N_29606,N_29506);
xor U30471 (N_30471,N_29853,N_29721);
xor U30472 (N_30472,N_29705,N_29985);
nor U30473 (N_30473,N_29984,N_29572);
nor U30474 (N_30474,N_29546,N_29794);
nand U30475 (N_30475,N_29910,N_29927);
and U30476 (N_30476,N_29520,N_29804);
xor U30477 (N_30477,N_29594,N_29576);
or U30478 (N_30478,N_29909,N_29866);
nand U30479 (N_30479,N_29820,N_29543);
or U30480 (N_30480,N_29968,N_29883);
nor U30481 (N_30481,N_29799,N_29903);
xnor U30482 (N_30482,N_29548,N_29555);
and U30483 (N_30483,N_29965,N_29863);
and U30484 (N_30484,N_29989,N_29946);
xnor U30485 (N_30485,N_29679,N_29795);
and U30486 (N_30486,N_29721,N_29695);
nor U30487 (N_30487,N_29607,N_29516);
or U30488 (N_30488,N_29995,N_29935);
nor U30489 (N_30489,N_29840,N_29673);
nand U30490 (N_30490,N_29853,N_29697);
nor U30491 (N_30491,N_29823,N_29782);
or U30492 (N_30492,N_29827,N_29771);
nor U30493 (N_30493,N_29545,N_29577);
nor U30494 (N_30494,N_29903,N_29653);
nand U30495 (N_30495,N_29502,N_29527);
xor U30496 (N_30496,N_29937,N_29728);
and U30497 (N_30497,N_29902,N_29502);
nand U30498 (N_30498,N_29930,N_29736);
nor U30499 (N_30499,N_29985,N_29989);
xnor U30500 (N_30500,N_30311,N_30404);
xor U30501 (N_30501,N_30450,N_30273);
xnor U30502 (N_30502,N_30353,N_30030);
or U30503 (N_30503,N_30033,N_30021);
or U30504 (N_30504,N_30206,N_30207);
and U30505 (N_30505,N_30413,N_30122);
or U30506 (N_30506,N_30189,N_30484);
or U30507 (N_30507,N_30110,N_30326);
nand U30508 (N_30508,N_30173,N_30023);
nand U30509 (N_30509,N_30071,N_30348);
nor U30510 (N_30510,N_30383,N_30292);
xor U30511 (N_30511,N_30460,N_30330);
or U30512 (N_30512,N_30366,N_30352);
and U30513 (N_30513,N_30014,N_30410);
nand U30514 (N_30514,N_30176,N_30082);
nand U30515 (N_30515,N_30276,N_30487);
or U30516 (N_30516,N_30191,N_30194);
or U30517 (N_30517,N_30163,N_30328);
nand U30518 (N_30518,N_30049,N_30092);
nand U30519 (N_30519,N_30474,N_30496);
xor U30520 (N_30520,N_30057,N_30318);
nor U30521 (N_30521,N_30284,N_30001);
or U30522 (N_30522,N_30044,N_30397);
or U30523 (N_30523,N_30103,N_30462);
or U30524 (N_30524,N_30425,N_30391);
and U30525 (N_30525,N_30296,N_30249);
nand U30526 (N_30526,N_30188,N_30196);
nand U30527 (N_30527,N_30275,N_30497);
xor U30528 (N_30528,N_30400,N_30406);
or U30529 (N_30529,N_30153,N_30038);
nand U30530 (N_30530,N_30449,N_30234);
or U30531 (N_30531,N_30323,N_30140);
or U30532 (N_30532,N_30079,N_30369);
nand U30533 (N_30533,N_30152,N_30015);
nand U30534 (N_30534,N_30494,N_30375);
nand U30535 (N_30535,N_30333,N_30144);
and U30536 (N_30536,N_30319,N_30068);
or U30537 (N_30537,N_30136,N_30228);
nand U30538 (N_30538,N_30016,N_30309);
nor U30539 (N_30539,N_30371,N_30358);
xor U30540 (N_30540,N_30491,N_30244);
nor U30541 (N_30541,N_30059,N_30324);
nor U30542 (N_30542,N_30133,N_30210);
or U30543 (N_30543,N_30243,N_30029);
xnor U30544 (N_30544,N_30213,N_30368);
nand U30545 (N_30545,N_30139,N_30004);
xor U30546 (N_30546,N_30074,N_30009);
and U30547 (N_30547,N_30350,N_30005);
nand U30548 (N_30548,N_30265,N_30047);
nor U30549 (N_30549,N_30347,N_30089);
xnor U30550 (N_30550,N_30381,N_30087);
or U30551 (N_30551,N_30086,N_30080);
and U30552 (N_30552,N_30149,N_30422);
xnor U30553 (N_30553,N_30257,N_30385);
xor U30554 (N_30554,N_30286,N_30129);
and U30555 (N_30555,N_30433,N_30409);
and U30556 (N_30556,N_30058,N_30392);
nand U30557 (N_30557,N_30499,N_30253);
and U30558 (N_30558,N_30341,N_30125);
nand U30559 (N_30559,N_30203,N_30126);
nor U30560 (N_30560,N_30495,N_30430);
or U30561 (N_30561,N_30380,N_30488);
and U30562 (N_30562,N_30280,N_30441);
or U30563 (N_30563,N_30221,N_30022);
and U30564 (N_30564,N_30003,N_30388);
xor U30565 (N_30565,N_30442,N_30008);
xor U30566 (N_30566,N_30032,N_30470);
or U30567 (N_30567,N_30377,N_30469);
xor U30568 (N_30568,N_30455,N_30065);
xnor U30569 (N_30569,N_30272,N_30060);
and U30570 (N_30570,N_30131,N_30482);
xnor U30571 (N_30571,N_30055,N_30012);
nand U30572 (N_30572,N_30112,N_30130);
and U30573 (N_30573,N_30317,N_30236);
nor U30574 (N_30574,N_30332,N_30048);
or U30575 (N_30575,N_30454,N_30389);
nand U30576 (N_30576,N_30204,N_30419);
nand U30577 (N_30577,N_30473,N_30282);
nand U30578 (N_30578,N_30148,N_30277);
xor U30579 (N_30579,N_30436,N_30002);
nand U30580 (N_30580,N_30100,N_30370);
nor U30581 (N_30581,N_30471,N_30254);
xnor U30582 (N_30582,N_30091,N_30486);
nor U30583 (N_30583,N_30235,N_30289);
and U30584 (N_30584,N_30160,N_30039);
or U30585 (N_30585,N_30246,N_30359);
nor U30586 (N_30586,N_30094,N_30155);
xnor U30587 (N_30587,N_30020,N_30314);
or U30588 (N_30588,N_30117,N_30424);
xnor U30589 (N_30589,N_30360,N_30240);
nand U30590 (N_30590,N_30143,N_30156);
or U30591 (N_30591,N_30171,N_30438);
xor U30592 (N_30592,N_30135,N_30159);
xnor U30593 (N_30593,N_30031,N_30172);
nor U30594 (N_30594,N_30247,N_30107);
nor U30595 (N_30595,N_30411,N_30342);
and U30596 (N_30596,N_30301,N_30337);
or U30597 (N_30597,N_30361,N_30278);
xnor U30598 (N_30598,N_30492,N_30354);
nand U30599 (N_30599,N_30017,N_30335);
xnor U30600 (N_30600,N_30298,N_30428);
nand U30601 (N_30601,N_30320,N_30043);
nor U30602 (N_30602,N_30439,N_30150);
nor U30603 (N_30603,N_30472,N_30480);
xor U30604 (N_30604,N_30034,N_30387);
or U30605 (N_30605,N_30024,N_30054);
or U30606 (N_30606,N_30279,N_30415);
and U30607 (N_30607,N_30281,N_30248);
or U30608 (N_30608,N_30013,N_30000);
and U30609 (N_30609,N_30178,N_30040);
nand U30610 (N_30610,N_30170,N_30215);
and U30611 (N_30611,N_30429,N_30050);
and U30612 (N_30612,N_30251,N_30205);
nor U30613 (N_30613,N_30175,N_30127);
and U30614 (N_30614,N_30432,N_30417);
nand U30615 (N_30615,N_30211,N_30293);
nand U30616 (N_30616,N_30336,N_30099);
nor U30617 (N_30617,N_30157,N_30443);
xor U30618 (N_30618,N_30457,N_30198);
nand U30619 (N_30619,N_30459,N_30230);
nor U30620 (N_30620,N_30476,N_30343);
nand U30621 (N_30621,N_30197,N_30313);
and U30622 (N_30622,N_30180,N_30285);
or U30623 (N_30623,N_30200,N_30104);
nand U30624 (N_30624,N_30372,N_30097);
and U30625 (N_30625,N_30090,N_30229);
nor U30626 (N_30626,N_30075,N_30305);
or U30627 (N_30627,N_30418,N_30339);
xor U30628 (N_30628,N_30056,N_30042);
and U30629 (N_30629,N_30493,N_30187);
nand U30630 (N_30630,N_30481,N_30477);
xnor U30631 (N_30631,N_30378,N_30299);
or U30632 (N_30632,N_30303,N_30220);
nand U30633 (N_30633,N_30349,N_30158);
and U30634 (N_30634,N_30363,N_30224);
nand U30635 (N_30635,N_30283,N_30255);
and U30636 (N_30636,N_30209,N_30475);
xnor U30637 (N_30637,N_30331,N_30468);
xnor U30638 (N_30638,N_30109,N_30183);
and U30639 (N_30639,N_30052,N_30241);
nand U30640 (N_30640,N_30452,N_30498);
nand U30641 (N_30641,N_30174,N_30365);
nand U30642 (N_30642,N_30227,N_30165);
nand U30643 (N_30643,N_30291,N_30357);
nor U30644 (N_30644,N_30238,N_30288);
and U30645 (N_30645,N_30062,N_30485);
nand U30646 (N_30646,N_30169,N_30222);
xnor U30647 (N_30647,N_30269,N_30111);
xor U30648 (N_30648,N_30223,N_30447);
nand U30649 (N_30649,N_30390,N_30212);
xor U30650 (N_30650,N_30088,N_30344);
nand U30651 (N_30651,N_30268,N_30479);
xor U30652 (N_30652,N_30258,N_30321);
nand U30653 (N_30653,N_30458,N_30478);
or U30654 (N_30654,N_30412,N_30408);
nor U30655 (N_30655,N_30217,N_30426);
and U30656 (N_30656,N_30019,N_30340);
nor U30657 (N_30657,N_30367,N_30010);
nand U30658 (N_30658,N_30297,N_30154);
and U30659 (N_30659,N_30451,N_30067);
or U30660 (N_30660,N_30446,N_30300);
or U30661 (N_30661,N_30434,N_30164);
and U30662 (N_30662,N_30242,N_30270);
and U30663 (N_30663,N_30114,N_30219);
nor U30664 (N_30664,N_30376,N_30036);
and U30665 (N_30665,N_30081,N_30395);
or U30666 (N_30666,N_30064,N_30128);
nand U30667 (N_30667,N_30355,N_30078);
xnor U30668 (N_30668,N_30231,N_30440);
and U30669 (N_30669,N_30134,N_30306);
or U30670 (N_30670,N_30098,N_30201);
nand U30671 (N_30671,N_30051,N_30066);
xor U30672 (N_30672,N_30364,N_30083);
xor U30673 (N_30673,N_30076,N_30421);
or U30674 (N_30674,N_30394,N_30489);
xor U30675 (N_30675,N_30199,N_30063);
nand U30676 (N_30676,N_30261,N_30445);
xnor U30677 (N_30677,N_30307,N_30167);
nand U30678 (N_30678,N_30399,N_30162);
and U30679 (N_30679,N_30356,N_30184);
and U30680 (N_30680,N_30264,N_30035);
nand U30681 (N_30681,N_30374,N_30262);
and U30682 (N_30682,N_30322,N_30393);
nor U30683 (N_30683,N_30302,N_30113);
and U30684 (N_30684,N_30329,N_30232);
nand U30685 (N_30685,N_30453,N_30093);
nor U30686 (N_30686,N_30414,N_30138);
and U30687 (N_30687,N_30026,N_30456);
nor U30688 (N_30688,N_30105,N_30386);
xnor U30689 (N_30689,N_30463,N_30084);
nor U30690 (N_30690,N_30037,N_30345);
nor U30691 (N_30691,N_30402,N_30327);
nor U30692 (N_30692,N_30085,N_30006);
or U30693 (N_30693,N_30202,N_30310);
nand U30694 (N_30694,N_30216,N_30007);
nand U30695 (N_30695,N_30053,N_30028);
nand U30696 (N_30696,N_30151,N_30259);
or U30697 (N_30697,N_30142,N_30226);
and U30698 (N_30698,N_30123,N_30192);
or U30699 (N_30699,N_30308,N_30132);
nor U30700 (N_30700,N_30405,N_30315);
nand U30701 (N_30701,N_30466,N_30362);
nor U30702 (N_30702,N_30271,N_30018);
nor U30703 (N_30703,N_30250,N_30423);
xor U30704 (N_30704,N_30420,N_30137);
xor U30705 (N_30705,N_30218,N_30483);
nand U30706 (N_30706,N_30403,N_30373);
nand U30707 (N_30707,N_30069,N_30168);
nor U30708 (N_30708,N_30116,N_30185);
and U30709 (N_30709,N_30045,N_30225);
or U30710 (N_30710,N_30011,N_30338);
nor U30711 (N_30711,N_30252,N_30431);
nand U30712 (N_30712,N_30181,N_30435);
or U30713 (N_30713,N_30193,N_30077);
nor U30714 (N_30714,N_30190,N_30464);
or U30715 (N_30715,N_30334,N_30427);
xor U30716 (N_30716,N_30263,N_30401);
xor U30717 (N_30717,N_30095,N_30108);
nand U30718 (N_30718,N_30312,N_30437);
or U30719 (N_30719,N_30416,N_30237);
and U30720 (N_30720,N_30396,N_30115);
nand U30721 (N_30721,N_30448,N_30179);
or U30722 (N_30722,N_30384,N_30146);
nand U30723 (N_30723,N_30120,N_30316);
or U30724 (N_30724,N_30072,N_30145);
nand U30725 (N_30725,N_30186,N_30274);
xor U30726 (N_30726,N_30398,N_30325);
nor U30727 (N_30727,N_30027,N_30304);
xnor U30728 (N_30728,N_30267,N_30096);
or U30729 (N_30729,N_30256,N_30287);
nor U30730 (N_30730,N_30106,N_30177);
and U30731 (N_30731,N_30260,N_30046);
or U30732 (N_30732,N_30266,N_30195);
xor U30733 (N_30733,N_30346,N_30245);
nand U30734 (N_30734,N_30166,N_30124);
xor U30735 (N_30735,N_30467,N_30407);
nand U30736 (N_30736,N_30118,N_30461);
nand U30737 (N_30737,N_30295,N_30025);
nand U30738 (N_30738,N_30208,N_30290);
xnor U30739 (N_30739,N_30161,N_30182);
and U30740 (N_30740,N_30121,N_30490);
or U30741 (N_30741,N_30101,N_30351);
nand U30742 (N_30742,N_30294,N_30233);
nor U30743 (N_30743,N_30214,N_30239);
or U30744 (N_30744,N_30465,N_30379);
xor U30745 (N_30745,N_30061,N_30070);
nor U30746 (N_30746,N_30119,N_30444);
xor U30747 (N_30747,N_30147,N_30141);
and U30748 (N_30748,N_30102,N_30382);
nand U30749 (N_30749,N_30073,N_30041);
or U30750 (N_30750,N_30452,N_30085);
or U30751 (N_30751,N_30231,N_30463);
and U30752 (N_30752,N_30145,N_30352);
xor U30753 (N_30753,N_30423,N_30251);
nor U30754 (N_30754,N_30292,N_30333);
and U30755 (N_30755,N_30441,N_30428);
nor U30756 (N_30756,N_30291,N_30404);
nor U30757 (N_30757,N_30057,N_30083);
nand U30758 (N_30758,N_30009,N_30061);
xor U30759 (N_30759,N_30115,N_30342);
or U30760 (N_30760,N_30374,N_30205);
nand U30761 (N_30761,N_30482,N_30165);
nor U30762 (N_30762,N_30222,N_30178);
or U30763 (N_30763,N_30227,N_30351);
xor U30764 (N_30764,N_30277,N_30373);
xnor U30765 (N_30765,N_30170,N_30053);
xnor U30766 (N_30766,N_30098,N_30023);
or U30767 (N_30767,N_30283,N_30329);
or U30768 (N_30768,N_30163,N_30380);
xnor U30769 (N_30769,N_30381,N_30063);
xnor U30770 (N_30770,N_30319,N_30081);
nor U30771 (N_30771,N_30416,N_30029);
xor U30772 (N_30772,N_30300,N_30427);
nand U30773 (N_30773,N_30295,N_30405);
xor U30774 (N_30774,N_30195,N_30261);
nor U30775 (N_30775,N_30146,N_30308);
nor U30776 (N_30776,N_30011,N_30411);
nand U30777 (N_30777,N_30499,N_30213);
nand U30778 (N_30778,N_30427,N_30171);
nor U30779 (N_30779,N_30018,N_30119);
or U30780 (N_30780,N_30027,N_30111);
nand U30781 (N_30781,N_30389,N_30059);
xor U30782 (N_30782,N_30282,N_30407);
xor U30783 (N_30783,N_30481,N_30116);
and U30784 (N_30784,N_30114,N_30266);
xnor U30785 (N_30785,N_30421,N_30190);
xnor U30786 (N_30786,N_30233,N_30353);
xor U30787 (N_30787,N_30248,N_30454);
and U30788 (N_30788,N_30305,N_30404);
xnor U30789 (N_30789,N_30315,N_30040);
xnor U30790 (N_30790,N_30023,N_30078);
nand U30791 (N_30791,N_30085,N_30009);
and U30792 (N_30792,N_30236,N_30367);
nand U30793 (N_30793,N_30137,N_30243);
or U30794 (N_30794,N_30348,N_30065);
xor U30795 (N_30795,N_30262,N_30354);
nand U30796 (N_30796,N_30416,N_30476);
nand U30797 (N_30797,N_30004,N_30421);
xnor U30798 (N_30798,N_30048,N_30098);
xnor U30799 (N_30799,N_30059,N_30021);
nand U30800 (N_30800,N_30479,N_30201);
and U30801 (N_30801,N_30125,N_30447);
or U30802 (N_30802,N_30336,N_30317);
xor U30803 (N_30803,N_30209,N_30486);
nand U30804 (N_30804,N_30066,N_30118);
and U30805 (N_30805,N_30048,N_30246);
nor U30806 (N_30806,N_30297,N_30453);
and U30807 (N_30807,N_30241,N_30071);
or U30808 (N_30808,N_30494,N_30404);
nand U30809 (N_30809,N_30281,N_30211);
xor U30810 (N_30810,N_30262,N_30290);
xnor U30811 (N_30811,N_30121,N_30164);
or U30812 (N_30812,N_30210,N_30231);
nor U30813 (N_30813,N_30025,N_30197);
nor U30814 (N_30814,N_30130,N_30429);
nor U30815 (N_30815,N_30324,N_30366);
nand U30816 (N_30816,N_30194,N_30285);
nand U30817 (N_30817,N_30050,N_30448);
nand U30818 (N_30818,N_30172,N_30192);
xnor U30819 (N_30819,N_30190,N_30325);
nand U30820 (N_30820,N_30213,N_30357);
and U30821 (N_30821,N_30243,N_30394);
xor U30822 (N_30822,N_30034,N_30358);
nor U30823 (N_30823,N_30455,N_30386);
xnor U30824 (N_30824,N_30028,N_30151);
nor U30825 (N_30825,N_30421,N_30337);
or U30826 (N_30826,N_30451,N_30488);
xnor U30827 (N_30827,N_30224,N_30222);
and U30828 (N_30828,N_30478,N_30111);
and U30829 (N_30829,N_30044,N_30383);
or U30830 (N_30830,N_30431,N_30065);
nand U30831 (N_30831,N_30005,N_30091);
xnor U30832 (N_30832,N_30239,N_30243);
nand U30833 (N_30833,N_30305,N_30332);
and U30834 (N_30834,N_30111,N_30098);
nand U30835 (N_30835,N_30253,N_30099);
nor U30836 (N_30836,N_30032,N_30371);
nor U30837 (N_30837,N_30376,N_30256);
nor U30838 (N_30838,N_30140,N_30237);
or U30839 (N_30839,N_30379,N_30194);
and U30840 (N_30840,N_30363,N_30407);
or U30841 (N_30841,N_30483,N_30458);
nand U30842 (N_30842,N_30432,N_30407);
nor U30843 (N_30843,N_30139,N_30422);
nor U30844 (N_30844,N_30045,N_30011);
and U30845 (N_30845,N_30126,N_30070);
nor U30846 (N_30846,N_30246,N_30291);
nor U30847 (N_30847,N_30216,N_30444);
xnor U30848 (N_30848,N_30028,N_30465);
and U30849 (N_30849,N_30192,N_30433);
or U30850 (N_30850,N_30044,N_30412);
and U30851 (N_30851,N_30202,N_30245);
and U30852 (N_30852,N_30318,N_30345);
xnor U30853 (N_30853,N_30205,N_30273);
and U30854 (N_30854,N_30264,N_30214);
xor U30855 (N_30855,N_30396,N_30180);
nor U30856 (N_30856,N_30495,N_30463);
or U30857 (N_30857,N_30142,N_30184);
or U30858 (N_30858,N_30190,N_30214);
and U30859 (N_30859,N_30379,N_30200);
nand U30860 (N_30860,N_30336,N_30129);
or U30861 (N_30861,N_30046,N_30018);
nor U30862 (N_30862,N_30102,N_30329);
nor U30863 (N_30863,N_30199,N_30374);
or U30864 (N_30864,N_30499,N_30401);
nand U30865 (N_30865,N_30227,N_30196);
and U30866 (N_30866,N_30410,N_30421);
nor U30867 (N_30867,N_30460,N_30204);
or U30868 (N_30868,N_30200,N_30384);
nand U30869 (N_30869,N_30218,N_30279);
nor U30870 (N_30870,N_30483,N_30479);
nand U30871 (N_30871,N_30159,N_30050);
xnor U30872 (N_30872,N_30031,N_30415);
nand U30873 (N_30873,N_30149,N_30427);
nand U30874 (N_30874,N_30093,N_30116);
or U30875 (N_30875,N_30246,N_30311);
nor U30876 (N_30876,N_30428,N_30123);
nand U30877 (N_30877,N_30162,N_30350);
nor U30878 (N_30878,N_30414,N_30289);
xnor U30879 (N_30879,N_30494,N_30170);
or U30880 (N_30880,N_30253,N_30033);
or U30881 (N_30881,N_30164,N_30194);
xor U30882 (N_30882,N_30210,N_30238);
nand U30883 (N_30883,N_30428,N_30430);
nand U30884 (N_30884,N_30320,N_30247);
or U30885 (N_30885,N_30126,N_30338);
nor U30886 (N_30886,N_30405,N_30234);
nor U30887 (N_30887,N_30482,N_30309);
or U30888 (N_30888,N_30437,N_30092);
or U30889 (N_30889,N_30454,N_30052);
and U30890 (N_30890,N_30398,N_30488);
nand U30891 (N_30891,N_30296,N_30122);
nor U30892 (N_30892,N_30031,N_30334);
xnor U30893 (N_30893,N_30166,N_30255);
and U30894 (N_30894,N_30491,N_30052);
and U30895 (N_30895,N_30419,N_30066);
or U30896 (N_30896,N_30425,N_30395);
nor U30897 (N_30897,N_30376,N_30367);
nand U30898 (N_30898,N_30456,N_30314);
and U30899 (N_30899,N_30032,N_30401);
and U30900 (N_30900,N_30081,N_30364);
nor U30901 (N_30901,N_30228,N_30180);
xor U30902 (N_30902,N_30371,N_30140);
xor U30903 (N_30903,N_30246,N_30118);
nor U30904 (N_30904,N_30256,N_30115);
and U30905 (N_30905,N_30258,N_30201);
and U30906 (N_30906,N_30272,N_30339);
and U30907 (N_30907,N_30116,N_30001);
or U30908 (N_30908,N_30182,N_30011);
nor U30909 (N_30909,N_30008,N_30131);
and U30910 (N_30910,N_30328,N_30198);
or U30911 (N_30911,N_30204,N_30467);
nand U30912 (N_30912,N_30006,N_30224);
or U30913 (N_30913,N_30132,N_30171);
and U30914 (N_30914,N_30316,N_30065);
nand U30915 (N_30915,N_30043,N_30388);
nand U30916 (N_30916,N_30402,N_30426);
nand U30917 (N_30917,N_30116,N_30266);
nand U30918 (N_30918,N_30205,N_30066);
and U30919 (N_30919,N_30244,N_30175);
nand U30920 (N_30920,N_30396,N_30083);
or U30921 (N_30921,N_30456,N_30422);
and U30922 (N_30922,N_30102,N_30420);
nand U30923 (N_30923,N_30420,N_30311);
and U30924 (N_30924,N_30045,N_30035);
or U30925 (N_30925,N_30430,N_30291);
and U30926 (N_30926,N_30454,N_30243);
or U30927 (N_30927,N_30056,N_30104);
or U30928 (N_30928,N_30103,N_30302);
xor U30929 (N_30929,N_30018,N_30042);
or U30930 (N_30930,N_30064,N_30437);
nand U30931 (N_30931,N_30345,N_30177);
nand U30932 (N_30932,N_30205,N_30270);
nand U30933 (N_30933,N_30454,N_30478);
xnor U30934 (N_30934,N_30218,N_30167);
and U30935 (N_30935,N_30480,N_30400);
nor U30936 (N_30936,N_30028,N_30459);
nor U30937 (N_30937,N_30305,N_30059);
nor U30938 (N_30938,N_30140,N_30401);
or U30939 (N_30939,N_30132,N_30183);
and U30940 (N_30940,N_30266,N_30193);
nor U30941 (N_30941,N_30359,N_30473);
nor U30942 (N_30942,N_30271,N_30255);
nor U30943 (N_30943,N_30099,N_30318);
nand U30944 (N_30944,N_30487,N_30144);
xor U30945 (N_30945,N_30070,N_30405);
nor U30946 (N_30946,N_30341,N_30074);
xnor U30947 (N_30947,N_30431,N_30420);
or U30948 (N_30948,N_30455,N_30003);
or U30949 (N_30949,N_30108,N_30489);
nand U30950 (N_30950,N_30177,N_30360);
nand U30951 (N_30951,N_30370,N_30472);
xor U30952 (N_30952,N_30161,N_30388);
xnor U30953 (N_30953,N_30088,N_30228);
or U30954 (N_30954,N_30364,N_30308);
xor U30955 (N_30955,N_30494,N_30155);
nand U30956 (N_30956,N_30307,N_30331);
xnor U30957 (N_30957,N_30428,N_30338);
nand U30958 (N_30958,N_30137,N_30337);
or U30959 (N_30959,N_30091,N_30351);
or U30960 (N_30960,N_30259,N_30136);
nand U30961 (N_30961,N_30049,N_30412);
nor U30962 (N_30962,N_30136,N_30256);
or U30963 (N_30963,N_30007,N_30142);
and U30964 (N_30964,N_30414,N_30244);
or U30965 (N_30965,N_30358,N_30289);
and U30966 (N_30966,N_30007,N_30176);
nor U30967 (N_30967,N_30047,N_30353);
xor U30968 (N_30968,N_30059,N_30245);
nor U30969 (N_30969,N_30133,N_30448);
xnor U30970 (N_30970,N_30185,N_30396);
or U30971 (N_30971,N_30002,N_30310);
and U30972 (N_30972,N_30077,N_30155);
or U30973 (N_30973,N_30098,N_30047);
xnor U30974 (N_30974,N_30357,N_30024);
nand U30975 (N_30975,N_30356,N_30140);
nor U30976 (N_30976,N_30053,N_30034);
nand U30977 (N_30977,N_30024,N_30111);
or U30978 (N_30978,N_30073,N_30210);
nor U30979 (N_30979,N_30248,N_30488);
or U30980 (N_30980,N_30012,N_30437);
xor U30981 (N_30981,N_30165,N_30323);
or U30982 (N_30982,N_30481,N_30170);
nand U30983 (N_30983,N_30266,N_30112);
or U30984 (N_30984,N_30374,N_30383);
or U30985 (N_30985,N_30043,N_30095);
or U30986 (N_30986,N_30066,N_30106);
and U30987 (N_30987,N_30235,N_30299);
and U30988 (N_30988,N_30310,N_30318);
nor U30989 (N_30989,N_30054,N_30343);
or U30990 (N_30990,N_30100,N_30372);
or U30991 (N_30991,N_30348,N_30130);
xnor U30992 (N_30992,N_30461,N_30268);
or U30993 (N_30993,N_30415,N_30026);
xnor U30994 (N_30994,N_30185,N_30449);
nand U30995 (N_30995,N_30315,N_30388);
and U30996 (N_30996,N_30467,N_30278);
or U30997 (N_30997,N_30051,N_30411);
nand U30998 (N_30998,N_30496,N_30297);
xor U30999 (N_30999,N_30252,N_30434);
and U31000 (N_31000,N_30766,N_30661);
or U31001 (N_31001,N_30991,N_30648);
and U31002 (N_31002,N_30935,N_30973);
nor U31003 (N_31003,N_30794,N_30587);
xor U31004 (N_31004,N_30781,N_30831);
nor U31005 (N_31005,N_30940,N_30590);
nand U31006 (N_31006,N_30697,N_30721);
or U31007 (N_31007,N_30681,N_30562);
or U31008 (N_31008,N_30568,N_30628);
xnor U31009 (N_31009,N_30775,N_30949);
xor U31010 (N_31010,N_30879,N_30951);
nor U31011 (N_31011,N_30680,N_30572);
or U31012 (N_31012,N_30863,N_30688);
and U31013 (N_31013,N_30578,N_30886);
or U31014 (N_31014,N_30666,N_30872);
or U31015 (N_31015,N_30686,N_30848);
xor U31016 (N_31016,N_30986,N_30868);
nor U31017 (N_31017,N_30747,N_30647);
and U31018 (N_31018,N_30699,N_30771);
nor U31019 (N_31019,N_30984,N_30751);
or U31020 (N_31020,N_30873,N_30615);
nand U31021 (N_31021,N_30535,N_30663);
nor U31022 (N_31022,N_30600,N_30575);
and U31023 (N_31023,N_30961,N_30825);
nor U31024 (N_31024,N_30630,N_30948);
or U31025 (N_31025,N_30701,N_30854);
or U31026 (N_31026,N_30524,N_30905);
xnor U31027 (N_31027,N_30977,N_30560);
or U31028 (N_31028,N_30542,N_30705);
nor U31029 (N_31029,N_30621,N_30637);
xor U31030 (N_31030,N_30574,N_30588);
or U31031 (N_31031,N_30727,N_30510);
nand U31032 (N_31032,N_30728,N_30513);
xnor U31033 (N_31033,N_30815,N_30658);
and U31034 (N_31034,N_30833,N_30812);
nand U31035 (N_31035,N_30683,N_30599);
and U31036 (N_31036,N_30618,N_30625);
nor U31037 (N_31037,N_30953,N_30736);
nor U31038 (N_31038,N_30821,N_30520);
and U31039 (N_31039,N_30678,N_30537);
nand U31040 (N_31040,N_30500,N_30957);
nor U31041 (N_31041,N_30938,N_30822);
xnor U31042 (N_31042,N_30906,N_30884);
nand U31043 (N_31043,N_30774,N_30853);
nand U31044 (N_31044,N_30911,N_30920);
nand U31045 (N_31045,N_30507,N_30895);
or U31046 (N_31046,N_30690,N_30960);
nor U31047 (N_31047,N_30750,N_30836);
and U31048 (N_31048,N_30577,N_30778);
nor U31049 (N_31049,N_30937,N_30689);
nor U31050 (N_31050,N_30692,N_30871);
xor U31051 (N_31051,N_30823,N_30660);
and U31052 (N_31052,N_30622,N_30624);
or U31053 (N_31053,N_30877,N_30931);
and U31054 (N_31054,N_30784,N_30936);
nor U31055 (N_31055,N_30662,N_30546);
and U31056 (N_31056,N_30726,N_30737);
xor U31057 (N_31057,N_30502,N_30539);
nand U31058 (N_31058,N_30764,N_30912);
nand U31059 (N_31059,N_30805,N_30841);
and U31060 (N_31060,N_30890,N_30566);
nor U31061 (N_31061,N_30965,N_30824);
and U31062 (N_31062,N_30846,N_30548);
or U31063 (N_31063,N_30640,N_30670);
nand U31064 (N_31064,N_30734,N_30564);
and U31065 (N_31065,N_30544,N_30753);
and U31066 (N_31066,N_30684,N_30643);
or U31067 (N_31067,N_30682,N_30667);
and U31068 (N_31068,N_30765,N_30669);
and U31069 (N_31069,N_30729,N_30858);
nor U31070 (N_31070,N_30988,N_30844);
nor U31071 (N_31071,N_30857,N_30547);
nand U31072 (N_31072,N_30992,N_30915);
or U31073 (N_31073,N_30767,N_30768);
xnor U31074 (N_31074,N_30816,N_30707);
nor U31075 (N_31075,N_30907,N_30832);
nor U31076 (N_31076,N_30793,N_30741);
or U31077 (N_31077,N_30800,N_30894);
nand U31078 (N_31078,N_30655,N_30749);
and U31079 (N_31079,N_30693,N_30602);
or U31080 (N_31080,N_30995,N_30806);
or U31081 (N_31081,N_30540,N_30555);
nor U31082 (N_31082,N_30604,N_30807);
xnor U31083 (N_31083,N_30606,N_30503);
or U31084 (N_31084,N_30875,N_30712);
and U31085 (N_31085,N_30665,N_30819);
xor U31086 (N_31086,N_30515,N_30934);
nor U31087 (N_31087,N_30921,N_30659);
nor U31088 (N_31088,N_30631,N_30717);
nand U31089 (N_31089,N_30942,N_30526);
nor U31090 (N_31090,N_30830,N_30508);
nor U31091 (N_31091,N_30976,N_30842);
and U31092 (N_31092,N_30914,N_30829);
and U31093 (N_31093,N_30870,N_30709);
nor U31094 (N_31094,N_30633,N_30714);
or U31095 (N_31095,N_30731,N_30855);
or U31096 (N_31096,N_30786,N_30592);
nand U31097 (N_31097,N_30964,N_30797);
or U31098 (N_31098,N_30638,N_30799);
nand U31099 (N_31099,N_30760,N_30913);
nand U31100 (N_31100,N_30791,N_30878);
or U31101 (N_31101,N_30543,N_30856);
nor U31102 (N_31102,N_30748,N_30803);
xnor U31103 (N_31103,N_30598,N_30571);
xnor U31104 (N_31104,N_30685,N_30967);
nor U31105 (N_31105,N_30504,N_30770);
xor U31106 (N_31106,N_30773,N_30772);
or U31107 (N_31107,N_30755,N_30917);
and U31108 (N_31108,N_30552,N_30835);
xor U31109 (N_31109,N_30601,N_30763);
xnor U31110 (N_31110,N_30530,N_30757);
nor U31111 (N_31111,N_30888,N_30919);
and U31112 (N_31112,N_30677,N_30759);
nor U31113 (N_31113,N_30541,N_30527);
nor U31114 (N_31114,N_30927,N_30987);
or U31115 (N_31115,N_30523,N_30933);
or U31116 (N_31116,N_30533,N_30923);
xor U31117 (N_31117,N_30881,N_30996);
nand U31118 (N_31118,N_30516,N_30865);
and U31119 (N_31119,N_30723,N_30597);
nand U31120 (N_31120,N_30904,N_30512);
nor U31121 (N_31121,N_30522,N_30596);
and U31122 (N_31122,N_30897,N_30792);
and U31123 (N_31123,N_30710,N_30534);
and U31124 (N_31124,N_30549,N_30553);
and U31125 (N_31125,N_30837,N_30946);
nand U31126 (N_31126,N_30673,N_30580);
xor U31127 (N_31127,N_30635,N_30817);
nor U31128 (N_31128,N_30617,N_30713);
and U31129 (N_31129,N_30595,N_30645);
nand U31130 (N_31130,N_30605,N_30758);
nand U31131 (N_31131,N_30959,N_30980);
nand U31132 (N_31132,N_30565,N_30899);
and U31133 (N_31133,N_30943,N_30963);
nand U31134 (N_31134,N_30909,N_30656);
or U31135 (N_31135,N_30834,N_30525);
nor U31136 (N_31136,N_30880,N_30809);
xor U31137 (N_31137,N_30889,N_30804);
nand U31138 (N_31138,N_30898,N_30627);
or U31139 (N_31139,N_30779,N_30859);
or U31140 (N_31140,N_30743,N_30756);
and U31141 (N_31141,N_30876,N_30982);
xor U31142 (N_31142,N_30573,N_30557);
xor U31143 (N_31143,N_30783,N_30653);
nand U31144 (N_31144,N_30703,N_30589);
nor U31145 (N_31145,N_30514,N_30827);
nand U31146 (N_31146,N_30929,N_30582);
nand U31147 (N_31147,N_30702,N_30867);
nor U31148 (N_31148,N_30509,N_30966);
nand U31149 (N_31149,N_30752,N_30972);
nor U31150 (N_31150,N_30922,N_30561);
nand U31151 (N_31151,N_30896,N_30820);
nand U31152 (N_31152,N_30607,N_30994);
xnor U31153 (N_31153,N_30802,N_30704);
xor U31154 (N_31154,N_30594,N_30744);
xnor U31155 (N_31155,N_30567,N_30671);
and U31156 (N_31156,N_30900,N_30970);
or U31157 (N_31157,N_30808,N_30614);
or U31158 (N_31158,N_30796,N_30777);
and U31159 (N_31159,N_30769,N_30887);
nor U31160 (N_31160,N_30950,N_30719);
xnor U31161 (N_31161,N_30551,N_30883);
nor U31162 (N_31162,N_30939,N_30696);
and U31163 (N_31163,N_30910,N_30732);
xnor U31164 (N_31164,N_30646,N_30538);
or U31165 (N_31165,N_30616,N_30612);
or U31166 (N_31166,N_30593,N_30828);
xnor U31167 (N_31167,N_30716,N_30990);
and U31168 (N_31168,N_30978,N_30632);
xor U31169 (N_31169,N_30885,N_30785);
and U31170 (N_31170,N_30609,N_30787);
nor U31171 (N_31171,N_30956,N_30583);
and U31172 (N_31172,N_30981,N_30619);
xnor U31173 (N_31173,N_30708,N_30695);
nor U31174 (N_31174,N_30584,N_30613);
and U31175 (N_31175,N_30652,N_30722);
and U31176 (N_31176,N_30916,N_30558);
or U31177 (N_31177,N_30556,N_30698);
nor U31178 (N_31178,N_30818,N_30790);
or U31179 (N_31179,N_30864,N_30610);
xor U31180 (N_31180,N_30813,N_30810);
or U31181 (N_31181,N_30754,N_30947);
xnor U31182 (N_31182,N_30672,N_30968);
nor U31183 (N_31183,N_30634,N_30739);
nor U31184 (N_31184,N_30985,N_30691);
xnor U31185 (N_31185,N_30891,N_30675);
or U31186 (N_31186,N_30706,N_30962);
xor U31187 (N_31187,N_30862,N_30814);
nand U31188 (N_31188,N_30811,N_30517);
nor U31189 (N_31189,N_30711,N_30776);
xor U31190 (N_31190,N_30901,N_30735);
nor U31191 (N_31191,N_30679,N_30528);
xor U31192 (N_31192,N_30840,N_30851);
and U31193 (N_31193,N_30536,N_30839);
and U31194 (N_31194,N_30559,N_30518);
and U31195 (N_31195,N_30586,N_30789);
nand U31196 (N_31196,N_30563,N_30850);
xnor U31197 (N_31197,N_30849,N_30958);
nand U31198 (N_31198,N_30893,N_30866);
nand U31199 (N_31199,N_30993,N_30997);
xnor U31200 (N_31200,N_30826,N_30932);
nand U31201 (N_31201,N_30843,N_30782);
xnor U31202 (N_31202,N_30801,N_30974);
nand U31203 (N_31203,N_30852,N_30550);
nand U31204 (N_31204,N_30944,N_30644);
xnor U31205 (N_31205,N_30746,N_30642);
xnor U31206 (N_31206,N_30989,N_30576);
and U31207 (N_31207,N_30745,N_30925);
nor U31208 (N_31208,N_30845,N_30569);
xnor U31209 (N_31209,N_30969,N_30952);
nand U31210 (N_31210,N_30506,N_30724);
nand U31211 (N_31211,N_30725,N_30694);
and U31212 (N_31212,N_30676,N_30579);
xnor U31213 (N_31213,N_30718,N_30521);
and U31214 (N_31214,N_30611,N_30545);
nor U31215 (N_31215,N_30674,N_30955);
nor U31216 (N_31216,N_30532,N_30930);
or U31217 (N_31217,N_30519,N_30908);
and U31218 (N_31218,N_30668,N_30874);
nand U31219 (N_31219,N_30636,N_30798);
nor U31220 (N_31220,N_30623,N_30738);
nand U31221 (N_31221,N_30975,N_30626);
or U31222 (N_31222,N_30861,N_30650);
nand U31223 (N_31223,N_30715,N_30902);
and U31224 (N_31224,N_30740,N_30945);
nand U31225 (N_31225,N_30654,N_30570);
xnor U31226 (N_31226,N_30581,N_30511);
nand U31227 (N_31227,N_30999,N_30591);
xnor U31228 (N_31228,N_30869,N_30838);
or U31229 (N_31229,N_30603,N_30687);
or U31230 (N_31230,N_30928,N_30585);
xnor U31231 (N_31231,N_30926,N_30941);
and U31232 (N_31232,N_30795,N_30882);
nor U31233 (N_31233,N_30529,N_30554);
nor U31234 (N_31234,N_30629,N_30860);
or U31235 (N_31235,N_30664,N_30720);
nand U31236 (N_31236,N_30971,N_30761);
xnor U31237 (N_31237,N_30847,N_30918);
and U31238 (N_31238,N_30979,N_30700);
and U31239 (N_31239,N_30780,N_30651);
nand U31240 (N_31240,N_30892,N_30903);
nand U31241 (N_31241,N_30730,N_30733);
nor U31242 (N_31242,N_30762,N_30924);
xnor U31243 (N_31243,N_30531,N_30505);
nand U31244 (N_31244,N_30998,N_30983);
or U31245 (N_31245,N_30641,N_30954);
and U31246 (N_31246,N_30649,N_30657);
or U31247 (N_31247,N_30639,N_30620);
or U31248 (N_31248,N_30742,N_30501);
and U31249 (N_31249,N_30788,N_30608);
or U31250 (N_31250,N_30933,N_30689);
nor U31251 (N_31251,N_30967,N_30973);
nand U31252 (N_31252,N_30833,N_30596);
xnor U31253 (N_31253,N_30980,N_30577);
xor U31254 (N_31254,N_30769,N_30807);
and U31255 (N_31255,N_30996,N_30800);
xnor U31256 (N_31256,N_30552,N_30798);
xnor U31257 (N_31257,N_30722,N_30587);
xor U31258 (N_31258,N_30655,N_30698);
xor U31259 (N_31259,N_30673,N_30697);
or U31260 (N_31260,N_30850,N_30651);
or U31261 (N_31261,N_30974,N_30750);
or U31262 (N_31262,N_30731,N_30858);
nand U31263 (N_31263,N_30508,N_30667);
nand U31264 (N_31264,N_30951,N_30859);
or U31265 (N_31265,N_30857,N_30701);
and U31266 (N_31266,N_30695,N_30624);
nor U31267 (N_31267,N_30824,N_30834);
nor U31268 (N_31268,N_30802,N_30721);
nor U31269 (N_31269,N_30920,N_30829);
xor U31270 (N_31270,N_30689,N_30870);
nor U31271 (N_31271,N_30565,N_30555);
nor U31272 (N_31272,N_30576,N_30962);
or U31273 (N_31273,N_30529,N_30505);
and U31274 (N_31274,N_30686,N_30633);
or U31275 (N_31275,N_30825,N_30881);
and U31276 (N_31276,N_30805,N_30759);
or U31277 (N_31277,N_30664,N_30911);
xnor U31278 (N_31278,N_30789,N_30507);
nand U31279 (N_31279,N_30729,N_30860);
nand U31280 (N_31280,N_30677,N_30988);
xor U31281 (N_31281,N_30682,N_30732);
and U31282 (N_31282,N_30903,N_30823);
nand U31283 (N_31283,N_30886,N_30611);
or U31284 (N_31284,N_30892,N_30967);
nor U31285 (N_31285,N_30931,N_30746);
xnor U31286 (N_31286,N_30685,N_30993);
nand U31287 (N_31287,N_30817,N_30946);
nand U31288 (N_31288,N_30787,N_30670);
or U31289 (N_31289,N_30799,N_30663);
or U31290 (N_31290,N_30845,N_30657);
nand U31291 (N_31291,N_30531,N_30976);
or U31292 (N_31292,N_30688,N_30508);
and U31293 (N_31293,N_30538,N_30847);
nand U31294 (N_31294,N_30504,N_30883);
or U31295 (N_31295,N_30649,N_30832);
nor U31296 (N_31296,N_30652,N_30574);
xor U31297 (N_31297,N_30659,N_30608);
and U31298 (N_31298,N_30628,N_30712);
and U31299 (N_31299,N_30719,N_30850);
nand U31300 (N_31300,N_30533,N_30714);
nor U31301 (N_31301,N_30808,N_30708);
xor U31302 (N_31302,N_30976,N_30505);
nand U31303 (N_31303,N_30516,N_30849);
nor U31304 (N_31304,N_30534,N_30830);
nand U31305 (N_31305,N_30805,N_30997);
xnor U31306 (N_31306,N_30741,N_30805);
xnor U31307 (N_31307,N_30524,N_30507);
and U31308 (N_31308,N_30742,N_30730);
nand U31309 (N_31309,N_30972,N_30714);
nor U31310 (N_31310,N_30965,N_30603);
nand U31311 (N_31311,N_30737,N_30697);
nor U31312 (N_31312,N_30606,N_30551);
xor U31313 (N_31313,N_30674,N_30722);
and U31314 (N_31314,N_30540,N_30744);
nand U31315 (N_31315,N_30594,N_30526);
nor U31316 (N_31316,N_30762,N_30868);
and U31317 (N_31317,N_30945,N_30586);
nor U31318 (N_31318,N_30769,N_30970);
xor U31319 (N_31319,N_30952,N_30673);
nor U31320 (N_31320,N_30912,N_30560);
or U31321 (N_31321,N_30878,N_30637);
nand U31322 (N_31322,N_30562,N_30726);
and U31323 (N_31323,N_30699,N_30726);
nor U31324 (N_31324,N_30929,N_30732);
nor U31325 (N_31325,N_30870,N_30794);
or U31326 (N_31326,N_30819,N_30778);
and U31327 (N_31327,N_30646,N_30521);
or U31328 (N_31328,N_30993,N_30751);
nand U31329 (N_31329,N_30728,N_30892);
and U31330 (N_31330,N_30921,N_30692);
xor U31331 (N_31331,N_30707,N_30985);
nand U31332 (N_31332,N_30547,N_30992);
or U31333 (N_31333,N_30686,N_30566);
or U31334 (N_31334,N_30813,N_30960);
or U31335 (N_31335,N_30627,N_30996);
nor U31336 (N_31336,N_30631,N_30635);
and U31337 (N_31337,N_30759,N_30685);
and U31338 (N_31338,N_30651,N_30783);
and U31339 (N_31339,N_30690,N_30863);
nand U31340 (N_31340,N_30953,N_30756);
and U31341 (N_31341,N_30608,N_30688);
nand U31342 (N_31342,N_30640,N_30579);
or U31343 (N_31343,N_30977,N_30879);
and U31344 (N_31344,N_30558,N_30949);
xnor U31345 (N_31345,N_30942,N_30930);
xor U31346 (N_31346,N_30904,N_30570);
xor U31347 (N_31347,N_30592,N_30513);
or U31348 (N_31348,N_30940,N_30974);
nand U31349 (N_31349,N_30729,N_30529);
nand U31350 (N_31350,N_30612,N_30711);
and U31351 (N_31351,N_30656,N_30825);
nor U31352 (N_31352,N_30760,N_30563);
nand U31353 (N_31353,N_30576,N_30947);
or U31354 (N_31354,N_30575,N_30653);
and U31355 (N_31355,N_30688,N_30606);
or U31356 (N_31356,N_30679,N_30862);
xnor U31357 (N_31357,N_30719,N_30595);
or U31358 (N_31358,N_30955,N_30526);
or U31359 (N_31359,N_30526,N_30545);
and U31360 (N_31360,N_30817,N_30653);
nor U31361 (N_31361,N_30507,N_30936);
nand U31362 (N_31362,N_30859,N_30892);
or U31363 (N_31363,N_30953,N_30987);
or U31364 (N_31364,N_30865,N_30788);
xor U31365 (N_31365,N_30987,N_30550);
or U31366 (N_31366,N_30602,N_30769);
nor U31367 (N_31367,N_30767,N_30660);
or U31368 (N_31368,N_30660,N_30609);
or U31369 (N_31369,N_30776,N_30832);
xor U31370 (N_31370,N_30661,N_30635);
nor U31371 (N_31371,N_30604,N_30865);
or U31372 (N_31372,N_30923,N_30878);
or U31373 (N_31373,N_30567,N_30865);
or U31374 (N_31374,N_30642,N_30767);
and U31375 (N_31375,N_30886,N_30553);
xnor U31376 (N_31376,N_30553,N_30934);
and U31377 (N_31377,N_30520,N_30835);
nor U31378 (N_31378,N_30526,N_30988);
nand U31379 (N_31379,N_30740,N_30715);
or U31380 (N_31380,N_30558,N_30684);
and U31381 (N_31381,N_30937,N_30539);
or U31382 (N_31382,N_30880,N_30710);
nor U31383 (N_31383,N_30979,N_30774);
and U31384 (N_31384,N_30738,N_30773);
and U31385 (N_31385,N_30602,N_30767);
or U31386 (N_31386,N_30859,N_30746);
xor U31387 (N_31387,N_30513,N_30666);
nor U31388 (N_31388,N_30600,N_30733);
nor U31389 (N_31389,N_30883,N_30533);
xnor U31390 (N_31390,N_30521,N_30911);
nor U31391 (N_31391,N_30658,N_30617);
xnor U31392 (N_31392,N_30896,N_30990);
nor U31393 (N_31393,N_30984,N_30938);
or U31394 (N_31394,N_30943,N_30974);
nor U31395 (N_31395,N_30871,N_30810);
or U31396 (N_31396,N_30789,N_30757);
and U31397 (N_31397,N_30978,N_30982);
or U31398 (N_31398,N_30824,N_30997);
nor U31399 (N_31399,N_30667,N_30769);
and U31400 (N_31400,N_30959,N_30783);
or U31401 (N_31401,N_30815,N_30918);
xnor U31402 (N_31402,N_30655,N_30602);
xnor U31403 (N_31403,N_30790,N_30572);
or U31404 (N_31404,N_30595,N_30684);
or U31405 (N_31405,N_30710,N_30690);
and U31406 (N_31406,N_30925,N_30693);
and U31407 (N_31407,N_30750,N_30630);
or U31408 (N_31408,N_30706,N_30719);
nand U31409 (N_31409,N_30825,N_30592);
and U31410 (N_31410,N_30636,N_30806);
and U31411 (N_31411,N_30569,N_30567);
and U31412 (N_31412,N_30679,N_30958);
nand U31413 (N_31413,N_30777,N_30577);
xor U31414 (N_31414,N_30923,N_30867);
nor U31415 (N_31415,N_30920,N_30755);
xor U31416 (N_31416,N_30790,N_30934);
nor U31417 (N_31417,N_30667,N_30920);
or U31418 (N_31418,N_30670,N_30825);
xnor U31419 (N_31419,N_30578,N_30810);
xnor U31420 (N_31420,N_30690,N_30936);
nor U31421 (N_31421,N_30518,N_30505);
xnor U31422 (N_31422,N_30606,N_30884);
nor U31423 (N_31423,N_30520,N_30525);
nand U31424 (N_31424,N_30943,N_30580);
nand U31425 (N_31425,N_30931,N_30736);
xor U31426 (N_31426,N_30681,N_30759);
xor U31427 (N_31427,N_30761,N_30767);
nor U31428 (N_31428,N_30716,N_30859);
or U31429 (N_31429,N_30758,N_30676);
nor U31430 (N_31430,N_30874,N_30860);
and U31431 (N_31431,N_30939,N_30631);
and U31432 (N_31432,N_30931,N_30637);
or U31433 (N_31433,N_30608,N_30922);
xnor U31434 (N_31434,N_30832,N_30506);
nor U31435 (N_31435,N_30796,N_30518);
nor U31436 (N_31436,N_30944,N_30776);
nand U31437 (N_31437,N_30703,N_30845);
nor U31438 (N_31438,N_30531,N_30812);
nand U31439 (N_31439,N_30985,N_30870);
nand U31440 (N_31440,N_30855,N_30554);
xnor U31441 (N_31441,N_30619,N_30904);
and U31442 (N_31442,N_30876,N_30649);
nor U31443 (N_31443,N_30731,N_30533);
or U31444 (N_31444,N_30800,N_30712);
and U31445 (N_31445,N_30753,N_30794);
xnor U31446 (N_31446,N_30735,N_30751);
nor U31447 (N_31447,N_30998,N_30718);
and U31448 (N_31448,N_30633,N_30705);
or U31449 (N_31449,N_30931,N_30733);
and U31450 (N_31450,N_30694,N_30563);
xnor U31451 (N_31451,N_30621,N_30726);
nor U31452 (N_31452,N_30692,N_30654);
xnor U31453 (N_31453,N_30969,N_30548);
or U31454 (N_31454,N_30955,N_30721);
xnor U31455 (N_31455,N_30917,N_30611);
xor U31456 (N_31456,N_30811,N_30966);
xnor U31457 (N_31457,N_30916,N_30880);
nand U31458 (N_31458,N_30683,N_30525);
or U31459 (N_31459,N_30848,N_30862);
nor U31460 (N_31460,N_30723,N_30570);
and U31461 (N_31461,N_30571,N_30871);
nand U31462 (N_31462,N_30856,N_30622);
xor U31463 (N_31463,N_30979,N_30659);
xnor U31464 (N_31464,N_30633,N_30609);
or U31465 (N_31465,N_30830,N_30737);
or U31466 (N_31466,N_30826,N_30588);
nand U31467 (N_31467,N_30992,N_30832);
xnor U31468 (N_31468,N_30816,N_30735);
xnor U31469 (N_31469,N_30838,N_30629);
nand U31470 (N_31470,N_30674,N_30773);
nor U31471 (N_31471,N_30564,N_30981);
xor U31472 (N_31472,N_30682,N_30871);
and U31473 (N_31473,N_30650,N_30799);
nand U31474 (N_31474,N_30593,N_30797);
xor U31475 (N_31475,N_30557,N_30506);
and U31476 (N_31476,N_30745,N_30853);
xnor U31477 (N_31477,N_30872,N_30878);
or U31478 (N_31478,N_30612,N_30783);
nor U31479 (N_31479,N_30980,N_30708);
and U31480 (N_31480,N_30617,N_30967);
nand U31481 (N_31481,N_30760,N_30564);
nor U31482 (N_31482,N_30821,N_30501);
nor U31483 (N_31483,N_30848,N_30913);
nor U31484 (N_31484,N_30515,N_30501);
nand U31485 (N_31485,N_30802,N_30531);
xor U31486 (N_31486,N_30927,N_30990);
nor U31487 (N_31487,N_30910,N_30985);
nand U31488 (N_31488,N_30592,N_30594);
and U31489 (N_31489,N_30695,N_30893);
xnor U31490 (N_31490,N_30926,N_30583);
and U31491 (N_31491,N_30784,N_30526);
nand U31492 (N_31492,N_30824,N_30808);
and U31493 (N_31493,N_30825,N_30737);
or U31494 (N_31494,N_30542,N_30832);
nand U31495 (N_31495,N_30655,N_30859);
and U31496 (N_31496,N_30954,N_30672);
and U31497 (N_31497,N_30847,N_30919);
nand U31498 (N_31498,N_30831,N_30717);
nand U31499 (N_31499,N_30898,N_30510);
or U31500 (N_31500,N_31060,N_31337);
nand U31501 (N_31501,N_31411,N_31353);
nand U31502 (N_31502,N_31229,N_31447);
or U31503 (N_31503,N_31101,N_31231);
or U31504 (N_31504,N_31368,N_31429);
nor U31505 (N_31505,N_31058,N_31405);
and U31506 (N_31506,N_31273,N_31010);
xnor U31507 (N_31507,N_31418,N_31174);
xnor U31508 (N_31508,N_31052,N_31410);
xnor U31509 (N_31509,N_31118,N_31059);
or U31510 (N_31510,N_31167,N_31239);
xor U31511 (N_31511,N_31201,N_31391);
xnor U31512 (N_31512,N_31164,N_31261);
or U31513 (N_31513,N_31298,N_31260);
nand U31514 (N_31514,N_31108,N_31212);
nand U31515 (N_31515,N_31233,N_31404);
nor U31516 (N_31516,N_31209,N_31104);
nor U31517 (N_31517,N_31308,N_31312);
xor U31518 (N_31518,N_31243,N_31445);
or U31519 (N_31519,N_31426,N_31251);
xnor U31520 (N_31520,N_31244,N_31439);
nand U31521 (N_31521,N_31181,N_31397);
xor U31522 (N_31522,N_31482,N_31131);
or U31523 (N_31523,N_31434,N_31035);
xnor U31524 (N_31524,N_31154,N_31462);
or U31525 (N_31525,N_31249,N_31143);
nand U31526 (N_31526,N_31012,N_31359);
and U31527 (N_31527,N_31489,N_31361);
or U31528 (N_31528,N_31223,N_31026);
nor U31529 (N_31529,N_31126,N_31471);
and U31530 (N_31530,N_31206,N_31088);
nor U31531 (N_31531,N_31316,N_31322);
and U31532 (N_31532,N_31307,N_31472);
nor U31533 (N_31533,N_31166,N_31175);
and U31534 (N_31534,N_31134,N_31013);
nor U31535 (N_31535,N_31494,N_31067);
and U31536 (N_31536,N_31050,N_31190);
nor U31537 (N_31537,N_31138,N_31480);
and U31538 (N_31538,N_31130,N_31215);
or U31539 (N_31539,N_31051,N_31449);
or U31540 (N_31540,N_31001,N_31037);
nand U31541 (N_31541,N_31333,N_31221);
nor U31542 (N_31542,N_31030,N_31412);
and U31543 (N_31543,N_31348,N_31269);
and U31544 (N_31544,N_31165,N_31022);
nand U31545 (N_31545,N_31485,N_31454);
nor U31546 (N_31546,N_31491,N_31474);
nand U31547 (N_31547,N_31219,N_31285);
xnor U31548 (N_31548,N_31265,N_31234);
nand U31549 (N_31549,N_31441,N_31179);
nand U31550 (N_31550,N_31087,N_31168);
nor U31551 (N_31551,N_31133,N_31171);
and U31552 (N_31552,N_31275,N_31458);
nor U31553 (N_31553,N_31198,N_31103);
or U31554 (N_31554,N_31369,N_31096);
xor U31555 (N_31555,N_31296,N_31237);
nand U31556 (N_31556,N_31325,N_31240);
nand U31557 (N_31557,N_31099,N_31204);
nand U31558 (N_31558,N_31072,N_31392);
or U31559 (N_31559,N_31173,N_31128);
or U31560 (N_31560,N_31289,N_31177);
nand U31561 (N_31561,N_31465,N_31015);
or U31562 (N_31562,N_31362,N_31250);
nand U31563 (N_31563,N_31347,N_31210);
or U31564 (N_31564,N_31342,N_31258);
xnor U31565 (N_31565,N_31195,N_31111);
xor U31566 (N_31566,N_31245,N_31406);
xnor U31567 (N_31567,N_31339,N_31176);
and U31568 (N_31568,N_31417,N_31033);
or U31569 (N_31569,N_31232,N_31194);
and U31570 (N_31570,N_31343,N_31425);
nand U31571 (N_31571,N_31490,N_31236);
nand U31572 (N_31572,N_31185,N_31414);
and U31573 (N_31573,N_31158,N_31427);
or U31574 (N_31574,N_31443,N_31467);
xor U31575 (N_31575,N_31302,N_31025);
and U31576 (N_31576,N_31129,N_31396);
or U31577 (N_31577,N_31428,N_31211);
nand U31578 (N_31578,N_31321,N_31469);
nor U31579 (N_31579,N_31303,N_31382);
or U31580 (N_31580,N_31123,N_31266);
or U31581 (N_31581,N_31057,N_31023);
nor U31582 (N_31582,N_31076,N_31120);
nand U31583 (N_31583,N_31358,N_31319);
or U31584 (N_31584,N_31300,N_31114);
xor U31585 (N_31585,N_31127,N_31438);
or U31586 (N_31586,N_31351,N_31378);
xor U31587 (N_31587,N_31079,N_31470);
nand U31588 (N_31588,N_31365,N_31460);
or U31589 (N_31589,N_31081,N_31376);
nor U31590 (N_31590,N_31180,N_31020);
nand U31591 (N_31591,N_31475,N_31323);
xnor U31592 (N_31592,N_31401,N_31301);
xnor U31593 (N_31593,N_31036,N_31218);
nand U31594 (N_31594,N_31207,N_31375);
and U31595 (N_31595,N_31446,N_31094);
and U31596 (N_31596,N_31197,N_31159);
nand U31597 (N_31597,N_31268,N_31436);
and U31598 (N_31598,N_31335,N_31297);
nor U31599 (N_31599,N_31373,N_31292);
and U31600 (N_31600,N_31242,N_31150);
and U31601 (N_31601,N_31422,N_31456);
xnor U31602 (N_31602,N_31355,N_31473);
or U31603 (N_31603,N_31336,N_31155);
and U31604 (N_31604,N_31077,N_31327);
or U31605 (N_31605,N_31157,N_31413);
and U31606 (N_31606,N_31043,N_31017);
or U31607 (N_31607,N_31091,N_31444);
nor U31608 (N_31608,N_31086,N_31383);
xor U31609 (N_31609,N_31332,N_31477);
or U31610 (N_31610,N_31069,N_31178);
nand U31611 (N_31611,N_31214,N_31016);
nand U31612 (N_31612,N_31487,N_31149);
nor U31613 (N_31613,N_31137,N_31125);
nand U31614 (N_31614,N_31281,N_31484);
and U31615 (N_31615,N_31113,N_31280);
xnor U31616 (N_31616,N_31254,N_31271);
nor U31617 (N_31617,N_31400,N_31070);
xnor U31618 (N_31618,N_31062,N_31027);
and U31619 (N_31619,N_31121,N_31419);
or U31620 (N_31620,N_31007,N_31220);
nand U31621 (N_31621,N_31082,N_31156);
and U31622 (N_31622,N_31151,N_31318);
nand U31623 (N_31623,N_31048,N_31442);
nand U31624 (N_31624,N_31424,N_31093);
and U31625 (N_31625,N_31450,N_31305);
nand U31626 (N_31626,N_31147,N_31196);
nand U31627 (N_31627,N_31056,N_31286);
nand U31628 (N_31628,N_31203,N_31064);
and U31629 (N_31629,N_31192,N_31235);
xnor U31630 (N_31630,N_31338,N_31109);
or U31631 (N_31631,N_31083,N_31119);
or U31632 (N_31632,N_31363,N_31183);
nor U31633 (N_31633,N_31011,N_31291);
nand U31634 (N_31634,N_31432,N_31344);
nor U31635 (N_31635,N_31047,N_31038);
nor U31636 (N_31636,N_31306,N_31481);
nand U31637 (N_31637,N_31049,N_31463);
nand U31638 (N_31638,N_31310,N_31352);
and U31639 (N_31639,N_31000,N_31388);
or U31640 (N_31640,N_31403,N_31409);
or U31641 (N_31641,N_31241,N_31092);
nand U31642 (N_31642,N_31205,N_31136);
and U31643 (N_31643,N_31357,N_31238);
xnor U31644 (N_31644,N_31466,N_31433);
and U31645 (N_31645,N_31097,N_31202);
xnor U31646 (N_31646,N_31153,N_31420);
nor U31647 (N_31647,N_31421,N_31372);
nor U31648 (N_31648,N_31112,N_31290);
and U31649 (N_31649,N_31430,N_31451);
and U31650 (N_31650,N_31374,N_31009);
nor U31651 (N_31651,N_31408,N_31386);
xor U31652 (N_31652,N_31063,N_31217);
and U31653 (N_31653,N_31457,N_31498);
nand U31654 (N_31654,N_31216,N_31334);
nand U31655 (N_31655,N_31499,N_31046);
and U31656 (N_31656,N_31106,N_31008);
or U31657 (N_31657,N_31073,N_31227);
xor U31658 (N_31658,N_31085,N_31315);
nand U31659 (N_31659,N_31452,N_31389);
and U31660 (N_31660,N_31304,N_31247);
or U31661 (N_31661,N_31478,N_31331);
nand U31662 (N_31662,N_31169,N_31019);
nor U31663 (N_31663,N_31287,N_31100);
and U31664 (N_31664,N_31170,N_31117);
nand U31665 (N_31665,N_31132,N_31055);
xor U31666 (N_31666,N_31222,N_31393);
xor U31667 (N_31667,N_31407,N_31071);
nor U31668 (N_31668,N_31225,N_31385);
or U31669 (N_31669,N_31399,N_31054);
nor U31670 (N_31670,N_31468,N_31142);
nand U31671 (N_31671,N_31040,N_31095);
nand U31672 (N_31672,N_31282,N_31279);
and U31673 (N_31673,N_31255,N_31492);
nor U31674 (N_31674,N_31380,N_31370);
or U31675 (N_31675,N_31431,N_31416);
xor U31676 (N_31676,N_31246,N_31116);
or U31677 (N_31677,N_31390,N_31288);
xor U31678 (N_31678,N_31395,N_31440);
xor U31679 (N_31679,N_31341,N_31213);
xnor U31680 (N_31680,N_31141,N_31146);
or U31681 (N_31681,N_31042,N_31188);
or U31682 (N_31682,N_31031,N_31329);
and U31683 (N_31683,N_31486,N_31224);
xor U31684 (N_31684,N_31311,N_31193);
nand U31685 (N_31685,N_31029,N_31002);
nor U31686 (N_31686,N_31264,N_31248);
nand U31687 (N_31687,N_31187,N_31263);
and U31688 (N_31688,N_31354,N_31488);
nor U31689 (N_31689,N_31018,N_31387);
nor U31690 (N_31690,N_31140,N_31004);
nand U31691 (N_31691,N_31186,N_31366);
nor U31692 (N_31692,N_31314,N_31084);
nand U31693 (N_31693,N_31024,N_31423);
xor U31694 (N_31694,N_31346,N_31496);
or U31695 (N_31695,N_31034,N_31272);
xnor U31696 (N_31696,N_31497,N_31252);
xnor U31697 (N_31697,N_31014,N_31461);
and U31698 (N_31698,N_31061,N_31283);
or U31699 (N_31699,N_31003,N_31299);
xor U31700 (N_31700,N_31415,N_31379);
or U31701 (N_31701,N_31045,N_31145);
nor U31702 (N_31702,N_31320,N_31278);
nand U31703 (N_31703,N_31356,N_31028);
nor U31704 (N_31704,N_31274,N_31367);
or U31705 (N_31705,N_31256,N_31191);
xor U31706 (N_31706,N_31074,N_31402);
and U31707 (N_31707,N_31144,N_31437);
and U31708 (N_31708,N_31350,N_31435);
nand U31709 (N_31709,N_31208,N_31345);
xnor U31710 (N_31710,N_31066,N_31453);
nor U31711 (N_31711,N_31039,N_31161);
nor U31712 (N_31712,N_31360,N_31078);
nor U31713 (N_31713,N_31182,N_31135);
and U31714 (N_31714,N_31276,N_31381);
and U31715 (N_31715,N_31162,N_31464);
and U31716 (N_31716,N_31006,N_31044);
nand U31717 (N_31717,N_31309,N_31495);
nand U31718 (N_31718,N_31340,N_31483);
nand U31719 (N_31719,N_31267,N_31102);
or U31720 (N_31720,N_31328,N_31277);
nor U31721 (N_31721,N_31021,N_31032);
nand U31722 (N_31722,N_31259,N_31160);
xor U31723 (N_31723,N_31326,N_31148);
and U31724 (N_31724,N_31448,N_31262);
xor U31725 (N_31725,N_31459,N_31493);
or U31726 (N_31726,N_31284,N_31172);
and U31727 (N_31727,N_31075,N_31317);
or U31728 (N_31728,N_31124,N_31349);
nand U31729 (N_31729,N_31199,N_31324);
nor U31730 (N_31730,N_31068,N_31455);
and U31731 (N_31731,N_31394,N_31122);
nand U31732 (N_31732,N_31139,N_31364);
nor U31733 (N_31733,N_31110,N_31041);
nand U31734 (N_31734,N_31295,N_31293);
nor U31735 (N_31735,N_31152,N_31115);
or U31736 (N_31736,N_31163,N_31189);
or U31737 (N_31737,N_31200,N_31270);
and U31738 (N_31738,N_31230,N_31294);
and U31739 (N_31739,N_31098,N_31080);
or U31740 (N_31740,N_31377,N_31398);
xor U31741 (N_31741,N_31228,N_31005);
or U31742 (N_31742,N_31257,N_31226);
nand U31743 (N_31743,N_31065,N_31384);
and U31744 (N_31744,N_31253,N_31313);
or U31745 (N_31745,N_31476,N_31330);
or U31746 (N_31746,N_31105,N_31090);
nand U31747 (N_31747,N_31371,N_31089);
or U31748 (N_31748,N_31053,N_31479);
xor U31749 (N_31749,N_31184,N_31107);
nor U31750 (N_31750,N_31310,N_31280);
or U31751 (N_31751,N_31494,N_31097);
nor U31752 (N_31752,N_31300,N_31474);
xor U31753 (N_31753,N_31218,N_31085);
or U31754 (N_31754,N_31325,N_31356);
xnor U31755 (N_31755,N_31468,N_31187);
nor U31756 (N_31756,N_31361,N_31112);
and U31757 (N_31757,N_31233,N_31151);
xnor U31758 (N_31758,N_31332,N_31465);
nor U31759 (N_31759,N_31012,N_31048);
or U31760 (N_31760,N_31488,N_31162);
nand U31761 (N_31761,N_31241,N_31207);
nand U31762 (N_31762,N_31175,N_31182);
nand U31763 (N_31763,N_31063,N_31169);
or U31764 (N_31764,N_31096,N_31336);
nand U31765 (N_31765,N_31327,N_31301);
nor U31766 (N_31766,N_31067,N_31196);
or U31767 (N_31767,N_31346,N_31166);
and U31768 (N_31768,N_31142,N_31473);
and U31769 (N_31769,N_31238,N_31421);
or U31770 (N_31770,N_31227,N_31372);
nor U31771 (N_31771,N_31317,N_31428);
xnor U31772 (N_31772,N_31165,N_31051);
nand U31773 (N_31773,N_31055,N_31246);
or U31774 (N_31774,N_31475,N_31187);
nor U31775 (N_31775,N_31038,N_31467);
nand U31776 (N_31776,N_31130,N_31125);
nand U31777 (N_31777,N_31131,N_31121);
nand U31778 (N_31778,N_31061,N_31176);
and U31779 (N_31779,N_31402,N_31025);
nor U31780 (N_31780,N_31137,N_31138);
nor U31781 (N_31781,N_31180,N_31434);
nand U31782 (N_31782,N_31124,N_31262);
or U31783 (N_31783,N_31065,N_31160);
nor U31784 (N_31784,N_31046,N_31076);
nand U31785 (N_31785,N_31087,N_31140);
nand U31786 (N_31786,N_31132,N_31445);
and U31787 (N_31787,N_31431,N_31434);
or U31788 (N_31788,N_31402,N_31290);
nor U31789 (N_31789,N_31182,N_31430);
xnor U31790 (N_31790,N_31163,N_31374);
xnor U31791 (N_31791,N_31359,N_31437);
or U31792 (N_31792,N_31498,N_31148);
or U31793 (N_31793,N_31451,N_31235);
nand U31794 (N_31794,N_31184,N_31145);
nand U31795 (N_31795,N_31129,N_31265);
nor U31796 (N_31796,N_31227,N_31049);
nand U31797 (N_31797,N_31135,N_31142);
or U31798 (N_31798,N_31390,N_31485);
and U31799 (N_31799,N_31064,N_31178);
nand U31800 (N_31800,N_31144,N_31200);
nand U31801 (N_31801,N_31096,N_31048);
nor U31802 (N_31802,N_31211,N_31003);
nor U31803 (N_31803,N_31122,N_31342);
xor U31804 (N_31804,N_31319,N_31079);
nor U31805 (N_31805,N_31217,N_31339);
and U31806 (N_31806,N_31160,N_31319);
or U31807 (N_31807,N_31470,N_31283);
and U31808 (N_31808,N_31058,N_31418);
or U31809 (N_31809,N_31234,N_31019);
nand U31810 (N_31810,N_31362,N_31288);
nand U31811 (N_31811,N_31298,N_31361);
nand U31812 (N_31812,N_31386,N_31198);
xnor U31813 (N_31813,N_31076,N_31363);
nor U31814 (N_31814,N_31332,N_31364);
nand U31815 (N_31815,N_31331,N_31106);
and U31816 (N_31816,N_31009,N_31196);
nor U31817 (N_31817,N_31185,N_31064);
nand U31818 (N_31818,N_31121,N_31284);
xor U31819 (N_31819,N_31400,N_31186);
nor U31820 (N_31820,N_31439,N_31309);
nor U31821 (N_31821,N_31449,N_31120);
nand U31822 (N_31822,N_31055,N_31007);
and U31823 (N_31823,N_31325,N_31285);
nand U31824 (N_31824,N_31173,N_31049);
nor U31825 (N_31825,N_31372,N_31441);
and U31826 (N_31826,N_31225,N_31496);
or U31827 (N_31827,N_31224,N_31042);
and U31828 (N_31828,N_31026,N_31391);
nand U31829 (N_31829,N_31458,N_31488);
nand U31830 (N_31830,N_31357,N_31354);
and U31831 (N_31831,N_31057,N_31234);
nor U31832 (N_31832,N_31413,N_31058);
or U31833 (N_31833,N_31195,N_31032);
or U31834 (N_31834,N_31149,N_31169);
nand U31835 (N_31835,N_31337,N_31486);
and U31836 (N_31836,N_31111,N_31077);
nand U31837 (N_31837,N_31404,N_31495);
xor U31838 (N_31838,N_31010,N_31395);
nor U31839 (N_31839,N_31254,N_31021);
nor U31840 (N_31840,N_31142,N_31343);
xor U31841 (N_31841,N_31273,N_31154);
xor U31842 (N_31842,N_31335,N_31372);
and U31843 (N_31843,N_31452,N_31399);
nor U31844 (N_31844,N_31128,N_31317);
xor U31845 (N_31845,N_31296,N_31423);
nor U31846 (N_31846,N_31165,N_31329);
nor U31847 (N_31847,N_31091,N_31137);
nand U31848 (N_31848,N_31023,N_31071);
or U31849 (N_31849,N_31420,N_31173);
and U31850 (N_31850,N_31069,N_31102);
and U31851 (N_31851,N_31470,N_31106);
nor U31852 (N_31852,N_31243,N_31074);
nand U31853 (N_31853,N_31398,N_31467);
nor U31854 (N_31854,N_31337,N_31368);
and U31855 (N_31855,N_31076,N_31078);
and U31856 (N_31856,N_31296,N_31245);
or U31857 (N_31857,N_31011,N_31430);
xor U31858 (N_31858,N_31466,N_31216);
or U31859 (N_31859,N_31240,N_31233);
xnor U31860 (N_31860,N_31093,N_31416);
xnor U31861 (N_31861,N_31420,N_31051);
xor U31862 (N_31862,N_31105,N_31389);
and U31863 (N_31863,N_31294,N_31347);
nand U31864 (N_31864,N_31060,N_31288);
or U31865 (N_31865,N_31350,N_31287);
nand U31866 (N_31866,N_31027,N_31475);
xor U31867 (N_31867,N_31253,N_31159);
and U31868 (N_31868,N_31238,N_31193);
nor U31869 (N_31869,N_31389,N_31399);
nand U31870 (N_31870,N_31017,N_31104);
or U31871 (N_31871,N_31387,N_31309);
or U31872 (N_31872,N_31255,N_31226);
nor U31873 (N_31873,N_31289,N_31008);
and U31874 (N_31874,N_31111,N_31042);
xor U31875 (N_31875,N_31228,N_31064);
or U31876 (N_31876,N_31350,N_31395);
nor U31877 (N_31877,N_31430,N_31360);
xor U31878 (N_31878,N_31305,N_31397);
and U31879 (N_31879,N_31214,N_31494);
nand U31880 (N_31880,N_31117,N_31317);
and U31881 (N_31881,N_31106,N_31231);
or U31882 (N_31882,N_31264,N_31022);
xnor U31883 (N_31883,N_31401,N_31118);
nand U31884 (N_31884,N_31433,N_31367);
or U31885 (N_31885,N_31169,N_31353);
and U31886 (N_31886,N_31484,N_31390);
or U31887 (N_31887,N_31447,N_31053);
nor U31888 (N_31888,N_31108,N_31160);
and U31889 (N_31889,N_31478,N_31240);
xnor U31890 (N_31890,N_31283,N_31262);
xnor U31891 (N_31891,N_31123,N_31172);
or U31892 (N_31892,N_31248,N_31321);
and U31893 (N_31893,N_31272,N_31441);
nand U31894 (N_31894,N_31075,N_31043);
nor U31895 (N_31895,N_31352,N_31495);
or U31896 (N_31896,N_31055,N_31260);
xor U31897 (N_31897,N_31209,N_31305);
and U31898 (N_31898,N_31404,N_31301);
nor U31899 (N_31899,N_31399,N_31240);
nand U31900 (N_31900,N_31263,N_31310);
nor U31901 (N_31901,N_31281,N_31429);
or U31902 (N_31902,N_31165,N_31116);
xnor U31903 (N_31903,N_31169,N_31066);
nor U31904 (N_31904,N_31064,N_31421);
and U31905 (N_31905,N_31303,N_31356);
nor U31906 (N_31906,N_31353,N_31126);
or U31907 (N_31907,N_31251,N_31345);
nand U31908 (N_31908,N_31478,N_31078);
and U31909 (N_31909,N_31283,N_31401);
xor U31910 (N_31910,N_31215,N_31125);
nor U31911 (N_31911,N_31038,N_31245);
and U31912 (N_31912,N_31445,N_31075);
and U31913 (N_31913,N_31166,N_31330);
nand U31914 (N_31914,N_31169,N_31227);
xor U31915 (N_31915,N_31469,N_31237);
nor U31916 (N_31916,N_31163,N_31256);
xor U31917 (N_31917,N_31149,N_31277);
nor U31918 (N_31918,N_31018,N_31155);
nor U31919 (N_31919,N_31043,N_31029);
nand U31920 (N_31920,N_31434,N_31355);
and U31921 (N_31921,N_31329,N_31003);
or U31922 (N_31922,N_31348,N_31061);
and U31923 (N_31923,N_31292,N_31074);
and U31924 (N_31924,N_31173,N_31131);
and U31925 (N_31925,N_31140,N_31161);
and U31926 (N_31926,N_31352,N_31028);
and U31927 (N_31927,N_31017,N_31444);
or U31928 (N_31928,N_31023,N_31172);
nor U31929 (N_31929,N_31472,N_31054);
and U31930 (N_31930,N_31025,N_31439);
or U31931 (N_31931,N_31309,N_31233);
xor U31932 (N_31932,N_31399,N_31442);
or U31933 (N_31933,N_31215,N_31445);
nand U31934 (N_31934,N_31010,N_31201);
nand U31935 (N_31935,N_31245,N_31250);
nor U31936 (N_31936,N_31469,N_31126);
nand U31937 (N_31937,N_31104,N_31185);
and U31938 (N_31938,N_31409,N_31033);
and U31939 (N_31939,N_31124,N_31116);
and U31940 (N_31940,N_31430,N_31282);
nand U31941 (N_31941,N_31142,N_31057);
and U31942 (N_31942,N_31139,N_31055);
nand U31943 (N_31943,N_31103,N_31121);
nor U31944 (N_31944,N_31062,N_31001);
nand U31945 (N_31945,N_31209,N_31077);
nor U31946 (N_31946,N_31406,N_31247);
and U31947 (N_31947,N_31374,N_31471);
xnor U31948 (N_31948,N_31327,N_31056);
or U31949 (N_31949,N_31435,N_31254);
nor U31950 (N_31950,N_31111,N_31019);
nor U31951 (N_31951,N_31489,N_31189);
xor U31952 (N_31952,N_31083,N_31186);
nor U31953 (N_31953,N_31081,N_31063);
and U31954 (N_31954,N_31329,N_31262);
nand U31955 (N_31955,N_31243,N_31228);
nor U31956 (N_31956,N_31266,N_31245);
or U31957 (N_31957,N_31149,N_31272);
or U31958 (N_31958,N_31294,N_31143);
and U31959 (N_31959,N_31443,N_31259);
nor U31960 (N_31960,N_31423,N_31345);
xor U31961 (N_31961,N_31042,N_31108);
xor U31962 (N_31962,N_31369,N_31201);
and U31963 (N_31963,N_31132,N_31082);
or U31964 (N_31964,N_31215,N_31376);
xnor U31965 (N_31965,N_31490,N_31093);
nand U31966 (N_31966,N_31121,N_31476);
and U31967 (N_31967,N_31145,N_31361);
nor U31968 (N_31968,N_31113,N_31479);
and U31969 (N_31969,N_31122,N_31108);
and U31970 (N_31970,N_31068,N_31333);
and U31971 (N_31971,N_31156,N_31403);
xnor U31972 (N_31972,N_31490,N_31402);
or U31973 (N_31973,N_31477,N_31131);
or U31974 (N_31974,N_31158,N_31414);
or U31975 (N_31975,N_31323,N_31041);
nor U31976 (N_31976,N_31020,N_31152);
or U31977 (N_31977,N_31333,N_31477);
and U31978 (N_31978,N_31265,N_31473);
nand U31979 (N_31979,N_31268,N_31312);
xor U31980 (N_31980,N_31050,N_31244);
or U31981 (N_31981,N_31182,N_31257);
and U31982 (N_31982,N_31080,N_31265);
nor U31983 (N_31983,N_31246,N_31214);
or U31984 (N_31984,N_31239,N_31116);
or U31985 (N_31985,N_31137,N_31077);
xnor U31986 (N_31986,N_31133,N_31381);
nand U31987 (N_31987,N_31493,N_31190);
nand U31988 (N_31988,N_31110,N_31205);
nand U31989 (N_31989,N_31376,N_31429);
xnor U31990 (N_31990,N_31410,N_31190);
or U31991 (N_31991,N_31401,N_31216);
xnor U31992 (N_31992,N_31205,N_31093);
or U31993 (N_31993,N_31200,N_31194);
xor U31994 (N_31994,N_31353,N_31091);
nand U31995 (N_31995,N_31194,N_31271);
nor U31996 (N_31996,N_31299,N_31121);
or U31997 (N_31997,N_31449,N_31388);
nand U31998 (N_31998,N_31026,N_31352);
xnor U31999 (N_31999,N_31231,N_31471);
and U32000 (N_32000,N_31764,N_31675);
and U32001 (N_32001,N_31527,N_31679);
or U32002 (N_32002,N_31597,N_31708);
and U32003 (N_32003,N_31676,N_31536);
xnor U32004 (N_32004,N_31530,N_31658);
nand U32005 (N_32005,N_31909,N_31517);
xor U32006 (N_32006,N_31816,N_31590);
xor U32007 (N_32007,N_31569,N_31721);
nand U32008 (N_32008,N_31800,N_31712);
nor U32009 (N_32009,N_31953,N_31626);
nand U32010 (N_32010,N_31524,N_31638);
xor U32011 (N_32011,N_31987,N_31560);
or U32012 (N_32012,N_31703,N_31904);
and U32013 (N_32013,N_31596,N_31557);
nand U32014 (N_32014,N_31746,N_31575);
or U32015 (N_32015,N_31965,N_31775);
nand U32016 (N_32016,N_31573,N_31635);
or U32017 (N_32017,N_31651,N_31821);
nand U32018 (N_32018,N_31879,N_31898);
or U32019 (N_32019,N_31755,N_31686);
nor U32020 (N_32020,N_31995,N_31789);
nor U32021 (N_32021,N_31641,N_31699);
or U32022 (N_32022,N_31839,N_31788);
nor U32023 (N_32023,N_31563,N_31790);
nor U32024 (N_32024,N_31678,N_31667);
or U32025 (N_32025,N_31897,N_31634);
and U32026 (N_32026,N_31617,N_31759);
nand U32027 (N_32027,N_31663,N_31750);
nand U32028 (N_32028,N_31916,N_31896);
nand U32029 (N_32029,N_31792,N_31691);
or U32030 (N_32030,N_31521,N_31911);
and U32031 (N_32031,N_31808,N_31562);
and U32032 (N_32032,N_31858,N_31594);
nor U32033 (N_32033,N_31545,N_31880);
nor U32034 (N_32034,N_31900,N_31556);
and U32035 (N_32035,N_31883,N_31811);
nor U32036 (N_32036,N_31551,N_31851);
nor U32037 (N_32037,N_31512,N_31528);
nand U32038 (N_32038,N_31623,N_31797);
nor U32039 (N_32039,N_31786,N_31662);
nand U32040 (N_32040,N_31720,N_31892);
or U32041 (N_32041,N_31829,N_31583);
xor U32042 (N_32042,N_31544,N_31922);
and U32043 (N_32043,N_31719,N_31985);
and U32044 (N_32044,N_31671,N_31571);
or U32045 (N_32045,N_31867,N_31624);
nor U32046 (N_32046,N_31593,N_31730);
nand U32047 (N_32047,N_31869,N_31749);
nand U32048 (N_32048,N_31606,N_31998);
xor U32049 (N_32049,N_31503,N_31502);
xnor U32050 (N_32050,N_31716,N_31710);
nand U32051 (N_32051,N_31983,N_31840);
xor U32052 (N_32052,N_31973,N_31768);
nand U32053 (N_32053,N_31625,N_31842);
nor U32054 (N_32054,N_31529,N_31933);
or U32055 (N_32055,N_31519,N_31516);
nor U32056 (N_32056,N_31866,N_31612);
and U32057 (N_32057,N_31872,N_31705);
or U32058 (N_32058,N_31543,N_31802);
and U32059 (N_32059,N_31685,N_31500);
nor U32060 (N_32060,N_31828,N_31784);
nand U32061 (N_32061,N_31632,N_31574);
xor U32062 (N_32062,N_31779,N_31853);
or U32063 (N_32063,N_31731,N_31567);
nor U32064 (N_32064,N_31857,N_31511);
and U32065 (N_32065,N_31780,N_31949);
or U32066 (N_32066,N_31628,N_31614);
nand U32067 (N_32067,N_31599,N_31548);
or U32068 (N_32068,N_31549,N_31694);
nor U32069 (N_32069,N_31927,N_31928);
xnor U32070 (N_32070,N_31656,N_31977);
and U32071 (N_32071,N_31868,N_31581);
xor U32072 (N_32072,N_31813,N_31728);
nor U32073 (N_32073,N_31837,N_31564);
nand U32074 (N_32074,N_31958,N_31974);
nor U32075 (N_32075,N_31769,N_31739);
xnor U32076 (N_32076,N_31706,N_31997);
and U32077 (N_32077,N_31937,N_31665);
and U32078 (N_32078,N_31627,N_31700);
or U32079 (N_32079,N_31893,N_31591);
xnor U32080 (N_32080,N_31696,N_31863);
or U32081 (N_32081,N_31946,N_31902);
or U32082 (N_32082,N_31692,N_31535);
nand U32083 (N_32083,N_31763,N_31538);
or U32084 (N_32084,N_31738,N_31752);
and U32085 (N_32085,N_31615,N_31670);
or U32086 (N_32086,N_31783,N_31920);
nor U32087 (N_32087,N_31558,N_31981);
nor U32088 (N_32088,N_31992,N_31772);
xnor U32089 (N_32089,N_31794,N_31509);
and U32090 (N_32090,N_31885,N_31602);
and U32091 (N_32091,N_31770,N_31709);
and U32092 (N_32092,N_31609,N_31773);
or U32093 (N_32093,N_31899,N_31585);
and U32094 (N_32094,N_31541,N_31537);
nor U32095 (N_32095,N_31774,N_31950);
or U32096 (N_32096,N_31723,N_31823);
or U32097 (N_32097,N_31669,N_31979);
and U32098 (N_32098,N_31849,N_31637);
or U32099 (N_32099,N_31994,N_31782);
or U32100 (N_32100,N_31832,N_31830);
xor U32101 (N_32101,N_31926,N_31865);
nor U32102 (N_32102,N_31835,N_31971);
nor U32103 (N_32103,N_31929,N_31912);
xor U32104 (N_32104,N_31781,N_31682);
and U32105 (N_32105,N_31684,N_31621);
xnor U32106 (N_32106,N_31807,N_31776);
nor U32107 (N_32107,N_31903,N_31777);
or U32108 (N_32108,N_31951,N_31742);
nor U32109 (N_32109,N_31827,N_31944);
and U32110 (N_32110,N_31955,N_31834);
and U32111 (N_32111,N_31598,N_31714);
and U32112 (N_32112,N_31673,N_31921);
xor U32113 (N_32113,N_31826,N_31644);
nand U32114 (N_32114,N_31841,N_31934);
and U32115 (N_32115,N_31613,N_31554);
xnor U32116 (N_32116,N_31646,N_31963);
xor U32117 (N_32117,N_31765,N_31859);
xnor U32118 (N_32118,N_31870,N_31622);
nand U32119 (N_32119,N_31724,N_31793);
or U32120 (N_32120,N_31999,N_31932);
and U32121 (N_32121,N_31820,N_31855);
nand U32122 (N_32122,N_31751,N_31910);
xor U32123 (N_32123,N_31578,N_31510);
nor U32124 (N_32124,N_31856,N_31532);
or U32125 (N_32125,N_31636,N_31603);
nand U32126 (N_32126,N_31861,N_31580);
or U32127 (N_32127,N_31570,N_31875);
and U32128 (N_32128,N_31520,N_31812);
or U32129 (N_32129,N_31822,N_31674);
xor U32130 (N_32130,N_31982,N_31889);
or U32131 (N_32131,N_31744,N_31843);
and U32132 (N_32132,N_31577,N_31975);
or U32133 (N_32133,N_31552,N_31639);
xnor U32134 (N_32134,N_31688,N_31559);
xor U32135 (N_32135,N_31931,N_31918);
xor U32136 (N_32136,N_31957,N_31796);
xor U32137 (N_32137,N_31905,N_31989);
or U32138 (N_32138,N_31605,N_31726);
nor U32139 (N_32139,N_31876,N_31846);
or U32140 (N_32140,N_31631,N_31653);
nor U32141 (N_32141,N_31972,N_31702);
nand U32142 (N_32142,N_31761,N_31962);
and U32143 (N_32143,N_31534,N_31546);
and U32144 (N_32144,N_31939,N_31745);
xnor U32145 (N_32145,N_31785,N_31589);
nand U32146 (N_32146,N_31514,N_31757);
nor U32147 (N_32147,N_31672,N_31533);
or U32148 (N_32148,N_31588,N_31791);
and U32149 (N_32149,N_31809,N_31566);
xor U32150 (N_32150,N_31988,N_31917);
xnor U32151 (N_32151,N_31649,N_31586);
nand U32152 (N_32152,N_31718,N_31758);
nor U32153 (N_32153,N_31592,N_31945);
nor U32154 (N_32154,N_31818,N_31683);
and U32155 (N_32155,N_31753,N_31923);
nor U32156 (N_32156,N_31938,N_31760);
and U32157 (N_32157,N_31930,N_31844);
xnor U32158 (N_32158,N_31640,N_31824);
nor U32159 (N_32159,N_31984,N_31762);
nor U32160 (N_32160,N_31801,N_31959);
xnor U32161 (N_32161,N_31711,N_31740);
nand U32162 (N_32162,N_31795,N_31831);
nor U32163 (N_32163,N_31991,N_31810);
and U32164 (N_32164,N_31687,N_31630);
or U32165 (N_32165,N_31970,N_31924);
and U32166 (N_32166,N_31913,N_31736);
nor U32167 (N_32167,N_31996,N_31864);
xor U32168 (N_32168,N_31664,N_31960);
or U32169 (N_32169,N_31969,N_31914);
nand U32170 (N_32170,N_31607,N_31819);
and U32171 (N_32171,N_31961,N_31715);
xor U32172 (N_32172,N_31778,N_31610);
nand U32173 (N_32173,N_31689,N_31704);
xnor U32174 (N_32174,N_31925,N_31964);
nor U32175 (N_32175,N_31659,N_31525);
or U32176 (N_32176,N_31803,N_31652);
or U32177 (N_32177,N_31815,N_31756);
or U32178 (N_32178,N_31513,N_31968);
nand U32179 (N_32179,N_31894,N_31884);
xor U32180 (N_32180,N_31542,N_31732);
or U32181 (N_32181,N_31978,N_31725);
and U32182 (N_32182,N_31854,N_31943);
and U32183 (N_32183,N_31619,N_31915);
xor U32184 (N_32184,N_31695,N_31547);
xor U32185 (N_32185,N_31572,N_31648);
and U32186 (N_32186,N_31729,N_31805);
nand U32187 (N_32187,N_31741,N_31845);
nand U32188 (N_32188,N_31947,N_31690);
xor U32189 (N_32189,N_31908,N_31936);
xor U32190 (N_32190,N_31806,N_31874);
nand U32191 (N_32191,N_31817,N_31666);
nor U32192 (N_32192,N_31655,N_31748);
or U32193 (N_32193,N_31647,N_31852);
xor U32194 (N_32194,N_31595,N_31515);
and U32195 (N_32195,N_31787,N_31713);
xor U32196 (N_32196,N_31941,N_31940);
nor U32197 (N_32197,N_31587,N_31661);
nor U32198 (N_32198,N_31561,N_31531);
nor U32199 (N_32199,N_31838,N_31501);
nand U32200 (N_32200,N_31507,N_31767);
nor U32201 (N_32201,N_31608,N_31919);
nor U32202 (N_32202,N_31717,N_31754);
nor U32203 (N_32203,N_31873,N_31871);
nand U32204 (N_32204,N_31901,N_31771);
and U32205 (N_32205,N_31954,N_31886);
nand U32206 (N_32206,N_31565,N_31860);
nand U32207 (N_32207,N_31747,N_31967);
xor U32208 (N_32208,N_31836,N_31798);
xor U32209 (N_32209,N_31727,N_31993);
nand U32210 (N_32210,N_31506,N_31660);
nand U32211 (N_32211,N_31743,N_31604);
and U32212 (N_32212,N_31518,N_31980);
and U32213 (N_32213,N_31707,N_31523);
nand U32214 (N_32214,N_31733,N_31877);
and U32215 (N_32215,N_31654,N_31956);
xor U32216 (N_32216,N_31847,N_31505);
and U32217 (N_32217,N_31701,N_31539);
and U32218 (N_32218,N_31633,N_31576);
nand U32219 (N_32219,N_31948,N_31553);
or U32220 (N_32220,N_31976,N_31555);
nor U32221 (N_32221,N_31526,N_31522);
nor U32222 (N_32222,N_31907,N_31722);
and U32223 (N_32223,N_31584,N_31906);
or U32224 (N_32224,N_31814,N_31890);
nand U32225 (N_32225,N_31881,N_31579);
and U32226 (N_32226,N_31986,N_31618);
xor U32227 (N_32227,N_31620,N_31766);
nor U32228 (N_32228,N_31887,N_31735);
xnor U32229 (N_32229,N_31650,N_31862);
xor U32230 (N_32230,N_31540,N_31850);
and U32231 (N_32231,N_31643,N_31833);
nor U32232 (N_32232,N_31990,N_31616);
nor U32233 (N_32233,N_31799,N_31966);
and U32234 (N_32234,N_31645,N_31878);
and U32235 (N_32235,N_31942,N_31600);
or U32236 (N_32236,N_31825,N_31601);
nand U32237 (N_32237,N_31737,N_31848);
nor U32238 (N_32238,N_31681,N_31952);
nand U32239 (N_32239,N_31677,N_31582);
xnor U32240 (N_32240,N_31504,N_31697);
xnor U32241 (N_32241,N_31895,N_31698);
nand U32242 (N_32242,N_31550,N_31804);
and U32243 (N_32243,N_31642,N_31629);
or U32244 (N_32244,N_31568,N_31891);
and U32245 (N_32245,N_31668,N_31611);
nand U32246 (N_32246,N_31935,N_31508);
or U32247 (N_32247,N_31680,N_31882);
or U32248 (N_32248,N_31734,N_31888);
nor U32249 (N_32249,N_31693,N_31657);
xnor U32250 (N_32250,N_31973,N_31821);
nand U32251 (N_32251,N_31657,N_31574);
xnor U32252 (N_32252,N_31648,N_31968);
xor U32253 (N_32253,N_31925,N_31672);
or U32254 (N_32254,N_31854,N_31550);
and U32255 (N_32255,N_31722,N_31662);
xnor U32256 (N_32256,N_31863,N_31924);
and U32257 (N_32257,N_31878,N_31917);
or U32258 (N_32258,N_31527,N_31723);
or U32259 (N_32259,N_31638,N_31964);
or U32260 (N_32260,N_31900,N_31743);
nor U32261 (N_32261,N_31925,N_31635);
xnor U32262 (N_32262,N_31798,N_31640);
nor U32263 (N_32263,N_31614,N_31804);
or U32264 (N_32264,N_31520,N_31761);
and U32265 (N_32265,N_31554,N_31758);
and U32266 (N_32266,N_31526,N_31930);
nor U32267 (N_32267,N_31578,N_31914);
or U32268 (N_32268,N_31583,N_31623);
nand U32269 (N_32269,N_31631,N_31904);
xnor U32270 (N_32270,N_31881,N_31529);
xor U32271 (N_32271,N_31666,N_31871);
xor U32272 (N_32272,N_31692,N_31887);
and U32273 (N_32273,N_31600,N_31924);
nand U32274 (N_32274,N_31910,N_31972);
xor U32275 (N_32275,N_31775,N_31506);
xnor U32276 (N_32276,N_31684,N_31562);
and U32277 (N_32277,N_31662,N_31724);
xnor U32278 (N_32278,N_31928,N_31820);
and U32279 (N_32279,N_31863,N_31543);
xnor U32280 (N_32280,N_31862,N_31928);
and U32281 (N_32281,N_31892,N_31845);
nand U32282 (N_32282,N_31746,N_31840);
nor U32283 (N_32283,N_31533,N_31980);
and U32284 (N_32284,N_31696,N_31588);
xnor U32285 (N_32285,N_31811,N_31544);
nor U32286 (N_32286,N_31682,N_31592);
xnor U32287 (N_32287,N_31644,N_31564);
or U32288 (N_32288,N_31809,N_31958);
xor U32289 (N_32289,N_31839,N_31560);
and U32290 (N_32290,N_31930,N_31847);
nor U32291 (N_32291,N_31509,N_31852);
xor U32292 (N_32292,N_31691,N_31512);
nand U32293 (N_32293,N_31578,N_31799);
nor U32294 (N_32294,N_31758,N_31660);
or U32295 (N_32295,N_31856,N_31528);
nor U32296 (N_32296,N_31666,N_31799);
or U32297 (N_32297,N_31730,N_31556);
and U32298 (N_32298,N_31819,N_31998);
or U32299 (N_32299,N_31866,N_31990);
or U32300 (N_32300,N_31921,N_31924);
nand U32301 (N_32301,N_31575,N_31629);
xor U32302 (N_32302,N_31926,N_31734);
nor U32303 (N_32303,N_31626,N_31639);
xor U32304 (N_32304,N_31791,N_31696);
and U32305 (N_32305,N_31728,N_31746);
and U32306 (N_32306,N_31505,N_31842);
nor U32307 (N_32307,N_31677,N_31902);
nor U32308 (N_32308,N_31506,N_31598);
nand U32309 (N_32309,N_31718,N_31741);
xor U32310 (N_32310,N_31504,N_31962);
and U32311 (N_32311,N_31588,N_31653);
and U32312 (N_32312,N_31792,N_31814);
and U32313 (N_32313,N_31882,N_31900);
xor U32314 (N_32314,N_31728,N_31847);
and U32315 (N_32315,N_31786,N_31543);
nand U32316 (N_32316,N_31978,N_31619);
nand U32317 (N_32317,N_31891,N_31941);
nor U32318 (N_32318,N_31558,N_31896);
xnor U32319 (N_32319,N_31664,N_31832);
nand U32320 (N_32320,N_31980,N_31896);
and U32321 (N_32321,N_31680,N_31879);
xnor U32322 (N_32322,N_31570,N_31907);
nor U32323 (N_32323,N_31593,N_31952);
nand U32324 (N_32324,N_31684,N_31532);
or U32325 (N_32325,N_31634,N_31787);
xnor U32326 (N_32326,N_31815,N_31508);
xor U32327 (N_32327,N_31817,N_31983);
and U32328 (N_32328,N_31960,N_31696);
or U32329 (N_32329,N_31611,N_31939);
and U32330 (N_32330,N_31586,N_31733);
or U32331 (N_32331,N_31875,N_31972);
or U32332 (N_32332,N_31762,N_31772);
xnor U32333 (N_32333,N_31866,N_31941);
xnor U32334 (N_32334,N_31777,N_31933);
xnor U32335 (N_32335,N_31931,N_31714);
nand U32336 (N_32336,N_31916,N_31901);
or U32337 (N_32337,N_31580,N_31522);
or U32338 (N_32338,N_31928,N_31745);
and U32339 (N_32339,N_31714,N_31799);
xor U32340 (N_32340,N_31901,N_31793);
and U32341 (N_32341,N_31808,N_31748);
xnor U32342 (N_32342,N_31822,N_31802);
xnor U32343 (N_32343,N_31902,N_31624);
xnor U32344 (N_32344,N_31718,N_31707);
or U32345 (N_32345,N_31913,N_31825);
or U32346 (N_32346,N_31891,N_31776);
nand U32347 (N_32347,N_31500,N_31697);
xor U32348 (N_32348,N_31573,N_31654);
and U32349 (N_32349,N_31698,N_31562);
xor U32350 (N_32350,N_31673,N_31651);
xnor U32351 (N_32351,N_31507,N_31868);
xor U32352 (N_32352,N_31683,N_31781);
nand U32353 (N_32353,N_31530,N_31883);
or U32354 (N_32354,N_31589,N_31515);
and U32355 (N_32355,N_31751,N_31795);
and U32356 (N_32356,N_31651,N_31848);
nor U32357 (N_32357,N_31845,N_31947);
and U32358 (N_32358,N_31955,N_31734);
xor U32359 (N_32359,N_31750,N_31714);
and U32360 (N_32360,N_31652,N_31632);
nand U32361 (N_32361,N_31783,N_31683);
xnor U32362 (N_32362,N_31545,N_31697);
nand U32363 (N_32363,N_31785,N_31502);
xor U32364 (N_32364,N_31816,N_31625);
nand U32365 (N_32365,N_31935,N_31820);
xnor U32366 (N_32366,N_31806,N_31696);
nor U32367 (N_32367,N_31579,N_31883);
or U32368 (N_32368,N_31909,N_31628);
nand U32369 (N_32369,N_31962,N_31804);
nor U32370 (N_32370,N_31743,N_31876);
xnor U32371 (N_32371,N_31898,N_31760);
nor U32372 (N_32372,N_31575,N_31983);
nand U32373 (N_32373,N_31799,N_31671);
xor U32374 (N_32374,N_31984,N_31780);
and U32375 (N_32375,N_31980,N_31620);
nand U32376 (N_32376,N_31644,N_31612);
or U32377 (N_32377,N_31878,N_31644);
xnor U32378 (N_32378,N_31680,N_31864);
nor U32379 (N_32379,N_31642,N_31588);
nand U32380 (N_32380,N_31681,N_31818);
and U32381 (N_32381,N_31507,N_31575);
nor U32382 (N_32382,N_31565,N_31952);
and U32383 (N_32383,N_31545,N_31930);
and U32384 (N_32384,N_31605,N_31505);
or U32385 (N_32385,N_31727,N_31520);
nor U32386 (N_32386,N_31620,N_31511);
nand U32387 (N_32387,N_31725,N_31950);
xor U32388 (N_32388,N_31760,N_31633);
or U32389 (N_32389,N_31516,N_31722);
or U32390 (N_32390,N_31821,N_31560);
or U32391 (N_32391,N_31749,N_31541);
or U32392 (N_32392,N_31788,N_31861);
nand U32393 (N_32393,N_31783,N_31735);
or U32394 (N_32394,N_31911,N_31656);
nand U32395 (N_32395,N_31507,N_31565);
or U32396 (N_32396,N_31835,N_31913);
xnor U32397 (N_32397,N_31531,N_31555);
and U32398 (N_32398,N_31942,N_31905);
xnor U32399 (N_32399,N_31829,N_31592);
or U32400 (N_32400,N_31975,N_31844);
xor U32401 (N_32401,N_31845,N_31792);
nand U32402 (N_32402,N_31698,N_31892);
nand U32403 (N_32403,N_31701,N_31557);
nor U32404 (N_32404,N_31515,N_31770);
or U32405 (N_32405,N_31688,N_31901);
xnor U32406 (N_32406,N_31810,N_31711);
and U32407 (N_32407,N_31887,N_31695);
nor U32408 (N_32408,N_31828,N_31568);
xor U32409 (N_32409,N_31540,N_31550);
or U32410 (N_32410,N_31856,N_31689);
or U32411 (N_32411,N_31733,N_31531);
or U32412 (N_32412,N_31913,N_31709);
nor U32413 (N_32413,N_31622,N_31789);
xor U32414 (N_32414,N_31966,N_31824);
nor U32415 (N_32415,N_31573,N_31870);
nor U32416 (N_32416,N_31952,N_31812);
nand U32417 (N_32417,N_31938,N_31851);
xor U32418 (N_32418,N_31770,N_31975);
nand U32419 (N_32419,N_31653,N_31996);
nand U32420 (N_32420,N_31734,N_31741);
xnor U32421 (N_32421,N_31916,N_31529);
nor U32422 (N_32422,N_31658,N_31854);
nand U32423 (N_32423,N_31722,N_31962);
and U32424 (N_32424,N_31960,N_31809);
xor U32425 (N_32425,N_31945,N_31675);
nand U32426 (N_32426,N_31994,N_31971);
or U32427 (N_32427,N_31736,N_31789);
nor U32428 (N_32428,N_31781,N_31950);
or U32429 (N_32429,N_31836,N_31714);
xor U32430 (N_32430,N_31701,N_31754);
nand U32431 (N_32431,N_31959,N_31889);
and U32432 (N_32432,N_31671,N_31973);
nor U32433 (N_32433,N_31805,N_31950);
xor U32434 (N_32434,N_31950,N_31843);
and U32435 (N_32435,N_31800,N_31923);
or U32436 (N_32436,N_31942,N_31790);
or U32437 (N_32437,N_31942,N_31634);
xor U32438 (N_32438,N_31917,N_31892);
and U32439 (N_32439,N_31580,N_31746);
nand U32440 (N_32440,N_31689,N_31555);
nor U32441 (N_32441,N_31980,N_31585);
nor U32442 (N_32442,N_31790,N_31545);
and U32443 (N_32443,N_31712,N_31770);
nor U32444 (N_32444,N_31912,N_31925);
nor U32445 (N_32445,N_31598,N_31749);
and U32446 (N_32446,N_31663,N_31628);
nand U32447 (N_32447,N_31700,N_31508);
nor U32448 (N_32448,N_31801,N_31501);
and U32449 (N_32449,N_31762,N_31638);
nand U32450 (N_32450,N_31552,N_31813);
and U32451 (N_32451,N_31640,N_31719);
nor U32452 (N_32452,N_31818,N_31674);
and U32453 (N_32453,N_31700,N_31699);
or U32454 (N_32454,N_31793,N_31624);
or U32455 (N_32455,N_31859,N_31887);
xor U32456 (N_32456,N_31888,N_31831);
and U32457 (N_32457,N_31759,N_31891);
xnor U32458 (N_32458,N_31982,N_31730);
xor U32459 (N_32459,N_31792,N_31681);
nand U32460 (N_32460,N_31548,N_31570);
xor U32461 (N_32461,N_31819,N_31726);
and U32462 (N_32462,N_31700,N_31889);
xor U32463 (N_32463,N_31765,N_31853);
or U32464 (N_32464,N_31789,N_31540);
nand U32465 (N_32465,N_31865,N_31975);
and U32466 (N_32466,N_31524,N_31939);
and U32467 (N_32467,N_31566,N_31553);
or U32468 (N_32468,N_31644,N_31502);
nand U32469 (N_32469,N_31904,N_31872);
nor U32470 (N_32470,N_31597,N_31580);
xor U32471 (N_32471,N_31800,N_31801);
nand U32472 (N_32472,N_31517,N_31775);
and U32473 (N_32473,N_31921,N_31731);
and U32474 (N_32474,N_31803,N_31799);
and U32475 (N_32475,N_31711,N_31738);
and U32476 (N_32476,N_31878,N_31584);
and U32477 (N_32477,N_31913,N_31886);
and U32478 (N_32478,N_31857,N_31956);
xnor U32479 (N_32479,N_31876,N_31999);
or U32480 (N_32480,N_31893,N_31808);
nor U32481 (N_32481,N_31919,N_31886);
nor U32482 (N_32482,N_31534,N_31953);
nand U32483 (N_32483,N_31770,N_31855);
nand U32484 (N_32484,N_31717,N_31869);
nand U32485 (N_32485,N_31604,N_31876);
nand U32486 (N_32486,N_31514,N_31583);
xnor U32487 (N_32487,N_31906,N_31992);
nor U32488 (N_32488,N_31981,N_31861);
or U32489 (N_32489,N_31651,N_31604);
nor U32490 (N_32490,N_31776,N_31932);
xor U32491 (N_32491,N_31935,N_31809);
nor U32492 (N_32492,N_31532,N_31521);
or U32493 (N_32493,N_31621,N_31783);
xnor U32494 (N_32494,N_31853,N_31661);
and U32495 (N_32495,N_31906,N_31522);
xor U32496 (N_32496,N_31675,N_31910);
or U32497 (N_32497,N_31862,N_31726);
and U32498 (N_32498,N_31876,N_31505);
and U32499 (N_32499,N_31795,N_31966);
xnor U32500 (N_32500,N_32273,N_32224);
and U32501 (N_32501,N_32263,N_32089);
nor U32502 (N_32502,N_32158,N_32452);
nand U32503 (N_32503,N_32043,N_32191);
nand U32504 (N_32504,N_32130,N_32105);
or U32505 (N_32505,N_32298,N_32335);
nand U32506 (N_32506,N_32355,N_32482);
xor U32507 (N_32507,N_32210,N_32127);
nor U32508 (N_32508,N_32258,N_32162);
nand U32509 (N_32509,N_32010,N_32341);
or U32510 (N_32510,N_32097,N_32337);
nand U32511 (N_32511,N_32112,N_32478);
nor U32512 (N_32512,N_32290,N_32294);
nand U32513 (N_32513,N_32124,N_32219);
or U32514 (N_32514,N_32070,N_32231);
nor U32515 (N_32515,N_32301,N_32033);
nand U32516 (N_32516,N_32011,N_32340);
nor U32517 (N_32517,N_32023,N_32152);
or U32518 (N_32518,N_32020,N_32206);
and U32519 (N_32519,N_32344,N_32437);
or U32520 (N_32520,N_32017,N_32411);
nand U32521 (N_32521,N_32026,N_32196);
nand U32522 (N_32522,N_32321,N_32299);
or U32523 (N_32523,N_32423,N_32410);
and U32524 (N_32524,N_32399,N_32087);
nor U32525 (N_32525,N_32433,N_32227);
and U32526 (N_32526,N_32028,N_32443);
xor U32527 (N_32527,N_32421,N_32350);
nand U32528 (N_32528,N_32018,N_32412);
xor U32529 (N_32529,N_32377,N_32141);
or U32530 (N_32530,N_32235,N_32498);
nor U32531 (N_32531,N_32048,N_32159);
nor U32532 (N_32532,N_32012,N_32046);
nor U32533 (N_32533,N_32123,N_32137);
xor U32534 (N_32534,N_32110,N_32244);
and U32535 (N_32535,N_32495,N_32040);
xnor U32536 (N_32536,N_32014,N_32462);
xor U32537 (N_32537,N_32236,N_32245);
and U32538 (N_32538,N_32195,N_32133);
or U32539 (N_32539,N_32333,N_32131);
nor U32540 (N_32540,N_32325,N_32115);
nor U32541 (N_32541,N_32473,N_32359);
nor U32542 (N_32542,N_32073,N_32183);
nor U32543 (N_32543,N_32047,N_32078);
nand U32544 (N_32544,N_32438,N_32367);
and U32545 (N_32545,N_32034,N_32042);
nand U32546 (N_32546,N_32172,N_32485);
nor U32547 (N_32547,N_32268,N_32233);
nand U32548 (N_32548,N_32054,N_32353);
xor U32549 (N_32549,N_32390,N_32328);
and U32550 (N_32550,N_32386,N_32025);
xnor U32551 (N_32551,N_32393,N_32487);
xor U32552 (N_32552,N_32488,N_32288);
or U32553 (N_32553,N_32055,N_32489);
xnor U32554 (N_32554,N_32365,N_32392);
nor U32555 (N_32555,N_32310,N_32007);
nor U32556 (N_32556,N_32375,N_32474);
and U32557 (N_32557,N_32378,N_32405);
and U32558 (N_32558,N_32356,N_32376);
and U32559 (N_32559,N_32218,N_32272);
xor U32560 (N_32560,N_32444,N_32456);
or U32561 (N_32561,N_32447,N_32471);
or U32562 (N_32562,N_32160,N_32332);
xnor U32563 (N_32563,N_32135,N_32029);
xnor U32564 (N_32564,N_32209,N_32214);
or U32565 (N_32565,N_32232,N_32429);
nor U32566 (N_32566,N_32408,N_32180);
nor U32567 (N_32567,N_32102,N_32119);
or U32568 (N_32568,N_32181,N_32417);
nand U32569 (N_32569,N_32352,N_32302);
nand U32570 (N_32570,N_32177,N_32414);
nand U32571 (N_32571,N_32292,N_32347);
nor U32572 (N_32572,N_32052,N_32213);
and U32573 (N_32573,N_32253,N_32274);
and U32574 (N_32574,N_32139,N_32212);
nor U32575 (N_32575,N_32469,N_32369);
or U32576 (N_32576,N_32169,N_32136);
nor U32577 (N_32577,N_32220,N_32116);
nand U32578 (N_32578,N_32419,N_32305);
xnor U32579 (N_32579,N_32016,N_32188);
and U32580 (N_32580,N_32389,N_32454);
xor U32581 (N_32581,N_32496,N_32256);
or U32582 (N_32582,N_32255,N_32401);
and U32583 (N_32583,N_32146,N_32458);
xor U32584 (N_32584,N_32186,N_32381);
nand U32585 (N_32585,N_32144,N_32450);
nand U32586 (N_32586,N_32416,N_32491);
or U32587 (N_32587,N_32320,N_32099);
or U32588 (N_32588,N_32430,N_32063);
nand U32589 (N_32589,N_32241,N_32472);
and U32590 (N_32590,N_32251,N_32431);
nand U32591 (N_32591,N_32391,N_32468);
and U32592 (N_32592,N_32126,N_32229);
xnor U32593 (N_32593,N_32327,N_32240);
or U32594 (N_32594,N_32334,N_32064);
and U32595 (N_32595,N_32314,N_32317);
xor U32596 (N_32596,N_32435,N_32051);
xnor U32597 (N_32597,N_32259,N_32326);
xnor U32598 (N_32598,N_32088,N_32425);
and U32599 (N_32599,N_32368,N_32291);
and U32600 (N_32600,N_32465,N_32154);
and U32601 (N_32601,N_32211,N_32217);
xnor U32602 (N_32602,N_32062,N_32380);
xor U32603 (N_32603,N_32164,N_32095);
nor U32604 (N_32604,N_32019,N_32374);
xor U32605 (N_32605,N_32413,N_32499);
nor U32606 (N_32606,N_32364,N_32187);
and U32607 (N_32607,N_32309,N_32013);
or U32608 (N_32608,N_32383,N_32284);
nor U32609 (N_32609,N_32304,N_32059);
xor U32610 (N_32610,N_32426,N_32289);
or U32611 (N_32611,N_32349,N_32319);
xnor U32612 (N_32612,N_32329,N_32009);
or U32613 (N_32613,N_32031,N_32362);
xor U32614 (N_32614,N_32001,N_32203);
or U32615 (N_32615,N_32216,N_32440);
and U32616 (N_32616,N_32202,N_32190);
or U32617 (N_32617,N_32120,N_32422);
or U32618 (N_32618,N_32486,N_32448);
or U32619 (N_32619,N_32453,N_32336);
xnor U32620 (N_32620,N_32371,N_32081);
or U32621 (N_32621,N_32032,N_32082);
or U32622 (N_32622,N_32185,N_32165);
xnor U32623 (N_32623,N_32207,N_32395);
nand U32624 (N_32624,N_32140,N_32113);
or U32625 (N_32625,N_32193,N_32324);
or U32626 (N_32626,N_32125,N_32483);
and U32627 (N_32627,N_32151,N_32134);
or U32628 (N_32628,N_32345,N_32179);
nor U32629 (N_32629,N_32153,N_32111);
xor U32630 (N_32630,N_32357,N_32297);
nor U32631 (N_32631,N_32281,N_32457);
or U32632 (N_32632,N_32295,N_32373);
xor U32633 (N_32633,N_32250,N_32163);
or U32634 (N_32634,N_32223,N_32303);
and U32635 (N_32635,N_32360,N_32024);
and U32636 (N_32636,N_32230,N_32092);
xor U32637 (N_32637,N_32286,N_32149);
and U32638 (N_32638,N_32083,N_32142);
nor U32639 (N_32639,N_32270,N_32418);
nand U32640 (N_32640,N_32323,N_32315);
nand U32641 (N_32641,N_32237,N_32050);
xnor U32642 (N_32642,N_32322,N_32398);
and U32643 (N_32643,N_32008,N_32276);
or U32644 (N_32644,N_32394,N_32293);
nand U32645 (N_32645,N_32461,N_32280);
nand U32646 (N_32646,N_32189,N_32173);
xnor U32647 (N_32647,N_32497,N_32204);
xnor U32648 (N_32648,N_32407,N_32313);
nor U32649 (N_32649,N_32174,N_32260);
or U32650 (N_32650,N_32311,N_32246);
nor U32651 (N_32651,N_32090,N_32198);
nand U32652 (N_32652,N_32106,N_32455);
nand U32653 (N_32653,N_32147,N_32184);
or U32654 (N_32654,N_32100,N_32037);
and U32655 (N_32655,N_32316,N_32069);
xor U32656 (N_32656,N_32201,N_32094);
and U32657 (N_32657,N_32300,N_32072);
xnor U32658 (N_32658,N_32138,N_32222);
xnor U32659 (N_32659,N_32442,N_32065);
nand U32660 (N_32660,N_32282,N_32428);
xnor U32661 (N_32661,N_32271,N_32096);
nand U32662 (N_32662,N_32379,N_32035);
nand U32663 (N_32663,N_32269,N_32058);
or U32664 (N_32664,N_32372,N_32030);
and U32665 (N_32665,N_32021,N_32403);
nand U32666 (N_32666,N_32308,N_32068);
nand U32667 (N_32667,N_32261,N_32118);
and U32668 (N_32668,N_32166,N_32467);
and U32669 (N_32669,N_32148,N_32006);
and U32670 (N_32670,N_32257,N_32117);
and U32671 (N_32671,N_32077,N_32307);
and U32672 (N_32672,N_32109,N_32225);
or U32673 (N_32673,N_32022,N_32346);
nand U32674 (N_32674,N_32348,N_32076);
and U32675 (N_32675,N_32121,N_32312);
or U32676 (N_32676,N_32415,N_32098);
and U32677 (N_32677,N_32406,N_32446);
or U32678 (N_32678,N_32306,N_32464);
nand U32679 (N_32679,N_32239,N_32036);
nand U32680 (N_32680,N_32279,N_32104);
xnor U32681 (N_32681,N_32388,N_32493);
nor U32682 (N_32682,N_32477,N_32404);
or U32683 (N_32683,N_32175,N_32432);
nand U32684 (N_32684,N_32150,N_32358);
or U32685 (N_32685,N_32484,N_32420);
nand U32686 (N_32686,N_32434,N_32242);
nor U32687 (N_32687,N_32132,N_32027);
nand U32688 (N_32688,N_32409,N_32114);
nor U32689 (N_32689,N_32397,N_32205);
nor U32690 (N_32690,N_32044,N_32000);
xnor U32691 (N_32691,N_32330,N_32161);
nand U32692 (N_32692,N_32238,N_32445);
nor U32693 (N_32693,N_32463,N_32157);
or U32694 (N_32694,N_32475,N_32004);
xor U32695 (N_32695,N_32400,N_32192);
nor U32696 (N_32696,N_32427,N_32066);
nor U32697 (N_32697,N_32075,N_32122);
nor U32698 (N_32698,N_32451,N_32003);
and U32699 (N_32699,N_32167,N_32128);
or U32700 (N_32700,N_32490,N_32296);
nand U32701 (N_32701,N_32176,N_32199);
nor U32702 (N_32702,N_32396,N_32366);
nand U32703 (N_32703,N_32277,N_32361);
nor U32704 (N_32704,N_32339,N_32285);
and U32705 (N_32705,N_32056,N_32178);
nor U32706 (N_32706,N_32226,N_32479);
xnor U32707 (N_32707,N_32424,N_32108);
nand U32708 (N_32708,N_32060,N_32171);
and U32709 (N_32709,N_32145,N_32264);
xor U32710 (N_32710,N_32200,N_32143);
and U32711 (N_32711,N_32079,N_32208);
xor U32712 (N_32712,N_32005,N_32170);
nand U32713 (N_32713,N_32283,N_32382);
nand U32714 (N_32714,N_32041,N_32038);
nand U32715 (N_32715,N_32074,N_32039);
xor U32716 (N_32716,N_32091,N_32459);
nand U32717 (N_32717,N_32370,N_32228);
nand U32718 (N_32718,N_32002,N_32387);
nand U32719 (N_32719,N_32182,N_32287);
nor U32720 (N_32720,N_32221,N_32278);
xor U32721 (N_32721,N_32338,N_32085);
nand U32722 (N_32722,N_32441,N_32103);
nor U32723 (N_32723,N_32266,N_32243);
nor U32724 (N_32724,N_32481,N_32234);
and U32725 (N_32725,N_32343,N_32086);
nand U32726 (N_32726,N_32057,N_32215);
nand U32727 (N_32727,N_32067,N_32331);
or U32728 (N_32728,N_32061,N_32053);
and U32729 (N_32729,N_32354,N_32107);
nor U32730 (N_32730,N_32249,N_32247);
and U32731 (N_32731,N_32470,N_32248);
nor U32732 (N_32732,N_32129,N_32480);
and U32733 (N_32733,N_32252,N_32080);
and U32734 (N_32734,N_32476,N_32197);
or U32735 (N_32735,N_32436,N_32084);
xor U32736 (N_32736,N_32015,N_32267);
xnor U32737 (N_32737,N_32194,N_32254);
nor U32738 (N_32738,N_32384,N_32049);
and U32739 (N_32739,N_32351,N_32439);
nand U32740 (N_32740,N_32460,N_32385);
and U32741 (N_32741,N_32466,N_32093);
or U32742 (N_32742,N_32071,N_32402);
nor U32743 (N_32743,N_32265,N_32492);
nand U32744 (N_32744,N_32342,N_32363);
nor U32745 (N_32745,N_32262,N_32155);
xor U32746 (N_32746,N_32168,N_32449);
and U32747 (N_32747,N_32275,N_32045);
and U32748 (N_32748,N_32156,N_32101);
xor U32749 (N_32749,N_32318,N_32494);
and U32750 (N_32750,N_32059,N_32041);
and U32751 (N_32751,N_32425,N_32285);
nand U32752 (N_32752,N_32441,N_32132);
or U32753 (N_32753,N_32468,N_32016);
xnor U32754 (N_32754,N_32263,N_32354);
xor U32755 (N_32755,N_32320,N_32054);
and U32756 (N_32756,N_32198,N_32037);
or U32757 (N_32757,N_32095,N_32273);
and U32758 (N_32758,N_32464,N_32378);
nor U32759 (N_32759,N_32152,N_32310);
nor U32760 (N_32760,N_32030,N_32203);
or U32761 (N_32761,N_32025,N_32413);
xnor U32762 (N_32762,N_32345,N_32288);
xnor U32763 (N_32763,N_32364,N_32352);
xor U32764 (N_32764,N_32300,N_32192);
nand U32765 (N_32765,N_32301,N_32455);
and U32766 (N_32766,N_32372,N_32287);
or U32767 (N_32767,N_32336,N_32063);
xnor U32768 (N_32768,N_32478,N_32135);
xor U32769 (N_32769,N_32255,N_32406);
and U32770 (N_32770,N_32188,N_32415);
and U32771 (N_32771,N_32427,N_32364);
and U32772 (N_32772,N_32243,N_32014);
nor U32773 (N_32773,N_32466,N_32357);
nor U32774 (N_32774,N_32271,N_32275);
xor U32775 (N_32775,N_32202,N_32295);
xor U32776 (N_32776,N_32484,N_32010);
nor U32777 (N_32777,N_32353,N_32430);
nand U32778 (N_32778,N_32162,N_32418);
xor U32779 (N_32779,N_32444,N_32451);
xnor U32780 (N_32780,N_32287,N_32220);
and U32781 (N_32781,N_32021,N_32387);
or U32782 (N_32782,N_32218,N_32216);
nand U32783 (N_32783,N_32172,N_32249);
nor U32784 (N_32784,N_32276,N_32428);
nand U32785 (N_32785,N_32481,N_32025);
or U32786 (N_32786,N_32100,N_32242);
and U32787 (N_32787,N_32055,N_32488);
nand U32788 (N_32788,N_32403,N_32427);
and U32789 (N_32789,N_32477,N_32378);
or U32790 (N_32790,N_32468,N_32321);
xor U32791 (N_32791,N_32151,N_32286);
xor U32792 (N_32792,N_32318,N_32042);
xor U32793 (N_32793,N_32125,N_32407);
or U32794 (N_32794,N_32178,N_32317);
and U32795 (N_32795,N_32423,N_32166);
and U32796 (N_32796,N_32233,N_32176);
nand U32797 (N_32797,N_32305,N_32492);
and U32798 (N_32798,N_32110,N_32264);
xor U32799 (N_32799,N_32448,N_32445);
or U32800 (N_32800,N_32266,N_32333);
or U32801 (N_32801,N_32046,N_32417);
or U32802 (N_32802,N_32217,N_32253);
xor U32803 (N_32803,N_32283,N_32197);
nor U32804 (N_32804,N_32259,N_32467);
xor U32805 (N_32805,N_32300,N_32151);
nor U32806 (N_32806,N_32058,N_32194);
or U32807 (N_32807,N_32402,N_32301);
nor U32808 (N_32808,N_32467,N_32363);
or U32809 (N_32809,N_32078,N_32081);
xnor U32810 (N_32810,N_32372,N_32430);
nand U32811 (N_32811,N_32449,N_32294);
nand U32812 (N_32812,N_32024,N_32211);
or U32813 (N_32813,N_32266,N_32364);
or U32814 (N_32814,N_32369,N_32432);
and U32815 (N_32815,N_32423,N_32418);
or U32816 (N_32816,N_32099,N_32179);
or U32817 (N_32817,N_32466,N_32342);
nand U32818 (N_32818,N_32406,N_32489);
or U32819 (N_32819,N_32334,N_32090);
or U32820 (N_32820,N_32125,N_32448);
nand U32821 (N_32821,N_32337,N_32466);
nor U32822 (N_32822,N_32049,N_32178);
nor U32823 (N_32823,N_32266,N_32442);
and U32824 (N_32824,N_32280,N_32222);
and U32825 (N_32825,N_32038,N_32457);
nand U32826 (N_32826,N_32449,N_32351);
nor U32827 (N_32827,N_32434,N_32120);
nand U32828 (N_32828,N_32353,N_32322);
or U32829 (N_32829,N_32271,N_32238);
nand U32830 (N_32830,N_32449,N_32148);
or U32831 (N_32831,N_32355,N_32122);
and U32832 (N_32832,N_32073,N_32262);
nand U32833 (N_32833,N_32440,N_32258);
or U32834 (N_32834,N_32400,N_32071);
and U32835 (N_32835,N_32109,N_32245);
and U32836 (N_32836,N_32209,N_32451);
nor U32837 (N_32837,N_32347,N_32498);
and U32838 (N_32838,N_32253,N_32300);
nand U32839 (N_32839,N_32338,N_32373);
nor U32840 (N_32840,N_32360,N_32410);
or U32841 (N_32841,N_32115,N_32445);
and U32842 (N_32842,N_32171,N_32116);
nor U32843 (N_32843,N_32009,N_32288);
nand U32844 (N_32844,N_32471,N_32085);
nand U32845 (N_32845,N_32265,N_32090);
nor U32846 (N_32846,N_32484,N_32341);
nor U32847 (N_32847,N_32188,N_32438);
or U32848 (N_32848,N_32396,N_32076);
xnor U32849 (N_32849,N_32259,N_32179);
xor U32850 (N_32850,N_32243,N_32101);
nand U32851 (N_32851,N_32047,N_32174);
nand U32852 (N_32852,N_32352,N_32008);
and U32853 (N_32853,N_32369,N_32447);
nor U32854 (N_32854,N_32284,N_32174);
xnor U32855 (N_32855,N_32430,N_32297);
xnor U32856 (N_32856,N_32469,N_32328);
xnor U32857 (N_32857,N_32229,N_32312);
or U32858 (N_32858,N_32032,N_32493);
nand U32859 (N_32859,N_32111,N_32004);
nand U32860 (N_32860,N_32495,N_32377);
and U32861 (N_32861,N_32031,N_32155);
nor U32862 (N_32862,N_32310,N_32395);
nand U32863 (N_32863,N_32479,N_32266);
nor U32864 (N_32864,N_32005,N_32086);
xor U32865 (N_32865,N_32380,N_32205);
nor U32866 (N_32866,N_32183,N_32163);
nand U32867 (N_32867,N_32461,N_32305);
nor U32868 (N_32868,N_32116,N_32085);
xor U32869 (N_32869,N_32389,N_32090);
nor U32870 (N_32870,N_32257,N_32358);
xnor U32871 (N_32871,N_32330,N_32409);
xor U32872 (N_32872,N_32211,N_32000);
xor U32873 (N_32873,N_32007,N_32136);
or U32874 (N_32874,N_32498,N_32205);
or U32875 (N_32875,N_32229,N_32172);
xnor U32876 (N_32876,N_32396,N_32041);
or U32877 (N_32877,N_32037,N_32230);
and U32878 (N_32878,N_32362,N_32049);
or U32879 (N_32879,N_32277,N_32172);
nand U32880 (N_32880,N_32309,N_32330);
xnor U32881 (N_32881,N_32268,N_32335);
nor U32882 (N_32882,N_32016,N_32341);
or U32883 (N_32883,N_32213,N_32220);
nor U32884 (N_32884,N_32369,N_32049);
nand U32885 (N_32885,N_32206,N_32243);
xor U32886 (N_32886,N_32249,N_32336);
and U32887 (N_32887,N_32329,N_32081);
nand U32888 (N_32888,N_32077,N_32102);
or U32889 (N_32889,N_32496,N_32393);
or U32890 (N_32890,N_32385,N_32410);
xnor U32891 (N_32891,N_32087,N_32412);
nor U32892 (N_32892,N_32009,N_32113);
xnor U32893 (N_32893,N_32268,N_32411);
nand U32894 (N_32894,N_32105,N_32071);
nand U32895 (N_32895,N_32300,N_32296);
and U32896 (N_32896,N_32033,N_32455);
nand U32897 (N_32897,N_32059,N_32397);
nand U32898 (N_32898,N_32475,N_32194);
xor U32899 (N_32899,N_32293,N_32224);
nor U32900 (N_32900,N_32070,N_32384);
nor U32901 (N_32901,N_32040,N_32375);
and U32902 (N_32902,N_32359,N_32028);
xnor U32903 (N_32903,N_32242,N_32295);
and U32904 (N_32904,N_32155,N_32405);
nand U32905 (N_32905,N_32064,N_32148);
and U32906 (N_32906,N_32132,N_32442);
or U32907 (N_32907,N_32130,N_32063);
nand U32908 (N_32908,N_32470,N_32028);
nand U32909 (N_32909,N_32428,N_32080);
or U32910 (N_32910,N_32192,N_32167);
nor U32911 (N_32911,N_32211,N_32089);
nor U32912 (N_32912,N_32238,N_32380);
and U32913 (N_32913,N_32349,N_32031);
nor U32914 (N_32914,N_32282,N_32413);
xor U32915 (N_32915,N_32159,N_32370);
nand U32916 (N_32916,N_32342,N_32256);
nor U32917 (N_32917,N_32281,N_32477);
and U32918 (N_32918,N_32490,N_32083);
and U32919 (N_32919,N_32089,N_32330);
and U32920 (N_32920,N_32027,N_32486);
and U32921 (N_32921,N_32208,N_32479);
or U32922 (N_32922,N_32077,N_32075);
or U32923 (N_32923,N_32063,N_32081);
or U32924 (N_32924,N_32087,N_32035);
nor U32925 (N_32925,N_32033,N_32322);
or U32926 (N_32926,N_32059,N_32156);
nor U32927 (N_32927,N_32359,N_32289);
xor U32928 (N_32928,N_32065,N_32110);
nor U32929 (N_32929,N_32320,N_32048);
nor U32930 (N_32930,N_32497,N_32215);
and U32931 (N_32931,N_32188,N_32257);
nor U32932 (N_32932,N_32431,N_32294);
and U32933 (N_32933,N_32430,N_32378);
and U32934 (N_32934,N_32353,N_32284);
nor U32935 (N_32935,N_32226,N_32441);
nand U32936 (N_32936,N_32300,N_32480);
nor U32937 (N_32937,N_32383,N_32260);
xnor U32938 (N_32938,N_32184,N_32405);
nor U32939 (N_32939,N_32206,N_32459);
nand U32940 (N_32940,N_32116,N_32392);
nor U32941 (N_32941,N_32232,N_32015);
or U32942 (N_32942,N_32198,N_32275);
nor U32943 (N_32943,N_32106,N_32119);
xor U32944 (N_32944,N_32303,N_32008);
nor U32945 (N_32945,N_32067,N_32269);
nand U32946 (N_32946,N_32456,N_32110);
nand U32947 (N_32947,N_32236,N_32046);
nand U32948 (N_32948,N_32463,N_32282);
xnor U32949 (N_32949,N_32490,N_32478);
and U32950 (N_32950,N_32266,N_32480);
nor U32951 (N_32951,N_32199,N_32104);
and U32952 (N_32952,N_32311,N_32180);
and U32953 (N_32953,N_32342,N_32423);
or U32954 (N_32954,N_32493,N_32332);
and U32955 (N_32955,N_32496,N_32171);
xnor U32956 (N_32956,N_32312,N_32231);
or U32957 (N_32957,N_32344,N_32302);
or U32958 (N_32958,N_32390,N_32242);
xor U32959 (N_32959,N_32334,N_32091);
xor U32960 (N_32960,N_32326,N_32126);
nand U32961 (N_32961,N_32169,N_32002);
or U32962 (N_32962,N_32478,N_32069);
nand U32963 (N_32963,N_32021,N_32293);
xor U32964 (N_32964,N_32381,N_32071);
nand U32965 (N_32965,N_32320,N_32094);
nor U32966 (N_32966,N_32384,N_32467);
nand U32967 (N_32967,N_32292,N_32152);
nor U32968 (N_32968,N_32250,N_32188);
nor U32969 (N_32969,N_32242,N_32417);
nand U32970 (N_32970,N_32307,N_32039);
and U32971 (N_32971,N_32330,N_32317);
and U32972 (N_32972,N_32469,N_32167);
nand U32973 (N_32973,N_32308,N_32298);
nor U32974 (N_32974,N_32020,N_32276);
nand U32975 (N_32975,N_32331,N_32076);
nand U32976 (N_32976,N_32025,N_32498);
nor U32977 (N_32977,N_32130,N_32155);
and U32978 (N_32978,N_32314,N_32285);
or U32979 (N_32979,N_32245,N_32372);
xor U32980 (N_32980,N_32043,N_32365);
nand U32981 (N_32981,N_32407,N_32048);
nand U32982 (N_32982,N_32212,N_32127);
nand U32983 (N_32983,N_32343,N_32265);
nand U32984 (N_32984,N_32240,N_32298);
or U32985 (N_32985,N_32449,N_32216);
xor U32986 (N_32986,N_32149,N_32252);
xor U32987 (N_32987,N_32278,N_32144);
nand U32988 (N_32988,N_32182,N_32051);
nor U32989 (N_32989,N_32440,N_32003);
xor U32990 (N_32990,N_32324,N_32080);
xnor U32991 (N_32991,N_32084,N_32018);
nand U32992 (N_32992,N_32413,N_32142);
or U32993 (N_32993,N_32105,N_32160);
nor U32994 (N_32994,N_32266,N_32444);
nand U32995 (N_32995,N_32141,N_32057);
nand U32996 (N_32996,N_32482,N_32392);
or U32997 (N_32997,N_32429,N_32443);
nor U32998 (N_32998,N_32462,N_32364);
xnor U32999 (N_32999,N_32471,N_32339);
nor U33000 (N_33000,N_32746,N_32725);
nor U33001 (N_33001,N_32567,N_32608);
xnor U33002 (N_33002,N_32989,N_32906);
xnor U33003 (N_33003,N_32855,N_32831);
and U33004 (N_33004,N_32687,N_32794);
xnor U33005 (N_33005,N_32867,N_32510);
xnor U33006 (N_33006,N_32557,N_32916);
xnor U33007 (N_33007,N_32684,N_32930);
nand U33008 (N_33008,N_32934,N_32620);
nand U33009 (N_33009,N_32627,N_32683);
or U33010 (N_33010,N_32897,N_32727);
xor U33011 (N_33011,N_32830,N_32880);
xnor U33012 (N_33012,N_32913,N_32709);
nor U33013 (N_33013,N_32730,N_32507);
or U33014 (N_33014,N_32543,N_32614);
or U33015 (N_33015,N_32811,N_32589);
or U33016 (N_33016,N_32740,N_32792);
nor U33017 (N_33017,N_32566,N_32766);
and U33018 (N_33018,N_32849,N_32938);
nand U33019 (N_33019,N_32999,N_32569);
or U33020 (N_33020,N_32837,N_32806);
xnor U33021 (N_33021,N_32739,N_32895);
nor U33022 (N_33022,N_32713,N_32749);
nand U33023 (N_33023,N_32904,N_32752);
nand U33024 (N_33024,N_32969,N_32685);
xnor U33025 (N_33025,N_32777,N_32733);
and U33026 (N_33026,N_32672,N_32692);
nor U33027 (N_33027,N_32943,N_32609);
nor U33028 (N_33028,N_32521,N_32558);
xor U33029 (N_33029,N_32563,N_32844);
nor U33030 (N_33030,N_32773,N_32705);
nand U33031 (N_33031,N_32535,N_32856);
xnor U33032 (N_33032,N_32581,N_32762);
and U33033 (N_33033,N_32861,N_32976);
or U33034 (N_33034,N_32908,N_32812);
xor U33035 (N_33035,N_32872,N_32869);
nand U33036 (N_33036,N_32610,N_32522);
and U33037 (N_33037,N_32808,N_32952);
xor U33038 (N_33038,N_32513,N_32530);
xor U33039 (N_33039,N_32506,N_32526);
nor U33040 (N_33040,N_32954,N_32886);
nor U33041 (N_33041,N_32742,N_32764);
nor U33042 (N_33042,N_32915,N_32681);
or U33043 (N_33043,N_32654,N_32927);
and U33044 (N_33044,N_32560,N_32774);
xnor U33045 (N_33045,N_32864,N_32926);
xnor U33046 (N_33046,N_32590,N_32673);
and U33047 (N_33047,N_32592,N_32997);
xnor U33048 (N_33048,N_32708,N_32508);
nor U33049 (N_33049,N_32720,N_32655);
nand U33050 (N_33050,N_32944,N_32760);
nand U33051 (N_33051,N_32948,N_32718);
or U33052 (N_33052,N_32652,N_32527);
nor U33053 (N_33053,N_32518,N_32755);
and U33054 (N_33054,N_32611,N_32647);
nor U33055 (N_33055,N_32584,N_32786);
xnor U33056 (N_33056,N_32676,N_32554);
and U33057 (N_33057,N_32981,N_32853);
xnor U33058 (N_33058,N_32545,N_32827);
nand U33059 (N_33059,N_32605,N_32975);
nor U33060 (N_33060,N_32784,N_32912);
nor U33061 (N_33061,N_32751,N_32795);
or U33062 (N_33062,N_32633,N_32631);
and U33063 (N_33063,N_32516,N_32588);
nor U33064 (N_33064,N_32628,N_32531);
xnor U33065 (N_33065,N_32556,N_32715);
or U33066 (N_33066,N_32754,N_32737);
xor U33067 (N_33067,N_32935,N_32859);
nor U33068 (N_33068,N_32818,N_32619);
nor U33069 (N_33069,N_32538,N_32578);
and U33070 (N_33070,N_32971,N_32962);
nand U33071 (N_33071,N_32559,N_32536);
and U33072 (N_33072,N_32911,N_32514);
nor U33073 (N_33073,N_32712,N_32781);
nand U33074 (N_33074,N_32960,N_32843);
or U33075 (N_33075,N_32940,N_32574);
and U33076 (N_33076,N_32591,N_32984);
nand U33077 (N_33077,N_32656,N_32579);
and U33078 (N_33078,N_32565,N_32642);
and U33079 (N_33079,N_32653,N_32788);
or U33080 (N_33080,N_32964,N_32729);
xnor U33081 (N_33081,N_32801,N_32947);
and U33082 (N_33082,N_32544,N_32779);
and U33083 (N_33083,N_32803,N_32946);
or U33084 (N_33084,N_32970,N_32957);
and U33085 (N_33085,N_32874,N_32929);
nand U33086 (N_33086,N_32896,N_32677);
or U33087 (N_33087,N_32887,N_32641);
xnor U33088 (N_33088,N_32866,N_32978);
xor U33089 (N_33089,N_32548,N_32520);
nor U33090 (N_33090,N_32986,N_32679);
nor U33091 (N_33091,N_32881,N_32601);
nor U33092 (N_33092,N_32695,N_32738);
nor U33093 (N_33093,N_32987,N_32840);
nand U33094 (N_33094,N_32992,N_32615);
xor U33095 (N_33095,N_32649,N_32778);
nor U33096 (N_33096,N_32731,N_32857);
xnor U33097 (N_33097,N_32595,N_32854);
and U33098 (N_33098,N_32748,N_32828);
and U33099 (N_33099,N_32898,N_32821);
or U33100 (N_33100,N_32597,N_32848);
nor U33101 (N_33101,N_32789,N_32838);
and U33102 (N_33102,N_32814,N_32763);
and U33103 (N_33103,N_32988,N_32757);
or U33104 (N_33104,N_32617,N_32686);
or U33105 (N_33105,N_32706,N_32575);
nor U33106 (N_33106,N_32734,N_32551);
nor U33107 (N_33107,N_32618,N_32674);
and U33108 (N_33108,N_32745,N_32953);
or U33109 (N_33109,N_32613,N_32793);
xnor U33110 (N_33110,N_32823,N_32502);
and U33111 (N_33111,N_32798,N_32753);
nor U33112 (N_33112,N_32555,N_32771);
or U33113 (N_33113,N_32638,N_32996);
nand U33114 (N_33114,N_32645,N_32723);
nor U33115 (N_33115,N_32825,N_32702);
or U33116 (N_33116,N_32782,N_32663);
or U33117 (N_33117,N_32750,N_32517);
and U33118 (N_33118,N_32961,N_32624);
or U33119 (N_33119,N_32657,N_32876);
or U33120 (N_33120,N_32743,N_32691);
or U33121 (N_33121,N_32602,N_32598);
xor U33122 (N_33122,N_32668,N_32509);
nor U33123 (N_33123,N_32758,N_32995);
nor U33124 (N_33124,N_32586,N_32888);
xnor U33125 (N_33125,N_32910,N_32503);
and U33126 (N_33126,N_32639,N_32650);
xor U33127 (N_33127,N_32918,N_32993);
nor U33128 (N_33128,N_32939,N_32634);
nor U33129 (N_33129,N_32907,N_32924);
xor U33130 (N_33130,N_32824,N_32860);
or U33131 (N_33131,N_32625,N_32770);
or U33132 (N_33132,N_32973,N_32928);
nor U33133 (N_33133,N_32549,N_32966);
nand U33134 (N_33134,N_32571,N_32902);
and U33135 (N_33135,N_32630,N_32768);
nor U33136 (N_33136,N_32726,N_32865);
nor U33137 (N_33137,N_32919,N_32846);
xor U33138 (N_33138,N_32863,N_32925);
or U33139 (N_33139,N_32658,N_32621);
nand U33140 (N_33140,N_32523,N_32796);
nand U33141 (N_33141,N_32802,N_32546);
or U33142 (N_33142,N_32659,N_32694);
or U33143 (N_33143,N_32921,N_32965);
xor U33144 (N_33144,N_32504,N_32985);
or U33145 (N_33145,N_32716,N_32599);
or U33146 (N_33146,N_32829,N_32807);
or U33147 (N_33147,N_32698,N_32660);
xnor U33148 (N_33148,N_32756,N_32537);
xnor U33149 (N_33149,N_32871,N_32607);
nor U33150 (N_33150,N_32622,N_32810);
xor U33151 (N_33151,N_32573,N_32682);
nand U33152 (N_33152,N_32553,N_32882);
nand U33153 (N_33153,N_32835,N_32878);
nor U33154 (N_33154,N_32815,N_32626);
or U33155 (N_33155,N_32552,N_32651);
or U33156 (N_33156,N_32822,N_32899);
and U33157 (N_33157,N_32524,N_32767);
xnor U33158 (N_33158,N_32665,N_32945);
nor U33159 (N_33159,N_32998,N_32532);
nand U33160 (N_33160,N_32923,N_32889);
xor U33161 (N_33161,N_32690,N_32805);
and U33162 (N_33162,N_32596,N_32670);
xor U33163 (N_33163,N_32955,N_32636);
xnor U33164 (N_33164,N_32703,N_32540);
and U33165 (N_33165,N_32977,N_32775);
nor U33166 (N_33166,N_32951,N_32879);
nor U33167 (N_33167,N_32847,N_32675);
and U33168 (N_33168,N_32759,N_32697);
nand U33169 (N_33169,N_32606,N_32547);
nor U33170 (N_33170,N_32950,N_32858);
or U33171 (N_33171,N_32600,N_32826);
and U33172 (N_33172,N_32900,N_32541);
or U33173 (N_33173,N_32862,N_32909);
or U33174 (N_33174,N_32587,N_32870);
xnor U33175 (N_33175,N_32505,N_32917);
or U33176 (N_33176,N_32983,N_32732);
or U33177 (N_33177,N_32834,N_32512);
xor U33178 (N_33178,N_32956,N_32972);
nor U33179 (N_33179,N_32920,N_32936);
or U33180 (N_33180,N_32582,N_32785);
nand U33181 (N_33181,N_32868,N_32696);
and U33182 (N_33182,N_32885,N_32688);
and U33183 (N_33183,N_32884,N_32680);
and U33184 (N_33184,N_32643,N_32741);
nor U33185 (N_33185,N_32851,N_32905);
and U33186 (N_33186,N_32577,N_32744);
xor U33187 (N_33187,N_32800,N_32721);
xnor U33188 (N_33188,N_32894,N_32850);
xor U33189 (N_33189,N_32875,N_32765);
and U33190 (N_33190,N_32903,N_32717);
xnor U33191 (N_33191,N_32772,N_32728);
nand U33192 (N_33192,N_32664,N_32883);
and U33193 (N_33193,N_32714,N_32736);
nor U33194 (N_33194,N_32817,N_32891);
xnor U33195 (N_33195,N_32809,N_32994);
or U33196 (N_33196,N_32699,N_32700);
nand U33197 (N_33197,N_32593,N_32932);
or U33198 (N_33198,N_32852,N_32667);
or U33199 (N_33199,N_32776,N_32949);
or U33200 (N_33200,N_32500,N_32790);
nand U33201 (N_33201,N_32974,N_32922);
nor U33202 (N_33202,N_32813,N_32635);
nand U33203 (N_33203,N_32542,N_32550);
nand U33204 (N_33204,N_32832,N_32933);
nand U33205 (N_33205,N_32991,N_32604);
nor U33206 (N_33206,N_32661,N_32515);
or U33207 (N_33207,N_32662,N_32982);
xor U33208 (N_33208,N_32724,N_32959);
nor U33209 (N_33209,N_32873,N_32761);
or U33210 (N_33210,N_32839,N_32570);
nand U33211 (N_33211,N_32511,N_32783);
or U33212 (N_33212,N_32845,N_32693);
nand U33213 (N_33213,N_32877,N_32958);
or U33214 (N_33214,N_32820,N_32722);
and U33215 (N_33215,N_32842,N_32890);
nand U33216 (N_33216,N_32678,N_32819);
nand U33217 (N_33217,N_32623,N_32564);
xor U33218 (N_33218,N_32735,N_32585);
xnor U33219 (N_33219,N_32594,N_32671);
and U33220 (N_33220,N_32640,N_32576);
nor U33221 (N_33221,N_32747,N_32704);
nor U33222 (N_33222,N_32804,N_32666);
xor U33223 (N_33223,N_32841,N_32787);
or U33224 (N_33224,N_32603,N_32769);
nor U33225 (N_33225,N_32968,N_32833);
xnor U33226 (N_33226,N_32963,N_32710);
or U33227 (N_33227,N_32616,N_32836);
xor U33228 (N_33228,N_32533,N_32701);
or U33229 (N_33229,N_32637,N_32632);
xnor U33230 (N_33230,N_32669,N_32525);
nand U33231 (N_33231,N_32561,N_32572);
or U33232 (N_33232,N_32980,N_32901);
nand U33233 (N_33233,N_32612,N_32914);
and U33234 (N_33234,N_32707,N_32501);
nor U33235 (N_33235,N_32937,N_32519);
xnor U33236 (N_33236,N_32629,N_32990);
xor U33237 (N_33237,N_32711,N_32797);
xor U33238 (N_33238,N_32799,N_32719);
nor U33239 (N_33239,N_32562,N_32791);
or U33240 (N_33240,N_32893,N_32942);
xnor U33241 (N_33241,N_32689,N_32580);
xnor U33242 (N_33242,N_32644,N_32967);
xnor U33243 (N_33243,N_32648,N_32529);
and U33244 (N_33244,N_32780,N_32931);
nor U33245 (N_33245,N_32583,N_32892);
nor U33246 (N_33246,N_32941,N_32979);
xnor U33247 (N_33247,N_32568,N_32528);
and U33248 (N_33248,N_32816,N_32534);
xor U33249 (N_33249,N_32646,N_32539);
nand U33250 (N_33250,N_32547,N_32509);
nand U33251 (N_33251,N_32953,N_32789);
nor U33252 (N_33252,N_32716,N_32649);
or U33253 (N_33253,N_32941,N_32812);
and U33254 (N_33254,N_32930,N_32949);
xnor U33255 (N_33255,N_32887,N_32875);
or U33256 (N_33256,N_32516,N_32795);
nor U33257 (N_33257,N_32761,N_32829);
nor U33258 (N_33258,N_32693,N_32748);
xor U33259 (N_33259,N_32837,N_32564);
and U33260 (N_33260,N_32682,N_32882);
or U33261 (N_33261,N_32721,N_32999);
or U33262 (N_33262,N_32735,N_32883);
xnor U33263 (N_33263,N_32669,N_32556);
xnor U33264 (N_33264,N_32990,N_32972);
or U33265 (N_33265,N_32888,N_32794);
xor U33266 (N_33266,N_32547,N_32926);
xnor U33267 (N_33267,N_32696,N_32939);
or U33268 (N_33268,N_32693,N_32777);
nor U33269 (N_33269,N_32521,N_32862);
and U33270 (N_33270,N_32722,N_32530);
nor U33271 (N_33271,N_32882,N_32797);
xor U33272 (N_33272,N_32849,N_32726);
or U33273 (N_33273,N_32764,N_32563);
nor U33274 (N_33274,N_32571,N_32857);
and U33275 (N_33275,N_32508,N_32866);
nand U33276 (N_33276,N_32991,N_32683);
nand U33277 (N_33277,N_32954,N_32743);
or U33278 (N_33278,N_32835,N_32904);
and U33279 (N_33279,N_32555,N_32641);
or U33280 (N_33280,N_32737,N_32986);
or U33281 (N_33281,N_32841,N_32595);
and U33282 (N_33282,N_32874,N_32940);
or U33283 (N_33283,N_32553,N_32509);
xor U33284 (N_33284,N_32942,N_32583);
nand U33285 (N_33285,N_32625,N_32693);
nor U33286 (N_33286,N_32808,N_32508);
nand U33287 (N_33287,N_32730,N_32566);
and U33288 (N_33288,N_32704,N_32680);
and U33289 (N_33289,N_32749,N_32695);
and U33290 (N_33290,N_32655,N_32928);
nor U33291 (N_33291,N_32816,N_32678);
nor U33292 (N_33292,N_32953,N_32604);
xnor U33293 (N_33293,N_32901,N_32804);
or U33294 (N_33294,N_32653,N_32892);
and U33295 (N_33295,N_32807,N_32874);
and U33296 (N_33296,N_32530,N_32578);
xnor U33297 (N_33297,N_32994,N_32713);
or U33298 (N_33298,N_32775,N_32979);
xor U33299 (N_33299,N_32739,N_32690);
xor U33300 (N_33300,N_32918,N_32924);
and U33301 (N_33301,N_32859,N_32996);
nand U33302 (N_33302,N_32551,N_32683);
and U33303 (N_33303,N_32920,N_32988);
nand U33304 (N_33304,N_32541,N_32998);
xor U33305 (N_33305,N_32793,N_32820);
nand U33306 (N_33306,N_32844,N_32961);
or U33307 (N_33307,N_32959,N_32682);
or U33308 (N_33308,N_32952,N_32843);
nand U33309 (N_33309,N_32771,N_32936);
or U33310 (N_33310,N_32874,N_32837);
or U33311 (N_33311,N_32606,N_32748);
or U33312 (N_33312,N_32545,N_32855);
nor U33313 (N_33313,N_32751,N_32880);
nand U33314 (N_33314,N_32650,N_32826);
or U33315 (N_33315,N_32863,N_32786);
nand U33316 (N_33316,N_32751,N_32827);
or U33317 (N_33317,N_32947,N_32886);
nand U33318 (N_33318,N_32915,N_32512);
and U33319 (N_33319,N_32721,N_32838);
xor U33320 (N_33320,N_32872,N_32959);
nor U33321 (N_33321,N_32726,N_32519);
nor U33322 (N_33322,N_32941,N_32673);
or U33323 (N_33323,N_32675,N_32808);
xor U33324 (N_33324,N_32691,N_32775);
and U33325 (N_33325,N_32861,N_32704);
nand U33326 (N_33326,N_32958,N_32529);
nand U33327 (N_33327,N_32582,N_32979);
xnor U33328 (N_33328,N_32735,N_32940);
nand U33329 (N_33329,N_32557,N_32744);
and U33330 (N_33330,N_32895,N_32622);
nor U33331 (N_33331,N_32955,N_32651);
or U33332 (N_33332,N_32598,N_32632);
nor U33333 (N_33333,N_32919,N_32931);
and U33334 (N_33334,N_32728,N_32536);
or U33335 (N_33335,N_32790,N_32900);
nor U33336 (N_33336,N_32923,N_32503);
nand U33337 (N_33337,N_32926,N_32561);
and U33338 (N_33338,N_32700,N_32694);
and U33339 (N_33339,N_32695,N_32505);
nand U33340 (N_33340,N_32702,N_32989);
and U33341 (N_33341,N_32635,N_32531);
nand U33342 (N_33342,N_32639,N_32950);
or U33343 (N_33343,N_32817,N_32834);
nor U33344 (N_33344,N_32940,N_32730);
nand U33345 (N_33345,N_32922,N_32637);
nand U33346 (N_33346,N_32517,N_32636);
and U33347 (N_33347,N_32545,N_32509);
or U33348 (N_33348,N_32825,N_32920);
and U33349 (N_33349,N_32878,N_32829);
nor U33350 (N_33350,N_32977,N_32794);
and U33351 (N_33351,N_32628,N_32728);
xor U33352 (N_33352,N_32699,N_32924);
xnor U33353 (N_33353,N_32865,N_32805);
nand U33354 (N_33354,N_32616,N_32571);
and U33355 (N_33355,N_32653,N_32829);
and U33356 (N_33356,N_32586,N_32606);
xor U33357 (N_33357,N_32532,N_32937);
or U33358 (N_33358,N_32985,N_32828);
nor U33359 (N_33359,N_32800,N_32774);
xnor U33360 (N_33360,N_32573,N_32537);
or U33361 (N_33361,N_32868,N_32573);
nand U33362 (N_33362,N_32948,N_32919);
nor U33363 (N_33363,N_32827,N_32671);
nor U33364 (N_33364,N_32557,N_32516);
xnor U33365 (N_33365,N_32827,N_32513);
and U33366 (N_33366,N_32912,N_32515);
and U33367 (N_33367,N_32834,N_32820);
nand U33368 (N_33368,N_32900,N_32700);
nand U33369 (N_33369,N_32994,N_32865);
and U33370 (N_33370,N_32696,N_32993);
and U33371 (N_33371,N_32895,N_32966);
or U33372 (N_33372,N_32671,N_32628);
nor U33373 (N_33373,N_32794,N_32825);
nand U33374 (N_33374,N_32997,N_32809);
or U33375 (N_33375,N_32800,N_32684);
or U33376 (N_33376,N_32654,N_32591);
nor U33377 (N_33377,N_32963,N_32783);
nor U33378 (N_33378,N_32605,N_32646);
nor U33379 (N_33379,N_32939,N_32661);
or U33380 (N_33380,N_32970,N_32935);
or U33381 (N_33381,N_32934,N_32979);
or U33382 (N_33382,N_32688,N_32916);
xor U33383 (N_33383,N_32514,N_32698);
or U33384 (N_33384,N_32995,N_32897);
or U33385 (N_33385,N_32518,N_32772);
nor U33386 (N_33386,N_32587,N_32829);
and U33387 (N_33387,N_32778,N_32887);
and U33388 (N_33388,N_32737,N_32548);
nand U33389 (N_33389,N_32696,N_32902);
nand U33390 (N_33390,N_32985,N_32623);
nand U33391 (N_33391,N_32923,N_32687);
nor U33392 (N_33392,N_32738,N_32994);
nand U33393 (N_33393,N_32751,N_32999);
nand U33394 (N_33394,N_32589,N_32805);
nand U33395 (N_33395,N_32550,N_32836);
nand U33396 (N_33396,N_32928,N_32678);
nand U33397 (N_33397,N_32624,N_32828);
nor U33398 (N_33398,N_32502,N_32509);
and U33399 (N_33399,N_32512,N_32989);
nand U33400 (N_33400,N_32625,N_32915);
nor U33401 (N_33401,N_32929,N_32530);
nand U33402 (N_33402,N_32744,N_32909);
xnor U33403 (N_33403,N_32878,N_32556);
nor U33404 (N_33404,N_32770,N_32577);
xnor U33405 (N_33405,N_32804,N_32983);
and U33406 (N_33406,N_32548,N_32876);
or U33407 (N_33407,N_32543,N_32749);
nand U33408 (N_33408,N_32781,N_32801);
nand U33409 (N_33409,N_32922,N_32765);
nor U33410 (N_33410,N_32835,N_32539);
xnor U33411 (N_33411,N_32634,N_32877);
or U33412 (N_33412,N_32515,N_32779);
nor U33413 (N_33413,N_32674,N_32766);
nand U33414 (N_33414,N_32675,N_32702);
nor U33415 (N_33415,N_32702,N_32691);
nand U33416 (N_33416,N_32718,N_32561);
and U33417 (N_33417,N_32874,N_32675);
or U33418 (N_33418,N_32923,N_32905);
nand U33419 (N_33419,N_32678,N_32746);
nor U33420 (N_33420,N_32943,N_32570);
or U33421 (N_33421,N_32995,N_32979);
nand U33422 (N_33422,N_32822,N_32859);
and U33423 (N_33423,N_32615,N_32623);
xor U33424 (N_33424,N_32835,N_32622);
or U33425 (N_33425,N_32882,N_32783);
xnor U33426 (N_33426,N_32831,N_32650);
or U33427 (N_33427,N_32518,N_32957);
and U33428 (N_33428,N_32683,N_32534);
xnor U33429 (N_33429,N_32746,N_32966);
or U33430 (N_33430,N_32992,N_32597);
xnor U33431 (N_33431,N_32655,N_32660);
xor U33432 (N_33432,N_32796,N_32965);
or U33433 (N_33433,N_32863,N_32681);
nand U33434 (N_33434,N_32749,N_32898);
xor U33435 (N_33435,N_32788,N_32709);
and U33436 (N_33436,N_32901,N_32787);
or U33437 (N_33437,N_32743,N_32848);
or U33438 (N_33438,N_32911,N_32873);
nor U33439 (N_33439,N_32833,N_32658);
nor U33440 (N_33440,N_32530,N_32660);
nand U33441 (N_33441,N_32594,N_32836);
nand U33442 (N_33442,N_32870,N_32864);
nand U33443 (N_33443,N_32509,N_32699);
nor U33444 (N_33444,N_32670,N_32569);
nor U33445 (N_33445,N_32861,N_32975);
nand U33446 (N_33446,N_32910,N_32513);
xor U33447 (N_33447,N_32950,N_32618);
xnor U33448 (N_33448,N_32746,N_32810);
or U33449 (N_33449,N_32612,N_32876);
nor U33450 (N_33450,N_32989,N_32933);
nor U33451 (N_33451,N_32976,N_32620);
xor U33452 (N_33452,N_32877,N_32856);
and U33453 (N_33453,N_32959,N_32856);
xor U33454 (N_33454,N_32576,N_32521);
and U33455 (N_33455,N_32514,N_32562);
and U33456 (N_33456,N_32821,N_32907);
nor U33457 (N_33457,N_32820,N_32905);
nor U33458 (N_33458,N_32796,N_32728);
or U33459 (N_33459,N_32926,N_32781);
nand U33460 (N_33460,N_32843,N_32637);
xnor U33461 (N_33461,N_32769,N_32758);
nor U33462 (N_33462,N_32658,N_32837);
and U33463 (N_33463,N_32855,N_32867);
xor U33464 (N_33464,N_32893,N_32769);
xnor U33465 (N_33465,N_32513,N_32856);
xor U33466 (N_33466,N_32967,N_32961);
nor U33467 (N_33467,N_32693,N_32535);
or U33468 (N_33468,N_32804,N_32980);
and U33469 (N_33469,N_32747,N_32634);
and U33470 (N_33470,N_32901,N_32956);
nand U33471 (N_33471,N_32795,N_32813);
nand U33472 (N_33472,N_32605,N_32594);
and U33473 (N_33473,N_32598,N_32537);
nor U33474 (N_33474,N_32672,N_32804);
nor U33475 (N_33475,N_32714,N_32842);
xnor U33476 (N_33476,N_32864,N_32568);
xor U33477 (N_33477,N_32837,N_32590);
nor U33478 (N_33478,N_32884,N_32542);
nand U33479 (N_33479,N_32990,N_32538);
nor U33480 (N_33480,N_32669,N_32973);
nor U33481 (N_33481,N_32520,N_32557);
and U33482 (N_33482,N_32775,N_32736);
nand U33483 (N_33483,N_32739,N_32708);
and U33484 (N_33484,N_32536,N_32657);
nand U33485 (N_33485,N_32980,N_32563);
nand U33486 (N_33486,N_32800,N_32751);
or U33487 (N_33487,N_32583,N_32566);
nor U33488 (N_33488,N_32965,N_32720);
nand U33489 (N_33489,N_32750,N_32955);
nor U33490 (N_33490,N_32729,N_32701);
and U33491 (N_33491,N_32654,N_32934);
xor U33492 (N_33492,N_32708,N_32869);
or U33493 (N_33493,N_32937,N_32604);
nand U33494 (N_33494,N_32616,N_32753);
or U33495 (N_33495,N_32783,N_32805);
or U33496 (N_33496,N_32959,N_32813);
and U33497 (N_33497,N_32538,N_32798);
xor U33498 (N_33498,N_32698,N_32738);
xor U33499 (N_33499,N_32995,N_32734);
and U33500 (N_33500,N_33147,N_33034);
xor U33501 (N_33501,N_33262,N_33291);
and U33502 (N_33502,N_33404,N_33430);
nand U33503 (N_33503,N_33072,N_33195);
nor U33504 (N_33504,N_33251,N_33422);
xnor U33505 (N_33505,N_33011,N_33379);
and U33506 (N_33506,N_33215,N_33161);
or U33507 (N_33507,N_33304,N_33051);
nor U33508 (N_33508,N_33055,N_33324);
xnor U33509 (N_33509,N_33470,N_33007);
and U33510 (N_33510,N_33057,N_33210);
xor U33511 (N_33511,N_33299,N_33157);
xor U33512 (N_33512,N_33335,N_33431);
nand U33513 (N_33513,N_33068,N_33280);
xor U33514 (N_33514,N_33120,N_33439);
and U33515 (N_33515,N_33252,N_33080);
and U33516 (N_33516,N_33248,N_33376);
nand U33517 (N_33517,N_33455,N_33006);
nand U33518 (N_33518,N_33010,N_33166);
and U33519 (N_33519,N_33468,N_33315);
nor U33520 (N_33520,N_33488,N_33014);
nand U33521 (N_33521,N_33040,N_33360);
or U33522 (N_33522,N_33241,N_33064);
nand U33523 (N_33523,N_33276,N_33222);
and U33524 (N_33524,N_33374,N_33037);
xnor U33525 (N_33525,N_33204,N_33485);
xnor U33526 (N_33526,N_33228,N_33473);
and U33527 (N_33527,N_33487,N_33388);
or U33528 (N_33528,N_33364,N_33044);
nand U33529 (N_33529,N_33085,N_33423);
nand U33530 (N_33530,N_33076,N_33476);
nand U33531 (N_33531,N_33395,N_33021);
nand U33532 (N_33532,N_33081,N_33174);
or U33533 (N_33533,N_33450,N_33296);
nor U33534 (N_33534,N_33109,N_33321);
nor U33535 (N_33535,N_33414,N_33428);
nand U33536 (N_33536,N_33329,N_33405);
nand U33537 (N_33537,N_33458,N_33005);
and U33538 (N_33538,N_33039,N_33119);
xor U33539 (N_33539,N_33460,N_33118);
or U33540 (N_33540,N_33145,N_33244);
xor U33541 (N_33541,N_33275,N_33362);
and U33542 (N_33542,N_33236,N_33350);
and U33543 (N_33543,N_33267,N_33142);
xnor U33544 (N_33544,N_33305,N_33392);
xor U33545 (N_33545,N_33060,N_33096);
nand U33546 (N_33546,N_33465,N_33383);
and U33547 (N_33547,N_33282,N_33486);
and U33548 (N_33548,N_33170,N_33406);
nor U33549 (N_33549,N_33151,N_33225);
and U33550 (N_33550,N_33095,N_33053);
xnor U33551 (N_33551,N_33012,N_33309);
and U33552 (N_33552,N_33424,N_33144);
nand U33553 (N_33553,N_33272,N_33330);
nand U33554 (N_33554,N_33004,N_33255);
nor U33555 (N_33555,N_33415,N_33246);
nand U33556 (N_33556,N_33483,N_33466);
nor U33557 (N_33557,N_33141,N_33198);
and U33558 (N_33558,N_33288,N_33314);
or U33559 (N_33559,N_33397,N_33219);
xnor U33560 (N_33560,N_33361,N_33365);
or U33561 (N_33561,N_33322,N_33290);
or U33562 (N_33562,N_33497,N_33347);
xnor U33563 (N_33563,N_33393,N_33363);
nand U33564 (N_33564,N_33054,N_33307);
xor U33565 (N_33565,N_33155,N_33443);
and U33566 (N_33566,N_33449,N_33352);
nand U33567 (N_33567,N_33094,N_33373);
and U33568 (N_33568,N_33162,N_33464);
nand U33569 (N_33569,N_33220,N_33201);
nand U33570 (N_33570,N_33143,N_33176);
xor U33571 (N_33571,N_33008,N_33092);
nor U33572 (N_33572,N_33384,N_33368);
nand U33573 (N_33573,N_33227,N_33213);
nor U33574 (N_33574,N_33442,N_33286);
and U33575 (N_33575,N_33190,N_33089);
and U33576 (N_33576,N_33242,N_33351);
and U33577 (N_33577,N_33075,N_33050);
nand U33578 (N_33578,N_33498,N_33130);
nand U33579 (N_33579,N_33214,N_33031);
or U33580 (N_33580,N_33371,N_33391);
xnor U33581 (N_33581,N_33325,N_33208);
xor U33582 (N_33582,N_33336,N_33292);
and U33583 (N_33583,N_33223,N_33418);
xnor U33584 (N_33584,N_33191,N_33293);
and U33585 (N_33585,N_33452,N_33038);
or U33586 (N_33586,N_33249,N_33110);
xor U33587 (N_33587,N_33029,N_33212);
and U33588 (N_33588,N_33394,N_33494);
xor U33589 (N_33589,N_33444,N_33359);
nand U33590 (N_33590,N_33186,N_33230);
xor U33591 (N_33591,N_33243,N_33387);
xor U33592 (N_33592,N_33357,N_33331);
and U33593 (N_33593,N_33066,N_33349);
nor U33594 (N_33594,N_33000,N_33104);
and U33595 (N_33595,N_33283,N_33375);
and U33596 (N_33596,N_33340,N_33160);
and U33597 (N_33597,N_33126,N_33149);
nor U33598 (N_33598,N_33049,N_33343);
nand U33599 (N_33599,N_33270,N_33348);
nand U33600 (N_33600,N_33226,N_33377);
and U33601 (N_33601,N_33328,N_33389);
or U33602 (N_33602,N_33199,N_33339);
or U33603 (N_33603,N_33015,N_33146);
nand U33604 (N_33604,N_33323,N_33217);
and U33605 (N_33605,N_33346,N_33457);
nand U33606 (N_33606,N_33074,N_33071);
nand U33607 (N_33607,N_33337,N_33193);
nor U33608 (N_33608,N_33203,N_33148);
or U33609 (N_33609,N_33052,N_33165);
nor U33610 (N_33610,N_33462,N_33491);
nor U33611 (N_33611,N_33107,N_33172);
nand U33612 (N_33612,N_33413,N_33002);
and U33613 (N_33613,N_33033,N_33035);
xor U33614 (N_33614,N_33344,N_33221);
nor U33615 (N_33615,N_33231,N_33420);
or U33616 (N_33616,N_33433,N_33396);
and U33617 (N_33617,N_33285,N_33023);
or U33618 (N_33618,N_33245,N_33234);
or U33619 (N_33619,N_33024,N_33438);
nor U33620 (N_33620,N_33202,N_33298);
nor U33621 (N_33621,N_33129,N_33065);
and U33622 (N_33622,N_33077,N_33097);
and U33623 (N_33623,N_33381,N_33209);
and U33624 (N_33624,N_33062,N_33279);
or U33625 (N_33625,N_33078,N_33232);
nand U33626 (N_33626,N_33237,N_33061);
nor U33627 (N_33627,N_33152,N_33326);
nand U33628 (N_33628,N_33451,N_33135);
or U33629 (N_33629,N_33009,N_33183);
nand U33630 (N_33630,N_33302,N_33284);
xnor U33631 (N_33631,N_33090,N_33271);
nor U33632 (N_33632,N_33372,N_33088);
xnor U33633 (N_33633,N_33278,N_33345);
xnor U33634 (N_33634,N_33171,N_33316);
and U33635 (N_33635,N_33312,N_33069);
xnor U33636 (N_33636,N_33434,N_33429);
and U33637 (N_33637,N_33131,N_33042);
nor U33638 (N_33638,N_33022,N_33206);
or U33639 (N_33639,N_33250,N_33093);
and U33640 (N_33640,N_33277,N_33269);
or U33641 (N_33641,N_33303,N_33103);
nor U33642 (N_33642,N_33492,N_33367);
nand U33643 (N_33643,N_33106,N_33259);
xor U33644 (N_33644,N_33479,N_33001);
xnor U33645 (N_33645,N_33308,N_33059);
and U33646 (N_33646,N_33099,N_33495);
or U33647 (N_33647,N_33318,N_33268);
or U33648 (N_33648,N_33447,N_33197);
nand U33649 (N_33649,N_33385,N_33378);
xnor U33650 (N_33650,N_33108,N_33184);
xor U33651 (N_33651,N_33264,N_33490);
nor U33652 (N_33652,N_33273,N_33224);
nand U33653 (N_33653,N_33086,N_33091);
nor U33654 (N_33654,N_33274,N_33432);
or U33655 (N_33655,N_33116,N_33056);
nor U33656 (N_33656,N_33113,N_33185);
and U33657 (N_33657,N_33254,N_33134);
nor U33658 (N_33658,N_33122,N_33489);
nand U33659 (N_33659,N_33453,N_33102);
nor U33660 (N_33660,N_33154,N_33358);
nor U33661 (N_33661,N_33137,N_33169);
or U33662 (N_33662,N_33063,N_33471);
or U33663 (N_33663,N_33140,N_33030);
and U33664 (N_33664,N_33111,N_33260);
nand U33665 (N_33665,N_33016,N_33334);
nand U33666 (N_33666,N_33207,N_33101);
and U33667 (N_33667,N_33425,N_33480);
nand U33668 (N_33668,N_33027,N_33180);
nand U33669 (N_33669,N_33426,N_33463);
and U33670 (N_33670,N_33353,N_33018);
nor U33671 (N_33671,N_33150,N_33182);
nor U33672 (N_33672,N_33370,N_33239);
nor U33673 (N_33673,N_33187,N_33300);
and U33674 (N_33674,N_33341,N_33205);
or U33675 (N_33675,N_33257,N_33445);
xnor U33676 (N_33676,N_33067,N_33416);
and U33677 (N_33677,N_33265,N_33019);
nand U33678 (N_33678,N_33295,N_33319);
or U33679 (N_33679,N_33164,N_33320);
or U33680 (N_33680,N_33200,N_33411);
xor U33681 (N_33681,N_33105,N_33047);
and U33682 (N_33682,N_33297,N_33013);
nor U33683 (N_33683,N_33459,N_33098);
xnor U33684 (N_33684,N_33117,N_33181);
nand U33685 (N_33685,N_33410,N_33263);
xnor U33686 (N_33686,N_33238,N_33070);
nor U33687 (N_33687,N_33448,N_33366);
or U33688 (N_33688,N_33356,N_33311);
nand U33689 (N_33689,N_33294,N_33258);
or U33690 (N_33690,N_33218,N_33369);
and U33691 (N_33691,N_33354,N_33382);
nor U33692 (N_33692,N_33178,N_33087);
or U33693 (N_33693,N_33261,N_33496);
xnor U33694 (N_33694,N_33437,N_33402);
and U33695 (N_33695,N_33233,N_33475);
nand U33696 (N_33696,N_33482,N_33127);
nor U33697 (N_33697,N_33082,N_33456);
xor U33698 (N_33698,N_33017,N_33036);
nor U33699 (N_33699,N_33412,N_33125);
nor U33700 (N_33700,N_33048,N_33454);
or U33701 (N_33701,N_33333,N_33159);
and U33702 (N_33702,N_33133,N_33441);
or U33703 (N_33703,N_33380,N_33121);
and U33704 (N_33704,N_33123,N_33058);
or U33705 (N_33705,N_33399,N_33240);
nand U33706 (N_33706,N_33287,N_33156);
nor U33707 (N_33707,N_33045,N_33073);
and U33708 (N_33708,N_33417,N_33083);
nand U33709 (N_33709,N_33313,N_33499);
nor U33710 (N_33710,N_33427,N_33211);
nor U33711 (N_33711,N_33446,N_33177);
and U33712 (N_33712,N_33216,N_33306);
xor U33713 (N_33713,N_33390,N_33253);
nor U33714 (N_33714,N_33079,N_33332);
and U33715 (N_33715,N_33175,N_33467);
or U33716 (N_33716,N_33189,N_33435);
and U33717 (N_33717,N_33043,N_33235);
xnor U33718 (N_33718,N_33179,N_33115);
xor U33719 (N_33719,N_33409,N_33493);
nor U33720 (N_33720,N_33484,N_33469);
or U33721 (N_33721,N_33400,N_33408);
nor U33722 (N_33722,N_33342,N_33167);
nand U33723 (N_33723,N_33138,N_33041);
xnor U33724 (N_33724,N_33124,N_33266);
nor U33725 (N_33725,N_33327,N_33003);
nor U33726 (N_33726,N_33153,N_33407);
and U33727 (N_33727,N_33128,N_33158);
and U33728 (N_33728,N_33338,N_33472);
xor U33729 (N_33729,N_33192,N_33477);
nor U33730 (N_33730,N_33168,N_33247);
and U33731 (N_33731,N_33421,N_33436);
or U33732 (N_33732,N_33132,N_33440);
nor U33733 (N_33733,N_33481,N_33310);
xnor U33734 (N_33734,N_33317,N_33478);
nor U33735 (N_33735,N_33301,N_33401);
nor U33736 (N_33736,N_33026,N_33419);
nand U33737 (N_33737,N_33163,N_33032);
and U33738 (N_33738,N_33046,N_33139);
nand U33739 (N_33739,N_33173,N_33474);
xnor U33740 (N_33740,N_33194,N_33136);
nand U33741 (N_33741,N_33289,N_33028);
xor U33742 (N_33742,N_33084,N_33229);
nor U33743 (N_33743,N_33025,N_33281);
and U33744 (N_33744,N_33100,N_33355);
and U33745 (N_33745,N_33020,N_33114);
or U33746 (N_33746,N_33188,N_33196);
nand U33747 (N_33747,N_33398,N_33461);
xor U33748 (N_33748,N_33403,N_33112);
xor U33749 (N_33749,N_33386,N_33256);
or U33750 (N_33750,N_33123,N_33240);
or U33751 (N_33751,N_33256,N_33372);
nand U33752 (N_33752,N_33135,N_33294);
nand U33753 (N_33753,N_33203,N_33184);
nor U33754 (N_33754,N_33175,N_33212);
and U33755 (N_33755,N_33194,N_33035);
and U33756 (N_33756,N_33380,N_33137);
nor U33757 (N_33757,N_33160,N_33199);
nor U33758 (N_33758,N_33468,N_33465);
nor U33759 (N_33759,N_33081,N_33272);
nor U33760 (N_33760,N_33336,N_33256);
or U33761 (N_33761,N_33290,N_33052);
and U33762 (N_33762,N_33009,N_33447);
nor U33763 (N_33763,N_33069,N_33465);
or U33764 (N_33764,N_33270,N_33402);
or U33765 (N_33765,N_33471,N_33145);
nand U33766 (N_33766,N_33159,N_33400);
nand U33767 (N_33767,N_33071,N_33141);
or U33768 (N_33768,N_33442,N_33208);
and U33769 (N_33769,N_33419,N_33094);
nand U33770 (N_33770,N_33467,N_33249);
xnor U33771 (N_33771,N_33169,N_33045);
and U33772 (N_33772,N_33462,N_33147);
or U33773 (N_33773,N_33137,N_33149);
xor U33774 (N_33774,N_33285,N_33276);
xor U33775 (N_33775,N_33088,N_33456);
nor U33776 (N_33776,N_33151,N_33401);
nor U33777 (N_33777,N_33495,N_33128);
and U33778 (N_33778,N_33443,N_33494);
nand U33779 (N_33779,N_33076,N_33153);
nand U33780 (N_33780,N_33217,N_33358);
xnor U33781 (N_33781,N_33398,N_33474);
xnor U33782 (N_33782,N_33170,N_33355);
nor U33783 (N_33783,N_33340,N_33386);
and U33784 (N_33784,N_33173,N_33238);
or U33785 (N_33785,N_33226,N_33101);
nor U33786 (N_33786,N_33321,N_33177);
xnor U33787 (N_33787,N_33495,N_33039);
or U33788 (N_33788,N_33242,N_33062);
nor U33789 (N_33789,N_33018,N_33101);
and U33790 (N_33790,N_33156,N_33204);
nor U33791 (N_33791,N_33482,N_33029);
and U33792 (N_33792,N_33475,N_33261);
and U33793 (N_33793,N_33392,N_33143);
xor U33794 (N_33794,N_33342,N_33131);
and U33795 (N_33795,N_33175,N_33466);
or U33796 (N_33796,N_33013,N_33223);
nand U33797 (N_33797,N_33241,N_33026);
nor U33798 (N_33798,N_33118,N_33364);
nand U33799 (N_33799,N_33448,N_33439);
nor U33800 (N_33800,N_33042,N_33171);
and U33801 (N_33801,N_33194,N_33291);
xor U33802 (N_33802,N_33158,N_33079);
nor U33803 (N_33803,N_33433,N_33236);
nor U33804 (N_33804,N_33122,N_33006);
xor U33805 (N_33805,N_33337,N_33271);
or U33806 (N_33806,N_33271,N_33209);
and U33807 (N_33807,N_33340,N_33457);
or U33808 (N_33808,N_33196,N_33159);
or U33809 (N_33809,N_33392,N_33141);
nor U33810 (N_33810,N_33358,N_33388);
or U33811 (N_33811,N_33372,N_33462);
and U33812 (N_33812,N_33433,N_33341);
nand U33813 (N_33813,N_33047,N_33205);
nand U33814 (N_33814,N_33268,N_33497);
xor U33815 (N_33815,N_33083,N_33149);
and U33816 (N_33816,N_33468,N_33076);
or U33817 (N_33817,N_33091,N_33206);
or U33818 (N_33818,N_33310,N_33382);
nor U33819 (N_33819,N_33465,N_33191);
and U33820 (N_33820,N_33412,N_33017);
and U33821 (N_33821,N_33091,N_33413);
and U33822 (N_33822,N_33252,N_33365);
or U33823 (N_33823,N_33157,N_33072);
nor U33824 (N_33824,N_33151,N_33172);
xor U33825 (N_33825,N_33078,N_33130);
or U33826 (N_33826,N_33213,N_33490);
and U33827 (N_33827,N_33034,N_33014);
and U33828 (N_33828,N_33232,N_33494);
xnor U33829 (N_33829,N_33044,N_33480);
or U33830 (N_33830,N_33497,N_33420);
nor U33831 (N_33831,N_33486,N_33225);
or U33832 (N_33832,N_33029,N_33081);
nand U33833 (N_33833,N_33035,N_33270);
and U33834 (N_33834,N_33126,N_33253);
and U33835 (N_33835,N_33264,N_33188);
nand U33836 (N_33836,N_33094,N_33049);
and U33837 (N_33837,N_33422,N_33163);
and U33838 (N_33838,N_33426,N_33311);
and U33839 (N_33839,N_33012,N_33444);
nand U33840 (N_33840,N_33329,N_33133);
xor U33841 (N_33841,N_33066,N_33293);
nor U33842 (N_33842,N_33064,N_33363);
nand U33843 (N_33843,N_33357,N_33375);
or U33844 (N_33844,N_33070,N_33208);
or U33845 (N_33845,N_33084,N_33048);
and U33846 (N_33846,N_33155,N_33490);
and U33847 (N_33847,N_33026,N_33495);
or U33848 (N_33848,N_33026,N_33273);
or U33849 (N_33849,N_33147,N_33375);
nand U33850 (N_33850,N_33019,N_33316);
nand U33851 (N_33851,N_33408,N_33280);
and U33852 (N_33852,N_33323,N_33025);
nand U33853 (N_33853,N_33348,N_33244);
or U33854 (N_33854,N_33235,N_33275);
and U33855 (N_33855,N_33323,N_33168);
or U33856 (N_33856,N_33263,N_33380);
nor U33857 (N_33857,N_33193,N_33208);
nand U33858 (N_33858,N_33093,N_33354);
xnor U33859 (N_33859,N_33099,N_33320);
xnor U33860 (N_33860,N_33412,N_33417);
nand U33861 (N_33861,N_33196,N_33043);
or U33862 (N_33862,N_33357,N_33430);
nand U33863 (N_33863,N_33336,N_33305);
xnor U33864 (N_33864,N_33433,N_33077);
xnor U33865 (N_33865,N_33278,N_33071);
or U33866 (N_33866,N_33394,N_33322);
xnor U33867 (N_33867,N_33138,N_33043);
nor U33868 (N_33868,N_33225,N_33289);
xnor U33869 (N_33869,N_33442,N_33488);
nor U33870 (N_33870,N_33443,N_33311);
nand U33871 (N_33871,N_33069,N_33414);
and U33872 (N_33872,N_33099,N_33131);
and U33873 (N_33873,N_33229,N_33094);
xnor U33874 (N_33874,N_33195,N_33158);
nor U33875 (N_33875,N_33319,N_33359);
xnor U33876 (N_33876,N_33317,N_33418);
nand U33877 (N_33877,N_33212,N_33196);
and U33878 (N_33878,N_33178,N_33464);
and U33879 (N_33879,N_33270,N_33440);
nand U33880 (N_33880,N_33381,N_33020);
and U33881 (N_33881,N_33331,N_33068);
nor U33882 (N_33882,N_33466,N_33359);
nand U33883 (N_33883,N_33490,N_33012);
nor U33884 (N_33884,N_33497,N_33480);
nor U33885 (N_33885,N_33491,N_33141);
xnor U33886 (N_33886,N_33273,N_33409);
xor U33887 (N_33887,N_33008,N_33223);
nor U33888 (N_33888,N_33378,N_33431);
xor U33889 (N_33889,N_33493,N_33117);
nor U33890 (N_33890,N_33006,N_33129);
nor U33891 (N_33891,N_33291,N_33075);
and U33892 (N_33892,N_33385,N_33483);
xor U33893 (N_33893,N_33426,N_33133);
xnor U33894 (N_33894,N_33084,N_33460);
nand U33895 (N_33895,N_33058,N_33280);
or U33896 (N_33896,N_33272,N_33176);
and U33897 (N_33897,N_33337,N_33071);
nand U33898 (N_33898,N_33030,N_33214);
or U33899 (N_33899,N_33350,N_33119);
or U33900 (N_33900,N_33129,N_33395);
or U33901 (N_33901,N_33166,N_33244);
or U33902 (N_33902,N_33189,N_33041);
xor U33903 (N_33903,N_33444,N_33034);
nand U33904 (N_33904,N_33347,N_33202);
nand U33905 (N_33905,N_33159,N_33348);
or U33906 (N_33906,N_33150,N_33360);
xor U33907 (N_33907,N_33432,N_33219);
xor U33908 (N_33908,N_33490,N_33485);
nor U33909 (N_33909,N_33389,N_33478);
xnor U33910 (N_33910,N_33435,N_33402);
nand U33911 (N_33911,N_33147,N_33156);
and U33912 (N_33912,N_33470,N_33289);
nand U33913 (N_33913,N_33272,N_33473);
or U33914 (N_33914,N_33158,N_33278);
xnor U33915 (N_33915,N_33339,N_33350);
xnor U33916 (N_33916,N_33180,N_33341);
or U33917 (N_33917,N_33128,N_33460);
or U33918 (N_33918,N_33220,N_33045);
or U33919 (N_33919,N_33196,N_33032);
xor U33920 (N_33920,N_33210,N_33195);
xnor U33921 (N_33921,N_33354,N_33185);
xor U33922 (N_33922,N_33433,N_33052);
or U33923 (N_33923,N_33028,N_33368);
xnor U33924 (N_33924,N_33153,N_33088);
or U33925 (N_33925,N_33012,N_33259);
xor U33926 (N_33926,N_33221,N_33309);
nor U33927 (N_33927,N_33169,N_33445);
nand U33928 (N_33928,N_33206,N_33266);
nand U33929 (N_33929,N_33173,N_33384);
or U33930 (N_33930,N_33238,N_33075);
nand U33931 (N_33931,N_33058,N_33304);
xor U33932 (N_33932,N_33286,N_33222);
xnor U33933 (N_33933,N_33111,N_33219);
nand U33934 (N_33934,N_33375,N_33039);
or U33935 (N_33935,N_33071,N_33243);
nand U33936 (N_33936,N_33312,N_33059);
nand U33937 (N_33937,N_33416,N_33161);
or U33938 (N_33938,N_33074,N_33029);
nor U33939 (N_33939,N_33432,N_33456);
and U33940 (N_33940,N_33151,N_33179);
nand U33941 (N_33941,N_33113,N_33355);
nor U33942 (N_33942,N_33327,N_33361);
xnor U33943 (N_33943,N_33485,N_33154);
nand U33944 (N_33944,N_33429,N_33054);
nand U33945 (N_33945,N_33382,N_33020);
xnor U33946 (N_33946,N_33498,N_33137);
xor U33947 (N_33947,N_33206,N_33306);
and U33948 (N_33948,N_33144,N_33433);
xnor U33949 (N_33949,N_33354,N_33303);
nor U33950 (N_33950,N_33237,N_33267);
nor U33951 (N_33951,N_33181,N_33084);
nor U33952 (N_33952,N_33070,N_33037);
nand U33953 (N_33953,N_33440,N_33459);
nand U33954 (N_33954,N_33005,N_33483);
or U33955 (N_33955,N_33166,N_33288);
nor U33956 (N_33956,N_33370,N_33140);
nor U33957 (N_33957,N_33421,N_33289);
nand U33958 (N_33958,N_33334,N_33215);
xor U33959 (N_33959,N_33096,N_33311);
xor U33960 (N_33960,N_33281,N_33048);
and U33961 (N_33961,N_33344,N_33043);
and U33962 (N_33962,N_33383,N_33174);
nand U33963 (N_33963,N_33402,N_33144);
nand U33964 (N_33964,N_33105,N_33489);
xor U33965 (N_33965,N_33098,N_33084);
xnor U33966 (N_33966,N_33265,N_33206);
nor U33967 (N_33967,N_33443,N_33498);
nand U33968 (N_33968,N_33194,N_33052);
nor U33969 (N_33969,N_33276,N_33025);
xnor U33970 (N_33970,N_33399,N_33494);
and U33971 (N_33971,N_33326,N_33359);
nand U33972 (N_33972,N_33040,N_33271);
and U33973 (N_33973,N_33271,N_33133);
nor U33974 (N_33974,N_33297,N_33488);
nand U33975 (N_33975,N_33114,N_33330);
xor U33976 (N_33976,N_33074,N_33037);
or U33977 (N_33977,N_33183,N_33117);
or U33978 (N_33978,N_33445,N_33004);
and U33979 (N_33979,N_33455,N_33155);
nand U33980 (N_33980,N_33401,N_33374);
xor U33981 (N_33981,N_33209,N_33064);
nor U33982 (N_33982,N_33050,N_33107);
xnor U33983 (N_33983,N_33324,N_33085);
nor U33984 (N_33984,N_33313,N_33336);
and U33985 (N_33985,N_33287,N_33268);
or U33986 (N_33986,N_33253,N_33381);
or U33987 (N_33987,N_33409,N_33030);
and U33988 (N_33988,N_33477,N_33424);
nand U33989 (N_33989,N_33214,N_33235);
nand U33990 (N_33990,N_33217,N_33288);
xor U33991 (N_33991,N_33163,N_33213);
and U33992 (N_33992,N_33304,N_33424);
nand U33993 (N_33993,N_33427,N_33379);
xor U33994 (N_33994,N_33361,N_33180);
or U33995 (N_33995,N_33369,N_33305);
nor U33996 (N_33996,N_33405,N_33491);
nand U33997 (N_33997,N_33383,N_33246);
nand U33998 (N_33998,N_33252,N_33444);
nand U33999 (N_33999,N_33178,N_33341);
xor U34000 (N_34000,N_33984,N_33521);
nor U34001 (N_34001,N_33856,N_33741);
nor U34002 (N_34002,N_33748,N_33925);
and U34003 (N_34003,N_33625,N_33956);
and U34004 (N_34004,N_33551,N_33908);
and U34005 (N_34005,N_33934,N_33791);
or U34006 (N_34006,N_33753,N_33800);
nand U34007 (N_34007,N_33536,N_33681);
xor U34008 (N_34008,N_33860,N_33605);
and U34009 (N_34009,N_33733,N_33718);
nand U34010 (N_34010,N_33990,N_33924);
xor U34011 (N_34011,N_33527,N_33634);
xnor U34012 (N_34012,N_33611,N_33994);
and U34013 (N_34013,N_33644,N_33998);
nand U34014 (N_34014,N_33651,N_33861);
xor U34015 (N_34015,N_33730,N_33722);
xnor U34016 (N_34016,N_33554,N_33729);
or U34017 (N_34017,N_33503,N_33633);
and U34018 (N_34018,N_33785,N_33824);
nand U34019 (N_34019,N_33576,N_33705);
xor U34020 (N_34020,N_33636,N_33547);
or U34021 (N_34021,N_33937,N_33737);
and U34022 (N_34022,N_33804,N_33706);
nor U34023 (N_34023,N_33889,N_33792);
or U34024 (N_34024,N_33794,N_33954);
xnor U34025 (N_34025,N_33936,N_33778);
xor U34026 (N_34026,N_33963,N_33784);
nor U34027 (N_34027,N_33827,N_33899);
nor U34028 (N_34028,N_33818,N_33606);
or U34029 (N_34029,N_33654,N_33969);
or U34030 (N_34030,N_33738,N_33915);
and U34031 (N_34031,N_33745,N_33630);
and U34032 (N_34032,N_33973,N_33906);
nand U34033 (N_34033,N_33702,N_33875);
nand U34034 (N_34034,N_33770,N_33689);
nor U34035 (N_34035,N_33996,N_33997);
nor U34036 (N_34036,N_33691,N_33767);
nand U34037 (N_34037,N_33945,N_33845);
xor U34038 (N_34038,N_33668,N_33789);
and U34039 (N_34039,N_33930,N_33768);
and U34040 (N_34040,N_33588,N_33764);
nand U34041 (N_34041,N_33658,N_33687);
nand U34042 (N_34042,N_33877,N_33568);
nand U34043 (N_34043,N_33574,N_33782);
or U34044 (N_34044,N_33762,N_33986);
or U34045 (N_34045,N_33869,N_33695);
or U34046 (N_34046,N_33892,N_33763);
xor U34047 (N_34047,N_33999,N_33585);
nor U34048 (N_34048,N_33571,N_33587);
or U34049 (N_34049,N_33978,N_33514);
or U34050 (N_34050,N_33834,N_33659);
xnor U34051 (N_34051,N_33679,N_33894);
nor U34052 (N_34052,N_33520,N_33720);
nand U34053 (N_34053,N_33885,N_33501);
nor U34054 (N_34054,N_33828,N_33858);
nand U34055 (N_34055,N_33874,N_33813);
or U34056 (N_34056,N_33913,N_33573);
and U34057 (N_34057,N_33979,N_33558);
nand U34058 (N_34058,N_33815,N_33697);
and U34059 (N_34059,N_33559,N_33935);
xnor U34060 (N_34060,N_33806,N_33816);
nand U34061 (N_34061,N_33970,N_33604);
nor U34062 (N_34062,N_33895,N_33656);
nand U34063 (N_34063,N_33927,N_33515);
and U34064 (N_34064,N_33591,N_33876);
nor U34065 (N_34065,N_33523,N_33678);
nand U34066 (N_34066,N_33534,N_33760);
xnor U34067 (N_34067,N_33629,N_33550);
nor U34068 (N_34068,N_33728,N_33731);
and U34069 (N_34069,N_33835,N_33953);
nand U34070 (N_34070,N_33504,N_33597);
nor U34071 (N_34071,N_33888,N_33739);
and U34072 (N_34072,N_33833,N_33972);
or U34073 (N_34073,N_33736,N_33788);
xnor U34074 (N_34074,N_33590,N_33796);
xor U34075 (N_34075,N_33980,N_33864);
and U34076 (N_34076,N_33616,N_33849);
and U34077 (N_34077,N_33982,N_33532);
or U34078 (N_34078,N_33964,N_33744);
xor U34079 (N_34079,N_33929,N_33840);
nor U34080 (N_34080,N_33583,N_33655);
xnor U34081 (N_34081,N_33623,N_33557);
or U34082 (N_34082,N_33732,N_33727);
xnor U34083 (N_34083,N_33923,N_33820);
xnor U34084 (N_34084,N_33992,N_33955);
and U34085 (N_34085,N_33988,N_33862);
nand U34086 (N_34086,N_33940,N_33593);
nor U34087 (N_34087,N_33901,N_33848);
nand U34088 (N_34088,N_33628,N_33653);
and U34089 (N_34089,N_33569,N_33620);
and U34090 (N_34090,N_33664,N_33939);
xor U34091 (N_34091,N_33805,N_33761);
nand U34092 (N_34092,N_33649,N_33635);
xor U34093 (N_34093,N_33841,N_33533);
or U34094 (N_34094,N_33867,N_33772);
nand U34095 (N_34095,N_33933,N_33638);
nor U34096 (N_34096,N_33803,N_33755);
and U34097 (N_34097,N_33952,N_33517);
or U34098 (N_34098,N_33563,N_33948);
nor U34099 (N_34099,N_33843,N_33713);
xor U34100 (N_34100,N_33809,N_33650);
nand U34101 (N_34101,N_33893,N_33540);
nor U34102 (N_34102,N_33844,N_33884);
xor U34103 (N_34103,N_33696,N_33910);
and U34104 (N_34104,N_33709,N_33811);
xnor U34105 (N_34105,N_33586,N_33707);
or U34106 (N_34106,N_33543,N_33661);
or U34107 (N_34107,N_33757,N_33526);
nand U34108 (N_34108,N_33688,N_33890);
nor U34109 (N_34109,N_33712,N_33759);
xnor U34110 (N_34110,N_33667,N_33613);
and U34111 (N_34111,N_33799,N_33662);
xnor U34112 (N_34112,N_33637,N_33962);
nor U34113 (N_34113,N_33795,N_33579);
nor U34114 (N_34114,N_33859,N_33842);
nand U34115 (N_34115,N_33565,N_33584);
xor U34116 (N_34116,N_33786,N_33823);
nor U34117 (N_34117,N_33631,N_33747);
xnor U34118 (N_34118,N_33643,N_33868);
or U34119 (N_34119,N_33989,N_33754);
nor U34120 (N_34120,N_33694,N_33938);
and U34121 (N_34121,N_33900,N_33983);
or U34122 (N_34122,N_33663,N_33993);
nor U34123 (N_34123,N_33821,N_33580);
nand U34124 (N_34124,N_33987,N_33529);
xnor U34125 (N_34125,N_33682,N_33595);
and U34126 (N_34126,N_33615,N_33909);
or U34127 (N_34127,N_33646,N_33780);
or U34128 (N_34128,N_33950,N_33609);
or U34129 (N_34129,N_33891,N_33775);
nor U34130 (N_34130,N_33798,N_33545);
nand U34131 (N_34131,N_33853,N_33510);
or U34132 (N_34132,N_33898,N_33581);
and U34133 (N_34133,N_33971,N_33807);
nor U34134 (N_34134,N_33850,N_33756);
and U34135 (N_34135,N_33854,N_33692);
xor U34136 (N_34136,N_33817,N_33947);
nor U34137 (N_34137,N_33704,N_33564);
nand U34138 (N_34138,N_33648,N_33690);
and U34139 (N_34139,N_33642,N_33814);
nor U34140 (N_34140,N_33836,N_33621);
nand U34141 (N_34141,N_33873,N_33944);
and U34142 (N_34142,N_33539,N_33887);
xnor U34143 (N_34143,N_33919,N_33716);
and U34144 (N_34144,N_33812,N_33645);
nor U34145 (N_34145,N_33671,N_33670);
xor U34146 (N_34146,N_33548,N_33535);
xnor U34147 (N_34147,N_33904,N_33566);
xnor U34148 (N_34148,N_33752,N_33619);
nor U34149 (N_34149,N_33603,N_33881);
nand U34150 (N_34150,N_33639,N_33880);
or U34151 (N_34151,N_33693,N_33610);
nand U34152 (N_34152,N_33830,N_33958);
and U34153 (N_34153,N_33657,N_33787);
xnor U34154 (N_34154,N_33560,N_33905);
xnor U34155 (N_34155,N_33832,N_33749);
nand U34156 (N_34156,N_33700,N_33897);
or U34157 (N_34157,N_33592,N_33669);
nand U34158 (N_34158,N_33556,N_33546);
or U34159 (N_34159,N_33522,N_33777);
and U34160 (N_34160,N_33949,N_33968);
nor U34161 (N_34161,N_33624,N_33672);
xnor U34162 (N_34162,N_33942,N_33544);
nor U34163 (N_34163,N_33740,N_33577);
or U34164 (N_34164,N_33685,N_33921);
and U34165 (N_34165,N_33734,N_33932);
or U34166 (N_34166,N_33721,N_33618);
or U34167 (N_34167,N_33525,N_33641);
and U34168 (N_34168,N_33911,N_33931);
and U34169 (N_34169,N_33528,N_33502);
and U34170 (N_34170,N_33974,N_33567);
xor U34171 (N_34171,N_33626,N_33505);
nand U34172 (N_34172,N_33516,N_33801);
and U34173 (N_34173,N_33724,N_33951);
and U34174 (N_34174,N_33710,N_33810);
or U34175 (N_34175,N_33882,N_33977);
nand U34176 (N_34176,N_33975,N_33866);
nor U34177 (N_34177,N_33647,N_33686);
nor U34178 (N_34178,N_33779,N_33781);
or U34179 (N_34179,N_33918,N_33596);
nand U34180 (N_34180,N_33676,N_33995);
nor U34181 (N_34181,N_33917,N_33500);
nor U34182 (N_34182,N_33549,N_33912);
xor U34183 (N_34183,N_33714,N_33617);
and U34184 (N_34184,N_33746,N_33839);
or U34185 (N_34185,N_33509,N_33965);
nor U34186 (N_34186,N_33766,N_33673);
xnor U34187 (N_34187,N_33666,N_33774);
nand U34188 (N_34188,N_33742,N_33808);
nor U34189 (N_34189,N_33561,N_33879);
or U34190 (N_34190,N_33758,N_33871);
or U34191 (N_34191,N_33765,N_33961);
or U34192 (N_34192,N_33793,N_33524);
or U34193 (N_34193,N_33507,N_33773);
nand U34194 (N_34194,N_33903,N_33914);
nand U34195 (N_34195,N_33957,N_33959);
or U34196 (N_34196,N_33941,N_33857);
and U34197 (N_34197,N_33920,N_33852);
and U34198 (N_34198,N_33872,N_33847);
nand U34199 (N_34199,N_33870,N_33640);
nor U34200 (N_34200,N_33723,N_33826);
or U34201 (N_34201,N_33599,N_33511);
or U34202 (N_34202,N_33614,N_33717);
nand U34203 (N_34203,N_33572,N_33594);
nor U34204 (N_34204,N_33976,N_33703);
and U34205 (N_34205,N_33769,N_33537);
nand U34206 (N_34206,N_33519,N_33675);
xor U34207 (N_34207,N_33582,N_33674);
nor U34208 (N_34208,N_33896,N_33902);
xor U34209 (N_34209,N_33837,N_33726);
xor U34210 (N_34210,N_33607,N_33797);
or U34211 (N_34211,N_33776,N_33846);
xnor U34212 (N_34212,N_33783,N_33531);
or U34213 (N_34213,N_33570,N_33589);
xnor U34214 (N_34214,N_33602,N_33665);
and U34215 (N_34215,N_33967,N_33966);
nand U34216 (N_34216,N_33513,N_33708);
or U34217 (N_34217,N_33922,N_33552);
nand U34218 (N_34218,N_33698,N_33829);
nor U34219 (N_34219,N_33508,N_33743);
or U34220 (N_34220,N_33802,N_33725);
or U34221 (N_34221,N_33916,N_33600);
nand U34222 (N_34222,N_33865,N_33627);
nand U34223 (N_34223,N_33553,N_33715);
nor U34224 (N_34224,N_33960,N_33991);
nor U34225 (N_34225,N_33863,N_33822);
nand U34226 (N_34226,N_33622,N_33886);
nor U34227 (N_34227,N_33684,N_33750);
nand U34228 (N_34228,N_33578,N_33612);
or U34229 (N_34229,N_33541,N_33719);
xnor U34230 (N_34230,N_33680,N_33771);
nand U34231 (N_34231,N_33981,N_33711);
or U34232 (N_34232,N_33699,N_33538);
nor U34233 (N_34233,N_33819,N_33562);
and U34234 (N_34234,N_33883,N_33751);
and U34235 (N_34235,N_33855,N_33518);
xnor U34236 (N_34236,N_33825,N_33506);
xnor U34237 (N_34237,N_33735,N_33926);
nand U34238 (N_34238,N_33652,N_33831);
xnor U34239 (N_34239,N_33701,N_33530);
nand U34240 (N_34240,N_33542,N_33660);
or U34241 (N_34241,N_33946,N_33555);
nand U34242 (N_34242,N_33851,N_33632);
or U34243 (N_34243,N_33677,N_33985);
nand U34244 (N_34244,N_33683,N_33598);
and U34245 (N_34245,N_33601,N_33512);
nor U34246 (N_34246,N_33878,N_33575);
xor U34247 (N_34247,N_33907,N_33838);
or U34248 (N_34248,N_33790,N_33608);
and U34249 (N_34249,N_33928,N_33943);
nor U34250 (N_34250,N_33829,N_33638);
xnor U34251 (N_34251,N_33864,N_33738);
or U34252 (N_34252,N_33555,N_33508);
or U34253 (N_34253,N_33859,N_33723);
nor U34254 (N_34254,N_33920,N_33587);
nand U34255 (N_34255,N_33706,N_33501);
nor U34256 (N_34256,N_33560,N_33824);
xnor U34257 (N_34257,N_33987,N_33955);
and U34258 (N_34258,N_33658,N_33791);
and U34259 (N_34259,N_33610,N_33919);
or U34260 (N_34260,N_33950,N_33928);
and U34261 (N_34261,N_33781,N_33655);
or U34262 (N_34262,N_33750,N_33501);
and U34263 (N_34263,N_33976,N_33593);
and U34264 (N_34264,N_33659,N_33726);
nor U34265 (N_34265,N_33555,N_33989);
nand U34266 (N_34266,N_33549,N_33648);
xor U34267 (N_34267,N_33711,N_33580);
or U34268 (N_34268,N_33995,N_33740);
xnor U34269 (N_34269,N_33997,N_33672);
and U34270 (N_34270,N_33672,N_33861);
or U34271 (N_34271,N_33801,N_33959);
xnor U34272 (N_34272,N_33932,N_33760);
nor U34273 (N_34273,N_33736,N_33567);
and U34274 (N_34274,N_33822,N_33799);
and U34275 (N_34275,N_33619,N_33775);
nand U34276 (N_34276,N_33665,N_33693);
and U34277 (N_34277,N_33914,N_33726);
nor U34278 (N_34278,N_33583,N_33854);
nand U34279 (N_34279,N_33876,N_33993);
nand U34280 (N_34280,N_33979,N_33942);
nand U34281 (N_34281,N_33510,N_33917);
nand U34282 (N_34282,N_33518,N_33719);
nand U34283 (N_34283,N_33849,N_33716);
and U34284 (N_34284,N_33692,N_33930);
and U34285 (N_34285,N_33719,N_33988);
or U34286 (N_34286,N_33984,N_33594);
xor U34287 (N_34287,N_33503,N_33864);
nor U34288 (N_34288,N_33520,N_33895);
nand U34289 (N_34289,N_33646,N_33623);
nand U34290 (N_34290,N_33533,N_33913);
and U34291 (N_34291,N_33804,N_33947);
and U34292 (N_34292,N_33996,N_33642);
or U34293 (N_34293,N_33926,N_33711);
and U34294 (N_34294,N_33554,N_33941);
and U34295 (N_34295,N_33969,N_33666);
nor U34296 (N_34296,N_33922,N_33997);
xnor U34297 (N_34297,N_33603,N_33737);
and U34298 (N_34298,N_33518,N_33636);
and U34299 (N_34299,N_33880,N_33811);
nor U34300 (N_34300,N_33604,N_33819);
nor U34301 (N_34301,N_33859,N_33958);
nor U34302 (N_34302,N_33525,N_33579);
and U34303 (N_34303,N_33629,N_33723);
and U34304 (N_34304,N_33748,N_33762);
nor U34305 (N_34305,N_33683,N_33722);
xor U34306 (N_34306,N_33556,N_33589);
or U34307 (N_34307,N_33552,N_33503);
xor U34308 (N_34308,N_33585,N_33936);
or U34309 (N_34309,N_33753,N_33811);
nor U34310 (N_34310,N_33865,N_33779);
and U34311 (N_34311,N_33931,N_33510);
nand U34312 (N_34312,N_33714,N_33593);
nand U34313 (N_34313,N_33906,N_33659);
and U34314 (N_34314,N_33671,N_33561);
nor U34315 (N_34315,N_33566,N_33778);
and U34316 (N_34316,N_33933,N_33588);
and U34317 (N_34317,N_33928,N_33584);
nor U34318 (N_34318,N_33868,N_33529);
xor U34319 (N_34319,N_33688,N_33950);
nand U34320 (N_34320,N_33662,N_33852);
or U34321 (N_34321,N_33506,N_33645);
xnor U34322 (N_34322,N_33905,N_33858);
nand U34323 (N_34323,N_33773,N_33670);
xor U34324 (N_34324,N_33533,N_33580);
xnor U34325 (N_34325,N_33791,N_33564);
nor U34326 (N_34326,N_33590,N_33848);
xor U34327 (N_34327,N_33940,N_33547);
nand U34328 (N_34328,N_33818,N_33663);
xor U34329 (N_34329,N_33581,N_33589);
xnor U34330 (N_34330,N_33600,N_33586);
xor U34331 (N_34331,N_33896,N_33750);
nand U34332 (N_34332,N_33664,N_33804);
nor U34333 (N_34333,N_33795,N_33897);
and U34334 (N_34334,N_33617,N_33720);
xnor U34335 (N_34335,N_33532,N_33640);
or U34336 (N_34336,N_33521,N_33930);
or U34337 (N_34337,N_33556,N_33767);
or U34338 (N_34338,N_33686,N_33596);
nor U34339 (N_34339,N_33504,N_33558);
and U34340 (N_34340,N_33722,N_33796);
nor U34341 (N_34341,N_33846,N_33888);
xnor U34342 (N_34342,N_33805,N_33641);
nand U34343 (N_34343,N_33740,N_33862);
xor U34344 (N_34344,N_33926,N_33912);
and U34345 (N_34345,N_33513,N_33610);
nor U34346 (N_34346,N_33586,N_33899);
nand U34347 (N_34347,N_33680,N_33545);
xor U34348 (N_34348,N_33796,N_33960);
or U34349 (N_34349,N_33626,N_33877);
or U34350 (N_34350,N_33589,N_33621);
nand U34351 (N_34351,N_33646,N_33895);
and U34352 (N_34352,N_33604,N_33600);
nor U34353 (N_34353,N_33922,N_33728);
and U34354 (N_34354,N_33617,N_33586);
nand U34355 (N_34355,N_33670,N_33504);
nand U34356 (N_34356,N_33652,N_33937);
xnor U34357 (N_34357,N_33719,N_33882);
nand U34358 (N_34358,N_33765,N_33855);
xor U34359 (N_34359,N_33885,N_33752);
xnor U34360 (N_34360,N_33658,N_33837);
or U34361 (N_34361,N_33843,N_33928);
or U34362 (N_34362,N_33663,N_33821);
and U34363 (N_34363,N_33900,N_33873);
and U34364 (N_34364,N_33956,N_33977);
nand U34365 (N_34365,N_33669,N_33943);
nand U34366 (N_34366,N_33878,N_33973);
xnor U34367 (N_34367,N_33819,N_33549);
nand U34368 (N_34368,N_33983,N_33920);
nand U34369 (N_34369,N_33861,N_33563);
xor U34370 (N_34370,N_33527,N_33783);
nor U34371 (N_34371,N_33740,N_33622);
or U34372 (N_34372,N_33703,N_33585);
xnor U34373 (N_34373,N_33513,N_33581);
xnor U34374 (N_34374,N_33831,N_33615);
or U34375 (N_34375,N_33778,N_33933);
and U34376 (N_34376,N_33845,N_33931);
nor U34377 (N_34377,N_33977,N_33692);
or U34378 (N_34378,N_33915,N_33803);
or U34379 (N_34379,N_33800,N_33658);
nand U34380 (N_34380,N_33936,N_33840);
xnor U34381 (N_34381,N_33531,N_33646);
nand U34382 (N_34382,N_33558,N_33789);
nand U34383 (N_34383,N_33984,N_33975);
or U34384 (N_34384,N_33647,N_33807);
nand U34385 (N_34385,N_33696,N_33513);
and U34386 (N_34386,N_33814,N_33971);
xnor U34387 (N_34387,N_33604,N_33984);
nor U34388 (N_34388,N_33943,N_33792);
or U34389 (N_34389,N_33838,N_33583);
or U34390 (N_34390,N_33811,N_33767);
nand U34391 (N_34391,N_33582,N_33877);
or U34392 (N_34392,N_33573,N_33656);
xor U34393 (N_34393,N_33756,N_33699);
nand U34394 (N_34394,N_33708,N_33609);
or U34395 (N_34395,N_33943,N_33768);
xnor U34396 (N_34396,N_33688,N_33698);
xnor U34397 (N_34397,N_33906,N_33619);
and U34398 (N_34398,N_33621,N_33913);
or U34399 (N_34399,N_33892,N_33679);
nor U34400 (N_34400,N_33865,N_33834);
and U34401 (N_34401,N_33706,N_33807);
and U34402 (N_34402,N_33711,N_33885);
or U34403 (N_34403,N_33848,N_33593);
nor U34404 (N_34404,N_33527,N_33824);
nand U34405 (N_34405,N_33864,N_33588);
xor U34406 (N_34406,N_33810,N_33820);
or U34407 (N_34407,N_33805,N_33980);
xnor U34408 (N_34408,N_33959,N_33624);
xor U34409 (N_34409,N_33561,N_33997);
xor U34410 (N_34410,N_33541,N_33931);
nand U34411 (N_34411,N_33809,N_33525);
or U34412 (N_34412,N_33555,N_33653);
or U34413 (N_34413,N_33637,N_33963);
or U34414 (N_34414,N_33897,N_33993);
or U34415 (N_34415,N_33722,N_33878);
or U34416 (N_34416,N_33971,N_33816);
nor U34417 (N_34417,N_33832,N_33973);
or U34418 (N_34418,N_33960,N_33643);
or U34419 (N_34419,N_33738,N_33657);
xor U34420 (N_34420,N_33958,N_33764);
and U34421 (N_34421,N_33836,N_33757);
nand U34422 (N_34422,N_33720,N_33978);
or U34423 (N_34423,N_33669,N_33788);
nand U34424 (N_34424,N_33730,N_33885);
nor U34425 (N_34425,N_33703,N_33636);
and U34426 (N_34426,N_33519,N_33791);
and U34427 (N_34427,N_33785,N_33650);
xor U34428 (N_34428,N_33721,N_33787);
xnor U34429 (N_34429,N_33672,N_33755);
nand U34430 (N_34430,N_33846,N_33682);
nand U34431 (N_34431,N_33671,N_33534);
or U34432 (N_34432,N_33514,N_33955);
xor U34433 (N_34433,N_33566,N_33849);
nor U34434 (N_34434,N_33864,N_33701);
nor U34435 (N_34435,N_33980,N_33755);
and U34436 (N_34436,N_33780,N_33724);
xnor U34437 (N_34437,N_33956,N_33578);
or U34438 (N_34438,N_33652,N_33920);
nand U34439 (N_34439,N_33574,N_33691);
xnor U34440 (N_34440,N_33908,N_33900);
nor U34441 (N_34441,N_33598,N_33788);
nand U34442 (N_34442,N_33693,N_33510);
or U34443 (N_34443,N_33917,N_33852);
or U34444 (N_34444,N_33832,N_33524);
nand U34445 (N_34445,N_33902,N_33968);
or U34446 (N_34446,N_33974,N_33660);
and U34447 (N_34447,N_33669,N_33913);
nand U34448 (N_34448,N_33850,N_33538);
nand U34449 (N_34449,N_33924,N_33886);
nand U34450 (N_34450,N_33640,N_33925);
nor U34451 (N_34451,N_33834,N_33985);
and U34452 (N_34452,N_33537,N_33767);
nand U34453 (N_34453,N_33971,N_33640);
nand U34454 (N_34454,N_33603,N_33785);
or U34455 (N_34455,N_33575,N_33507);
nor U34456 (N_34456,N_33896,N_33546);
and U34457 (N_34457,N_33666,N_33949);
and U34458 (N_34458,N_33942,N_33948);
xor U34459 (N_34459,N_33544,N_33533);
or U34460 (N_34460,N_33936,N_33961);
or U34461 (N_34461,N_33696,N_33561);
nand U34462 (N_34462,N_33699,N_33905);
nor U34463 (N_34463,N_33964,N_33815);
nor U34464 (N_34464,N_33809,N_33643);
or U34465 (N_34465,N_33723,N_33793);
xor U34466 (N_34466,N_33724,N_33694);
xor U34467 (N_34467,N_33982,N_33850);
nand U34468 (N_34468,N_33624,N_33921);
nor U34469 (N_34469,N_33653,N_33946);
xor U34470 (N_34470,N_33549,N_33804);
xor U34471 (N_34471,N_33993,N_33587);
nand U34472 (N_34472,N_33655,N_33521);
and U34473 (N_34473,N_33901,N_33933);
nor U34474 (N_34474,N_33832,N_33697);
or U34475 (N_34475,N_33819,N_33532);
nand U34476 (N_34476,N_33556,N_33823);
xor U34477 (N_34477,N_33826,N_33947);
nand U34478 (N_34478,N_33897,N_33623);
or U34479 (N_34479,N_33639,N_33809);
nor U34480 (N_34480,N_33916,N_33672);
or U34481 (N_34481,N_33975,N_33571);
and U34482 (N_34482,N_33517,N_33662);
nor U34483 (N_34483,N_33906,N_33527);
nand U34484 (N_34484,N_33986,N_33528);
nand U34485 (N_34485,N_33926,N_33583);
or U34486 (N_34486,N_33529,N_33862);
nor U34487 (N_34487,N_33578,N_33781);
and U34488 (N_34488,N_33565,N_33609);
xnor U34489 (N_34489,N_33761,N_33688);
and U34490 (N_34490,N_33561,N_33983);
and U34491 (N_34491,N_33746,N_33714);
or U34492 (N_34492,N_33934,N_33745);
nand U34493 (N_34493,N_33935,N_33908);
nand U34494 (N_34494,N_33669,N_33582);
nor U34495 (N_34495,N_33544,N_33999);
or U34496 (N_34496,N_33815,N_33788);
or U34497 (N_34497,N_33663,N_33612);
and U34498 (N_34498,N_33740,N_33776);
nand U34499 (N_34499,N_33650,N_33605);
nand U34500 (N_34500,N_34332,N_34003);
nand U34501 (N_34501,N_34253,N_34152);
and U34502 (N_34502,N_34281,N_34130);
or U34503 (N_34503,N_34464,N_34167);
and U34504 (N_34504,N_34475,N_34462);
or U34505 (N_34505,N_34151,N_34461);
or U34506 (N_34506,N_34233,N_34055);
nor U34507 (N_34507,N_34449,N_34329);
xnor U34508 (N_34508,N_34368,N_34010);
and U34509 (N_34509,N_34221,N_34319);
or U34510 (N_34510,N_34135,N_34433);
xor U34511 (N_34511,N_34430,N_34350);
nand U34512 (N_34512,N_34246,N_34285);
or U34513 (N_34513,N_34089,N_34240);
nand U34514 (N_34514,N_34238,N_34157);
xor U34515 (N_34515,N_34176,N_34218);
and U34516 (N_34516,N_34195,N_34208);
xnor U34517 (N_34517,N_34276,N_34473);
or U34518 (N_34518,N_34123,N_34125);
or U34519 (N_34519,N_34407,N_34244);
xor U34520 (N_34520,N_34408,N_34096);
nor U34521 (N_34521,N_34297,N_34439);
or U34522 (N_34522,N_34454,N_34267);
or U34523 (N_34523,N_34339,N_34302);
or U34524 (N_34524,N_34043,N_34259);
and U34525 (N_34525,N_34357,N_34292);
nand U34526 (N_34526,N_34274,N_34242);
xnor U34527 (N_34527,N_34039,N_34250);
or U34528 (N_34528,N_34134,N_34248);
nor U34529 (N_34529,N_34049,N_34009);
or U34530 (N_34530,N_34303,N_34088);
nor U34531 (N_34531,N_34066,N_34149);
and U34532 (N_34532,N_34442,N_34094);
or U34533 (N_34533,N_34306,N_34150);
nor U34534 (N_34534,N_34204,N_34323);
nor U34535 (N_34535,N_34298,N_34355);
or U34536 (N_34536,N_34405,N_34166);
nor U34537 (N_34537,N_34177,N_34024);
nand U34538 (N_34538,N_34075,N_34227);
nor U34539 (N_34539,N_34359,N_34448);
xor U34540 (N_34540,N_34373,N_34018);
nor U34541 (N_34541,N_34162,N_34182);
nor U34542 (N_34542,N_34370,N_34211);
xnor U34543 (N_34543,N_34365,N_34158);
nand U34544 (N_34544,N_34418,N_34087);
nor U34545 (N_34545,N_34327,N_34366);
nand U34546 (N_34546,N_34005,N_34097);
nor U34547 (N_34547,N_34065,N_34443);
or U34548 (N_34548,N_34169,N_34254);
nor U34549 (N_34549,N_34232,N_34121);
nor U34550 (N_34550,N_34498,N_34262);
xnor U34551 (N_34551,N_34495,N_34452);
nor U34552 (N_34552,N_34266,N_34273);
xor U34553 (N_34553,N_34189,N_34423);
xnor U34554 (N_34554,N_34004,N_34174);
and U34555 (N_34555,N_34496,N_34386);
xnor U34556 (N_34556,N_34404,N_34336);
and U34557 (N_34557,N_34059,N_34489);
and U34558 (N_34558,N_34234,N_34201);
nand U34559 (N_34559,N_34486,N_34098);
xor U34560 (N_34560,N_34388,N_34035);
nor U34561 (N_34561,N_34426,N_34138);
or U34562 (N_34562,N_34184,N_34132);
nand U34563 (N_34563,N_34012,N_34385);
nor U34564 (N_34564,N_34367,N_34160);
nand U34565 (N_34565,N_34422,N_34105);
nor U34566 (N_34566,N_34054,N_34406);
and U34567 (N_34567,N_34395,N_34110);
xor U34568 (N_34568,N_34450,N_34057);
and U34569 (N_34569,N_34076,N_34081);
xor U34570 (N_34570,N_34399,N_34068);
xor U34571 (N_34571,N_34341,N_34223);
xnor U34572 (N_34572,N_34008,N_34164);
nand U34573 (N_34573,N_34456,N_34324);
nor U34574 (N_34574,N_34479,N_34095);
and U34575 (N_34575,N_34375,N_34356);
xor U34576 (N_34576,N_34237,N_34256);
xor U34577 (N_34577,N_34251,N_34014);
or U34578 (N_34578,N_34497,N_34316);
nor U34579 (N_34579,N_34052,N_34222);
or U34580 (N_34580,N_34340,N_34435);
or U34581 (N_34581,N_34212,N_34192);
xor U34582 (N_34582,N_34457,N_34128);
nand U34583 (N_34583,N_34438,N_34447);
and U34584 (N_34584,N_34321,N_34277);
nor U34585 (N_34585,N_34265,N_34021);
nand U34586 (N_34586,N_34213,N_34133);
and U34587 (N_34587,N_34330,N_34136);
nand U34588 (N_34588,N_34034,N_34451);
or U34589 (N_34589,N_34137,N_34016);
nor U34590 (N_34590,N_34352,N_34427);
nor U34591 (N_34591,N_34038,N_34112);
xnor U34592 (N_34592,N_34127,N_34476);
and U34593 (N_34593,N_34307,N_34113);
nor U34594 (N_34594,N_34117,N_34187);
and U34595 (N_34595,N_34129,N_34459);
nor U34596 (N_34596,N_34353,N_34190);
or U34597 (N_34597,N_34420,N_34317);
or U34598 (N_34598,N_34069,N_34205);
and U34599 (N_34599,N_34348,N_34022);
xor U34600 (N_34600,N_34286,N_34171);
or U34601 (N_34601,N_34255,N_34122);
and U34602 (N_34602,N_34284,N_34280);
xor U34603 (N_34603,N_34453,N_34301);
or U34604 (N_34604,N_34031,N_34421);
nor U34605 (N_34605,N_34020,N_34002);
xor U34606 (N_34606,N_34099,N_34109);
and U34607 (N_34607,N_34384,N_34100);
and U34608 (N_34608,N_34419,N_34156);
and U34609 (N_34609,N_34436,N_34261);
nor U34610 (N_34610,N_34119,N_34041);
nand U34611 (N_34611,N_34104,N_34376);
xnor U34612 (N_34612,N_34397,N_34230);
or U34613 (N_34613,N_34334,N_34092);
and U34614 (N_34614,N_34379,N_34102);
or U34615 (N_34615,N_34412,N_34007);
nand U34616 (N_34616,N_34252,N_34091);
and U34617 (N_34617,N_34207,N_34358);
or U34618 (N_34618,N_34155,N_34432);
nand U34619 (N_34619,N_34175,N_34070);
xor U34620 (N_34620,N_34260,N_34470);
and U34621 (N_34621,N_34465,N_34165);
and U34622 (N_34622,N_34268,N_34335);
nor U34623 (N_34623,N_34484,N_34483);
and U34624 (N_34624,N_34377,N_34120);
nand U34625 (N_34625,N_34400,N_34090);
nand U34626 (N_34626,N_34445,N_34061);
xnor U34627 (N_34627,N_34325,N_34383);
or U34628 (N_34628,N_34172,N_34338);
nand U34629 (N_34629,N_34111,N_34173);
or U34630 (N_34630,N_34460,N_34093);
nor U34631 (N_34631,N_34401,N_34351);
nor U34632 (N_34632,N_34142,N_34387);
and U34633 (N_34633,N_34314,N_34344);
or U34634 (N_34634,N_34469,N_34287);
or U34635 (N_34635,N_34296,N_34243);
nor U34636 (N_34636,N_34131,N_34163);
or U34637 (N_34637,N_34214,N_34179);
xor U34638 (N_34638,N_34369,N_34310);
nor U34639 (N_34639,N_34033,N_34200);
and U34640 (N_34640,N_34393,N_34074);
xnor U34641 (N_34641,N_34145,N_34029);
xnor U34642 (N_34642,N_34343,N_34019);
or U34643 (N_34643,N_34288,N_34312);
and U34644 (N_34644,N_34275,N_34488);
nand U34645 (N_34645,N_34360,N_34047);
nor U34646 (N_34646,N_34032,N_34236);
or U34647 (N_34647,N_34026,N_34382);
or U34648 (N_34648,N_34023,N_34493);
nor U34649 (N_34649,N_34206,N_34231);
nand U34650 (N_34650,N_34101,N_34185);
and U34651 (N_34651,N_34264,N_34381);
nand U34652 (N_34652,N_34467,N_34389);
and U34653 (N_34653,N_34478,N_34417);
and U34654 (N_34654,N_34115,N_34114);
xnor U34655 (N_34655,N_34084,N_34154);
nor U34656 (N_34656,N_34180,N_34202);
or U34657 (N_34657,N_34108,N_34271);
and U34658 (N_34658,N_34082,N_34027);
nor U34659 (N_34659,N_34300,N_34245);
nor U34660 (N_34660,N_34337,N_34079);
or U34661 (N_34661,N_34073,N_34148);
or U34662 (N_34662,N_34028,N_34001);
or U34663 (N_34663,N_34000,N_34153);
nor U34664 (N_34664,N_34224,N_34394);
nand U34665 (N_34665,N_34485,N_34480);
nand U34666 (N_34666,N_34402,N_34235);
nand U34667 (N_34667,N_34146,N_34058);
nand U34668 (N_34668,N_34015,N_34072);
nand U34669 (N_34669,N_34046,N_34116);
nand U34670 (N_34670,N_34295,N_34416);
and U34671 (N_34671,N_34067,N_34311);
xor U34672 (N_34672,N_34144,N_34309);
and U34673 (N_34673,N_34396,N_34168);
nand U34674 (N_34674,N_34203,N_34025);
xor U34675 (N_34675,N_34198,N_34499);
nor U34676 (N_34676,N_34282,N_34345);
nor U34677 (N_34677,N_34291,N_34143);
and U34678 (N_34678,N_34491,N_34354);
or U34679 (N_34679,N_34349,N_34380);
and U34680 (N_34680,N_34414,N_34077);
nand U34681 (N_34681,N_34347,N_34210);
or U34682 (N_34682,N_34037,N_34147);
or U34683 (N_34683,N_34318,N_34126);
xor U34684 (N_34684,N_34225,N_34279);
nor U34685 (N_34685,N_34036,N_34362);
nand U34686 (N_34686,N_34342,N_34371);
and U34687 (N_34687,N_34216,N_34424);
nor U34688 (N_34688,N_34322,N_34199);
xor U34689 (N_34689,N_34328,N_34263);
xnor U34690 (N_34690,N_34410,N_34378);
or U34691 (N_34691,N_34006,N_34346);
and U34692 (N_34692,N_34080,N_34429);
nand U34693 (N_34693,N_34425,N_34051);
nor U34694 (N_34694,N_34183,N_34226);
and U34695 (N_34695,N_34188,N_34209);
nor U34696 (N_34696,N_34060,N_34477);
or U34697 (N_34697,N_34078,N_34299);
or U34698 (N_34698,N_34444,N_34392);
or U34699 (N_34699,N_34186,N_34331);
and U34700 (N_34700,N_34124,N_34490);
xnor U34701 (N_34701,N_34494,N_34159);
xor U34702 (N_34702,N_34305,N_34220);
and U34703 (N_34703,N_34468,N_34103);
and U34704 (N_34704,N_34178,N_34455);
nand U34705 (N_34705,N_34118,N_34215);
nor U34706 (N_34706,N_34193,N_34239);
xnor U34707 (N_34707,N_34481,N_34106);
xor U34708 (N_34708,N_34217,N_34161);
or U34709 (N_34709,N_34030,N_34283);
and U34710 (N_34710,N_34403,N_34441);
xor U34711 (N_34711,N_34472,N_34063);
and U34712 (N_34712,N_34413,N_34017);
and U34713 (N_34713,N_34170,N_34290);
or U34714 (N_34714,N_34040,N_34482);
xnor U34715 (N_34715,N_34466,N_34042);
nand U34716 (N_34716,N_34431,N_34194);
and U34717 (N_34717,N_34440,N_34411);
nand U34718 (N_34718,N_34249,N_34071);
and U34719 (N_34719,N_34278,N_34053);
or U34720 (N_34720,N_34241,N_34308);
and U34721 (N_34721,N_34247,N_34333);
nand U34722 (N_34722,N_34196,N_34228);
xor U34723 (N_34723,N_34409,N_34013);
xor U34724 (N_34724,N_34056,N_34269);
xor U34725 (N_34725,N_34458,N_34086);
or U34726 (N_34726,N_34229,N_34390);
nor U34727 (N_34727,N_34320,N_34391);
or U34728 (N_34728,N_34107,N_34304);
and U34729 (N_34729,N_34374,N_34257);
nor U34730 (N_34730,N_34258,N_34045);
or U34731 (N_34731,N_34474,N_34083);
xnor U34732 (N_34732,N_34313,N_34398);
nor U34733 (N_34733,N_34050,N_34294);
and U34734 (N_34734,N_34181,N_34270);
xnor U34735 (N_34735,N_34141,N_34062);
nand U34736 (N_34736,N_34492,N_34487);
or U34737 (N_34737,N_34363,N_34372);
or U34738 (N_34738,N_34463,N_34434);
nand U34739 (N_34739,N_34140,N_34044);
and U34740 (N_34740,N_34085,N_34415);
xnor U34741 (N_34741,N_34437,N_34064);
xor U34742 (N_34742,N_34361,N_34293);
xor U34743 (N_34743,N_34139,N_34315);
nor U34744 (N_34744,N_34272,N_34428);
nand U34745 (N_34745,N_34191,N_34364);
nand U34746 (N_34746,N_34048,N_34219);
xnor U34747 (N_34747,N_34011,N_34326);
or U34748 (N_34748,N_34197,N_34289);
and U34749 (N_34749,N_34446,N_34471);
nand U34750 (N_34750,N_34385,N_34013);
or U34751 (N_34751,N_34255,N_34421);
nor U34752 (N_34752,N_34028,N_34179);
xor U34753 (N_34753,N_34222,N_34289);
or U34754 (N_34754,N_34463,N_34432);
or U34755 (N_34755,N_34306,N_34358);
nor U34756 (N_34756,N_34412,N_34110);
nor U34757 (N_34757,N_34168,N_34250);
xnor U34758 (N_34758,N_34103,N_34498);
and U34759 (N_34759,N_34463,N_34400);
and U34760 (N_34760,N_34367,N_34306);
and U34761 (N_34761,N_34267,N_34473);
nor U34762 (N_34762,N_34172,N_34240);
nor U34763 (N_34763,N_34211,N_34001);
nor U34764 (N_34764,N_34006,N_34297);
nand U34765 (N_34765,N_34384,N_34483);
nand U34766 (N_34766,N_34135,N_34224);
nor U34767 (N_34767,N_34387,N_34013);
nand U34768 (N_34768,N_34150,N_34464);
nor U34769 (N_34769,N_34247,N_34039);
and U34770 (N_34770,N_34243,N_34149);
and U34771 (N_34771,N_34389,N_34143);
or U34772 (N_34772,N_34246,N_34383);
nor U34773 (N_34773,N_34090,N_34357);
nand U34774 (N_34774,N_34224,N_34002);
or U34775 (N_34775,N_34130,N_34147);
or U34776 (N_34776,N_34425,N_34139);
xnor U34777 (N_34777,N_34413,N_34215);
and U34778 (N_34778,N_34413,N_34284);
xor U34779 (N_34779,N_34445,N_34007);
nor U34780 (N_34780,N_34173,N_34276);
xor U34781 (N_34781,N_34295,N_34160);
or U34782 (N_34782,N_34472,N_34197);
nor U34783 (N_34783,N_34425,N_34213);
and U34784 (N_34784,N_34317,N_34352);
nand U34785 (N_34785,N_34345,N_34429);
or U34786 (N_34786,N_34063,N_34214);
and U34787 (N_34787,N_34414,N_34078);
nand U34788 (N_34788,N_34193,N_34348);
or U34789 (N_34789,N_34267,N_34363);
or U34790 (N_34790,N_34233,N_34330);
and U34791 (N_34791,N_34312,N_34461);
nor U34792 (N_34792,N_34234,N_34065);
and U34793 (N_34793,N_34327,N_34352);
or U34794 (N_34794,N_34336,N_34416);
nand U34795 (N_34795,N_34077,N_34388);
or U34796 (N_34796,N_34243,N_34133);
xor U34797 (N_34797,N_34291,N_34321);
or U34798 (N_34798,N_34443,N_34335);
xor U34799 (N_34799,N_34232,N_34153);
and U34800 (N_34800,N_34433,N_34353);
nand U34801 (N_34801,N_34431,N_34449);
and U34802 (N_34802,N_34082,N_34400);
nand U34803 (N_34803,N_34263,N_34408);
or U34804 (N_34804,N_34262,N_34461);
nand U34805 (N_34805,N_34329,N_34419);
nand U34806 (N_34806,N_34100,N_34406);
xnor U34807 (N_34807,N_34172,N_34281);
xor U34808 (N_34808,N_34037,N_34349);
nand U34809 (N_34809,N_34433,N_34004);
or U34810 (N_34810,N_34141,N_34491);
nor U34811 (N_34811,N_34412,N_34481);
or U34812 (N_34812,N_34313,N_34032);
nor U34813 (N_34813,N_34090,N_34427);
xnor U34814 (N_34814,N_34196,N_34062);
nor U34815 (N_34815,N_34342,N_34162);
and U34816 (N_34816,N_34051,N_34237);
or U34817 (N_34817,N_34013,N_34281);
xnor U34818 (N_34818,N_34046,N_34212);
nor U34819 (N_34819,N_34482,N_34385);
nand U34820 (N_34820,N_34093,N_34438);
xnor U34821 (N_34821,N_34241,N_34003);
nand U34822 (N_34822,N_34481,N_34388);
and U34823 (N_34823,N_34277,N_34108);
xnor U34824 (N_34824,N_34134,N_34307);
and U34825 (N_34825,N_34058,N_34028);
nand U34826 (N_34826,N_34066,N_34222);
nand U34827 (N_34827,N_34398,N_34266);
and U34828 (N_34828,N_34084,N_34436);
nand U34829 (N_34829,N_34334,N_34082);
xor U34830 (N_34830,N_34118,N_34496);
and U34831 (N_34831,N_34401,N_34499);
and U34832 (N_34832,N_34062,N_34087);
and U34833 (N_34833,N_34269,N_34355);
nand U34834 (N_34834,N_34065,N_34000);
nand U34835 (N_34835,N_34393,N_34245);
xor U34836 (N_34836,N_34156,N_34144);
nand U34837 (N_34837,N_34362,N_34122);
or U34838 (N_34838,N_34051,N_34246);
nand U34839 (N_34839,N_34237,N_34308);
xnor U34840 (N_34840,N_34295,N_34069);
nor U34841 (N_34841,N_34352,N_34238);
nand U34842 (N_34842,N_34136,N_34441);
or U34843 (N_34843,N_34453,N_34465);
nor U34844 (N_34844,N_34037,N_34446);
or U34845 (N_34845,N_34407,N_34032);
nand U34846 (N_34846,N_34371,N_34443);
nor U34847 (N_34847,N_34235,N_34055);
nor U34848 (N_34848,N_34319,N_34344);
and U34849 (N_34849,N_34082,N_34338);
nor U34850 (N_34850,N_34103,N_34288);
or U34851 (N_34851,N_34362,N_34059);
and U34852 (N_34852,N_34488,N_34343);
or U34853 (N_34853,N_34254,N_34039);
nand U34854 (N_34854,N_34269,N_34311);
nor U34855 (N_34855,N_34459,N_34445);
xnor U34856 (N_34856,N_34331,N_34362);
nor U34857 (N_34857,N_34134,N_34428);
nor U34858 (N_34858,N_34138,N_34389);
nand U34859 (N_34859,N_34154,N_34065);
and U34860 (N_34860,N_34351,N_34211);
nor U34861 (N_34861,N_34410,N_34131);
and U34862 (N_34862,N_34068,N_34184);
nor U34863 (N_34863,N_34182,N_34469);
and U34864 (N_34864,N_34255,N_34240);
nand U34865 (N_34865,N_34067,N_34101);
and U34866 (N_34866,N_34498,N_34453);
or U34867 (N_34867,N_34278,N_34154);
or U34868 (N_34868,N_34470,N_34116);
nand U34869 (N_34869,N_34099,N_34288);
or U34870 (N_34870,N_34211,N_34373);
nor U34871 (N_34871,N_34229,N_34322);
nand U34872 (N_34872,N_34041,N_34127);
and U34873 (N_34873,N_34006,N_34210);
and U34874 (N_34874,N_34427,N_34103);
or U34875 (N_34875,N_34203,N_34040);
nor U34876 (N_34876,N_34179,N_34392);
or U34877 (N_34877,N_34286,N_34419);
or U34878 (N_34878,N_34106,N_34475);
or U34879 (N_34879,N_34022,N_34139);
xor U34880 (N_34880,N_34423,N_34406);
nor U34881 (N_34881,N_34497,N_34007);
and U34882 (N_34882,N_34225,N_34442);
nand U34883 (N_34883,N_34359,N_34181);
nand U34884 (N_34884,N_34284,N_34463);
nand U34885 (N_34885,N_34315,N_34134);
or U34886 (N_34886,N_34099,N_34122);
or U34887 (N_34887,N_34411,N_34347);
nand U34888 (N_34888,N_34453,N_34206);
and U34889 (N_34889,N_34136,N_34127);
or U34890 (N_34890,N_34325,N_34280);
or U34891 (N_34891,N_34404,N_34432);
and U34892 (N_34892,N_34452,N_34146);
or U34893 (N_34893,N_34480,N_34241);
or U34894 (N_34894,N_34387,N_34190);
xor U34895 (N_34895,N_34315,N_34235);
nand U34896 (N_34896,N_34295,N_34320);
nand U34897 (N_34897,N_34397,N_34338);
or U34898 (N_34898,N_34061,N_34209);
xor U34899 (N_34899,N_34368,N_34373);
and U34900 (N_34900,N_34417,N_34242);
xor U34901 (N_34901,N_34037,N_34295);
and U34902 (N_34902,N_34309,N_34182);
nand U34903 (N_34903,N_34037,N_34376);
nand U34904 (N_34904,N_34060,N_34063);
and U34905 (N_34905,N_34431,N_34236);
nand U34906 (N_34906,N_34312,N_34371);
nor U34907 (N_34907,N_34406,N_34097);
or U34908 (N_34908,N_34160,N_34380);
nand U34909 (N_34909,N_34229,N_34495);
nand U34910 (N_34910,N_34184,N_34379);
xor U34911 (N_34911,N_34297,N_34320);
or U34912 (N_34912,N_34257,N_34132);
xnor U34913 (N_34913,N_34497,N_34213);
and U34914 (N_34914,N_34413,N_34333);
nand U34915 (N_34915,N_34412,N_34301);
nand U34916 (N_34916,N_34483,N_34493);
nand U34917 (N_34917,N_34216,N_34488);
and U34918 (N_34918,N_34173,N_34458);
nand U34919 (N_34919,N_34403,N_34205);
xnor U34920 (N_34920,N_34376,N_34270);
and U34921 (N_34921,N_34216,N_34099);
nand U34922 (N_34922,N_34370,N_34167);
and U34923 (N_34923,N_34053,N_34363);
nor U34924 (N_34924,N_34405,N_34230);
nor U34925 (N_34925,N_34418,N_34310);
or U34926 (N_34926,N_34023,N_34083);
xnor U34927 (N_34927,N_34253,N_34162);
nor U34928 (N_34928,N_34180,N_34482);
nand U34929 (N_34929,N_34002,N_34100);
and U34930 (N_34930,N_34250,N_34420);
xnor U34931 (N_34931,N_34441,N_34475);
nor U34932 (N_34932,N_34485,N_34093);
nor U34933 (N_34933,N_34317,N_34048);
and U34934 (N_34934,N_34084,N_34415);
nand U34935 (N_34935,N_34299,N_34381);
or U34936 (N_34936,N_34478,N_34314);
or U34937 (N_34937,N_34312,N_34069);
nand U34938 (N_34938,N_34413,N_34157);
nor U34939 (N_34939,N_34135,N_34497);
nor U34940 (N_34940,N_34369,N_34182);
nor U34941 (N_34941,N_34159,N_34276);
or U34942 (N_34942,N_34360,N_34448);
and U34943 (N_34943,N_34457,N_34476);
xor U34944 (N_34944,N_34192,N_34385);
nor U34945 (N_34945,N_34076,N_34126);
or U34946 (N_34946,N_34237,N_34312);
nand U34947 (N_34947,N_34204,N_34111);
xnor U34948 (N_34948,N_34179,N_34030);
nand U34949 (N_34949,N_34405,N_34315);
nand U34950 (N_34950,N_34057,N_34294);
nand U34951 (N_34951,N_34173,N_34196);
and U34952 (N_34952,N_34265,N_34217);
nor U34953 (N_34953,N_34133,N_34186);
or U34954 (N_34954,N_34447,N_34078);
and U34955 (N_34955,N_34498,N_34239);
nor U34956 (N_34956,N_34154,N_34197);
or U34957 (N_34957,N_34331,N_34279);
nor U34958 (N_34958,N_34387,N_34304);
and U34959 (N_34959,N_34246,N_34300);
nand U34960 (N_34960,N_34442,N_34049);
nor U34961 (N_34961,N_34247,N_34394);
nand U34962 (N_34962,N_34451,N_34420);
nor U34963 (N_34963,N_34192,N_34012);
and U34964 (N_34964,N_34300,N_34019);
nand U34965 (N_34965,N_34119,N_34204);
or U34966 (N_34966,N_34171,N_34085);
and U34967 (N_34967,N_34403,N_34201);
xnor U34968 (N_34968,N_34057,N_34251);
nor U34969 (N_34969,N_34133,N_34222);
or U34970 (N_34970,N_34327,N_34485);
nand U34971 (N_34971,N_34437,N_34024);
or U34972 (N_34972,N_34146,N_34095);
or U34973 (N_34973,N_34446,N_34447);
and U34974 (N_34974,N_34122,N_34023);
and U34975 (N_34975,N_34443,N_34368);
or U34976 (N_34976,N_34472,N_34285);
or U34977 (N_34977,N_34276,N_34306);
nor U34978 (N_34978,N_34469,N_34322);
xnor U34979 (N_34979,N_34243,N_34439);
nor U34980 (N_34980,N_34001,N_34279);
and U34981 (N_34981,N_34054,N_34466);
nor U34982 (N_34982,N_34059,N_34192);
or U34983 (N_34983,N_34188,N_34035);
nand U34984 (N_34984,N_34057,N_34152);
xor U34985 (N_34985,N_34208,N_34157);
xnor U34986 (N_34986,N_34454,N_34496);
nand U34987 (N_34987,N_34089,N_34235);
nor U34988 (N_34988,N_34168,N_34307);
or U34989 (N_34989,N_34142,N_34029);
xnor U34990 (N_34990,N_34006,N_34172);
and U34991 (N_34991,N_34033,N_34437);
nor U34992 (N_34992,N_34335,N_34295);
or U34993 (N_34993,N_34065,N_34097);
nand U34994 (N_34994,N_34186,N_34378);
nor U34995 (N_34995,N_34023,N_34191);
nand U34996 (N_34996,N_34292,N_34029);
nand U34997 (N_34997,N_34370,N_34343);
nor U34998 (N_34998,N_34168,N_34047);
and U34999 (N_34999,N_34316,N_34142);
or U35000 (N_35000,N_34834,N_34773);
nand U35001 (N_35001,N_34591,N_34764);
and U35002 (N_35002,N_34806,N_34813);
or U35003 (N_35003,N_34787,N_34845);
nand U35004 (N_35004,N_34724,N_34723);
nand U35005 (N_35005,N_34730,N_34585);
xnor U35006 (N_35006,N_34652,N_34857);
nand U35007 (N_35007,N_34877,N_34866);
and U35008 (N_35008,N_34710,N_34781);
nand U35009 (N_35009,N_34627,N_34970);
or U35010 (N_35010,N_34955,N_34913);
xnor U35011 (N_35011,N_34717,N_34934);
and U35012 (N_35012,N_34986,N_34611);
xor U35013 (N_35013,N_34725,N_34975);
nor U35014 (N_35014,N_34782,N_34729);
or U35015 (N_35015,N_34509,N_34593);
or U35016 (N_35016,N_34543,N_34912);
xnor U35017 (N_35017,N_34742,N_34830);
or U35018 (N_35018,N_34760,N_34969);
nor U35019 (N_35019,N_34529,N_34979);
or U35020 (N_35020,N_34902,N_34553);
nor U35021 (N_35021,N_34536,N_34985);
nand U35022 (N_35022,N_34793,N_34949);
xor U35023 (N_35023,N_34511,N_34897);
nand U35024 (N_35024,N_34712,N_34868);
or U35025 (N_35025,N_34768,N_34967);
or U35026 (N_35026,N_34847,N_34735);
nand U35027 (N_35027,N_34844,N_34798);
nand U35028 (N_35028,N_34719,N_34555);
xnor U35029 (N_35029,N_34930,N_34921);
nand U35030 (N_35030,N_34636,N_34508);
xnor U35031 (N_35031,N_34947,N_34524);
nand U35032 (N_35032,N_34637,N_34523);
xor U35033 (N_35033,N_34766,N_34562);
or U35034 (N_35034,N_34968,N_34561);
and U35035 (N_35035,N_34993,N_34681);
and U35036 (N_35036,N_34859,N_34563);
nand U35037 (N_35037,N_34937,N_34978);
xor U35038 (N_35038,N_34948,N_34505);
or U35039 (N_35039,N_34858,N_34926);
and U35040 (N_35040,N_34596,N_34905);
or U35041 (N_35041,N_34595,N_34989);
nand U35042 (N_35042,N_34670,N_34738);
nor U35043 (N_35043,N_34826,N_34500);
xor U35044 (N_35044,N_34884,N_34539);
nor U35045 (N_35045,N_34871,N_34656);
nand U35046 (N_35046,N_34842,N_34833);
nor U35047 (N_35047,N_34927,N_34588);
xnor U35048 (N_35048,N_34966,N_34657);
xor U35049 (N_35049,N_34513,N_34982);
xnor U35050 (N_35050,N_34522,N_34566);
xor U35051 (N_35051,N_34882,N_34554);
xor U35052 (N_35052,N_34914,N_34852);
and U35053 (N_35053,N_34853,N_34686);
xnor U35054 (N_35054,N_34574,N_34805);
and U35055 (N_35055,N_34936,N_34518);
xor U35056 (N_35056,N_34503,N_34980);
xnor U35057 (N_35057,N_34890,N_34922);
nand U35058 (N_35058,N_34789,N_34706);
xor U35059 (N_35059,N_34716,N_34749);
xnor U35060 (N_35060,N_34808,N_34869);
xor U35061 (N_35061,N_34973,N_34722);
and U35062 (N_35062,N_34942,N_34624);
xnor U35063 (N_35063,N_34567,N_34786);
nor U35064 (N_35064,N_34707,N_34771);
and U35065 (N_35065,N_34501,N_34647);
xnor U35066 (N_35066,N_34759,N_34795);
xnor U35067 (N_35067,N_34824,N_34526);
or U35068 (N_35068,N_34514,N_34662);
nand U35069 (N_35069,N_34661,N_34642);
xor U35070 (N_35070,N_34996,N_34675);
xor U35071 (N_35071,N_34639,N_34770);
nand U35072 (N_35072,N_34757,N_34878);
and U35073 (N_35073,N_34856,N_34872);
nor U35074 (N_35074,N_34812,N_34739);
and U35075 (N_35075,N_34688,N_34690);
nand U35076 (N_35076,N_34635,N_34676);
or U35077 (N_35077,N_34630,N_34646);
nor U35078 (N_35078,N_34836,N_34535);
nor U35079 (N_35079,N_34840,N_34888);
nand U35080 (N_35080,N_34744,N_34849);
xnor U35081 (N_35081,N_34791,N_34964);
and U35082 (N_35082,N_34557,N_34817);
xor U35083 (N_35083,N_34677,N_34577);
and U35084 (N_35084,N_34838,N_34565);
nand U35085 (N_35085,N_34599,N_34792);
nor U35086 (N_35086,N_34820,N_34620);
nor U35087 (N_35087,N_34909,N_34622);
xnor U35088 (N_35088,N_34659,N_34552);
and U35089 (N_35089,N_34579,N_34850);
nor U35090 (N_35090,N_34726,N_34831);
or U35091 (N_35091,N_34648,N_34502);
xor U35092 (N_35092,N_34765,N_34545);
xor U35093 (N_35093,N_34976,N_34504);
xor U35094 (N_35094,N_34899,N_34740);
and U35095 (N_35095,N_34772,N_34959);
nor U35096 (N_35096,N_34816,N_34821);
and U35097 (N_35097,N_34839,N_34667);
or U35098 (N_35098,N_34741,N_34633);
nand U35099 (N_35099,N_34860,N_34533);
or U35100 (N_35100,N_34713,N_34534);
nor U35101 (N_35101,N_34699,N_34705);
nand U35102 (N_35102,N_34783,N_34893);
and U35103 (N_35103,N_34923,N_34758);
nand U35104 (N_35104,N_34907,N_34779);
or U35105 (N_35105,N_34692,N_34972);
nor U35106 (N_35106,N_34924,N_34837);
and U35107 (N_35107,N_34752,N_34901);
nand U35108 (N_35108,N_34804,N_34682);
and U35109 (N_35109,N_34754,N_34544);
nor U35110 (N_35110,N_34977,N_34651);
or U35111 (N_35111,N_34800,N_34687);
or U35112 (N_35112,N_34775,N_34672);
or U35113 (N_35113,N_34634,N_34721);
nor U35114 (N_35114,N_34874,N_34887);
or U35115 (N_35115,N_34896,N_34917);
nor U35116 (N_35116,N_34586,N_34680);
xnor U35117 (N_35117,N_34609,N_34911);
nand U35118 (N_35118,N_34932,N_34701);
or U35119 (N_35119,N_34568,N_34892);
xor U35120 (N_35120,N_34929,N_34540);
and U35121 (N_35121,N_34573,N_34548);
nand U35122 (N_35122,N_34731,N_34650);
and U35123 (N_35123,N_34815,N_34935);
nand U35124 (N_35124,N_34718,N_34698);
nand U35125 (N_35125,N_34530,N_34835);
xor U35126 (N_35126,N_34691,N_34547);
nand U35127 (N_35127,N_34875,N_34737);
nor U35128 (N_35128,N_34617,N_34963);
or U35129 (N_35129,N_34525,N_34537);
xnor U35130 (N_35130,N_34843,N_34974);
xor U35131 (N_35131,N_34761,N_34998);
and U35132 (N_35132,N_34928,N_34623);
xor U35133 (N_35133,N_34751,N_34981);
and U35134 (N_35134,N_34931,N_34769);
or U35135 (N_35135,N_34632,N_34891);
xor U35136 (N_35136,N_34876,N_34714);
xor U35137 (N_35137,N_34753,N_34863);
or U35138 (N_35138,N_34983,N_34668);
xor U35139 (N_35139,N_34580,N_34546);
and U35140 (N_35140,N_34910,N_34736);
xor U35141 (N_35141,N_34994,N_34810);
or U35142 (N_35142,N_34908,N_34696);
xor U35143 (N_35143,N_34818,N_34621);
xor U35144 (N_35144,N_34743,N_34802);
xor U35145 (N_35145,N_34702,N_34576);
nor U35146 (N_35146,N_34885,N_34645);
nand U35147 (N_35147,N_34814,N_34569);
or U35148 (N_35148,N_34987,N_34946);
nand U35149 (N_35149,N_34861,N_34697);
nand U35150 (N_35150,N_34807,N_34660);
nand U35151 (N_35151,N_34822,N_34532);
and U35152 (N_35152,N_34515,N_34704);
xnor U35153 (N_35153,N_34803,N_34665);
nor U35154 (N_35154,N_34747,N_34506);
nor U35155 (N_35155,N_34819,N_34711);
and U35156 (N_35156,N_34708,N_34799);
and U35157 (N_35157,N_34767,N_34828);
nor U35158 (N_35158,N_34797,N_34578);
nor U35159 (N_35159,N_34538,N_34776);
or U35160 (N_35160,N_34616,N_34965);
nor U35161 (N_35161,N_34894,N_34572);
or U35162 (N_35162,N_34881,N_34763);
or U35163 (N_35163,N_34825,N_34658);
nand U35164 (N_35164,N_34631,N_34582);
xor U35165 (N_35165,N_34794,N_34683);
or U35166 (N_35166,N_34862,N_34939);
or U35167 (N_35167,N_34956,N_34558);
nor U35168 (N_35168,N_34746,N_34906);
nand U35169 (N_35169,N_34614,N_34715);
and U35170 (N_35170,N_34777,N_34755);
and U35171 (N_35171,N_34694,N_34610);
or U35172 (N_35172,N_34733,N_34748);
and U35173 (N_35173,N_34603,N_34619);
and U35174 (N_35174,N_34678,N_34612);
nand U35175 (N_35175,N_34879,N_34564);
and U35176 (N_35176,N_34602,N_34527);
or U35177 (N_35177,N_34531,N_34992);
and U35178 (N_35178,N_34867,N_34541);
nand U35179 (N_35179,N_34643,N_34679);
xnor U35180 (N_35180,N_34517,N_34615);
nand U35181 (N_35181,N_34920,N_34734);
or U35182 (N_35182,N_34957,N_34629);
xor U35183 (N_35183,N_34550,N_34542);
xnor U35184 (N_35184,N_34883,N_34709);
xor U35185 (N_35185,N_34832,N_34960);
xnor U35186 (N_35186,N_34940,N_34961);
xnor U35187 (N_35187,N_34841,N_34570);
and U35188 (N_35188,N_34951,N_34933);
nand U35189 (N_35189,N_34870,N_34811);
and U35190 (N_35190,N_34848,N_34915);
and U35191 (N_35191,N_34944,N_34809);
nor U35192 (N_35192,N_34594,N_34598);
nand U35193 (N_35193,N_34575,N_34606);
nand U35194 (N_35194,N_34674,N_34851);
and U35195 (N_35195,N_34995,N_34886);
or U35196 (N_35196,N_34762,N_34512);
nor U35197 (N_35197,N_34903,N_34855);
and U35198 (N_35198,N_34516,N_34549);
xnor U35199 (N_35199,N_34780,N_34666);
and U35200 (N_35200,N_34919,N_34790);
nor U35201 (N_35201,N_34589,N_34601);
nor U35202 (N_35202,N_34916,N_34590);
xnor U35203 (N_35203,N_34641,N_34519);
or U35204 (N_35204,N_34685,N_34954);
nor U35205 (N_35205,N_34990,N_34953);
nand U35206 (N_35206,N_34785,N_34663);
nor U35207 (N_35207,N_34607,N_34654);
and U35208 (N_35208,N_34664,N_34655);
or U35209 (N_35209,N_34900,N_34640);
xnor U35210 (N_35210,N_34774,N_34560);
nor U35211 (N_35211,N_34925,N_34988);
nor U35212 (N_35212,N_34823,N_34829);
nand U35213 (N_35213,N_34784,N_34991);
xnor U35214 (N_35214,N_34684,N_34618);
and U35215 (N_35215,N_34628,N_34626);
nor U35216 (N_35216,N_34669,N_34695);
or U35217 (N_35217,N_34984,N_34999);
nor U35218 (N_35218,N_34571,N_34520);
nor U35219 (N_35219,N_34703,N_34605);
nand U35220 (N_35220,N_34962,N_34649);
xor U35221 (N_35221,N_34581,N_34952);
xor U35222 (N_35222,N_34644,N_34689);
nand U35223 (N_35223,N_34559,N_34889);
and U35224 (N_35224,N_34904,N_34918);
or U35225 (N_35225,N_34827,N_34895);
nand U35226 (N_35226,N_34854,N_34958);
nor U35227 (N_35227,N_34671,N_34584);
xor U35228 (N_35228,N_34608,N_34778);
and U35229 (N_35229,N_34700,N_34938);
nor U35230 (N_35230,N_34750,N_34727);
and U35231 (N_35231,N_34943,N_34510);
xnor U35232 (N_35232,N_34880,N_34673);
nor U35233 (N_35233,N_34613,N_34600);
or U35234 (N_35234,N_34950,N_34604);
xnor U35235 (N_35235,N_34720,N_34728);
and U35236 (N_35236,N_34864,N_34846);
and U35237 (N_35237,N_34971,N_34583);
or U35238 (N_35238,N_34521,N_34732);
and U35239 (N_35239,N_34801,N_34756);
nor U35240 (N_35240,N_34625,N_34865);
nand U35241 (N_35241,N_34788,N_34528);
nand U35242 (N_35242,N_34587,N_34597);
and U35243 (N_35243,N_34551,N_34745);
nand U35244 (N_35244,N_34997,N_34796);
or U35245 (N_35245,N_34898,N_34873);
or U35246 (N_35246,N_34693,N_34507);
nand U35247 (N_35247,N_34638,N_34556);
or U35248 (N_35248,N_34945,N_34941);
xnor U35249 (N_35249,N_34653,N_34592);
or U35250 (N_35250,N_34777,N_34596);
nor U35251 (N_35251,N_34766,N_34987);
or U35252 (N_35252,N_34806,N_34884);
xor U35253 (N_35253,N_34821,N_34703);
xnor U35254 (N_35254,N_34616,N_34752);
nand U35255 (N_35255,N_34713,N_34995);
or U35256 (N_35256,N_34586,N_34880);
or U35257 (N_35257,N_34700,N_34725);
nand U35258 (N_35258,N_34664,N_34724);
and U35259 (N_35259,N_34889,N_34960);
nand U35260 (N_35260,N_34557,N_34578);
nand U35261 (N_35261,N_34619,N_34662);
nand U35262 (N_35262,N_34874,N_34611);
nand U35263 (N_35263,N_34666,N_34746);
xnor U35264 (N_35264,N_34949,N_34786);
nor U35265 (N_35265,N_34604,N_34620);
and U35266 (N_35266,N_34756,N_34704);
nor U35267 (N_35267,N_34733,N_34742);
xnor U35268 (N_35268,N_34613,N_34932);
or U35269 (N_35269,N_34858,N_34730);
nand U35270 (N_35270,N_34970,N_34554);
nor U35271 (N_35271,N_34893,N_34860);
nand U35272 (N_35272,N_34963,N_34655);
and U35273 (N_35273,N_34973,N_34677);
nand U35274 (N_35274,N_34952,N_34610);
and U35275 (N_35275,N_34930,N_34937);
and U35276 (N_35276,N_34650,N_34543);
nor U35277 (N_35277,N_34667,N_34729);
or U35278 (N_35278,N_34806,N_34649);
nor U35279 (N_35279,N_34657,N_34615);
nand U35280 (N_35280,N_34958,N_34522);
nor U35281 (N_35281,N_34818,N_34876);
or U35282 (N_35282,N_34567,N_34690);
nand U35283 (N_35283,N_34777,N_34574);
xor U35284 (N_35284,N_34808,N_34630);
and U35285 (N_35285,N_34731,N_34533);
xor U35286 (N_35286,N_34879,N_34868);
or U35287 (N_35287,N_34751,N_34888);
nor U35288 (N_35288,N_34609,N_34836);
nand U35289 (N_35289,N_34995,N_34601);
nand U35290 (N_35290,N_34749,N_34835);
nor U35291 (N_35291,N_34785,N_34694);
nor U35292 (N_35292,N_34637,N_34941);
xnor U35293 (N_35293,N_34804,N_34548);
and U35294 (N_35294,N_34842,N_34688);
or U35295 (N_35295,N_34829,N_34882);
nand U35296 (N_35296,N_34739,N_34795);
nand U35297 (N_35297,N_34632,N_34570);
and U35298 (N_35298,N_34764,N_34905);
and U35299 (N_35299,N_34894,N_34927);
nand U35300 (N_35300,N_34962,N_34674);
or U35301 (N_35301,N_34864,N_34777);
nor U35302 (N_35302,N_34768,N_34637);
nand U35303 (N_35303,N_34653,N_34940);
and U35304 (N_35304,N_34562,N_34591);
xor U35305 (N_35305,N_34806,N_34935);
nand U35306 (N_35306,N_34797,N_34770);
nand U35307 (N_35307,N_34890,N_34578);
and U35308 (N_35308,N_34785,N_34754);
xor U35309 (N_35309,N_34888,N_34971);
xor U35310 (N_35310,N_34859,N_34702);
and U35311 (N_35311,N_34846,N_34935);
xor U35312 (N_35312,N_34933,N_34813);
or U35313 (N_35313,N_34542,N_34834);
xnor U35314 (N_35314,N_34624,N_34993);
nor U35315 (N_35315,N_34655,N_34785);
and U35316 (N_35316,N_34591,N_34908);
or U35317 (N_35317,N_34532,N_34891);
nor U35318 (N_35318,N_34557,N_34766);
or U35319 (N_35319,N_34813,N_34792);
nand U35320 (N_35320,N_34857,N_34609);
xnor U35321 (N_35321,N_34813,N_34978);
nand U35322 (N_35322,N_34686,N_34955);
xnor U35323 (N_35323,N_34807,N_34742);
or U35324 (N_35324,N_34544,N_34913);
nand U35325 (N_35325,N_34691,N_34573);
or U35326 (N_35326,N_34664,N_34650);
xnor U35327 (N_35327,N_34714,N_34743);
xor U35328 (N_35328,N_34567,N_34706);
xnor U35329 (N_35329,N_34996,N_34518);
xnor U35330 (N_35330,N_34505,N_34635);
and U35331 (N_35331,N_34533,N_34780);
or U35332 (N_35332,N_34930,N_34919);
nand U35333 (N_35333,N_34874,N_34749);
and U35334 (N_35334,N_34505,N_34839);
xnor U35335 (N_35335,N_34913,N_34698);
nand U35336 (N_35336,N_34718,N_34797);
and U35337 (N_35337,N_34661,N_34971);
xnor U35338 (N_35338,N_34783,N_34810);
and U35339 (N_35339,N_34571,N_34905);
or U35340 (N_35340,N_34701,N_34703);
nand U35341 (N_35341,N_34828,N_34845);
xnor U35342 (N_35342,N_34825,N_34510);
or U35343 (N_35343,N_34769,N_34695);
xor U35344 (N_35344,N_34762,N_34808);
xor U35345 (N_35345,N_34864,N_34861);
nand U35346 (N_35346,N_34841,N_34645);
xor U35347 (N_35347,N_34773,N_34638);
or U35348 (N_35348,N_34700,N_34905);
and U35349 (N_35349,N_34652,N_34832);
nor U35350 (N_35350,N_34860,N_34711);
nor U35351 (N_35351,N_34817,N_34965);
xor U35352 (N_35352,N_34990,N_34505);
or U35353 (N_35353,N_34934,N_34903);
xor U35354 (N_35354,N_34545,N_34858);
and U35355 (N_35355,N_34545,N_34896);
xor U35356 (N_35356,N_34802,N_34772);
and U35357 (N_35357,N_34714,N_34751);
and U35358 (N_35358,N_34785,N_34616);
nand U35359 (N_35359,N_34980,N_34757);
and U35360 (N_35360,N_34752,N_34837);
or U35361 (N_35361,N_34621,N_34595);
or U35362 (N_35362,N_34581,N_34568);
nand U35363 (N_35363,N_34508,N_34830);
nand U35364 (N_35364,N_34629,N_34646);
nor U35365 (N_35365,N_34779,N_34696);
nor U35366 (N_35366,N_34854,N_34516);
or U35367 (N_35367,N_34580,N_34840);
or U35368 (N_35368,N_34772,N_34716);
or U35369 (N_35369,N_34758,N_34614);
nor U35370 (N_35370,N_34968,N_34843);
and U35371 (N_35371,N_34738,N_34819);
xor U35372 (N_35372,N_34965,N_34542);
nand U35373 (N_35373,N_34829,N_34530);
or U35374 (N_35374,N_34691,N_34669);
nor U35375 (N_35375,N_34926,N_34884);
or U35376 (N_35376,N_34962,N_34896);
xor U35377 (N_35377,N_34698,N_34606);
xor U35378 (N_35378,N_34700,N_34598);
or U35379 (N_35379,N_34859,N_34604);
or U35380 (N_35380,N_34936,N_34649);
or U35381 (N_35381,N_34540,N_34588);
or U35382 (N_35382,N_34860,N_34650);
or U35383 (N_35383,N_34783,N_34509);
and U35384 (N_35384,N_34580,N_34505);
nor U35385 (N_35385,N_34770,N_34870);
and U35386 (N_35386,N_34624,N_34867);
nand U35387 (N_35387,N_34602,N_34777);
or U35388 (N_35388,N_34757,N_34746);
xnor U35389 (N_35389,N_34762,N_34635);
nor U35390 (N_35390,N_34811,N_34830);
nor U35391 (N_35391,N_34656,N_34936);
xnor U35392 (N_35392,N_34715,N_34761);
or U35393 (N_35393,N_34861,N_34931);
or U35394 (N_35394,N_34771,N_34584);
nand U35395 (N_35395,N_34652,N_34904);
nor U35396 (N_35396,N_34567,N_34795);
or U35397 (N_35397,N_34868,N_34532);
nor U35398 (N_35398,N_34594,N_34990);
nor U35399 (N_35399,N_34897,N_34703);
xnor U35400 (N_35400,N_34907,N_34650);
and U35401 (N_35401,N_34815,N_34525);
and U35402 (N_35402,N_34595,N_34901);
nand U35403 (N_35403,N_34887,N_34826);
or U35404 (N_35404,N_34503,N_34601);
or U35405 (N_35405,N_34729,N_34831);
nor U35406 (N_35406,N_34777,N_34801);
xor U35407 (N_35407,N_34601,N_34843);
nand U35408 (N_35408,N_34500,N_34501);
and U35409 (N_35409,N_34502,N_34786);
nor U35410 (N_35410,N_34715,N_34899);
nand U35411 (N_35411,N_34886,N_34571);
or U35412 (N_35412,N_34520,N_34976);
nand U35413 (N_35413,N_34836,N_34746);
nand U35414 (N_35414,N_34817,N_34789);
or U35415 (N_35415,N_34699,N_34604);
and U35416 (N_35416,N_34900,N_34971);
nand U35417 (N_35417,N_34644,N_34620);
and U35418 (N_35418,N_34547,N_34618);
or U35419 (N_35419,N_34619,N_34883);
or U35420 (N_35420,N_34744,N_34641);
nor U35421 (N_35421,N_34616,N_34598);
or U35422 (N_35422,N_34852,N_34633);
nor U35423 (N_35423,N_34808,N_34625);
nor U35424 (N_35424,N_34596,N_34722);
or U35425 (N_35425,N_34638,N_34996);
or U35426 (N_35426,N_34636,N_34502);
or U35427 (N_35427,N_34613,N_34815);
nor U35428 (N_35428,N_34614,N_34727);
xnor U35429 (N_35429,N_34645,N_34951);
or U35430 (N_35430,N_34839,N_34707);
or U35431 (N_35431,N_34601,N_34570);
or U35432 (N_35432,N_34742,N_34857);
xor U35433 (N_35433,N_34925,N_34599);
nand U35434 (N_35434,N_34954,N_34599);
and U35435 (N_35435,N_34526,N_34650);
nor U35436 (N_35436,N_34700,N_34662);
nand U35437 (N_35437,N_34865,N_34791);
or U35438 (N_35438,N_34601,N_34764);
or U35439 (N_35439,N_34773,N_34679);
xnor U35440 (N_35440,N_34748,N_34766);
and U35441 (N_35441,N_34669,N_34641);
nand U35442 (N_35442,N_34557,N_34812);
nand U35443 (N_35443,N_34992,N_34711);
or U35444 (N_35444,N_34878,N_34812);
xor U35445 (N_35445,N_34700,N_34748);
or U35446 (N_35446,N_34501,N_34991);
or U35447 (N_35447,N_34536,N_34530);
nor U35448 (N_35448,N_34645,N_34773);
xnor U35449 (N_35449,N_34848,N_34772);
xor U35450 (N_35450,N_34754,N_34579);
xnor U35451 (N_35451,N_34840,N_34600);
nand U35452 (N_35452,N_34808,N_34934);
xnor U35453 (N_35453,N_34560,N_34591);
and U35454 (N_35454,N_34779,N_34506);
nor U35455 (N_35455,N_34515,N_34649);
nor U35456 (N_35456,N_34758,N_34650);
xnor U35457 (N_35457,N_34912,N_34895);
or U35458 (N_35458,N_34805,N_34644);
or U35459 (N_35459,N_34742,N_34877);
nor U35460 (N_35460,N_34887,N_34589);
nor U35461 (N_35461,N_34865,N_34666);
nor U35462 (N_35462,N_34575,N_34586);
xor U35463 (N_35463,N_34514,N_34667);
nor U35464 (N_35464,N_34827,N_34673);
nor U35465 (N_35465,N_34557,N_34610);
xnor U35466 (N_35466,N_34874,N_34521);
and U35467 (N_35467,N_34735,N_34701);
xnor U35468 (N_35468,N_34630,N_34743);
nor U35469 (N_35469,N_34702,N_34990);
nor U35470 (N_35470,N_34503,N_34952);
xnor U35471 (N_35471,N_34778,N_34539);
nor U35472 (N_35472,N_34605,N_34861);
nand U35473 (N_35473,N_34708,N_34922);
nor U35474 (N_35474,N_34763,N_34513);
nor U35475 (N_35475,N_34733,N_34768);
xnor U35476 (N_35476,N_34953,N_34606);
xnor U35477 (N_35477,N_34966,N_34900);
or U35478 (N_35478,N_34614,N_34539);
nand U35479 (N_35479,N_34866,N_34715);
nand U35480 (N_35480,N_34971,N_34930);
nor U35481 (N_35481,N_34563,N_34822);
nor U35482 (N_35482,N_34506,N_34567);
and U35483 (N_35483,N_34567,N_34631);
or U35484 (N_35484,N_34764,N_34746);
or U35485 (N_35485,N_34672,N_34665);
and U35486 (N_35486,N_34865,N_34710);
xnor U35487 (N_35487,N_34777,N_34734);
xnor U35488 (N_35488,N_34544,N_34903);
and U35489 (N_35489,N_34957,N_34680);
or U35490 (N_35490,N_34800,N_34974);
nand U35491 (N_35491,N_34758,N_34922);
and U35492 (N_35492,N_34886,N_34581);
nand U35493 (N_35493,N_34541,N_34958);
xnor U35494 (N_35494,N_34861,N_34842);
nand U35495 (N_35495,N_34562,N_34600);
nand U35496 (N_35496,N_34865,N_34834);
and U35497 (N_35497,N_34912,N_34753);
nor U35498 (N_35498,N_34804,N_34514);
and U35499 (N_35499,N_34744,N_34911);
nor U35500 (N_35500,N_35190,N_35153);
and U35501 (N_35501,N_35428,N_35060);
or U35502 (N_35502,N_35346,N_35298);
or U35503 (N_35503,N_35336,N_35418);
or U35504 (N_35504,N_35465,N_35053);
and U35505 (N_35505,N_35441,N_35163);
xnor U35506 (N_35506,N_35084,N_35301);
and U35507 (N_35507,N_35366,N_35055);
nand U35508 (N_35508,N_35120,N_35310);
xor U35509 (N_35509,N_35064,N_35121);
xnor U35510 (N_35510,N_35089,N_35252);
and U35511 (N_35511,N_35265,N_35221);
nor U35512 (N_35512,N_35041,N_35056);
xor U35513 (N_35513,N_35202,N_35168);
and U35514 (N_35514,N_35050,N_35086);
and U35515 (N_35515,N_35091,N_35297);
nor U35516 (N_35516,N_35494,N_35144);
nand U35517 (N_35517,N_35139,N_35430);
xnor U35518 (N_35518,N_35278,N_35447);
xnor U35519 (N_35519,N_35328,N_35090);
or U35520 (N_35520,N_35167,N_35087);
nand U35521 (N_35521,N_35002,N_35195);
nor U35522 (N_35522,N_35427,N_35098);
nor U35523 (N_35523,N_35484,N_35466);
and U35524 (N_35524,N_35044,N_35017);
and U35525 (N_35525,N_35407,N_35130);
nor U35526 (N_35526,N_35245,N_35377);
xor U35527 (N_35527,N_35429,N_35173);
and U35528 (N_35528,N_35450,N_35077);
or U35529 (N_35529,N_35423,N_35454);
nand U35530 (N_35530,N_35287,N_35443);
and U35531 (N_35531,N_35473,N_35231);
nor U35532 (N_35532,N_35286,N_35256);
xnor U35533 (N_35533,N_35391,N_35141);
nand U35534 (N_35534,N_35078,N_35235);
nand U35535 (N_35535,N_35290,N_35400);
nor U35536 (N_35536,N_35420,N_35203);
nor U35537 (N_35537,N_35421,N_35350);
nor U35538 (N_35538,N_35355,N_35489);
nand U35539 (N_35539,N_35257,N_35174);
nor U35540 (N_35540,N_35157,N_35289);
or U35541 (N_35541,N_35474,N_35412);
and U35542 (N_35542,N_35455,N_35183);
nor U35543 (N_35543,N_35281,N_35342);
and U35544 (N_35544,N_35300,N_35228);
and U35545 (N_35545,N_35057,N_35205);
or U35546 (N_35546,N_35325,N_35048);
xor U35547 (N_35547,N_35131,N_35137);
and U35548 (N_35548,N_35357,N_35248);
xor U35549 (N_35549,N_35011,N_35013);
and U35550 (N_35550,N_35379,N_35415);
xnor U35551 (N_35551,N_35476,N_35007);
nand U35552 (N_35552,N_35499,N_35004);
xnor U35553 (N_35553,N_35399,N_35213);
and U35554 (N_35554,N_35497,N_35171);
nor U35555 (N_35555,N_35065,N_35107);
and U35556 (N_35556,N_35025,N_35304);
xnor U35557 (N_35557,N_35234,N_35179);
xor U35558 (N_35558,N_35291,N_35339);
and U35559 (N_35559,N_35285,N_35193);
nor U35560 (N_35560,N_35424,N_35480);
nor U35561 (N_35561,N_35269,N_35200);
nand U35562 (N_35562,N_35255,N_35394);
or U35563 (N_35563,N_35438,N_35305);
nor U35564 (N_35564,N_35496,N_35416);
nor U35565 (N_35565,N_35270,N_35401);
nor U35566 (N_35566,N_35225,N_35222);
or U35567 (N_35567,N_35068,N_35075);
or U35568 (N_35568,N_35197,N_35276);
nor U35569 (N_35569,N_35442,N_35437);
nand U35570 (N_35570,N_35322,N_35206);
and U35571 (N_35571,N_35329,N_35343);
nand U35572 (N_35572,N_35023,N_35099);
nand U35573 (N_35573,N_35127,N_35467);
or U35574 (N_35574,N_35259,N_35176);
xor U35575 (N_35575,N_35299,N_35295);
or U35576 (N_35576,N_35150,N_35101);
nand U35577 (N_35577,N_35129,N_35324);
and U35578 (N_35578,N_35178,N_35326);
nor U35579 (N_35579,N_35170,N_35122);
nand U35580 (N_35580,N_35364,N_35188);
nor U35581 (N_35581,N_35132,N_35273);
nor U35582 (N_35582,N_35340,N_35277);
nand U35583 (N_35583,N_35334,N_35102);
and U35584 (N_35584,N_35406,N_35397);
xnor U35585 (N_35585,N_35094,N_35146);
nor U35586 (N_35586,N_35124,N_35463);
nand U35587 (N_35587,N_35232,N_35477);
xor U35588 (N_35588,N_35061,N_35363);
nor U35589 (N_35589,N_35279,N_35368);
and U35590 (N_35590,N_35338,N_35396);
nor U35591 (N_35591,N_35076,N_35151);
and U35592 (N_35592,N_35220,N_35172);
nor U35593 (N_35593,N_35229,N_35296);
xnor U35594 (N_35594,N_35373,N_35148);
nand U35595 (N_35595,N_35405,N_35417);
nand U35596 (N_35596,N_35003,N_35387);
nand U35597 (N_35597,N_35106,N_35143);
nand U35598 (N_35598,N_35026,N_35046);
or U35599 (N_35599,N_35319,N_35470);
and U35600 (N_35600,N_35419,N_35062);
nand U35601 (N_35601,N_35408,N_35481);
nor U35602 (N_35602,N_35006,N_35311);
and U35603 (N_35603,N_35010,N_35095);
xnor U35604 (N_35604,N_35258,N_35027);
and U35605 (N_35605,N_35495,N_35035);
nor U35606 (N_35606,N_35116,N_35110);
or U35607 (N_35607,N_35054,N_35199);
xnor U35608 (N_35608,N_35337,N_35436);
or U35609 (N_35609,N_35136,N_35254);
or U35610 (N_35610,N_35092,N_35487);
or U35611 (N_35611,N_35260,N_35492);
nand U35612 (N_35612,N_35113,N_35214);
nand U35613 (N_35613,N_35135,N_35196);
or U35614 (N_35614,N_35280,N_35316);
nor U35615 (N_35615,N_35453,N_35482);
xnor U35616 (N_35616,N_35460,N_35112);
or U35617 (N_35617,N_35445,N_35021);
nand U35618 (N_35618,N_35126,N_35320);
nor U35619 (N_35619,N_35045,N_35294);
xnor U35620 (N_35620,N_35082,N_35052);
or U35621 (N_35621,N_35382,N_35272);
nand U35622 (N_35622,N_35372,N_35493);
and U35623 (N_35623,N_35241,N_35018);
or U35624 (N_35624,N_35093,N_35250);
nor U35625 (N_35625,N_35081,N_35083);
nor U35626 (N_35626,N_35426,N_35347);
nor U35627 (N_35627,N_35029,N_35485);
and U35628 (N_35628,N_35177,N_35165);
nand U35629 (N_35629,N_35016,N_35264);
nand U35630 (N_35630,N_35066,N_35376);
nor U35631 (N_35631,N_35108,N_35244);
and U35632 (N_35632,N_35145,N_35303);
or U35633 (N_35633,N_35464,N_35069);
and U35634 (N_35634,N_35262,N_35348);
xnor U35635 (N_35635,N_35293,N_35240);
and U35636 (N_35636,N_35103,N_35440);
or U35637 (N_35637,N_35491,N_35020);
or U35638 (N_35638,N_35096,N_35133);
nand U35639 (N_35639,N_35111,N_35247);
nand U35640 (N_35640,N_35393,N_35384);
or U35641 (N_35641,N_35446,N_35362);
or U35642 (N_35642,N_35404,N_35209);
nand U35643 (N_35643,N_35433,N_35284);
and U35644 (N_35644,N_35243,N_35201);
nand U35645 (N_35645,N_35351,N_35282);
nand U35646 (N_35646,N_35472,N_35216);
or U35647 (N_35647,N_35331,N_35274);
nor U35648 (N_35648,N_35388,N_35341);
or U35649 (N_35649,N_35034,N_35283);
and U35650 (N_35650,N_35204,N_35097);
nand U35651 (N_35651,N_35344,N_35236);
nand U35652 (N_35652,N_35215,N_35125);
xnor U35653 (N_35653,N_35211,N_35080);
nor U35654 (N_35654,N_35317,N_35439);
nor U35655 (N_35655,N_35224,N_35067);
xor U35656 (N_35656,N_35115,N_35239);
xnor U35657 (N_35657,N_35181,N_35198);
and U35658 (N_35658,N_35488,N_35217);
xnor U35659 (N_35659,N_35128,N_35271);
or U35660 (N_35660,N_35227,N_35070);
nor U35661 (N_35661,N_35457,N_35022);
nand U35662 (N_35662,N_35327,N_35458);
nand U35663 (N_35663,N_35074,N_35088);
nand U35664 (N_35664,N_35267,N_35333);
nor U35665 (N_35665,N_35469,N_35251);
or U35666 (N_35666,N_35313,N_35071);
nor U35667 (N_35667,N_35383,N_35425);
nor U35668 (N_35668,N_35422,N_35330);
and U35669 (N_35669,N_35237,N_35014);
xor U35670 (N_35670,N_35402,N_35370);
xor U35671 (N_35671,N_35123,N_35140);
nand U35672 (N_35672,N_35390,N_35315);
nand U35673 (N_35673,N_35043,N_35085);
and U35674 (N_35674,N_35005,N_35411);
and U35675 (N_35675,N_35036,N_35169);
or U35676 (N_35676,N_35134,N_35185);
and U35677 (N_35677,N_35352,N_35359);
and U35678 (N_35678,N_35307,N_35212);
or U35679 (N_35679,N_35318,N_35154);
and U35680 (N_35680,N_35226,N_35180);
nor U35681 (N_35681,N_35038,N_35142);
xnor U35682 (N_35682,N_35024,N_35354);
nand U35683 (N_35683,N_35490,N_35161);
and U35684 (N_35684,N_35246,N_35238);
nor U35685 (N_35685,N_35186,N_35335);
xnor U35686 (N_35686,N_35403,N_35312);
nor U35687 (N_35687,N_35028,N_35332);
and U35688 (N_35688,N_35449,N_35263);
and U35689 (N_35689,N_35105,N_35037);
or U35690 (N_35690,N_35166,N_35031);
and U35691 (N_35691,N_35192,N_35219);
or U35692 (N_35692,N_35398,N_35308);
nor U35693 (N_35693,N_35147,N_35478);
and U35694 (N_35694,N_35156,N_35009);
xor U35695 (N_35695,N_35249,N_35321);
xor U35696 (N_35696,N_35242,N_35385);
and U35697 (N_35697,N_35375,N_35008);
and U35698 (N_35698,N_35019,N_35162);
and U35699 (N_35699,N_35288,N_35042);
and U35700 (N_35700,N_35435,N_35389);
nor U35701 (N_35701,N_35386,N_35253);
nor U35702 (N_35702,N_35155,N_35040);
nand U35703 (N_35703,N_35033,N_35323);
xor U35704 (N_35704,N_35306,N_35152);
nand U35705 (N_35705,N_35413,N_35345);
and U35706 (N_35706,N_35261,N_35461);
nand U35707 (N_35707,N_35302,N_35479);
and U35708 (N_35708,N_35072,N_35266);
xnor U35709 (N_35709,N_35063,N_35182);
and U35710 (N_35710,N_35149,N_35468);
nand U35711 (N_35711,N_35015,N_35309);
nor U35712 (N_35712,N_35358,N_35432);
and U35713 (N_35713,N_35360,N_35349);
xnor U35714 (N_35714,N_35456,N_35059);
nand U35715 (N_35715,N_35374,N_35118);
and U35716 (N_35716,N_35223,N_35452);
nor U35717 (N_35717,N_35314,N_35100);
nand U35718 (N_35718,N_35268,N_35194);
or U35719 (N_35719,N_35208,N_35459);
xor U35720 (N_35720,N_35000,N_35462);
and U35721 (N_35721,N_35032,N_35371);
nor U35722 (N_35722,N_35109,N_35051);
and U35723 (N_35723,N_35207,N_35104);
nand U35724 (N_35724,N_35365,N_35210);
or U35725 (N_35725,N_35353,N_35369);
nor U35726 (N_35726,N_35119,N_35187);
nand U35727 (N_35727,N_35378,N_35475);
nand U35728 (N_35728,N_35073,N_35039);
nor U35729 (N_35729,N_35292,N_35483);
and U35730 (N_35730,N_35191,N_35395);
xnor U35731 (N_35731,N_35079,N_35159);
or U35732 (N_35732,N_35160,N_35380);
xnor U35733 (N_35733,N_35409,N_35218);
or U35734 (N_35734,N_35030,N_35434);
or U35735 (N_35735,N_35356,N_35392);
or U35736 (N_35736,N_35138,N_35381);
and U35737 (N_35737,N_35012,N_35058);
xnor U35738 (N_35738,N_35001,N_35444);
nor U35739 (N_35739,N_35471,N_35047);
nand U35740 (N_35740,N_35175,N_35448);
or U35741 (N_35741,N_35410,N_35498);
and U35742 (N_35742,N_35414,N_35184);
nor U35743 (N_35743,N_35189,N_35275);
nand U35744 (N_35744,N_35431,N_35158);
nor U35745 (N_35745,N_35117,N_35361);
or U35746 (N_35746,N_35233,N_35049);
nand U35747 (N_35747,N_35230,N_35164);
xor U35748 (N_35748,N_35114,N_35451);
xor U35749 (N_35749,N_35367,N_35486);
or U35750 (N_35750,N_35354,N_35283);
or U35751 (N_35751,N_35044,N_35270);
or U35752 (N_35752,N_35228,N_35206);
xnor U35753 (N_35753,N_35378,N_35237);
nor U35754 (N_35754,N_35454,N_35360);
or U35755 (N_35755,N_35467,N_35112);
nand U35756 (N_35756,N_35295,N_35323);
nor U35757 (N_35757,N_35357,N_35337);
nor U35758 (N_35758,N_35026,N_35348);
and U35759 (N_35759,N_35353,N_35265);
nand U35760 (N_35760,N_35464,N_35403);
or U35761 (N_35761,N_35491,N_35100);
or U35762 (N_35762,N_35283,N_35404);
or U35763 (N_35763,N_35138,N_35199);
nand U35764 (N_35764,N_35076,N_35028);
nor U35765 (N_35765,N_35383,N_35233);
xnor U35766 (N_35766,N_35392,N_35288);
xnor U35767 (N_35767,N_35185,N_35370);
nand U35768 (N_35768,N_35262,N_35435);
and U35769 (N_35769,N_35086,N_35314);
nor U35770 (N_35770,N_35409,N_35296);
nor U35771 (N_35771,N_35454,N_35110);
nand U35772 (N_35772,N_35394,N_35420);
and U35773 (N_35773,N_35013,N_35430);
and U35774 (N_35774,N_35130,N_35412);
and U35775 (N_35775,N_35466,N_35434);
and U35776 (N_35776,N_35189,N_35042);
xnor U35777 (N_35777,N_35277,N_35315);
or U35778 (N_35778,N_35349,N_35457);
or U35779 (N_35779,N_35481,N_35419);
and U35780 (N_35780,N_35003,N_35306);
xor U35781 (N_35781,N_35421,N_35232);
nor U35782 (N_35782,N_35133,N_35139);
or U35783 (N_35783,N_35099,N_35360);
or U35784 (N_35784,N_35248,N_35163);
and U35785 (N_35785,N_35393,N_35451);
or U35786 (N_35786,N_35166,N_35223);
nand U35787 (N_35787,N_35131,N_35173);
or U35788 (N_35788,N_35163,N_35413);
or U35789 (N_35789,N_35385,N_35350);
and U35790 (N_35790,N_35380,N_35456);
or U35791 (N_35791,N_35196,N_35309);
nand U35792 (N_35792,N_35486,N_35170);
nor U35793 (N_35793,N_35380,N_35251);
or U35794 (N_35794,N_35225,N_35053);
nand U35795 (N_35795,N_35285,N_35195);
and U35796 (N_35796,N_35450,N_35363);
and U35797 (N_35797,N_35020,N_35010);
and U35798 (N_35798,N_35113,N_35352);
nor U35799 (N_35799,N_35226,N_35409);
and U35800 (N_35800,N_35309,N_35014);
nand U35801 (N_35801,N_35212,N_35202);
nor U35802 (N_35802,N_35221,N_35394);
xor U35803 (N_35803,N_35496,N_35221);
xor U35804 (N_35804,N_35196,N_35167);
xnor U35805 (N_35805,N_35095,N_35362);
nand U35806 (N_35806,N_35030,N_35092);
and U35807 (N_35807,N_35420,N_35383);
and U35808 (N_35808,N_35168,N_35071);
xor U35809 (N_35809,N_35138,N_35123);
or U35810 (N_35810,N_35330,N_35498);
and U35811 (N_35811,N_35497,N_35206);
and U35812 (N_35812,N_35211,N_35062);
nor U35813 (N_35813,N_35071,N_35459);
xnor U35814 (N_35814,N_35420,N_35364);
and U35815 (N_35815,N_35262,N_35223);
xnor U35816 (N_35816,N_35007,N_35122);
xor U35817 (N_35817,N_35403,N_35441);
nand U35818 (N_35818,N_35377,N_35107);
xor U35819 (N_35819,N_35200,N_35480);
or U35820 (N_35820,N_35322,N_35161);
and U35821 (N_35821,N_35135,N_35433);
nand U35822 (N_35822,N_35054,N_35175);
xor U35823 (N_35823,N_35043,N_35241);
or U35824 (N_35824,N_35063,N_35253);
and U35825 (N_35825,N_35282,N_35200);
nor U35826 (N_35826,N_35132,N_35468);
nand U35827 (N_35827,N_35010,N_35449);
nand U35828 (N_35828,N_35379,N_35145);
nor U35829 (N_35829,N_35343,N_35063);
and U35830 (N_35830,N_35017,N_35126);
xor U35831 (N_35831,N_35094,N_35307);
xnor U35832 (N_35832,N_35435,N_35233);
and U35833 (N_35833,N_35339,N_35454);
or U35834 (N_35834,N_35275,N_35473);
or U35835 (N_35835,N_35390,N_35003);
xor U35836 (N_35836,N_35199,N_35204);
or U35837 (N_35837,N_35049,N_35076);
nand U35838 (N_35838,N_35245,N_35006);
xor U35839 (N_35839,N_35477,N_35069);
xor U35840 (N_35840,N_35370,N_35080);
or U35841 (N_35841,N_35202,N_35276);
or U35842 (N_35842,N_35275,N_35280);
nand U35843 (N_35843,N_35435,N_35207);
xnor U35844 (N_35844,N_35039,N_35199);
nand U35845 (N_35845,N_35351,N_35068);
or U35846 (N_35846,N_35235,N_35400);
nor U35847 (N_35847,N_35155,N_35331);
xor U35848 (N_35848,N_35284,N_35470);
xor U35849 (N_35849,N_35051,N_35321);
and U35850 (N_35850,N_35338,N_35075);
xor U35851 (N_35851,N_35390,N_35142);
nor U35852 (N_35852,N_35096,N_35052);
nand U35853 (N_35853,N_35224,N_35118);
nor U35854 (N_35854,N_35076,N_35356);
xor U35855 (N_35855,N_35332,N_35233);
or U35856 (N_35856,N_35004,N_35337);
nor U35857 (N_35857,N_35130,N_35254);
xnor U35858 (N_35858,N_35375,N_35104);
nand U35859 (N_35859,N_35157,N_35179);
nand U35860 (N_35860,N_35293,N_35393);
and U35861 (N_35861,N_35261,N_35371);
or U35862 (N_35862,N_35201,N_35275);
nand U35863 (N_35863,N_35462,N_35486);
nor U35864 (N_35864,N_35409,N_35095);
xor U35865 (N_35865,N_35479,N_35416);
and U35866 (N_35866,N_35381,N_35426);
xor U35867 (N_35867,N_35283,N_35269);
or U35868 (N_35868,N_35228,N_35342);
and U35869 (N_35869,N_35125,N_35420);
and U35870 (N_35870,N_35025,N_35346);
nor U35871 (N_35871,N_35444,N_35490);
and U35872 (N_35872,N_35445,N_35466);
nand U35873 (N_35873,N_35435,N_35409);
nand U35874 (N_35874,N_35288,N_35026);
nand U35875 (N_35875,N_35012,N_35329);
or U35876 (N_35876,N_35027,N_35491);
nand U35877 (N_35877,N_35453,N_35427);
nand U35878 (N_35878,N_35082,N_35390);
nor U35879 (N_35879,N_35386,N_35261);
xnor U35880 (N_35880,N_35183,N_35490);
nand U35881 (N_35881,N_35029,N_35362);
nand U35882 (N_35882,N_35119,N_35110);
or U35883 (N_35883,N_35333,N_35238);
and U35884 (N_35884,N_35116,N_35196);
or U35885 (N_35885,N_35292,N_35076);
or U35886 (N_35886,N_35348,N_35060);
or U35887 (N_35887,N_35310,N_35116);
or U35888 (N_35888,N_35377,N_35408);
nand U35889 (N_35889,N_35159,N_35063);
xor U35890 (N_35890,N_35484,N_35252);
and U35891 (N_35891,N_35164,N_35358);
or U35892 (N_35892,N_35092,N_35136);
nor U35893 (N_35893,N_35432,N_35200);
or U35894 (N_35894,N_35230,N_35104);
or U35895 (N_35895,N_35452,N_35108);
xnor U35896 (N_35896,N_35103,N_35057);
nor U35897 (N_35897,N_35431,N_35419);
nand U35898 (N_35898,N_35305,N_35434);
nand U35899 (N_35899,N_35263,N_35351);
and U35900 (N_35900,N_35122,N_35455);
and U35901 (N_35901,N_35041,N_35180);
and U35902 (N_35902,N_35240,N_35146);
nand U35903 (N_35903,N_35465,N_35081);
xor U35904 (N_35904,N_35046,N_35429);
and U35905 (N_35905,N_35260,N_35103);
nor U35906 (N_35906,N_35256,N_35146);
or U35907 (N_35907,N_35371,N_35080);
nand U35908 (N_35908,N_35214,N_35478);
xnor U35909 (N_35909,N_35203,N_35370);
nand U35910 (N_35910,N_35426,N_35194);
nor U35911 (N_35911,N_35369,N_35069);
and U35912 (N_35912,N_35479,N_35262);
nor U35913 (N_35913,N_35202,N_35107);
nand U35914 (N_35914,N_35325,N_35340);
or U35915 (N_35915,N_35001,N_35417);
xor U35916 (N_35916,N_35292,N_35254);
xor U35917 (N_35917,N_35450,N_35349);
xnor U35918 (N_35918,N_35278,N_35045);
or U35919 (N_35919,N_35373,N_35164);
nor U35920 (N_35920,N_35027,N_35216);
and U35921 (N_35921,N_35240,N_35301);
nor U35922 (N_35922,N_35154,N_35232);
nand U35923 (N_35923,N_35363,N_35120);
or U35924 (N_35924,N_35269,N_35381);
nand U35925 (N_35925,N_35099,N_35205);
nand U35926 (N_35926,N_35127,N_35100);
or U35927 (N_35927,N_35485,N_35497);
and U35928 (N_35928,N_35169,N_35353);
or U35929 (N_35929,N_35233,N_35498);
nor U35930 (N_35930,N_35409,N_35294);
nand U35931 (N_35931,N_35141,N_35078);
xnor U35932 (N_35932,N_35402,N_35118);
or U35933 (N_35933,N_35077,N_35176);
nor U35934 (N_35934,N_35169,N_35348);
nor U35935 (N_35935,N_35240,N_35349);
nor U35936 (N_35936,N_35116,N_35296);
xnor U35937 (N_35937,N_35351,N_35485);
or U35938 (N_35938,N_35365,N_35096);
nand U35939 (N_35939,N_35440,N_35181);
xnor U35940 (N_35940,N_35271,N_35446);
and U35941 (N_35941,N_35044,N_35350);
or U35942 (N_35942,N_35417,N_35497);
xnor U35943 (N_35943,N_35192,N_35227);
nor U35944 (N_35944,N_35401,N_35316);
and U35945 (N_35945,N_35311,N_35421);
nor U35946 (N_35946,N_35493,N_35377);
xnor U35947 (N_35947,N_35365,N_35138);
xor U35948 (N_35948,N_35245,N_35068);
nor U35949 (N_35949,N_35354,N_35191);
nor U35950 (N_35950,N_35082,N_35135);
and U35951 (N_35951,N_35070,N_35303);
nand U35952 (N_35952,N_35105,N_35343);
nand U35953 (N_35953,N_35340,N_35264);
nor U35954 (N_35954,N_35201,N_35279);
and U35955 (N_35955,N_35363,N_35496);
nor U35956 (N_35956,N_35309,N_35216);
nor U35957 (N_35957,N_35313,N_35237);
nand U35958 (N_35958,N_35287,N_35181);
nor U35959 (N_35959,N_35447,N_35314);
or U35960 (N_35960,N_35351,N_35043);
xnor U35961 (N_35961,N_35088,N_35279);
or U35962 (N_35962,N_35247,N_35431);
nor U35963 (N_35963,N_35384,N_35445);
nor U35964 (N_35964,N_35150,N_35272);
xor U35965 (N_35965,N_35452,N_35135);
nand U35966 (N_35966,N_35290,N_35100);
xnor U35967 (N_35967,N_35439,N_35303);
nor U35968 (N_35968,N_35185,N_35453);
nor U35969 (N_35969,N_35060,N_35359);
and U35970 (N_35970,N_35220,N_35095);
nor U35971 (N_35971,N_35150,N_35355);
xnor U35972 (N_35972,N_35189,N_35141);
nand U35973 (N_35973,N_35456,N_35429);
or U35974 (N_35974,N_35407,N_35155);
or U35975 (N_35975,N_35151,N_35488);
xor U35976 (N_35976,N_35297,N_35419);
nor U35977 (N_35977,N_35021,N_35260);
nor U35978 (N_35978,N_35365,N_35320);
nand U35979 (N_35979,N_35486,N_35299);
or U35980 (N_35980,N_35360,N_35258);
xnor U35981 (N_35981,N_35436,N_35214);
or U35982 (N_35982,N_35354,N_35090);
xnor U35983 (N_35983,N_35002,N_35423);
xnor U35984 (N_35984,N_35445,N_35234);
and U35985 (N_35985,N_35413,N_35357);
nand U35986 (N_35986,N_35009,N_35390);
nor U35987 (N_35987,N_35384,N_35008);
nor U35988 (N_35988,N_35235,N_35241);
and U35989 (N_35989,N_35321,N_35284);
and U35990 (N_35990,N_35123,N_35281);
xnor U35991 (N_35991,N_35355,N_35186);
nand U35992 (N_35992,N_35429,N_35280);
xor U35993 (N_35993,N_35292,N_35072);
xor U35994 (N_35994,N_35244,N_35015);
and U35995 (N_35995,N_35255,N_35121);
and U35996 (N_35996,N_35022,N_35363);
xor U35997 (N_35997,N_35430,N_35148);
xor U35998 (N_35998,N_35451,N_35294);
or U35999 (N_35999,N_35099,N_35286);
xnor U36000 (N_36000,N_35873,N_35555);
xnor U36001 (N_36001,N_35839,N_35789);
xnor U36002 (N_36002,N_35500,N_35558);
nand U36003 (N_36003,N_35728,N_35653);
and U36004 (N_36004,N_35816,N_35949);
nand U36005 (N_36005,N_35512,N_35510);
nor U36006 (N_36006,N_35651,N_35610);
nand U36007 (N_36007,N_35745,N_35544);
nor U36008 (N_36008,N_35724,N_35755);
and U36009 (N_36009,N_35998,N_35842);
or U36010 (N_36010,N_35895,N_35813);
nand U36011 (N_36011,N_35913,N_35975);
xor U36012 (N_36012,N_35658,N_35621);
nand U36013 (N_36013,N_35678,N_35853);
nand U36014 (N_36014,N_35821,N_35573);
nor U36015 (N_36015,N_35561,N_35657);
or U36016 (N_36016,N_35877,N_35707);
and U36017 (N_36017,N_35684,N_35847);
xor U36018 (N_36018,N_35704,N_35675);
or U36019 (N_36019,N_35885,N_35922);
or U36020 (N_36020,N_35982,N_35629);
nor U36021 (N_36021,N_35624,N_35959);
or U36022 (N_36022,N_35669,N_35995);
and U36023 (N_36023,N_35576,N_35862);
xor U36024 (N_36024,N_35616,N_35851);
nand U36025 (N_36025,N_35923,N_35615);
xnor U36026 (N_36026,N_35664,N_35918);
nor U36027 (N_36027,N_35825,N_35860);
and U36028 (N_36028,N_35593,N_35981);
nor U36029 (N_36029,N_35794,N_35973);
nor U36030 (N_36030,N_35891,N_35690);
nand U36031 (N_36031,N_35562,N_35868);
xor U36032 (N_36032,N_35545,N_35606);
and U36033 (N_36033,N_35970,N_35686);
or U36034 (N_36034,N_35683,N_35772);
nor U36035 (N_36035,N_35598,N_35680);
and U36036 (N_36036,N_35647,N_35566);
or U36037 (N_36037,N_35737,N_35726);
nand U36038 (N_36038,N_35894,N_35809);
and U36039 (N_36039,N_35964,N_35687);
nand U36040 (N_36040,N_35521,N_35990);
nand U36041 (N_36041,N_35650,N_35915);
nor U36042 (N_36042,N_35822,N_35713);
nor U36043 (N_36043,N_35831,N_35546);
nand U36044 (N_36044,N_35820,N_35908);
xnor U36045 (N_36045,N_35954,N_35854);
nor U36046 (N_36046,N_35698,N_35681);
nor U36047 (N_36047,N_35695,N_35953);
and U36048 (N_36048,N_35708,N_35799);
and U36049 (N_36049,N_35987,N_35869);
nor U36050 (N_36050,N_35641,N_35957);
and U36051 (N_36051,N_35778,N_35926);
nor U36052 (N_36052,N_35575,N_35955);
and U36053 (N_36053,N_35517,N_35670);
or U36054 (N_36054,N_35829,N_35516);
xor U36055 (N_36055,N_35817,N_35793);
nor U36056 (N_36056,N_35974,N_35927);
and U36057 (N_36057,N_35667,N_35925);
and U36058 (N_36058,N_35983,N_35589);
or U36059 (N_36059,N_35884,N_35557);
nand U36060 (N_36060,N_35688,N_35504);
nor U36061 (N_36061,N_35945,N_35733);
nand U36062 (N_36062,N_35592,N_35832);
nand U36063 (N_36063,N_35689,N_35966);
nand U36064 (N_36064,N_35752,N_35883);
nor U36065 (N_36065,N_35731,N_35694);
nand U36066 (N_36066,N_35897,N_35880);
nor U36067 (N_36067,N_35844,N_35760);
and U36068 (N_36068,N_35819,N_35612);
or U36069 (N_36069,N_35919,N_35547);
nor U36070 (N_36070,N_35900,N_35596);
and U36071 (N_36071,N_35608,N_35586);
or U36072 (N_36072,N_35852,N_35828);
nor U36073 (N_36073,N_35846,N_35725);
nand U36074 (N_36074,N_35734,N_35655);
or U36075 (N_36075,N_35739,N_35985);
and U36076 (N_36076,N_35746,N_35934);
nand U36077 (N_36077,N_35933,N_35812);
xnor U36078 (N_36078,N_35924,N_35888);
and U36079 (N_36079,N_35767,N_35786);
and U36080 (N_36080,N_35766,N_35764);
and U36081 (N_36081,N_35867,N_35743);
or U36082 (N_36082,N_35942,N_35505);
nand U36083 (N_36083,N_35787,N_35602);
nand U36084 (N_36084,N_35859,N_35721);
nand U36085 (N_36085,N_35879,N_35774);
xnor U36086 (N_36086,N_35785,N_35824);
and U36087 (N_36087,N_35588,N_35634);
nand U36088 (N_36088,N_35798,N_35783);
or U36089 (N_36089,N_35501,N_35930);
nand U36090 (N_36090,N_35635,N_35951);
or U36091 (N_36091,N_35511,N_35958);
and U36092 (N_36092,N_35814,N_35674);
or U36093 (N_36093,N_35578,N_35795);
or U36094 (N_36094,N_35685,N_35549);
nand U36095 (N_36095,N_35903,N_35636);
nor U36096 (N_36096,N_35991,N_35528);
xnor U36097 (N_36097,N_35570,N_35600);
xor U36098 (N_36098,N_35758,N_35972);
and U36099 (N_36099,N_35866,N_35940);
nand U36100 (N_36100,N_35630,N_35780);
nand U36101 (N_36101,N_35763,N_35980);
xnor U36102 (N_36102,N_35941,N_35841);
or U36103 (N_36103,N_35776,N_35762);
nand U36104 (N_36104,N_35865,N_35723);
xor U36105 (N_36105,N_35568,N_35863);
and U36106 (N_36106,N_35542,N_35572);
nand U36107 (N_36107,N_35878,N_35673);
nand U36108 (N_36108,N_35911,N_35902);
xnor U36109 (N_36109,N_35692,N_35645);
and U36110 (N_36110,N_35929,N_35916);
nand U36111 (N_36111,N_35585,N_35599);
nand U36112 (N_36112,N_35808,N_35803);
and U36113 (N_36113,N_35648,N_35912);
nand U36114 (N_36114,N_35882,N_35715);
nor U36115 (N_36115,N_35525,N_35909);
nor U36116 (N_36116,N_35997,N_35579);
nand U36117 (N_36117,N_35649,N_35875);
nor U36118 (N_36118,N_35666,N_35782);
xnor U36119 (N_36119,N_35534,N_35693);
or U36120 (N_36120,N_35718,N_35976);
and U36121 (N_36121,N_35805,N_35550);
and U36122 (N_36122,N_35748,N_35871);
nor U36123 (N_36123,N_35671,N_35857);
nor U36124 (N_36124,N_35740,N_35773);
nand U36125 (N_36125,N_35967,N_35849);
nor U36126 (N_36126,N_35896,N_35810);
or U36127 (N_36127,N_35910,N_35656);
or U36128 (N_36128,N_35892,N_35637);
and U36129 (N_36129,N_35503,N_35939);
nor U36130 (N_36130,N_35580,N_35705);
and U36131 (N_36131,N_35899,N_35567);
xor U36132 (N_36132,N_35551,N_35701);
and U36133 (N_36133,N_35646,N_35577);
nand U36134 (N_36134,N_35652,N_35747);
nand U36135 (N_36135,N_35887,N_35548);
xor U36136 (N_36136,N_35617,N_35917);
nand U36137 (N_36137,N_35597,N_35533);
nor U36138 (N_36138,N_35946,N_35947);
and U36139 (N_36139,N_35697,N_35898);
xor U36140 (N_36140,N_35965,N_35827);
nor U36141 (N_36141,N_35770,N_35623);
or U36142 (N_36142,N_35639,N_35727);
nand U36143 (N_36143,N_35559,N_35523);
xnor U36144 (N_36144,N_35749,N_35977);
and U36145 (N_36145,N_35696,N_35881);
xnor U36146 (N_36146,N_35971,N_35514);
or U36147 (N_36147,N_35775,N_35631);
or U36148 (N_36148,N_35565,N_35754);
and U36149 (N_36149,N_35948,N_35906);
nand U36150 (N_36150,N_35907,N_35604);
or U36151 (N_36151,N_35537,N_35700);
nor U36152 (N_36152,N_35717,N_35732);
nand U36153 (N_36153,N_35936,N_35984);
or U36154 (N_36154,N_35571,N_35638);
nand U36155 (N_36155,N_35931,N_35595);
xor U36156 (N_36156,N_35937,N_35796);
nor U36157 (N_36157,N_35761,N_35513);
xnor U36158 (N_36158,N_35642,N_35890);
and U36159 (N_36159,N_35855,N_35823);
and U36160 (N_36160,N_35711,N_35836);
nor U36161 (N_36161,N_35759,N_35797);
nand U36162 (N_36162,N_35515,N_35886);
and U36163 (N_36163,N_35952,N_35611);
nand U36164 (N_36164,N_35583,N_35781);
nand U36165 (N_36165,N_35950,N_35502);
nand U36166 (N_36166,N_35543,N_35730);
or U36167 (N_36167,N_35679,N_35554);
nand U36168 (N_36168,N_35963,N_35607);
nor U36169 (N_36169,N_35712,N_35535);
nand U36170 (N_36170,N_35714,N_35626);
and U36171 (N_36171,N_35800,N_35999);
xnor U36172 (N_36172,N_35552,N_35811);
nand U36173 (N_36173,N_35751,N_35938);
nor U36174 (N_36174,N_35720,N_35806);
and U36175 (N_36175,N_35845,N_35756);
or U36176 (N_36176,N_35969,N_35662);
and U36177 (N_36177,N_35807,N_35591);
or U36178 (N_36178,N_35663,N_35614);
or U36179 (N_36179,N_35703,N_35914);
and U36180 (N_36180,N_35757,N_35790);
xor U36181 (N_36181,N_35861,N_35553);
and U36182 (N_36182,N_35584,N_35876);
nand U36183 (N_36183,N_35628,N_35676);
xnor U36184 (N_36184,N_35590,N_35702);
or U36185 (N_36185,N_35750,N_35709);
xnor U36186 (N_36186,N_35979,N_35856);
xnor U36187 (N_36187,N_35618,N_35654);
and U36188 (N_36188,N_35777,N_35509);
or U36189 (N_36189,N_35527,N_35582);
or U36190 (N_36190,N_35815,N_35706);
nor U36191 (N_36191,N_35769,N_35935);
nand U36192 (N_36192,N_35932,N_35835);
nand U36193 (N_36193,N_35802,N_35870);
nand U36194 (N_36194,N_35519,N_35901);
or U36195 (N_36195,N_35569,N_35874);
or U36196 (N_36196,N_35536,N_35986);
xor U36197 (N_36197,N_35729,N_35644);
nand U36198 (N_36198,N_35771,N_35837);
nor U36199 (N_36199,N_35864,N_35668);
or U36200 (N_36200,N_35665,N_35840);
nand U36201 (N_36201,N_35921,N_35538);
xor U36202 (N_36202,N_35633,N_35742);
nand U36203 (N_36203,N_35904,N_35826);
nand U36204 (N_36204,N_35735,N_35978);
or U36205 (N_36205,N_35858,N_35529);
xor U36206 (N_36206,N_35526,N_35603);
and U36207 (N_36207,N_35830,N_35574);
or U36208 (N_36208,N_35632,N_35928);
xor U36209 (N_36209,N_35539,N_35677);
xnor U36210 (N_36210,N_35556,N_35765);
and U36211 (N_36211,N_35944,N_35850);
nand U36212 (N_36212,N_35992,N_35682);
or U36213 (N_36213,N_35619,N_35779);
nand U36214 (N_36214,N_35993,N_35601);
nor U36215 (N_36215,N_35956,N_35560);
xnor U36216 (N_36216,N_35640,N_35744);
xnor U36217 (N_36217,N_35563,N_35843);
nor U36218 (N_36218,N_35920,N_35962);
nor U36219 (N_36219,N_35620,N_35625);
nand U36220 (N_36220,N_35719,N_35710);
nor U36221 (N_36221,N_35834,N_35672);
or U36222 (N_36222,N_35889,N_35507);
nand U36223 (N_36223,N_35524,N_35988);
or U36224 (N_36224,N_35893,N_35753);
and U36225 (N_36225,N_35660,N_35848);
and U36226 (N_36226,N_35587,N_35613);
nand U36227 (N_36227,N_35508,N_35961);
nor U36228 (N_36228,N_35989,N_35792);
nand U36229 (N_36229,N_35609,N_35661);
nand U36230 (N_36230,N_35520,N_35994);
nand U36231 (N_36231,N_35738,N_35818);
nand U36232 (N_36232,N_35801,N_35872);
or U36233 (N_36233,N_35943,N_35532);
nand U36234 (N_36234,N_35905,N_35564);
or U36235 (N_36235,N_35960,N_35622);
xnor U36236 (N_36236,N_35736,N_35791);
or U36237 (N_36237,N_35659,N_35627);
or U36238 (N_36238,N_35699,N_35643);
nand U36239 (N_36239,N_35605,N_35522);
nor U36240 (N_36240,N_35804,N_35540);
and U36241 (N_36241,N_35716,N_35788);
and U36242 (N_36242,N_35541,N_35691);
and U36243 (N_36243,N_35996,N_35722);
and U36244 (N_36244,N_35518,N_35530);
nand U36245 (N_36245,N_35581,N_35741);
or U36246 (N_36246,N_35768,N_35968);
nand U36247 (N_36247,N_35838,N_35594);
nor U36248 (N_36248,N_35833,N_35531);
xor U36249 (N_36249,N_35506,N_35784);
and U36250 (N_36250,N_35521,N_35563);
nor U36251 (N_36251,N_35649,N_35706);
nand U36252 (N_36252,N_35541,N_35514);
nand U36253 (N_36253,N_35629,N_35734);
nand U36254 (N_36254,N_35509,N_35697);
nor U36255 (N_36255,N_35942,N_35567);
and U36256 (N_36256,N_35908,N_35844);
nand U36257 (N_36257,N_35618,N_35661);
and U36258 (N_36258,N_35776,N_35933);
xnor U36259 (N_36259,N_35901,N_35582);
nand U36260 (N_36260,N_35782,N_35817);
and U36261 (N_36261,N_35882,N_35834);
or U36262 (N_36262,N_35599,N_35644);
and U36263 (N_36263,N_35677,N_35626);
nand U36264 (N_36264,N_35992,N_35613);
nand U36265 (N_36265,N_35510,N_35874);
or U36266 (N_36266,N_35538,N_35752);
or U36267 (N_36267,N_35567,N_35958);
and U36268 (N_36268,N_35727,N_35658);
or U36269 (N_36269,N_35994,N_35628);
nor U36270 (N_36270,N_35730,N_35819);
nor U36271 (N_36271,N_35950,N_35708);
or U36272 (N_36272,N_35891,N_35964);
or U36273 (N_36273,N_35513,N_35809);
xor U36274 (N_36274,N_35860,N_35563);
nand U36275 (N_36275,N_35728,N_35580);
nor U36276 (N_36276,N_35695,N_35734);
and U36277 (N_36277,N_35784,N_35726);
and U36278 (N_36278,N_35913,N_35645);
xnor U36279 (N_36279,N_35606,N_35557);
or U36280 (N_36280,N_35651,N_35807);
or U36281 (N_36281,N_35657,N_35537);
xor U36282 (N_36282,N_35891,N_35954);
and U36283 (N_36283,N_35833,N_35766);
and U36284 (N_36284,N_35553,N_35502);
or U36285 (N_36285,N_35727,N_35513);
and U36286 (N_36286,N_35847,N_35886);
or U36287 (N_36287,N_35506,N_35923);
and U36288 (N_36288,N_35957,N_35879);
nor U36289 (N_36289,N_35543,N_35589);
xnor U36290 (N_36290,N_35858,N_35956);
and U36291 (N_36291,N_35712,N_35627);
and U36292 (N_36292,N_35672,N_35669);
or U36293 (N_36293,N_35554,N_35930);
and U36294 (N_36294,N_35808,N_35592);
nand U36295 (N_36295,N_35655,N_35843);
or U36296 (N_36296,N_35790,N_35853);
xor U36297 (N_36297,N_35780,N_35836);
xor U36298 (N_36298,N_35843,N_35893);
nor U36299 (N_36299,N_35764,N_35904);
nor U36300 (N_36300,N_35957,N_35985);
and U36301 (N_36301,N_35513,N_35892);
or U36302 (N_36302,N_35724,N_35847);
xor U36303 (N_36303,N_35978,N_35503);
xnor U36304 (N_36304,N_35916,N_35535);
xnor U36305 (N_36305,N_35913,N_35861);
or U36306 (N_36306,N_35723,N_35563);
nor U36307 (N_36307,N_35916,N_35562);
nor U36308 (N_36308,N_35978,N_35806);
nand U36309 (N_36309,N_35836,N_35611);
xnor U36310 (N_36310,N_35717,N_35639);
and U36311 (N_36311,N_35765,N_35910);
nor U36312 (N_36312,N_35950,N_35965);
nand U36313 (N_36313,N_35578,N_35840);
and U36314 (N_36314,N_35788,N_35783);
nand U36315 (N_36315,N_35505,N_35925);
nand U36316 (N_36316,N_35862,N_35504);
xor U36317 (N_36317,N_35971,N_35960);
nand U36318 (N_36318,N_35534,N_35602);
nor U36319 (N_36319,N_35967,N_35656);
nand U36320 (N_36320,N_35567,N_35809);
nand U36321 (N_36321,N_35986,N_35647);
xor U36322 (N_36322,N_35735,N_35727);
nor U36323 (N_36323,N_35582,N_35994);
xnor U36324 (N_36324,N_35872,N_35686);
or U36325 (N_36325,N_35629,N_35508);
nor U36326 (N_36326,N_35632,N_35800);
and U36327 (N_36327,N_35791,N_35678);
nor U36328 (N_36328,N_35931,N_35817);
or U36329 (N_36329,N_35824,N_35965);
nand U36330 (N_36330,N_35996,N_35906);
and U36331 (N_36331,N_35559,N_35618);
or U36332 (N_36332,N_35934,N_35972);
xnor U36333 (N_36333,N_35994,N_35552);
nor U36334 (N_36334,N_35981,N_35951);
or U36335 (N_36335,N_35848,N_35670);
xnor U36336 (N_36336,N_35778,N_35969);
or U36337 (N_36337,N_35708,N_35892);
or U36338 (N_36338,N_35704,N_35832);
and U36339 (N_36339,N_35879,N_35842);
and U36340 (N_36340,N_35569,N_35752);
nor U36341 (N_36341,N_35508,N_35884);
and U36342 (N_36342,N_35532,N_35866);
nand U36343 (N_36343,N_35656,N_35840);
nand U36344 (N_36344,N_35866,N_35993);
or U36345 (N_36345,N_35916,N_35993);
and U36346 (N_36346,N_35634,N_35524);
xor U36347 (N_36347,N_35779,N_35754);
or U36348 (N_36348,N_35578,N_35568);
nand U36349 (N_36349,N_35768,N_35870);
or U36350 (N_36350,N_35633,N_35521);
or U36351 (N_36351,N_35687,N_35734);
xnor U36352 (N_36352,N_35803,N_35635);
or U36353 (N_36353,N_35962,N_35627);
and U36354 (N_36354,N_35517,N_35643);
xnor U36355 (N_36355,N_35789,N_35794);
nand U36356 (N_36356,N_35744,N_35980);
nand U36357 (N_36357,N_35555,N_35952);
xnor U36358 (N_36358,N_35631,N_35618);
xor U36359 (N_36359,N_35807,N_35620);
or U36360 (N_36360,N_35722,N_35529);
xnor U36361 (N_36361,N_35918,N_35794);
nand U36362 (N_36362,N_35682,N_35716);
nand U36363 (N_36363,N_35775,N_35960);
nor U36364 (N_36364,N_35759,N_35667);
xor U36365 (N_36365,N_35974,N_35801);
nor U36366 (N_36366,N_35799,N_35620);
and U36367 (N_36367,N_35530,N_35570);
and U36368 (N_36368,N_35669,N_35633);
or U36369 (N_36369,N_35875,N_35591);
nor U36370 (N_36370,N_35722,N_35915);
or U36371 (N_36371,N_35998,N_35728);
or U36372 (N_36372,N_35614,N_35943);
nor U36373 (N_36373,N_35781,N_35680);
or U36374 (N_36374,N_35718,N_35774);
and U36375 (N_36375,N_35994,N_35574);
and U36376 (N_36376,N_35752,N_35637);
and U36377 (N_36377,N_35964,N_35999);
nor U36378 (N_36378,N_35881,N_35711);
nand U36379 (N_36379,N_35939,N_35938);
and U36380 (N_36380,N_35773,N_35702);
xnor U36381 (N_36381,N_35560,N_35984);
or U36382 (N_36382,N_35576,N_35654);
and U36383 (N_36383,N_35571,N_35726);
xor U36384 (N_36384,N_35588,N_35770);
nand U36385 (N_36385,N_35953,N_35878);
xnor U36386 (N_36386,N_35577,N_35710);
or U36387 (N_36387,N_35711,N_35805);
nor U36388 (N_36388,N_35548,N_35929);
nor U36389 (N_36389,N_35502,N_35739);
nand U36390 (N_36390,N_35934,N_35821);
xnor U36391 (N_36391,N_35912,N_35524);
xor U36392 (N_36392,N_35964,N_35875);
or U36393 (N_36393,N_35640,N_35620);
nand U36394 (N_36394,N_35577,N_35766);
nor U36395 (N_36395,N_35735,N_35749);
nand U36396 (N_36396,N_35945,N_35795);
nor U36397 (N_36397,N_35653,N_35610);
nand U36398 (N_36398,N_35595,N_35937);
nand U36399 (N_36399,N_35877,N_35818);
xor U36400 (N_36400,N_35875,N_35807);
or U36401 (N_36401,N_35817,N_35566);
or U36402 (N_36402,N_35629,N_35880);
or U36403 (N_36403,N_35854,N_35740);
nor U36404 (N_36404,N_35738,N_35925);
or U36405 (N_36405,N_35886,N_35754);
xnor U36406 (N_36406,N_35603,N_35501);
nor U36407 (N_36407,N_35829,N_35907);
nand U36408 (N_36408,N_35623,N_35764);
nor U36409 (N_36409,N_35960,N_35801);
or U36410 (N_36410,N_35964,N_35726);
xnor U36411 (N_36411,N_35858,N_35743);
nand U36412 (N_36412,N_35985,N_35692);
and U36413 (N_36413,N_35678,N_35699);
nor U36414 (N_36414,N_35522,N_35937);
and U36415 (N_36415,N_35987,N_35679);
nand U36416 (N_36416,N_35579,N_35729);
nor U36417 (N_36417,N_35697,N_35738);
and U36418 (N_36418,N_35743,N_35878);
or U36419 (N_36419,N_35579,N_35961);
xor U36420 (N_36420,N_35835,N_35842);
nor U36421 (N_36421,N_35877,N_35974);
nor U36422 (N_36422,N_35605,N_35975);
nand U36423 (N_36423,N_35671,N_35757);
nor U36424 (N_36424,N_35746,N_35745);
xnor U36425 (N_36425,N_35962,N_35671);
nand U36426 (N_36426,N_35620,N_35597);
xnor U36427 (N_36427,N_35663,N_35542);
xnor U36428 (N_36428,N_35909,N_35615);
and U36429 (N_36429,N_35748,N_35570);
xnor U36430 (N_36430,N_35808,N_35607);
nand U36431 (N_36431,N_35910,N_35896);
nand U36432 (N_36432,N_35941,N_35750);
and U36433 (N_36433,N_35887,N_35999);
nand U36434 (N_36434,N_35861,N_35942);
and U36435 (N_36435,N_35555,N_35754);
or U36436 (N_36436,N_35768,N_35648);
nand U36437 (N_36437,N_35992,N_35839);
and U36438 (N_36438,N_35632,N_35919);
or U36439 (N_36439,N_35737,N_35591);
nand U36440 (N_36440,N_35620,N_35877);
or U36441 (N_36441,N_35894,N_35974);
nor U36442 (N_36442,N_35657,N_35689);
nor U36443 (N_36443,N_35626,N_35569);
nand U36444 (N_36444,N_35850,N_35940);
xnor U36445 (N_36445,N_35539,N_35788);
and U36446 (N_36446,N_35789,N_35872);
and U36447 (N_36447,N_35987,N_35588);
or U36448 (N_36448,N_35896,N_35543);
and U36449 (N_36449,N_35552,N_35539);
nand U36450 (N_36450,N_35832,N_35632);
nor U36451 (N_36451,N_35670,N_35649);
or U36452 (N_36452,N_35616,N_35693);
or U36453 (N_36453,N_35767,N_35626);
or U36454 (N_36454,N_35970,N_35912);
and U36455 (N_36455,N_35611,N_35795);
xnor U36456 (N_36456,N_35822,N_35796);
nor U36457 (N_36457,N_35839,N_35893);
and U36458 (N_36458,N_35589,N_35931);
nor U36459 (N_36459,N_35855,N_35508);
nor U36460 (N_36460,N_35607,N_35664);
nand U36461 (N_36461,N_35692,N_35731);
nor U36462 (N_36462,N_35602,N_35641);
xor U36463 (N_36463,N_35775,N_35704);
nor U36464 (N_36464,N_35904,N_35884);
nor U36465 (N_36465,N_35622,N_35828);
xor U36466 (N_36466,N_35683,N_35604);
and U36467 (N_36467,N_35959,N_35722);
and U36468 (N_36468,N_35966,N_35568);
nor U36469 (N_36469,N_35972,N_35559);
nor U36470 (N_36470,N_35565,N_35929);
xor U36471 (N_36471,N_35604,N_35712);
nand U36472 (N_36472,N_35584,N_35949);
and U36473 (N_36473,N_35763,N_35707);
or U36474 (N_36474,N_35549,N_35900);
nor U36475 (N_36475,N_35578,N_35883);
and U36476 (N_36476,N_35787,N_35508);
or U36477 (N_36477,N_35844,N_35835);
nand U36478 (N_36478,N_35825,N_35823);
nand U36479 (N_36479,N_35765,N_35906);
nor U36480 (N_36480,N_35795,N_35940);
or U36481 (N_36481,N_35886,N_35769);
nand U36482 (N_36482,N_35785,N_35609);
or U36483 (N_36483,N_35559,N_35510);
or U36484 (N_36484,N_35948,N_35563);
xor U36485 (N_36485,N_35633,N_35771);
nand U36486 (N_36486,N_35655,N_35662);
nand U36487 (N_36487,N_35904,N_35711);
nand U36488 (N_36488,N_35981,N_35870);
and U36489 (N_36489,N_35510,N_35961);
xor U36490 (N_36490,N_35719,N_35913);
nor U36491 (N_36491,N_35553,N_35701);
and U36492 (N_36492,N_35852,N_35732);
nor U36493 (N_36493,N_35959,N_35998);
or U36494 (N_36494,N_35700,N_35996);
nor U36495 (N_36495,N_35518,N_35763);
nor U36496 (N_36496,N_35734,N_35665);
and U36497 (N_36497,N_35810,N_35634);
xnor U36498 (N_36498,N_35711,N_35810);
and U36499 (N_36499,N_35511,N_35663);
xnor U36500 (N_36500,N_36382,N_36434);
or U36501 (N_36501,N_36172,N_36432);
xnor U36502 (N_36502,N_36031,N_36210);
and U36503 (N_36503,N_36343,N_36356);
nor U36504 (N_36504,N_36049,N_36179);
nand U36505 (N_36505,N_36133,N_36467);
or U36506 (N_36506,N_36389,N_36020);
xnor U36507 (N_36507,N_36483,N_36392);
or U36508 (N_36508,N_36140,N_36315);
and U36509 (N_36509,N_36366,N_36066);
and U36510 (N_36510,N_36162,N_36428);
nand U36511 (N_36511,N_36163,N_36156);
xor U36512 (N_36512,N_36150,N_36387);
xnor U36513 (N_36513,N_36285,N_36202);
nand U36514 (N_36514,N_36470,N_36121);
or U36515 (N_36515,N_36201,N_36021);
or U36516 (N_36516,N_36253,N_36209);
and U36517 (N_36517,N_36318,N_36427);
and U36518 (N_36518,N_36265,N_36192);
nor U36519 (N_36519,N_36166,N_36440);
or U36520 (N_36520,N_36301,N_36498);
nor U36521 (N_36521,N_36426,N_36365);
and U36522 (N_36522,N_36293,N_36085);
and U36523 (N_36523,N_36272,N_36204);
nand U36524 (N_36524,N_36221,N_36290);
xor U36525 (N_36525,N_36369,N_36271);
and U36526 (N_36526,N_36231,N_36118);
nor U36527 (N_36527,N_36082,N_36357);
xnor U36528 (N_36528,N_36276,N_36193);
nand U36529 (N_36529,N_36003,N_36386);
and U36530 (N_36530,N_36174,N_36284);
nand U36531 (N_36531,N_36393,N_36263);
and U36532 (N_36532,N_36060,N_36072);
nor U36533 (N_36533,N_36466,N_36308);
or U36534 (N_36534,N_36041,N_36362);
nor U36535 (N_36535,N_36168,N_36354);
nor U36536 (N_36536,N_36149,N_36252);
and U36537 (N_36537,N_36295,N_36421);
or U36538 (N_36538,N_36216,N_36348);
and U36539 (N_36539,N_36171,N_36442);
xor U36540 (N_36540,N_36316,N_36227);
nand U36541 (N_36541,N_36310,N_36262);
nand U36542 (N_36542,N_36092,N_36079);
xor U36543 (N_36543,N_36414,N_36061);
xnor U36544 (N_36544,N_36230,N_36329);
or U36545 (N_36545,N_36496,N_36321);
nor U36546 (N_36546,N_36019,N_36489);
xnor U36547 (N_36547,N_36388,N_36036);
nor U36548 (N_36548,N_36159,N_36096);
xnor U36549 (N_36549,N_36224,N_36142);
xor U36550 (N_36550,N_36304,N_36016);
xor U36551 (N_36551,N_36220,N_36303);
nand U36552 (N_36552,N_36347,N_36103);
and U36553 (N_36553,N_36111,N_36346);
nor U36554 (N_36554,N_36311,N_36146);
or U36555 (N_36555,N_36420,N_36257);
nand U36556 (N_36556,N_36051,N_36007);
xor U36557 (N_36557,N_36360,N_36338);
nand U36558 (N_36558,N_36323,N_36234);
xnor U36559 (N_36559,N_36244,N_36377);
nand U36560 (N_36560,N_36006,N_36232);
nor U36561 (N_36561,N_36353,N_36009);
and U36562 (N_36562,N_36412,N_36050);
nand U36563 (N_36563,N_36010,N_36475);
nor U36564 (N_36564,N_36023,N_36469);
nand U36565 (N_36565,N_36274,N_36270);
nor U36566 (N_36566,N_36494,N_36451);
nor U36567 (N_36567,N_36395,N_36110);
nor U36568 (N_36568,N_36076,N_36029);
or U36569 (N_36569,N_36298,N_36151);
or U36570 (N_36570,N_36409,N_36206);
or U36571 (N_36571,N_36012,N_36098);
nor U36572 (N_36572,N_36207,N_36008);
nor U36573 (N_36573,N_36297,N_36047);
xor U36574 (N_36574,N_36044,N_36190);
nor U36575 (N_36575,N_36139,N_36144);
nand U36576 (N_36576,N_36260,N_36283);
nor U36577 (N_36577,N_36336,N_36312);
and U36578 (N_36578,N_36344,N_36045);
and U36579 (N_36579,N_36198,N_36127);
or U36580 (N_36580,N_36450,N_36130);
nor U36581 (N_36581,N_36436,N_36390);
xor U36582 (N_36582,N_36239,N_36477);
nor U36583 (N_36583,N_36355,N_36246);
and U36584 (N_36584,N_36170,N_36117);
or U36585 (N_36585,N_36183,N_36138);
and U36586 (N_36586,N_36141,N_36238);
nand U36587 (N_36587,N_36471,N_36363);
or U36588 (N_36588,N_36018,N_36487);
or U36589 (N_36589,N_36030,N_36034);
nand U36590 (N_36590,N_36175,N_36408);
nor U36591 (N_36591,N_36435,N_36474);
and U36592 (N_36592,N_36129,N_36225);
or U36593 (N_36593,N_36067,N_36431);
xnor U36594 (N_36594,N_36148,N_36267);
and U36595 (N_36595,N_36430,N_36385);
or U36596 (N_36596,N_36481,N_36482);
nor U36597 (N_36597,N_36119,N_36102);
or U36598 (N_36598,N_36215,N_36070);
nor U36599 (N_36599,N_36203,N_36286);
and U36600 (N_36600,N_36078,N_36397);
nand U36601 (N_36601,N_36399,N_36320);
nand U36602 (N_36602,N_36465,N_36281);
or U36603 (N_36603,N_36074,N_36378);
and U36604 (N_36604,N_36370,N_36058);
nor U36605 (N_36605,N_36017,N_36123);
nor U36606 (N_36606,N_36278,N_36268);
or U36607 (N_36607,N_36473,N_36056);
or U36608 (N_36608,N_36247,N_36306);
or U36609 (N_36609,N_36439,N_36379);
nand U36610 (N_36610,N_36359,N_36188);
nand U36611 (N_36611,N_36187,N_36059);
nor U36612 (N_36612,N_36122,N_36341);
or U36613 (N_36613,N_36404,N_36120);
nand U36614 (N_36614,N_36052,N_36196);
and U36615 (N_36615,N_36277,N_36240);
nand U36616 (N_36616,N_36063,N_36033);
nor U36617 (N_36617,N_36014,N_36124);
and U36618 (N_36618,N_36180,N_36364);
nor U36619 (N_36619,N_36212,N_36037);
xor U36620 (N_36620,N_36128,N_36453);
xor U36621 (N_36621,N_36410,N_36068);
and U36622 (N_36622,N_36419,N_36415);
or U36623 (N_36623,N_36089,N_36333);
or U36624 (N_36624,N_36376,N_36229);
nand U36625 (N_36625,N_36241,N_36391);
nand U36626 (N_36626,N_36396,N_36446);
and U36627 (N_36627,N_36279,N_36444);
and U36628 (N_36628,N_36090,N_36373);
or U36629 (N_36629,N_36147,N_36005);
and U36630 (N_36630,N_36449,N_36400);
nor U36631 (N_36631,N_36112,N_36328);
and U36632 (N_36632,N_36282,N_36189);
nor U36633 (N_36633,N_36332,N_36136);
and U36634 (N_36634,N_36035,N_36491);
xnor U36635 (N_36635,N_36292,N_36228);
nand U36636 (N_36636,N_36406,N_36087);
or U36637 (N_36637,N_36108,N_36027);
xor U36638 (N_36638,N_36307,N_36046);
or U36639 (N_36639,N_36235,N_36083);
nor U36640 (N_36640,N_36157,N_36184);
xnor U36641 (N_36641,N_36104,N_36368);
nor U36642 (N_36642,N_36326,N_36349);
nand U36643 (N_36643,N_36476,N_36381);
nand U36644 (N_36644,N_36043,N_36197);
nand U36645 (N_36645,N_36024,N_36053);
nand U36646 (N_36646,N_36407,N_36275);
and U36647 (N_36647,N_36086,N_36266);
nor U36648 (N_36648,N_36445,N_36114);
or U36649 (N_36649,N_36334,N_36411);
xor U36650 (N_36650,N_36495,N_36222);
nand U36651 (N_36651,N_36422,N_36401);
nand U36652 (N_36652,N_36080,N_36134);
nor U36653 (N_36653,N_36248,N_36398);
or U36654 (N_36654,N_36186,N_36468);
or U36655 (N_36655,N_36459,N_36182);
nor U36656 (N_36656,N_36462,N_36094);
or U36657 (N_36657,N_36004,N_36062);
nor U36658 (N_36658,N_36223,N_36345);
and U36659 (N_36659,N_36001,N_36423);
xnor U36660 (N_36660,N_36109,N_36093);
nor U36661 (N_36661,N_36317,N_36296);
xnor U36662 (N_36662,N_36280,N_36342);
or U36663 (N_36663,N_36013,N_36461);
and U36664 (N_36664,N_36161,N_36164);
and U36665 (N_36665,N_36038,N_36456);
or U36666 (N_36666,N_36490,N_36106);
nand U36667 (N_36667,N_36075,N_36219);
nor U36668 (N_36668,N_36107,N_36250);
xnor U36669 (N_36669,N_36335,N_36361);
and U36670 (N_36670,N_36438,N_36300);
and U36671 (N_36671,N_36177,N_36330);
nand U36672 (N_36672,N_36199,N_36135);
or U36673 (N_36673,N_36394,N_36403);
and U36674 (N_36674,N_36288,N_36371);
and U36675 (N_36675,N_36126,N_36026);
or U36676 (N_36676,N_36145,N_36479);
and U36677 (N_36677,N_36251,N_36226);
nand U36678 (N_36678,N_36113,N_36367);
or U36679 (N_36679,N_36493,N_36057);
nor U36680 (N_36680,N_36443,N_36425);
nor U36681 (N_36681,N_36217,N_36327);
nand U36682 (N_36682,N_36294,N_36042);
nor U36683 (N_36683,N_36088,N_36191);
xor U36684 (N_36684,N_36181,N_36350);
xor U36685 (N_36685,N_36319,N_36302);
nor U36686 (N_36686,N_36492,N_36165);
and U36687 (N_36687,N_36256,N_36314);
and U36688 (N_36688,N_36132,N_36417);
xor U36689 (N_36689,N_36287,N_36313);
and U36690 (N_36690,N_36485,N_36131);
or U36691 (N_36691,N_36173,N_36464);
nand U36692 (N_36692,N_36213,N_36325);
nand U36693 (N_36693,N_36424,N_36324);
and U36694 (N_36694,N_36116,N_36488);
and U36695 (N_36695,N_36243,N_36071);
nor U36696 (N_36696,N_36084,N_36264);
or U36697 (N_36697,N_36039,N_36069);
and U36698 (N_36698,N_36153,N_36454);
nand U36699 (N_36699,N_36155,N_36374);
or U36700 (N_36700,N_36299,N_36486);
nor U36701 (N_36701,N_36405,N_36457);
or U36702 (N_36702,N_36205,N_36384);
and U36703 (N_36703,N_36040,N_36402);
nand U36704 (N_36704,N_36322,N_36291);
or U36705 (N_36705,N_36022,N_36077);
and U36706 (N_36706,N_36011,N_36375);
nor U36707 (N_36707,N_36337,N_36380);
xnor U36708 (N_36708,N_36211,N_36358);
or U36709 (N_36709,N_36169,N_36289);
or U36710 (N_36710,N_36447,N_36158);
nor U36711 (N_36711,N_36480,N_36242);
or U36712 (N_36712,N_36478,N_36340);
nand U36713 (N_36713,N_36383,N_36249);
nor U36714 (N_36714,N_36460,N_36437);
xnor U36715 (N_36715,N_36002,N_36097);
nor U36716 (N_36716,N_36000,N_36055);
xor U36717 (N_36717,N_36015,N_36214);
and U36718 (N_36718,N_36448,N_36305);
or U36719 (N_36719,N_36233,N_36455);
nor U36720 (N_36720,N_36048,N_36458);
nand U36721 (N_36721,N_36125,N_36105);
and U36722 (N_36722,N_36218,N_36054);
nand U36723 (N_36723,N_36237,N_36115);
nor U36724 (N_36724,N_36452,N_36463);
nor U36725 (N_36725,N_36259,N_36154);
nand U36726 (N_36726,N_36269,N_36194);
nand U36727 (N_36727,N_36472,N_36100);
nor U36728 (N_36728,N_36429,N_36160);
xor U36729 (N_36729,N_36413,N_36236);
or U36730 (N_36730,N_36025,N_36261);
nand U36731 (N_36731,N_36273,N_36195);
or U36732 (N_36732,N_36095,N_36143);
or U36733 (N_36733,N_36254,N_36351);
nor U36734 (N_36734,N_36028,N_36200);
and U36735 (N_36735,N_36416,N_36064);
nand U36736 (N_36736,N_36185,N_36339);
or U36737 (N_36737,N_36081,N_36245);
nand U36738 (N_36738,N_36176,N_36101);
and U36739 (N_36739,N_36099,N_36309);
xor U36740 (N_36740,N_36137,N_36441);
or U36741 (N_36741,N_36167,N_36258);
and U36742 (N_36742,N_36208,N_36499);
nor U36743 (N_36743,N_36073,N_36178);
or U36744 (N_36744,N_36418,N_36091);
nand U36745 (N_36745,N_36352,N_36497);
and U36746 (N_36746,N_36484,N_36255);
nor U36747 (N_36747,N_36433,N_36152);
xor U36748 (N_36748,N_36065,N_36372);
nand U36749 (N_36749,N_36032,N_36331);
and U36750 (N_36750,N_36273,N_36052);
or U36751 (N_36751,N_36028,N_36352);
and U36752 (N_36752,N_36113,N_36365);
and U36753 (N_36753,N_36170,N_36383);
xor U36754 (N_36754,N_36366,N_36412);
nand U36755 (N_36755,N_36479,N_36207);
and U36756 (N_36756,N_36346,N_36206);
xor U36757 (N_36757,N_36260,N_36356);
and U36758 (N_36758,N_36169,N_36115);
nor U36759 (N_36759,N_36434,N_36455);
xnor U36760 (N_36760,N_36347,N_36472);
and U36761 (N_36761,N_36338,N_36424);
or U36762 (N_36762,N_36347,N_36096);
xor U36763 (N_36763,N_36093,N_36278);
nand U36764 (N_36764,N_36240,N_36348);
or U36765 (N_36765,N_36325,N_36003);
nand U36766 (N_36766,N_36144,N_36472);
or U36767 (N_36767,N_36291,N_36198);
or U36768 (N_36768,N_36088,N_36220);
and U36769 (N_36769,N_36055,N_36496);
and U36770 (N_36770,N_36105,N_36259);
and U36771 (N_36771,N_36476,N_36146);
or U36772 (N_36772,N_36222,N_36284);
and U36773 (N_36773,N_36398,N_36138);
or U36774 (N_36774,N_36393,N_36465);
nor U36775 (N_36775,N_36155,N_36246);
and U36776 (N_36776,N_36168,N_36317);
and U36777 (N_36777,N_36297,N_36281);
nor U36778 (N_36778,N_36454,N_36412);
nor U36779 (N_36779,N_36171,N_36070);
xnor U36780 (N_36780,N_36482,N_36328);
or U36781 (N_36781,N_36204,N_36260);
nand U36782 (N_36782,N_36370,N_36453);
nor U36783 (N_36783,N_36147,N_36328);
nor U36784 (N_36784,N_36319,N_36005);
nand U36785 (N_36785,N_36253,N_36242);
nand U36786 (N_36786,N_36463,N_36127);
nor U36787 (N_36787,N_36314,N_36327);
or U36788 (N_36788,N_36365,N_36224);
nor U36789 (N_36789,N_36349,N_36455);
nand U36790 (N_36790,N_36153,N_36227);
or U36791 (N_36791,N_36480,N_36324);
nor U36792 (N_36792,N_36259,N_36133);
nand U36793 (N_36793,N_36341,N_36054);
xnor U36794 (N_36794,N_36426,N_36252);
nand U36795 (N_36795,N_36335,N_36430);
nor U36796 (N_36796,N_36436,N_36308);
or U36797 (N_36797,N_36201,N_36450);
nand U36798 (N_36798,N_36349,N_36330);
and U36799 (N_36799,N_36090,N_36216);
and U36800 (N_36800,N_36273,N_36432);
nand U36801 (N_36801,N_36144,N_36043);
nor U36802 (N_36802,N_36259,N_36112);
nand U36803 (N_36803,N_36417,N_36228);
nor U36804 (N_36804,N_36037,N_36416);
nand U36805 (N_36805,N_36146,N_36454);
and U36806 (N_36806,N_36384,N_36217);
or U36807 (N_36807,N_36227,N_36025);
nand U36808 (N_36808,N_36073,N_36309);
xor U36809 (N_36809,N_36415,N_36343);
nand U36810 (N_36810,N_36252,N_36154);
nand U36811 (N_36811,N_36344,N_36176);
nand U36812 (N_36812,N_36241,N_36413);
xor U36813 (N_36813,N_36013,N_36375);
nor U36814 (N_36814,N_36284,N_36306);
xor U36815 (N_36815,N_36081,N_36194);
or U36816 (N_36816,N_36491,N_36146);
nand U36817 (N_36817,N_36157,N_36496);
xnor U36818 (N_36818,N_36028,N_36009);
nor U36819 (N_36819,N_36162,N_36327);
or U36820 (N_36820,N_36111,N_36493);
or U36821 (N_36821,N_36401,N_36366);
nand U36822 (N_36822,N_36119,N_36298);
nor U36823 (N_36823,N_36337,N_36397);
nand U36824 (N_36824,N_36322,N_36440);
nand U36825 (N_36825,N_36165,N_36094);
and U36826 (N_36826,N_36201,N_36234);
nor U36827 (N_36827,N_36136,N_36309);
nor U36828 (N_36828,N_36466,N_36172);
or U36829 (N_36829,N_36320,N_36400);
nand U36830 (N_36830,N_36183,N_36184);
nand U36831 (N_36831,N_36009,N_36018);
nand U36832 (N_36832,N_36432,N_36371);
or U36833 (N_36833,N_36244,N_36128);
nor U36834 (N_36834,N_36432,N_36400);
nor U36835 (N_36835,N_36331,N_36330);
or U36836 (N_36836,N_36388,N_36168);
or U36837 (N_36837,N_36398,N_36105);
or U36838 (N_36838,N_36173,N_36041);
and U36839 (N_36839,N_36057,N_36275);
xnor U36840 (N_36840,N_36301,N_36323);
xnor U36841 (N_36841,N_36387,N_36228);
nor U36842 (N_36842,N_36214,N_36028);
and U36843 (N_36843,N_36293,N_36357);
and U36844 (N_36844,N_36136,N_36140);
nor U36845 (N_36845,N_36379,N_36303);
nor U36846 (N_36846,N_36485,N_36196);
and U36847 (N_36847,N_36072,N_36351);
nand U36848 (N_36848,N_36099,N_36402);
or U36849 (N_36849,N_36325,N_36006);
nor U36850 (N_36850,N_36285,N_36209);
or U36851 (N_36851,N_36213,N_36364);
or U36852 (N_36852,N_36384,N_36066);
and U36853 (N_36853,N_36294,N_36176);
nor U36854 (N_36854,N_36370,N_36338);
or U36855 (N_36855,N_36337,N_36474);
and U36856 (N_36856,N_36480,N_36445);
and U36857 (N_36857,N_36352,N_36366);
nand U36858 (N_36858,N_36341,N_36117);
or U36859 (N_36859,N_36153,N_36066);
nor U36860 (N_36860,N_36133,N_36206);
and U36861 (N_36861,N_36229,N_36173);
xnor U36862 (N_36862,N_36373,N_36324);
nand U36863 (N_36863,N_36006,N_36181);
or U36864 (N_36864,N_36455,N_36227);
xnor U36865 (N_36865,N_36350,N_36125);
xnor U36866 (N_36866,N_36363,N_36423);
and U36867 (N_36867,N_36138,N_36175);
or U36868 (N_36868,N_36106,N_36225);
and U36869 (N_36869,N_36337,N_36187);
or U36870 (N_36870,N_36426,N_36015);
or U36871 (N_36871,N_36251,N_36028);
or U36872 (N_36872,N_36196,N_36376);
or U36873 (N_36873,N_36369,N_36178);
nand U36874 (N_36874,N_36111,N_36451);
and U36875 (N_36875,N_36352,N_36250);
nand U36876 (N_36876,N_36112,N_36160);
and U36877 (N_36877,N_36011,N_36349);
and U36878 (N_36878,N_36216,N_36418);
nand U36879 (N_36879,N_36411,N_36274);
and U36880 (N_36880,N_36194,N_36327);
or U36881 (N_36881,N_36444,N_36053);
nor U36882 (N_36882,N_36014,N_36425);
nand U36883 (N_36883,N_36339,N_36064);
or U36884 (N_36884,N_36480,N_36463);
and U36885 (N_36885,N_36037,N_36482);
xor U36886 (N_36886,N_36429,N_36274);
or U36887 (N_36887,N_36219,N_36054);
nand U36888 (N_36888,N_36447,N_36213);
or U36889 (N_36889,N_36480,N_36201);
and U36890 (N_36890,N_36144,N_36312);
nor U36891 (N_36891,N_36282,N_36225);
xnor U36892 (N_36892,N_36349,N_36428);
nand U36893 (N_36893,N_36272,N_36375);
and U36894 (N_36894,N_36141,N_36140);
or U36895 (N_36895,N_36259,N_36380);
nor U36896 (N_36896,N_36397,N_36237);
nand U36897 (N_36897,N_36135,N_36324);
and U36898 (N_36898,N_36413,N_36045);
and U36899 (N_36899,N_36437,N_36414);
or U36900 (N_36900,N_36141,N_36347);
nand U36901 (N_36901,N_36494,N_36163);
and U36902 (N_36902,N_36488,N_36182);
nand U36903 (N_36903,N_36022,N_36080);
and U36904 (N_36904,N_36114,N_36080);
xnor U36905 (N_36905,N_36191,N_36110);
nand U36906 (N_36906,N_36030,N_36009);
xnor U36907 (N_36907,N_36434,N_36041);
nor U36908 (N_36908,N_36142,N_36305);
and U36909 (N_36909,N_36317,N_36409);
and U36910 (N_36910,N_36390,N_36321);
nand U36911 (N_36911,N_36245,N_36301);
or U36912 (N_36912,N_36203,N_36247);
nand U36913 (N_36913,N_36072,N_36304);
nand U36914 (N_36914,N_36150,N_36421);
and U36915 (N_36915,N_36080,N_36478);
nor U36916 (N_36916,N_36130,N_36175);
or U36917 (N_36917,N_36219,N_36134);
nor U36918 (N_36918,N_36023,N_36107);
nor U36919 (N_36919,N_36340,N_36010);
nand U36920 (N_36920,N_36072,N_36271);
or U36921 (N_36921,N_36073,N_36267);
and U36922 (N_36922,N_36042,N_36030);
xnor U36923 (N_36923,N_36192,N_36021);
nand U36924 (N_36924,N_36427,N_36388);
nor U36925 (N_36925,N_36336,N_36041);
nor U36926 (N_36926,N_36111,N_36099);
xor U36927 (N_36927,N_36473,N_36251);
nand U36928 (N_36928,N_36266,N_36485);
xnor U36929 (N_36929,N_36380,N_36335);
and U36930 (N_36930,N_36299,N_36151);
nand U36931 (N_36931,N_36337,N_36358);
nor U36932 (N_36932,N_36190,N_36399);
or U36933 (N_36933,N_36052,N_36276);
and U36934 (N_36934,N_36253,N_36493);
nand U36935 (N_36935,N_36445,N_36459);
nor U36936 (N_36936,N_36232,N_36428);
and U36937 (N_36937,N_36243,N_36210);
nor U36938 (N_36938,N_36160,N_36153);
and U36939 (N_36939,N_36453,N_36014);
nor U36940 (N_36940,N_36275,N_36319);
nand U36941 (N_36941,N_36071,N_36444);
and U36942 (N_36942,N_36172,N_36341);
or U36943 (N_36943,N_36266,N_36048);
or U36944 (N_36944,N_36246,N_36272);
xnor U36945 (N_36945,N_36199,N_36214);
and U36946 (N_36946,N_36074,N_36008);
nor U36947 (N_36947,N_36379,N_36053);
nand U36948 (N_36948,N_36203,N_36447);
and U36949 (N_36949,N_36194,N_36395);
and U36950 (N_36950,N_36465,N_36163);
nand U36951 (N_36951,N_36319,N_36134);
nor U36952 (N_36952,N_36236,N_36357);
and U36953 (N_36953,N_36371,N_36192);
xor U36954 (N_36954,N_36473,N_36217);
nor U36955 (N_36955,N_36496,N_36258);
or U36956 (N_36956,N_36028,N_36061);
and U36957 (N_36957,N_36370,N_36004);
and U36958 (N_36958,N_36229,N_36260);
nand U36959 (N_36959,N_36423,N_36118);
nand U36960 (N_36960,N_36163,N_36295);
xnor U36961 (N_36961,N_36425,N_36221);
and U36962 (N_36962,N_36413,N_36327);
and U36963 (N_36963,N_36421,N_36027);
xnor U36964 (N_36964,N_36083,N_36106);
and U36965 (N_36965,N_36060,N_36277);
and U36966 (N_36966,N_36326,N_36190);
xnor U36967 (N_36967,N_36209,N_36346);
or U36968 (N_36968,N_36365,N_36229);
and U36969 (N_36969,N_36265,N_36427);
nand U36970 (N_36970,N_36094,N_36124);
xnor U36971 (N_36971,N_36395,N_36370);
xnor U36972 (N_36972,N_36473,N_36033);
and U36973 (N_36973,N_36021,N_36471);
or U36974 (N_36974,N_36223,N_36003);
nor U36975 (N_36975,N_36398,N_36448);
nand U36976 (N_36976,N_36269,N_36499);
and U36977 (N_36977,N_36145,N_36433);
xor U36978 (N_36978,N_36054,N_36165);
nand U36979 (N_36979,N_36434,N_36144);
xor U36980 (N_36980,N_36417,N_36375);
nor U36981 (N_36981,N_36266,N_36329);
nand U36982 (N_36982,N_36212,N_36299);
nand U36983 (N_36983,N_36410,N_36402);
nand U36984 (N_36984,N_36415,N_36389);
and U36985 (N_36985,N_36089,N_36457);
and U36986 (N_36986,N_36329,N_36497);
and U36987 (N_36987,N_36344,N_36249);
nor U36988 (N_36988,N_36143,N_36159);
or U36989 (N_36989,N_36495,N_36205);
or U36990 (N_36990,N_36237,N_36036);
xnor U36991 (N_36991,N_36339,N_36134);
and U36992 (N_36992,N_36354,N_36469);
nand U36993 (N_36993,N_36347,N_36291);
or U36994 (N_36994,N_36254,N_36023);
xnor U36995 (N_36995,N_36435,N_36051);
and U36996 (N_36996,N_36370,N_36331);
xnor U36997 (N_36997,N_36141,N_36300);
or U36998 (N_36998,N_36336,N_36089);
nand U36999 (N_36999,N_36113,N_36423);
xnor U37000 (N_37000,N_36867,N_36687);
and U37001 (N_37001,N_36723,N_36879);
and U37002 (N_37002,N_36794,N_36681);
or U37003 (N_37003,N_36851,N_36539);
or U37004 (N_37004,N_36501,N_36581);
and U37005 (N_37005,N_36657,N_36656);
nor U37006 (N_37006,N_36947,N_36719);
xnor U37007 (N_37007,N_36802,N_36934);
nand U37008 (N_37008,N_36998,N_36958);
and U37009 (N_37009,N_36908,N_36840);
nand U37010 (N_37010,N_36905,N_36798);
and U37011 (N_37011,N_36860,N_36974);
and U37012 (N_37012,N_36627,N_36817);
or U37013 (N_37013,N_36756,N_36510);
xnor U37014 (N_37014,N_36877,N_36910);
nor U37015 (N_37015,N_36674,N_36781);
or U37016 (N_37016,N_36869,N_36861);
or U37017 (N_37017,N_36536,N_36560);
and U37018 (N_37018,N_36976,N_36729);
nand U37019 (N_37019,N_36982,N_36739);
and U37020 (N_37020,N_36952,N_36738);
nand U37021 (N_37021,N_36913,N_36873);
nand U37022 (N_37022,N_36697,N_36830);
or U37023 (N_37023,N_36874,N_36927);
and U37024 (N_37024,N_36928,N_36748);
or U37025 (N_37025,N_36994,N_36638);
or U37026 (N_37026,N_36610,N_36646);
nand U37027 (N_37027,N_36534,N_36871);
nand U37028 (N_37028,N_36891,N_36550);
xor U37029 (N_37029,N_36561,N_36774);
nor U37030 (N_37030,N_36569,N_36537);
and U37031 (N_37031,N_36834,N_36589);
nand U37032 (N_37032,N_36615,N_36829);
and U37033 (N_37033,N_36660,N_36972);
or U37034 (N_37034,N_36975,N_36990);
and U37035 (N_37035,N_36682,N_36895);
or U37036 (N_37036,N_36992,N_36619);
or U37037 (N_37037,N_36700,N_36898);
xnor U37038 (N_37038,N_36606,N_36547);
nand U37039 (N_37039,N_36936,N_36985);
nor U37040 (N_37040,N_36944,N_36528);
or U37041 (N_37041,N_36587,N_36991);
nand U37042 (N_37042,N_36644,N_36800);
and U37043 (N_37043,N_36916,N_36590);
nand U37044 (N_37044,N_36541,N_36698);
nor U37045 (N_37045,N_36814,N_36937);
xnor U37046 (N_37046,N_36556,N_36647);
nor U37047 (N_37047,N_36592,N_36758);
or U37048 (N_37048,N_36866,N_36940);
xnor U37049 (N_37049,N_36710,N_36848);
and U37050 (N_37050,N_36618,N_36977);
xor U37051 (N_37051,N_36742,N_36961);
xor U37052 (N_37052,N_36765,N_36902);
or U37053 (N_37053,N_36813,N_36837);
xnor U37054 (N_37054,N_36938,N_36515);
xor U37055 (N_37055,N_36987,N_36533);
nor U37056 (N_37056,N_36669,N_36683);
nor U37057 (N_37057,N_36875,N_36918);
nor U37058 (N_37058,N_36633,N_36588);
or U37059 (N_37059,N_36704,N_36708);
nand U37060 (N_37060,N_36744,N_36612);
or U37061 (N_37061,N_36816,N_36582);
and U37062 (N_37062,N_36625,N_36551);
or U37063 (N_37063,N_36962,N_36750);
and U37064 (N_37064,N_36822,N_36711);
xor U37065 (N_37065,N_36764,N_36929);
and U37066 (N_37066,N_36931,N_36825);
nor U37067 (N_37067,N_36542,N_36519);
nand U37068 (N_37068,N_36526,N_36824);
and U37069 (N_37069,N_36703,N_36770);
and U37070 (N_37070,N_36686,N_36917);
or U37071 (N_37071,N_36522,N_36695);
nand U37072 (N_37072,N_36752,N_36773);
xnor U37073 (N_37073,N_36768,N_36964);
or U37074 (N_37074,N_36671,N_36844);
nor U37075 (N_37075,N_36585,N_36663);
xnor U37076 (N_37076,N_36573,N_36901);
xnor U37077 (N_37077,N_36602,N_36552);
nor U37078 (N_37078,N_36999,N_36933);
or U37079 (N_37079,N_36523,N_36926);
and U37080 (N_37080,N_36521,N_36838);
xor U37081 (N_37081,N_36562,N_36736);
xnor U37082 (N_37082,N_36776,N_36771);
nand U37083 (N_37083,N_36543,N_36568);
nor U37084 (N_37084,N_36661,N_36850);
nand U37085 (N_37085,N_36572,N_36804);
and U37086 (N_37086,N_36922,N_36823);
or U37087 (N_37087,N_36544,N_36948);
xnor U37088 (N_37088,N_36614,N_36761);
nand U37089 (N_37089,N_36720,N_36833);
xnor U37090 (N_37090,N_36970,N_36932);
xnor U37091 (N_37091,N_36574,N_36580);
or U37092 (N_37092,N_36733,N_36705);
xor U37093 (N_37093,N_36880,N_36864);
xnor U37094 (N_37094,N_36531,N_36503);
xor U37095 (N_37095,N_36524,N_36688);
or U37096 (N_37096,N_36907,N_36951);
nand U37097 (N_37097,N_36731,N_36870);
nand U37098 (N_37098,N_36603,N_36511);
nand U37099 (N_37099,N_36699,N_36535);
or U37100 (N_37100,N_36769,N_36759);
nor U37101 (N_37101,N_36616,N_36514);
or U37102 (N_37102,N_36668,N_36826);
or U37103 (N_37103,N_36712,N_36530);
and U37104 (N_37104,N_36702,N_36617);
or U37105 (N_37105,N_36784,N_36689);
or U37106 (N_37106,N_36753,N_36664);
or U37107 (N_37107,N_36788,N_36591);
xor U37108 (N_37108,N_36713,N_36696);
and U37109 (N_37109,N_36507,N_36676);
or U37110 (N_37110,N_36728,N_36604);
and U37111 (N_37111,N_36717,N_36821);
nand U37112 (N_37112,N_36649,N_36903);
and U37113 (N_37113,N_36807,N_36853);
and U37114 (N_37114,N_36892,N_36596);
nand U37115 (N_37115,N_36808,N_36760);
nand U37116 (N_37116,N_36988,N_36805);
xor U37117 (N_37117,N_36594,N_36797);
or U37118 (N_37118,N_36854,N_36500);
nor U37119 (N_37119,N_36645,N_36899);
and U37120 (N_37120,N_36971,N_36577);
xor U37121 (N_37121,N_36741,N_36734);
nand U37122 (N_37122,N_36783,N_36775);
xnor U37123 (N_37123,N_36896,N_36836);
and U37124 (N_37124,N_36925,N_36652);
nor U37125 (N_37125,N_36843,N_36942);
and U37126 (N_37126,N_36642,N_36984);
xor U37127 (N_37127,N_36754,N_36924);
nand U37128 (N_37128,N_36631,N_36815);
and U37129 (N_37129,N_36540,N_36803);
nor U37130 (N_37130,N_36692,N_36502);
nand U37131 (N_37131,N_36949,N_36780);
or U37132 (N_37132,N_36886,N_36716);
xnor U37133 (N_37133,N_36659,N_36595);
or U37134 (N_37134,N_36986,N_36557);
or U37135 (N_37135,N_36505,N_36620);
xor U37136 (N_37136,N_36890,N_36651);
nor U37137 (N_37137,N_36762,N_36790);
xor U37138 (N_37138,N_36767,N_36513);
nand U37139 (N_37139,N_36506,N_36737);
or U37140 (N_37140,N_36584,N_36641);
nand U37141 (N_37141,N_36923,N_36832);
xor U37142 (N_37142,N_36921,N_36583);
nor U37143 (N_37143,N_36546,N_36565);
nor U37144 (N_37144,N_36956,N_36529);
and U37145 (N_37145,N_36778,N_36946);
or U37146 (N_37146,N_36554,N_36662);
and U37147 (N_37147,N_36629,N_36576);
xor U37148 (N_37148,N_36632,N_36555);
nor U37149 (N_37149,N_36623,N_36959);
xor U37150 (N_37150,N_36912,N_36791);
or U37151 (N_37151,N_36724,N_36978);
nor U37152 (N_37152,N_36607,N_36667);
nor U37153 (N_37153,N_36885,N_36878);
nor U37154 (N_37154,N_36801,N_36613);
and U37155 (N_37155,N_36611,N_36810);
or U37156 (N_37156,N_36520,N_36673);
and U37157 (N_37157,N_36893,N_36745);
nand U37158 (N_37158,N_36709,N_36714);
nor U37159 (N_37159,N_36512,N_36548);
nor U37160 (N_37160,N_36835,N_36706);
and U37161 (N_37161,N_36725,N_36969);
xnor U37162 (N_37162,N_36599,N_36943);
nand U37163 (N_37163,N_36549,N_36578);
nor U37164 (N_37164,N_36564,N_36665);
or U37165 (N_37165,N_36570,N_36693);
or U37166 (N_37166,N_36796,N_36967);
nor U37167 (N_37167,N_36650,N_36532);
nor U37168 (N_37168,N_36635,N_36881);
nor U37169 (N_37169,N_36636,N_36980);
or U37170 (N_37170,N_36571,N_36882);
nor U37171 (N_37171,N_36666,N_36820);
xnor U37172 (N_37172,N_36997,N_36919);
nand U37173 (N_37173,N_36966,N_36605);
or U37174 (N_37174,N_36558,N_36621);
and U37175 (N_37175,N_36701,N_36960);
and U37176 (N_37176,N_36841,N_36852);
nor U37177 (N_37177,N_36965,N_36637);
or U37178 (N_37178,N_36566,N_36670);
nand U37179 (N_37179,N_36849,N_36600);
or U37180 (N_37180,N_36643,N_36579);
or U37181 (N_37181,N_36679,N_36690);
nor U37182 (N_37182,N_36626,N_36954);
nand U37183 (N_37183,N_36538,N_36883);
nand U37184 (N_37184,N_36996,N_36812);
or U37185 (N_37185,N_36939,N_36658);
nor U37186 (N_37186,N_36757,N_36622);
or U37187 (N_37187,N_36887,N_36504);
nor U37188 (N_37188,N_36779,N_36862);
nor U37189 (N_37189,N_36935,N_36653);
xnor U37190 (N_37190,N_36545,N_36787);
or U37191 (N_37191,N_36845,N_36684);
nor U37192 (N_37192,N_36735,N_36598);
nand U37193 (N_37193,N_36597,N_36819);
xor U37194 (N_37194,N_36955,N_36755);
nand U37195 (N_37195,N_36868,N_36553);
and U37196 (N_37196,N_36527,N_36675);
or U37197 (N_37197,N_36718,N_36945);
or U37198 (N_37198,N_36586,N_36648);
nand U37199 (N_37199,N_36909,N_36715);
nor U37200 (N_37200,N_36847,N_36827);
nand U37201 (N_37201,N_36727,N_36973);
nand U37202 (N_37202,N_36884,N_36915);
xnor U37203 (N_37203,N_36792,N_36857);
nand U37204 (N_37204,N_36559,N_36624);
nand U37205 (N_37205,N_36677,N_36567);
xor U37206 (N_37206,N_36842,N_36865);
xnor U37207 (N_37207,N_36672,N_36806);
xor U37208 (N_37208,N_36856,N_36981);
nand U37209 (N_37209,N_36872,N_36811);
nand U37210 (N_37210,N_36889,N_36517);
nand U37211 (N_37211,N_36608,N_36730);
and U37212 (N_37212,N_36930,N_36876);
or U37213 (N_37213,N_36763,N_36721);
nor U37214 (N_37214,N_36751,N_36609);
or U37215 (N_37215,N_36839,N_36846);
xnor U37216 (N_37216,N_36772,N_36601);
nor U37217 (N_37217,N_36563,N_36894);
or U37218 (N_37218,N_36963,N_36749);
nand U37219 (N_37219,N_36640,N_36685);
nor U37220 (N_37220,N_36516,N_36799);
nor U37221 (N_37221,N_36518,N_36979);
nand U37222 (N_37222,N_36680,N_36508);
or U37223 (N_37223,N_36654,N_36818);
nor U37224 (N_37224,N_36707,N_36904);
nand U37225 (N_37225,N_36914,N_36782);
or U37226 (N_37226,N_36509,N_36989);
xor U37227 (N_37227,N_36828,N_36855);
or U37228 (N_37228,N_36777,N_36793);
xor U37229 (N_37229,N_36911,N_36525);
xnor U37230 (N_37230,N_36630,N_36795);
and U37231 (N_37231,N_36993,N_36941);
nand U37232 (N_37232,N_36694,N_36920);
nand U37233 (N_37233,N_36786,N_36888);
or U37234 (N_37234,N_36995,N_36746);
and U37235 (N_37235,N_36906,N_36766);
and U37236 (N_37236,N_36858,N_36950);
nor U37237 (N_37237,N_36831,N_36785);
and U37238 (N_37238,N_36726,N_36628);
xnor U37239 (N_37239,N_36747,N_36634);
or U37240 (N_37240,N_36900,N_36575);
nand U37241 (N_37241,N_36740,N_36863);
nand U37242 (N_37242,N_36789,N_36639);
xor U37243 (N_37243,N_36655,N_36732);
and U37244 (N_37244,N_36953,N_36859);
nor U37245 (N_37245,N_36983,N_36968);
or U37246 (N_37246,N_36593,N_36722);
xnor U37247 (N_37247,N_36897,N_36691);
or U37248 (N_37248,N_36809,N_36957);
xnor U37249 (N_37249,N_36743,N_36678);
or U37250 (N_37250,N_36842,N_36945);
and U37251 (N_37251,N_36882,N_36852);
and U37252 (N_37252,N_36901,N_36730);
nor U37253 (N_37253,N_36799,N_36635);
or U37254 (N_37254,N_36914,N_36951);
or U37255 (N_37255,N_36806,N_36750);
xor U37256 (N_37256,N_36965,N_36996);
and U37257 (N_37257,N_36961,N_36753);
xnor U37258 (N_37258,N_36815,N_36976);
nor U37259 (N_37259,N_36669,N_36795);
or U37260 (N_37260,N_36987,N_36963);
and U37261 (N_37261,N_36697,N_36658);
xor U37262 (N_37262,N_36939,N_36746);
nand U37263 (N_37263,N_36967,N_36768);
and U37264 (N_37264,N_36803,N_36976);
nand U37265 (N_37265,N_36906,N_36908);
and U37266 (N_37266,N_36718,N_36746);
and U37267 (N_37267,N_36505,N_36697);
and U37268 (N_37268,N_36698,N_36660);
nor U37269 (N_37269,N_36635,N_36990);
xor U37270 (N_37270,N_36940,N_36768);
xnor U37271 (N_37271,N_36814,N_36610);
or U37272 (N_37272,N_36779,N_36902);
xor U37273 (N_37273,N_36540,N_36507);
or U37274 (N_37274,N_36840,N_36953);
xnor U37275 (N_37275,N_36805,N_36810);
and U37276 (N_37276,N_36705,N_36671);
and U37277 (N_37277,N_36641,N_36675);
nor U37278 (N_37278,N_36685,N_36652);
nor U37279 (N_37279,N_36518,N_36672);
xnor U37280 (N_37280,N_36535,N_36662);
or U37281 (N_37281,N_36905,N_36821);
nand U37282 (N_37282,N_36766,N_36576);
xor U37283 (N_37283,N_36958,N_36739);
nand U37284 (N_37284,N_36761,N_36611);
and U37285 (N_37285,N_36614,N_36910);
nand U37286 (N_37286,N_36984,N_36559);
xor U37287 (N_37287,N_36675,N_36504);
nand U37288 (N_37288,N_36844,N_36984);
or U37289 (N_37289,N_36530,N_36534);
nor U37290 (N_37290,N_36999,N_36510);
nand U37291 (N_37291,N_36925,N_36671);
nor U37292 (N_37292,N_36592,N_36774);
or U37293 (N_37293,N_36730,N_36551);
nor U37294 (N_37294,N_36532,N_36817);
xnor U37295 (N_37295,N_36565,N_36878);
nand U37296 (N_37296,N_36508,N_36948);
or U37297 (N_37297,N_36557,N_36868);
nand U37298 (N_37298,N_36680,N_36977);
and U37299 (N_37299,N_36642,N_36627);
nor U37300 (N_37300,N_36524,N_36735);
and U37301 (N_37301,N_36731,N_36863);
xor U37302 (N_37302,N_36842,N_36807);
xnor U37303 (N_37303,N_36932,N_36533);
nand U37304 (N_37304,N_36630,N_36584);
nand U37305 (N_37305,N_36807,N_36616);
xor U37306 (N_37306,N_36822,N_36818);
nor U37307 (N_37307,N_36826,N_36638);
or U37308 (N_37308,N_36995,N_36655);
and U37309 (N_37309,N_36878,N_36631);
nand U37310 (N_37310,N_36592,N_36827);
or U37311 (N_37311,N_36728,N_36843);
and U37312 (N_37312,N_36799,N_36890);
xor U37313 (N_37313,N_36529,N_36942);
nor U37314 (N_37314,N_36927,N_36696);
or U37315 (N_37315,N_36699,N_36945);
xnor U37316 (N_37316,N_36866,N_36613);
nor U37317 (N_37317,N_36539,N_36623);
or U37318 (N_37318,N_36597,N_36542);
or U37319 (N_37319,N_36949,N_36690);
nor U37320 (N_37320,N_36967,N_36531);
nand U37321 (N_37321,N_36760,N_36919);
or U37322 (N_37322,N_36676,N_36630);
nand U37323 (N_37323,N_36662,N_36978);
or U37324 (N_37324,N_36694,N_36687);
nor U37325 (N_37325,N_36711,N_36543);
xor U37326 (N_37326,N_36913,N_36690);
xnor U37327 (N_37327,N_36747,N_36578);
xor U37328 (N_37328,N_36777,N_36603);
and U37329 (N_37329,N_36727,N_36929);
and U37330 (N_37330,N_36618,N_36669);
nor U37331 (N_37331,N_36863,N_36531);
xor U37332 (N_37332,N_36772,N_36630);
and U37333 (N_37333,N_36957,N_36516);
xor U37334 (N_37334,N_36577,N_36890);
nand U37335 (N_37335,N_36859,N_36602);
and U37336 (N_37336,N_36512,N_36963);
and U37337 (N_37337,N_36953,N_36930);
xor U37338 (N_37338,N_36653,N_36593);
nand U37339 (N_37339,N_36858,N_36650);
nor U37340 (N_37340,N_36594,N_36616);
nand U37341 (N_37341,N_36810,N_36701);
nor U37342 (N_37342,N_36801,N_36524);
and U37343 (N_37343,N_36671,N_36702);
and U37344 (N_37344,N_36834,N_36962);
xor U37345 (N_37345,N_36585,N_36904);
nor U37346 (N_37346,N_36878,N_36802);
nand U37347 (N_37347,N_36765,N_36556);
nand U37348 (N_37348,N_36882,N_36986);
xor U37349 (N_37349,N_36583,N_36866);
nand U37350 (N_37350,N_36786,N_36904);
and U37351 (N_37351,N_36552,N_36956);
or U37352 (N_37352,N_36765,N_36712);
or U37353 (N_37353,N_36869,N_36718);
xor U37354 (N_37354,N_36836,N_36906);
xor U37355 (N_37355,N_36992,N_36768);
and U37356 (N_37356,N_36815,N_36807);
nand U37357 (N_37357,N_36677,N_36863);
and U37358 (N_37358,N_36745,N_36548);
and U37359 (N_37359,N_36557,N_36890);
nand U37360 (N_37360,N_36744,N_36900);
xnor U37361 (N_37361,N_36746,N_36749);
xor U37362 (N_37362,N_36789,N_36876);
xor U37363 (N_37363,N_36588,N_36761);
or U37364 (N_37364,N_36726,N_36773);
nor U37365 (N_37365,N_36836,N_36939);
nor U37366 (N_37366,N_36517,N_36512);
xor U37367 (N_37367,N_36685,N_36633);
xor U37368 (N_37368,N_36722,N_36956);
nor U37369 (N_37369,N_36810,N_36979);
and U37370 (N_37370,N_36525,N_36910);
and U37371 (N_37371,N_36789,N_36538);
xnor U37372 (N_37372,N_36955,N_36981);
xnor U37373 (N_37373,N_36680,N_36705);
and U37374 (N_37374,N_36804,N_36947);
nor U37375 (N_37375,N_36776,N_36931);
nor U37376 (N_37376,N_36511,N_36696);
nor U37377 (N_37377,N_36998,N_36757);
and U37378 (N_37378,N_36635,N_36538);
and U37379 (N_37379,N_36678,N_36681);
or U37380 (N_37380,N_36959,N_36820);
and U37381 (N_37381,N_36577,N_36628);
and U37382 (N_37382,N_36553,N_36544);
nor U37383 (N_37383,N_36964,N_36547);
xor U37384 (N_37384,N_36680,N_36969);
nor U37385 (N_37385,N_36981,N_36768);
nand U37386 (N_37386,N_36907,N_36754);
or U37387 (N_37387,N_36759,N_36693);
nand U37388 (N_37388,N_36765,N_36975);
nor U37389 (N_37389,N_36945,N_36534);
and U37390 (N_37390,N_36621,N_36868);
nor U37391 (N_37391,N_36507,N_36559);
and U37392 (N_37392,N_36996,N_36691);
nor U37393 (N_37393,N_36865,N_36701);
or U37394 (N_37394,N_36508,N_36885);
xor U37395 (N_37395,N_36603,N_36946);
or U37396 (N_37396,N_36779,N_36514);
or U37397 (N_37397,N_36644,N_36926);
nor U37398 (N_37398,N_36903,N_36555);
or U37399 (N_37399,N_36899,N_36640);
and U37400 (N_37400,N_36650,N_36831);
nor U37401 (N_37401,N_36987,N_36876);
or U37402 (N_37402,N_36905,N_36548);
and U37403 (N_37403,N_36785,N_36586);
nor U37404 (N_37404,N_36778,N_36934);
nor U37405 (N_37405,N_36762,N_36606);
nand U37406 (N_37406,N_36884,N_36516);
nor U37407 (N_37407,N_36639,N_36760);
and U37408 (N_37408,N_36625,N_36942);
or U37409 (N_37409,N_36818,N_36509);
xnor U37410 (N_37410,N_36720,N_36706);
nand U37411 (N_37411,N_36566,N_36695);
nand U37412 (N_37412,N_36793,N_36756);
nand U37413 (N_37413,N_36871,N_36783);
and U37414 (N_37414,N_36983,N_36579);
xnor U37415 (N_37415,N_36794,N_36862);
xnor U37416 (N_37416,N_36770,N_36707);
and U37417 (N_37417,N_36963,N_36603);
or U37418 (N_37418,N_36832,N_36921);
or U37419 (N_37419,N_36600,N_36855);
and U37420 (N_37420,N_36841,N_36539);
xnor U37421 (N_37421,N_36711,N_36776);
nand U37422 (N_37422,N_36795,N_36636);
xor U37423 (N_37423,N_36586,N_36804);
and U37424 (N_37424,N_36927,N_36637);
nand U37425 (N_37425,N_36908,N_36661);
nor U37426 (N_37426,N_36508,N_36994);
xnor U37427 (N_37427,N_36734,N_36781);
nand U37428 (N_37428,N_36808,N_36588);
nor U37429 (N_37429,N_36819,N_36813);
xor U37430 (N_37430,N_36608,N_36569);
and U37431 (N_37431,N_36517,N_36798);
and U37432 (N_37432,N_36988,N_36840);
nand U37433 (N_37433,N_36781,N_36950);
nor U37434 (N_37434,N_36986,N_36899);
xnor U37435 (N_37435,N_36945,N_36652);
and U37436 (N_37436,N_36731,N_36872);
xnor U37437 (N_37437,N_36537,N_36504);
xnor U37438 (N_37438,N_36938,N_36874);
nor U37439 (N_37439,N_36965,N_36998);
nor U37440 (N_37440,N_36511,N_36843);
nor U37441 (N_37441,N_36834,N_36820);
nor U37442 (N_37442,N_36820,N_36897);
nor U37443 (N_37443,N_36989,N_36689);
nand U37444 (N_37444,N_36637,N_36894);
or U37445 (N_37445,N_36880,N_36781);
nor U37446 (N_37446,N_36575,N_36929);
nor U37447 (N_37447,N_36852,N_36903);
or U37448 (N_37448,N_36942,N_36956);
nor U37449 (N_37449,N_36525,N_36763);
or U37450 (N_37450,N_36591,N_36804);
xor U37451 (N_37451,N_36760,N_36579);
and U37452 (N_37452,N_36501,N_36861);
xnor U37453 (N_37453,N_36676,N_36819);
nor U37454 (N_37454,N_36815,N_36709);
xor U37455 (N_37455,N_36978,N_36858);
or U37456 (N_37456,N_36757,N_36755);
and U37457 (N_37457,N_36781,N_36744);
nor U37458 (N_37458,N_36913,N_36969);
nand U37459 (N_37459,N_36547,N_36676);
xnor U37460 (N_37460,N_36651,N_36874);
and U37461 (N_37461,N_36536,N_36558);
nor U37462 (N_37462,N_36648,N_36789);
and U37463 (N_37463,N_36661,N_36790);
or U37464 (N_37464,N_36790,N_36793);
and U37465 (N_37465,N_36634,N_36655);
and U37466 (N_37466,N_36741,N_36630);
or U37467 (N_37467,N_36573,N_36905);
or U37468 (N_37468,N_36851,N_36742);
nor U37469 (N_37469,N_36612,N_36696);
xor U37470 (N_37470,N_36865,N_36661);
nand U37471 (N_37471,N_36819,N_36623);
xor U37472 (N_37472,N_36955,N_36623);
nor U37473 (N_37473,N_36500,N_36678);
xnor U37474 (N_37474,N_36620,N_36766);
nand U37475 (N_37475,N_36939,N_36799);
xor U37476 (N_37476,N_36666,N_36838);
nand U37477 (N_37477,N_36900,N_36587);
nand U37478 (N_37478,N_36923,N_36862);
or U37479 (N_37479,N_36816,N_36702);
and U37480 (N_37480,N_36519,N_36907);
nor U37481 (N_37481,N_36750,N_36901);
xnor U37482 (N_37482,N_36594,N_36962);
and U37483 (N_37483,N_36593,N_36740);
or U37484 (N_37484,N_36647,N_36632);
nor U37485 (N_37485,N_36633,N_36946);
or U37486 (N_37486,N_36905,N_36572);
or U37487 (N_37487,N_36533,N_36556);
and U37488 (N_37488,N_36867,N_36618);
nand U37489 (N_37489,N_36501,N_36616);
nand U37490 (N_37490,N_36850,N_36788);
and U37491 (N_37491,N_36573,N_36781);
or U37492 (N_37492,N_36567,N_36526);
nand U37493 (N_37493,N_36744,N_36546);
nand U37494 (N_37494,N_36717,N_36953);
nor U37495 (N_37495,N_36610,N_36980);
nor U37496 (N_37496,N_36734,N_36539);
and U37497 (N_37497,N_36524,N_36747);
nand U37498 (N_37498,N_36733,N_36894);
nor U37499 (N_37499,N_36673,N_36619);
xnor U37500 (N_37500,N_37447,N_37451);
nand U37501 (N_37501,N_37148,N_37416);
and U37502 (N_37502,N_37220,N_37246);
xor U37503 (N_37503,N_37428,N_37151);
nor U37504 (N_37504,N_37215,N_37064);
nor U37505 (N_37505,N_37418,N_37390);
or U37506 (N_37506,N_37166,N_37441);
and U37507 (N_37507,N_37065,N_37020);
nor U37508 (N_37508,N_37238,N_37352);
xor U37509 (N_37509,N_37409,N_37046);
nor U37510 (N_37510,N_37406,N_37131);
nor U37511 (N_37511,N_37021,N_37184);
and U37512 (N_37512,N_37124,N_37324);
nor U37513 (N_37513,N_37004,N_37030);
and U37514 (N_37514,N_37189,N_37367);
or U37515 (N_37515,N_37171,N_37116);
or U37516 (N_37516,N_37387,N_37008);
xnor U37517 (N_37517,N_37186,N_37015);
nor U37518 (N_37518,N_37107,N_37162);
nand U37519 (N_37519,N_37373,N_37152);
nor U37520 (N_37520,N_37319,N_37351);
or U37521 (N_37521,N_37488,N_37476);
or U37522 (N_37522,N_37233,N_37368);
nor U37523 (N_37523,N_37049,N_37132);
xnor U37524 (N_37524,N_37334,N_37169);
nand U37525 (N_37525,N_37011,N_37484);
xnor U37526 (N_37526,N_37307,N_37435);
and U37527 (N_37527,N_37417,N_37332);
xnor U37528 (N_37528,N_37341,N_37330);
or U37529 (N_37529,N_37028,N_37159);
and U37530 (N_37530,N_37002,N_37266);
nor U37531 (N_37531,N_37265,N_37336);
nand U37532 (N_37532,N_37185,N_37092);
and U37533 (N_37533,N_37261,N_37258);
or U37534 (N_37534,N_37455,N_37420);
nand U37535 (N_37535,N_37267,N_37288);
and U37536 (N_37536,N_37344,N_37232);
or U37537 (N_37537,N_37262,N_37048);
xnor U37538 (N_37538,N_37144,N_37391);
and U37539 (N_37539,N_37143,N_37006);
nand U37540 (N_37540,N_37437,N_37173);
xor U37541 (N_37541,N_37491,N_37123);
nand U37542 (N_37542,N_37063,N_37083);
nand U37543 (N_37543,N_37154,N_37000);
nand U37544 (N_37544,N_37242,N_37157);
nand U37545 (N_37545,N_37062,N_37110);
nor U37546 (N_37546,N_37342,N_37041);
nand U37547 (N_37547,N_37084,N_37458);
and U37548 (N_37548,N_37408,N_37038);
nor U37549 (N_37549,N_37419,N_37378);
nor U37550 (N_37550,N_37308,N_37045);
or U37551 (N_37551,N_37252,N_37466);
nor U37552 (N_37552,N_37198,N_37013);
xor U37553 (N_37553,N_37089,N_37163);
and U37554 (N_37554,N_37073,N_37257);
or U37555 (N_37555,N_37379,N_37053);
nand U37556 (N_37556,N_37389,N_37106);
nand U37557 (N_37557,N_37457,N_37005);
or U37558 (N_37558,N_37462,N_37088);
and U37559 (N_37559,N_37199,N_37472);
nor U37560 (N_37560,N_37290,N_37424);
xnor U37561 (N_37561,N_37253,N_37034);
and U37562 (N_37562,N_37313,N_37235);
nand U37563 (N_37563,N_37204,N_37090);
nor U37564 (N_37564,N_37179,N_37353);
nand U37565 (N_37565,N_37297,N_37432);
and U37566 (N_37566,N_37438,N_37365);
or U37567 (N_37567,N_37100,N_37209);
xor U37568 (N_37568,N_37474,N_37450);
and U37569 (N_37569,N_37206,N_37347);
or U37570 (N_37570,N_37118,N_37029);
xor U37571 (N_37571,N_37079,N_37395);
xnor U37572 (N_37572,N_37058,N_37135);
nor U37573 (N_37573,N_37475,N_37150);
xnor U37574 (N_37574,N_37282,N_37172);
or U37575 (N_37575,N_37480,N_37369);
and U37576 (N_37576,N_37454,N_37385);
nor U37577 (N_37577,N_37093,N_37374);
xnor U37578 (N_37578,N_37111,N_37176);
nand U37579 (N_37579,N_37244,N_37249);
nor U37580 (N_37580,N_37104,N_37156);
nand U37581 (N_37581,N_37141,N_37305);
or U37582 (N_37582,N_37200,N_37444);
and U37583 (N_37583,N_37335,N_37227);
nor U37584 (N_37584,N_37228,N_37280);
and U37585 (N_37585,N_37214,N_37337);
or U37586 (N_37586,N_37033,N_37278);
nand U37587 (N_37587,N_37229,N_37032);
nor U37588 (N_37588,N_37237,N_37178);
nand U37589 (N_37589,N_37328,N_37481);
or U37590 (N_37590,N_37130,N_37255);
nor U37591 (N_37591,N_37294,N_37259);
or U37592 (N_37592,N_37260,N_37477);
and U37593 (N_37593,N_37027,N_37216);
xnor U37594 (N_37594,N_37161,N_37310);
and U37595 (N_37595,N_37165,N_37375);
xor U37596 (N_37596,N_37098,N_37298);
nand U37597 (N_37597,N_37051,N_37007);
nand U37598 (N_37598,N_37471,N_37354);
xnor U37599 (N_37599,N_37421,N_37291);
or U37600 (N_37600,N_37326,N_37001);
and U37601 (N_37601,N_37213,N_37309);
and U37602 (N_37602,N_37443,N_37434);
nand U37603 (N_37603,N_37318,N_37212);
nor U37604 (N_37604,N_37182,N_37348);
nor U37605 (N_37605,N_37277,N_37296);
nand U37606 (N_37606,N_37254,N_37145);
xor U37607 (N_37607,N_37464,N_37263);
nand U37608 (N_37608,N_37251,N_37174);
or U37609 (N_37609,N_37139,N_37483);
xor U37610 (N_37610,N_37393,N_37219);
nand U37611 (N_37611,N_37289,N_37137);
and U37612 (N_37612,N_37453,N_37306);
nand U37613 (N_37613,N_37300,N_37413);
or U37614 (N_37614,N_37105,N_37039);
nor U37615 (N_37615,N_37091,N_37155);
or U37616 (N_37616,N_37205,N_37356);
nand U37617 (N_37617,N_37146,N_37114);
or U37618 (N_37618,N_37180,N_37134);
or U37619 (N_37619,N_37312,N_37066);
and U37620 (N_37620,N_37014,N_37470);
nand U37621 (N_37621,N_37400,N_37321);
and U37622 (N_37622,N_37372,N_37388);
and U37623 (N_37623,N_37115,N_37059);
nor U37624 (N_37624,N_37167,N_37061);
nand U37625 (N_37625,N_37234,N_37175);
or U37626 (N_37626,N_37327,N_37264);
nor U37627 (N_37627,N_37201,N_37412);
xnor U37628 (N_37628,N_37009,N_37362);
and U37629 (N_37629,N_37188,N_37274);
xnor U37630 (N_37630,N_37386,N_37316);
xnor U37631 (N_37631,N_37380,N_37397);
or U37632 (N_37632,N_37446,N_37128);
xnor U37633 (N_37633,N_37448,N_37325);
nand U37634 (N_37634,N_37074,N_37398);
and U37635 (N_37635,N_37010,N_37269);
xor U37636 (N_37636,N_37486,N_37044);
nor U37637 (N_37637,N_37054,N_37355);
nor U37638 (N_37638,N_37121,N_37024);
nor U37639 (N_37639,N_37460,N_37050);
or U37640 (N_37640,N_37493,N_37301);
and U37641 (N_37641,N_37340,N_37097);
xnor U37642 (N_37642,N_37218,N_37404);
and U37643 (N_37643,N_37022,N_37025);
and U37644 (N_37644,N_37425,N_37056);
xnor U37645 (N_37645,N_37320,N_37197);
and U37646 (N_37646,N_37445,N_37381);
or U37647 (N_37647,N_37192,N_37482);
nand U37648 (N_37648,N_37339,N_37170);
and U37649 (N_37649,N_37211,N_37067);
nand U37650 (N_37650,N_37485,N_37075);
or U37651 (N_37651,N_37099,N_37346);
nand U37652 (N_37652,N_37236,N_37060);
xor U37653 (N_37653,N_37479,N_37279);
and U37654 (N_37654,N_37012,N_37338);
or U37655 (N_37655,N_37456,N_37019);
or U37656 (N_37656,N_37031,N_37195);
and U37657 (N_37657,N_37222,N_37323);
nor U37658 (N_37658,N_37069,N_37394);
and U37659 (N_37659,N_37377,N_37042);
and U37660 (N_37660,N_37431,N_37129);
nor U37661 (N_37661,N_37489,N_37411);
or U37662 (N_37662,N_37497,N_37103);
nand U37663 (N_37663,N_37256,N_37343);
nor U37664 (N_37664,N_37401,N_37096);
nor U37665 (N_37665,N_37226,N_37314);
xnor U37666 (N_37666,N_37271,N_37183);
xor U37667 (N_37667,N_37017,N_37383);
nand U37668 (N_37668,N_37125,N_37452);
and U37669 (N_37669,N_37072,N_37361);
and U37670 (N_37670,N_37275,N_37371);
or U37671 (N_37671,N_37345,N_37284);
or U37672 (N_37672,N_37499,N_37126);
nor U37673 (N_37673,N_37360,N_37018);
xnor U37674 (N_37674,N_37392,N_37191);
and U37675 (N_37675,N_37230,N_37317);
xnor U37676 (N_37676,N_37109,N_37293);
nor U37677 (N_37677,N_37463,N_37403);
or U37678 (N_37678,N_37080,N_37496);
and U37679 (N_37679,N_37490,N_37459);
nand U37680 (N_37680,N_37405,N_37133);
or U37681 (N_37681,N_37112,N_37268);
xnor U37682 (N_37682,N_37187,N_37076);
nor U37683 (N_37683,N_37240,N_37026);
nor U37684 (N_37684,N_37329,N_37248);
nand U37685 (N_37685,N_37245,N_37193);
xnor U37686 (N_37686,N_37086,N_37283);
or U37687 (N_37687,N_37467,N_37057);
and U37688 (N_37688,N_37085,N_37429);
xnor U37689 (N_37689,N_37016,N_37158);
nor U37690 (N_37690,N_37160,N_37247);
nand U37691 (N_37691,N_37070,N_37207);
nand U37692 (N_37692,N_37358,N_37492);
nor U37693 (N_37693,N_37402,N_37225);
nand U37694 (N_37694,N_37302,N_37035);
nand U37695 (N_37695,N_37440,N_37498);
or U37696 (N_37696,N_37196,N_37468);
nand U37697 (N_37697,N_37250,N_37023);
nor U37698 (N_37698,N_37040,N_37071);
and U37699 (N_37699,N_37370,N_37427);
nor U37700 (N_37700,N_37315,N_37164);
nor U37701 (N_37701,N_37350,N_37117);
nor U37702 (N_37702,N_37449,N_37068);
or U37703 (N_37703,N_37177,N_37077);
xnor U37704 (N_37704,N_37399,N_37469);
or U37705 (N_37705,N_37494,N_37149);
or U37706 (N_37706,N_37430,N_37078);
and U37707 (N_37707,N_37243,N_37473);
xnor U37708 (N_37708,N_37410,N_37101);
or U37709 (N_37709,N_37120,N_37357);
nand U37710 (N_37710,N_37363,N_37210);
and U37711 (N_37711,N_37407,N_37359);
nor U37712 (N_37712,N_37081,N_37415);
nand U37713 (N_37713,N_37217,N_37426);
nand U37714 (N_37714,N_37303,N_37037);
and U37715 (N_37715,N_37231,N_37181);
nand U37716 (N_37716,N_37433,N_37119);
or U37717 (N_37717,N_37423,N_37366);
nor U37718 (N_37718,N_37190,N_37436);
nand U37719 (N_37719,N_37304,N_37422);
and U37720 (N_37720,N_37292,N_37495);
and U37721 (N_37721,N_37382,N_37333);
nand U37722 (N_37722,N_37287,N_37384);
and U37723 (N_37723,N_37094,N_37036);
nand U37724 (N_37724,N_37276,N_37087);
xor U37725 (N_37725,N_37478,N_37364);
and U37726 (N_37726,N_37043,N_37122);
and U37727 (N_37727,N_37465,N_37322);
nand U37728 (N_37728,N_37272,N_37208);
or U37729 (N_37729,N_37349,N_37052);
and U37730 (N_37730,N_37376,N_37142);
xnor U37731 (N_37731,N_37127,N_37082);
nor U37732 (N_37732,N_37224,N_37203);
and U37733 (N_37733,N_37396,N_37140);
and U37734 (N_37734,N_37108,N_37003);
nand U37735 (N_37735,N_37102,N_37194);
or U37736 (N_37736,N_37273,N_37442);
nor U37737 (N_37737,N_37461,N_37414);
nor U37738 (N_37738,N_37223,N_37487);
xor U37739 (N_37739,N_37299,N_37153);
nor U37740 (N_37740,N_37047,N_37270);
nor U37741 (N_37741,N_37439,N_37055);
nor U37742 (N_37742,N_37138,N_37113);
nor U37743 (N_37743,N_37285,N_37286);
or U37744 (N_37744,N_37202,N_37281);
xor U37745 (N_37745,N_37168,N_37311);
nor U37746 (N_37746,N_37095,N_37295);
nand U37747 (N_37747,N_37241,N_37331);
and U37748 (N_37748,N_37136,N_37221);
nand U37749 (N_37749,N_37147,N_37239);
nor U37750 (N_37750,N_37469,N_37195);
and U37751 (N_37751,N_37424,N_37262);
and U37752 (N_37752,N_37069,N_37216);
or U37753 (N_37753,N_37133,N_37415);
xnor U37754 (N_37754,N_37295,N_37385);
and U37755 (N_37755,N_37026,N_37473);
and U37756 (N_37756,N_37142,N_37109);
or U37757 (N_37757,N_37404,N_37149);
or U37758 (N_37758,N_37182,N_37239);
xor U37759 (N_37759,N_37423,N_37020);
nor U37760 (N_37760,N_37365,N_37472);
xnor U37761 (N_37761,N_37405,N_37180);
or U37762 (N_37762,N_37297,N_37070);
nor U37763 (N_37763,N_37497,N_37259);
xor U37764 (N_37764,N_37051,N_37059);
xor U37765 (N_37765,N_37398,N_37219);
or U37766 (N_37766,N_37050,N_37002);
xor U37767 (N_37767,N_37353,N_37173);
nor U37768 (N_37768,N_37255,N_37126);
nand U37769 (N_37769,N_37064,N_37073);
xor U37770 (N_37770,N_37212,N_37293);
and U37771 (N_37771,N_37367,N_37403);
nor U37772 (N_37772,N_37173,N_37138);
or U37773 (N_37773,N_37061,N_37325);
nand U37774 (N_37774,N_37263,N_37401);
nand U37775 (N_37775,N_37340,N_37332);
nand U37776 (N_37776,N_37024,N_37094);
nand U37777 (N_37777,N_37206,N_37031);
or U37778 (N_37778,N_37324,N_37426);
or U37779 (N_37779,N_37349,N_37191);
or U37780 (N_37780,N_37141,N_37142);
nand U37781 (N_37781,N_37225,N_37051);
nand U37782 (N_37782,N_37420,N_37197);
nand U37783 (N_37783,N_37153,N_37250);
and U37784 (N_37784,N_37458,N_37011);
nor U37785 (N_37785,N_37232,N_37193);
nor U37786 (N_37786,N_37003,N_37379);
nand U37787 (N_37787,N_37042,N_37406);
and U37788 (N_37788,N_37131,N_37253);
nand U37789 (N_37789,N_37388,N_37025);
nand U37790 (N_37790,N_37476,N_37179);
and U37791 (N_37791,N_37322,N_37150);
xor U37792 (N_37792,N_37061,N_37363);
and U37793 (N_37793,N_37133,N_37142);
nand U37794 (N_37794,N_37207,N_37418);
or U37795 (N_37795,N_37103,N_37112);
xor U37796 (N_37796,N_37065,N_37455);
or U37797 (N_37797,N_37166,N_37262);
xnor U37798 (N_37798,N_37336,N_37292);
nor U37799 (N_37799,N_37181,N_37020);
or U37800 (N_37800,N_37212,N_37452);
nand U37801 (N_37801,N_37368,N_37422);
and U37802 (N_37802,N_37304,N_37178);
nor U37803 (N_37803,N_37404,N_37367);
nor U37804 (N_37804,N_37408,N_37134);
or U37805 (N_37805,N_37389,N_37203);
nand U37806 (N_37806,N_37093,N_37430);
xnor U37807 (N_37807,N_37327,N_37365);
nor U37808 (N_37808,N_37481,N_37056);
nand U37809 (N_37809,N_37166,N_37123);
xor U37810 (N_37810,N_37452,N_37170);
nor U37811 (N_37811,N_37365,N_37482);
or U37812 (N_37812,N_37148,N_37139);
xnor U37813 (N_37813,N_37334,N_37298);
and U37814 (N_37814,N_37169,N_37408);
nand U37815 (N_37815,N_37292,N_37268);
nand U37816 (N_37816,N_37364,N_37228);
nor U37817 (N_37817,N_37207,N_37390);
or U37818 (N_37818,N_37166,N_37150);
and U37819 (N_37819,N_37121,N_37398);
or U37820 (N_37820,N_37035,N_37125);
and U37821 (N_37821,N_37345,N_37176);
nand U37822 (N_37822,N_37412,N_37258);
nand U37823 (N_37823,N_37496,N_37036);
or U37824 (N_37824,N_37443,N_37206);
nor U37825 (N_37825,N_37001,N_37071);
and U37826 (N_37826,N_37398,N_37312);
nor U37827 (N_37827,N_37034,N_37385);
or U37828 (N_37828,N_37083,N_37482);
xor U37829 (N_37829,N_37200,N_37230);
or U37830 (N_37830,N_37389,N_37366);
nand U37831 (N_37831,N_37108,N_37061);
nor U37832 (N_37832,N_37366,N_37444);
nor U37833 (N_37833,N_37211,N_37291);
xnor U37834 (N_37834,N_37075,N_37108);
nor U37835 (N_37835,N_37488,N_37070);
and U37836 (N_37836,N_37024,N_37202);
nand U37837 (N_37837,N_37118,N_37202);
xnor U37838 (N_37838,N_37436,N_37483);
nor U37839 (N_37839,N_37067,N_37089);
nand U37840 (N_37840,N_37326,N_37412);
or U37841 (N_37841,N_37131,N_37092);
and U37842 (N_37842,N_37378,N_37090);
nand U37843 (N_37843,N_37069,N_37344);
and U37844 (N_37844,N_37489,N_37327);
xor U37845 (N_37845,N_37426,N_37369);
nor U37846 (N_37846,N_37067,N_37393);
and U37847 (N_37847,N_37223,N_37198);
xor U37848 (N_37848,N_37458,N_37002);
or U37849 (N_37849,N_37480,N_37302);
and U37850 (N_37850,N_37450,N_37331);
nor U37851 (N_37851,N_37431,N_37217);
or U37852 (N_37852,N_37489,N_37086);
or U37853 (N_37853,N_37267,N_37156);
and U37854 (N_37854,N_37112,N_37435);
nand U37855 (N_37855,N_37002,N_37275);
or U37856 (N_37856,N_37247,N_37382);
and U37857 (N_37857,N_37090,N_37255);
and U37858 (N_37858,N_37006,N_37285);
nand U37859 (N_37859,N_37181,N_37057);
nor U37860 (N_37860,N_37015,N_37463);
xor U37861 (N_37861,N_37097,N_37343);
and U37862 (N_37862,N_37369,N_37259);
and U37863 (N_37863,N_37497,N_37349);
nand U37864 (N_37864,N_37116,N_37179);
or U37865 (N_37865,N_37467,N_37101);
nor U37866 (N_37866,N_37252,N_37268);
xor U37867 (N_37867,N_37193,N_37285);
or U37868 (N_37868,N_37020,N_37252);
and U37869 (N_37869,N_37318,N_37088);
and U37870 (N_37870,N_37198,N_37450);
nor U37871 (N_37871,N_37098,N_37345);
nand U37872 (N_37872,N_37006,N_37222);
xnor U37873 (N_37873,N_37366,N_37112);
and U37874 (N_37874,N_37137,N_37485);
nand U37875 (N_37875,N_37120,N_37291);
and U37876 (N_37876,N_37199,N_37337);
nand U37877 (N_37877,N_37081,N_37357);
xor U37878 (N_37878,N_37233,N_37306);
xor U37879 (N_37879,N_37381,N_37172);
and U37880 (N_37880,N_37113,N_37297);
nor U37881 (N_37881,N_37066,N_37262);
and U37882 (N_37882,N_37275,N_37014);
and U37883 (N_37883,N_37417,N_37103);
xor U37884 (N_37884,N_37144,N_37115);
xnor U37885 (N_37885,N_37308,N_37157);
nand U37886 (N_37886,N_37493,N_37022);
nand U37887 (N_37887,N_37053,N_37122);
or U37888 (N_37888,N_37187,N_37148);
nor U37889 (N_37889,N_37033,N_37313);
nor U37890 (N_37890,N_37052,N_37497);
nand U37891 (N_37891,N_37294,N_37129);
nand U37892 (N_37892,N_37441,N_37342);
or U37893 (N_37893,N_37349,N_37353);
or U37894 (N_37894,N_37037,N_37085);
nand U37895 (N_37895,N_37345,N_37332);
xor U37896 (N_37896,N_37482,N_37490);
xnor U37897 (N_37897,N_37029,N_37181);
nor U37898 (N_37898,N_37053,N_37200);
and U37899 (N_37899,N_37200,N_37428);
or U37900 (N_37900,N_37198,N_37480);
nor U37901 (N_37901,N_37491,N_37245);
and U37902 (N_37902,N_37174,N_37318);
xor U37903 (N_37903,N_37006,N_37027);
nand U37904 (N_37904,N_37322,N_37388);
nand U37905 (N_37905,N_37087,N_37484);
nand U37906 (N_37906,N_37163,N_37347);
or U37907 (N_37907,N_37017,N_37305);
or U37908 (N_37908,N_37216,N_37361);
or U37909 (N_37909,N_37443,N_37024);
nor U37910 (N_37910,N_37250,N_37382);
nor U37911 (N_37911,N_37227,N_37083);
nor U37912 (N_37912,N_37032,N_37471);
xor U37913 (N_37913,N_37367,N_37323);
and U37914 (N_37914,N_37226,N_37049);
nor U37915 (N_37915,N_37236,N_37030);
nand U37916 (N_37916,N_37133,N_37223);
nor U37917 (N_37917,N_37497,N_37198);
xor U37918 (N_37918,N_37307,N_37493);
xor U37919 (N_37919,N_37072,N_37005);
nor U37920 (N_37920,N_37283,N_37152);
xnor U37921 (N_37921,N_37408,N_37439);
nor U37922 (N_37922,N_37298,N_37308);
nor U37923 (N_37923,N_37217,N_37081);
or U37924 (N_37924,N_37406,N_37454);
xnor U37925 (N_37925,N_37047,N_37318);
nor U37926 (N_37926,N_37202,N_37043);
nand U37927 (N_37927,N_37021,N_37009);
and U37928 (N_37928,N_37116,N_37322);
nand U37929 (N_37929,N_37208,N_37047);
nor U37930 (N_37930,N_37013,N_37155);
nor U37931 (N_37931,N_37491,N_37044);
nand U37932 (N_37932,N_37134,N_37173);
nor U37933 (N_37933,N_37402,N_37101);
nand U37934 (N_37934,N_37237,N_37134);
nand U37935 (N_37935,N_37312,N_37107);
nor U37936 (N_37936,N_37169,N_37397);
xor U37937 (N_37937,N_37137,N_37346);
nand U37938 (N_37938,N_37408,N_37205);
nor U37939 (N_37939,N_37032,N_37186);
and U37940 (N_37940,N_37142,N_37113);
or U37941 (N_37941,N_37159,N_37123);
and U37942 (N_37942,N_37152,N_37199);
or U37943 (N_37943,N_37120,N_37448);
nand U37944 (N_37944,N_37297,N_37279);
or U37945 (N_37945,N_37400,N_37235);
nor U37946 (N_37946,N_37301,N_37351);
nand U37947 (N_37947,N_37496,N_37129);
xnor U37948 (N_37948,N_37388,N_37391);
nor U37949 (N_37949,N_37388,N_37163);
nor U37950 (N_37950,N_37421,N_37458);
and U37951 (N_37951,N_37225,N_37329);
nor U37952 (N_37952,N_37448,N_37206);
nand U37953 (N_37953,N_37146,N_37419);
nand U37954 (N_37954,N_37130,N_37413);
and U37955 (N_37955,N_37297,N_37189);
xnor U37956 (N_37956,N_37025,N_37061);
nand U37957 (N_37957,N_37293,N_37011);
xnor U37958 (N_37958,N_37152,N_37051);
xnor U37959 (N_37959,N_37424,N_37476);
xor U37960 (N_37960,N_37486,N_37488);
or U37961 (N_37961,N_37061,N_37292);
or U37962 (N_37962,N_37270,N_37362);
and U37963 (N_37963,N_37033,N_37148);
nand U37964 (N_37964,N_37141,N_37282);
nand U37965 (N_37965,N_37021,N_37460);
and U37966 (N_37966,N_37447,N_37392);
xor U37967 (N_37967,N_37207,N_37416);
nand U37968 (N_37968,N_37403,N_37190);
nor U37969 (N_37969,N_37052,N_37070);
or U37970 (N_37970,N_37216,N_37330);
and U37971 (N_37971,N_37264,N_37388);
nand U37972 (N_37972,N_37214,N_37416);
xnor U37973 (N_37973,N_37076,N_37166);
nor U37974 (N_37974,N_37360,N_37472);
xor U37975 (N_37975,N_37083,N_37205);
nor U37976 (N_37976,N_37096,N_37496);
nor U37977 (N_37977,N_37100,N_37364);
xor U37978 (N_37978,N_37469,N_37046);
nand U37979 (N_37979,N_37229,N_37289);
and U37980 (N_37980,N_37105,N_37303);
nand U37981 (N_37981,N_37343,N_37483);
nand U37982 (N_37982,N_37149,N_37345);
or U37983 (N_37983,N_37172,N_37112);
nand U37984 (N_37984,N_37293,N_37034);
or U37985 (N_37985,N_37070,N_37394);
nor U37986 (N_37986,N_37005,N_37057);
nand U37987 (N_37987,N_37300,N_37312);
nor U37988 (N_37988,N_37277,N_37014);
nand U37989 (N_37989,N_37266,N_37045);
or U37990 (N_37990,N_37125,N_37434);
nand U37991 (N_37991,N_37453,N_37020);
nor U37992 (N_37992,N_37182,N_37094);
xnor U37993 (N_37993,N_37030,N_37162);
xnor U37994 (N_37994,N_37033,N_37052);
or U37995 (N_37995,N_37003,N_37032);
nand U37996 (N_37996,N_37485,N_37009);
and U37997 (N_37997,N_37253,N_37085);
and U37998 (N_37998,N_37008,N_37468);
and U37999 (N_37999,N_37212,N_37480);
or U38000 (N_38000,N_37930,N_37770);
nor U38001 (N_38001,N_37679,N_37720);
or U38002 (N_38002,N_37558,N_37963);
nor U38003 (N_38003,N_37813,N_37611);
nor U38004 (N_38004,N_37879,N_37956);
nor U38005 (N_38005,N_37683,N_37772);
xor U38006 (N_38006,N_37723,N_37912);
xor U38007 (N_38007,N_37844,N_37917);
nor U38008 (N_38008,N_37985,N_37767);
and U38009 (N_38009,N_37977,N_37549);
xnor U38010 (N_38010,N_37906,N_37633);
xor U38011 (N_38011,N_37916,N_37808);
nand U38012 (N_38012,N_37730,N_37557);
and U38013 (N_38013,N_37714,N_37654);
nor U38014 (N_38014,N_37957,N_37626);
nand U38015 (N_38015,N_37920,N_37617);
or U38016 (N_38016,N_37527,N_37729);
xnor U38017 (N_38017,N_37867,N_37817);
xnor U38018 (N_38018,N_37843,N_37888);
and U38019 (N_38019,N_37555,N_37775);
nand U38020 (N_38020,N_37990,N_37783);
nor U38021 (N_38021,N_37933,N_37700);
nand U38022 (N_38022,N_37824,N_37809);
xor U38023 (N_38023,N_37771,N_37741);
or U38024 (N_38024,N_37885,N_37588);
nand U38025 (N_38025,N_37690,N_37810);
or U38026 (N_38026,N_37955,N_37922);
or U38027 (N_38027,N_37797,N_37623);
nor U38028 (N_38028,N_37900,N_37951);
nand U38029 (N_38029,N_37925,N_37876);
or U38030 (N_38030,N_37711,N_37836);
and U38031 (N_38031,N_37942,N_37508);
xnor U38032 (N_38032,N_37969,N_37758);
nor U38033 (N_38033,N_37596,N_37866);
or U38034 (N_38034,N_37560,N_37796);
or U38035 (N_38035,N_37563,N_37791);
nand U38036 (N_38036,N_37535,N_37891);
and U38037 (N_38037,N_37948,N_37822);
xnor U38038 (N_38038,N_37570,N_37649);
nor U38039 (N_38039,N_37832,N_37864);
and U38040 (N_38040,N_37890,N_37859);
xnor U38041 (N_38041,N_37695,N_37556);
nand U38042 (N_38042,N_37537,N_37904);
nor U38043 (N_38043,N_37503,N_37637);
nand U38044 (N_38044,N_37678,N_37785);
and U38045 (N_38045,N_37505,N_37657);
or U38046 (N_38046,N_37840,N_37681);
nor U38047 (N_38047,N_37782,N_37786);
nand U38048 (N_38048,N_37950,N_37574);
or U38049 (N_38049,N_37746,N_37788);
nand U38050 (N_38050,N_37874,N_37708);
or U38051 (N_38051,N_37510,N_37940);
nor U38052 (N_38052,N_37567,N_37697);
or U38053 (N_38053,N_37909,N_37754);
nor U38054 (N_38054,N_37982,N_37965);
xnor U38055 (N_38055,N_37750,N_37628);
or U38056 (N_38056,N_37924,N_37938);
or U38057 (N_38057,N_37725,N_37554);
nand U38058 (N_38058,N_37576,N_37845);
nand U38059 (N_38059,N_37870,N_37862);
and U38060 (N_38060,N_37854,N_37531);
nor U38061 (N_38061,N_37997,N_37581);
nand U38062 (N_38062,N_37675,N_37651);
or U38063 (N_38063,N_37835,N_37523);
and U38064 (N_38064,N_37639,N_37993);
or U38065 (N_38065,N_37768,N_37937);
nor U38066 (N_38066,N_37525,N_37911);
and U38067 (N_38067,N_37672,N_37552);
xor U38068 (N_38068,N_37826,N_37949);
xnor U38069 (N_38069,N_37934,N_37850);
nor U38070 (N_38070,N_37627,N_37605);
nand U38071 (N_38071,N_37773,N_37636);
nand U38072 (N_38072,N_37536,N_37595);
nor U38073 (N_38073,N_37702,N_37842);
nand U38074 (N_38074,N_37829,N_37670);
nor U38075 (N_38075,N_37550,N_37910);
xnor U38076 (N_38076,N_37926,N_37717);
or U38077 (N_38077,N_37721,N_37971);
nand U38078 (N_38078,N_37852,N_37919);
xnor U38079 (N_38079,N_37787,N_37841);
or U38080 (N_38080,N_37865,N_37684);
nor U38081 (N_38081,N_37590,N_37763);
nor U38082 (N_38082,N_37792,N_37929);
nand U38083 (N_38083,N_37507,N_37784);
nor U38084 (N_38084,N_37533,N_37582);
nor U38085 (N_38085,N_37954,N_37722);
or U38086 (N_38086,N_37502,N_37812);
nor U38087 (N_38087,N_37846,N_37914);
nand U38088 (N_38088,N_37968,N_37984);
nand U38089 (N_38089,N_37749,N_37551);
xor U38090 (N_38090,N_37814,N_37794);
nand U38091 (N_38091,N_37534,N_37587);
nor U38092 (N_38092,N_37732,N_37903);
nand U38093 (N_38093,N_37935,N_37540);
nor U38094 (N_38094,N_37641,N_37830);
and U38095 (N_38095,N_37674,N_37882);
or U38096 (N_38096,N_37710,N_37779);
nor U38097 (N_38097,N_37728,N_37789);
and U38098 (N_38098,N_37542,N_37652);
nor U38099 (N_38099,N_37855,N_37894);
xor U38100 (N_38100,N_37622,N_37584);
nor U38101 (N_38101,N_37631,N_37868);
nand U38102 (N_38102,N_37774,N_37851);
xnor U38103 (N_38103,N_37877,N_37757);
or U38104 (N_38104,N_37946,N_37705);
nand U38105 (N_38105,N_37593,N_37665);
nand U38106 (N_38106,N_37734,N_37802);
nor U38107 (N_38107,N_37673,N_37528);
nor U38108 (N_38108,N_37943,N_37878);
and U38109 (N_38109,N_37765,N_37983);
and U38110 (N_38110,N_37875,N_37820);
or U38111 (N_38111,N_37823,N_37513);
nor U38112 (N_38112,N_37847,N_37941);
xnor U38113 (N_38113,N_37514,N_37953);
and U38114 (N_38114,N_37889,N_37501);
or U38115 (N_38115,N_37667,N_37966);
nand U38116 (N_38116,N_37518,N_37693);
and U38117 (N_38117,N_37837,N_37669);
nor U38118 (N_38118,N_37543,N_37892);
nand U38119 (N_38119,N_37902,N_37987);
nor U38120 (N_38120,N_37530,N_37908);
or U38121 (N_38121,N_37973,N_37995);
nor U38122 (N_38122,N_37572,N_37872);
nand U38123 (N_38123,N_37740,N_37566);
nand U38124 (N_38124,N_37539,N_37704);
or U38125 (N_38125,N_37603,N_37524);
nand U38126 (N_38126,N_37992,N_37896);
and U38127 (N_38127,N_37688,N_37568);
xnor U38128 (N_38128,N_37660,N_37629);
and U38129 (N_38129,N_37585,N_37819);
xnor U38130 (N_38130,N_37577,N_37806);
nand U38131 (N_38131,N_37613,N_37610);
nor U38132 (N_38132,N_37517,N_37959);
and U38133 (N_38133,N_37805,N_37803);
and U38134 (N_38134,N_37743,N_37994);
and U38135 (N_38135,N_37532,N_37913);
nand U38136 (N_38136,N_37619,N_37759);
nand U38137 (N_38137,N_37547,N_37664);
nor U38138 (N_38138,N_37893,N_37918);
xnor U38139 (N_38139,N_37860,N_37962);
or U38140 (N_38140,N_37591,N_37668);
and U38141 (N_38141,N_37856,N_37831);
xor U38142 (N_38142,N_37635,N_37607);
nor U38143 (N_38143,N_37761,N_37748);
nor U38144 (N_38144,N_37696,N_37927);
nand U38145 (N_38145,N_37816,N_37762);
nor U38146 (N_38146,N_37907,N_37975);
xnor U38147 (N_38147,N_37998,N_37601);
or U38148 (N_38148,N_37663,N_37811);
xor U38149 (N_38149,N_37932,N_37515);
nand U38150 (N_38150,N_37931,N_37905);
and U38151 (N_38151,N_37646,N_37602);
nor U38152 (N_38152,N_37545,N_37519);
nand U38153 (N_38153,N_37511,N_37978);
nand U38154 (N_38154,N_37839,N_37571);
nand U38155 (N_38155,N_37790,N_37915);
nand U38156 (N_38156,N_37724,N_37769);
xnor U38157 (N_38157,N_37945,N_37682);
nor U38158 (N_38158,N_37658,N_37884);
and U38159 (N_38159,N_37939,N_37686);
xnor U38160 (N_38160,N_37541,N_37974);
xor U38161 (N_38161,N_37716,N_37947);
and U38162 (N_38162,N_37642,N_37742);
nor U38163 (N_38163,N_37726,N_37707);
xor U38164 (N_38164,N_37638,N_37731);
nor U38165 (N_38165,N_37881,N_37827);
nor U38166 (N_38166,N_37921,N_37592);
xnor U38167 (N_38167,N_37848,N_37701);
or U38168 (N_38168,N_37579,N_37739);
nand U38169 (N_38169,N_37640,N_37899);
xor U38170 (N_38170,N_37880,N_37575);
xnor U38171 (N_38171,N_37718,N_37834);
xor U38172 (N_38172,N_37544,N_37871);
nand U38173 (N_38173,N_37516,N_37586);
nand U38174 (N_38174,N_37677,N_37719);
nand U38175 (N_38175,N_37793,N_37744);
xnor U38176 (N_38176,N_37996,N_37818);
and U38177 (N_38177,N_37777,N_37833);
xnor U38178 (N_38178,N_37751,N_37869);
nor U38179 (N_38179,N_37624,N_37546);
nand U38180 (N_38180,N_37647,N_37807);
nor U38181 (N_38181,N_37618,N_37764);
xnor U38182 (N_38182,N_37952,N_37600);
xor U38183 (N_38183,N_37801,N_37760);
nor U38184 (N_38184,N_37804,N_37800);
or U38185 (N_38185,N_37615,N_37895);
or U38186 (N_38186,N_37573,N_37736);
xnor U38187 (N_38187,N_37979,N_37778);
or U38188 (N_38188,N_37713,N_37561);
nand U38189 (N_38189,N_37632,N_37653);
xor U38190 (N_38190,N_37897,N_37662);
xor U38191 (N_38191,N_37529,N_37861);
nor U38192 (N_38192,N_37815,N_37825);
nor U38193 (N_38193,N_37886,N_37564);
or U38194 (N_38194,N_37659,N_37597);
and U38195 (N_38195,N_37691,N_37648);
nor U38196 (N_38196,N_37616,N_37988);
nand U38197 (N_38197,N_37614,N_37901);
nor U38198 (N_38198,N_37512,N_37689);
or U38199 (N_38199,N_37735,N_37620);
or U38200 (N_38200,N_37509,N_37526);
and U38201 (N_38201,N_37500,N_37521);
nor U38202 (N_38202,N_37655,N_37604);
nand U38203 (N_38203,N_37752,N_37583);
or U38204 (N_38204,N_37780,N_37980);
nand U38205 (N_38205,N_37643,N_37853);
nand U38206 (N_38206,N_37928,N_37863);
xnor U38207 (N_38207,N_37766,N_37709);
or U38208 (N_38208,N_37873,N_37589);
or U38209 (N_38209,N_37504,N_37645);
or U38210 (N_38210,N_37733,N_37828);
nor U38211 (N_38211,N_37599,N_37999);
and U38212 (N_38212,N_37738,N_37976);
nor U38213 (N_38213,N_37676,N_37961);
xnor U38214 (N_38214,N_37661,N_37644);
and U38215 (N_38215,N_37548,N_37737);
nand U38216 (N_38216,N_37795,N_37578);
nand U38217 (N_38217,N_37506,N_37609);
nand U38218 (N_38218,N_37522,N_37703);
and U38219 (N_38219,N_37612,N_37964);
or U38220 (N_38220,N_37608,N_37821);
nor U38221 (N_38221,N_37944,N_37650);
nor U38222 (N_38222,N_37630,N_37656);
nand U38223 (N_38223,N_37598,N_37569);
xor U38224 (N_38224,N_37958,N_37680);
nand U38225 (N_38225,N_37936,N_37967);
nand U38226 (N_38226,N_37986,N_37747);
nor U38227 (N_38227,N_37685,N_37755);
nor U38228 (N_38228,N_37692,N_37606);
nand U38229 (N_38229,N_37520,N_37923);
xor U38230 (N_38230,N_37671,N_37666);
nor U38231 (N_38231,N_37960,N_37857);
or U38232 (N_38232,N_37756,N_37991);
xor U38233 (N_38233,N_37553,N_37883);
nand U38234 (N_38234,N_37687,N_37972);
nand U38235 (N_38235,N_37799,N_37849);
and U38236 (N_38236,N_37699,N_37981);
xor U38237 (N_38237,N_37580,N_37565);
xnor U38238 (N_38238,N_37776,N_37798);
or U38239 (N_38239,N_37745,N_37727);
or U38240 (N_38240,N_37753,N_37559);
nand U38241 (N_38241,N_37781,N_37898);
and U38242 (N_38242,N_37694,N_37594);
and U38243 (N_38243,N_37887,N_37706);
nand U38244 (N_38244,N_37634,N_37838);
or U38245 (N_38245,N_37625,N_37989);
xnor U38246 (N_38246,N_37621,N_37698);
nand U38247 (N_38247,N_37562,N_37858);
xor U38248 (N_38248,N_37715,N_37538);
or U38249 (N_38249,N_37970,N_37712);
nand U38250 (N_38250,N_37743,N_37990);
or U38251 (N_38251,N_37734,N_37888);
or U38252 (N_38252,N_37567,N_37680);
and U38253 (N_38253,N_37524,N_37573);
and U38254 (N_38254,N_37708,N_37886);
nand U38255 (N_38255,N_37849,N_37522);
or U38256 (N_38256,N_37728,N_37824);
nand U38257 (N_38257,N_37785,N_37806);
xor U38258 (N_38258,N_37924,N_37761);
nor U38259 (N_38259,N_37904,N_37834);
nand U38260 (N_38260,N_37600,N_37875);
and U38261 (N_38261,N_37537,N_37955);
and U38262 (N_38262,N_37975,N_37839);
xor U38263 (N_38263,N_37765,N_37976);
xnor U38264 (N_38264,N_37518,N_37543);
or U38265 (N_38265,N_37545,N_37647);
or U38266 (N_38266,N_37847,N_37893);
xnor U38267 (N_38267,N_37634,N_37608);
xnor U38268 (N_38268,N_37997,N_37641);
nor U38269 (N_38269,N_37634,N_37540);
xor U38270 (N_38270,N_37925,N_37995);
nand U38271 (N_38271,N_37565,N_37726);
and U38272 (N_38272,N_37534,N_37589);
and U38273 (N_38273,N_37626,N_37664);
xnor U38274 (N_38274,N_37849,N_37587);
or U38275 (N_38275,N_37570,N_37863);
or U38276 (N_38276,N_37884,N_37628);
xnor U38277 (N_38277,N_37505,N_37927);
nor U38278 (N_38278,N_37950,N_37544);
nand U38279 (N_38279,N_37736,N_37745);
nor U38280 (N_38280,N_37553,N_37550);
nand U38281 (N_38281,N_37687,N_37994);
or U38282 (N_38282,N_37644,N_37881);
and U38283 (N_38283,N_37712,N_37741);
and U38284 (N_38284,N_37803,N_37500);
or U38285 (N_38285,N_37701,N_37863);
xnor U38286 (N_38286,N_37565,N_37746);
or U38287 (N_38287,N_37882,N_37782);
nor U38288 (N_38288,N_37931,N_37996);
and U38289 (N_38289,N_37879,N_37746);
xor U38290 (N_38290,N_37518,N_37818);
and U38291 (N_38291,N_37845,N_37659);
and U38292 (N_38292,N_37507,N_37669);
nor U38293 (N_38293,N_37594,N_37569);
or U38294 (N_38294,N_37713,N_37959);
or U38295 (N_38295,N_37722,N_37781);
or U38296 (N_38296,N_37870,N_37636);
and U38297 (N_38297,N_37978,N_37968);
nand U38298 (N_38298,N_37738,N_37971);
xor U38299 (N_38299,N_37888,N_37953);
or U38300 (N_38300,N_37940,N_37712);
or U38301 (N_38301,N_37892,N_37648);
xnor U38302 (N_38302,N_37762,N_37740);
nor U38303 (N_38303,N_37896,N_37779);
or U38304 (N_38304,N_37771,N_37513);
nand U38305 (N_38305,N_37991,N_37967);
nand U38306 (N_38306,N_37803,N_37971);
or U38307 (N_38307,N_37841,N_37825);
nor U38308 (N_38308,N_37590,N_37662);
or U38309 (N_38309,N_37693,N_37952);
nor U38310 (N_38310,N_37750,N_37944);
and U38311 (N_38311,N_37774,N_37602);
xnor U38312 (N_38312,N_37545,N_37882);
or U38313 (N_38313,N_37522,N_37978);
xnor U38314 (N_38314,N_37783,N_37958);
and U38315 (N_38315,N_37905,N_37681);
and U38316 (N_38316,N_37869,N_37573);
xnor U38317 (N_38317,N_37576,N_37822);
or U38318 (N_38318,N_37769,N_37664);
nand U38319 (N_38319,N_37814,N_37658);
and U38320 (N_38320,N_37664,N_37562);
xnor U38321 (N_38321,N_37522,N_37783);
nor U38322 (N_38322,N_37634,N_37668);
and U38323 (N_38323,N_37872,N_37833);
and U38324 (N_38324,N_37699,N_37674);
xnor U38325 (N_38325,N_37576,N_37511);
and U38326 (N_38326,N_37932,N_37518);
nand U38327 (N_38327,N_37652,N_37608);
and U38328 (N_38328,N_37741,N_37579);
xnor U38329 (N_38329,N_37606,N_37919);
or U38330 (N_38330,N_37951,N_37741);
nand U38331 (N_38331,N_37946,N_37837);
xor U38332 (N_38332,N_37997,N_37743);
nor U38333 (N_38333,N_37660,N_37822);
and U38334 (N_38334,N_37850,N_37735);
or U38335 (N_38335,N_37988,N_37964);
nand U38336 (N_38336,N_37667,N_37829);
xnor U38337 (N_38337,N_37852,N_37992);
nand U38338 (N_38338,N_37718,N_37661);
nand U38339 (N_38339,N_37724,N_37752);
and U38340 (N_38340,N_37689,N_37633);
nand U38341 (N_38341,N_37994,N_37790);
and U38342 (N_38342,N_37809,N_37745);
xor U38343 (N_38343,N_37925,N_37637);
or U38344 (N_38344,N_37965,N_37685);
and U38345 (N_38345,N_37882,N_37886);
and U38346 (N_38346,N_37780,N_37994);
xor U38347 (N_38347,N_37766,N_37594);
nor U38348 (N_38348,N_37669,N_37805);
and U38349 (N_38349,N_37546,N_37531);
xnor U38350 (N_38350,N_37856,N_37745);
nor U38351 (N_38351,N_37741,N_37855);
nand U38352 (N_38352,N_37610,N_37639);
xnor U38353 (N_38353,N_37727,N_37721);
xor U38354 (N_38354,N_37961,N_37577);
nor U38355 (N_38355,N_37769,N_37803);
or U38356 (N_38356,N_37662,N_37875);
nor U38357 (N_38357,N_37734,N_37883);
nand U38358 (N_38358,N_37833,N_37691);
nor U38359 (N_38359,N_37613,N_37707);
xnor U38360 (N_38360,N_37534,N_37912);
nand U38361 (N_38361,N_37530,N_37590);
nand U38362 (N_38362,N_37932,N_37912);
nor U38363 (N_38363,N_37880,N_37980);
nor U38364 (N_38364,N_37690,N_37660);
or U38365 (N_38365,N_37545,N_37913);
and U38366 (N_38366,N_37543,N_37810);
and U38367 (N_38367,N_37686,N_37942);
nand U38368 (N_38368,N_37914,N_37706);
nor U38369 (N_38369,N_37814,N_37534);
nor U38370 (N_38370,N_37897,N_37946);
xnor U38371 (N_38371,N_37858,N_37976);
nand U38372 (N_38372,N_37666,N_37817);
nand U38373 (N_38373,N_37806,N_37815);
or U38374 (N_38374,N_37828,N_37740);
nand U38375 (N_38375,N_37761,N_37662);
or U38376 (N_38376,N_37546,N_37618);
nand U38377 (N_38377,N_37673,N_37971);
or U38378 (N_38378,N_37597,N_37808);
or U38379 (N_38379,N_37610,N_37859);
nand U38380 (N_38380,N_37859,N_37559);
nand U38381 (N_38381,N_37714,N_37743);
nand U38382 (N_38382,N_37730,N_37713);
nor U38383 (N_38383,N_37701,N_37657);
xnor U38384 (N_38384,N_37750,N_37780);
xnor U38385 (N_38385,N_37771,N_37573);
nor U38386 (N_38386,N_37992,N_37915);
xor U38387 (N_38387,N_37997,N_37705);
nand U38388 (N_38388,N_37993,N_37890);
and U38389 (N_38389,N_37716,N_37637);
or U38390 (N_38390,N_37794,N_37546);
xnor U38391 (N_38391,N_37593,N_37837);
xor U38392 (N_38392,N_37877,N_37928);
nand U38393 (N_38393,N_37713,N_37722);
or U38394 (N_38394,N_37779,N_37667);
nor U38395 (N_38395,N_37621,N_37816);
xnor U38396 (N_38396,N_37998,N_37744);
nand U38397 (N_38397,N_37551,N_37670);
and U38398 (N_38398,N_37966,N_37936);
xnor U38399 (N_38399,N_37842,N_37633);
and U38400 (N_38400,N_37537,N_37916);
nand U38401 (N_38401,N_37930,N_37631);
or U38402 (N_38402,N_37609,N_37678);
or U38403 (N_38403,N_37504,N_37789);
nand U38404 (N_38404,N_37655,N_37660);
nor U38405 (N_38405,N_37976,N_37552);
and U38406 (N_38406,N_37848,N_37875);
and U38407 (N_38407,N_37562,N_37805);
xor U38408 (N_38408,N_37865,N_37761);
and U38409 (N_38409,N_37659,N_37580);
or U38410 (N_38410,N_37888,N_37871);
nor U38411 (N_38411,N_37600,N_37804);
and U38412 (N_38412,N_37641,N_37714);
or U38413 (N_38413,N_37633,N_37650);
xor U38414 (N_38414,N_37700,N_37895);
nand U38415 (N_38415,N_37923,N_37546);
nor U38416 (N_38416,N_37868,N_37763);
nor U38417 (N_38417,N_37792,N_37963);
or U38418 (N_38418,N_37633,N_37988);
xnor U38419 (N_38419,N_37900,N_37727);
nand U38420 (N_38420,N_37841,N_37635);
xnor U38421 (N_38421,N_37879,N_37925);
or U38422 (N_38422,N_37508,N_37832);
and U38423 (N_38423,N_37807,N_37976);
nor U38424 (N_38424,N_37627,N_37838);
nand U38425 (N_38425,N_37951,N_37516);
and U38426 (N_38426,N_37629,N_37845);
nor U38427 (N_38427,N_37719,N_37932);
or U38428 (N_38428,N_37722,N_37770);
xnor U38429 (N_38429,N_37765,N_37941);
and U38430 (N_38430,N_37751,N_37735);
or U38431 (N_38431,N_37693,N_37656);
or U38432 (N_38432,N_37970,N_37798);
or U38433 (N_38433,N_37863,N_37908);
and U38434 (N_38434,N_37815,N_37999);
and U38435 (N_38435,N_37516,N_37735);
nor U38436 (N_38436,N_37513,N_37602);
and U38437 (N_38437,N_37628,N_37607);
xnor U38438 (N_38438,N_37705,N_37837);
nand U38439 (N_38439,N_37610,N_37989);
nand U38440 (N_38440,N_37934,N_37809);
nand U38441 (N_38441,N_37541,N_37996);
nor U38442 (N_38442,N_37738,N_37641);
nor U38443 (N_38443,N_37652,N_37897);
and U38444 (N_38444,N_37508,N_37673);
xor U38445 (N_38445,N_37954,N_37911);
or U38446 (N_38446,N_37657,N_37937);
and U38447 (N_38447,N_37635,N_37719);
and U38448 (N_38448,N_37753,N_37828);
and U38449 (N_38449,N_37775,N_37677);
and U38450 (N_38450,N_37702,N_37972);
nand U38451 (N_38451,N_37510,N_37847);
xnor U38452 (N_38452,N_37971,N_37550);
xor U38453 (N_38453,N_37822,N_37611);
xor U38454 (N_38454,N_37662,N_37673);
or U38455 (N_38455,N_37904,N_37586);
nand U38456 (N_38456,N_37822,N_37689);
and U38457 (N_38457,N_37848,N_37572);
nand U38458 (N_38458,N_37650,N_37643);
nor U38459 (N_38459,N_37965,N_37859);
and U38460 (N_38460,N_37677,N_37653);
xor U38461 (N_38461,N_37737,N_37826);
nor U38462 (N_38462,N_37606,N_37826);
and U38463 (N_38463,N_37752,N_37888);
nor U38464 (N_38464,N_37767,N_37586);
xnor U38465 (N_38465,N_37792,N_37946);
and U38466 (N_38466,N_37956,N_37773);
nand U38467 (N_38467,N_37776,N_37757);
nand U38468 (N_38468,N_37957,N_37967);
nand U38469 (N_38469,N_37559,N_37745);
and U38470 (N_38470,N_37922,N_37923);
and U38471 (N_38471,N_37994,N_37699);
nor U38472 (N_38472,N_37953,N_37722);
and U38473 (N_38473,N_37770,N_37880);
or U38474 (N_38474,N_37703,N_37805);
or U38475 (N_38475,N_37857,N_37941);
nor U38476 (N_38476,N_37945,N_37870);
nor U38477 (N_38477,N_37916,N_37965);
or U38478 (N_38478,N_37678,N_37737);
or U38479 (N_38479,N_37595,N_37919);
or U38480 (N_38480,N_37595,N_37836);
xor U38481 (N_38481,N_37582,N_37605);
and U38482 (N_38482,N_37632,N_37773);
xnor U38483 (N_38483,N_37915,N_37787);
or U38484 (N_38484,N_37611,N_37673);
nand U38485 (N_38485,N_37879,N_37906);
xor U38486 (N_38486,N_37690,N_37806);
nand U38487 (N_38487,N_37713,N_37726);
xnor U38488 (N_38488,N_37814,N_37751);
and U38489 (N_38489,N_37685,N_37811);
or U38490 (N_38490,N_37912,N_37572);
xor U38491 (N_38491,N_37540,N_37589);
nor U38492 (N_38492,N_37579,N_37972);
xnor U38493 (N_38493,N_37791,N_37997);
nor U38494 (N_38494,N_37641,N_37585);
or U38495 (N_38495,N_37633,N_37622);
nand U38496 (N_38496,N_37898,N_37584);
xnor U38497 (N_38497,N_37911,N_37625);
or U38498 (N_38498,N_37923,N_37537);
nand U38499 (N_38499,N_37603,N_37714);
nor U38500 (N_38500,N_38321,N_38394);
xnor U38501 (N_38501,N_38352,N_38258);
nor U38502 (N_38502,N_38081,N_38220);
xnor U38503 (N_38503,N_38201,N_38048);
and U38504 (N_38504,N_38218,N_38168);
and U38505 (N_38505,N_38059,N_38298);
and U38506 (N_38506,N_38024,N_38358);
nor U38507 (N_38507,N_38290,N_38291);
or U38508 (N_38508,N_38406,N_38126);
xnor U38509 (N_38509,N_38134,N_38245);
nor U38510 (N_38510,N_38075,N_38392);
or U38511 (N_38511,N_38409,N_38431);
or U38512 (N_38512,N_38163,N_38248);
nor U38513 (N_38513,N_38100,N_38178);
nor U38514 (N_38514,N_38139,N_38354);
nor U38515 (N_38515,N_38181,N_38198);
nand U38516 (N_38516,N_38088,N_38050);
xnor U38517 (N_38517,N_38491,N_38019);
nor U38518 (N_38518,N_38222,N_38403);
xnor U38519 (N_38519,N_38451,N_38240);
nor U38520 (N_38520,N_38383,N_38343);
or U38521 (N_38521,N_38293,N_38184);
nor U38522 (N_38522,N_38195,N_38459);
or U38523 (N_38523,N_38113,N_38123);
and U38524 (N_38524,N_38225,N_38111);
nor U38525 (N_38525,N_38033,N_38242);
or U38526 (N_38526,N_38036,N_38216);
and U38527 (N_38527,N_38094,N_38040);
nor U38528 (N_38528,N_38210,N_38294);
nor U38529 (N_38529,N_38250,N_38054);
xnor U38530 (N_38530,N_38212,N_38109);
nor U38531 (N_38531,N_38327,N_38000);
nor U38532 (N_38532,N_38344,N_38364);
and U38533 (N_38533,N_38389,N_38132);
nand U38534 (N_38534,N_38331,N_38230);
or U38535 (N_38535,N_38027,N_38122);
xnor U38536 (N_38536,N_38265,N_38428);
or U38537 (N_38537,N_38485,N_38009);
xor U38538 (N_38538,N_38297,N_38053);
and U38539 (N_38539,N_38227,N_38481);
nand U38540 (N_38540,N_38467,N_38118);
or U38541 (N_38541,N_38234,N_38158);
and U38542 (N_38542,N_38285,N_38275);
or U38543 (N_38543,N_38056,N_38253);
nor U38544 (N_38544,N_38270,N_38474);
xnor U38545 (N_38545,N_38315,N_38464);
nand U38546 (N_38546,N_38175,N_38317);
and U38547 (N_38547,N_38404,N_38420);
nor U38548 (N_38548,N_38470,N_38278);
nand U38549 (N_38549,N_38399,N_38269);
or U38550 (N_38550,N_38255,N_38400);
and U38551 (N_38551,N_38271,N_38351);
nor U38552 (N_38552,N_38076,N_38260);
nand U38553 (N_38553,N_38197,N_38486);
nor U38554 (N_38554,N_38267,N_38412);
and U38555 (N_38555,N_38207,N_38105);
nor U38556 (N_38556,N_38396,N_38405);
nand U38557 (N_38557,N_38476,N_38487);
xor U38558 (N_38558,N_38376,N_38146);
and U38559 (N_38559,N_38098,N_38356);
or U38560 (N_38560,N_38115,N_38429);
or U38561 (N_38561,N_38078,N_38068);
nor U38562 (N_38562,N_38138,N_38127);
xnor U38563 (N_38563,N_38017,N_38092);
nand U38564 (N_38564,N_38208,N_38183);
or U38565 (N_38565,N_38103,N_38243);
and U38566 (N_38566,N_38339,N_38030);
nand U38567 (N_38567,N_38016,N_38455);
nor U38568 (N_38568,N_38223,N_38147);
or U38569 (N_38569,N_38211,N_38273);
nand U38570 (N_38570,N_38203,N_38161);
or U38571 (N_38571,N_38277,N_38005);
nor U38572 (N_38572,N_38087,N_38137);
nand U38573 (N_38573,N_38112,N_38292);
xnor U38574 (N_38574,N_38148,N_38438);
and U38575 (N_38575,N_38437,N_38155);
xor U38576 (N_38576,N_38488,N_38099);
xor U38577 (N_38577,N_38104,N_38310);
and U38578 (N_38578,N_38414,N_38397);
and U38579 (N_38579,N_38282,N_38046);
xnor U38580 (N_38580,N_38280,N_38346);
xnor U38581 (N_38581,N_38372,N_38492);
and U38582 (N_38582,N_38300,N_38002);
xor U38583 (N_38583,N_38173,N_38261);
nor U38584 (N_38584,N_38215,N_38468);
nand U38585 (N_38585,N_38170,N_38106);
and U38586 (N_38586,N_38417,N_38375);
and U38587 (N_38587,N_38365,N_38171);
nand U38588 (N_38588,N_38257,N_38043);
xor U38589 (N_38589,N_38453,N_38164);
nand U38590 (N_38590,N_38249,N_38499);
or U38591 (N_38591,N_38482,N_38107);
and U38592 (N_38592,N_38169,N_38373);
nand U38593 (N_38593,N_38345,N_38001);
nand U38594 (N_38594,N_38086,N_38286);
nor U38595 (N_38595,N_38469,N_38239);
and U38596 (N_38596,N_38384,N_38303);
nor U38597 (N_38597,N_38237,N_38456);
nor U38598 (N_38598,N_38063,N_38312);
or U38599 (N_38599,N_38313,N_38307);
xor U38600 (N_38600,N_38185,N_38496);
xor U38601 (N_38601,N_38039,N_38125);
nand U38602 (N_38602,N_38135,N_38333);
nor U38603 (N_38603,N_38288,N_38308);
nand U38604 (N_38604,N_38374,N_38415);
nor U38605 (N_38605,N_38199,N_38334);
nor U38606 (N_38606,N_38196,N_38316);
nand U38607 (N_38607,N_38152,N_38419);
nand U38608 (N_38608,N_38348,N_38436);
nand U38609 (N_38609,N_38318,N_38435);
xor U38610 (N_38610,N_38247,N_38091);
or U38611 (N_38611,N_38241,N_38069);
nand U38612 (N_38612,N_38390,N_38445);
or U38613 (N_38613,N_38079,N_38149);
and U38614 (N_38614,N_38205,N_38131);
and U38615 (N_38615,N_38160,N_38110);
and U38616 (N_38616,N_38304,N_38309);
nor U38617 (N_38617,N_38336,N_38454);
or U38618 (N_38618,N_38073,N_38153);
nand U38619 (N_38619,N_38363,N_38264);
nor U38620 (N_38620,N_38055,N_38355);
and U38621 (N_38621,N_38129,N_38187);
nor U38622 (N_38622,N_38366,N_38433);
xnor U38623 (N_38623,N_38130,N_38449);
and U38624 (N_38624,N_38461,N_38434);
and U38625 (N_38625,N_38335,N_38095);
nand U38626 (N_38626,N_38026,N_38402);
xor U38627 (N_38627,N_38289,N_38179);
or U38628 (N_38628,N_38012,N_38480);
xnor U38629 (N_38629,N_38314,N_38357);
xnor U38630 (N_38630,N_38121,N_38359);
xnor U38631 (N_38631,N_38497,N_38188);
and U38632 (N_38632,N_38176,N_38219);
nand U38633 (N_38633,N_38042,N_38066);
and U38634 (N_38634,N_38368,N_38200);
nor U38635 (N_38635,N_38256,N_38159);
and U38636 (N_38636,N_38157,N_38064);
or U38637 (N_38637,N_38395,N_38360);
xor U38638 (N_38638,N_38154,N_38263);
and U38639 (N_38639,N_38254,N_38114);
and U38640 (N_38640,N_38031,N_38057);
and U38641 (N_38641,N_38302,N_38432);
or U38642 (N_38642,N_38167,N_38072);
nor U38643 (N_38643,N_38025,N_38180);
and U38644 (N_38644,N_38077,N_38172);
nand U38645 (N_38645,N_38022,N_38462);
or U38646 (N_38646,N_38332,N_38477);
and U38647 (N_38647,N_38259,N_38382);
or U38648 (N_38648,N_38003,N_38466);
nor U38649 (N_38649,N_38371,N_38388);
or U38650 (N_38650,N_38440,N_38349);
nand U38651 (N_38651,N_38401,N_38380);
nand U38652 (N_38652,N_38150,N_38323);
nand U38653 (N_38653,N_38423,N_38191);
or U38654 (N_38654,N_38051,N_38194);
xor U38655 (N_38655,N_38136,N_38301);
nand U38656 (N_38656,N_38108,N_38165);
xnor U38657 (N_38657,N_38441,N_38284);
nor U38658 (N_38658,N_38119,N_38274);
nor U38659 (N_38659,N_38463,N_38037);
or U38660 (N_38660,N_38221,N_38029);
nand U38661 (N_38661,N_38279,N_38452);
nand U38662 (N_38662,N_38007,N_38299);
or U38663 (N_38663,N_38350,N_38262);
or U38664 (N_38664,N_38329,N_38411);
and U38665 (N_38665,N_38319,N_38447);
nor U38666 (N_38666,N_38224,N_38296);
nand U38667 (N_38667,N_38341,N_38479);
nor U38668 (N_38668,N_38228,N_38166);
nand U38669 (N_38669,N_38272,N_38306);
or U38670 (N_38670,N_38338,N_38337);
nand U38671 (N_38671,N_38326,N_38044);
or U38672 (N_38672,N_38379,N_38023);
nand U38673 (N_38673,N_38393,N_38231);
and U38674 (N_38674,N_38067,N_38151);
nor U38675 (N_38675,N_38142,N_38071);
and U38676 (N_38676,N_38252,N_38028);
and U38677 (N_38677,N_38013,N_38421);
and U38678 (N_38678,N_38324,N_38322);
nor U38679 (N_38679,N_38116,N_38102);
and U38680 (N_38680,N_38035,N_38233);
nand U38681 (N_38681,N_38448,N_38268);
or U38682 (N_38682,N_38425,N_38266);
xor U38683 (N_38683,N_38038,N_38192);
xor U38684 (N_38684,N_38422,N_38177);
xnor U38685 (N_38685,N_38101,N_38182);
and U38686 (N_38686,N_38143,N_38353);
or U38687 (N_38687,N_38124,N_38325);
and U38688 (N_38688,N_38251,N_38320);
nor U38689 (N_38689,N_38416,N_38439);
xnor U38690 (N_38690,N_38032,N_38473);
or U38691 (N_38691,N_38156,N_38082);
or U38692 (N_38692,N_38049,N_38287);
xor U38693 (N_38693,N_38213,N_38494);
xor U38694 (N_38694,N_38186,N_38133);
nand U38695 (N_38695,N_38204,N_38045);
and U38696 (N_38696,N_38090,N_38120);
and U38697 (N_38697,N_38483,N_38209);
nand U38698 (N_38698,N_38006,N_38471);
and U38699 (N_38699,N_38342,N_38021);
or U38700 (N_38700,N_38174,N_38229);
nor U38701 (N_38701,N_38189,N_38085);
nor U38702 (N_38702,N_38475,N_38235);
nor U38703 (N_38703,N_38141,N_38232);
nand U38704 (N_38704,N_38460,N_38408);
and U38705 (N_38705,N_38295,N_38244);
or U38706 (N_38706,N_38465,N_38472);
nor U38707 (N_38707,N_38206,N_38442);
xor U38708 (N_38708,N_38093,N_38145);
or U38709 (N_38709,N_38398,N_38387);
nor U38710 (N_38710,N_38238,N_38080);
xor U38711 (N_38711,N_38010,N_38236);
nand U38712 (N_38712,N_38498,N_38061);
and U38713 (N_38713,N_38430,N_38386);
nor U38714 (N_38714,N_38193,N_38281);
or U38715 (N_38715,N_38283,N_38034);
xor U38716 (N_38716,N_38443,N_38015);
nand U38717 (N_38717,N_38381,N_38427);
nor U38718 (N_38718,N_38128,N_38014);
xnor U38719 (N_38719,N_38446,N_38385);
nor U38720 (N_38720,N_38450,N_38089);
or U38721 (N_38721,N_38047,N_38011);
xor U38722 (N_38722,N_38378,N_38495);
or U38723 (N_38723,N_38490,N_38370);
or U38724 (N_38724,N_38484,N_38413);
or U38725 (N_38725,N_38276,N_38020);
or U38726 (N_38726,N_38117,N_38424);
xnor U38727 (N_38727,N_38202,N_38162);
xnor U38728 (N_38728,N_38004,N_38377);
xnor U38729 (N_38729,N_38074,N_38305);
nand U38730 (N_38730,N_38426,N_38362);
and U38731 (N_38731,N_38190,N_38083);
xnor U38732 (N_38732,N_38065,N_38458);
and U38733 (N_38733,N_38391,N_38407);
nand U38734 (N_38734,N_38367,N_38493);
xnor U38735 (N_38735,N_38144,N_38489);
and U38736 (N_38736,N_38361,N_38347);
nor U38737 (N_38737,N_38018,N_38052);
nor U38738 (N_38738,N_38140,N_38478);
nand U38739 (N_38739,N_38097,N_38008);
and U38740 (N_38740,N_38311,N_38084);
xor U38741 (N_38741,N_38070,N_38217);
and U38742 (N_38742,N_38444,N_38330);
xnor U38743 (N_38743,N_38226,N_38062);
xnor U38744 (N_38744,N_38410,N_38060);
or U38745 (N_38745,N_38041,N_38246);
nand U38746 (N_38746,N_38418,N_38058);
nand U38747 (N_38747,N_38340,N_38328);
nand U38748 (N_38748,N_38096,N_38214);
or U38749 (N_38749,N_38369,N_38457);
and U38750 (N_38750,N_38046,N_38469);
or U38751 (N_38751,N_38291,N_38111);
nor U38752 (N_38752,N_38275,N_38318);
or U38753 (N_38753,N_38226,N_38232);
nor U38754 (N_38754,N_38037,N_38160);
nor U38755 (N_38755,N_38447,N_38402);
or U38756 (N_38756,N_38045,N_38305);
xnor U38757 (N_38757,N_38479,N_38192);
nand U38758 (N_38758,N_38393,N_38427);
or U38759 (N_38759,N_38327,N_38354);
and U38760 (N_38760,N_38350,N_38209);
nand U38761 (N_38761,N_38496,N_38446);
xor U38762 (N_38762,N_38081,N_38323);
nor U38763 (N_38763,N_38108,N_38386);
and U38764 (N_38764,N_38097,N_38373);
nand U38765 (N_38765,N_38053,N_38141);
nor U38766 (N_38766,N_38427,N_38465);
or U38767 (N_38767,N_38212,N_38387);
or U38768 (N_38768,N_38106,N_38406);
nor U38769 (N_38769,N_38382,N_38373);
nor U38770 (N_38770,N_38017,N_38386);
nand U38771 (N_38771,N_38412,N_38107);
xor U38772 (N_38772,N_38471,N_38317);
nand U38773 (N_38773,N_38078,N_38417);
nand U38774 (N_38774,N_38408,N_38026);
or U38775 (N_38775,N_38322,N_38078);
nor U38776 (N_38776,N_38367,N_38252);
or U38777 (N_38777,N_38068,N_38278);
or U38778 (N_38778,N_38368,N_38310);
and U38779 (N_38779,N_38056,N_38093);
nand U38780 (N_38780,N_38382,N_38292);
xor U38781 (N_38781,N_38441,N_38185);
or U38782 (N_38782,N_38262,N_38135);
and U38783 (N_38783,N_38181,N_38398);
and U38784 (N_38784,N_38152,N_38359);
and U38785 (N_38785,N_38141,N_38210);
and U38786 (N_38786,N_38157,N_38387);
nor U38787 (N_38787,N_38318,N_38052);
nand U38788 (N_38788,N_38337,N_38284);
nand U38789 (N_38789,N_38472,N_38096);
nor U38790 (N_38790,N_38153,N_38385);
nor U38791 (N_38791,N_38299,N_38459);
or U38792 (N_38792,N_38212,N_38014);
nor U38793 (N_38793,N_38091,N_38451);
and U38794 (N_38794,N_38251,N_38157);
or U38795 (N_38795,N_38487,N_38230);
xor U38796 (N_38796,N_38180,N_38061);
xor U38797 (N_38797,N_38162,N_38265);
nand U38798 (N_38798,N_38033,N_38082);
xor U38799 (N_38799,N_38169,N_38448);
nand U38800 (N_38800,N_38130,N_38457);
or U38801 (N_38801,N_38454,N_38414);
xor U38802 (N_38802,N_38275,N_38303);
or U38803 (N_38803,N_38464,N_38007);
and U38804 (N_38804,N_38070,N_38109);
nand U38805 (N_38805,N_38209,N_38062);
xor U38806 (N_38806,N_38480,N_38436);
nor U38807 (N_38807,N_38430,N_38288);
or U38808 (N_38808,N_38473,N_38149);
nand U38809 (N_38809,N_38479,N_38417);
and U38810 (N_38810,N_38247,N_38388);
nand U38811 (N_38811,N_38267,N_38215);
nor U38812 (N_38812,N_38181,N_38413);
and U38813 (N_38813,N_38437,N_38008);
or U38814 (N_38814,N_38390,N_38243);
xor U38815 (N_38815,N_38117,N_38299);
nor U38816 (N_38816,N_38435,N_38100);
nor U38817 (N_38817,N_38033,N_38477);
nor U38818 (N_38818,N_38022,N_38031);
xor U38819 (N_38819,N_38026,N_38031);
and U38820 (N_38820,N_38162,N_38136);
xor U38821 (N_38821,N_38346,N_38489);
xnor U38822 (N_38822,N_38166,N_38424);
or U38823 (N_38823,N_38226,N_38325);
and U38824 (N_38824,N_38152,N_38215);
xnor U38825 (N_38825,N_38314,N_38372);
and U38826 (N_38826,N_38279,N_38417);
xnor U38827 (N_38827,N_38219,N_38308);
nor U38828 (N_38828,N_38038,N_38379);
or U38829 (N_38829,N_38323,N_38420);
nor U38830 (N_38830,N_38131,N_38425);
nand U38831 (N_38831,N_38071,N_38020);
xnor U38832 (N_38832,N_38366,N_38213);
nand U38833 (N_38833,N_38113,N_38483);
nor U38834 (N_38834,N_38308,N_38395);
or U38835 (N_38835,N_38160,N_38284);
nand U38836 (N_38836,N_38414,N_38262);
and U38837 (N_38837,N_38428,N_38124);
nand U38838 (N_38838,N_38064,N_38180);
and U38839 (N_38839,N_38474,N_38286);
xnor U38840 (N_38840,N_38132,N_38347);
xor U38841 (N_38841,N_38177,N_38388);
and U38842 (N_38842,N_38257,N_38434);
xor U38843 (N_38843,N_38415,N_38289);
and U38844 (N_38844,N_38135,N_38201);
nand U38845 (N_38845,N_38382,N_38486);
nand U38846 (N_38846,N_38118,N_38155);
nand U38847 (N_38847,N_38338,N_38481);
nand U38848 (N_38848,N_38440,N_38127);
xor U38849 (N_38849,N_38010,N_38053);
nand U38850 (N_38850,N_38247,N_38047);
and U38851 (N_38851,N_38129,N_38333);
and U38852 (N_38852,N_38471,N_38386);
nand U38853 (N_38853,N_38050,N_38222);
nor U38854 (N_38854,N_38363,N_38472);
or U38855 (N_38855,N_38075,N_38187);
nand U38856 (N_38856,N_38460,N_38480);
or U38857 (N_38857,N_38056,N_38276);
and U38858 (N_38858,N_38293,N_38270);
nand U38859 (N_38859,N_38397,N_38367);
xnor U38860 (N_38860,N_38063,N_38094);
or U38861 (N_38861,N_38408,N_38134);
and U38862 (N_38862,N_38441,N_38140);
nand U38863 (N_38863,N_38427,N_38303);
or U38864 (N_38864,N_38090,N_38020);
nand U38865 (N_38865,N_38173,N_38001);
nor U38866 (N_38866,N_38130,N_38071);
nand U38867 (N_38867,N_38044,N_38299);
xor U38868 (N_38868,N_38066,N_38117);
xor U38869 (N_38869,N_38287,N_38447);
or U38870 (N_38870,N_38100,N_38241);
or U38871 (N_38871,N_38215,N_38384);
nor U38872 (N_38872,N_38453,N_38348);
and U38873 (N_38873,N_38067,N_38328);
and U38874 (N_38874,N_38074,N_38213);
nand U38875 (N_38875,N_38064,N_38085);
or U38876 (N_38876,N_38389,N_38004);
xnor U38877 (N_38877,N_38410,N_38356);
nor U38878 (N_38878,N_38429,N_38171);
xnor U38879 (N_38879,N_38181,N_38268);
and U38880 (N_38880,N_38392,N_38190);
and U38881 (N_38881,N_38400,N_38404);
xnor U38882 (N_38882,N_38267,N_38220);
nor U38883 (N_38883,N_38315,N_38011);
nor U38884 (N_38884,N_38420,N_38002);
nand U38885 (N_38885,N_38148,N_38296);
nor U38886 (N_38886,N_38498,N_38309);
xor U38887 (N_38887,N_38398,N_38392);
nor U38888 (N_38888,N_38293,N_38210);
nand U38889 (N_38889,N_38427,N_38202);
and U38890 (N_38890,N_38428,N_38488);
or U38891 (N_38891,N_38402,N_38439);
or U38892 (N_38892,N_38001,N_38188);
nand U38893 (N_38893,N_38401,N_38321);
and U38894 (N_38894,N_38196,N_38129);
xnor U38895 (N_38895,N_38090,N_38144);
nand U38896 (N_38896,N_38288,N_38361);
and U38897 (N_38897,N_38114,N_38225);
nand U38898 (N_38898,N_38243,N_38240);
xnor U38899 (N_38899,N_38458,N_38230);
nand U38900 (N_38900,N_38371,N_38153);
xnor U38901 (N_38901,N_38319,N_38499);
nor U38902 (N_38902,N_38216,N_38294);
xor U38903 (N_38903,N_38267,N_38321);
or U38904 (N_38904,N_38093,N_38222);
nor U38905 (N_38905,N_38013,N_38335);
xor U38906 (N_38906,N_38021,N_38026);
xnor U38907 (N_38907,N_38269,N_38442);
and U38908 (N_38908,N_38162,N_38010);
nor U38909 (N_38909,N_38161,N_38430);
or U38910 (N_38910,N_38129,N_38338);
nand U38911 (N_38911,N_38370,N_38079);
nor U38912 (N_38912,N_38118,N_38100);
or U38913 (N_38913,N_38394,N_38179);
xnor U38914 (N_38914,N_38450,N_38286);
or U38915 (N_38915,N_38238,N_38301);
xnor U38916 (N_38916,N_38289,N_38429);
nand U38917 (N_38917,N_38374,N_38255);
or U38918 (N_38918,N_38431,N_38203);
nor U38919 (N_38919,N_38235,N_38410);
and U38920 (N_38920,N_38001,N_38165);
nor U38921 (N_38921,N_38297,N_38136);
and U38922 (N_38922,N_38115,N_38104);
or U38923 (N_38923,N_38259,N_38234);
nor U38924 (N_38924,N_38289,N_38241);
xor U38925 (N_38925,N_38167,N_38141);
nor U38926 (N_38926,N_38084,N_38070);
xor U38927 (N_38927,N_38162,N_38398);
and U38928 (N_38928,N_38457,N_38458);
and U38929 (N_38929,N_38284,N_38328);
xnor U38930 (N_38930,N_38459,N_38251);
nand U38931 (N_38931,N_38114,N_38125);
and U38932 (N_38932,N_38048,N_38246);
nor U38933 (N_38933,N_38290,N_38279);
xnor U38934 (N_38934,N_38464,N_38252);
or U38935 (N_38935,N_38112,N_38188);
and U38936 (N_38936,N_38347,N_38333);
xnor U38937 (N_38937,N_38316,N_38145);
nand U38938 (N_38938,N_38277,N_38319);
or U38939 (N_38939,N_38184,N_38281);
or U38940 (N_38940,N_38469,N_38269);
or U38941 (N_38941,N_38212,N_38328);
or U38942 (N_38942,N_38437,N_38294);
nand U38943 (N_38943,N_38241,N_38094);
and U38944 (N_38944,N_38394,N_38056);
and U38945 (N_38945,N_38261,N_38162);
xor U38946 (N_38946,N_38480,N_38193);
nand U38947 (N_38947,N_38299,N_38297);
nand U38948 (N_38948,N_38201,N_38357);
and U38949 (N_38949,N_38432,N_38359);
nor U38950 (N_38950,N_38273,N_38218);
nor U38951 (N_38951,N_38482,N_38005);
nor U38952 (N_38952,N_38038,N_38153);
xor U38953 (N_38953,N_38331,N_38300);
xnor U38954 (N_38954,N_38489,N_38172);
nor U38955 (N_38955,N_38387,N_38426);
or U38956 (N_38956,N_38087,N_38446);
xor U38957 (N_38957,N_38415,N_38270);
nor U38958 (N_38958,N_38331,N_38118);
nand U38959 (N_38959,N_38443,N_38093);
nor U38960 (N_38960,N_38420,N_38122);
xnor U38961 (N_38961,N_38438,N_38495);
and U38962 (N_38962,N_38385,N_38476);
and U38963 (N_38963,N_38208,N_38364);
nor U38964 (N_38964,N_38121,N_38249);
nand U38965 (N_38965,N_38063,N_38309);
xor U38966 (N_38966,N_38029,N_38305);
nand U38967 (N_38967,N_38317,N_38003);
nor U38968 (N_38968,N_38151,N_38092);
xor U38969 (N_38969,N_38290,N_38064);
nor U38970 (N_38970,N_38192,N_38413);
and U38971 (N_38971,N_38318,N_38332);
xor U38972 (N_38972,N_38453,N_38369);
and U38973 (N_38973,N_38059,N_38490);
or U38974 (N_38974,N_38155,N_38472);
nand U38975 (N_38975,N_38351,N_38155);
nor U38976 (N_38976,N_38456,N_38197);
or U38977 (N_38977,N_38340,N_38069);
xnor U38978 (N_38978,N_38107,N_38013);
or U38979 (N_38979,N_38417,N_38242);
nor U38980 (N_38980,N_38024,N_38211);
or U38981 (N_38981,N_38073,N_38275);
or U38982 (N_38982,N_38228,N_38318);
or U38983 (N_38983,N_38215,N_38377);
or U38984 (N_38984,N_38447,N_38483);
xnor U38985 (N_38985,N_38253,N_38021);
nand U38986 (N_38986,N_38317,N_38203);
xor U38987 (N_38987,N_38141,N_38414);
xor U38988 (N_38988,N_38251,N_38103);
xor U38989 (N_38989,N_38188,N_38430);
or U38990 (N_38990,N_38152,N_38146);
nor U38991 (N_38991,N_38381,N_38475);
and U38992 (N_38992,N_38201,N_38129);
and U38993 (N_38993,N_38380,N_38354);
xor U38994 (N_38994,N_38231,N_38071);
nand U38995 (N_38995,N_38103,N_38152);
nand U38996 (N_38996,N_38050,N_38140);
and U38997 (N_38997,N_38142,N_38470);
or U38998 (N_38998,N_38203,N_38424);
nor U38999 (N_38999,N_38359,N_38263);
or U39000 (N_39000,N_38928,N_38844);
nor U39001 (N_39001,N_38957,N_38505);
xnor U39002 (N_39002,N_38801,N_38823);
nor U39003 (N_39003,N_38591,N_38831);
xnor U39004 (N_39004,N_38767,N_38960);
xor U39005 (N_39005,N_38795,N_38619);
or U39006 (N_39006,N_38506,N_38908);
and U39007 (N_39007,N_38738,N_38569);
and U39008 (N_39008,N_38897,N_38710);
nand U39009 (N_39009,N_38907,N_38624);
and U39010 (N_39010,N_38816,N_38670);
nor U39011 (N_39011,N_38627,N_38990);
and U39012 (N_39012,N_38744,N_38768);
xor U39013 (N_39013,N_38789,N_38980);
xnor U39014 (N_39014,N_38708,N_38514);
and U39015 (N_39015,N_38689,N_38838);
and U39016 (N_39016,N_38618,N_38771);
or U39017 (N_39017,N_38631,N_38724);
xor U39018 (N_39018,N_38994,N_38553);
and U39019 (N_39019,N_38582,N_38676);
nor U39020 (N_39020,N_38938,N_38589);
or U39021 (N_39021,N_38750,N_38502);
nor U39022 (N_39022,N_38895,N_38829);
xor U39023 (N_39023,N_38544,N_38772);
xor U39024 (N_39024,N_38586,N_38934);
nand U39025 (N_39025,N_38731,N_38892);
nand U39026 (N_39026,N_38828,N_38715);
xor U39027 (N_39027,N_38688,N_38930);
nor U39028 (N_39028,N_38728,N_38597);
nor U39029 (N_39029,N_38570,N_38786);
nand U39030 (N_39030,N_38763,N_38971);
and U39031 (N_39031,N_38882,N_38920);
xnor U39032 (N_39032,N_38626,N_38848);
or U39033 (N_39033,N_38587,N_38565);
nand U39034 (N_39034,N_38739,N_38593);
nor U39035 (N_39035,N_38655,N_38966);
and U39036 (N_39036,N_38691,N_38923);
nor U39037 (N_39037,N_38600,N_38913);
nor U39038 (N_39038,N_38769,N_38953);
nor U39039 (N_39039,N_38815,N_38975);
nor U39040 (N_39040,N_38775,N_38555);
and U39041 (N_39041,N_38515,N_38543);
and U39042 (N_39042,N_38978,N_38947);
or U39043 (N_39043,N_38699,N_38945);
xnor U39044 (N_39044,N_38664,N_38770);
nor U39045 (N_39045,N_38940,N_38900);
xor U39046 (N_39046,N_38937,N_38893);
and U39047 (N_39047,N_38636,N_38736);
nor U39048 (N_39048,N_38509,N_38683);
and U39049 (N_39049,N_38722,N_38566);
and U39050 (N_39050,N_38981,N_38824);
and U39051 (N_39051,N_38922,N_38813);
nor U39052 (N_39052,N_38573,N_38564);
xor U39053 (N_39053,N_38554,N_38741);
nand U39054 (N_39054,N_38927,N_38579);
nor U39055 (N_39055,N_38692,N_38518);
or U39056 (N_39056,N_38610,N_38756);
nand U39057 (N_39057,N_38754,N_38899);
and U39058 (N_39058,N_38866,N_38915);
and U39059 (N_39059,N_38718,N_38791);
nand U39060 (N_39060,N_38540,N_38519);
nor U39061 (N_39061,N_38865,N_38825);
and U39062 (N_39062,N_38864,N_38651);
xor U39063 (N_39063,N_38751,N_38881);
or U39064 (N_39064,N_38721,N_38942);
or U39065 (N_39065,N_38758,N_38808);
xnor U39066 (N_39066,N_38991,N_38997);
and U39067 (N_39067,N_38740,N_38605);
or U39068 (N_39068,N_38842,N_38834);
nand U39069 (N_39069,N_38604,N_38603);
or U39070 (N_39070,N_38633,N_38711);
nor U39071 (N_39071,N_38964,N_38985);
xnor U39072 (N_39072,N_38525,N_38551);
xnor U39073 (N_39073,N_38870,N_38625);
or U39074 (N_39074,N_38935,N_38986);
nand U39075 (N_39075,N_38561,N_38800);
nand U39076 (N_39076,N_38698,N_38989);
or U39077 (N_39077,N_38617,N_38678);
and U39078 (N_39078,N_38556,N_38716);
or U39079 (N_39079,N_38988,N_38963);
nand U39080 (N_39080,N_38622,N_38863);
xor U39081 (N_39081,N_38837,N_38684);
xnor U39082 (N_39082,N_38941,N_38658);
nand U39083 (N_39083,N_38712,N_38668);
nand U39084 (N_39084,N_38861,N_38950);
xor U39085 (N_39085,N_38512,N_38681);
xor U39086 (N_39086,N_38644,N_38727);
and U39087 (N_39087,N_38694,N_38803);
and U39088 (N_39088,N_38933,N_38675);
xor U39089 (N_39089,N_38919,N_38798);
xor U39090 (N_39090,N_38623,N_38806);
and U39091 (N_39091,N_38890,N_38733);
nor U39092 (N_39092,N_38535,N_38832);
nor U39093 (N_39093,N_38608,N_38601);
nor U39094 (N_39094,N_38585,N_38542);
xnor U39095 (N_39095,N_38620,N_38883);
xor U39096 (N_39096,N_38993,N_38752);
and U39097 (N_39097,N_38562,N_38807);
or U39098 (N_39098,N_38876,N_38647);
nor U39099 (N_39099,N_38707,N_38958);
nand U39100 (N_39100,N_38705,N_38560);
and U39101 (N_39101,N_38507,N_38719);
or U39102 (N_39102,N_38969,N_38677);
xnor U39103 (N_39103,N_38697,N_38590);
nand U39104 (N_39104,N_38547,N_38583);
nand U39105 (N_39105,N_38851,N_38827);
or U39106 (N_39106,N_38745,N_38599);
nor U39107 (N_39107,N_38530,N_38878);
and U39108 (N_39108,N_38634,N_38730);
nor U39109 (N_39109,N_38517,N_38850);
nor U39110 (N_39110,N_38725,N_38536);
nor U39111 (N_39111,N_38999,N_38541);
and U39112 (N_39112,N_38594,N_38679);
nor U39113 (N_39113,N_38792,N_38630);
xnor U39114 (N_39114,N_38615,N_38787);
or U39115 (N_39115,N_38962,N_38672);
and U39116 (N_39116,N_38932,N_38901);
or U39117 (N_39117,N_38819,N_38671);
xnor U39118 (N_39118,N_38797,N_38654);
nand U39119 (N_39119,N_38918,N_38635);
xnor U39120 (N_39120,N_38737,N_38812);
xnor U39121 (N_39121,N_38785,N_38885);
nor U39122 (N_39122,N_38760,N_38793);
xnor U39123 (N_39123,N_38805,N_38898);
nor U39124 (N_39124,N_38952,N_38779);
or U39125 (N_39125,N_38550,N_38529);
xor U39126 (N_39126,N_38916,N_38944);
xor U39127 (N_39127,N_38537,N_38880);
nor U39128 (N_39128,N_38538,N_38977);
xnor U39129 (N_39129,N_38955,N_38926);
and U39130 (N_39130,N_38656,N_38931);
nand U39131 (N_39131,N_38784,N_38503);
nor U39132 (N_39132,N_38743,N_38821);
xor U39133 (N_39133,N_38777,N_38875);
or U39134 (N_39134,N_38528,N_38577);
xnor U39135 (N_39135,N_38735,N_38835);
and U39136 (N_39136,N_38888,N_38765);
nor U39137 (N_39137,N_38889,N_38840);
and U39138 (N_39138,N_38961,N_38500);
nand U39139 (N_39139,N_38841,N_38959);
nand U39140 (N_39140,N_38661,N_38778);
xnor U39141 (N_39141,N_38637,N_38902);
and U39142 (N_39142,N_38584,N_38510);
xor U39143 (N_39143,N_38965,N_38501);
nand U39144 (N_39144,N_38996,N_38896);
nand U39145 (N_39145,N_38749,N_38723);
xor U39146 (N_39146,N_38968,N_38660);
nand U39147 (N_39147,N_38886,N_38817);
or U39148 (N_39148,N_38820,N_38726);
and U39149 (N_39149,N_38979,N_38649);
or U39150 (N_39150,N_38859,N_38527);
or U39151 (N_39151,N_38904,N_38970);
or U39152 (N_39152,N_38917,N_38685);
nor U39153 (N_39153,N_38911,N_38909);
nand U39154 (N_39154,N_38759,N_38845);
and U39155 (N_39155,N_38532,N_38894);
xnor U39156 (N_39156,N_38729,N_38983);
xor U39157 (N_39157,N_38648,N_38954);
nor U39158 (N_39158,N_38906,N_38612);
xor U39159 (N_39159,N_38874,N_38642);
or U39160 (N_39160,N_38891,N_38621);
nor U39161 (N_39161,N_38690,N_38860);
xor U39162 (N_39162,N_38910,N_38967);
nor U39163 (N_39163,N_38905,N_38616);
xnor U39164 (N_39164,N_38869,N_38513);
xnor U39165 (N_39165,N_38575,N_38521);
nor U39166 (N_39166,N_38511,N_38628);
and U39167 (N_39167,N_38984,N_38774);
nand U39168 (N_39168,N_38534,N_38508);
nor U39169 (N_39169,N_38558,N_38696);
nand U39170 (N_39170,N_38666,N_38549);
xnor U39171 (N_39171,N_38973,N_38662);
or U39172 (N_39172,N_38761,N_38526);
xor U39173 (N_39173,N_38833,N_38714);
nand U39174 (N_39174,N_38602,N_38693);
and U39175 (N_39175,N_38706,N_38747);
or U39176 (N_39176,N_38847,N_38790);
xor U39177 (N_39177,N_38814,N_38686);
xor U39178 (N_39178,N_38643,N_38520);
nor U39179 (N_39179,N_38855,N_38734);
or U39180 (N_39180,N_38871,N_38924);
nand U39181 (N_39181,N_38852,N_38946);
xor U39182 (N_39182,N_38703,N_38925);
or U39183 (N_39183,N_38780,N_38929);
xnor U39184 (N_39184,N_38663,N_38887);
or U39185 (N_39185,N_38987,N_38638);
xor U39186 (N_39186,N_38516,N_38879);
nor U39187 (N_39187,N_38559,N_38856);
nor U39188 (N_39188,N_38802,N_38606);
and U39189 (N_39189,N_38552,N_38742);
nand U39190 (N_39190,N_38588,N_38571);
nor U39191 (N_39191,N_38781,N_38748);
nand U39192 (N_39192,N_38794,N_38609);
nor U39193 (N_39193,N_38607,N_38545);
nor U39194 (N_39194,N_38854,N_38598);
or U39195 (N_39195,N_38653,N_38667);
nor U39196 (N_39196,N_38581,N_38868);
or U39197 (N_39197,N_38641,N_38921);
xor U39198 (N_39198,N_38843,N_38611);
nand U39199 (N_39199,N_38873,N_38914);
or U39200 (N_39200,N_38912,N_38673);
xor U39201 (N_39201,N_38523,N_38773);
nand U39202 (N_39202,N_38949,N_38563);
xnor U39203 (N_39203,N_38657,N_38939);
and U39204 (N_39204,N_38640,N_38755);
nor U39205 (N_39205,N_38700,N_38809);
and U39206 (N_39206,N_38646,N_38717);
nor U39207 (N_39207,N_38783,N_38596);
nand U39208 (N_39208,N_38867,N_38639);
nor U39209 (N_39209,N_38504,N_38974);
and U39210 (N_39210,N_38862,N_38982);
nand U39211 (N_39211,N_38546,N_38872);
and U39212 (N_39212,N_38595,N_38674);
and U39213 (N_39213,N_38522,N_38757);
nor U39214 (N_39214,N_38614,N_38613);
xor U39215 (N_39215,N_38695,N_38548);
xnor U39216 (N_39216,N_38948,N_38704);
xor U39217 (N_39217,N_38857,N_38574);
nand U39218 (N_39218,N_38884,N_38669);
nor U39219 (N_39219,N_38645,N_38766);
nor U39220 (N_39220,N_38652,N_38632);
and U39221 (N_39221,N_38804,N_38903);
nor U39222 (N_39222,N_38998,N_38702);
and U39223 (N_39223,N_38682,N_38956);
or U39224 (N_39224,N_38972,N_38858);
or U39225 (N_39225,N_38687,N_38951);
or U39226 (N_39226,N_38568,N_38531);
nand U39227 (N_39227,N_38796,N_38753);
nor U39228 (N_39228,N_38680,N_38830);
and U39229 (N_39229,N_38746,N_38853);
xnor U39230 (N_39230,N_38557,N_38818);
xnor U39231 (N_39231,N_38788,N_38592);
or U39232 (N_39232,N_38762,N_38839);
xor U39233 (N_39233,N_38578,N_38580);
xor U39234 (N_39234,N_38764,N_38836);
nor U39235 (N_39235,N_38846,N_38811);
nand U39236 (N_39236,N_38720,N_38877);
nand U39237 (N_39237,N_38782,N_38799);
nor U39238 (N_39238,N_38665,N_38539);
or U39239 (N_39239,N_38576,N_38849);
nor U39240 (N_39240,N_38629,N_38533);
nand U39241 (N_39241,N_38713,N_38650);
nor U39242 (N_39242,N_38659,N_38822);
nor U39243 (N_39243,N_38936,N_38567);
xnor U39244 (N_39244,N_38572,N_38776);
or U39245 (N_39245,N_38524,N_38709);
xor U39246 (N_39246,N_38732,N_38701);
nor U39247 (N_39247,N_38976,N_38992);
or U39248 (N_39248,N_38810,N_38826);
nor U39249 (N_39249,N_38995,N_38943);
or U39250 (N_39250,N_38592,N_38881);
nand U39251 (N_39251,N_38593,N_38859);
and U39252 (N_39252,N_38921,N_38560);
nor U39253 (N_39253,N_38853,N_38703);
nor U39254 (N_39254,N_38564,N_38986);
or U39255 (N_39255,N_38783,N_38802);
and U39256 (N_39256,N_38640,N_38871);
xor U39257 (N_39257,N_38702,N_38502);
nor U39258 (N_39258,N_38884,N_38695);
nor U39259 (N_39259,N_38790,N_38752);
xor U39260 (N_39260,N_38625,N_38939);
nor U39261 (N_39261,N_38745,N_38758);
xnor U39262 (N_39262,N_38590,N_38513);
or U39263 (N_39263,N_38541,N_38507);
nand U39264 (N_39264,N_38738,N_38870);
xor U39265 (N_39265,N_38689,N_38704);
and U39266 (N_39266,N_38801,N_38953);
nor U39267 (N_39267,N_38551,N_38812);
xor U39268 (N_39268,N_38964,N_38904);
nand U39269 (N_39269,N_38914,N_38747);
or U39270 (N_39270,N_38763,N_38605);
xnor U39271 (N_39271,N_38835,N_38915);
and U39272 (N_39272,N_38998,N_38962);
or U39273 (N_39273,N_38514,N_38676);
and U39274 (N_39274,N_38664,N_38515);
and U39275 (N_39275,N_38974,N_38900);
and U39276 (N_39276,N_38596,N_38603);
xor U39277 (N_39277,N_38737,N_38621);
or U39278 (N_39278,N_38708,N_38987);
and U39279 (N_39279,N_38596,N_38920);
nand U39280 (N_39280,N_38882,N_38859);
nand U39281 (N_39281,N_38593,N_38926);
xor U39282 (N_39282,N_38919,N_38580);
and U39283 (N_39283,N_38626,N_38992);
and U39284 (N_39284,N_38919,N_38753);
nor U39285 (N_39285,N_38727,N_38753);
nand U39286 (N_39286,N_38744,N_38570);
nand U39287 (N_39287,N_38874,N_38737);
nand U39288 (N_39288,N_38707,N_38919);
and U39289 (N_39289,N_38887,N_38906);
and U39290 (N_39290,N_38556,N_38607);
and U39291 (N_39291,N_38907,N_38529);
and U39292 (N_39292,N_38917,N_38865);
xor U39293 (N_39293,N_38852,N_38571);
or U39294 (N_39294,N_38524,N_38732);
or U39295 (N_39295,N_38688,N_38532);
nand U39296 (N_39296,N_38680,N_38625);
or U39297 (N_39297,N_38601,N_38906);
and U39298 (N_39298,N_38822,N_38683);
xor U39299 (N_39299,N_38848,N_38634);
nand U39300 (N_39300,N_38670,N_38599);
xor U39301 (N_39301,N_38745,N_38828);
and U39302 (N_39302,N_38534,N_38593);
xnor U39303 (N_39303,N_38912,N_38777);
or U39304 (N_39304,N_38574,N_38809);
or U39305 (N_39305,N_38760,N_38986);
nor U39306 (N_39306,N_38566,N_38843);
nor U39307 (N_39307,N_38814,N_38867);
nand U39308 (N_39308,N_38811,N_38776);
or U39309 (N_39309,N_38862,N_38514);
nand U39310 (N_39310,N_38530,N_38918);
xor U39311 (N_39311,N_38667,N_38946);
or U39312 (N_39312,N_38527,N_38921);
nor U39313 (N_39313,N_38545,N_38629);
xor U39314 (N_39314,N_38899,N_38624);
or U39315 (N_39315,N_38834,N_38818);
xor U39316 (N_39316,N_38673,N_38896);
nor U39317 (N_39317,N_38802,N_38666);
nand U39318 (N_39318,N_38728,N_38834);
nand U39319 (N_39319,N_38918,N_38746);
nor U39320 (N_39320,N_38996,N_38629);
nand U39321 (N_39321,N_38985,N_38734);
xor U39322 (N_39322,N_38892,N_38695);
or U39323 (N_39323,N_38554,N_38719);
nand U39324 (N_39324,N_38993,N_38584);
xor U39325 (N_39325,N_38983,N_38957);
nand U39326 (N_39326,N_38914,N_38814);
or U39327 (N_39327,N_38798,N_38523);
nand U39328 (N_39328,N_38528,N_38616);
xnor U39329 (N_39329,N_38660,N_38900);
xor U39330 (N_39330,N_38841,N_38862);
xnor U39331 (N_39331,N_38662,N_38573);
or U39332 (N_39332,N_38934,N_38549);
and U39333 (N_39333,N_38885,N_38603);
or U39334 (N_39334,N_38672,N_38633);
nand U39335 (N_39335,N_38967,N_38546);
nor U39336 (N_39336,N_38718,N_38587);
nor U39337 (N_39337,N_38781,N_38589);
or U39338 (N_39338,N_38961,N_38601);
or U39339 (N_39339,N_38668,N_38991);
nor U39340 (N_39340,N_38846,N_38699);
or U39341 (N_39341,N_38581,N_38923);
and U39342 (N_39342,N_38541,N_38603);
nand U39343 (N_39343,N_38588,N_38887);
and U39344 (N_39344,N_38975,N_38902);
or U39345 (N_39345,N_38504,N_38828);
nand U39346 (N_39346,N_38610,N_38710);
nand U39347 (N_39347,N_38639,N_38657);
nand U39348 (N_39348,N_38553,N_38572);
nor U39349 (N_39349,N_38767,N_38844);
and U39350 (N_39350,N_38985,N_38991);
nand U39351 (N_39351,N_38990,N_38599);
xnor U39352 (N_39352,N_38955,N_38552);
or U39353 (N_39353,N_38922,N_38893);
or U39354 (N_39354,N_38791,N_38729);
nor U39355 (N_39355,N_38736,N_38750);
nor U39356 (N_39356,N_38666,N_38805);
xor U39357 (N_39357,N_38607,N_38655);
nand U39358 (N_39358,N_38717,N_38997);
nor U39359 (N_39359,N_38906,N_38602);
nor U39360 (N_39360,N_38581,N_38517);
and U39361 (N_39361,N_38971,N_38959);
nor U39362 (N_39362,N_38509,N_38759);
nand U39363 (N_39363,N_38981,N_38909);
and U39364 (N_39364,N_38879,N_38637);
nand U39365 (N_39365,N_38976,N_38749);
and U39366 (N_39366,N_38763,N_38698);
xnor U39367 (N_39367,N_38913,N_38540);
and U39368 (N_39368,N_38759,N_38967);
xor U39369 (N_39369,N_38971,N_38673);
xor U39370 (N_39370,N_38807,N_38701);
xor U39371 (N_39371,N_38640,N_38973);
nor U39372 (N_39372,N_38974,N_38957);
and U39373 (N_39373,N_38546,N_38827);
or U39374 (N_39374,N_38903,N_38736);
or U39375 (N_39375,N_38918,N_38640);
nor U39376 (N_39376,N_38818,N_38964);
nand U39377 (N_39377,N_38514,N_38829);
nor U39378 (N_39378,N_38733,N_38886);
nor U39379 (N_39379,N_38641,N_38797);
or U39380 (N_39380,N_38911,N_38662);
or U39381 (N_39381,N_38899,N_38914);
and U39382 (N_39382,N_38892,N_38516);
and U39383 (N_39383,N_38547,N_38788);
or U39384 (N_39384,N_38626,N_38961);
nor U39385 (N_39385,N_38636,N_38961);
xnor U39386 (N_39386,N_38918,N_38576);
nor U39387 (N_39387,N_38840,N_38725);
or U39388 (N_39388,N_38647,N_38680);
nand U39389 (N_39389,N_38692,N_38561);
and U39390 (N_39390,N_38614,N_38668);
nor U39391 (N_39391,N_38843,N_38669);
nand U39392 (N_39392,N_38585,N_38667);
xor U39393 (N_39393,N_38812,N_38870);
nand U39394 (N_39394,N_38706,N_38764);
nor U39395 (N_39395,N_38997,N_38900);
or U39396 (N_39396,N_38730,N_38727);
or U39397 (N_39397,N_38826,N_38583);
and U39398 (N_39398,N_38726,N_38511);
xnor U39399 (N_39399,N_38770,N_38702);
nor U39400 (N_39400,N_38836,N_38610);
xnor U39401 (N_39401,N_38963,N_38955);
and U39402 (N_39402,N_38529,N_38815);
or U39403 (N_39403,N_38769,N_38896);
nand U39404 (N_39404,N_38729,N_38780);
nand U39405 (N_39405,N_38987,N_38581);
nor U39406 (N_39406,N_38568,N_38923);
nor U39407 (N_39407,N_38515,N_38542);
or U39408 (N_39408,N_38648,N_38959);
and U39409 (N_39409,N_38659,N_38572);
or U39410 (N_39410,N_38756,N_38977);
nor U39411 (N_39411,N_38726,N_38649);
or U39412 (N_39412,N_38625,N_38531);
and U39413 (N_39413,N_38906,N_38890);
and U39414 (N_39414,N_38716,N_38631);
nor U39415 (N_39415,N_38681,N_38871);
nor U39416 (N_39416,N_38631,N_38882);
nand U39417 (N_39417,N_38656,N_38960);
or U39418 (N_39418,N_38728,N_38577);
nor U39419 (N_39419,N_38798,N_38986);
nor U39420 (N_39420,N_38952,N_38913);
or U39421 (N_39421,N_38792,N_38782);
or U39422 (N_39422,N_38734,N_38942);
or U39423 (N_39423,N_38791,N_38615);
or U39424 (N_39424,N_38986,N_38776);
nor U39425 (N_39425,N_38955,N_38715);
xor U39426 (N_39426,N_38657,N_38917);
or U39427 (N_39427,N_38536,N_38661);
xor U39428 (N_39428,N_38627,N_38966);
xnor U39429 (N_39429,N_38873,N_38769);
xnor U39430 (N_39430,N_38696,N_38848);
and U39431 (N_39431,N_38990,N_38840);
or U39432 (N_39432,N_38973,N_38835);
and U39433 (N_39433,N_38908,N_38964);
or U39434 (N_39434,N_38726,N_38532);
or U39435 (N_39435,N_38957,N_38788);
xnor U39436 (N_39436,N_38975,N_38623);
xnor U39437 (N_39437,N_38547,N_38656);
nor U39438 (N_39438,N_38992,N_38541);
nand U39439 (N_39439,N_38826,N_38608);
nand U39440 (N_39440,N_38869,N_38734);
or U39441 (N_39441,N_38796,N_38959);
or U39442 (N_39442,N_38590,N_38879);
or U39443 (N_39443,N_38916,N_38752);
nand U39444 (N_39444,N_38776,N_38602);
xnor U39445 (N_39445,N_38750,N_38529);
or U39446 (N_39446,N_38529,N_38629);
or U39447 (N_39447,N_38923,N_38513);
or U39448 (N_39448,N_38956,N_38711);
xnor U39449 (N_39449,N_38654,N_38816);
and U39450 (N_39450,N_38990,N_38964);
xor U39451 (N_39451,N_38959,N_38715);
nor U39452 (N_39452,N_38817,N_38877);
nand U39453 (N_39453,N_38534,N_38661);
xnor U39454 (N_39454,N_38913,N_38681);
or U39455 (N_39455,N_38869,N_38720);
nor U39456 (N_39456,N_38629,N_38574);
nand U39457 (N_39457,N_38921,N_38509);
nand U39458 (N_39458,N_38591,N_38668);
nand U39459 (N_39459,N_38634,N_38545);
nor U39460 (N_39460,N_38570,N_38730);
and U39461 (N_39461,N_38584,N_38805);
nor U39462 (N_39462,N_38900,N_38700);
nand U39463 (N_39463,N_38510,N_38778);
xnor U39464 (N_39464,N_38657,N_38580);
xor U39465 (N_39465,N_38788,N_38559);
or U39466 (N_39466,N_38618,N_38564);
xnor U39467 (N_39467,N_38759,N_38930);
xor U39468 (N_39468,N_38842,N_38723);
nand U39469 (N_39469,N_38830,N_38958);
or U39470 (N_39470,N_38544,N_38942);
nand U39471 (N_39471,N_38752,N_38624);
xor U39472 (N_39472,N_38729,N_38866);
or U39473 (N_39473,N_38927,N_38765);
and U39474 (N_39474,N_38746,N_38609);
nand U39475 (N_39475,N_38573,N_38884);
xnor U39476 (N_39476,N_38629,N_38897);
or U39477 (N_39477,N_38888,N_38539);
nand U39478 (N_39478,N_38505,N_38567);
and U39479 (N_39479,N_38765,N_38664);
xor U39480 (N_39480,N_38897,N_38973);
xor U39481 (N_39481,N_38939,N_38922);
xor U39482 (N_39482,N_38678,N_38790);
xor U39483 (N_39483,N_38547,N_38640);
or U39484 (N_39484,N_38709,N_38796);
nor U39485 (N_39485,N_38875,N_38745);
xnor U39486 (N_39486,N_38989,N_38622);
xor U39487 (N_39487,N_38791,N_38595);
or U39488 (N_39488,N_38754,N_38974);
nand U39489 (N_39489,N_38563,N_38553);
or U39490 (N_39490,N_38604,N_38537);
nand U39491 (N_39491,N_38806,N_38519);
xor U39492 (N_39492,N_38817,N_38718);
nand U39493 (N_39493,N_38602,N_38505);
or U39494 (N_39494,N_38555,N_38701);
nor U39495 (N_39495,N_38854,N_38743);
and U39496 (N_39496,N_38647,N_38511);
and U39497 (N_39497,N_38651,N_38816);
or U39498 (N_39498,N_38731,N_38841);
nor U39499 (N_39499,N_38639,N_38646);
or U39500 (N_39500,N_39441,N_39424);
nand U39501 (N_39501,N_39497,N_39064);
and U39502 (N_39502,N_39013,N_39232);
and U39503 (N_39503,N_39173,N_39422);
or U39504 (N_39504,N_39371,N_39140);
nor U39505 (N_39505,N_39162,N_39434);
xnor U39506 (N_39506,N_39458,N_39443);
xnor U39507 (N_39507,N_39100,N_39348);
and U39508 (N_39508,N_39143,N_39386);
xnor U39509 (N_39509,N_39242,N_39224);
nor U39510 (N_39510,N_39350,N_39022);
and U39511 (N_39511,N_39270,N_39264);
nand U39512 (N_39512,N_39410,N_39156);
or U39513 (N_39513,N_39356,N_39402);
or U39514 (N_39514,N_39090,N_39414);
xor U39515 (N_39515,N_39228,N_39212);
nor U39516 (N_39516,N_39210,N_39052);
nor U39517 (N_39517,N_39225,N_39235);
or U39518 (N_39518,N_39428,N_39080);
nand U39519 (N_39519,N_39044,N_39359);
nand U39520 (N_39520,N_39248,N_39189);
or U39521 (N_39521,N_39184,N_39439);
xor U39522 (N_39522,N_39020,N_39385);
xor U39523 (N_39523,N_39009,N_39286);
or U39524 (N_39524,N_39318,N_39357);
xor U39525 (N_39525,N_39055,N_39272);
xor U39526 (N_39526,N_39281,N_39244);
and U39527 (N_39527,N_39153,N_39499);
nand U39528 (N_39528,N_39099,N_39193);
xnor U39529 (N_39529,N_39250,N_39398);
nor U39530 (N_39530,N_39030,N_39132);
nor U39531 (N_39531,N_39086,N_39262);
or U39532 (N_39532,N_39331,N_39365);
xor U39533 (N_39533,N_39310,N_39074);
and U39534 (N_39534,N_39484,N_39457);
or U39535 (N_39535,N_39034,N_39195);
nand U39536 (N_39536,N_39444,N_39130);
nand U39537 (N_39537,N_39368,N_39054);
nand U39538 (N_39538,N_39245,N_39101);
or U39539 (N_39539,N_39289,N_39008);
nand U39540 (N_39540,N_39349,N_39107);
nor U39541 (N_39541,N_39389,N_39121);
xnor U39542 (N_39542,N_39294,N_39141);
xor U39543 (N_39543,N_39026,N_39023);
xor U39544 (N_39544,N_39291,N_39137);
or U39545 (N_39545,N_39450,N_39072);
and U39546 (N_39546,N_39406,N_39154);
nand U39547 (N_39547,N_39133,N_39394);
xnor U39548 (N_39548,N_39115,N_39255);
nor U39549 (N_39549,N_39062,N_39351);
nor U39550 (N_39550,N_39098,N_39461);
or U39551 (N_39551,N_39078,N_39126);
nor U39552 (N_39552,N_39185,N_39113);
nor U39553 (N_39553,N_39324,N_39307);
xor U39554 (N_39554,N_39222,N_39011);
nand U39555 (N_39555,N_39227,N_39215);
xor U39556 (N_39556,N_39373,N_39199);
or U39557 (N_39557,N_39313,N_39489);
nand U39558 (N_39558,N_39437,N_39093);
nor U39559 (N_39559,N_39241,N_39483);
nand U39560 (N_39560,N_39000,N_39150);
or U39561 (N_39561,N_39495,N_39338);
or U39562 (N_39562,N_39071,N_39257);
and U39563 (N_39563,N_39089,N_39380);
xnor U39564 (N_39564,N_39178,N_39165);
xnor U39565 (N_39565,N_39298,N_39271);
nand U39566 (N_39566,N_39267,N_39025);
or U39567 (N_39567,N_39112,N_39278);
nor U39568 (N_39568,N_39122,N_39019);
and U39569 (N_39569,N_39149,N_39092);
and U39570 (N_39570,N_39181,N_39363);
nand U39571 (N_39571,N_39028,N_39367);
and U39572 (N_39572,N_39161,N_39436);
xnor U39573 (N_39573,N_39430,N_39075);
and U39574 (N_39574,N_39105,N_39172);
nor U39575 (N_39575,N_39218,N_39216);
nand U39576 (N_39576,N_39312,N_39076);
xor U39577 (N_39577,N_39183,N_39079);
and U39578 (N_39578,N_39304,N_39236);
nor U39579 (N_39579,N_39038,N_39413);
or U39580 (N_39580,N_39012,N_39401);
nor U39581 (N_39581,N_39192,N_39411);
xor U39582 (N_39582,N_39306,N_39238);
and U39583 (N_39583,N_39087,N_39277);
or U39584 (N_39584,N_39360,N_39016);
xnor U39585 (N_39585,N_39015,N_39301);
xor U39586 (N_39586,N_39221,N_39332);
xnor U39587 (N_39587,N_39040,N_39207);
xor U39588 (N_39588,N_39491,N_39382);
xor U39589 (N_39589,N_39418,N_39314);
and U39590 (N_39590,N_39104,N_39018);
or U39591 (N_39591,N_39202,N_39326);
nor U39592 (N_39592,N_39471,N_39152);
and U39593 (N_39593,N_39157,N_39120);
and U39594 (N_39594,N_39010,N_39472);
xor U39595 (N_39595,N_39285,N_39231);
and U39596 (N_39596,N_39396,N_39252);
nor U39597 (N_39597,N_39256,N_39174);
nor U39598 (N_39598,N_39266,N_39213);
or U39599 (N_39599,N_39415,N_39387);
xor U39600 (N_39600,N_39138,N_39223);
nand U39601 (N_39601,N_39493,N_39005);
nor U39602 (N_39602,N_39325,N_39167);
or U39603 (N_39603,N_39136,N_39240);
xor U39604 (N_39604,N_39375,N_39194);
or U39605 (N_39605,N_39377,N_39454);
nand U39606 (N_39606,N_39106,N_39187);
nand U39607 (N_39607,N_39200,N_39408);
and U39608 (N_39608,N_39283,N_39317);
nand U39609 (N_39609,N_39345,N_39473);
nand U39610 (N_39610,N_39036,N_39311);
nand U39611 (N_39611,N_39364,N_39327);
nor U39612 (N_39612,N_39229,N_39391);
nand U39613 (N_39613,N_39094,N_39102);
and U39614 (N_39614,N_39388,N_39209);
nor U39615 (N_39615,N_39147,N_39070);
or U39616 (N_39616,N_39449,N_39372);
and U39617 (N_39617,N_39151,N_39081);
xnor U39618 (N_39618,N_39061,N_39065);
and U39619 (N_39619,N_39417,N_39186);
nand U39620 (N_39620,N_39333,N_39452);
nand U39621 (N_39621,N_39180,N_39467);
or U39622 (N_39622,N_39171,N_39051);
or U39623 (N_39623,N_39407,N_39003);
or U39624 (N_39624,N_39226,N_39247);
nand U39625 (N_39625,N_39427,N_39239);
xor U39626 (N_39626,N_39142,N_39383);
and U39627 (N_39627,N_39487,N_39128);
or U39628 (N_39628,N_39336,N_39399);
and U39629 (N_39629,N_39145,N_39276);
nand U39630 (N_39630,N_39084,N_39343);
nor U39631 (N_39631,N_39297,N_39485);
nor U39632 (N_39632,N_39384,N_39395);
nor U39633 (N_39633,N_39004,N_39303);
nand U39634 (N_39634,N_39131,N_39259);
nand U39635 (N_39635,N_39263,N_39447);
and U39636 (N_39636,N_39230,N_39042);
or U39637 (N_39637,N_39127,N_39056);
or U39638 (N_39638,N_39108,N_39246);
and U39639 (N_39639,N_39296,N_39197);
or U39640 (N_39640,N_39035,N_39279);
and U39641 (N_39641,N_39243,N_39319);
or U39642 (N_39642,N_39159,N_39305);
nor U39643 (N_39643,N_39006,N_39299);
xor U39644 (N_39644,N_39366,N_39091);
and U39645 (N_39645,N_39046,N_39486);
nand U39646 (N_39646,N_39217,N_39021);
nand U39647 (N_39647,N_39329,N_39488);
and U39648 (N_39648,N_39117,N_39435);
nor U39649 (N_39649,N_39456,N_39198);
xnor U39650 (N_39650,N_39166,N_39374);
xor U39651 (N_39651,N_39060,N_39125);
nor U39652 (N_39652,N_39459,N_39322);
nand U39653 (N_39653,N_39433,N_39169);
xor U39654 (N_39654,N_39460,N_39116);
and U39655 (N_39655,N_39290,N_39144);
or U39656 (N_39656,N_39354,N_39423);
or U39657 (N_39657,N_39347,N_39481);
xnor U39658 (N_39658,N_39109,N_39047);
xnor U39659 (N_39659,N_39308,N_39474);
and U39660 (N_39660,N_39369,N_39017);
nand U39661 (N_39661,N_39273,N_39067);
and U39662 (N_39662,N_39158,N_39492);
or U39663 (N_39663,N_39292,N_39249);
xor U39664 (N_39664,N_39479,N_39082);
nor U39665 (N_39665,N_39045,N_39376);
or U39666 (N_39666,N_39111,N_39463);
nor U39667 (N_39667,N_39426,N_39315);
xnor U39668 (N_39668,N_39204,N_39440);
or U39669 (N_39669,N_39465,N_39334);
and U39670 (N_39670,N_39288,N_39177);
xnor U39671 (N_39671,N_39088,N_39103);
or U39672 (N_39672,N_39258,N_39068);
xor U39673 (N_39673,N_39342,N_39274);
xor U39674 (N_39674,N_39182,N_39420);
and U39675 (N_39675,N_39251,N_39265);
nand U39676 (N_39676,N_39269,N_39405);
nor U39677 (N_39677,N_39069,N_39124);
nor U39678 (N_39678,N_39490,N_39059);
and U39679 (N_39679,N_39477,N_39393);
and U39680 (N_39680,N_39470,N_39464);
and U39681 (N_39681,N_39220,N_39438);
and U39682 (N_39682,N_39118,N_39237);
and U39683 (N_39683,N_39341,N_39361);
nand U39684 (N_39684,N_39431,N_39233);
xnor U39685 (N_39685,N_39191,N_39024);
nand U39686 (N_39686,N_39190,N_39451);
and U39687 (N_39687,N_39073,N_39077);
xor U39688 (N_39688,N_39429,N_39164);
xnor U39689 (N_39689,N_39057,N_39032);
xnor U39690 (N_39690,N_39260,N_39063);
or U39691 (N_39691,N_39445,N_39362);
or U39692 (N_39692,N_39287,N_39358);
nand U39693 (N_39693,N_39280,N_39392);
and U39694 (N_39694,N_39001,N_39390);
nor U39695 (N_39695,N_39346,N_39085);
or U39696 (N_39696,N_39275,N_39397);
nand U39697 (N_39697,N_39039,N_39300);
or U39698 (N_39698,N_39400,N_39114);
nand U39699 (N_39699,N_39196,N_39176);
nand U39700 (N_39700,N_39321,N_39494);
nand U39701 (N_39701,N_39442,N_39097);
xor U39702 (N_39702,N_39110,N_39432);
and U39703 (N_39703,N_39482,N_39160);
nand U39704 (N_39704,N_39496,N_39188);
and U39705 (N_39705,N_39353,N_39337);
nand U39706 (N_39706,N_39425,N_39095);
nand U39707 (N_39707,N_39048,N_39119);
xor U39708 (N_39708,N_39293,N_39404);
nand U39709 (N_39709,N_39253,N_39175);
or U39710 (N_39710,N_39049,N_39409);
or U39711 (N_39711,N_39254,N_39146);
or U39712 (N_39712,N_39135,N_39170);
xor U39713 (N_39713,N_39478,N_39448);
nor U39714 (N_39714,N_39352,N_39208);
nand U39715 (N_39715,N_39344,N_39284);
or U39716 (N_39716,N_39309,N_39480);
nand U39717 (N_39717,N_39261,N_39066);
or U39718 (N_39718,N_39211,N_39029);
and U39719 (N_39719,N_39206,N_39498);
and U39720 (N_39720,N_39295,N_39058);
or U39721 (N_39721,N_39053,N_39014);
or U39722 (N_39722,N_39050,N_39002);
nand U39723 (N_39723,N_39219,N_39031);
xnor U39724 (N_39724,N_39370,N_39139);
or U39725 (N_39725,N_39379,N_39340);
nand U39726 (N_39726,N_39041,N_39201);
xor U39727 (N_39727,N_39033,N_39455);
xor U39728 (N_39728,N_39328,N_39421);
nor U39729 (N_39729,N_39037,N_39214);
xnor U39730 (N_39730,N_39419,N_39163);
nor U39731 (N_39731,N_39027,N_39083);
nand U39732 (N_39732,N_39475,N_39282);
xor U39733 (N_39733,N_39203,N_39466);
xnor U39734 (N_39734,N_39330,N_39320);
nor U39735 (N_39735,N_39462,N_39205);
nor U39736 (N_39736,N_39381,N_39446);
or U39737 (N_39737,N_39416,N_39123);
nor U39738 (N_39738,N_39043,N_39335);
nor U39739 (N_39739,N_39468,N_39148);
nor U39740 (N_39740,N_39168,N_39453);
or U39741 (N_39741,N_39155,N_39007);
nor U39742 (N_39742,N_39476,N_39339);
nand U39743 (N_39743,N_39268,N_39323);
or U39744 (N_39744,N_39412,N_39096);
nand U39745 (N_39745,N_39179,N_39403);
xor U39746 (N_39746,N_39316,N_39134);
nor U39747 (N_39747,N_39234,N_39378);
nor U39748 (N_39748,N_39129,N_39469);
and U39749 (N_39749,N_39355,N_39302);
nor U39750 (N_39750,N_39033,N_39293);
nor U39751 (N_39751,N_39274,N_39162);
nand U39752 (N_39752,N_39096,N_39336);
nand U39753 (N_39753,N_39182,N_39303);
xnor U39754 (N_39754,N_39142,N_39153);
nand U39755 (N_39755,N_39106,N_39398);
nor U39756 (N_39756,N_39458,N_39408);
nand U39757 (N_39757,N_39433,N_39012);
nand U39758 (N_39758,N_39066,N_39077);
nor U39759 (N_39759,N_39108,N_39340);
xor U39760 (N_39760,N_39330,N_39221);
nand U39761 (N_39761,N_39434,N_39296);
or U39762 (N_39762,N_39333,N_39090);
nand U39763 (N_39763,N_39031,N_39374);
or U39764 (N_39764,N_39281,N_39330);
nor U39765 (N_39765,N_39389,N_39168);
xnor U39766 (N_39766,N_39199,N_39239);
nor U39767 (N_39767,N_39174,N_39226);
nor U39768 (N_39768,N_39052,N_39492);
nand U39769 (N_39769,N_39462,N_39155);
xor U39770 (N_39770,N_39142,N_39181);
and U39771 (N_39771,N_39079,N_39228);
or U39772 (N_39772,N_39393,N_39419);
nor U39773 (N_39773,N_39059,N_39249);
and U39774 (N_39774,N_39158,N_39437);
nor U39775 (N_39775,N_39212,N_39246);
nor U39776 (N_39776,N_39005,N_39427);
nand U39777 (N_39777,N_39268,N_39257);
or U39778 (N_39778,N_39311,N_39461);
nor U39779 (N_39779,N_39061,N_39370);
xnor U39780 (N_39780,N_39344,N_39309);
or U39781 (N_39781,N_39113,N_39038);
xor U39782 (N_39782,N_39049,N_39251);
or U39783 (N_39783,N_39079,N_39373);
and U39784 (N_39784,N_39003,N_39087);
nand U39785 (N_39785,N_39411,N_39466);
or U39786 (N_39786,N_39425,N_39401);
nor U39787 (N_39787,N_39358,N_39044);
and U39788 (N_39788,N_39288,N_39111);
nor U39789 (N_39789,N_39097,N_39263);
nor U39790 (N_39790,N_39199,N_39279);
or U39791 (N_39791,N_39476,N_39186);
nand U39792 (N_39792,N_39381,N_39012);
nand U39793 (N_39793,N_39228,N_39217);
xor U39794 (N_39794,N_39424,N_39001);
and U39795 (N_39795,N_39251,N_39468);
xor U39796 (N_39796,N_39369,N_39429);
xnor U39797 (N_39797,N_39159,N_39448);
xor U39798 (N_39798,N_39037,N_39002);
nand U39799 (N_39799,N_39429,N_39248);
or U39800 (N_39800,N_39482,N_39156);
nor U39801 (N_39801,N_39061,N_39415);
or U39802 (N_39802,N_39086,N_39372);
nand U39803 (N_39803,N_39487,N_39059);
or U39804 (N_39804,N_39429,N_39288);
nor U39805 (N_39805,N_39322,N_39056);
xor U39806 (N_39806,N_39274,N_39468);
and U39807 (N_39807,N_39263,N_39406);
xor U39808 (N_39808,N_39170,N_39358);
or U39809 (N_39809,N_39350,N_39204);
nor U39810 (N_39810,N_39438,N_39325);
xor U39811 (N_39811,N_39040,N_39427);
or U39812 (N_39812,N_39210,N_39126);
and U39813 (N_39813,N_39057,N_39434);
nor U39814 (N_39814,N_39174,N_39361);
nand U39815 (N_39815,N_39491,N_39085);
or U39816 (N_39816,N_39449,N_39488);
nor U39817 (N_39817,N_39201,N_39316);
nor U39818 (N_39818,N_39117,N_39239);
nor U39819 (N_39819,N_39122,N_39154);
nand U39820 (N_39820,N_39333,N_39113);
nand U39821 (N_39821,N_39480,N_39028);
nand U39822 (N_39822,N_39219,N_39497);
nand U39823 (N_39823,N_39339,N_39107);
or U39824 (N_39824,N_39160,N_39431);
xor U39825 (N_39825,N_39023,N_39161);
and U39826 (N_39826,N_39441,N_39391);
or U39827 (N_39827,N_39022,N_39107);
or U39828 (N_39828,N_39271,N_39418);
nor U39829 (N_39829,N_39068,N_39411);
xor U39830 (N_39830,N_39072,N_39273);
nor U39831 (N_39831,N_39032,N_39308);
nand U39832 (N_39832,N_39279,N_39249);
nand U39833 (N_39833,N_39068,N_39432);
nor U39834 (N_39834,N_39234,N_39482);
nand U39835 (N_39835,N_39154,N_39272);
nor U39836 (N_39836,N_39227,N_39051);
xor U39837 (N_39837,N_39170,N_39371);
or U39838 (N_39838,N_39081,N_39148);
and U39839 (N_39839,N_39094,N_39276);
xor U39840 (N_39840,N_39178,N_39389);
and U39841 (N_39841,N_39293,N_39383);
nand U39842 (N_39842,N_39364,N_39468);
nand U39843 (N_39843,N_39189,N_39291);
xnor U39844 (N_39844,N_39016,N_39056);
or U39845 (N_39845,N_39162,N_39489);
nand U39846 (N_39846,N_39174,N_39486);
xnor U39847 (N_39847,N_39459,N_39324);
nor U39848 (N_39848,N_39372,N_39040);
nor U39849 (N_39849,N_39481,N_39275);
nor U39850 (N_39850,N_39086,N_39388);
nand U39851 (N_39851,N_39358,N_39480);
and U39852 (N_39852,N_39067,N_39245);
nand U39853 (N_39853,N_39133,N_39201);
nor U39854 (N_39854,N_39377,N_39450);
nand U39855 (N_39855,N_39276,N_39084);
or U39856 (N_39856,N_39261,N_39212);
xor U39857 (N_39857,N_39332,N_39107);
or U39858 (N_39858,N_39129,N_39088);
nand U39859 (N_39859,N_39364,N_39356);
xor U39860 (N_39860,N_39429,N_39196);
or U39861 (N_39861,N_39496,N_39465);
nand U39862 (N_39862,N_39108,N_39456);
xnor U39863 (N_39863,N_39049,N_39092);
nand U39864 (N_39864,N_39432,N_39440);
nor U39865 (N_39865,N_39498,N_39459);
xnor U39866 (N_39866,N_39456,N_39243);
or U39867 (N_39867,N_39417,N_39483);
nor U39868 (N_39868,N_39089,N_39096);
and U39869 (N_39869,N_39098,N_39302);
and U39870 (N_39870,N_39370,N_39224);
nand U39871 (N_39871,N_39424,N_39282);
nor U39872 (N_39872,N_39011,N_39021);
and U39873 (N_39873,N_39189,N_39260);
nor U39874 (N_39874,N_39220,N_39275);
nand U39875 (N_39875,N_39395,N_39120);
and U39876 (N_39876,N_39348,N_39347);
nor U39877 (N_39877,N_39329,N_39386);
nor U39878 (N_39878,N_39125,N_39310);
xor U39879 (N_39879,N_39376,N_39371);
xnor U39880 (N_39880,N_39097,N_39130);
xnor U39881 (N_39881,N_39193,N_39058);
nand U39882 (N_39882,N_39088,N_39347);
and U39883 (N_39883,N_39481,N_39147);
nand U39884 (N_39884,N_39333,N_39168);
or U39885 (N_39885,N_39317,N_39027);
and U39886 (N_39886,N_39400,N_39067);
nand U39887 (N_39887,N_39378,N_39228);
or U39888 (N_39888,N_39117,N_39030);
xor U39889 (N_39889,N_39466,N_39422);
and U39890 (N_39890,N_39056,N_39128);
or U39891 (N_39891,N_39008,N_39349);
and U39892 (N_39892,N_39100,N_39165);
nor U39893 (N_39893,N_39322,N_39120);
xnor U39894 (N_39894,N_39364,N_39407);
nand U39895 (N_39895,N_39096,N_39280);
xnor U39896 (N_39896,N_39128,N_39463);
and U39897 (N_39897,N_39482,N_39492);
nand U39898 (N_39898,N_39312,N_39046);
or U39899 (N_39899,N_39210,N_39245);
xnor U39900 (N_39900,N_39010,N_39473);
and U39901 (N_39901,N_39150,N_39450);
nand U39902 (N_39902,N_39425,N_39450);
or U39903 (N_39903,N_39075,N_39127);
xor U39904 (N_39904,N_39110,N_39480);
nand U39905 (N_39905,N_39117,N_39004);
nand U39906 (N_39906,N_39155,N_39048);
nor U39907 (N_39907,N_39033,N_39046);
xor U39908 (N_39908,N_39215,N_39108);
xor U39909 (N_39909,N_39184,N_39316);
and U39910 (N_39910,N_39499,N_39462);
and U39911 (N_39911,N_39303,N_39242);
nand U39912 (N_39912,N_39114,N_39133);
and U39913 (N_39913,N_39192,N_39162);
xnor U39914 (N_39914,N_39382,N_39171);
or U39915 (N_39915,N_39228,N_39151);
nand U39916 (N_39916,N_39086,N_39095);
nand U39917 (N_39917,N_39274,N_39251);
and U39918 (N_39918,N_39094,N_39428);
nor U39919 (N_39919,N_39032,N_39257);
and U39920 (N_39920,N_39395,N_39011);
and U39921 (N_39921,N_39044,N_39179);
xor U39922 (N_39922,N_39050,N_39279);
or U39923 (N_39923,N_39177,N_39483);
or U39924 (N_39924,N_39026,N_39440);
or U39925 (N_39925,N_39403,N_39003);
nor U39926 (N_39926,N_39068,N_39490);
nand U39927 (N_39927,N_39057,N_39491);
or U39928 (N_39928,N_39237,N_39020);
or U39929 (N_39929,N_39425,N_39257);
nor U39930 (N_39930,N_39334,N_39119);
nand U39931 (N_39931,N_39445,N_39442);
and U39932 (N_39932,N_39284,N_39221);
xnor U39933 (N_39933,N_39435,N_39224);
xor U39934 (N_39934,N_39225,N_39275);
xor U39935 (N_39935,N_39099,N_39323);
nor U39936 (N_39936,N_39171,N_39446);
or U39937 (N_39937,N_39288,N_39053);
nor U39938 (N_39938,N_39182,N_39123);
nand U39939 (N_39939,N_39157,N_39116);
nand U39940 (N_39940,N_39132,N_39492);
or U39941 (N_39941,N_39486,N_39363);
or U39942 (N_39942,N_39113,N_39220);
nand U39943 (N_39943,N_39425,N_39260);
nor U39944 (N_39944,N_39447,N_39332);
nor U39945 (N_39945,N_39271,N_39194);
nand U39946 (N_39946,N_39333,N_39233);
nand U39947 (N_39947,N_39200,N_39282);
or U39948 (N_39948,N_39236,N_39177);
xnor U39949 (N_39949,N_39114,N_39136);
nand U39950 (N_39950,N_39389,N_39132);
and U39951 (N_39951,N_39250,N_39139);
or U39952 (N_39952,N_39226,N_39156);
or U39953 (N_39953,N_39181,N_39337);
and U39954 (N_39954,N_39449,N_39096);
nand U39955 (N_39955,N_39041,N_39294);
nor U39956 (N_39956,N_39024,N_39083);
nor U39957 (N_39957,N_39302,N_39074);
or U39958 (N_39958,N_39462,N_39147);
nand U39959 (N_39959,N_39440,N_39453);
or U39960 (N_39960,N_39096,N_39176);
or U39961 (N_39961,N_39432,N_39276);
and U39962 (N_39962,N_39106,N_39165);
nand U39963 (N_39963,N_39113,N_39011);
nor U39964 (N_39964,N_39206,N_39029);
and U39965 (N_39965,N_39210,N_39004);
xor U39966 (N_39966,N_39335,N_39034);
or U39967 (N_39967,N_39204,N_39231);
xnor U39968 (N_39968,N_39388,N_39248);
xnor U39969 (N_39969,N_39165,N_39248);
nor U39970 (N_39970,N_39221,N_39154);
nand U39971 (N_39971,N_39104,N_39334);
nand U39972 (N_39972,N_39249,N_39075);
nor U39973 (N_39973,N_39248,N_39255);
nand U39974 (N_39974,N_39262,N_39173);
nor U39975 (N_39975,N_39451,N_39101);
xnor U39976 (N_39976,N_39496,N_39034);
xnor U39977 (N_39977,N_39291,N_39191);
and U39978 (N_39978,N_39032,N_39262);
nor U39979 (N_39979,N_39254,N_39499);
xor U39980 (N_39980,N_39424,N_39167);
and U39981 (N_39981,N_39202,N_39325);
xor U39982 (N_39982,N_39211,N_39395);
xor U39983 (N_39983,N_39463,N_39060);
and U39984 (N_39984,N_39092,N_39174);
and U39985 (N_39985,N_39128,N_39204);
nand U39986 (N_39986,N_39438,N_39487);
nor U39987 (N_39987,N_39353,N_39469);
and U39988 (N_39988,N_39428,N_39090);
nor U39989 (N_39989,N_39424,N_39461);
nor U39990 (N_39990,N_39275,N_39449);
or U39991 (N_39991,N_39332,N_39093);
nand U39992 (N_39992,N_39390,N_39137);
xor U39993 (N_39993,N_39391,N_39404);
nand U39994 (N_39994,N_39304,N_39300);
nor U39995 (N_39995,N_39031,N_39153);
nand U39996 (N_39996,N_39480,N_39271);
or U39997 (N_39997,N_39447,N_39053);
and U39998 (N_39998,N_39278,N_39243);
and U39999 (N_39999,N_39317,N_39478);
or U40000 (N_40000,N_39664,N_39972);
nor U40001 (N_40001,N_39812,N_39714);
or U40002 (N_40002,N_39640,N_39822);
and U40003 (N_40003,N_39795,N_39775);
or U40004 (N_40004,N_39747,N_39741);
or U40005 (N_40005,N_39927,N_39763);
or U40006 (N_40006,N_39978,N_39666);
and U40007 (N_40007,N_39758,N_39627);
xor U40008 (N_40008,N_39790,N_39751);
or U40009 (N_40009,N_39556,N_39702);
or U40010 (N_40010,N_39860,N_39639);
xnor U40011 (N_40011,N_39936,N_39571);
xnor U40012 (N_40012,N_39574,N_39833);
nand U40013 (N_40013,N_39510,N_39817);
and U40014 (N_40014,N_39944,N_39625);
nand U40015 (N_40015,N_39748,N_39724);
xnor U40016 (N_40016,N_39548,N_39593);
and U40017 (N_40017,N_39622,N_39628);
or U40018 (N_40018,N_39608,N_39695);
xnor U40019 (N_40019,N_39541,N_39513);
xnor U40020 (N_40020,N_39791,N_39709);
nor U40021 (N_40021,N_39713,N_39655);
nand U40022 (N_40022,N_39585,N_39559);
nand U40023 (N_40023,N_39769,N_39965);
or U40024 (N_40024,N_39918,N_39783);
and U40025 (N_40025,N_39850,N_39911);
nand U40026 (N_40026,N_39659,N_39777);
or U40027 (N_40027,N_39813,N_39983);
or U40028 (N_40028,N_39858,N_39715);
nor U40029 (N_40029,N_39598,N_39945);
nor U40030 (N_40030,N_39583,N_39752);
nand U40031 (N_40031,N_39973,N_39700);
nand U40032 (N_40032,N_39685,N_39515);
nand U40033 (N_40033,N_39996,N_39674);
and U40034 (N_40034,N_39867,N_39594);
nand U40035 (N_40035,N_39681,N_39624);
nor U40036 (N_40036,N_39638,N_39810);
xnor U40037 (N_40037,N_39785,N_39566);
and U40038 (N_40038,N_39511,N_39660);
nor U40039 (N_40039,N_39634,N_39756);
xnor U40040 (N_40040,N_39731,N_39919);
or U40041 (N_40041,N_39696,N_39900);
nand U40042 (N_40042,N_39669,N_39917);
nand U40043 (N_40043,N_39505,N_39975);
nand U40044 (N_40044,N_39619,N_39806);
xnor U40045 (N_40045,N_39939,N_39727);
nor U40046 (N_40046,N_39668,N_39636);
nand U40047 (N_40047,N_39932,N_39597);
xor U40048 (N_40048,N_39509,N_39537);
nor U40049 (N_40049,N_39504,N_39542);
or U40050 (N_40050,N_39605,N_39779);
xnor U40051 (N_40051,N_39689,N_39591);
nand U40052 (N_40052,N_39798,N_39652);
or U40053 (N_40053,N_39837,N_39877);
nor U40054 (N_40054,N_39573,N_39831);
nor U40055 (N_40055,N_39637,N_39601);
or U40056 (N_40056,N_39815,N_39930);
or U40057 (N_40057,N_39976,N_39672);
nand U40058 (N_40058,N_39746,N_39768);
or U40059 (N_40059,N_39916,N_39926);
xor U40060 (N_40060,N_39992,N_39550);
or U40061 (N_40061,N_39662,N_39915);
nand U40062 (N_40062,N_39914,N_39921);
nand U40063 (N_40063,N_39698,N_39765);
or U40064 (N_40064,N_39596,N_39892);
and U40065 (N_40065,N_39907,N_39694);
or U40066 (N_40066,N_39502,N_39712);
xnor U40067 (N_40067,N_39545,N_39683);
or U40068 (N_40068,N_39567,N_39909);
xor U40069 (N_40069,N_39611,N_39667);
and U40070 (N_40070,N_39990,N_39985);
xor U40071 (N_40071,N_39897,N_39869);
xnor U40072 (N_40072,N_39552,N_39839);
or U40073 (N_40073,N_39923,N_39863);
xnor U40074 (N_40074,N_39943,N_39687);
nor U40075 (N_40075,N_39508,N_39893);
nor U40076 (N_40076,N_39979,N_39725);
nand U40077 (N_40077,N_39680,N_39635);
nand U40078 (N_40078,N_39692,N_39717);
nor U40079 (N_40079,N_39762,N_39761);
and U40080 (N_40080,N_39631,N_39814);
and U40081 (N_40081,N_39517,N_39564);
nand U40082 (N_40082,N_39739,N_39974);
and U40083 (N_40083,N_39544,N_39609);
nand U40084 (N_40084,N_39723,N_39966);
nand U40085 (N_40085,N_39531,N_39633);
nor U40086 (N_40086,N_39843,N_39898);
or U40087 (N_40087,N_39707,N_39568);
nand U40088 (N_40088,N_39658,N_39961);
or U40089 (N_40089,N_39824,N_39728);
and U40090 (N_40090,N_39830,N_39957);
or U40091 (N_40091,N_39697,N_39778);
xor U40092 (N_40092,N_39857,N_39520);
nand U40093 (N_40093,N_39686,N_39522);
or U40094 (N_40094,N_39629,N_39711);
nor U40095 (N_40095,N_39630,N_39844);
xor U40096 (N_40096,N_39587,N_39940);
nor U40097 (N_40097,N_39721,N_39562);
and U40098 (N_40098,N_39941,N_39704);
nand U40099 (N_40099,N_39745,N_39967);
nor U40100 (N_40100,N_39870,N_39617);
or U40101 (N_40101,N_39586,N_39665);
nand U40102 (N_40102,N_39993,N_39950);
nand U40103 (N_40103,N_39754,N_39736);
xor U40104 (N_40104,N_39895,N_39786);
nand U40105 (N_40105,N_39871,N_39928);
and U40106 (N_40106,N_39887,N_39773);
xnor U40107 (N_40107,N_39935,N_39670);
and U40108 (N_40108,N_39538,N_39836);
nor U40109 (N_40109,N_39565,N_39653);
xnor U40110 (N_40110,N_39523,N_39570);
xnor U40111 (N_40111,N_39690,N_39614);
or U40112 (N_40112,N_39811,N_39507);
or U40113 (N_40113,N_39656,N_39533);
and U40114 (N_40114,N_39521,N_39924);
and U40115 (N_40115,N_39876,N_39535);
nor U40116 (N_40116,N_39755,N_39874);
xnor U40117 (N_40117,N_39582,N_39873);
nor U40118 (N_40118,N_39543,N_39904);
and U40119 (N_40119,N_39995,N_39807);
or U40120 (N_40120,N_39988,N_39557);
nor U40121 (N_40121,N_39896,N_39906);
xor U40122 (N_40122,N_39767,N_39612);
and U40123 (N_40123,N_39500,N_39820);
and U40124 (N_40124,N_39821,N_39766);
xor U40125 (N_40125,N_39792,N_39977);
nand U40126 (N_40126,N_39528,N_39514);
nor U40127 (N_40127,N_39551,N_39829);
and U40128 (N_40128,N_39952,N_39626);
xor U40129 (N_40129,N_39726,N_39949);
nand U40130 (N_40130,N_39827,N_39722);
xor U40131 (N_40131,N_39708,N_39580);
nor U40132 (N_40132,N_39803,N_39616);
or U40133 (N_40133,N_39991,N_39800);
nor U40134 (N_40134,N_39749,N_39980);
xor U40135 (N_40135,N_39555,N_39645);
nor U40136 (N_40136,N_39506,N_39632);
or U40137 (N_40137,N_39960,N_39663);
nor U40138 (N_40138,N_39592,N_39536);
xnor U40139 (N_40139,N_39782,N_39641);
or U40140 (N_40140,N_39529,N_39615);
nor U40141 (N_40141,N_39787,N_39735);
nand U40142 (N_40142,N_39770,N_39699);
xnor U40143 (N_40143,N_39678,N_39883);
xnor U40144 (N_40144,N_39826,N_39901);
and U40145 (N_40145,N_39642,N_39651);
nand U40146 (N_40146,N_39584,N_39872);
or U40147 (N_40147,N_39676,N_39938);
or U40148 (N_40148,N_39679,N_39801);
and U40149 (N_40149,N_39524,N_39759);
or U40150 (N_40150,N_39643,N_39693);
or U40151 (N_40151,N_39740,N_39621);
or U40152 (N_40152,N_39981,N_39716);
or U40153 (N_40153,N_39920,N_39856);
xnor U40154 (N_40154,N_39738,N_39620);
or U40155 (N_40155,N_39518,N_39933);
nor U40156 (N_40156,N_39793,N_39646);
nor U40157 (N_40157,N_39847,N_39908);
nor U40158 (N_40158,N_39899,N_39772);
xnor U40159 (N_40159,N_39606,N_39547);
nand U40160 (N_40160,N_39563,N_39931);
and U40161 (N_40161,N_39675,N_39789);
xnor U40162 (N_40162,N_39841,N_39982);
or U40163 (N_40163,N_39885,N_39743);
and U40164 (N_40164,N_39554,N_39677);
nand U40165 (N_40165,N_39588,N_39828);
and U40166 (N_40166,N_39947,N_39880);
xor U40167 (N_40167,N_39809,N_39881);
and U40168 (N_40168,N_39825,N_39956);
nand U40169 (N_40169,N_39710,N_39737);
and U40170 (N_40170,N_39838,N_39618);
or U40171 (N_40171,N_39561,N_39742);
or U40172 (N_40172,N_39703,N_39999);
or U40173 (N_40173,N_39845,N_39818);
nand U40174 (N_40174,N_39942,N_39834);
or U40175 (N_40175,N_39623,N_39540);
and U40176 (N_40176,N_39730,N_39953);
xor U40177 (N_40177,N_39516,N_39684);
or U40178 (N_40178,N_39971,N_39846);
nor U40179 (N_40179,N_39534,N_39569);
xor U40180 (N_40180,N_39913,N_39650);
xnor U40181 (N_40181,N_39613,N_39600);
nor U40182 (N_40182,N_39577,N_39576);
nor U40183 (N_40183,N_39854,N_39862);
and U40184 (N_40184,N_39861,N_39603);
xnor U40185 (N_40185,N_39802,N_39774);
nand U40186 (N_40186,N_39610,N_39835);
or U40187 (N_40187,N_39578,N_39997);
nand U40188 (N_40188,N_39954,N_39889);
or U40189 (N_40189,N_39503,N_39832);
and U40190 (N_40190,N_39888,N_39910);
nand U40191 (N_40191,N_39905,N_39903);
nand U40192 (N_40192,N_39705,N_39969);
nand U40193 (N_40193,N_39512,N_39816);
nand U40194 (N_40194,N_39602,N_39501);
nand U40195 (N_40195,N_39925,N_39855);
or U40196 (N_40196,N_39912,N_39706);
or U40197 (N_40197,N_39875,N_39859);
and U40198 (N_40198,N_39780,N_39849);
and U40199 (N_40199,N_39922,N_39719);
nand U40200 (N_40200,N_39648,N_39553);
nor U40201 (N_40201,N_39937,N_39804);
and U40202 (N_40202,N_39671,N_39994);
xnor U40203 (N_40203,N_39929,N_39744);
or U40204 (N_40204,N_39842,N_39720);
nand U40205 (N_40205,N_39878,N_39946);
nand U40206 (N_40206,N_39819,N_39851);
nand U40207 (N_40207,N_39691,N_39776);
and U40208 (N_40208,N_39868,N_39866);
nand U40209 (N_40209,N_39579,N_39549);
nand U40210 (N_40210,N_39964,N_39891);
or U40211 (N_40211,N_39647,N_39558);
nand U40212 (N_40212,N_39958,N_39853);
xor U40213 (N_40213,N_39948,N_39519);
and U40214 (N_40214,N_39753,N_39886);
or U40215 (N_40215,N_39968,N_39654);
and U40216 (N_40216,N_39771,N_39530);
nor U40217 (N_40217,N_39840,N_39823);
or U40218 (N_40218,N_39984,N_39955);
nand U40219 (N_40219,N_39607,N_39788);
nand U40220 (N_40220,N_39526,N_39595);
xor U40221 (N_40221,N_39890,N_39581);
nand U40222 (N_40222,N_39808,N_39989);
nor U40223 (N_40223,N_39797,N_39539);
xor U40224 (N_40224,N_39688,N_39527);
and U40225 (N_40225,N_39560,N_39934);
nor U40226 (N_40226,N_39718,N_39963);
nor U40227 (N_40227,N_39733,N_39657);
nor U40228 (N_40228,N_39852,N_39987);
xor U40229 (N_40229,N_39764,N_39532);
xor U40230 (N_40230,N_39864,N_39750);
nand U40231 (N_40231,N_39951,N_39734);
or U40232 (N_40232,N_39546,N_39732);
or U40233 (N_40233,N_39649,N_39599);
nor U40234 (N_40234,N_39589,N_39781);
xnor U40235 (N_40235,N_39805,N_39590);
and U40236 (N_40236,N_39959,N_39882);
xor U40237 (N_40237,N_39604,N_39757);
nand U40238 (N_40238,N_39799,N_39572);
and U40239 (N_40239,N_39644,N_39884);
nand U40240 (N_40240,N_39794,N_39902);
nor U40241 (N_40241,N_39682,N_39865);
and U40242 (N_40242,N_39760,N_39575);
nor U40243 (N_40243,N_39701,N_39879);
nor U40244 (N_40244,N_39661,N_39998);
or U40245 (N_40245,N_39673,N_39796);
xor U40246 (N_40246,N_39525,N_39986);
nor U40247 (N_40247,N_39962,N_39784);
xnor U40248 (N_40248,N_39894,N_39729);
and U40249 (N_40249,N_39970,N_39848);
or U40250 (N_40250,N_39571,N_39678);
nand U40251 (N_40251,N_39743,N_39564);
xnor U40252 (N_40252,N_39761,N_39834);
xnor U40253 (N_40253,N_39787,N_39583);
nand U40254 (N_40254,N_39892,N_39521);
xor U40255 (N_40255,N_39815,N_39625);
and U40256 (N_40256,N_39658,N_39800);
nor U40257 (N_40257,N_39515,N_39890);
and U40258 (N_40258,N_39830,N_39607);
xor U40259 (N_40259,N_39578,N_39691);
nor U40260 (N_40260,N_39635,N_39687);
xnor U40261 (N_40261,N_39960,N_39559);
or U40262 (N_40262,N_39767,N_39706);
nand U40263 (N_40263,N_39801,N_39738);
nor U40264 (N_40264,N_39682,N_39518);
nor U40265 (N_40265,N_39962,N_39677);
and U40266 (N_40266,N_39761,N_39644);
nor U40267 (N_40267,N_39505,N_39624);
nand U40268 (N_40268,N_39852,N_39686);
nor U40269 (N_40269,N_39578,N_39917);
nand U40270 (N_40270,N_39673,N_39731);
or U40271 (N_40271,N_39949,N_39510);
nor U40272 (N_40272,N_39920,N_39786);
and U40273 (N_40273,N_39614,N_39963);
or U40274 (N_40274,N_39633,N_39573);
nand U40275 (N_40275,N_39641,N_39840);
or U40276 (N_40276,N_39572,N_39995);
xnor U40277 (N_40277,N_39776,N_39679);
xor U40278 (N_40278,N_39973,N_39904);
and U40279 (N_40279,N_39969,N_39897);
nor U40280 (N_40280,N_39676,N_39977);
and U40281 (N_40281,N_39707,N_39609);
nor U40282 (N_40282,N_39863,N_39654);
xnor U40283 (N_40283,N_39692,N_39956);
and U40284 (N_40284,N_39836,N_39912);
or U40285 (N_40285,N_39627,N_39816);
nand U40286 (N_40286,N_39716,N_39917);
nor U40287 (N_40287,N_39781,N_39572);
nor U40288 (N_40288,N_39760,N_39872);
nand U40289 (N_40289,N_39831,N_39749);
nor U40290 (N_40290,N_39931,N_39786);
nand U40291 (N_40291,N_39986,N_39577);
nor U40292 (N_40292,N_39782,N_39954);
or U40293 (N_40293,N_39844,N_39610);
nand U40294 (N_40294,N_39576,N_39925);
xor U40295 (N_40295,N_39730,N_39877);
and U40296 (N_40296,N_39652,N_39801);
nand U40297 (N_40297,N_39875,N_39701);
nand U40298 (N_40298,N_39539,N_39607);
nand U40299 (N_40299,N_39934,N_39569);
nand U40300 (N_40300,N_39541,N_39995);
nand U40301 (N_40301,N_39920,N_39982);
nor U40302 (N_40302,N_39687,N_39735);
or U40303 (N_40303,N_39977,N_39811);
or U40304 (N_40304,N_39841,N_39809);
nor U40305 (N_40305,N_39797,N_39757);
xnor U40306 (N_40306,N_39777,N_39735);
and U40307 (N_40307,N_39891,N_39853);
and U40308 (N_40308,N_39535,N_39773);
xnor U40309 (N_40309,N_39706,N_39631);
and U40310 (N_40310,N_39774,N_39656);
and U40311 (N_40311,N_39930,N_39571);
and U40312 (N_40312,N_39872,N_39831);
nand U40313 (N_40313,N_39778,N_39504);
xnor U40314 (N_40314,N_39840,N_39604);
xnor U40315 (N_40315,N_39672,N_39770);
and U40316 (N_40316,N_39619,N_39799);
nor U40317 (N_40317,N_39667,N_39967);
and U40318 (N_40318,N_39968,N_39616);
nand U40319 (N_40319,N_39545,N_39968);
nand U40320 (N_40320,N_39773,N_39963);
nand U40321 (N_40321,N_39606,N_39590);
xnor U40322 (N_40322,N_39637,N_39509);
or U40323 (N_40323,N_39515,N_39792);
nand U40324 (N_40324,N_39823,N_39577);
xor U40325 (N_40325,N_39898,N_39823);
or U40326 (N_40326,N_39596,N_39986);
nand U40327 (N_40327,N_39527,N_39814);
and U40328 (N_40328,N_39807,N_39562);
xor U40329 (N_40329,N_39753,N_39637);
nand U40330 (N_40330,N_39804,N_39754);
xor U40331 (N_40331,N_39515,N_39940);
and U40332 (N_40332,N_39777,N_39949);
and U40333 (N_40333,N_39602,N_39683);
and U40334 (N_40334,N_39936,N_39924);
nand U40335 (N_40335,N_39819,N_39621);
and U40336 (N_40336,N_39891,N_39510);
or U40337 (N_40337,N_39826,N_39986);
and U40338 (N_40338,N_39902,N_39566);
xor U40339 (N_40339,N_39516,N_39815);
nand U40340 (N_40340,N_39670,N_39575);
xor U40341 (N_40341,N_39983,N_39525);
or U40342 (N_40342,N_39977,N_39766);
or U40343 (N_40343,N_39604,N_39928);
or U40344 (N_40344,N_39841,N_39987);
nand U40345 (N_40345,N_39555,N_39698);
xor U40346 (N_40346,N_39894,N_39687);
nand U40347 (N_40347,N_39831,N_39723);
nand U40348 (N_40348,N_39665,N_39541);
xnor U40349 (N_40349,N_39544,N_39946);
nand U40350 (N_40350,N_39542,N_39768);
nor U40351 (N_40351,N_39833,N_39795);
xor U40352 (N_40352,N_39667,N_39846);
xor U40353 (N_40353,N_39592,N_39936);
and U40354 (N_40354,N_39906,N_39520);
and U40355 (N_40355,N_39626,N_39872);
xor U40356 (N_40356,N_39983,N_39518);
nor U40357 (N_40357,N_39703,N_39894);
xor U40358 (N_40358,N_39933,N_39763);
nor U40359 (N_40359,N_39786,N_39867);
or U40360 (N_40360,N_39619,N_39816);
nor U40361 (N_40361,N_39581,N_39521);
and U40362 (N_40362,N_39561,N_39709);
or U40363 (N_40363,N_39725,N_39936);
nand U40364 (N_40364,N_39797,N_39698);
nand U40365 (N_40365,N_39535,N_39696);
or U40366 (N_40366,N_39536,N_39532);
nand U40367 (N_40367,N_39755,N_39660);
nor U40368 (N_40368,N_39642,N_39837);
nand U40369 (N_40369,N_39919,N_39730);
or U40370 (N_40370,N_39832,N_39833);
xnor U40371 (N_40371,N_39513,N_39843);
xnor U40372 (N_40372,N_39606,N_39594);
xnor U40373 (N_40373,N_39866,N_39725);
or U40374 (N_40374,N_39921,N_39522);
and U40375 (N_40375,N_39613,N_39907);
nand U40376 (N_40376,N_39721,N_39871);
and U40377 (N_40377,N_39807,N_39708);
nor U40378 (N_40378,N_39581,N_39673);
or U40379 (N_40379,N_39842,N_39512);
nand U40380 (N_40380,N_39925,N_39951);
or U40381 (N_40381,N_39913,N_39853);
or U40382 (N_40382,N_39949,N_39816);
or U40383 (N_40383,N_39950,N_39612);
nor U40384 (N_40384,N_39512,N_39762);
nand U40385 (N_40385,N_39617,N_39624);
xor U40386 (N_40386,N_39824,N_39754);
nand U40387 (N_40387,N_39749,N_39681);
or U40388 (N_40388,N_39904,N_39505);
nand U40389 (N_40389,N_39927,N_39863);
and U40390 (N_40390,N_39864,N_39500);
xnor U40391 (N_40391,N_39882,N_39626);
or U40392 (N_40392,N_39583,N_39595);
xor U40393 (N_40393,N_39964,N_39769);
nand U40394 (N_40394,N_39717,N_39631);
or U40395 (N_40395,N_39856,N_39673);
nand U40396 (N_40396,N_39838,N_39948);
xor U40397 (N_40397,N_39734,N_39700);
or U40398 (N_40398,N_39784,N_39723);
and U40399 (N_40399,N_39895,N_39735);
xnor U40400 (N_40400,N_39685,N_39574);
and U40401 (N_40401,N_39967,N_39579);
xnor U40402 (N_40402,N_39997,N_39896);
nor U40403 (N_40403,N_39503,N_39897);
xnor U40404 (N_40404,N_39885,N_39872);
nor U40405 (N_40405,N_39758,N_39571);
xor U40406 (N_40406,N_39712,N_39679);
or U40407 (N_40407,N_39765,N_39569);
or U40408 (N_40408,N_39665,N_39675);
nand U40409 (N_40409,N_39719,N_39816);
and U40410 (N_40410,N_39913,N_39831);
nand U40411 (N_40411,N_39508,N_39987);
or U40412 (N_40412,N_39913,N_39787);
or U40413 (N_40413,N_39831,N_39758);
nor U40414 (N_40414,N_39859,N_39817);
or U40415 (N_40415,N_39838,N_39827);
and U40416 (N_40416,N_39900,N_39924);
nand U40417 (N_40417,N_39973,N_39985);
nor U40418 (N_40418,N_39675,N_39551);
nor U40419 (N_40419,N_39515,N_39896);
nand U40420 (N_40420,N_39987,N_39850);
xnor U40421 (N_40421,N_39783,N_39566);
or U40422 (N_40422,N_39523,N_39623);
xnor U40423 (N_40423,N_39995,N_39757);
nor U40424 (N_40424,N_39521,N_39633);
or U40425 (N_40425,N_39982,N_39825);
or U40426 (N_40426,N_39743,N_39965);
or U40427 (N_40427,N_39987,N_39898);
xor U40428 (N_40428,N_39562,N_39537);
xnor U40429 (N_40429,N_39578,N_39731);
nand U40430 (N_40430,N_39973,N_39594);
xnor U40431 (N_40431,N_39839,N_39746);
nor U40432 (N_40432,N_39768,N_39519);
nand U40433 (N_40433,N_39791,N_39986);
xnor U40434 (N_40434,N_39918,N_39998);
xnor U40435 (N_40435,N_39673,N_39750);
nand U40436 (N_40436,N_39581,N_39642);
and U40437 (N_40437,N_39545,N_39982);
xnor U40438 (N_40438,N_39553,N_39757);
nand U40439 (N_40439,N_39974,N_39708);
nor U40440 (N_40440,N_39704,N_39730);
nand U40441 (N_40441,N_39831,N_39641);
nor U40442 (N_40442,N_39744,N_39847);
and U40443 (N_40443,N_39974,N_39562);
xor U40444 (N_40444,N_39589,N_39510);
xnor U40445 (N_40445,N_39778,N_39531);
nor U40446 (N_40446,N_39960,N_39856);
or U40447 (N_40447,N_39641,N_39875);
xor U40448 (N_40448,N_39787,N_39526);
nor U40449 (N_40449,N_39870,N_39705);
and U40450 (N_40450,N_39830,N_39638);
xor U40451 (N_40451,N_39585,N_39645);
or U40452 (N_40452,N_39892,N_39798);
and U40453 (N_40453,N_39653,N_39591);
or U40454 (N_40454,N_39776,N_39999);
nand U40455 (N_40455,N_39713,N_39612);
xnor U40456 (N_40456,N_39641,N_39612);
and U40457 (N_40457,N_39536,N_39697);
nor U40458 (N_40458,N_39978,N_39920);
and U40459 (N_40459,N_39832,N_39848);
nor U40460 (N_40460,N_39866,N_39500);
xnor U40461 (N_40461,N_39553,N_39915);
and U40462 (N_40462,N_39965,N_39682);
or U40463 (N_40463,N_39848,N_39570);
nor U40464 (N_40464,N_39938,N_39516);
nor U40465 (N_40465,N_39647,N_39881);
nor U40466 (N_40466,N_39906,N_39725);
nand U40467 (N_40467,N_39675,N_39691);
nor U40468 (N_40468,N_39913,N_39715);
nand U40469 (N_40469,N_39997,N_39607);
and U40470 (N_40470,N_39601,N_39926);
or U40471 (N_40471,N_39832,N_39772);
and U40472 (N_40472,N_39696,N_39583);
nor U40473 (N_40473,N_39596,N_39669);
nor U40474 (N_40474,N_39654,N_39925);
and U40475 (N_40475,N_39727,N_39925);
or U40476 (N_40476,N_39824,N_39500);
xor U40477 (N_40477,N_39961,N_39509);
or U40478 (N_40478,N_39822,N_39977);
nor U40479 (N_40479,N_39602,N_39975);
and U40480 (N_40480,N_39801,N_39823);
xnor U40481 (N_40481,N_39586,N_39690);
nand U40482 (N_40482,N_39731,N_39648);
or U40483 (N_40483,N_39843,N_39885);
or U40484 (N_40484,N_39757,N_39581);
nor U40485 (N_40485,N_39718,N_39872);
nor U40486 (N_40486,N_39911,N_39558);
and U40487 (N_40487,N_39864,N_39724);
and U40488 (N_40488,N_39913,N_39779);
and U40489 (N_40489,N_39638,N_39725);
and U40490 (N_40490,N_39759,N_39772);
xor U40491 (N_40491,N_39761,N_39786);
or U40492 (N_40492,N_39885,N_39528);
nor U40493 (N_40493,N_39837,N_39715);
nor U40494 (N_40494,N_39533,N_39580);
or U40495 (N_40495,N_39522,N_39876);
xor U40496 (N_40496,N_39828,N_39798);
and U40497 (N_40497,N_39735,N_39740);
nor U40498 (N_40498,N_39648,N_39953);
nor U40499 (N_40499,N_39733,N_39777);
nand U40500 (N_40500,N_40212,N_40353);
xnor U40501 (N_40501,N_40097,N_40211);
nor U40502 (N_40502,N_40448,N_40465);
or U40503 (N_40503,N_40366,N_40352);
xnor U40504 (N_40504,N_40390,N_40089);
nor U40505 (N_40505,N_40490,N_40110);
xor U40506 (N_40506,N_40179,N_40299);
xnor U40507 (N_40507,N_40162,N_40153);
xor U40508 (N_40508,N_40106,N_40358);
xor U40509 (N_40509,N_40269,N_40165);
xor U40510 (N_40510,N_40345,N_40234);
xnor U40511 (N_40511,N_40334,N_40317);
nand U40512 (N_40512,N_40099,N_40157);
or U40513 (N_40513,N_40050,N_40458);
nor U40514 (N_40514,N_40046,N_40113);
nand U40515 (N_40515,N_40047,N_40178);
nand U40516 (N_40516,N_40237,N_40004);
or U40517 (N_40517,N_40051,N_40218);
nand U40518 (N_40518,N_40067,N_40470);
and U40519 (N_40519,N_40138,N_40032);
and U40520 (N_40520,N_40406,N_40336);
nand U40521 (N_40521,N_40284,N_40319);
nor U40522 (N_40522,N_40135,N_40104);
nand U40523 (N_40523,N_40363,N_40360);
nand U40524 (N_40524,N_40452,N_40308);
nand U40525 (N_40525,N_40100,N_40441);
nor U40526 (N_40526,N_40320,N_40231);
xor U40527 (N_40527,N_40484,N_40028);
nand U40528 (N_40528,N_40226,N_40344);
and U40529 (N_40529,N_40103,N_40027);
or U40530 (N_40530,N_40161,N_40139);
nand U40531 (N_40531,N_40025,N_40467);
or U40532 (N_40532,N_40393,N_40164);
or U40533 (N_40533,N_40193,N_40439);
nor U40534 (N_40534,N_40418,N_40070);
and U40535 (N_40535,N_40453,N_40267);
xor U40536 (N_40536,N_40496,N_40488);
or U40537 (N_40537,N_40374,N_40029);
or U40538 (N_40538,N_40222,N_40447);
or U40539 (N_40539,N_40213,N_40313);
nand U40540 (N_40540,N_40365,N_40183);
or U40541 (N_40541,N_40065,N_40119);
or U40542 (N_40542,N_40301,N_40391);
nand U40543 (N_40543,N_40235,N_40400);
or U40544 (N_40544,N_40056,N_40274);
and U40545 (N_40545,N_40087,N_40117);
nand U40546 (N_40546,N_40483,N_40149);
or U40547 (N_40547,N_40300,N_40081);
xnor U40548 (N_40548,N_40209,N_40294);
nand U40549 (N_40549,N_40464,N_40159);
nand U40550 (N_40550,N_40475,N_40482);
nand U40551 (N_40551,N_40250,N_40077);
nand U40552 (N_40552,N_40037,N_40187);
nor U40553 (N_40553,N_40380,N_40480);
nor U40554 (N_40554,N_40023,N_40341);
or U40555 (N_40555,N_40287,N_40128);
nor U40556 (N_40556,N_40392,N_40039);
nand U40557 (N_40557,N_40463,N_40355);
nor U40558 (N_40558,N_40134,N_40206);
and U40559 (N_40559,N_40003,N_40262);
nand U40560 (N_40560,N_40002,N_40474);
nand U40561 (N_40561,N_40421,N_40411);
or U40562 (N_40562,N_40306,N_40182);
or U40563 (N_40563,N_40019,N_40361);
nand U40564 (N_40564,N_40498,N_40455);
and U40565 (N_40565,N_40381,N_40057);
and U40566 (N_40566,N_40090,N_40265);
xnor U40567 (N_40567,N_40072,N_40438);
or U40568 (N_40568,N_40216,N_40412);
nor U40569 (N_40569,N_40220,N_40311);
or U40570 (N_40570,N_40066,N_40275);
xor U40571 (N_40571,N_40401,N_40131);
xnor U40572 (N_40572,N_40395,N_40091);
and U40573 (N_40573,N_40342,N_40232);
xor U40574 (N_40574,N_40196,N_40052);
nor U40575 (N_40575,N_40180,N_40174);
nor U40576 (N_40576,N_40230,N_40102);
nor U40577 (N_40577,N_40433,N_40410);
nor U40578 (N_40578,N_40095,N_40170);
and U40579 (N_40579,N_40279,N_40315);
nor U40580 (N_40580,N_40442,N_40325);
nand U40581 (N_40581,N_40141,N_40191);
nand U40582 (N_40582,N_40307,N_40053);
nand U40583 (N_40583,N_40327,N_40258);
nand U40584 (N_40584,N_40343,N_40350);
nor U40585 (N_40585,N_40322,N_40396);
or U40586 (N_40586,N_40010,N_40451);
xnor U40587 (N_40587,N_40389,N_40324);
nor U40588 (N_40588,N_40477,N_40449);
and U40589 (N_40589,N_40120,N_40469);
and U40590 (N_40590,N_40473,N_40253);
nor U40591 (N_40591,N_40125,N_40219);
or U40592 (N_40592,N_40247,N_40198);
xor U40593 (N_40593,N_40368,N_40493);
or U40594 (N_40594,N_40166,N_40036);
xor U40595 (N_40595,N_40064,N_40257);
and U40596 (N_40596,N_40001,N_40085);
nor U40597 (N_40597,N_40491,N_40338);
nor U40598 (N_40598,N_40163,N_40351);
and U40599 (N_40599,N_40158,N_40414);
nor U40600 (N_40600,N_40116,N_40271);
nor U40601 (N_40601,N_40244,N_40446);
nor U40602 (N_40602,N_40186,N_40487);
or U40603 (N_40603,N_40243,N_40321);
nand U40604 (N_40604,N_40238,N_40098);
or U40605 (N_40605,N_40378,N_40424);
xnor U40606 (N_40606,N_40478,N_40221);
nor U40607 (N_40607,N_40015,N_40362);
or U40608 (N_40608,N_40370,N_40031);
nor U40609 (N_40609,N_40118,N_40172);
or U40610 (N_40610,N_40335,N_40021);
nand U40611 (N_40611,N_40202,N_40022);
nand U40612 (N_40612,N_40248,N_40073);
nand U40613 (N_40613,N_40115,N_40006);
and U40614 (N_40614,N_40456,N_40086);
nand U40615 (N_40615,N_40160,N_40429);
nor U40616 (N_40616,N_40318,N_40249);
and U40617 (N_40617,N_40376,N_40282);
nand U40618 (N_40618,N_40111,N_40379);
nor U40619 (N_40619,N_40286,N_40194);
nand U40620 (N_40620,N_40304,N_40397);
or U40621 (N_40621,N_40024,N_40328);
and U40622 (N_40622,N_40215,N_40330);
and U40623 (N_40623,N_40356,N_40444);
or U40624 (N_40624,N_40228,N_40137);
nand U40625 (N_40625,N_40289,N_40144);
nor U40626 (N_40626,N_40074,N_40233);
xnor U40627 (N_40627,N_40489,N_40101);
or U40628 (N_40628,N_40272,N_40079);
xnor U40629 (N_40629,N_40476,N_40388);
and U40630 (N_40630,N_40254,N_40096);
or U40631 (N_40631,N_40405,N_40428);
or U40632 (N_40632,N_40075,N_40359);
and U40633 (N_40633,N_40434,N_40340);
nand U40634 (N_40634,N_40154,N_40329);
nand U40635 (N_40635,N_40246,N_40078);
nand U40636 (N_40636,N_40305,N_40485);
nand U40637 (N_40637,N_40038,N_40255);
xnor U40638 (N_40638,N_40277,N_40176);
or U40639 (N_40639,N_40092,N_40309);
or U40640 (N_40640,N_40200,N_40132);
nand U40641 (N_40641,N_40020,N_40285);
xnor U40642 (N_40642,N_40175,N_40084);
xor U40643 (N_40643,N_40142,N_40382);
and U40644 (N_40644,N_40152,N_40059);
nor U40645 (N_40645,N_40109,N_40454);
nand U40646 (N_40646,N_40492,N_40008);
and U40647 (N_40647,N_40012,N_40018);
xnor U40648 (N_40648,N_40207,N_40346);
and U40649 (N_40649,N_40331,N_40369);
nand U40650 (N_40650,N_40189,N_40416);
nand U40651 (N_40651,N_40326,N_40042);
xnor U40652 (N_40652,N_40303,N_40017);
or U40653 (N_40653,N_40204,N_40140);
or U40654 (N_40654,N_40419,N_40167);
and U40655 (N_40655,N_40208,N_40143);
nor U40656 (N_40656,N_40133,N_40423);
or U40657 (N_40657,N_40339,N_40443);
xnor U40658 (N_40658,N_40403,N_40290);
xnor U40659 (N_40659,N_40188,N_40121);
nand U40660 (N_40660,N_40385,N_40241);
nand U40661 (N_40661,N_40043,N_40124);
xor U40662 (N_40662,N_40147,N_40045);
and U40663 (N_40663,N_40227,N_40136);
nor U40664 (N_40664,N_40058,N_40192);
nand U40665 (N_40665,N_40375,N_40432);
xnor U40666 (N_40666,N_40151,N_40472);
or U40667 (N_40667,N_40349,N_40276);
nand U40668 (N_40668,N_40377,N_40127);
xnor U40669 (N_40669,N_40150,N_40223);
nand U40670 (N_40670,N_40011,N_40060);
or U40671 (N_40671,N_40460,N_40259);
nor U40672 (N_40672,N_40314,N_40291);
nor U40673 (N_40673,N_40016,N_40114);
xnor U40674 (N_40674,N_40364,N_40417);
or U40675 (N_40675,N_40076,N_40061);
xnor U40676 (N_40676,N_40148,N_40394);
xor U40677 (N_40677,N_40214,N_40422);
xnor U40678 (N_40678,N_40486,N_40499);
xor U40679 (N_40679,N_40190,N_40281);
nor U40680 (N_40680,N_40252,N_40266);
or U40681 (N_40681,N_40445,N_40431);
nor U40682 (N_40682,N_40122,N_40278);
and U40683 (N_40683,N_40000,N_40040);
or U40684 (N_40684,N_40312,N_40479);
nand U40685 (N_40685,N_40229,N_40173);
nor U40686 (N_40686,N_40013,N_40203);
xnor U40687 (N_40687,N_40112,N_40415);
or U40688 (N_40688,N_40145,N_40270);
nand U40689 (N_40689,N_40014,N_40156);
and U40690 (N_40690,N_40195,N_40407);
xnor U40691 (N_40691,N_40373,N_40034);
nand U40692 (N_40692,N_40261,N_40386);
xor U40693 (N_40693,N_40387,N_40168);
or U40694 (N_40694,N_40372,N_40129);
nor U40695 (N_40695,N_40055,N_40199);
nor U40696 (N_40696,N_40080,N_40332);
nor U40697 (N_40697,N_40466,N_40384);
and U40698 (N_40698,N_40177,N_40296);
and U40699 (N_40699,N_40041,N_40107);
and U40700 (N_40700,N_40030,N_40273);
nand U40701 (N_40701,N_40297,N_40316);
nand U40702 (N_40702,N_40408,N_40007);
or U40703 (N_40703,N_40044,N_40093);
nand U40704 (N_40704,N_40048,N_40054);
nor U40705 (N_40705,N_40242,N_40437);
xor U40706 (N_40706,N_40292,N_40409);
nand U40707 (N_40707,N_40399,N_40201);
or U40708 (N_40708,N_40240,N_40283);
nor U40709 (N_40709,N_40383,N_40123);
or U40710 (N_40710,N_40197,N_40413);
and U40711 (N_40711,N_40181,N_40217);
xor U40712 (N_40712,N_40298,N_40459);
and U40713 (N_40713,N_40239,N_40302);
and U40714 (N_40714,N_40425,N_40251);
or U40715 (N_40715,N_40426,N_40481);
nor U40716 (N_40716,N_40268,N_40462);
or U40717 (N_40717,N_40371,N_40169);
or U40718 (N_40718,N_40062,N_40310);
and U40719 (N_40719,N_40436,N_40069);
and U40720 (N_40720,N_40185,N_40468);
xor U40721 (N_40721,N_40357,N_40071);
or U40722 (N_40722,N_40404,N_40005);
nor U40723 (N_40723,N_40494,N_40224);
xor U40724 (N_40724,N_40260,N_40348);
nand U40725 (N_40725,N_40323,N_40427);
and U40726 (N_40726,N_40367,N_40094);
xor U40727 (N_40727,N_40009,N_40245);
or U40728 (N_40728,N_40126,N_40402);
nor U40729 (N_40729,N_40295,N_40457);
or U40730 (N_40730,N_40264,N_40347);
and U40731 (N_40731,N_40184,N_40105);
or U40732 (N_40732,N_40435,N_40263);
xor U40733 (N_40733,N_40450,N_40280);
nand U40734 (N_40734,N_40430,N_40083);
nor U40735 (N_40735,N_40236,N_40063);
xor U40736 (N_40736,N_40497,N_40225);
nand U40737 (N_40737,N_40398,N_40440);
nand U40738 (N_40738,N_40256,N_40068);
or U40739 (N_40739,N_40155,N_40471);
and U40740 (N_40740,N_40495,N_40108);
xor U40741 (N_40741,N_40026,N_40146);
or U40742 (N_40742,N_40205,N_40035);
and U40743 (N_40743,N_40420,N_40171);
xor U40744 (N_40744,N_40049,N_40288);
and U40745 (N_40745,N_40461,N_40337);
nor U40746 (N_40746,N_40082,N_40293);
nand U40747 (N_40747,N_40354,N_40210);
xor U40748 (N_40748,N_40130,N_40088);
and U40749 (N_40749,N_40333,N_40033);
nor U40750 (N_40750,N_40150,N_40246);
nand U40751 (N_40751,N_40118,N_40432);
xnor U40752 (N_40752,N_40064,N_40402);
xnor U40753 (N_40753,N_40024,N_40352);
or U40754 (N_40754,N_40048,N_40257);
nor U40755 (N_40755,N_40216,N_40105);
nand U40756 (N_40756,N_40165,N_40137);
and U40757 (N_40757,N_40165,N_40429);
or U40758 (N_40758,N_40029,N_40302);
or U40759 (N_40759,N_40498,N_40465);
xnor U40760 (N_40760,N_40088,N_40169);
or U40761 (N_40761,N_40402,N_40356);
or U40762 (N_40762,N_40295,N_40337);
nor U40763 (N_40763,N_40461,N_40182);
nand U40764 (N_40764,N_40185,N_40323);
nor U40765 (N_40765,N_40453,N_40435);
nor U40766 (N_40766,N_40221,N_40302);
nor U40767 (N_40767,N_40146,N_40200);
nand U40768 (N_40768,N_40187,N_40156);
nand U40769 (N_40769,N_40203,N_40043);
or U40770 (N_40770,N_40302,N_40018);
and U40771 (N_40771,N_40026,N_40375);
or U40772 (N_40772,N_40248,N_40127);
or U40773 (N_40773,N_40475,N_40418);
or U40774 (N_40774,N_40228,N_40066);
or U40775 (N_40775,N_40254,N_40111);
xor U40776 (N_40776,N_40369,N_40278);
nand U40777 (N_40777,N_40023,N_40227);
nor U40778 (N_40778,N_40080,N_40168);
nor U40779 (N_40779,N_40300,N_40173);
nor U40780 (N_40780,N_40087,N_40449);
or U40781 (N_40781,N_40245,N_40110);
nand U40782 (N_40782,N_40351,N_40277);
xor U40783 (N_40783,N_40177,N_40141);
xor U40784 (N_40784,N_40448,N_40307);
and U40785 (N_40785,N_40024,N_40468);
nand U40786 (N_40786,N_40357,N_40118);
xor U40787 (N_40787,N_40295,N_40244);
and U40788 (N_40788,N_40410,N_40251);
nor U40789 (N_40789,N_40262,N_40112);
nor U40790 (N_40790,N_40493,N_40320);
xnor U40791 (N_40791,N_40082,N_40201);
and U40792 (N_40792,N_40243,N_40016);
and U40793 (N_40793,N_40398,N_40084);
and U40794 (N_40794,N_40415,N_40490);
nor U40795 (N_40795,N_40175,N_40310);
nor U40796 (N_40796,N_40106,N_40129);
and U40797 (N_40797,N_40251,N_40063);
or U40798 (N_40798,N_40297,N_40198);
nor U40799 (N_40799,N_40293,N_40160);
xnor U40800 (N_40800,N_40360,N_40119);
nand U40801 (N_40801,N_40196,N_40475);
nand U40802 (N_40802,N_40003,N_40110);
and U40803 (N_40803,N_40328,N_40394);
and U40804 (N_40804,N_40192,N_40122);
xor U40805 (N_40805,N_40225,N_40006);
or U40806 (N_40806,N_40063,N_40395);
nor U40807 (N_40807,N_40422,N_40425);
or U40808 (N_40808,N_40117,N_40276);
or U40809 (N_40809,N_40363,N_40140);
xnor U40810 (N_40810,N_40371,N_40396);
and U40811 (N_40811,N_40461,N_40397);
or U40812 (N_40812,N_40073,N_40127);
xor U40813 (N_40813,N_40175,N_40471);
nor U40814 (N_40814,N_40213,N_40167);
nand U40815 (N_40815,N_40067,N_40115);
xor U40816 (N_40816,N_40173,N_40480);
xor U40817 (N_40817,N_40408,N_40138);
nor U40818 (N_40818,N_40430,N_40136);
and U40819 (N_40819,N_40433,N_40058);
xnor U40820 (N_40820,N_40413,N_40418);
nor U40821 (N_40821,N_40257,N_40074);
xor U40822 (N_40822,N_40365,N_40495);
and U40823 (N_40823,N_40225,N_40458);
and U40824 (N_40824,N_40378,N_40461);
nor U40825 (N_40825,N_40182,N_40126);
xnor U40826 (N_40826,N_40108,N_40004);
nand U40827 (N_40827,N_40477,N_40067);
or U40828 (N_40828,N_40313,N_40193);
and U40829 (N_40829,N_40433,N_40005);
nor U40830 (N_40830,N_40229,N_40035);
and U40831 (N_40831,N_40095,N_40160);
xnor U40832 (N_40832,N_40330,N_40463);
nand U40833 (N_40833,N_40111,N_40449);
xor U40834 (N_40834,N_40240,N_40063);
nor U40835 (N_40835,N_40228,N_40063);
xor U40836 (N_40836,N_40478,N_40276);
nor U40837 (N_40837,N_40077,N_40260);
and U40838 (N_40838,N_40179,N_40442);
and U40839 (N_40839,N_40449,N_40156);
nor U40840 (N_40840,N_40102,N_40190);
or U40841 (N_40841,N_40356,N_40243);
or U40842 (N_40842,N_40042,N_40256);
and U40843 (N_40843,N_40143,N_40020);
and U40844 (N_40844,N_40241,N_40214);
and U40845 (N_40845,N_40209,N_40359);
nand U40846 (N_40846,N_40156,N_40127);
xor U40847 (N_40847,N_40430,N_40247);
xor U40848 (N_40848,N_40409,N_40358);
and U40849 (N_40849,N_40160,N_40332);
nand U40850 (N_40850,N_40057,N_40369);
xor U40851 (N_40851,N_40087,N_40351);
or U40852 (N_40852,N_40152,N_40145);
nor U40853 (N_40853,N_40104,N_40377);
nor U40854 (N_40854,N_40066,N_40366);
or U40855 (N_40855,N_40247,N_40485);
xor U40856 (N_40856,N_40069,N_40196);
nand U40857 (N_40857,N_40282,N_40338);
xnor U40858 (N_40858,N_40290,N_40309);
xnor U40859 (N_40859,N_40055,N_40407);
and U40860 (N_40860,N_40313,N_40229);
or U40861 (N_40861,N_40399,N_40080);
and U40862 (N_40862,N_40404,N_40200);
xor U40863 (N_40863,N_40217,N_40078);
and U40864 (N_40864,N_40046,N_40070);
nor U40865 (N_40865,N_40413,N_40309);
nor U40866 (N_40866,N_40146,N_40213);
nand U40867 (N_40867,N_40069,N_40255);
and U40868 (N_40868,N_40374,N_40453);
nand U40869 (N_40869,N_40378,N_40074);
xor U40870 (N_40870,N_40140,N_40406);
nand U40871 (N_40871,N_40064,N_40179);
xor U40872 (N_40872,N_40215,N_40154);
xnor U40873 (N_40873,N_40126,N_40325);
and U40874 (N_40874,N_40007,N_40282);
nor U40875 (N_40875,N_40077,N_40274);
or U40876 (N_40876,N_40131,N_40306);
xor U40877 (N_40877,N_40385,N_40331);
and U40878 (N_40878,N_40130,N_40423);
nor U40879 (N_40879,N_40166,N_40161);
nand U40880 (N_40880,N_40270,N_40435);
nand U40881 (N_40881,N_40262,N_40276);
or U40882 (N_40882,N_40394,N_40065);
nand U40883 (N_40883,N_40257,N_40015);
or U40884 (N_40884,N_40373,N_40343);
nor U40885 (N_40885,N_40110,N_40099);
nor U40886 (N_40886,N_40337,N_40205);
nand U40887 (N_40887,N_40355,N_40497);
nand U40888 (N_40888,N_40057,N_40396);
nand U40889 (N_40889,N_40241,N_40149);
xnor U40890 (N_40890,N_40392,N_40024);
or U40891 (N_40891,N_40398,N_40162);
nand U40892 (N_40892,N_40183,N_40250);
and U40893 (N_40893,N_40183,N_40198);
and U40894 (N_40894,N_40078,N_40327);
and U40895 (N_40895,N_40311,N_40487);
nand U40896 (N_40896,N_40181,N_40030);
or U40897 (N_40897,N_40432,N_40039);
and U40898 (N_40898,N_40129,N_40060);
or U40899 (N_40899,N_40160,N_40210);
nor U40900 (N_40900,N_40234,N_40323);
nand U40901 (N_40901,N_40327,N_40063);
nand U40902 (N_40902,N_40106,N_40303);
nand U40903 (N_40903,N_40327,N_40143);
or U40904 (N_40904,N_40301,N_40072);
or U40905 (N_40905,N_40437,N_40448);
and U40906 (N_40906,N_40101,N_40054);
nor U40907 (N_40907,N_40259,N_40177);
and U40908 (N_40908,N_40201,N_40303);
xnor U40909 (N_40909,N_40292,N_40023);
nor U40910 (N_40910,N_40342,N_40368);
or U40911 (N_40911,N_40054,N_40226);
nand U40912 (N_40912,N_40075,N_40003);
nor U40913 (N_40913,N_40023,N_40219);
xor U40914 (N_40914,N_40272,N_40194);
nor U40915 (N_40915,N_40012,N_40438);
and U40916 (N_40916,N_40274,N_40286);
xnor U40917 (N_40917,N_40267,N_40026);
nor U40918 (N_40918,N_40224,N_40068);
xor U40919 (N_40919,N_40444,N_40180);
and U40920 (N_40920,N_40034,N_40107);
xnor U40921 (N_40921,N_40436,N_40124);
and U40922 (N_40922,N_40445,N_40007);
or U40923 (N_40923,N_40067,N_40136);
xor U40924 (N_40924,N_40396,N_40279);
or U40925 (N_40925,N_40484,N_40264);
xor U40926 (N_40926,N_40214,N_40187);
nand U40927 (N_40927,N_40225,N_40209);
nor U40928 (N_40928,N_40267,N_40169);
or U40929 (N_40929,N_40232,N_40206);
xnor U40930 (N_40930,N_40085,N_40021);
xnor U40931 (N_40931,N_40149,N_40218);
or U40932 (N_40932,N_40021,N_40447);
or U40933 (N_40933,N_40134,N_40463);
nor U40934 (N_40934,N_40389,N_40318);
nor U40935 (N_40935,N_40357,N_40160);
or U40936 (N_40936,N_40415,N_40199);
and U40937 (N_40937,N_40285,N_40360);
or U40938 (N_40938,N_40258,N_40420);
or U40939 (N_40939,N_40025,N_40372);
nand U40940 (N_40940,N_40194,N_40439);
nand U40941 (N_40941,N_40216,N_40081);
nand U40942 (N_40942,N_40085,N_40064);
nor U40943 (N_40943,N_40267,N_40190);
and U40944 (N_40944,N_40429,N_40010);
and U40945 (N_40945,N_40098,N_40249);
nand U40946 (N_40946,N_40173,N_40499);
and U40947 (N_40947,N_40145,N_40213);
or U40948 (N_40948,N_40385,N_40229);
or U40949 (N_40949,N_40370,N_40098);
xnor U40950 (N_40950,N_40132,N_40256);
or U40951 (N_40951,N_40344,N_40496);
nand U40952 (N_40952,N_40221,N_40045);
nor U40953 (N_40953,N_40391,N_40324);
xor U40954 (N_40954,N_40074,N_40259);
or U40955 (N_40955,N_40048,N_40206);
nand U40956 (N_40956,N_40299,N_40055);
nor U40957 (N_40957,N_40272,N_40474);
and U40958 (N_40958,N_40412,N_40135);
and U40959 (N_40959,N_40380,N_40250);
and U40960 (N_40960,N_40370,N_40190);
and U40961 (N_40961,N_40176,N_40073);
and U40962 (N_40962,N_40305,N_40492);
xnor U40963 (N_40963,N_40358,N_40283);
nand U40964 (N_40964,N_40169,N_40460);
nor U40965 (N_40965,N_40400,N_40041);
nor U40966 (N_40966,N_40049,N_40138);
or U40967 (N_40967,N_40074,N_40129);
or U40968 (N_40968,N_40045,N_40105);
nor U40969 (N_40969,N_40069,N_40330);
or U40970 (N_40970,N_40362,N_40452);
and U40971 (N_40971,N_40036,N_40263);
nor U40972 (N_40972,N_40487,N_40302);
nand U40973 (N_40973,N_40287,N_40309);
or U40974 (N_40974,N_40489,N_40139);
xnor U40975 (N_40975,N_40342,N_40050);
xor U40976 (N_40976,N_40212,N_40166);
and U40977 (N_40977,N_40162,N_40058);
nor U40978 (N_40978,N_40423,N_40230);
xor U40979 (N_40979,N_40450,N_40112);
nand U40980 (N_40980,N_40135,N_40297);
or U40981 (N_40981,N_40299,N_40472);
xnor U40982 (N_40982,N_40411,N_40007);
nand U40983 (N_40983,N_40198,N_40306);
nor U40984 (N_40984,N_40322,N_40466);
xor U40985 (N_40985,N_40124,N_40163);
nand U40986 (N_40986,N_40459,N_40359);
nand U40987 (N_40987,N_40419,N_40324);
or U40988 (N_40988,N_40146,N_40051);
or U40989 (N_40989,N_40417,N_40343);
and U40990 (N_40990,N_40449,N_40359);
nand U40991 (N_40991,N_40070,N_40165);
nand U40992 (N_40992,N_40436,N_40315);
nor U40993 (N_40993,N_40247,N_40320);
nand U40994 (N_40994,N_40150,N_40276);
or U40995 (N_40995,N_40009,N_40082);
nand U40996 (N_40996,N_40266,N_40428);
xor U40997 (N_40997,N_40135,N_40304);
or U40998 (N_40998,N_40121,N_40093);
nand U40999 (N_40999,N_40054,N_40234);
or U41000 (N_41000,N_40591,N_40869);
xor U41001 (N_41001,N_40642,N_40758);
nand U41002 (N_41002,N_40941,N_40977);
and U41003 (N_41003,N_40601,N_40722);
nor U41004 (N_41004,N_40626,N_40937);
xnor U41005 (N_41005,N_40650,N_40654);
and U41006 (N_41006,N_40605,N_40594);
nor U41007 (N_41007,N_40628,N_40533);
or U41008 (N_41008,N_40567,N_40677);
xnor U41009 (N_41009,N_40645,N_40939);
or U41010 (N_41010,N_40715,N_40827);
xnor U41011 (N_41011,N_40515,N_40788);
xnor U41012 (N_41012,N_40978,N_40948);
xnor U41013 (N_41013,N_40706,N_40569);
nand U41014 (N_41014,N_40551,N_40570);
and U41015 (N_41015,N_40519,N_40998);
nand U41016 (N_41016,N_40882,N_40621);
and U41017 (N_41017,N_40709,N_40790);
nor U41018 (N_41018,N_40683,N_40983);
xnor U41019 (N_41019,N_40846,N_40700);
nand U41020 (N_41020,N_40714,N_40997);
xor U41021 (N_41021,N_40611,N_40680);
nand U41022 (N_41022,N_40742,N_40878);
or U41023 (N_41023,N_40564,N_40552);
or U41024 (N_41024,N_40877,N_40961);
xor U41025 (N_41025,N_40529,N_40746);
xor U41026 (N_41026,N_40968,N_40546);
xor U41027 (N_41027,N_40837,N_40644);
nand U41028 (N_41028,N_40696,N_40867);
xnor U41029 (N_41029,N_40737,N_40951);
and U41030 (N_41030,N_40610,N_40549);
nand U41031 (N_41031,N_40632,N_40864);
nor U41032 (N_41032,N_40634,N_40576);
nand U41033 (N_41033,N_40749,N_40729);
and U41034 (N_41034,N_40776,N_40606);
nor U41035 (N_41035,N_40883,N_40915);
or U41036 (N_41036,N_40833,N_40684);
nand U41037 (N_41037,N_40592,N_40822);
nand U41038 (N_41038,N_40741,N_40624);
xnor U41039 (N_41039,N_40526,N_40586);
and U41040 (N_41040,N_40676,N_40618);
nor U41041 (N_41041,N_40510,N_40779);
and U41042 (N_41042,N_40902,N_40687);
nand U41043 (N_41043,N_40970,N_40809);
or U41044 (N_41044,N_40555,N_40752);
and U41045 (N_41045,N_40988,N_40958);
or U41046 (N_41046,N_40842,N_40585);
nand U41047 (N_41047,N_40795,N_40971);
nand U41048 (N_41048,N_40732,N_40685);
nand U41049 (N_41049,N_40995,N_40792);
nor U41050 (N_41050,N_40747,N_40571);
nor U41051 (N_41051,N_40659,N_40782);
and U41052 (N_41052,N_40879,N_40553);
and U41053 (N_41053,N_40872,N_40641);
or U41054 (N_41054,N_40565,N_40542);
nand U41055 (N_41055,N_40996,N_40853);
xnor U41056 (N_41056,N_40774,N_40717);
xnor U41057 (N_41057,N_40960,N_40731);
nand U41058 (N_41058,N_40893,N_40789);
xor U41059 (N_41059,N_40554,N_40914);
xor U41060 (N_41060,N_40568,N_40697);
xnor U41061 (N_41061,N_40537,N_40518);
xnor U41062 (N_41062,N_40969,N_40686);
or U41063 (N_41063,N_40578,N_40777);
nor U41064 (N_41064,N_40698,N_40723);
and U41065 (N_41065,N_40656,N_40938);
and U41066 (N_41066,N_40539,N_40658);
nor U41067 (N_41067,N_40620,N_40799);
nor U41068 (N_41068,N_40726,N_40859);
or U41069 (N_41069,N_40973,N_40875);
xor U41070 (N_41070,N_40891,N_40817);
nor U41071 (N_41071,N_40811,N_40734);
and U41072 (N_41072,N_40798,N_40984);
or U41073 (N_41073,N_40922,N_40794);
and U41074 (N_41074,N_40652,N_40963);
or U41075 (N_41075,N_40534,N_40587);
or U41076 (N_41076,N_40524,N_40761);
and U41077 (N_41077,N_40679,N_40655);
nand U41078 (N_41078,N_40544,N_40807);
or U41079 (N_41079,N_40540,N_40716);
or U41080 (N_41080,N_40735,N_40849);
nand U41081 (N_41081,N_40695,N_40974);
or U41082 (N_41082,N_40959,N_40770);
and U41083 (N_41083,N_40919,N_40901);
or U41084 (N_41084,N_40943,N_40952);
and U41085 (N_41085,N_40885,N_40991);
nand U41086 (N_41086,N_40511,N_40981);
and U41087 (N_41087,N_40665,N_40574);
and U41088 (N_41088,N_40816,N_40953);
nor U41089 (N_41089,N_40913,N_40661);
xor U41090 (N_41090,N_40692,N_40517);
or U41091 (N_41091,N_40613,N_40506);
nor U41092 (N_41092,N_40603,N_40556);
nor U41093 (N_41093,N_40589,N_40593);
nor U41094 (N_41094,N_40688,N_40616);
and U41095 (N_41095,N_40630,N_40625);
nand U41096 (N_41096,N_40845,N_40850);
nor U41097 (N_41097,N_40608,N_40775);
nor U41098 (N_41098,N_40813,N_40824);
nor U41099 (N_41099,N_40828,N_40886);
nand U41100 (N_41100,N_40595,N_40590);
and U41101 (N_41101,N_40762,N_40609);
nand U41102 (N_41102,N_40651,N_40797);
xnor U41103 (N_41103,N_40711,N_40965);
nand U41104 (N_41104,N_40884,N_40989);
nand U41105 (N_41105,N_40986,N_40523);
xor U41106 (N_41106,N_40823,N_40636);
and U41107 (N_41107,N_40838,N_40990);
xnor U41108 (N_41108,N_40583,N_40946);
or U41109 (N_41109,N_40964,N_40821);
or U41110 (N_41110,N_40619,N_40721);
nand U41111 (N_41111,N_40667,N_40892);
nand U41112 (N_41112,N_40736,N_40547);
nand U41113 (N_41113,N_40707,N_40623);
nand U41114 (N_41114,N_40681,N_40559);
and U41115 (N_41115,N_40844,N_40934);
nand U41116 (N_41116,N_40784,N_40600);
xor U41117 (N_41117,N_40785,N_40643);
nand U41118 (N_41118,N_40500,N_40814);
nor U41119 (N_41119,N_40670,N_40504);
and U41120 (N_41120,N_40803,N_40501);
and U41121 (N_41121,N_40648,N_40710);
xor U41122 (N_41122,N_40631,N_40724);
xor U41123 (N_41123,N_40704,N_40855);
and U41124 (N_41124,N_40744,N_40771);
and U41125 (N_41125,N_40992,N_40614);
nand U41126 (N_41126,N_40808,N_40834);
nand U41127 (N_41127,N_40725,N_40905);
and U41128 (N_41128,N_40873,N_40532);
xnor U41129 (N_41129,N_40513,N_40733);
nor U41130 (N_41130,N_40745,N_40617);
and U41131 (N_41131,N_40750,N_40701);
xor U41132 (N_41132,N_40982,N_40548);
xor U41133 (N_41133,N_40773,N_40929);
nor U41134 (N_41134,N_40760,N_40691);
xnor U41135 (N_41135,N_40512,N_40694);
or U41136 (N_41136,N_40503,N_40932);
nand U41137 (N_41137,N_40581,N_40566);
and U41138 (N_41138,N_40507,N_40543);
nand U41139 (N_41139,N_40979,N_40975);
xnor U41140 (N_41140,N_40930,N_40881);
nand U41141 (N_41141,N_40836,N_40640);
nand U41142 (N_41142,N_40847,N_40928);
or U41143 (N_41143,N_40753,N_40604);
or U41144 (N_41144,N_40718,N_40527);
or U41145 (N_41145,N_40525,N_40588);
nor U41146 (N_41146,N_40856,N_40528);
or U41147 (N_41147,N_40839,N_40682);
or U41148 (N_41148,N_40861,N_40865);
xor U41149 (N_41149,N_40976,N_40740);
nand U41150 (N_41150,N_40728,N_40629);
and U41151 (N_41151,N_40896,N_40805);
or U41152 (N_41152,N_40787,N_40545);
or U41153 (N_41153,N_40906,N_40806);
nor U41154 (N_41154,N_40947,N_40646);
nor U41155 (N_41155,N_40825,N_40759);
nand U41156 (N_41156,N_40597,N_40582);
or U41157 (N_41157,N_40739,N_40763);
xnor U41158 (N_41158,N_40622,N_40927);
and U41159 (N_41159,N_40780,N_40521);
and U41160 (N_41160,N_40942,N_40920);
nor U41161 (N_41161,N_40921,N_40888);
or U41162 (N_41162,N_40854,N_40520);
nand U41163 (N_41163,N_40756,N_40820);
or U41164 (N_41164,N_40508,N_40857);
nor U41165 (N_41165,N_40898,N_40933);
xnor U41166 (N_41166,N_40899,N_40638);
xnor U41167 (N_41167,N_40669,N_40832);
xnor U41168 (N_41168,N_40751,N_40829);
or U41169 (N_41169,N_40730,N_40781);
xor U41170 (N_41170,N_40944,N_40972);
nand U41171 (N_41171,N_40866,N_40900);
and U41172 (N_41172,N_40563,N_40802);
nor U41173 (N_41173,N_40871,N_40666);
and U41174 (N_41174,N_40599,N_40674);
or U41175 (N_41175,N_40719,N_40675);
nand U41176 (N_41176,N_40598,N_40840);
or U41177 (N_41177,N_40931,N_40573);
nand U41178 (N_41178,N_40580,N_40936);
or U41179 (N_41179,N_40572,N_40671);
or U41180 (N_41180,N_40502,N_40908);
and U41181 (N_41181,N_40967,N_40673);
and U41182 (N_41182,N_40690,N_40509);
or U41183 (N_41183,N_40577,N_40815);
nand U41184 (N_41184,N_40705,N_40767);
and U41185 (N_41185,N_40800,N_40678);
nand U41186 (N_41186,N_40764,N_40607);
nand U41187 (N_41187,N_40627,N_40538);
and U41188 (N_41188,N_40657,N_40560);
and U41189 (N_41189,N_40912,N_40999);
xnor U41190 (N_41190,N_40870,N_40765);
or U41191 (N_41191,N_40505,N_40708);
or U41192 (N_41192,N_40950,N_40649);
and U41193 (N_41193,N_40858,N_40615);
nand U41194 (N_41194,N_40664,N_40635);
nand U41195 (N_41195,N_40584,N_40575);
nand U41196 (N_41196,N_40703,N_40949);
nor U41197 (N_41197,N_40876,N_40917);
nand U41198 (N_41198,N_40935,N_40647);
xnor U41199 (N_41199,N_40812,N_40907);
nor U41200 (N_41200,N_40993,N_40956);
nor U41201 (N_41201,N_40754,N_40522);
or U41202 (N_41202,N_40874,N_40755);
nand U41203 (N_41203,N_40897,N_40924);
xor U41204 (N_41204,N_40772,N_40769);
or U41205 (N_41205,N_40962,N_40804);
xnor U41206 (N_41206,N_40910,N_40994);
nand U41207 (N_41207,N_40596,N_40660);
and U41208 (N_41208,N_40957,N_40925);
nor U41209 (N_41209,N_40639,N_40841);
and U41210 (N_41210,N_40904,N_40766);
nor U41211 (N_41211,N_40557,N_40830);
and U41212 (N_41212,N_40668,N_40954);
nor U41213 (N_41213,N_40550,N_40757);
nand U41214 (N_41214,N_40980,N_40535);
nand U41215 (N_41215,N_40848,N_40778);
and U41216 (N_41216,N_40713,N_40653);
nor U41217 (N_41217,N_40727,N_40791);
or U41218 (N_41218,N_40743,N_40890);
nor U41219 (N_41219,N_40793,N_40783);
and U41220 (N_41220,N_40862,N_40633);
xnor U41221 (N_41221,N_40662,N_40768);
and U41222 (N_41222,N_40955,N_40851);
nand U41223 (N_41223,N_40672,N_40530);
nor U41224 (N_41224,N_40786,N_40923);
xnor U41225 (N_41225,N_40693,N_40868);
nor U41226 (N_41226,N_40810,N_40916);
xnor U41227 (N_41227,N_40796,N_40966);
nand U41228 (N_41228,N_40940,N_40602);
or U41229 (N_41229,N_40516,N_40562);
nor U41230 (N_41230,N_40738,N_40835);
xnor U41231 (N_41231,N_40987,N_40558);
and U41232 (N_41232,N_40985,N_40831);
xor U41233 (N_41233,N_40637,N_40880);
nor U41234 (N_41234,N_40712,N_40720);
or U41235 (N_41235,N_40843,N_40945);
nand U41236 (N_41236,N_40541,N_40860);
xor U41237 (N_41237,N_40663,N_40612);
nand U41238 (N_41238,N_40889,N_40748);
or U41239 (N_41239,N_40702,N_40561);
nand U41240 (N_41240,N_40514,N_40699);
or U41241 (N_41241,N_40852,N_40801);
and U41242 (N_41242,N_40909,N_40689);
nand U41243 (N_41243,N_40911,N_40819);
nand U41244 (N_41244,N_40863,N_40903);
and U41245 (N_41245,N_40887,N_40536);
nand U41246 (N_41246,N_40826,N_40926);
or U41247 (N_41247,N_40894,N_40531);
or U41248 (N_41248,N_40818,N_40579);
and U41249 (N_41249,N_40918,N_40895);
nand U41250 (N_41250,N_40517,N_40640);
and U41251 (N_41251,N_40801,N_40892);
nand U41252 (N_41252,N_40640,N_40724);
or U41253 (N_41253,N_40793,N_40557);
nor U41254 (N_41254,N_40816,N_40569);
xor U41255 (N_41255,N_40598,N_40761);
nand U41256 (N_41256,N_40579,N_40711);
nand U41257 (N_41257,N_40595,N_40970);
nor U41258 (N_41258,N_40616,N_40951);
and U41259 (N_41259,N_40912,N_40879);
or U41260 (N_41260,N_40897,N_40908);
nand U41261 (N_41261,N_40962,N_40996);
xor U41262 (N_41262,N_40931,N_40732);
xor U41263 (N_41263,N_40909,N_40991);
and U41264 (N_41264,N_40603,N_40989);
nand U41265 (N_41265,N_40512,N_40517);
nor U41266 (N_41266,N_40856,N_40861);
nor U41267 (N_41267,N_40964,N_40931);
and U41268 (N_41268,N_40806,N_40715);
nand U41269 (N_41269,N_40802,N_40531);
xor U41270 (N_41270,N_40877,N_40829);
nand U41271 (N_41271,N_40635,N_40782);
xnor U41272 (N_41272,N_40987,N_40584);
xnor U41273 (N_41273,N_40777,N_40600);
xor U41274 (N_41274,N_40706,N_40806);
nand U41275 (N_41275,N_40617,N_40826);
nor U41276 (N_41276,N_40553,N_40599);
xnor U41277 (N_41277,N_40550,N_40745);
and U41278 (N_41278,N_40824,N_40564);
xnor U41279 (N_41279,N_40982,N_40557);
or U41280 (N_41280,N_40801,N_40555);
or U41281 (N_41281,N_40877,N_40633);
nand U41282 (N_41282,N_40566,N_40892);
xnor U41283 (N_41283,N_40836,N_40502);
or U41284 (N_41284,N_40821,N_40797);
nand U41285 (N_41285,N_40954,N_40842);
xnor U41286 (N_41286,N_40729,N_40747);
nor U41287 (N_41287,N_40761,N_40591);
or U41288 (N_41288,N_40895,N_40849);
nor U41289 (N_41289,N_40896,N_40984);
or U41290 (N_41290,N_40925,N_40672);
and U41291 (N_41291,N_40782,N_40758);
nor U41292 (N_41292,N_40641,N_40822);
or U41293 (N_41293,N_40566,N_40558);
or U41294 (N_41294,N_40959,N_40845);
nor U41295 (N_41295,N_40989,N_40637);
nand U41296 (N_41296,N_40726,N_40705);
nor U41297 (N_41297,N_40556,N_40593);
and U41298 (N_41298,N_40808,N_40830);
xor U41299 (N_41299,N_40670,N_40956);
or U41300 (N_41300,N_40943,N_40826);
and U41301 (N_41301,N_40815,N_40682);
xor U41302 (N_41302,N_40907,N_40702);
and U41303 (N_41303,N_40623,N_40580);
or U41304 (N_41304,N_40640,N_40951);
and U41305 (N_41305,N_40742,N_40847);
or U41306 (N_41306,N_40687,N_40554);
nor U41307 (N_41307,N_40806,N_40591);
and U41308 (N_41308,N_40714,N_40851);
nor U41309 (N_41309,N_40893,N_40751);
or U41310 (N_41310,N_40764,N_40916);
xor U41311 (N_41311,N_40571,N_40874);
nor U41312 (N_41312,N_40674,N_40590);
xor U41313 (N_41313,N_40567,N_40884);
nand U41314 (N_41314,N_40932,N_40593);
nor U41315 (N_41315,N_40890,N_40632);
xor U41316 (N_41316,N_40515,N_40590);
or U41317 (N_41317,N_40937,N_40620);
and U41318 (N_41318,N_40829,N_40644);
or U41319 (N_41319,N_40810,N_40726);
or U41320 (N_41320,N_40882,N_40890);
nand U41321 (N_41321,N_40928,N_40961);
and U41322 (N_41322,N_40510,N_40731);
and U41323 (N_41323,N_40534,N_40890);
nor U41324 (N_41324,N_40520,N_40959);
xnor U41325 (N_41325,N_40989,N_40924);
xnor U41326 (N_41326,N_40535,N_40611);
nand U41327 (N_41327,N_40524,N_40657);
nor U41328 (N_41328,N_40792,N_40603);
nor U41329 (N_41329,N_40528,N_40702);
or U41330 (N_41330,N_40980,N_40578);
xor U41331 (N_41331,N_40828,N_40647);
or U41332 (N_41332,N_40976,N_40818);
and U41333 (N_41333,N_40542,N_40573);
nand U41334 (N_41334,N_40839,N_40571);
nor U41335 (N_41335,N_40584,N_40843);
and U41336 (N_41336,N_40595,N_40784);
nor U41337 (N_41337,N_40981,N_40999);
nor U41338 (N_41338,N_40772,N_40786);
and U41339 (N_41339,N_40975,N_40545);
xor U41340 (N_41340,N_40534,N_40640);
nand U41341 (N_41341,N_40500,N_40903);
nand U41342 (N_41342,N_40770,N_40657);
and U41343 (N_41343,N_40755,N_40549);
and U41344 (N_41344,N_40505,N_40862);
nand U41345 (N_41345,N_40826,N_40705);
and U41346 (N_41346,N_40599,N_40676);
xor U41347 (N_41347,N_40557,N_40973);
and U41348 (N_41348,N_40557,N_40910);
and U41349 (N_41349,N_40539,N_40779);
nand U41350 (N_41350,N_40941,N_40961);
and U41351 (N_41351,N_40753,N_40711);
nor U41352 (N_41352,N_40934,N_40614);
or U41353 (N_41353,N_40612,N_40883);
and U41354 (N_41354,N_40808,N_40975);
nor U41355 (N_41355,N_40667,N_40525);
or U41356 (N_41356,N_40717,N_40545);
xnor U41357 (N_41357,N_40917,N_40991);
nor U41358 (N_41358,N_40544,N_40974);
nor U41359 (N_41359,N_40635,N_40559);
nor U41360 (N_41360,N_40722,N_40527);
xnor U41361 (N_41361,N_40608,N_40999);
xor U41362 (N_41362,N_40789,N_40690);
and U41363 (N_41363,N_40680,N_40689);
and U41364 (N_41364,N_40971,N_40564);
and U41365 (N_41365,N_40937,N_40969);
or U41366 (N_41366,N_40822,N_40808);
and U41367 (N_41367,N_40638,N_40826);
nand U41368 (N_41368,N_40617,N_40647);
xor U41369 (N_41369,N_40592,N_40559);
and U41370 (N_41370,N_40971,N_40551);
or U41371 (N_41371,N_40875,N_40611);
xor U41372 (N_41372,N_40673,N_40793);
nand U41373 (N_41373,N_40597,N_40645);
xor U41374 (N_41374,N_40975,N_40980);
nand U41375 (N_41375,N_40980,N_40722);
xor U41376 (N_41376,N_40529,N_40950);
nand U41377 (N_41377,N_40767,N_40879);
nor U41378 (N_41378,N_40616,N_40690);
nor U41379 (N_41379,N_40574,N_40632);
nand U41380 (N_41380,N_40640,N_40678);
nand U41381 (N_41381,N_40694,N_40908);
or U41382 (N_41382,N_40621,N_40915);
nand U41383 (N_41383,N_40966,N_40679);
or U41384 (N_41384,N_40877,N_40500);
xnor U41385 (N_41385,N_40808,N_40595);
nand U41386 (N_41386,N_40506,N_40866);
nor U41387 (N_41387,N_40906,N_40711);
and U41388 (N_41388,N_40585,N_40661);
nand U41389 (N_41389,N_40939,N_40858);
nand U41390 (N_41390,N_40651,N_40857);
nor U41391 (N_41391,N_40893,N_40728);
or U41392 (N_41392,N_40997,N_40585);
or U41393 (N_41393,N_40704,N_40927);
nand U41394 (N_41394,N_40798,N_40642);
and U41395 (N_41395,N_40575,N_40681);
and U41396 (N_41396,N_40552,N_40911);
and U41397 (N_41397,N_40845,N_40862);
and U41398 (N_41398,N_40643,N_40911);
and U41399 (N_41399,N_40977,N_40525);
and U41400 (N_41400,N_40835,N_40971);
xnor U41401 (N_41401,N_40578,N_40935);
nor U41402 (N_41402,N_40893,N_40509);
xnor U41403 (N_41403,N_40563,N_40770);
nand U41404 (N_41404,N_40856,N_40730);
or U41405 (N_41405,N_40866,N_40694);
nor U41406 (N_41406,N_40712,N_40895);
or U41407 (N_41407,N_40704,N_40830);
nand U41408 (N_41408,N_40869,N_40832);
nand U41409 (N_41409,N_40911,N_40886);
xnor U41410 (N_41410,N_40650,N_40810);
or U41411 (N_41411,N_40977,N_40513);
xnor U41412 (N_41412,N_40924,N_40976);
nand U41413 (N_41413,N_40809,N_40751);
xnor U41414 (N_41414,N_40934,N_40824);
nor U41415 (N_41415,N_40572,N_40863);
and U41416 (N_41416,N_40566,N_40924);
nand U41417 (N_41417,N_40716,N_40573);
nor U41418 (N_41418,N_40944,N_40507);
xnor U41419 (N_41419,N_40879,N_40663);
nand U41420 (N_41420,N_40540,N_40740);
or U41421 (N_41421,N_40542,N_40523);
or U41422 (N_41422,N_40587,N_40773);
xor U41423 (N_41423,N_40803,N_40937);
xnor U41424 (N_41424,N_40990,N_40905);
and U41425 (N_41425,N_40858,N_40809);
and U41426 (N_41426,N_40909,N_40518);
or U41427 (N_41427,N_40967,N_40757);
or U41428 (N_41428,N_40792,N_40599);
xor U41429 (N_41429,N_40814,N_40578);
nor U41430 (N_41430,N_40513,N_40547);
and U41431 (N_41431,N_40766,N_40990);
nor U41432 (N_41432,N_40857,N_40859);
nor U41433 (N_41433,N_40853,N_40959);
xor U41434 (N_41434,N_40786,N_40865);
nor U41435 (N_41435,N_40646,N_40851);
nor U41436 (N_41436,N_40897,N_40836);
nor U41437 (N_41437,N_40950,N_40609);
nand U41438 (N_41438,N_40900,N_40751);
nor U41439 (N_41439,N_40584,N_40656);
xnor U41440 (N_41440,N_40684,N_40755);
and U41441 (N_41441,N_40801,N_40667);
nand U41442 (N_41442,N_40602,N_40671);
or U41443 (N_41443,N_40855,N_40944);
or U41444 (N_41444,N_40593,N_40945);
and U41445 (N_41445,N_40646,N_40815);
nand U41446 (N_41446,N_40800,N_40718);
xor U41447 (N_41447,N_40595,N_40540);
and U41448 (N_41448,N_40749,N_40642);
or U41449 (N_41449,N_40750,N_40666);
nand U41450 (N_41450,N_40623,N_40918);
xor U41451 (N_41451,N_40624,N_40857);
nand U41452 (N_41452,N_40778,N_40667);
or U41453 (N_41453,N_40736,N_40662);
and U41454 (N_41454,N_40925,N_40973);
nand U41455 (N_41455,N_40734,N_40747);
or U41456 (N_41456,N_40639,N_40629);
nand U41457 (N_41457,N_40739,N_40526);
or U41458 (N_41458,N_40530,N_40553);
nand U41459 (N_41459,N_40598,N_40970);
nand U41460 (N_41460,N_40732,N_40874);
xor U41461 (N_41461,N_40940,N_40699);
nand U41462 (N_41462,N_40543,N_40945);
nand U41463 (N_41463,N_40763,N_40717);
nor U41464 (N_41464,N_40610,N_40611);
or U41465 (N_41465,N_40902,N_40946);
nand U41466 (N_41466,N_40772,N_40917);
nand U41467 (N_41467,N_40930,N_40642);
nand U41468 (N_41468,N_40983,N_40539);
nand U41469 (N_41469,N_40843,N_40907);
nand U41470 (N_41470,N_40502,N_40703);
nor U41471 (N_41471,N_40841,N_40838);
nor U41472 (N_41472,N_40953,N_40646);
nor U41473 (N_41473,N_40677,N_40595);
nor U41474 (N_41474,N_40642,N_40564);
and U41475 (N_41475,N_40671,N_40576);
xor U41476 (N_41476,N_40663,N_40662);
nor U41477 (N_41477,N_40835,N_40876);
and U41478 (N_41478,N_40632,N_40812);
or U41479 (N_41479,N_40778,N_40723);
or U41480 (N_41480,N_40725,N_40622);
nor U41481 (N_41481,N_40999,N_40838);
or U41482 (N_41482,N_40809,N_40696);
xnor U41483 (N_41483,N_40720,N_40677);
nand U41484 (N_41484,N_40748,N_40536);
nor U41485 (N_41485,N_40918,N_40753);
and U41486 (N_41486,N_40970,N_40813);
and U41487 (N_41487,N_40686,N_40926);
nor U41488 (N_41488,N_40860,N_40803);
or U41489 (N_41489,N_40873,N_40817);
and U41490 (N_41490,N_40863,N_40911);
xor U41491 (N_41491,N_40866,N_40999);
nand U41492 (N_41492,N_40549,N_40970);
and U41493 (N_41493,N_40597,N_40563);
and U41494 (N_41494,N_40536,N_40835);
xnor U41495 (N_41495,N_40667,N_40580);
nor U41496 (N_41496,N_40928,N_40568);
xor U41497 (N_41497,N_40877,N_40786);
and U41498 (N_41498,N_40764,N_40902);
and U41499 (N_41499,N_40559,N_40940);
nor U41500 (N_41500,N_41470,N_41437);
nor U41501 (N_41501,N_41064,N_41364);
xor U41502 (N_41502,N_41233,N_41001);
or U41503 (N_41503,N_41319,N_41394);
nor U41504 (N_41504,N_41229,N_41373);
nor U41505 (N_41505,N_41215,N_41357);
nand U41506 (N_41506,N_41368,N_41492);
nand U41507 (N_41507,N_41339,N_41162);
and U41508 (N_41508,N_41268,N_41234);
xnor U41509 (N_41509,N_41487,N_41451);
xor U41510 (N_41510,N_41236,N_41243);
and U41511 (N_41511,N_41404,N_41214);
nand U41512 (N_41512,N_41167,N_41479);
nor U41513 (N_41513,N_41353,N_41189);
xor U41514 (N_41514,N_41021,N_41408);
nand U41515 (N_41515,N_41293,N_41129);
and U41516 (N_41516,N_41410,N_41178);
nand U41517 (N_41517,N_41332,N_41193);
nand U41518 (N_41518,N_41059,N_41011);
nand U41519 (N_41519,N_41484,N_41247);
nand U41520 (N_41520,N_41421,N_41081);
xnor U41521 (N_41521,N_41005,N_41305);
nor U41522 (N_41522,N_41087,N_41209);
xnor U41523 (N_41523,N_41086,N_41230);
nor U41524 (N_41524,N_41418,N_41388);
and U41525 (N_41525,N_41221,N_41448);
nor U41526 (N_41526,N_41267,N_41093);
nand U41527 (N_41527,N_41100,N_41245);
nor U41528 (N_41528,N_41184,N_41442);
nand U41529 (N_41529,N_41401,N_41318);
xnor U41530 (N_41530,N_41058,N_41226);
nor U41531 (N_41531,N_41483,N_41307);
nand U41532 (N_41532,N_41458,N_41375);
xor U41533 (N_41533,N_41037,N_41459);
xnor U41534 (N_41534,N_41420,N_41187);
nor U41535 (N_41535,N_41258,N_41083);
nor U41536 (N_41536,N_41429,N_41321);
xnor U41537 (N_41537,N_41118,N_41140);
nor U41538 (N_41538,N_41407,N_41195);
and U41539 (N_41539,N_41128,N_41327);
nor U41540 (N_41540,N_41350,N_41445);
and U41541 (N_41541,N_41467,N_41428);
nor U41542 (N_41542,N_41281,N_41109);
xnor U41543 (N_41543,N_41228,N_41395);
and U41544 (N_41544,N_41126,N_41406);
xnor U41545 (N_41545,N_41251,N_41491);
nor U41546 (N_41546,N_41453,N_41485);
or U41547 (N_41547,N_41155,N_41272);
xnor U41548 (N_41548,N_41134,N_41440);
nor U41549 (N_41549,N_41363,N_41117);
nand U41550 (N_41550,N_41441,N_41029);
or U41551 (N_41551,N_41146,N_41351);
or U41552 (N_41552,N_41142,N_41066);
nand U41553 (N_41553,N_41466,N_41259);
xnor U41554 (N_41554,N_41302,N_41360);
xor U41555 (N_41555,N_41220,N_41172);
and U41556 (N_41556,N_41211,N_41174);
nor U41557 (N_41557,N_41398,N_41417);
and U41558 (N_41558,N_41053,N_41004);
or U41559 (N_41559,N_41488,N_41284);
nor U41560 (N_41560,N_41385,N_41337);
nor U41561 (N_41561,N_41113,N_41106);
xor U41562 (N_41562,N_41208,N_41182);
nand U41563 (N_41563,N_41238,N_41099);
xnor U41564 (N_41564,N_41008,N_41468);
xor U41565 (N_41565,N_41203,N_41108);
nand U41566 (N_41566,N_41256,N_41196);
nor U41567 (N_41567,N_41202,N_41124);
nor U41568 (N_41568,N_41443,N_41012);
and U41569 (N_41569,N_41380,N_41300);
xor U41570 (N_41570,N_41206,N_41063);
xor U41571 (N_41571,N_41003,N_41378);
or U41572 (N_41572,N_41158,N_41347);
or U41573 (N_41573,N_41323,N_41292);
nor U41574 (N_41574,N_41069,N_41250);
nor U41575 (N_41575,N_41370,N_41263);
nor U41576 (N_41576,N_41160,N_41377);
and U41577 (N_41577,N_41316,N_41328);
xor U41578 (N_41578,N_41496,N_41057);
xor U41579 (N_41579,N_41463,N_41200);
and U41580 (N_41580,N_41077,N_41120);
and U41581 (N_41581,N_41369,N_41179);
and U41582 (N_41582,N_41153,N_41315);
nand U41583 (N_41583,N_41168,N_41449);
xor U41584 (N_41584,N_41218,N_41232);
nor U41585 (N_41585,N_41414,N_41499);
nor U41586 (N_41586,N_41283,N_41255);
nand U41587 (N_41587,N_41006,N_41047);
nand U41588 (N_41588,N_41102,N_41030);
or U41589 (N_41589,N_41405,N_41239);
or U41590 (N_41590,N_41469,N_41461);
and U41591 (N_41591,N_41186,N_41169);
xor U41592 (N_41592,N_41345,N_41205);
xnor U41593 (N_41593,N_41489,N_41291);
xor U41594 (N_41594,N_41391,N_41055);
and U41595 (N_41595,N_41389,N_41261);
and U41596 (N_41596,N_41139,N_41240);
or U41597 (N_41597,N_41144,N_41269);
xor U41598 (N_41598,N_41254,N_41276);
and U41599 (N_41599,N_41010,N_41076);
nor U41600 (N_41600,N_41159,N_41136);
xnor U41601 (N_41601,N_41403,N_41040);
or U41602 (N_41602,N_41143,N_41296);
nor U41603 (N_41603,N_41450,N_41181);
nor U41604 (N_41604,N_41114,N_41304);
nand U41605 (N_41605,N_41299,N_41311);
or U41606 (N_41606,N_41456,N_41257);
xor U41607 (N_41607,N_41183,N_41045);
nand U41608 (N_41608,N_41265,N_41361);
nor U41609 (N_41609,N_41138,N_41065);
nor U41610 (N_41610,N_41016,N_41125);
xor U41611 (N_41611,N_41036,N_41101);
and U41612 (N_41612,N_41435,N_41362);
nor U41613 (N_41613,N_41018,N_41297);
nand U41614 (N_41614,N_41325,N_41156);
nand U41615 (N_41615,N_41048,N_41349);
nor U41616 (N_41616,N_41049,N_41032);
nand U41617 (N_41617,N_41041,N_41175);
nand U41618 (N_41618,N_41022,N_41014);
and U41619 (N_41619,N_41348,N_41072);
nand U41620 (N_41620,N_41285,N_41324);
or U41621 (N_41621,N_41460,N_41434);
or U41622 (N_41622,N_41400,N_41015);
and U41623 (N_41623,N_41201,N_41024);
and U41624 (N_41624,N_41116,N_41366);
and U41625 (N_41625,N_41260,N_41397);
and U41626 (N_41626,N_41242,N_41330);
nand U41627 (N_41627,N_41147,N_41294);
or U41628 (N_41628,N_41079,N_41062);
and U41629 (N_41629,N_41473,N_41249);
or U41630 (N_41630,N_41413,N_41080);
xnor U41631 (N_41631,N_41344,N_41033);
and U41632 (N_41632,N_41303,N_41137);
nand U41633 (N_41633,N_41280,N_41119);
nand U41634 (N_41634,N_41198,N_41402);
xnor U41635 (N_41635,N_41122,N_41490);
nor U41636 (N_41636,N_41068,N_41390);
or U41637 (N_41637,N_41223,N_41170);
xnor U41638 (N_41638,N_41415,N_41084);
or U41639 (N_41639,N_41056,N_41498);
nor U41640 (N_41640,N_41180,N_41075);
nor U41641 (N_41641,N_41096,N_41384);
xor U41642 (N_41642,N_41043,N_41431);
nor U41643 (N_41643,N_41224,N_41409);
or U41644 (N_41644,N_41246,N_41145);
and U41645 (N_41645,N_41191,N_41071);
nand U41646 (N_41646,N_41392,N_41475);
xor U41647 (N_41647,N_41343,N_41210);
or U41648 (N_41648,N_41301,N_41141);
xor U41649 (N_41649,N_41161,N_41121);
nor U41650 (N_41650,N_41322,N_41481);
or U41651 (N_41651,N_41457,N_41264);
or U41652 (N_41652,N_41217,N_41165);
and U41653 (N_41653,N_41219,N_41237);
xor U41654 (N_41654,N_41317,N_41314);
xnor U41655 (N_41655,N_41090,N_41038);
or U41656 (N_41656,N_41358,N_41354);
nand U41657 (N_41657,N_41082,N_41110);
nor U41658 (N_41658,N_41341,N_41497);
and U41659 (N_41659,N_41157,N_41430);
or U41660 (N_41660,N_41042,N_41149);
xnor U41661 (N_41661,N_41286,N_41235);
and U41662 (N_41662,N_41130,N_41356);
and U41663 (N_41663,N_41287,N_41477);
nor U41664 (N_41664,N_41288,N_41188);
or U41665 (N_41665,N_41070,N_41098);
xor U41666 (N_41666,N_41371,N_41054);
xor U41667 (N_41667,N_41306,N_41432);
or U41668 (N_41668,N_41131,N_41416);
xnor U41669 (N_41669,N_41212,N_41009);
and U41670 (N_41670,N_41073,N_41455);
and U41671 (N_41671,N_41092,N_41094);
nor U41672 (N_41672,N_41424,N_41173);
xnor U41673 (N_41673,N_41277,N_41381);
nor U41674 (N_41674,N_41383,N_41355);
xor U41675 (N_41675,N_41061,N_41034);
and U41676 (N_41676,N_41279,N_41197);
nor U41677 (N_41677,N_41309,N_41225);
xnor U41678 (N_41678,N_41091,N_41308);
and U41679 (N_41679,N_41436,N_41213);
or U41680 (N_41680,N_41493,N_41231);
nor U41681 (N_41681,N_41089,N_41227);
xor U41682 (N_41682,N_41482,N_41019);
nand U41683 (N_41683,N_41310,N_41273);
nor U41684 (N_41684,N_41000,N_41326);
and U41685 (N_41685,N_41152,N_41123);
and U41686 (N_41686,N_41386,N_41433);
nand U41687 (N_41687,N_41190,N_41244);
nand U41688 (N_41688,N_41039,N_41035);
xor U41689 (N_41689,N_41185,N_41447);
nand U41690 (N_41690,N_41248,N_41338);
nand U41691 (N_41691,N_41112,N_41336);
xnor U41692 (N_41692,N_41177,N_41204);
xnor U41693 (N_41693,N_41312,N_41411);
or U41694 (N_41694,N_41111,N_41271);
or U41695 (N_41695,N_41320,N_41164);
nand U41696 (N_41696,N_41444,N_41207);
xnor U41697 (N_41697,N_41060,N_41222);
nor U41698 (N_41698,N_41495,N_41046);
nor U41699 (N_41699,N_41333,N_41331);
xor U41700 (N_41700,N_41472,N_41298);
nor U41701 (N_41701,N_41115,N_41253);
or U41702 (N_41702,N_41422,N_41199);
and U41703 (N_41703,N_41067,N_41027);
and U41704 (N_41704,N_41379,N_41266);
xor U41705 (N_41705,N_41278,N_41399);
nor U41706 (N_41706,N_41192,N_41166);
xor U41707 (N_41707,N_41252,N_41216);
nand U41708 (N_41708,N_41313,N_41270);
and U41709 (N_41709,N_41340,N_41132);
or U41710 (N_41710,N_41474,N_41154);
and U41711 (N_41711,N_41171,N_41013);
and U41712 (N_41712,N_41103,N_41088);
and U41713 (N_41713,N_41454,N_41023);
nand U41714 (N_41714,N_41026,N_41085);
or U41715 (N_41715,N_41097,N_41464);
nand U41716 (N_41716,N_41376,N_41241);
or U41717 (N_41717,N_41367,N_41439);
nor U41718 (N_41718,N_41150,N_41107);
and U41719 (N_41719,N_41105,N_41476);
nor U41720 (N_41720,N_41028,N_41274);
xor U41721 (N_41721,N_41352,N_41289);
nor U41722 (N_41722,N_41163,N_41486);
and U41723 (N_41723,N_41471,N_41044);
or U41724 (N_41724,N_41050,N_41412);
nand U41725 (N_41725,N_41020,N_41426);
or U41726 (N_41726,N_41478,N_41282);
nor U41727 (N_41727,N_41051,N_41382);
or U41728 (N_41728,N_41342,N_41295);
or U41729 (N_41729,N_41095,N_41127);
or U41730 (N_41730,N_41465,N_41151);
nand U41731 (N_41731,N_41133,N_41365);
and U41732 (N_41732,N_41275,N_41335);
nor U41733 (N_41733,N_41078,N_41194);
and U41734 (N_41734,N_41446,N_41462);
xnor U41735 (N_41735,N_41359,N_41176);
and U41736 (N_41736,N_41425,N_41427);
xor U41737 (N_41737,N_41346,N_41494);
nor U41738 (N_41738,N_41419,N_41031);
or U41739 (N_41739,N_41148,N_41396);
xor U41740 (N_41740,N_41423,N_41002);
xor U41741 (N_41741,N_41290,N_41374);
nand U41742 (N_41742,N_41135,N_41074);
xnor U41743 (N_41743,N_41387,N_41334);
or U41744 (N_41744,N_41052,N_41104);
nand U41745 (N_41745,N_41480,N_41017);
xnor U41746 (N_41746,N_41329,N_41438);
nand U41747 (N_41747,N_41393,N_41452);
xnor U41748 (N_41748,N_41007,N_41025);
nand U41749 (N_41749,N_41372,N_41262);
nand U41750 (N_41750,N_41371,N_41457);
nand U41751 (N_41751,N_41063,N_41386);
or U41752 (N_41752,N_41266,N_41311);
xnor U41753 (N_41753,N_41195,N_41218);
nor U41754 (N_41754,N_41288,N_41287);
xnor U41755 (N_41755,N_41424,N_41172);
nor U41756 (N_41756,N_41283,N_41186);
and U41757 (N_41757,N_41229,N_41184);
or U41758 (N_41758,N_41019,N_41418);
nand U41759 (N_41759,N_41436,N_41469);
and U41760 (N_41760,N_41370,N_41355);
xor U41761 (N_41761,N_41365,N_41271);
nor U41762 (N_41762,N_41434,N_41051);
xor U41763 (N_41763,N_41092,N_41242);
or U41764 (N_41764,N_41409,N_41447);
xor U41765 (N_41765,N_41225,N_41138);
nor U41766 (N_41766,N_41299,N_41079);
nand U41767 (N_41767,N_41133,N_41220);
xor U41768 (N_41768,N_41389,N_41430);
nor U41769 (N_41769,N_41095,N_41111);
nor U41770 (N_41770,N_41143,N_41085);
or U41771 (N_41771,N_41468,N_41372);
nand U41772 (N_41772,N_41003,N_41288);
or U41773 (N_41773,N_41071,N_41337);
nand U41774 (N_41774,N_41417,N_41345);
nor U41775 (N_41775,N_41468,N_41152);
nand U41776 (N_41776,N_41129,N_41047);
and U41777 (N_41777,N_41200,N_41480);
nor U41778 (N_41778,N_41485,N_41114);
and U41779 (N_41779,N_41264,N_41190);
nor U41780 (N_41780,N_41362,N_41254);
xnor U41781 (N_41781,N_41331,N_41348);
xnor U41782 (N_41782,N_41054,N_41272);
xor U41783 (N_41783,N_41077,N_41116);
xnor U41784 (N_41784,N_41029,N_41493);
or U41785 (N_41785,N_41389,N_41314);
nor U41786 (N_41786,N_41008,N_41154);
or U41787 (N_41787,N_41368,N_41146);
xnor U41788 (N_41788,N_41002,N_41006);
and U41789 (N_41789,N_41058,N_41002);
and U41790 (N_41790,N_41391,N_41082);
or U41791 (N_41791,N_41054,N_41451);
or U41792 (N_41792,N_41357,N_41460);
or U41793 (N_41793,N_41486,N_41435);
xnor U41794 (N_41794,N_41409,N_41014);
nand U41795 (N_41795,N_41026,N_41379);
nand U41796 (N_41796,N_41206,N_41272);
or U41797 (N_41797,N_41223,N_41004);
nor U41798 (N_41798,N_41235,N_41417);
nor U41799 (N_41799,N_41425,N_41305);
nand U41800 (N_41800,N_41296,N_41298);
nand U41801 (N_41801,N_41403,N_41370);
or U41802 (N_41802,N_41436,N_41109);
and U41803 (N_41803,N_41092,N_41464);
nor U41804 (N_41804,N_41041,N_41075);
or U41805 (N_41805,N_41174,N_41341);
xnor U41806 (N_41806,N_41248,N_41190);
and U41807 (N_41807,N_41423,N_41026);
or U41808 (N_41808,N_41497,N_41178);
or U41809 (N_41809,N_41187,N_41492);
or U41810 (N_41810,N_41308,N_41331);
nand U41811 (N_41811,N_41227,N_41180);
nand U41812 (N_41812,N_41432,N_41371);
nor U41813 (N_41813,N_41008,N_41409);
and U41814 (N_41814,N_41283,N_41084);
nand U41815 (N_41815,N_41444,N_41042);
and U41816 (N_41816,N_41128,N_41291);
nand U41817 (N_41817,N_41112,N_41005);
and U41818 (N_41818,N_41117,N_41448);
nor U41819 (N_41819,N_41016,N_41433);
or U41820 (N_41820,N_41330,N_41282);
and U41821 (N_41821,N_41217,N_41096);
nor U41822 (N_41822,N_41322,N_41433);
or U41823 (N_41823,N_41131,N_41211);
xnor U41824 (N_41824,N_41195,N_41215);
nor U41825 (N_41825,N_41282,N_41186);
nand U41826 (N_41826,N_41460,N_41334);
xnor U41827 (N_41827,N_41296,N_41263);
and U41828 (N_41828,N_41000,N_41247);
and U41829 (N_41829,N_41055,N_41240);
and U41830 (N_41830,N_41179,N_41475);
xor U41831 (N_41831,N_41414,N_41138);
or U41832 (N_41832,N_41318,N_41263);
xnor U41833 (N_41833,N_41401,N_41093);
nand U41834 (N_41834,N_41455,N_41117);
and U41835 (N_41835,N_41137,N_41441);
and U41836 (N_41836,N_41417,N_41219);
xor U41837 (N_41837,N_41397,N_41272);
xor U41838 (N_41838,N_41494,N_41388);
xnor U41839 (N_41839,N_41274,N_41408);
and U41840 (N_41840,N_41048,N_41420);
or U41841 (N_41841,N_41390,N_41347);
and U41842 (N_41842,N_41027,N_41449);
nand U41843 (N_41843,N_41301,N_41409);
xor U41844 (N_41844,N_41459,N_41405);
or U41845 (N_41845,N_41350,N_41344);
xor U41846 (N_41846,N_41310,N_41271);
nand U41847 (N_41847,N_41406,N_41455);
nand U41848 (N_41848,N_41465,N_41338);
and U41849 (N_41849,N_41125,N_41127);
nand U41850 (N_41850,N_41204,N_41255);
xor U41851 (N_41851,N_41168,N_41268);
nand U41852 (N_41852,N_41174,N_41266);
nand U41853 (N_41853,N_41129,N_41318);
and U41854 (N_41854,N_41337,N_41246);
and U41855 (N_41855,N_41116,N_41430);
and U41856 (N_41856,N_41256,N_41057);
nor U41857 (N_41857,N_41162,N_41216);
nand U41858 (N_41858,N_41452,N_41396);
and U41859 (N_41859,N_41086,N_41276);
xor U41860 (N_41860,N_41042,N_41361);
or U41861 (N_41861,N_41240,N_41062);
or U41862 (N_41862,N_41248,N_41160);
xnor U41863 (N_41863,N_41289,N_41229);
and U41864 (N_41864,N_41229,N_41053);
or U41865 (N_41865,N_41215,N_41106);
and U41866 (N_41866,N_41334,N_41247);
nand U41867 (N_41867,N_41291,N_41072);
nor U41868 (N_41868,N_41336,N_41300);
nor U41869 (N_41869,N_41415,N_41483);
and U41870 (N_41870,N_41455,N_41150);
nand U41871 (N_41871,N_41191,N_41200);
nor U41872 (N_41872,N_41007,N_41385);
nor U41873 (N_41873,N_41305,N_41245);
xor U41874 (N_41874,N_41284,N_41134);
nand U41875 (N_41875,N_41342,N_41122);
nand U41876 (N_41876,N_41434,N_41278);
and U41877 (N_41877,N_41493,N_41124);
nand U41878 (N_41878,N_41132,N_41331);
nor U41879 (N_41879,N_41382,N_41462);
or U41880 (N_41880,N_41160,N_41279);
nand U41881 (N_41881,N_41056,N_41200);
xnor U41882 (N_41882,N_41443,N_41289);
and U41883 (N_41883,N_41473,N_41210);
xor U41884 (N_41884,N_41443,N_41048);
nor U41885 (N_41885,N_41423,N_41464);
or U41886 (N_41886,N_41375,N_41489);
nor U41887 (N_41887,N_41386,N_41067);
nor U41888 (N_41888,N_41064,N_41239);
xnor U41889 (N_41889,N_41455,N_41377);
and U41890 (N_41890,N_41499,N_41383);
or U41891 (N_41891,N_41496,N_41133);
nor U41892 (N_41892,N_41374,N_41402);
nor U41893 (N_41893,N_41392,N_41177);
nand U41894 (N_41894,N_41081,N_41390);
and U41895 (N_41895,N_41240,N_41470);
xnor U41896 (N_41896,N_41378,N_41065);
or U41897 (N_41897,N_41335,N_41296);
xor U41898 (N_41898,N_41033,N_41236);
xnor U41899 (N_41899,N_41298,N_41476);
or U41900 (N_41900,N_41432,N_41414);
and U41901 (N_41901,N_41111,N_41432);
xnor U41902 (N_41902,N_41129,N_41479);
nor U41903 (N_41903,N_41412,N_41496);
nand U41904 (N_41904,N_41372,N_41426);
and U41905 (N_41905,N_41472,N_41345);
nor U41906 (N_41906,N_41080,N_41448);
nor U41907 (N_41907,N_41458,N_41312);
or U41908 (N_41908,N_41145,N_41350);
nand U41909 (N_41909,N_41091,N_41255);
nand U41910 (N_41910,N_41192,N_41044);
xor U41911 (N_41911,N_41130,N_41015);
xor U41912 (N_41912,N_41304,N_41094);
or U41913 (N_41913,N_41437,N_41235);
xor U41914 (N_41914,N_41103,N_41420);
nor U41915 (N_41915,N_41089,N_41012);
and U41916 (N_41916,N_41133,N_41337);
or U41917 (N_41917,N_41123,N_41483);
and U41918 (N_41918,N_41057,N_41266);
nor U41919 (N_41919,N_41490,N_41418);
nor U41920 (N_41920,N_41322,N_41334);
or U41921 (N_41921,N_41448,N_41361);
nor U41922 (N_41922,N_41403,N_41382);
nor U41923 (N_41923,N_41482,N_41045);
or U41924 (N_41924,N_41272,N_41436);
nor U41925 (N_41925,N_41370,N_41458);
xor U41926 (N_41926,N_41022,N_41467);
and U41927 (N_41927,N_41213,N_41482);
or U41928 (N_41928,N_41286,N_41241);
nand U41929 (N_41929,N_41224,N_41119);
or U41930 (N_41930,N_41291,N_41286);
nand U41931 (N_41931,N_41268,N_41129);
nor U41932 (N_41932,N_41143,N_41209);
and U41933 (N_41933,N_41433,N_41259);
or U41934 (N_41934,N_41372,N_41438);
nand U41935 (N_41935,N_41001,N_41062);
xnor U41936 (N_41936,N_41209,N_41139);
and U41937 (N_41937,N_41336,N_41194);
xor U41938 (N_41938,N_41159,N_41486);
and U41939 (N_41939,N_41276,N_41321);
nand U41940 (N_41940,N_41058,N_41345);
nor U41941 (N_41941,N_41232,N_41035);
nand U41942 (N_41942,N_41218,N_41298);
xor U41943 (N_41943,N_41121,N_41200);
xor U41944 (N_41944,N_41324,N_41464);
nor U41945 (N_41945,N_41411,N_41058);
and U41946 (N_41946,N_41159,N_41330);
and U41947 (N_41947,N_41283,N_41444);
xnor U41948 (N_41948,N_41015,N_41191);
nand U41949 (N_41949,N_41372,N_41400);
nor U41950 (N_41950,N_41081,N_41208);
xor U41951 (N_41951,N_41049,N_41297);
or U41952 (N_41952,N_41401,N_41372);
nand U41953 (N_41953,N_41367,N_41141);
or U41954 (N_41954,N_41262,N_41475);
and U41955 (N_41955,N_41140,N_41185);
nor U41956 (N_41956,N_41112,N_41255);
nand U41957 (N_41957,N_41231,N_41138);
nor U41958 (N_41958,N_41336,N_41248);
or U41959 (N_41959,N_41218,N_41481);
nor U41960 (N_41960,N_41052,N_41441);
xnor U41961 (N_41961,N_41295,N_41206);
nor U41962 (N_41962,N_41007,N_41186);
nand U41963 (N_41963,N_41032,N_41345);
and U41964 (N_41964,N_41004,N_41015);
nor U41965 (N_41965,N_41182,N_41122);
nand U41966 (N_41966,N_41075,N_41069);
nor U41967 (N_41967,N_41406,N_41172);
and U41968 (N_41968,N_41214,N_41036);
nand U41969 (N_41969,N_41317,N_41276);
nor U41970 (N_41970,N_41000,N_41133);
xnor U41971 (N_41971,N_41372,N_41419);
xnor U41972 (N_41972,N_41320,N_41306);
nor U41973 (N_41973,N_41137,N_41180);
nand U41974 (N_41974,N_41370,N_41207);
nor U41975 (N_41975,N_41152,N_41139);
nor U41976 (N_41976,N_41002,N_41409);
nand U41977 (N_41977,N_41097,N_41368);
and U41978 (N_41978,N_41074,N_41451);
xor U41979 (N_41979,N_41178,N_41332);
or U41980 (N_41980,N_41103,N_41122);
and U41981 (N_41981,N_41275,N_41363);
nand U41982 (N_41982,N_41138,N_41284);
xnor U41983 (N_41983,N_41351,N_41323);
xnor U41984 (N_41984,N_41328,N_41330);
nor U41985 (N_41985,N_41110,N_41431);
xor U41986 (N_41986,N_41052,N_41210);
nor U41987 (N_41987,N_41145,N_41042);
or U41988 (N_41988,N_41236,N_41355);
nand U41989 (N_41989,N_41385,N_41070);
and U41990 (N_41990,N_41207,N_41423);
xnor U41991 (N_41991,N_41312,N_41262);
xnor U41992 (N_41992,N_41358,N_41363);
nor U41993 (N_41993,N_41432,N_41405);
or U41994 (N_41994,N_41111,N_41194);
nor U41995 (N_41995,N_41206,N_41056);
xnor U41996 (N_41996,N_41459,N_41290);
and U41997 (N_41997,N_41260,N_41121);
nor U41998 (N_41998,N_41392,N_41288);
or U41999 (N_41999,N_41203,N_41321);
and U42000 (N_42000,N_41988,N_41984);
nand U42001 (N_42001,N_41766,N_41667);
or U42002 (N_42002,N_41728,N_41790);
nor U42003 (N_42003,N_41929,N_41737);
or U42004 (N_42004,N_41755,N_41581);
xnor U42005 (N_42005,N_41877,N_41845);
xor U42006 (N_42006,N_41522,N_41865);
xor U42007 (N_42007,N_41926,N_41770);
nand U42008 (N_42008,N_41509,N_41889);
nor U42009 (N_42009,N_41527,N_41678);
nand U42010 (N_42010,N_41894,N_41746);
and U42011 (N_42011,N_41860,N_41679);
nor U42012 (N_42012,N_41725,N_41780);
nor U42013 (N_42013,N_41838,N_41973);
or U42014 (N_42014,N_41714,N_41673);
xnor U42015 (N_42015,N_41761,N_41918);
and U42016 (N_42016,N_41552,N_41551);
nor U42017 (N_42017,N_41597,N_41813);
nor U42018 (N_42018,N_41645,N_41979);
xnor U42019 (N_42019,N_41570,N_41966);
and U42020 (N_42020,N_41646,N_41594);
xnor U42021 (N_42021,N_41974,N_41821);
nand U42022 (N_42022,N_41914,N_41978);
nor U42023 (N_42023,N_41520,N_41639);
nor U42024 (N_42024,N_41716,N_41789);
and U42025 (N_42025,N_41818,N_41610);
xnor U42026 (N_42026,N_41642,N_41700);
or U42027 (N_42027,N_41738,N_41992);
or U42028 (N_42028,N_41618,N_41536);
xnor U42029 (N_42029,N_41593,N_41732);
nor U42030 (N_42030,N_41830,N_41874);
nand U42031 (N_42031,N_41945,N_41632);
nand U42032 (N_42032,N_41547,N_41799);
and U42033 (N_42033,N_41612,N_41924);
xnor U42034 (N_42034,N_41814,N_41649);
or U42035 (N_42035,N_41751,N_41694);
or U42036 (N_42036,N_41868,N_41937);
xor U42037 (N_42037,N_41827,N_41934);
nand U42038 (N_42038,N_41582,N_41604);
and U42039 (N_42039,N_41898,N_41505);
or U42040 (N_42040,N_41909,N_41895);
xor U42041 (N_42041,N_41638,N_41576);
or U42042 (N_42042,N_41983,N_41772);
xor U42043 (N_42043,N_41599,N_41788);
or U42044 (N_42044,N_41968,N_41869);
nand U42045 (N_42045,N_41670,N_41685);
nand U42046 (N_42046,N_41933,N_41990);
xor U42047 (N_42047,N_41574,N_41923);
and U42048 (N_42048,N_41995,N_41785);
and U42049 (N_42049,N_41784,N_41840);
xnor U42050 (N_42050,N_41952,N_41820);
xor U42051 (N_42051,N_41857,N_41598);
and U42052 (N_42052,N_41851,N_41702);
nand U42053 (N_42053,N_41504,N_41880);
nand U42054 (N_42054,N_41940,N_41502);
and U42055 (N_42055,N_41807,N_41873);
nand U42056 (N_42056,N_41546,N_41579);
nor U42057 (N_42057,N_41887,N_41861);
xnor U42058 (N_42058,N_41657,N_41805);
nand U42059 (N_42059,N_41796,N_41613);
nor U42060 (N_42060,N_41823,N_41743);
and U42061 (N_42061,N_41883,N_41519);
nand U42062 (N_42062,N_41765,N_41764);
xor U42063 (N_42063,N_41524,N_41689);
nand U42064 (N_42064,N_41659,N_41580);
or U42065 (N_42065,N_41938,N_41916);
and U42066 (N_42066,N_41614,N_41943);
nor U42067 (N_42067,N_41927,N_41757);
and U42068 (N_42068,N_41710,N_41740);
xnor U42069 (N_42069,N_41588,N_41915);
nor U42070 (N_42070,N_41816,N_41782);
nor U42071 (N_42071,N_41779,N_41711);
nor U42072 (N_42072,N_41666,N_41615);
nor U42073 (N_42073,N_41822,N_41800);
nor U42074 (N_42074,N_41925,N_41953);
and U42075 (N_42075,N_41585,N_41787);
and U42076 (N_42076,N_41629,N_41681);
nor U42077 (N_42077,N_41921,N_41712);
or U42078 (N_42078,N_41882,N_41825);
and U42079 (N_42079,N_41809,N_41797);
and U42080 (N_42080,N_41786,N_41986);
nor U42081 (N_42081,N_41683,N_41864);
xnor U42082 (N_42082,N_41571,N_41900);
nand U42083 (N_42083,N_41719,N_41724);
and U42084 (N_42084,N_41549,N_41885);
nand U42085 (N_42085,N_41961,N_41733);
nor U42086 (N_42086,N_41695,N_41903);
xor U42087 (N_42087,N_41977,N_41723);
nand U42088 (N_42088,N_41950,N_41993);
xnor U42089 (N_42089,N_41867,N_41542);
nand U42090 (N_42090,N_41967,N_41939);
or U42091 (N_42091,N_41508,N_41703);
or U42092 (N_42092,N_41619,N_41890);
and U42093 (N_42093,N_41798,N_41901);
xnor U42094 (N_42094,N_41562,N_41976);
or U42095 (N_42095,N_41662,N_41843);
nor U42096 (N_42096,N_41781,N_41587);
or U42097 (N_42097,N_41727,N_41637);
nand U42098 (N_42098,N_41565,N_41688);
or U42099 (N_42099,N_41652,N_41592);
or U42100 (N_42100,N_41875,N_41741);
xnor U42101 (N_42101,N_41928,N_41611);
nand U42102 (N_42102,N_41932,N_41503);
xnor U42103 (N_42103,N_41791,N_41532);
and U42104 (N_42104,N_41775,N_41617);
xor U42105 (N_42105,N_41590,N_41578);
xnor U42106 (N_42106,N_41960,N_41686);
or U42107 (N_42107,N_41841,N_41668);
xor U42108 (N_42108,N_41963,N_41858);
nor U42109 (N_42109,N_41623,N_41713);
nor U42110 (N_42110,N_41989,N_41706);
nor U42111 (N_42111,N_41601,N_41540);
nand U42112 (N_42112,N_41935,N_41958);
xnor U42113 (N_42113,N_41630,N_41653);
nor U42114 (N_42114,N_41987,N_41512);
and U42115 (N_42115,N_41535,N_41949);
nand U42116 (N_42116,N_41690,N_41720);
or U42117 (N_42117,N_41815,N_41920);
nand U42118 (N_42118,N_41811,N_41904);
xnor U42119 (N_42119,N_41705,N_41866);
nand U42120 (N_42120,N_41525,N_41817);
xor U42121 (N_42121,N_41831,N_41586);
or U42122 (N_42122,N_41626,N_41819);
and U42123 (N_42123,N_41910,N_41651);
nor U42124 (N_42124,N_41803,N_41734);
or U42125 (N_42125,N_41654,N_41517);
xnor U42126 (N_42126,N_41844,N_41852);
nand U42127 (N_42127,N_41533,N_41650);
nand U42128 (N_42128,N_41804,N_41763);
and U42129 (N_42129,N_41687,N_41768);
or U42130 (N_42130,N_41559,N_41944);
nor U42131 (N_42131,N_41769,N_41906);
or U42132 (N_42132,N_41554,N_41715);
nand U42133 (N_42133,N_41523,N_41507);
nand U42134 (N_42134,N_41628,N_41607);
xor U42135 (N_42135,N_41828,N_41564);
or U42136 (N_42136,N_41892,N_41528);
xnor U42137 (N_42137,N_41709,N_41876);
and U42138 (N_42138,N_41731,N_41671);
or U42139 (N_42139,N_41862,N_41998);
nand U42140 (N_42140,N_41842,N_41539);
or U42141 (N_42141,N_41930,N_41948);
or U42142 (N_42142,N_41839,N_41881);
nand U42143 (N_42143,N_41665,N_41606);
xor U42144 (N_42144,N_41534,N_41631);
nand U42145 (N_42145,N_41985,N_41812);
xnor U42146 (N_42146,N_41980,N_41962);
and U42147 (N_42147,N_41891,N_41936);
and U42148 (N_42148,N_41975,N_41893);
nand U42149 (N_42149,N_41946,N_41931);
xnor U42150 (N_42150,N_41555,N_41501);
and U42151 (N_42151,N_41633,N_41793);
nand U42152 (N_42152,N_41531,N_41698);
and U42153 (N_42153,N_41749,N_41513);
or U42154 (N_42154,N_41955,N_41941);
nor U42155 (N_42155,N_41558,N_41691);
nand U42156 (N_42156,N_41742,N_41641);
nand U42157 (N_42157,N_41767,N_41942);
nand U42158 (N_42158,N_41643,N_41569);
and U42159 (N_42159,N_41999,N_41640);
and U42160 (N_42160,N_41577,N_41954);
nand U42161 (N_42161,N_41773,N_41635);
or U42162 (N_42162,N_41506,N_41584);
nand U42163 (N_42163,N_41545,N_41634);
or U42164 (N_42164,N_41829,N_41693);
or U42165 (N_42165,N_41810,N_41835);
nor U42166 (N_42166,N_41735,N_41658);
xnor U42167 (N_42167,N_41660,N_41675);
xor U42168 (N_42168,N_41721,N_41756);
xnor U42169 (N_42169,N_41661,N_41648);
nor U42170 (N_42170,N_41622,N_41872);
or U42171 (N_42171,N_41981,N_41616);
or U42172 (N_42172,N_41808,N_41996);
nand U42173 (N_42173,N_41856,N_41556);
xnor U42174 (N_42174,N_41972,N_41568);
and U42175 (N_42175,N_41824,N_41991);
nand U42176 (N_42176,N_41956,N_41959);
or U42177 (N_42177,N_41951,N_41905);
nand U42178 (N_42178,N_41526,N_41701);
or U42179 (N_42179,N_41621,N_41853);
or U42180 (N_42180,N_41777,N_41870);
nor U42181 (N_42181,N_41833,N_41538);
or U42182 (N_42182,N_41674,N_41848);
nand U42183 (N_42183,N_41664,N_41888);
nand U42184 (N_42184,N_41682,N_41573);
nand U42185 (N_42185,N_41997,N_41837);
or U42186 (N_42186,N_41669,N_41596);
or U42187 (N_42187,N_41567,N_41969);
xnor U42188 (N_42188,N_41913,N_41663);
nor U42189 (N_42189,N_41699,N_41744);
or U42190 (N_42190,N_41550,N_41537);
xnor U42191 (N_42191,N_41970,N_41871);
or U42192 (N_42192,N_41620,N_41672);
nand U42193 (N_42193,N_41500,N_41850);
nand U42194 (N_42194,N_41521,N_41855);
nor U42195 (N_42195,N_41863,N_41908);
nor U42196 (N_42196,N_41912,N_41692);
or U42197 (N_42197,N_41947,N_41510);
xnor U42198 (N_42198,N_41717,N_41776);
xor U42199 (N_42199,N_41529,N_41514);
nand U42200 (N_42200,N_41748,N_41783);
or U42201 (N_42201,N_41544,N_41603);
or U42202 (N_42202,N_41902,N_41707);
or U42203 (N_42203,N_41879,N_41849);
and U42204 (N_42204,N_41730,N_41655);
or U42205 (N_42205,N_41696,N_41899);
and U42206 (N_42206,N_41575,N_41964);
nor U42207 (N_42207,N_41836,N_41718);
and U42208 (N_42208,N_41557,N_41530);
nand U42209 (N_42209,N_41736,N_41676);
nand U42210 (N_42210,N_41794,N_41760);
nor U42211 (N_42211,N_41560,N_41726);
nand U42212 (N_42212,N_41774,N_41854);
nand U42213 (N_42213,N_41605,N_41589);
nor U42214 (N_42214,N_41806,N_41553);
nand U42215 (N_42215,N_41680,N_41792);
xor U42216 (N_42216,N_41566,N_41515);
and U42217 (N_42217,N_41982,N_41801);
and U42218 (N_42218,N_41957,N_41543);
nand U42219 (N_42219,N_41750,N_41518);
and U42220 (N_42220,N_41884,N_41745);
nand U42221 (N_42221,N_41922,N_41802);
and U42222 (N_42222,N_41747,N_41911);
or U42223 (N_42223,N_41625,N_41739);
xnor U42224 (N_42224,N_41759,N_41994);
nor U42225 (N_42225,N_41896,N_41753);
and U42226 (N_42226,N_41886,N_41656);
nand U42227 (N_42227,N_41826,N_41624);
nand U42228 (N_42228,N_41846,N_41572);
nor U42229 (N_42229,N_41697,N_41561);
or U42230 (N_42230,N_41771,N_41762);
xor U42231 (N_42231,N_41919,N_41644);
nor U42232 (N_42232,N_41965,N_41677);
or U42233 (N_42233,N_41627,N_41971);
nor U42234 (N_42234,N_41602,N_41832);
xor U42235 (N_42235,N_41541,N_41583);
and U42236 (N_42236,N_41758,N_41563);
nor U42237 (N_42237,N_41859,N_41834);
xnor U42238 (N_42238,N_41708,N_41591);
and U42239 (N_42239,N_41516,N_41907);
nor U42240 (N_42240,N_41684,N_41778);
nor U42241 (N_42241,N_41636,N_41897);
xor U42242 (N_42242,N_41609,N_41548);
nor U42243 (N_42243,N_41511,N_41608);
nand U42244 (N_42244,N_41729,N_41704);
xnor U42245 (N_42245,N_41595,N_41847);
nand U42246 (N_42246,N_41795,N_41878);
or U42247 (N_42247,N_41647,N_41917);
or U42248 (N_42248,N_41722,N_41600);
or U42249 (N_42249,N_41754,N_41752);
nand U42250 (N_42250,N_41583,N_41762);
or U42251 (N_42251,N_41568,N_41917);
and U42252 (N_42252,N_41972,N_41726);
nand U42253 (N_42253,N_41884,N_41910);
nand U42254 (N_42254,N_41584,N_41965);
xnor U42255 (N_42255,N_41937,N_41863);
or U42256 (N_42256,N_41803,N_41917);
and U42257 (N_42257,N_41612,N_41952);
and U42258 (N_42258,N_41830,N_41728);
or U42259 (N_42259,N_41960,N_41534);
or U42260 (N_42260,N_41920,N_41845);
nor U42261 (N_42261,N_41979,N_41972);
or U42262 (N_42262,N_41991,N_41709);
and U42263 (N_42263,N_41647,N_41530);
or U42264 (N_42264,N_41680,N_41945);
or U42265 (N_42265,N_41928,N_41724);
and U42266 (N_42266,N_41715,N_41613);
nand U42267 (N_42267,N_41938,N_41873);
and U42268 (N_42268,N_41748,N_41913);
or U42269 (N_42269,N_41788,N_41944);
nand U42270 (N_42270,N_41510,N_41878);
and U42271 (N_42271,N_41887,N_41906);
or U42272 (N_42272,N_41744,N_41715);
and U42273 (N_42273,N_41904,N_41926);
or U42274 (N_42274,N_41706,N_41860);
nor U42275 (N_42275,N_41940,N_41718);
or U42276 (N_42276,N_41597,N_41791);
xor U42277 (N_42277,N_41821,N_41880);
nor U42278 (N_42278,N_41765,N_41811);
nor U42279 (N_42279,N_41944,N_41896);
xor U42280 (N_42280,N_41916,N_41715);
and U42281 (N_42281,N_41908,N_41616);
or U42282 (N_42282,N_41804,N_41959);
nor U42283 (N_42283,N_41976,N_41791);
xor U42284 (N_42284,N_41695,N_41724);
nor U42285 (N_42285,N_41975,N_41950);
nand U42286 (N_42286,N_41992,N_41507);
nor U42287 (N_42287,N_41699,N_41718);
and U42288 (N_42288,N_41792,N_41575);
xor U42289 (N_42289,N_41687,N_41724);
nand U42290 (N_42290,N_41641,N_41870);
nor U42291 (N_42291,N_41993,N_41519);
xnor U42292 (N_42292,N_41984,N_41911);
and U42293 (N_42293,N_41997,N_41500);
xnor U42294 (N_42294,N_41562,N_41630);
nor U42295 (N_42295,N_41666,N_41860);
and U42296 (N_42296,N_41934,N_41663);
nor U42297 (N_42297,N_41759,N_41767);
or U42298 (N_42298,N_41568,N_41975);
xnor U42299 (N_42299,N_41998,N_41760);
xor U42300 (N_42300,N_41665,N_41939);
nand U42301 (N_42301,N_41726,N_41545);
nand U42302 (N_42302,N_41754,N_41771);
xor U42303 (N_42303,N_41520,N_41738);
or U42304 (N_42304,N_41874,N_41639);
nand U42305 (N_42305,N_41776,N_41644);
xnor U42306 (N_42306,N_41710,N_41928);
xor U42307 (N_42307,N_41909,N_41948);
xnor U42308 (N_42308,N_41936,N_41999);
nor U42309 (N_42309,N_41620,N_41890);
nor U42310 (N_42310,N_41509,N_41844);
and U42311 (N_42311,N_41726,N_41762);
and U42312 (N_42312,N_41736,N_41646);
and U42313 (N_42313,N_41582,N_41636);
nand U42314 (N_42314,N_41708,N_41602);
and U42315 (N_42315,N_41641,N_41556);
and U42316 (N_42316,N_41909,N_41530);
xor U42317 (N_42317,N_41920,N_41773);
or U42318 (N_42318,N_41972,N_41954);
and U42319 (N_42319,N_41716,N_41924);
xor U42320 (N_42320,N_41905,N_41800);
nor U42321 (N_42321,N_41738,N_41809);
xnor U42322 (N_42322,N_41881,N_41810);
nor U42323 (N_42323,N_41976,N_41898);
xnor U42324 (N_42324,N_41992,N_41983);
nand U42325 (N_42325,N_41761,N_41797);
nand U42326 (N_42326,N_41601,N_41510);
xor U42327 (N_42327,N_41558,N_41554);
and U42328 (N_42328,N_41778,N_41591);
and U42329 (N_42329,N_41682,N_41762);
or U42330 (N_42330,N_41828,N_41596);
xor U42331 (N_42331,N_41637,N_41575);
xor U42332 (N_42332,N_41789,N_41666);
nor U42333 (N_42333,N_41539,N_41646);
xnor U42334 (N_42334,N_41733,N_41652);
nor U42335 (N_42335,N_41887,N_41822);
and U42336 (N_42336,N_41840,N_41708);
or U42337 (N_42337,N_41688,N_41785);
nor U42338 (N_42338,N_41866,N_41762);
xor U42339 (N_42339,N_41522,N_41776);
and U42340 (N_42340,N_41700,N_41677);
xor U42341 (N_42341,N_41713,N_41983);
and U42342 (N_42342,N_41509,N_41823);
nand U42343 (N_42343,N_41782,N_41500);
xnor U42344 (N_42344,N_41539,N_41550);
or U42345 (N_42345,N_41527,N_41855);
or U42346 (N_42346,N_41543,N_41548);
or U42347 (N_42347,N_41510,N_41867);
nand U42348 (N_42348,N_41577,N_41879);
xnor U42349 (N_42349,N_41611,N_41592);
nand U42350 (N_42350,N_41564,N_41657);
and U42351 (N_42351,N_41723,N_41914);
nor U42352 (N_42352,N_41632,N_41643);
or U42353 (N_42353,N_41680,N_41655);
nor U42354 (N_42354,N_41715,N_41837);
or U42355 (N_42355,N_41882,N_41717);
or U42356 (N_42356,N_41700,N_41587);
nand U42357 (N_42357,N_41556,N_41793);
and U42358 (N_42358,N_41557,N_41856);
nor U42359 (N_42359,N_41629,N_41714);
xnor U42360 (N_42360,N_41615,N_41636);
xor U42361 (N_42361,N_41825,N_41527);
nor U42362 (N_42362,N_41663,N_41639);
nor U42363 (N_42363,N_41613,N_41787);
and U42364 (N_42364,N_41899,N_41945);
nand U42365 (N_42365,N_41764,N_41844);
or U42366 (N_42366,N_41908,N_41776);
xnor U42367 (N_42367,N_41759,N_41966);
nand U42368 (N_42368,N_41744,N_41785);
nor U42369 (N_42369,N_41797,N_41619);
and U42370 (N_42370,N_41898,N_41815);
and U42371 (N_42371,N_41776,N_41681);
and U42372 (N_42372,N_41677,N_41865);
nor U42373 (N_42373,N_41510,N_41731);
nand U42374 (N_42374,N_41688,N_41502);
and U42375 (N_42375,N_41554,N_41533);
or U42376 (N_42376,N_41935,N_41821);
xnor U42377 (N_42377,N_41835,N_41886);
xor U42378 (N_42378,N_41819,N_41953);
or U42379 (N_42379,N_41624,N_41581);
nand U42380 (N_42380,N_41695,N_41514);
nand U42381 (N_42381,N_41982,N_41808);
nand U42382 (N_42382,N_41525,N_41985);
nor U42383 (N_42383,N_41595,N_41533);
and U42384 (N_42384,N_41967,N_41946);
and U42385 (N_42385,N_41988,N_41561);
or U42386 (N_42386,N_41600,N_41823);
xor U42387 (N_42387,N_41563,N_41879);
or U42388 (N_42388,N_41793,N_41908);
nor U42389 (N_42389,N_41722,N_41763);
or U42390 (N_42390,N_41729,N_41890);
and U42391 (N_42391,N_41583,N_41883);
and U42392 (N_42392,N_41844,N_41935);
xnor U42393 (N_42393,N_41568,N_41591);
nor U42394 (N_42394,N_41931,N_41978);
nand U42395 (N_42395,N_41614,N_41539);
nand U42396 (N_42396,N_41599,N_41809);
xnor U42397 (N_42397,N_41781,N_41880);
nand U42398 (N_42398,N_41785,N_41984);
nor U42399 (N_42399,N_41822,N_41819);
nand U42400 (N_42400,N_41508,N_41962);
xor U42401 (N_42401,N_41629,N_41531);
and U42402 (N_42402,N_41806,N_41937);
xnor U42403 (N_42403,N_41837,N_41964);
and U42404 (N_42404,N_41842,N_41896);
xor U42405 (N_42405,N_41927,N_41935);
nand U42406 (N_42406,N_41712,N_41527);
nor U42407 (N_42407,N_41546,N_41720);
and U42408 (N_42408,N_41935,N_41803);
xor U42409 (N_42409,N_41881,N_41863);
or U42410 (N_42410,N_41931,N_41554);
xnor U42411 (N_42411,N_41811,N_41599);
nand U42412 (N_42412,N_41753,N_41685);
or U42413 (N_42413,N_41858,N_41992);
and U42414 (N_42414,N_41973,N_41504);
and U42415 (N_42415,N_41708,N_41874);
and U42416 (N_42416,N_41861,N_41554);
nor U42417 (N_42417,N_41590,N_41994);
and U42418 (N_42418,N_41819,N_41898);
xnor U42419 (N_42419,N_41679,N_41673);
and U42420 (N_42420,N_41533,N_41837);
xor U42421 (N_42421,N_41946,N_41795);
and U42422 (N_42422,N_41811,N_41659);
and U42423 (N_42423,N_41983,N_41720);
or U42424 (N_42424,N_41718,N_41819);
nor U42425 (N_42425,N_41583,N_41993);
nand U42426 (N_42426,N_41816,N_41913);
nor U42427 (N_42427,N_41750,N_41752);
or U42428 (N_42428,N_41769,N_41911);
and U42429 (N_42429,N_41662,N_41710);
xnor U42430 (N_42430,N_41868,N_41531);
or U42431 (N_42431,N_41667,N_41787);
xor U42432 (N_42432,N_41698,N_41819);
nand U42433 (N_42433,N_41532,N_41523);
nor U42434 (N_42434,N_41639,N_41918);
and U42435 (N_42435,N_41817,N_41848);
or U42436 (N_42436,N_41623,N_41731);
nand U42437 (N_42437,N_41650,N_41945);
or U42438 (N_42438,N_41527,N_41736);
and U42439 (N_42439,N_41558,N_41580);
nand U42440 (N_42440,N_41671,N_41785);
nor U42441 (N_42441,N_41580,N_41823);
nand U42442 (N_42442,N_41791,N_41613);
nor U42443 (N_42443,N_41613,N_41735);
or U42444 (N_42444,N_41783,N_41892);
and U42445 (N_42445,N_41764,N_41536);
and U42446 (N_42446,N_41834,N_41752);
nor U42447 (N_42447,N_41541,N_41897);
nor U42448 (N_42448,N_41986,N_41811);
and U42449 (N_42449,N_41947,N_41910);
nor U42450 (N_42450,N_41761,N_41882);
xnor U42451 (N_42451,N_41985,N_41688);
nand U42452 (N_42452,N_41544,N_41501);
and U42453 (N_42453,N_41796,N_41556);
and U42454 (N_42454,N_41685,N_41739);
or U42455 (N_42455,N_41868,N_41708);
nand U42456 (N_42456,N_41512,N_41695);
nor U42457 (N_42457,N_41757,N_41959);
and U42458 (N_42458,N_41941,N_41631);
xnor U42459 (N_42459,N_41871,N_41695);
nor U42460 (N_42460,N_41976,N_41714);
nor U42461 (N_42461,N_41556,N_41766);
nand U42462 (N_42462,N_41707,N_41596);
or U42463 (N_42463,N_41812,N_41789);
and U42464 (N_42464,N_41826,N_41553);
or U42465 (N_42465,N_41596,N_41558);
nor U42466 (N_42466,N_41988,N_41636);
nor U42467 (N_42467,N_41739,N_41936);
nor U42468 (N_42468,N_41739,N_41814);
and U42469 (N_42469,N_41896,N_41612);
or U42470 (N_42470,N_41886,N_41942);
or U42471 (N_42471,N_41887,N_41842);
or U42472 (N_42472,N_41690,N_41646);
and U42473 (N_42473,N_41764,N_41613);
xor U42474 (N_42474,N_41675,N_41688);
and U42475 (N_42475,N_41582,N_41895);
and U42476 (N_42476,N_41598,N_41700);
nand U42477 (N_42477,N_41654,N_41796);
and U42478 (N_42478,N_41916,N_41825);
and U42479 (N_42479,N_41832,N_41979);
nor U42480 (N_42480,N_41977,N_41901);
xor U42481 (N_42481,N_41829,N_41830);
xnor U42482 (N_42482,N_41676,N_41623);
and U42483 (N_42483,N_41723,N_41649);
xnor U42484 (N_42484,N_41683,N_41877);
nand U42485 (N_42485,N_41896,N_41845);
xor U42486 (N_42486,N_41582,N_41782);
nand U42487 (N_42487,N_41762,N_41686);
nor U42488 (N_42488,N_41569,N_41656);
or U42489 (N_42489,N_41945,N_41526);
nand U42490 (N_42490,N_41604,N_41629);
nand U42491 (N_42491,N_41641,N_41885);
nor U42492 (N_42492,N_41558,N_41683);
nand U42493 (N_42493,N_41874,N_41779);
nand U42494 (N_42494,N_41745,N_41825);
and U42495 (N_42495,N_41535,N_41582);
and U42496 (N_42496,N_41978,N_41865);
and U42497 (N_42497,N_41657,N_41999);
nand U42498 (N_42498,N_41651,N_41675);
nand U42499 (N_42499,N_41938,N_41930);
and U42500 (N_42500,N_42273,N_42227);
or U42501 (N_42501,N_42162,N_42037);
nor U42502 (N_42502,N_42336,N_42422);
nor U42503 (N_42503,N_42113,N_42197);
or U42504 (N_42504,N_42428,N_42215);
nand U42505 (N_42505,N_42109,N_42119);
nor U42506 (N_42506,N_42298,N_42414);
nand U42507 (N_42507,N_42387,N_42258);
nor U42508 (N_42508,N_42405,N_42398);
nand U42509 (N_42509,N_42150,N_42321);
nor U42510 (N_42510,N_42304,N_42168);
or U42511 (N_42511,N_42324,N_42021);
or U42512 (N_42512,N_42261,N_42346);
or U42513 (N_42513,N_42341,N_42266);
and U42514 (N_42514,N_42093,N_42272);
and U42515 (N_42515,N_42016,N_42138);
or U42516 (N_42516,N_42161,N_42471);
xnor U42517 (N_42517,N_42046,N_42112);
or U42518 (N_42518,N_42107,N_42061);
xor U42519 (N_42519,N_42404,N_42050);
xnor U42520 (N_42520,N_42207,N_42169);
and U42521 (N_42521,N_42262,N_42089);
xnor U42522 (N_42522,N_42314,N_42320);
nor U42523 (N_42523,N_42310,N_42449);
xor U42524 (N_42524,N_42147,N_42388);
nor U42525 (N_42525,N_42146,N_42313);
nor U42526 (N_42526,N_42250,N_42182);
nand U42527 (N_42527,N_42458,N_42069);
and U42528 (N_42528,N_42438,N_42493);
nand U42529 (N_42529,N_42189,N_42277);
nand U42530 (N_42530,N_42305,N_42049);
xnor U42531 (N_42531,N_42319,N_42437);
nand U42532 (N_42532,N_42027,N_42203);
or U42533 (N_42533,N_42470,N_42008);
and U42534 (N_42534,N_42199,N_42009);
nor U42535 (N_42535,N_42245,N_42148);
xnor U42536 (N_42536,N_42483,N_42095);
or U42537 (N_42537,N_42312,N_42073);
xnor U42538 (N_42538,N_42303,N_42022);
xor U42539 (N_42539,N_42209,N_42097);
nor U42540 (N_42540,N_42126,N_42395);
xnor U42541 (N_42541,N_42407,N_42263);
xor U42542 (N_42542,N_42375,N_42447);
nand U42543 (N_42543,N_42391,N_42122);
nand U42544 (N_42544,N_42415,N_42159);
nand U42545 (N_42545,N_42251,N_42482);
and U42546 (N_42546,N_42006,N_42397);
xnor U42547 (N_42547,N_42334,N_42323);
and U42548 (N_42548,N_42165,N_42475);
nand U42549 (N_42549,N_42408,N_42418);
nor U42550 (N_42550,N_42038,N_42004);
nand U42551 (N_42551,N_42284,N_42176);
and U42552 (N_42552,N_42390,N_42079);
nand U42553 (N_42553,N_42456,N_42130);
nor U42554 (N_42554,N_42005,N_42469);
and U42555 (N_42555,N_42379,N_42349);
and U42556 (N_42556,N_42236,N_42246);
or U42557 (N_42557,N_42143,N_42208);
nand U42558 (N_42558,N_42317,N_42108);
nor U42559 (N_42559,N_42115,N_42059);
xnor U42560 (N_42560,N_42386,N_42232);
or U42561 (N_42561,N_42043,N_42399);
nor U42562 (N_42562,N_42274,N_42139);
or U42563 (N_42563,N_42023,N_42025);
xor U42564 (N_42564,N_42366,N_42413);
and U42565 (N_42565,N_42171,N_42100);
nor U42566 (N_42566,N_42243,N_42495);
or U42567 (N_42567,N_42219,N_42497);
nor U42568 (N_42568,N_42459,N_42098);
or U42569 (N_42569,N_42256,N_42344);
xor U42570 (N_42570,N_42086,N_42400);
and U42571 (N_42571,N_42218,N_42087);
nor U42572 (N_42572,N_42491,N_42091);
xnor U42573 (N_42573,N_42178,N_42442);
and U42574 (N_42574,N_42354,N_42014);
and U42575 (N_42575,N_42393,N_42105);
nand U42576 (N_42576,N_42235,N_42396);
xor U42577 (N_42577,N_42142,N_42081);
xor U42578 (N_42578,N_42292,N_42015);
xor U42579 (N_42579,N_42440,N_42071);
nor U42580 (N_42580,N_42350,N_42177);
and U42581 (N_42581,N_42315,N_42196);
nand U42582 (N_42582,N_42231,N_42496);
and U42583 (N_42583,N_42034,N_42260);
xor U42584 (N_42584,N_42096,N_42289);
or U42585 (N_42585,N_42134,N_42441);
xnor U42586 (N_42586,N_42020,N_42193);
nor U42587 (N_42587,N_42200,N_42247);
xor U42588 (N_42588,N_42052,N_42402);
xnor U42589 (N_42589,N_42233,N_42474);
nor U42590 (N_42590,N_42392,N_42488);
nand U42591 (N_42591,N_42352,N_42360);
xor U42592 (N_42592,N_42286,N_42181);
and U42593 (N_42593,N_42160,N_42299);
or U42594 (N_42594,N_42135,N_42282);
nand U42595 (N_42595,N_42378,N_42296);
xor U42596 (N_42596,N_42187,N_42367);
nand U42597 (N_42597,N_42270,N_42033);
xor U42598 (N_42598,N_42088,N_42190);
nor U42599 (N_42599,N_42464,N_42267);
and U42600 (N_42600,N_42028,N_42067);
or U42601 (N_42601,N_42424,N_42291);
nand U42602 (N_42602,N_42467,N_42104);
xor U42603 (N_42603,N_42127,N_42311);
nor U42604 (N_42604,N_42452,N_42080);
xnor U42605 (N_42605,N_42363,N_42412);
xnor U42606 (N_42606,N_42044,N_42094);
and U42607 (N_42607,N_42255,N_42013);
nor U42608 (N_42608,N_42372,N_42191);
and U42609 (N_42609,N_42487,N_42380);
nor U42610 (N_42610,N_42185,N_42241);
xnor U42611 (N_42611,N_42252,N_42430);
nand U42612 (N_42612,N_42417,N_42448);
nor U42613 (N_42613,N_42056,N_42129);
and U42614 (N_42614,N_42318,N_42478);
nand U42615 (N_42615,N_42221,N_42362);
xor U42616 (N_42616,N_42342,N_42382);
and U42617 (N_42617,N_42431,N_42206);
nor U42618 (N_42618,N_42410,N_42217);
nor U42619 (N_42619,N_42123,N_42268);
nor U42620 (N_42620,N_42198,N_42293);
xor U42621 (N_42621,N_42460,N_42133);
xor U42622 (N_42622,N_42288,N_42225);
or U42623 (N_42623,N_42085,N_42180);
xor U42624 (N_42624,N_42099,N_42216);
or U42625 (N_42625,N_42394,N_42083);
xnor U42626 (N_42626,N_42144,N_42204);
nor U42627 (N_42627,N_42423,N_42429);
nor U42628 (N_42628,N_42007,N_42163);
nor U42629 (N_42629,N_42019,N_42030);
nand U42630 (N_42630,N_42121,N_42285);
nand U42631 (N_42631,N_42457,N_42173);
xnor U42632 (N_42632,N_42017,N_42172);
nor U42633 (N_42633,N_42103,N_42347);
nand U42634 (N_42634,N_42276,N_42444);
nor U42635 (N_42635,N_42090,N_42371);
xnor U42636 (N_42636,N_42331,N_42157);
nand U42637 (N_42637,N_42051,N_42077);
and U42638 (N_42638,N_42114,N_42041);
nor U42639 (N_42639,N_42329,N_42443);
nand U42640 (N_42640,N_42461,N_42082);
and U42641 (N_42641,N_42434,N_42477);
nor U42642 (N_42642,N_42365,N_42158);
nand U42643 (N_42643,N_42222,N_42253);
or U42644 (N_42644,N_42128,N_42340);
nand U42645 (N_42645,N_42377,N_42136);
xnor U42646 (N_42646,N_42226,N_42368);
or U42647 (N_42647,N_42132,N_42381);
nand U42648 (N_42648,N_42409,N_42376);
xor U42649 (N_42649,N_42401,N_42295);
and U42650 (N_42650,N_42029,N_42358);
and U42651 (N_42651,N_42140,N_42453);
xor U42652 (N_42652,N_42472,N_42339);
nand U42653 (N_42653,N_42244,N_42152);
nand U42654 (N_42654,N_42271,N_42047);
nand U42655 (N_42655,N_42151,N_42445);
xnor U42656 (N_42656,N_42118,N_42306);
xnor U42657 (N_42657,N_42433,N_42308);
xor U42658 (N_42658,N_42058,N_42205);
and U42659 (N_42659,N_42063,N_42045);
nand U42660 (N_42660,N_42384,N_42489);
nor U42661 (N_42661,N_42283,N_42195);
xor U42662 (N_42662,N_42454,N_42072);
xnor U42663 (N_42663,N_42137,N_42359);
nor U42664 (N_42664,N_42290,N_42055);
nor U42665 (N_42665,N_42175,N_42463);
and U42666 (N_42666,N_42210,N_42435);
xor U42667 (N_42667,N_42436,N_42111);
nand U42668 (N_42668,N_42337,N_42057);
and U42669 (N_42669,N_42468,N_42242);
or U42670 (N_42670,N_42326,N_42498);
and U42671 (N_42671,N_42476,N_42214);
nand U42672 (N_42672,N_42068,N_42343);
or U42673 (N_42673,N_42026,N_42145);
and U42674 (N_42674,N_42066,N_42345);
xor U42675 (N_42675,N_42070,N_42425);
and U42676 (N_42676,N_42076,N_42333);
nor U42677 (N_42677,N_42439,N_42383);
and U42678 (N_42678,N_42092,N_42064);
xor U42679 (N_42679,N_42330,N_42328);
nand U42680 (N_42680,N_42054,N_42278);
nand U42681 (N_42681,N_42300,N_42212);
xnor U42682 (N_42682,N_42240,N_42325);
nor U42683 (N_42683,N_42265,N_42234);
or U42684 (N_42684,N_42010,N_42406);
and U42685 (N_42685,N_42238,N_42389);
and U42686 (N_42686,N_42364,N_42355);
and U42687 (N_42687,N_42174,N_42213);
nor U42688 (N_42688,N_42228,N_42031);
xor U42689 (N_42689,N_42124,N_42248);
nand U42690 (N_42690,N_42155,N_42116);
xor U42691 (N_42691,N_42322,N_42403);
xnor U42692 (N_42692,N_42229,N_42451);
xor U42693 (N_42693,N_42426,N_42184);
and U42694 (N_42694,N_42421,N_42110);
or U42695 (N_42695,N_42281,N_42164);
and U42696 (N_42696,N_42060,N_42192);
nor U42697 (N_42697,N_42040,N_42356);
and U42698 (N_42698,N_42032,N_42149);
nor U42699 (N_42699,N_42125,N_42369);
or U42700 (N_42700,N_42279,N_42194);
nand U42701 (N_42701,N_42301,N_42280);
xor U42702 (N_42702,N_42494,N_42042);
and U42703 (N_42703,N_42183,N_42332);
or U42704 (N_42704,N_42074,N_42370);
or U42705 (N_42705,N_42230,N_42499);
nand U42706 (N_42706,N_42078,N_42361);
or U42707 (N_42707,N_42201,N_42338);
or U42708 (N_42708,N_42327,N_42167);
and U42709 (N_42709,N_42154,N_42465);
nor U42710 (N_42710,N_42224,N_42257);
or U42711 (N_42711,N_42202,N_42486);
xor U42712 (N_42712,N_42259,N_42120);
xnor U42713 (N_42713,N_42170,N_42102);
nand U42714 (N_42714,N_42012,N_42188);
and U42715 (N_42715,N_42053,N_42481);
and U42716 (N_42716,N_42039,N_42294);
xnor U42717 (N_42717,N_42000,N_42353);
or U42718 (N_42718,N_42075,N_42351);
nor U42719 (N_42719,N_42141,N_42264);
nor U42720 (N_42720,N_42275,N_42335);
xor U42721 (N_42721,N_42237,N_42357);
nor U42722 (N_42722,N_42411,N_42419);
xnor U42723 (N_42723,N_42416,N_42001);
xnor U42724 (N_42724,N_42062,N_42309);
nor U42725 (N_42725,N_42287,N_42024);
nor U42726 (N_42726,N_42490,N_42427);
or U42727 (N_42727,N_42035,N_42269);
nand U42728 (N_42728,N_42153,N_42374);
or U42729 (N_42729,N_42084,N_42131);
nor U42730 (N_42730,N_42462,N_42156);
nor U42731 (N_42731,N_42011,N_42307);
nand U42732 (N_42732,N_42223,N_42065);
nor U42733 (N_42733,N_42249,N_42479);
or U42734 (N_42734,N_42466,N_42450);
nand U42735 (N_42735,N_42446,N_42220);
xor U42736 (N_42736,N_42117,N_42048);
nand U42737 (N_42737,N_42385,N_42003);
or U42738 (N_42738,N_42373,N_42179);
or U42739 (N_42739,N_42036,N_42239);
nor U42740 (N_42740,N_42316,N_42302);
and U42741 (N_42741,N_42432,N_42473);
or U42742 (N_42742,N_42492,N_42485);
nor U42743 (N_42743,N_42254,N_42348);
xnor U42744 (N_42744,N_42106,N_42018);
xor U42745 (N_42745,N_42002,N_42186);
and U42746 (N_42746,N_42166,N_42211);
xnor U42747 (N_42747,N_42484,N_42480);
nor U42748 (N_42748,N_42455,N_42297);
or U42749 (N_42749,N_42420,N_42101);
and U42750 (N_42750,N_42169,N_42368);
nand U42751 (N_42751,N_42262,N_42342);
xnor U42752 (N_42752,N_42323,N_42496);
nand U42753 (N_42753,N_42112,N_42324);
or U42754 (N_42754,N_42430,N_42388);
and U42755 (N_42755,N_42256,N_42198);
nor U42756 (N_42756,N_42011,N_42319);
nand U42757 (N_42757,N_42003,N_42118);
xor U42758 (N_42758,N_42457,N_42288);
nor U42759 (N_42759,N_42464,N_42044);
nand U42760 (N_42760,N_42319,N_42340);
or U42761 (N_42761,N_42188,N_42304);
and U42762 (N_42762,N_42116,N_42343);
or U42763 (N_42763,N_42167,N_42350);
and U42764 (N_42764,N_42371,N_42208);
xor U42765 (N_42765,N_42202,N_42183);
nor U42766 (N_42766,N_42240,N_42362);
and U42767 (N_42767,N_42226,N_42439);
nor U42768 (N_42768,N_42068,N_42147);
xnor U42769 (N_42769,N_42491,N_42205);
nor U42770 (N_42770,N_42080,N_42177);
nor U42771 (N_42771,N_42090,N_42238);
nand U42772 (N_42772,N_42371,N_42232);
nor U42773 (N_42773,N_42075,N_42456);
nor U42774 (N_42774,N_42172,N_42055);
or U42775 (N_42775,N_42199,N_42428);
and U42776 (N_42776,N_42345,N_42266);
or U42777 (N_42777,N_42002,N_42128);
nand U42778 (N_42778,N_42125,N_42042);
xor U42779 (N_42779,N_42441,N_42232);
nand U42780 (N_42780,N_42078,N_42039);
xnor U42781 (N_42781,N_42120,N_42169);
or U42782 (N_42782,N_42423,N_42023);
nor U42783 (N_42783,N_42040,N_42104);
nand U42784 (N_42784,N_42384,N_42102);
and U42785 (N_42785,N_42040,N_42033);
nor U42786 (N_42786,N_42167,N_42157);
and U42787 (N_42787,N_42033,N_42103);
and U42788 (N_42788,N_42063,N_42064);
or U42789 (N_42789,N_42099,N_42247);
nor U42790 (N_42790,N_42336,N_42143);
nand U42791 (N_42791,N_42449,N_42370);
nor U42792 (N_42792,N_42007,N_42299);
or U42793 (N_42793,N_42336,N_42433);
xor U42794 (N_42794,N_42443,N_42438);
nor U42795 (N_42795,N_42490,N_42208);
xor U42796 (N_42796,N_42314,N_42048);
nand U42797 (N_42797,N_42120,N_42181);
nand U42798 (N_42798,N_42392,N_42487);
xor U42799 (N_42799,N_42482,N_42389);
nand U42800 (N_42800,N_42469,N_42157);
nand U42801 (N_42801,N_42304,N_42108);
nand U42802 (N_42802,N_42020,N_42036);
nand U42803 (N_42803,N_42283,N_42088);
and U42804 (N_42804,N_42129,N_42391);
xnor U42805 (N_42805,N_42219,N_42088);
nor U42806 (N_42806,N_42140,N_42046);
nand U42807 (N_42807,N_42303,N_42188);
or U42808 (N_42808,N_42248,N_42020);
nor U42809 (N_42809,N_42273,N_42464);
nor U42810 (N_42810,N_42363,N_42494);
nand U42811 (N_42811,N_42443,N_42204);
or U42812 (N_42812,N_42014,N_42270);
nand U42813 (N_42813,N_42460,N_42408);
nor U42814 (N_42814,N_42494,N_42290);
xor U42815 (N_42815,N_42089,N_42308);
or U42816 (N_42816,N_42003,N_42005);
and U42817 (N_42817,N_42476,N_42071);
nor U42818 (N_42818,N_42469,N_42179);
nand U42819 (N_42819,N_42481,N_42200);
or U42820 (N_42820,N_42278,N_42437);
nor U42821 (N_42821,N_42216,N_42038);
and U42822 (N_42822,N_42485,N_42072);
or U42823 (N_42823,N_42093,N_42176);
nor U42824 (N_42824,N_42280,N_42383);
and U42825 (N_42825,N_42028,N_42190);
xor U42826 (N_42826,N_42449,N_42337);
or U42827 (N_42827,N_42419,N_42106);
nor U42828 (N_42828,N_42483,N_42409);
nand U42829 (N_42829,N_42343,N_42468);
nor U42830 (N_42830,N_42287,N_42318);
xnor U42831 (N_42831,N_42044,N_42018);
nand U42832 (N_42832,N_42373,N_42042);
or U42833 (N_42833,N_42013,N_42021);
or U42834 (N_42834,N_42374,N_42074);
nor U42835 (N_42835,N_42384,N_42097);
xor U42836 (N_42836,N_42252,N_42024);
or U42837 (N_42837,N_42437,N_42311);
nand U42838 (N_42838,N_42340,N_42135);
or U42839 (N_42839,N_42252,N_42224);
or U42840 (N_42840,N_42188,N_42142);
or U42841 (N_42841,N_42002,N_42172);
or U42842 (N_42842,N_42043,N_42334);
and U42843 (N_42843,N_42353,N_42162);
nor U42844 (N_42844,N_42128,N_42263);
nor U42845 (N_42845,N_42416,N_42089);
xor U42846 (N_42846,N_42159,N_42289);
or U42847 (N_42847,N_42431,N_42421);
and U42848 (N_42848,N_42284,N_42209);
or U42849 (N_42849,N_42006,N_42149);
or U42850 (N_42850,N_42414,N_42342);
or U42851 (N_42851,N_42206,N_42145);
xor U42852 (N_42852,N_42326,N_42353);
or U42853 (N_42853,N_42285,N_42493);
nand U42854 (N_42854,N_42203,N_42021);
or U42855 (N_42855,N_42451,N_42499);
xnor U42856 (N_42856,N_42400,N_42035);
nand U42857 (N_42857,N_42417,N_42457);
xor U42858 (N_42858,N_42104,N_42253);
xnor U42859 (N_42859,N_42364,N_42220);
nand U42860 (N_42860,N_42033,N_42422);
or U42861 (N_42861,N_42099,N_42173);
xor U42862 (N_42862,N_42449,N_42403);
and U42863 (N_42863,N_42159,N_42382);
xnor U42864 (N_42864,N_42341,N_42304);
nand U42865 (N_42865,N_42428,N_42342);
xnor U42866 (N_42866,N_42113,N_42404);
or U42867 (N_42867,N_42235,N_42429);
nand U42868 (N_42868,N_42279,N_42438);
or U42869 (N_42869,N_42016,N_42304);
and U42870 (N_42870,N_42301,N_42202);
xnor U42871 (N_42871,N_42074,N_42301);
nor U42872 (N_42872,N_42028,N_42025);
or U42873 (N_42873,N_42221,N_42384);
or U42874 (N_42874,N_42494,N_42283);
and U42875 (N_42875,N_42326,N_42106);
and U42876 (N_42876,N_42420,N_42451);
nand U42877 (N_42877,N_42421,N_42141);
nor U42878 (N_42878,N_42401,N_42025);
xor U42879 (N_42879,N_42228,N_42326);
nand U42880 (N_42880,N_42375,N_42187);
nand U42881 (N_42881,N_42413,N_42280);
or U42882 (N_42882,N_42219,N_42456);
nand U42883 (N_42883,N_42271,N_42496);
nor U42884 (N_42884,N_42361,N_42005);
nor U42885 (N_42885,N_42344,N_42243);
nand U42886 (N_42886,N_42319,N_42254);
nor U42887 (N_42887,N_42242,N_42344);
nor U42888 (N_42888,N_42428,N_42376);
and U42889 (N_42889,N_42212,N_42210);
xor U42890 (N_42890,N_42395,N_42030);
xnor U42891 (N_42891,N_42038,N_42397);
nand U42892 (N_42892,N_42080,N_42354);
nand U42893 (N_42893,N_42121,N_42415);
and U42894 (N_42894,N_42444,N_42074);
xnor U42895 (N_42895,N_42151,N_42369);
or U42896 (N_42896,N_42337,N_42293);
or U42897 (N_42897,N_42450,N_42003);
and U42898 (N_42898,N_42110,N_42277);
nand U42899 (N_42899,N_42218,N_42197);
xor U42900 (N_42900,N_42419,N_42308);
xnor U42901 (N_42901,N_42105,N_42494);
nor U42902 (N_42902,N_42060,N_42062);
nor U42903 (N_42903,N_42104,N_42109);
nor U42904 (N_42904,N_42112,N_42330);
nand U42905 (N_42905,N_42246,N_42151);
nand U42906 (N_42906,N_42087,N_42037);
nand U42907 (N_42907,N_42063,N_42231);
or U42908 (N_42908,N_42150,N_42335);
xor U42909 (N_42909,N_42082,N_42450);
or U42910 (N_42910,N_42326,N_42217);
nor U42911 (N_42911,N_42068,N_42271);
or U42912 (N_42912,N_42358,N_42474);
and U42913 (N_42913,N_42188,N_42368);
xor U42914 (N_42914,N_42395,N_42135);
nor U42915 (N_42915,N_42224,N_42290);
and U42916 (N_42916,N_42498,N_42106);
or U42917 (N_42917,N_42313,N_42252);
and U42918 (N_42918,N_42423,N_42411);
xnor U42919 (N_42919,N_42150,N_42124);
nor U42920 (N_42920,N_42292,N_42128);
and U42921 (N_42921,N_42284,N_42135);
and U42922 (N_42922,N_42258,N_42305);
and U42923 (N_42923,N_42117,N_42272);
nor U42924 (N_42924,N_42366,N_42323);
nand U42925 (N_42925,N_42127,N_42331);
nor U42926 (N_42926,N_42336,N_42156);
and U42927 (N_42927,N_42279,N_42391);
nand U42928 (N_42928,N_42464,N_42013);
xnor U42929 (N_42929,N_42275,N_42201);
and U42930 (N_42930,N_42141,N_42032);
and U42931 (N_42931,N_42014,N_42113);
or U42932 (N_42932,N_42287,N_42221);
xnor U42933 (N_42933,N_42107,N_42388);
nand U42934 (N_42934,N_42401,N_42019);
nand U42935 (N_42935,N_42098,N_42192);
or U42936 (N_42936,N_42146,N_42371);
and U42937 (N_42937,N_42238,N_42230);
or U42938 (N_42938,N_42059,N_42498);
xnor U42939 (N_42939,N_42165,N_42111);
xor U42940 (N_42940,N_42063,N_42232);
nor U42941 (N_42941,N_42427,N_42288);
or U42942 (N_42942,N_42071,N_42315);
and U42943 (N_42943,N_42164,N_42123);
xnor U42944 (N_42944,N_42319,N_42449);
nor U42945 (N_42945,N_42253,N_42496);
or U42946 (N_42946,N_42097,N_42193);
and U42947 (N_42947,N_42246,N_42076);
or U42948 (N_42948,N_42463,N_42489);
nand U42949 (N_42949,N_42216,N_42024);
nor U42950 (N_42950,N_42440,N_42465);
nand U42951 (N_42951,N_42499,N_42432);
xnor U42952 (N_42952,N_42499,N_42138);
nor U42953 (N_42953,N_42286,N_42287);
or U42954 (N_42954,N_42162,N_42115);
nor U42955 (N_42955,N_42365,N_42364);
and U42956 (N_42956,N_42451,N_42128);
nand U42957 (N_42957,N_42065,N_42362);
nand U42958 (N_42958,N_42245,N_42322);
and U42959 (N_42959,N_42332,N_42224);
nand U42960 (N_42960,N_42101,N_42182);
or U42961 (N_42961,N_42243,N_42474);
and U42962 (N_42962,N_42136,N_42457);
and U42963 (N_42963,N_42271,N_42127);
nand U42964 (N_42964,N_42017,N_42099);
nor U42965 (N_42965,N_42260,N_42054);
and U42966 (N_42966,N_42228,N_42493);
or U42967 (N_42967,N_42281,N_42254);
and U42968 (N_42968,N_42396,N_42297);
nand U42969 (N_42969,N_42257,N_42176);
nand U42970 (N_42970,N_42487,N_42284);
or U42971 (N_42971,N_42279,N_42368);
nor U42972 (N_42972,N_42134,N_42477);
or U42973 (N_42973,N_42383,N_42031);
or U42974 (N_42974,N_42280,N_42487);
and U42975 (N_42975,N_42158,N_42326);
or U42976 (N_42976,N_42040,N_42463);
xor U42977 (N_42977,N_42452,N_42225);
nor U42978 (N_42978,N_42331,N_42325);
and U42979 (N_42979,N_42379,N_42184);
nand U42980 (N_42980,N_42237,N_42263);
and U42981 (N_42981,N_42161,N_42383);
xnor U42982 (N_42982,N_42491,N_42366);
nor U42983 (N_42983,N_42428,N_42203);
xor U42984 (N_42984,N_42353,N_42498);
and U42985 (N_42985,N_42197,N_42426);
xor U42986 (N_42986,N_42047,N_42329);
and U42987 (N_42987,N_42186,N_42423);
xor U42988 (N_42988,N_42217,N_42485);
nand U42989 (N_42989,N_42061,N_42366);
and U42990 (N_42990,N_42263,N_42138);
nor U42991 (N_42991,N_42371,N_42408);
nand U42992 (N_42992,N_42313,N_42224);
nand U42993 (N_42993,N_42357,N_42452);
or U42994 (N_42994,N_42076,N_42012);
or U42995 (N_42995,N_42240,N_42262);
or U42996 (N_42996,N_42037,N_42459);
and U42997 (N_42997,N_42217,N_42053);
nand U42998 (N_42998,N_42222,N_42389);
nor U42999 (N_42999,N_42271,N_42202);
or U43000 (N_43000,N_42968,N_42662);
and U43001 (N_43001,N_42514,N_42617);
xor U43002 (N_43002,N_42725,N_42945);
nand U43003 (N_43003,N_42831,N_42929);
and U43004 (N_43004,N_42598,N_42814);
or U43005 (N_43005,N_42600,N_42592);
nand U43006 (N_43006,N_42848,N_42665);
and U43007 (N_43007,N_42791,N_42888);
xor U43008 (N_43008,N_42918,N_42944);
nand U43009 (N_43009,N_42841,N_42533);
nand U43010 (N_43010,N_42647,N_42842);
or U43011 (N_43011,N_42840,N_42671);
and U43012 (N_43012,N_42556,N_42534);
nand U43013 (N_43013,N_42790,N_42737);
nand U43014 (N_43014,N_42891,N_42905);
nand U43015 (N_43015,N_42864,N_42988);
or U43016 (N_43016,N_42626,N_42717);
nand U43017 (N_43017,N_42588,N_42693);
xnor U43018 (N_43018,N_42974,N_42750);
and U43019 (N_43019,N_42937,N_42976);
nand U43020 (N_43020,N_42505,N_42604);
xnor U43021 (N_43021,N_42874,N_42913);
nor U43022 (N_43022,N_42501,N_42923);
nand U43023 (N_43023,N_42813,N_42981);
or U43024 (N_43024,N_42773,N_42922);
xnor U43025 (N_43025,N_42759,N_42729);
or U43026 (N_43026,N_42704,N_42557);
xor U43027 (N_43027,N_42771,N_42743);
and U43028 (N_43028,N_42719,N_42889);
nor U43029 (N_43029,N_42690,N_42881);
or U43030 (N_43030,N_42825,N_42712);
nor U43031 (N_43031,N_42837,N_42979);
nor U43032 (N_43032,N_42832,N_42894);
xnor U43033 (N_43033,N_42769,N_42628);
and U43034 (N_43034,N_42518,N_42836);
or U43035 (N_43035,N_42839,N_42637);
nor U43036 (N_43036,N_42555,N_42686);
nor U43037 (N_43037,N_42632,N_42609);
nor U43038 (N_43038,N_42576,N_42614);
or U43039 (N_43039,N_42795,N_42920);
nand U43040 (N_43040,N_42833,N_42957);
or U43041 (N_43041,N_42644,N_42776);
nor U43042 (N_43042,N_42823,N_42596);
xor U43043 (N_43043,N_42511,N_42990);
or U43044 (N_43044,N_42789,N_42910);
nand U43045 (N_43045,N_42544,N_42897);
nand U43046 (N_43046,N_42765,N_42901);
or U43047 (N_43047,N_42784,N_42932);
or U43048 (N_43048,N_42657,N_42992);
and U43049 (N_43049,N_42969,N_42744);
or U43050 (N_43050,N_42740,N_42512);
xnor U43051 (N_43051,N_42540,N_42618);
xnor U43052 (N_43052,N_42579,N_42653);
xnor U43053 (N_43053,N_42735,N_42568);
nand U43054 (N_43054,N_42782,N_42705);
xnor U43055 (N_43055,N_42654,N_42925);
and U43056 (N_43056,N_42786,N_42589);
nor U43057 (N_43057,N_42955,N_42800);
nand U43058 (N_43058,N_42687,N_42503);
nor U43059 (N_43059,N_42681,N_42629);
and U43060 (N_43060,N_42890,N_42953);
xnor U43061 (N_43061,N_42973,N_42797);
or U43062 (N_43062,N_42940,N_42636);
xor U43063 (N_43063,N_42933,N_42870);
nor U43064 (N_43064,N_42631,N_42633);
nor U43065 (N_43065,N_42767,N_42846);
xnor U43066 (N_43066,N_42573,N_42746);
xor U43067 (N_43067,N_42536,N_42710);
nand U43068 (N_43068,N_42983,N_42865);
nand U43069 (N_43069,N_42569,N_42678);
xnor U43070 (N_43070,N_42612,N_42639);
and U43071 (N_43071,N_42853,N_42886);
nor U43072 (N_43072,N_42748,N_42819);
and U43073 (N_43073,N_42741,N_42707);
and U43074 (N_43074,N_42630,N_42802);
xnor U43075 (N_43075,N_42532,N_42542);
nor U43076 (N_43076,N_42545,N_42702);
nand U43077 (N_43077,N_42752,N_42818);
and U43078 (N_43078,N_42727,N_42779);
nand U43079 (N_43079,N_42561,N_42673);
or U43080 (N_43080,N_42547,N_42978);
nor U43081 (N_43081,N_42745,N_42620);
or U43082 (N_43082,N_42904,N_42691);
nand U43083 (N_43083,N_42896,N_42971);
xnor U43084 (N_43084,N_42772,N_42621);
or U43085 (N_43085,N_42715,N_42515);
nand U43086 (N_43086,N_42851,N_42924);
or U43087 (N_43087,N_42638,N_42875);
or U43088 (N_43088,N_42793,N_42844);
and U43089 (N_43089,N_42543,N_42849);
nor U43090 (N_43090,N_42783,N_42694);
xnor U43091 (N_43091,N_42649,N_42724);
or U43092 (N_43092,N_42997,N_42607);
nor U43093 (N_43093,N_42525,N_42838);
nor U43094 (N_43094,N_42854,N_42634);
xor U43095 (N_43095,N_42720,N_42706);
and U43096 (N_43096,N_42655,N_42930);
or U43097 (N_43097,N_42943,N_42811);
xnor U43098 (N_43098,N_42882,N_42527);
and U43099 (N_43099,N_42946,N_42987);
nand U43100 (N_43100,N_42663,N_42726);
and U43101 (N_43101,N_42591,N_42575);
or U43102 (N_43102,N_42510,N_42764);
nand U43103 (N_43103,N_42857,N_42850);
or U43104 (N_43104,N_42909,N_42766);
nand U43105 (N_43105,N_42577,N_42986);
and U43106 (N_43106,N_42787,N_42883);
and U43107 (N_43107,N_42615,N_42822);
nand U43108 (N_43108,N_42961,N_42587);
nor U43109 (N_43109,N_42834,N_42778);
and U43110 (N_43110,N_42869,N_42756);
and U43111 (N_43111,N_42739,N_42893);
xor U43112 (N_43112,N_42852,N_42926);
or U43113 (N_43113,N_42826,N_42954);
xnor U43114 (N_43114,N_42770,N_42939);
or U43115 (N_43115,N_42661,N_42581);
or U43116 (N_43116,N_42680,N_42794);
xor U43117 (N_43117,N_42696,N_42967);
xor U43118 (N_43118,N_42703,N_42516);
xor U43119 (N_43119,N_42760,N_42754);
or U43120 (N_43120,N_42755,N_42892);
xor U43121 (N_43121,N_42664,N_42574);
and U43122 (N_43122,N_42985,N_42963);
or U43123 (N_43123,N_42669,N_42659);
nor U43124 (N_43124,N_42911,N_42613);
and U43125 (N_43125,N_42816,N_42860);
or U43126 (N_43126,N_42535,N_42935);
nand U43127 (N_43127,N_42677,N_42572);
or U43128 (N_43128,N_42872,N_42716);
nand U43129 (N_43129,N_42975,N_42502);
nor U43130 (N_43130,N_42845,N_42606);
nand U43131 (N_43131,N_42551,N_42879);
and U43132 (N_43132,N_42627,N_42683);
xor U43133 (N_43133,N_42698,N_42984);
or U43134 (N_43134,N_42898,N_42648);
nor U43135 (N_43135,N_42919,N_42597);
and U43136 (N_43136,N_42762,N_42820);
xor U43137 (N_43137,N_42642,N_42711);
xor U43138 (N_43138,N_42936,N_42734);
xnor U43139 (N_43139,N_42517,N_42830);
nor U43140 (N_43140,N_42768,N_42803);
xor U43141 (N_43141,N_42611,N_42810);
nor U43142 (N_43142,N_42582,N_42538);
xnor U43143 (N_43143,N_42950,N_42513);
and U43144 (N_43144,N_42991,N_42774);
nand U43145 (N_43145,N_42580,N_42646);
xnor U43146 (N_43146,N_42829,N_42880);
nand U43147 (N_43147,N_42733,N_42956);
or U43148 (N_43148,N_42796,N_42804);
and U43149 (N_43149,N_42567,N_42812);
nor U43150 (N_43150,N_42623,N_42558);
xor U43151 (N_43151,N_42858,N_42566);
and U43152 (N_43152,N_42722,N_42996);
or U43153 (N_43153,N_42520,N_42578);
xnor U43154 (N_43154,N_42895,N_42709);
or U43155 (N_43155,N_42824,N_42656);
or U43156 (N_43156,N_42993,N_42721);
and U43157 (N_43157,N_42676,N_42785);
nor U43158 (N_43158,N_42625,N_42900);
and U43159 (N_43159,N_42738,N_42624);
and U43160 (N_43160,N_42757,N_42554);
xnor U43161 (N_43161,N_42807,N_42708);
xnor U43162 (N_43162,N_42714,N_42552);
and U43163 (N_43163,N_42941,N_42643);
xnor U43164 (N_43164,N_42583,N_42563);
and U43165 (N_43165,N_42828,N_42989);
xor U43166 (N_43166,N_42885,N_42539);
nand U43167 (N_43167,N_42862,N_42861);
nor U43168 (N_43168,N_42622,N_42966);
nand U43169 (N_43169,N_42522,N_42747);
or U43170 (N_43170,N_42749,N_42934);
xnor U43171 (N_43171,N_42640,N_42641);
and U43172 (N_43172,N_42602,N_42692);
xor U43173 (N_43173,N_42560,N_42524);
nor U43174 (N_43174,N_42777,N_42808);
or U43175 (N_43175,N_42668,N_42675);
xnor U43176 (N_43176,N_42679,N_42856);
nand U43177 (N_43177,N_42601,N_42603);
and U43178 (N_43178,N_42780,N_42541);
or U43179 (N_43179,N_42562,N_42876);
xnor U43180 (N_43180,N_42723,N_42590);
nand U43181 (N_43181,N_42564,N_42938);
xor U43182 (N_43182,N_42610,N_42593);
xnor U43183 (N_43183,N_42763,N_42942);
and U43184 (N_43184,N_42594,N_42994);
and U43185 (N_43185,N_42827,N_42928);
nor U43186 (N_43186,N_42902,N_42847);
xor U43187 (N_43187,N_42866,N_42660);
or U43188 (N_43188,N_42713,N_42507);
or U43189 (N_43189,N_42958,N_42670);
xnor U43190 (N_43190,N_42731,N_42921);
xnor U43191 (N_43191,N_42916,N_42899);
or U43192 (N_43192,N_42500,N_42537);
or U43193 (N_43193,N_42742,N_42521);
and U43194 (N_43194,N_42873,N_42799);
nor U43195 (N_43195,N_42871,N_42700);
nor U43196 (N_43196,N_42565,N_42549);
nand U43197 (N_43197,N_42951,N_42931);
xor U43198 (N_43198,N_42528,N_42666);
nand U43199 (N_43199,N_42753,N_42998);
xor U43200 (N_43200,N_42652,N_42689);
and U43201 (N_43201,N_42509,N_42867);
nand U43202 (N_43202,N_42868,N_42608);
and U43203 (N_43203,N_42728,N_42798);
nor U43204 (N_43204,N_42688,N_42927);
and U43205 (N_43205,N_42605,N_42775);
xor U43206 (N_43206,N_42781,N_42908);
and U43207 (N_43207,N_42571,N_42972);
xnor U43208 (N_43208,N_42685,N_42965);
xnor U43209 (N_43209,N_42506,N_42806);
nand U43210 (N_43210,N_42761,N_42585);
xor U43211 (N_43211,N_42529,N_42736);
nand U43212 (N_43212,N_42599,N_42995);
or U43213 (N_43213,N_42672,N_42977);
and U43214 (N_43214,N_42809,N_42948);
nand U43215 (N_43215,N_42877,N_42699);
nand U43216 (N_43216,N_42907,N_42682);
nand U43217 (N_43217,N_42651,N_42964);
nor U43218 (N_43218,N_42863,N_42697);
and U43219 (N_43219,N_42586,N_42550);
nor U43220 (N_43220,N_42667,N_42674);
nor U43221 (N_43221,N_42805,N_42732);
nand U43222 (N_43222,N_42962,N_42792);
and U43223 (N_43223,N_42982,N_42595);
nor U43224 (N_43224,N_42835,N_42949);
xnor U43225 (N_43225,N_42553,N_42815);
or U43226 (N_43226,N_42619,N_42788);
and U43227 (N_43227,N_42960,N_42616);
nor U43228 (N_43228,N_42584,N_42695);
nand U43229 (N_43229,N_42859,N_42801);
nor U43230 (N_43230,N_42887,N_42504);
and U43231 (N_43231,N_42508,N_42912);
and U43232 (N_43232,N_42906,N_42855);
and U43233 (N_43233,N_42635,N_42730);
xnor U43234 (N_43234,N_42523,N_42645);
or U43235 (N_43235,N_42718,N_42570);
nor U43236 (N_43236,N_42531,N_42650);
nor U43237 (N_43237,N_42548,N_42884);
and U43238 (N_43238,N_42821,N_42526);
and U43239 (N_43239,N_42980,N_42970);
or U43240 (N_43240,N_42917,N_42658);
or U43241 (N_43241,N_42947,N_42701);
nor U43242 (N_43242,N_42559,N_42915);
nand U43243 (N_43243,N_42952,N_42751);
nand U43244 (N_43244,N_42878,N_42519);
nor U43245 (N_43245,N_42758,N_42843);
and U43246 (N_43246,N_42999,N_42530);
xor U43247 (N_43247,N_42903,N_42817);
nor U43248 (N_43248,N_42546,N_42959);
nor U43249 (N_43249,N_42914,N_42684);
or U43250 (N_43250,N_42787,N_42888);
and U43251 (N_43251,N_42996,N_42660);
xnor U43252 (N_43252,N_42811,N_42973);
and U43253 (N_43253,N_42694,N_42511);
nand U43254 (N_43254,N_42723,N_42512);
nor U43255 (N_43255,N_42766,N_42763);
and U43256 (N_43256,N_42974,N_42567);
and U43257 (N_43257,N_42586,N_42546);
nor U43258 (N_43258,N_42952,N_42934);
xnor U43259 (N_43259,N_42659,N_42792);
xnor U43260 (N_43260,N_42558,N_42865);
nand U43261 (N_43261,N_42930,N_42514);
nor U43262 (N_43262,N_42600,N_42655);
and U43263 (N_43263,N_42692,N_42985);
nor U43264 (N_43264,N_42657,N_42623);
and U43265 (N_43265,N_42728,N_42889);
and U43266 (N_43266,N_42645,N_42726);
and U43267 (N_43267,N_42674,N_42848);
and U43268 (N_43268,N_42946,N_42552);
nor U43269 (N_43269,N_42506,N_42641);
xor U43270 (N_43270,N_42591,N_42568);
xor U43271 (N_43271,N_42740,N_42774);
nand U43272 (N_43272,N_42892,N_42636);
and U43273 (N_43273,N_42696,N_42912);
or U43274 (N_43274,N_42645,N_42826);
and U43275 (N_43275,N_42904,N_42708);
nand U43276 (N_43276,N_42694,N_42548);
xor U43277 (N_43277,N_42920,N_42676);
nand U43278 (N_43278,N_42775,N_42668);
or U43279 (N_43279,N_42706,N_42748);
xor U43280 (N_43280,N_42686,N_42848);
nand U43281 (N_43281,N_42872,N_42884);
nor U43282 (N_43282,N_42561,N_42586);
and U43283 (N_43283,N_42974,N_42546);
or U43284 (N_43284,N_42566,N_42532);
or U43285 (N_43285,N_42772,N_42698);
and U43286 (N_43286,N_42865,N_42883);
xnor U43287 (N_43287,N_42996,N_42868);
nand U43288 (N_43288,N_42751,N_42723);
nor U43289 (N_43289,N_42721,N_42931);
nor U43290 (N_43290,N_42891,N_42774);
nand U43291 (N_43291,N_42743,N_42916);
xor U43292 (N_43292,N_42720,N_42772);
nand U43293 (N_43293,N_42568,N_42777);
or U43294 (N_43294,N_42690,N_42650);
or U43295 (N_43295,N_42819,N_42650);
nand U43296 (N_43296,N_42545,N_42782);
and U43297 (N_43297,N_42986,N_42991);
xor U43298 (N_43298,N_42963,N_42955);
xor U43299 (N_43299,N_42691,N_42962);
xnor U43300 (N_43300,N_42641,N_42847);
nor U43301 (N_43301,N_42522,N_42532);
nand U43302 (N_43302,N_42960,N_42865);
nor U43303 (N_43303,N_42501,N_42731);
or U43304 (N_43304,N_42872,N_42623);
or U43305 (N_43305,N_42566,N_42743);
nor U43306 (N_43306,N_42703,N_42665);
and U43307 (N_43307,N_42598,N_42664);
xnor U43308 (N_43308,N_42963,N_42757);
nor U43309 (N_43309,N_42585,N_42934);
or U43310 (N_43310,N_42882,N_42859);
xnor U43311 (N_43311,N_42840,N_42890);
xor U43312 (N_43312,N_42880,N_42571);
nand U43313 (N_43313,N_42568,N_42862);
xnor U43314 (N_43314,N_42993,N_42672);
or U43315 (N_43315,N_42567,N_42679);
nor U43316 (N_43316,N_42685,N_42802);
nand U43317 (N_43317,N_42782,N_42564);
nand U43318 (N_43318,N_42625,N_42768);
xor U43319 (N_43319,N_42752,N_42873);
nand U43320 (N_43320,N_42542,N_42836);
xor U43321 (N_43321,N_42619,N_42845);
xnor U43322 (N_43322,N_42597,N_42677);
xnor U43323 (N_43323,N_42607,N_42748);
xnor U43324 (N_43324,N_42568,N_42540);
nand U43325 (N_43325,N_42760,N_42743);
and U43326 (N_43326,N_42794,N_42550);
or U43327 (N_43327,N_42712,N_42600);
xnor U43328 (N_43328,N_42947,N_42656);
nor U43329 (N_43329,N_42725,N_42595);
and U43330 (N_43330,N_42650,N_42885);
xor U43331 (N_43331,N_42999,N_42575);
and U43332 (N_43332,N_42659,N_42911);
xnor U43333 (N_43333,N_42535,N_42505);
or U43334 (N_43334,N_42544,N_42506);
nor U43335 (N_43335,N_42584,N_42747);
nor U43336 (N_43336,N_42640,N_42506);
or U43337 (N_43337,N_42920,N_42567);
or U43338 (N_43338,N_42755,N_42523);
xnor U43339 (N_43339,N_42563,N_42946);
nand U43340 (N_43340,N_42722,N_42675);
xor U43341 (N_43341,N_42705,N_42870);
and U43342 (N_43342,N_42684,N_42635);
and U43343 (N_43343,N_42692,N_42638);
and U43344 (N_43344,N_42805,N_42502);
nand U43345 (N_43345,N_42876,N_42546);
or U43346 (N_43346,N_42872,N_42639);
and U43347 (N_43347,N_42747,N_42890);
or U43348 (N_43348,N_42566,N_42919);
nor U43349 (N_43349,N_42826,N_42600);
xor U43350 (N_43350,N_42755,N_42714);
or U43351 (N_43351,N_42843,N_42741);
nor U43352 (N_43352,N_42800,N_42762);
or U43353 (N_43353,N_42960,N_42932);
and U43354 (N_43354,N_42839,N_42985);
and U43355 (N_43355,N_42756,N_42859);
and U43356 (N_43356,N_42590,N_42838);
nand U43357 (N_43357,N_42573,N_42807);
and U43358 (N_43358,N_42609,N_42900);
nor U43359 (N_43359,N_42562,N_42929);
nor U43360 (N_43360,N_42732,N_42596);
and U43361 (N_43361,N_42602,N_42950);
and U43362 (N_43362,N_42786,N_42666);
nor U43363 (N_43363,N_42558,N_42741);
xor U43364 (N_43364,N_42953,N_42669);
nand U43365 (N_43365,N_42796,N_42562);
nor U43366 (N_43366,N_42903,N_42856);
nand U43367 (N_43367,N_42528,N_42581);
nand U43368 (N_43368,N_42874,N_42818);
or U43369 (N_43369,N_42688,N_42520);
or U43370 (N_43370,N_42762,N_42795);
nand U43371 (N_43371,N_42855,N_42988);
and U43372 (N_43372,N_42681,N_42715);
nor U43373 (N_43373,N_42537,N_42898);
or U43374 (N_43374,N_42995,N_42854);
and U43375 (N_43375,N_42739,N_42652);
nor U43376 (N_43376,N_42849,N_42972);
or U43377 (N_43377,N_42551,N_42754);
and U43378 (N_43378,N_42753,N_42969);
and U43379 (N_43379,N_42651,N_42937);
nand U43380 (N_43380,N_42874,N_42599);
and U43381 (N_43381,N_42932,N_42612);
and U43382 (N_43382,N_42769,N_42728);
nor U43383 (N_43383,N_42994,N_42794);
nor U43384 (N_43384,N_42740,N_42683);
nand U43385 (N_43385,N_42895,N_42633);
nand U43386 (N_43386,N_42502,N_42685);
nor U43387 (N_43387,N_42887,N_42737);
xor U43388 (N_43388,N_42532,N_42844);
nand U43389 (N_43389,N_42594,N_42736);
nor U43390 (N_43390,N_42654,N_42665);
xor U43391 (N_43391,N_42910,N_42942);
and U43392 (N_43392,N_42973,N_42673);
xnor U43393 (N_43393,N_42645,N_42792);
and U43394 (N_43394,N_42810,N_42831);
nor U43395 (N_43395,N_42646,N_42850);
xor U43396 (N_43396,N_42827,N_42858);
nor U43397 (N_43397,N_42857,N_42509);
nand U43398 (N_43398,N_42827,N_42775);
xor U43399 (N_43399,N_42896,N_42897);
nor U43400 (N_43400,N_42613,N_42599);
nand U43401 (N_43401,N_42791,N_42973);
nor U43402 (N_43402,N_42590,N_42622);
xnor U43403 (N_43403,N_42595,N_42708);
nand U43404 (N_43404,N_42616,N_42820);
or U43405 (N_43405,N_42806,N_42757);
nor U43406 (N_43406,N_42519,N_42760);
and U43407 (N_43407,N_42607,N_42634);
nand U43408 (N_43408,N_42764,N_42615);
or U43409 (N_43409,N_42888,N_42899);
nand U43410 (N_43410,N_42785,N_42610);
or U43411 (N_43411,N_42768,N_42789);
or U43412 (N_43412,N_42613,N_42537);
nand U43413 (N_43413,N_42923,N_42788);
and U43414 (N_43414,N_42671,N_42645);
nand U43415 (N_43415,N_42647,N_42580);
nor U43416 (N_43416,N_42636,N_42965);
nor U43417 (N_43417,N_42865,N_42520);
nand U43418 (N_43418,N_42952,N_42704);
nor U43419 (N_43419,N_42974,N_42561);
or U43420 (N_43420,N_42676,N_42619);
xnor U43421 (N_43421,N_42630,N_42870);
or U43422 (N_43422,N_42624,N_42960);
xor U43423 (N_43423,N_42991,N_42538);
nor U43424 (N_43424,N_42803,N_42655);
or U43425 (N_43425,N_42979,N_42666);
xnor U43426 (N_43426,N_42621,N_42518);
or U43427 (N_43427,N_42501,N_42939);
or U43428 (N_43428,N_42564,N_42667);
nor U43429 (N_43429,N_42874,N_42654);
and U43430 (N_43430,N_42910,N_42818);
nor U43431 (N_43431,N_42510,N_42714);
nand U43432 (N_43432,N_42570,N_42541);
and U43433 (N_43433,N_42916,N_42865);
and U43434 (N_43434,N_42889,N_42886);
or U43435 (N_43435,N_42832,N_42926);
xnor U43436 (N_43436,N_42884,N_42895);
nor U43437 (N_43437,N_42566,N_42541);
and U43438 (N_43438,N_42695,N_42777);
or U43439 (N_43439,N_42602,N_42641);
or U43440 (N_43440,N_42889,N_42682);
nor U43441 (N_43441,N_42906,N_42784);
nor U43442 (N_43442,N_42661,N_42794);
xor U43443 (N_43443,N_42529,N_42907);
xor U43444 (N_43444,N_42938,N_42809);
nor U43445 (N_43445,N_42925,N_42714);
xor U43446 (N_43446,N_42974,N_42597);
nand U43447 (N_43447,N_42767,N_42815);
nor U43448 (N_43448,N_42821,N_42834);
and U43449 (N_43449,N_42595,N_42543);
or U43450 (N_43450,N_42575,N_42735);
nand U43451 (N_43451,N_42797,N_42985);
and U43452 (N_43452,N_42907,N_42554);
nor U43453 (N_43453,N_42623,N_42844);
and U43454 (N_43454,N_42519,N_42962);
and U43455 (N_43455,N_42980,N_42561);
nor U43456 (N_43456,N_42665,N_42534);
or U43457 (N_43457,N_42784,N_42806);
or U43458 (N_43458,N_42616,N_42831);
and U43459 (N_43459,N_42702,N_42905);
or U43460 (N_43460,N_42554,N_42815);
nor U43461 (N_43461,N_42612,N_42844);
xnor U43462 (N_43462,N_42779,N_42830);
xor U43463 (N_43463,N_42797,N_42895);
nor U43464 (N_43464,N_42697,N_42854);
nand U43465 (N_43465,N_42996,N_42865);
xor U43466 (N_43466,N_42627,N_42563);
nand U43467 (N_43467,N_42908,N_42868);
and U43468 (N_43468,N_42689,N_42982);
and U43469 (N_43469,N_42949,N_42873);
xor U43470 (N_43470,N_42614,N_42704);
nand U43471 (N_43471,N_42551,N_42793);
or U43472 (N_43472,N_42541,N_42705);
or U43473 (N_43473,N_42567,N_42738);
or U43474 (N_43474,N_42869,N_42981);
or U43475 (N_43475,N_42526,N_42561);
nor U43476 (N_43476,N_42529,N_42508);
nand U43477 (N_43477,N_42718,N_42534);
xnor U43478 (N_43478,N_42699,N_42601);
xnor U43479 (N_43479,N_42905,N_42710);
nor U43480 (N_43480,N_42590,N_42669);
and U43481 (N_43481,N_42723,N_42818);
and U43482 (N_43482,N_42600,N_42558);
or U43483 (N_43483,N_42750,N_42924);
or U43484 (N_43484,N_42590,N_42948);
nor U43485 (N_43485,N_42868,N_42579);
nand U43486 (N_43486,N_42999,N_42923);
nand U43487 (N_43487,N_42539,N_42553);
nand U43488 (N_43488,N_42693,N_42912);
and U43489 (N_43489,N_42815,N_42512);
or U43490 (N_43490,N_42527,N_42638);
nand U43491 (N_43491,N_42873,N_42690);
xnor U43492 (N_43492,N_42996,N_42696);
and U43493 (N_43493,N_42750,N_42833);
and U43494 (N_43494,N_42520,N_42506);
nand U43495 (N_43495,N_42730,N_42694);
and U43496 (N_43496,N_42518,N_42540);
xor U43497 (N_43497,N_42552,N_42997);
or U43498 (N_43498,N_42803,N_42834);
and U43499 (N_43499,N_42919,N_42605);
xnor U43500 (N_43500,N_43191,N_43014);
nand U43501 (N_43501,N_43017,N_43371);
nand U43502 (N_43502,N_43060,N_43296);
nor U43503 (N_43503,N_43265,N_43161);
or U43504 (N_43504,N_43271,N_43001);
or U43505 (N_43505,N_43426,N_43402);
or U43506 (N_43506,N_43247,N_43368);
xor U43507 (N_43507,N_43420,N_43338);
nor U43508 (N_43508,N_43168,N_43477);
nor U43509 (N_43509,N_43388,N_43107);
nand U43510 (N_43510,N_43150,N_43479);
nand U43511 (N_43511,N_43429,N_43404);
and U43512 (N_43512,N_43092,N_43074);
xnor U43513 (N_43513,N_43177,N_43389);
nand U43514 (N_43514,N_43323,N_43185);
nor U43515 (N_43515,N_43039,N_43237);
nor U43516 (N_43516,N_43147,N_43026);
and U43517 (N_43517,N_43085,N_43448);
nor U43518 (N_43518,N_43197,N_43311);
or U43519 (N_43519,N_43061,N_43236);
xnor U43520 (N_43520,N_43469,N_43254);
nand U43521 (N_43521,N_43359,N_43342);
nor U43522 (N_43522,N_43041,N_43360);
nand U43523 (N_43523,N_43203,N_43437);
or U43524 (N_43524,N_43210,N_43123);
and U43525 (N_43525,N_43332,N_43183);
or U43526 (N_43526,N_43385,N_43246);
nor U43527 (N_43527,N_43013,N_43187);
xor U43528 (N_43528,N_43459,N_43294);
nand U43529 (N_43529,N_43053,N_43347);
and U43530 (N_43530,N_43225,N_43489);
nor U43531 (N_43531,N_43495,N_43078);
or U43532 (N_43532,N_43252,N_43015);
xor U43533 (N_43533,N_43467,N_43021);
and U43534 (N_43534,N_43255,N_43005);
and U43535 (N_43535,N_43067,N_43444);
nand U43536 (N_43536,N_43029,N_43488);
nand U43537 (N_43537,N_43322,N_43240);
nor U43538 (N_43538,N_43214,N_43220);
or U43539 (N_43539,N_43167,N_43233);
or U43540 (N_43540,N_43358,N_43414);
and U43541 (N_43541,N_43163,N_43179);
nand U43542 (N_43542,N_43372,N_43059);
nand U43543 (N_43543,N_43226,N_43186);
nor U43544 (N_43544,N_43086,N_43139);
and U43545 (N_43545,N_43260,N_43160);
and U43546 (N_43546,N_43111,N_43457);
and U43547 (N_43547,N_43090,N_43124);
or U43548 (N_43548,N_43058,N_43280);
or U43549 (N_43549,N_43416,N_43082);
or U43550 (N_43550,N_43487,N_43242);
xor U43551 (N_43551,N_43312,N_43142);
xnor U43552 (N_43552,N_43284,N_43266);
xor U43553 (N_43553,N_43480,N_43386);
xnor U43554 (N_43554,N_43004,N_43132);
nand U43555 (N_43555,N_43096,N_43496);
xor U43556 (N_43556,N_43317,N_43106);
nor U43557 (N_43557,N_43138,N_43318);
nor U43558 (N_43558,N_43439,N_43465);
or U43559 (N_43559,N_43057,N_43498);
xnor U43560 (N_43560,N_43329,N_43049);
or U43561 (N_43561,N_43178,N_43116);
or U43562 (N_43562,N_43434,N_43171);
and U43563 (N_43563,N_43355,N_43063);
or U43564 (N_43564,N_43016,N_43231);
and U43565 (N_43565,N_43308,N_43449);
or U43566 (N_43566,N_43056,N_43069);
and U43567 (N_43567,N_43095,N_43274);
nor U43568 (N_43568,N_43070,N_43158);
xnor U43569 (N_43569,N_43114,N_43065);
and U43570 (N_43570,N_43129,N_43042);
and U43571 (N_43571,N_43257,N_43390);
nand U43572 (N_43572,N_43451,N_43102);
xnor U43573 (N_43573,N_43028,N_43412);
and U43574 (N_43574,N_43267,N_43230);
nor U43575 (N_43575,N_43221,N_43273);
nand U43576 (N_43576,N_43201,N_43173);
xnor U43577 (N_43577,N_43241,N_43346);
nand U43578 (N_43578,N_43364,N_43224);
nand U43579 (N_43579,N_43184,N_43165);
xnor U43580 (N_43580,N_43394,N_43407);
xnor U43581 (N_43581,N_43409,N_43403);
nand U43582 (N_43582,N_43418,N_43339);
nor U43583 (N_43583,N_43471,N_43034);
and U43584 (N_43584,N_43120,N_43227);
or U43585 (N_43585,N_43464,N_43326);
nor U43586 (N_43586,N_43204,N_43283);
or U43587 (N_43587,N_43245,N_43474);
and U43588 (N_43588,N_43356,N_43345);
or U43589 (N_43589,N_43212,N_43126);
xnor U43590 (N_43590,N_43192,N_43431);
xnor U43591 (N_43591,N_43277,N_43103);
or U43592 (N_43592,N_43009,N_43081);
or U43593 (N_43593,N_43232,N_43239);
and U43594 (N_43594,N_43045,N_43417);
or U43595 (N_43595,N_43050,N_43478);
nor U43596 (N_43596,N_43482,N_43238);
nor U43597 (N_43597,N_43020,N_43046);
or U43598 (N_43598,N_43286,N_43316);
nor U43599 (N_43599,N_43290,N_43335);
and U43600 (N_43600,N_43089,N_43181);
nand U43601 (N_43601,N_43441,N_43458);
nand U43602 (N_43602,N_43195,N_43327);
xnor U43603 (N_43603,N_43475,N_43117);
nand U43604 (N_43604,N_43091,N_43052);
nand U43605 (N_43605,N_43189,N_43164);
or U43606 (N_43606,N_43098,N_43032);
xnor U43607 (N_43607,N_43401,N_43313);
nand U43608 (N_43608,N_43218,N_43293);
or U43609 (N_43609,N_43456,N_43024);
xor U43610 (N_43610,N_43405,N_43300);
nand U43611 (N_43611,N_43397,N_43235);
nand U43612 (N_43612,N_43447,N_43190);
and U43613 (N_43613,N_43208,N_43250);
nor U43614 (N_43614,N_43440,N_43248);
nand U43615 (N_43615,N_43154,N_43331);
xnor U43616 (N_43616,N_43088,N_43199);
xor U43617 (N_43617,N_43392,N_43118);
nor U43618 (N_43618,N_43442,N_43380);
nor U43619 (N_43619,N_43149,N_43217);
nor U43620 (N_43620,N_43051,N_43262);
or U43621 (N_43621,N_43193,N_43310);
nand U43622 (N_43622,N_43428,N_43320);
nand U43623 (N_43623,N_43472,N_43340);
or U43624 (N_43624,N_43100,N_43087);
nand U43625 (N_43625,N_43206,N_43383);
or U43626 (N_43626,N_43152,N_43258);
or U43627 (N_43627,N_43452,N_43337);
nand U43628 (N_43628,N_43194,N_43130);
or U43629 (N_43629,N_43427,N_43175);
or U43630 (N_43630,N_43443,N_43270);
nor U43631 (N_43631,N_43170,N_43490);
xor U43632 (N_43632,N_43162,N_43373);
nand U43633 (N_43633,N_43446,N_43285);
or U43634 (N_43634,N_43291,N_43297);
or U43635 (N_43635,N_43330,N_43461);
nor U43636 (N_43636,N_43476,N_43068);
xor U43637 (N_43637,N_43011,N_43148);
or U43638 (N_43638,N_43319,N_43146);
nor U43639 (N_43639,N_43127,N_43044);
nor U43640 (N_43640,N_43176,N_43137);
nor U43641 (N_43641,N_43205,N_43494);
and U43642 (N_43642,N_43104,N_43305);
nand U43643 (N_43643,N_43048,N_43083);
and U43644 (N_43644,N_43306,N_43351);
nor U43645 (N_43645,N_43419,N_43307);
xor U43646 (N_43646,N_43315,N_43435);
nand U43647 (N_43647,N_43491,N_43309);
nor U43648 (N_43648,N_43462,N_43415);
and U43649 (N_43649,N_43492,N_43037);
nand U43650 (N_43650,N_43282,N_43030);
nor U43651 (N_43651,N_43425,N_43357);
or U43652 (N_43652,N_43387,N_43354);
and U43653 (N_43653,N_43002,N_43486);
xor U43654 (N_43654,N_43157,N_43134);
and U43655 (N_43655,N_43093,N_43097);
nand U43656 (N_43656,N_43349,N_43400);
and U43657 (N_43657,N_43122,N_43279);
nand U43658 (N_43658,N_43314,N_43003);
nand U43659 (N_43659,N_43408,N_43369);
nor U43660 (N_43660,N_43376,N_43450);
and U43661 (N_43661,N_43196,N_43244);
nand U43662 (N_43662,N_43382,N_43151);
or U43663 (N_43663,N_43341,N_43207);
nand U43664 (N_43664,N_43343,N_43430);
nand U43665 (N_43665,N_43144,N_43406);
nor U43666 (N_43666,N_43396,N_43422);
nand U43667 (N_43667,N_43047,N_43135);
and U43668 (N_43668,N_43384,N_43010);
nor U43669 (N_43669,N_43287,N_43366);
or U43670 (N_43670,N_43333,N_43453);
and U43671 (N_43671,N_43054,N_43182);
nand U43672 (N_43672,N_43423,N_43027);
xnor U43673 (N_43673,N_43460,N_43229);
nand U43674 (N_43674,N_43038,N_43302);
nor U43675 (N_43675,N_43136,N_43261);
and U43676 (N_43676,N_43370,N_43121);
nand U43677 (N_43677,N_43140,N_43075);
or U43678 (N_43678,N_43499,N_43363);
xor U43679 (N_43679,N_43421,N_43484);
and U43680 (N_43680,N_43145,N_43399);
nor U43681 (N_43681,N_43361,N_43278);
and U43682 (N_43682,N_43473,N_43115);
or U43683 (N_43683,N_43200,N_43012);
nor U43684 (N_43684,N_43172,N_43379);
nor U43685 (N_43685,N_43295,N_43253);
nand U43686 (N_43686,N_43216,N_43497);
xnor U43687 (N_43687,N_43481,N_43128);
nor U43688 (N_43688,N_43375,N_43228);
nand U43689 (N_43689,N_43485,N_43299);
xor U43690 (N_43690,N_43256,N_43019);
nor U43691 (N_43691,N_43289,N_43031);
or U43692 (N_43692,N_43022,N_43040);
xor U43693 (N_43693,N_43259,N_43143);
nand U43694 (N_43694,N_43395,N_43410);
nand U43695 (N_43695,N_43109,N_43432);
nand U43696 (N_43696,N_43378,N_43202);
or U43697 (N_43697,N_43119,N_43105);
nand U43698 (N_43698,N_43209,N_43094);
xor U43699 (N_43699,N_43281,N_43080);
nor U43700 (N_43700,N_43374,N_43263);
xnor U43701 (N_43701,N_43141,N_43264);
xnor U43702 (N_43702,N_43324,N_43269);
and U43703 (N_43703,N_43188,N_43398);
or U43704 (N_43704,N_43072,N_43219);
and U43705 (N_43705,N_43084,N_43159);
or U43706 (N_43706,N_43073,N_43077);
xor U43707 (N_43707,N_43099,N_43303);
nand U43708 (N_43708,N_43362,N_43234);
xnor U43709 (N_43709,N_43468,N_43463);
nand U43710 (N_43710,N_43352,N_43301);
xnor U43711 (N_43711,N_43025,N_43125);
nand U43712 (N_43712,N_43008,N_43445);
and U43713 (N_43713,N_43292,N_43062);
or U43714 (N_43714,N_43043,N_43079);
nor U43715 (N_43715,N_43064,N_43391);
and U43716 (N_43716,N_43156,N_43174);
and U43717 (N_43717,N_43466,N_43036);
and U43718 (N_43718,N_43436,N_43413);
nand U43719 (N_43719,N_43493,N_43000);
or U43720 (N_43720,N_43424,N_43275);
nor U43721 (N_43721,N_43110,N_43006);
nand U43722 (N_43722,N_43033,N_43298);
nor U43723 (N_43723,N_43113,N_43433);
or U43724 (N_43724,N_43411,N_43344);
nand U43725 (N_43725,N_43334,N_43243);
or U43726 (N_43726,N_43350,N_43018);
nand U43727 (N_43727,N_43223,N_43325);
and U43728 (N_43728,N_43288,N_43076);
or U43729 (N_43729,N_43055,N_43071);
nand U43730 (N_43730,N_43249,N_43169);
nor U43731 (N_43731,N_43365,N_43023);
or U43732 (N_43732,N_43454,N_43348);
xor U43733 (N_43733,N_43166,N_43381);
xnor U43734 (N_43734,N_43066,N_43268);
xor U43735 (N_43735,N_43215,N_43377);
nor U43736 (N_43736,N_43108,N_43213);
and U43737 (N_43737,N_43035,N_43101);
nand U43738 (N_43738,N_43483,N_43198);
and U43739 (N_43739,N_43211,N_43455);
and U43740 (N_43740,N_43393,N_43112);
nand U43741 (N_43741,N_43133,N_43276);
nor U43742 (N_43742,N_43180,N_43155);
nand U43743 (N_43743,N_43367,N_43321);
xnor U43744 (N_43744,N_43328,N_43353);
xnor U43745 (N_43745,N_43251,N_43131);
and U43746 (N_43746,N_43272,N_43304);
or U43747 (N_43747,N_43470,N_43153);
xor U43748 (N_43748,N_43438,N_43007);
nand U43749 (N_43749,N_43336,N_43222);
or U43750 (N_43750,N_43281,N_43129);
nor U43751 (N_43751,N_43277,N_43172);
nand U43752 (N_43752,N_43055,N_43037);
nor U43753 (N_43753,N_43022,N_43138);
nor U43754 (N_43754,N_43083,N_43284);
and U43755 (N_43755,N_43258,N_43246);
or U43756 (N_43756,N_43460,N_43250);
xnor U43757 (N_43757,N_43430,N_43348);
or U43758 (N_43758,N_43027,N_43343);
nor U43759 (N_43759,N_43177,N_43181);
nand U43760 (N_43760,N_43290,N_43378);
xnor U43761 (N_43761,N_43146,N_43404);
and U43762 (N_43762,N_43312,N_43082);
or U43763 (N_43763,N_43256,N_43311);
nor U43764 (N_43764,N_43124,N_43285);
nand U43765 (N_43765,N_43497,N_43275);
nand U43766 (N_43766,N_43073,N_43268);
and U43767 (N_43767,N_43153,N_43499);
or U43768 (N_43768,N_43331,N_43487);
nor U43769 (N_43769,N_43237,N_43236);
nor U43770 (N_43770,N_43270,N_43205);
or U43771 (N_43771,N_43230,N_43436);
xnor U43772 (N_43772,N_43466,N_43025);
or U43773 (N_43773,N_43036,N_43271);
nor U43774 (N_43774,N_43258,N_43232);
or U43775 (N_43775,N_43452,N_43165);
xnor U43776 (N_43776,N_43182,N_43488);
xor U43777 (N_43777,N_43041,N_43014);
nand U43778 (N_43778,N_43135,N_43054);
xnor U43779 (N_43779,N_43096,N_43081);
nor U43780 (N_43780,N_43198,N_43495);
or U43781 (N_43781,N_43404,N_43224);
xnor U43782 (N_43782,N_43169,N_43308);
or U43783 (N_43783,N_43113,N_43363);
xor U43784 (N_43784,N_43142,N_43161);
and U43785 (N_43785,N_43224,N_43342);
and U43786 (N_43786,N_43224,N_43353);
nand U43787 (N_43787,N_43022,N_43122);
and U43788 (N_43788,N_43305,N_43288);
nand U43789 (N_43789,N_43054,N_43077);
nor U43790 (N_43790,N_43452,N_43403);
or U43791 (N_43791,N_43368,N_43417);
nand U43792 (N_43792,N_43296,N_43349);
or U43793 (N_43793,N_43313,N_43438);
or U43794 (N_43794,N_43457,N_43301);
and U43795 (N_43795,N_43007,N_43424);
nand U43796 (N_43796,N_43370,N_43419);
nand U43797 (N_43797,N_43023,N_43367);
nor U43798 (N_43798,N_43452,N_43245);
nand U43799 (N_43799,N_43357,N_43187);
and U43800 (N_43800,N_43084,N_43379);
nor U43801 (N_43801,N_43200,N_43281);
xor U43802 (N_43802,N_43320,N_43200);
nand U43803 (N_43803,N_43462,N_43410);
nor U43804 (N_43804,N_43436,N_43466);
or U43805 (N_43805,N_43171,N_43320);
nand U43806 (N_43806,N_43239,N_43495);
nand U43807 (N_43807,N_43186,N_43401);
nor U43808 (N_43808,N_43356,N_43273);
nor U43809 (N_43809,N_43115,N_43340);
nor U43810 (N_43810,N_43396,N_43065);
and U43811 (N_43811,N_43309,N_43378);
nor U43812 (N_43812,N_43324,N_43086);
or U43813 (N_43813,N_43090,N_43253);
and U43814 (N_43814,N_43076,N_43400);
and U43815 (N_43815,N_43232,N_43181);
nand U43816 (N_43816,N_43476,N_43411);
nand U43817 (N_43817,N_43442,N_43497);
nand U43818 (N_43818,N_43045,N_43181);
or U43819 (N_43819,N_43209,N_43138);
nand U43820 (N_43820,N_43130,N_43198);
nor U43821 (N_43821,N_43165,N_43025);
and U43822 (N_43822,N_43123,N_43147);
nor U43823 (N_43823,N_43219,N_43117);
nand U43824 (N_43824,N_43211,N_43320);
nor U43825 (N_43825,N_43297,N_43056);
xor U43826 (N_43826,N_43034,N_43210);
nand U43827 (N_43827,N_43405,N_43250);
and U43828 (N_43828,N_43221,N_43082);
nor U43829 (N_43829,N_43399,N_43483);
or U43830 (N_43830,N_43436,N_43074);
xor U43831 (N_43831,N_43416,N_43466);
nor U43832 (N_43832,N_43402,N_43131);
nand U43833 (N_43833,N_43059,N_43480);
and U43834 (N_43834,N_43100,N_43386);
xnor U43835 (N_43835,N_43269,N_43353);
nor U43836 (N_43836,N_43037,N_43345);
xor U43837 (N_43837,N_43033,N_43016);
xor U43838 (N_43838,N_43037,N_43042);
and U43839 (N_43839,N_43125,N_43213);
and U43840 (N_43840,N_43143,N_43198);
or U43841 (N_43841,N_43499,N_43221);
nand U43842 (N_43842,N_43089,N_43211);
nand U43843 (N_43843,N_43367,N_43287);
xor U43844 (N_43844,N_43299,N_43164);
and U43845 (N_43845,N_43362,N_43096);
or U43846 (N_43846,N_43178,N_43107);
xnor U43847 (N_43847,N_43248,N_43081);
nand U43848 (N_43848,N_43247,N_43374);
nor U43849 (N_43849,N_43333,N_43003);
nand U43850 (N_43850,N_43106,N_43143);
nor U43851 (N_43851,N_43448,N_43141);
or U43852 (N_43852,N_43093,N_43008);
nor U43853 (N_43853,N_43086,N_43140);
and U43854 (N_43854,N_43200,N_43475);
nand U43855 (N_43855,N_43480,N_43094);
xor U43856 (N_43856,N_43085,N_43017);
xor U43857 (N_43857,N_43087,N_43289);
or U43858 (N_43858,N_43424,N_43025);
and U43859 (N_43859,N_43168,N_43321);
nand U43860 (N_43860,N_43108,N_43036);
nor U43861 (N_43861,N_43178,N_43434);
or U43862 (N_43862,N_43460,N_43043);
nor U43863 (N_43863,N_43037,N_43224);
xnor U43864 (N_43864,N_43459,N_43088);
nor U43865 (N_43865,N_43303,N_43313);
nand U43866 (N_43866,N_43454,N_43269);
and U43867 (N_43867,N_43150,N_43363);
nor U43868 (N_43868,N_43156,N_43238);
or U43869 (N_43869,N_43043,N_43230);
nor U43870 (N_43870,N_43188,N_43299);
xor U43871 (N_43871,N_43275,N_43487);
nor U43872 (N_43872,N_43488,N_43020);
xor U43873 (N_43873,N_43461,N_43312);
nand U43874 (N_43874,N_43456,N_43207);
nor U43875 (N_43875,N_43102,N_43014);
nand U43876 (N_43876,N_43098,N_43311);
nor U43877 (N_43877,N_43449,N_43004);
and U43878 (N_43878,N_43104,N_43103);
or U43879 (N_43879,N_43284,N_43305);
xor U43880 (N_43880,N_43490,N_43210);
and U43881 (N_43881,N_43366,N_43046);
or U43882 (N_43882,N_43220,N_43467);
nand U43883 (N_43883,N_43245,N_43353);
xnor U43884 (N_43884,N_43171,N_43325);
xnor U43885 (N_43885,N_43389,N_43330);
and U43886 (N_43886,N_43487,N_43258);
nor U43887 (N_43887,N_43389,N_43139);
xnor U43888 (N_43888,N_43002,N_43462);
or U43889 (N_43889,N_43126,N_43362);
and U43890 (N_43890,N_43444,N_43325);
nor U43891 (N_43891,N_43434,N_43072);
or U43892 (N_43892,N_43108,N_43469);
or U43893 (N_43893,N_43154,N_43327);
nand U43894 (N_43894,N_43405,N_43034);
or U43895 (N_43895,N_43290,N_43047);
nand U43896 (N_43896,N_43482,N_43220);
nor U43897 (N_43897,N_43405,N_43198);
nor U43898 (N_43898,N_43416,N_43377);
and U43899 (N_43899,N_43436,N_43143);
and U43900 (N_43900,N_43137,N_43073);
and U43901 (N_43901,N_43218,N_43448);
or U43902 (N_43902,N_43175,N_43064);
xor U43903 (N_43903,N_43473,N_43072);
nor U43904 (N_43904,N_43258,N_43073);
nor U43905 (N_43905,N_43395,N_43102);
nand U43906 (N_43906,N_43103,N_43419);
nand U43907 (N_43907,N_43376,N_43192);
or U43908 (N_43908,N_43227,N_43398);
nand U43909 (N_43909,N_43310,N_43420);
or U43910 (N_43910,N_43281,N_43440);
xnor U43911 (N_43911,N_43093,N_43204);
or U43912 (N_43912,N_43470,N_43485);
xor U43913 (N_43913,N_43040,N_43225);
and U43914 (N_43914,N_43282,N_43250);
or U43915 (N_43915,N_43391,N_43483);
nor U43916 (N_43916,N_43038,N_43089);
nand U43917 (N_43917,N_43109,N_43134);
nand U43918 (N_43918,N_43136,N_43277);
nand U43919 (N_43919,N_43247,N_43443);
xor U43920 (N_43920,N_43090,N_43293);
nand U43921 (N_43921,N_43009,N_43256);
and U43922 (N_43922,N_43167,N_43253);
xor U43923 (N_43923,N_43414,N_43115);
xor U43924 (N_43924,N_43474,N_43134);
and U43925 (N_43925,N_43200,N_43313);
nand U43926 (N_43926,N_43105,N_43358);
and U43927 (N_43927,N_43227,N_43239);
and U43928 (N_43928,N_43242,N_43074);
nand U43929 (N_43929,N_43418,N_43092);
or U43930 (N_43930,N_43342,N_43117);
or U43931 (N_43931,N_43350,N_43397);
or U43932 (N_43932,N_43165,N_43417);
nor U43933 (N_43933,N_43167,N_43440);
or U43934 (N_43934,N_43117,N_43441);
nand U43935 (N_43935,N_43415,N_43178);
nor U43936 (N_43936,N_43350,N_43224);
and U43937 (N_43937,N_43306,N_43143);
xnor U43938 (N_43938,N_43267,N_43314);
nand U43939 (N_43939,N_43343,N_43063);
xnor U43940 (N_43940,N_43157,N_43003);
nor U43941 (N_43941,N_43267,N_43019);
xnor U43942 (N_43942,N_43055,N_43118);
xor U43943 (N_43943,N_43452,N_43353);
xor U43944 (N_43944,N_43287,N_43029);
nor U43945 (N_43945,N_43457,N_43497);
nor U43946 (N_43946,N_43389,N_43266);
xnor U43947 (N_43947,N_43003,N_43286);
or U43948 (N_43948,N_43309,N_43077);
nand U43949 (N_43949,N_43378,N_43457);
nor U43950 (N_43950,N_43273,N_43334);
nor U43951 (N_43951,N_43323,N_43199);
or U43952 (N_43952,N_43171,N_43218);
xnor U43953 (N_43953,N_43482,N_43182);
or U43954 (N_43954,N_43160,N_43375);
nand U43955 (N_43955,N_43288,N_43336);
or U43956 (N_43956,N_43079,N_43447);
or U43957 (N_43957,N_43052,N_43323);
nand U43958 (N_43958,N_43125,N_43244);
and U43959 (N_43959,N_43495,N_43301);
and U43960 (N_43960,N_43414,N_43274);
nor U43961 (N_43961,N_43305,N_43018);
nand U43962 (N_43962,N_43172,N_43161);
xor U43963 (N_43963,N_43139,N_43253);
and U43964 (N_43964,N_43238,N_43235);
xor U43965 (N_43965,N_43424,N_43124);
nor U43966 (N_43966,N_43101,N_43380);
nand U43967 (N_43967,N_43391,N_43301);
nand U43968 (N_43968,N_43267,N_43453);
xnor U43969 (N_43969,N_43449,N_43002);
nor U43970 (N_43970,N_43218,N_43388);
nand U43971 (N_43971,N_43108,N_43386);
nand U43972 (N_43972,N_43040,N_43070);
nand U43973 (N_43973,N_43154,N_43422);
nand U43974 (N_43974,N_43212,N_43333);
xor U43975 (N_43975,N_43402,N_43310);
nor U43976 (N_43976,N_43133,N_43012);
nor U43977 (N_43977,N_43156,N_43109);
and U43978 (N_43978,N_43140,N_43456);
or U43979 (N_43979,N_43278,N_43284);
nor U43980 (N_43980,N_43344,N_43270);
xnor U43981 (N_43981,N_43418,N_43036);
and U43982 (N_43982,N_43237,N_43235);
nand U43983 (N_43983,N_43445,N_43408);
nor U43984 (N_43984,N_43455,N_43497);
and U43985 (N_43985,N_43486,N_43354);
and U43986 (N_43986,N_43041,N_43402);
xor U43987 (N_43987,N_43054,N_43311);
or U43988 (N_43988,N_43430,N_43173);
nor U43989 (N_43989,N_43099,N_43179);
and U43990 (N_43990,N_43370,N_43474);
nor U43991 (N_43991,N_43149,N_43330);
xnor U43992 (N_43992,N_43113,N_43121);
or U43993 (N_43993,N_43105,N_43169);
xnor U43994 (N_43994,N_43326,N_43052);
nor U43995 (N_43995,N_43267,N_43290);
and U43996 (N_43996,N_43216,N_43116);
nand U43997 (N_43997,N_43300,N_43238);
nor U43998 (N_43998,N_43240,N_43133);
nor U43999 (N_43999,N_43083,N_43070);
or U44000 (N_44000,N_43748,N_43755);
nand U44001 (N_44001,N_43749,N_43840);
or U44002 (N_44002,N_43837,N_43998);
xnor U44003 (N_44003,N_43954,N_43574);
xor U44004 (N_44004,N_43780,N_43508);
and U44005 (N_44005,N_43532,N_43902);
or U44006 (N_44006,N_43945,N_43856);
and U44007 (N_44007,N_43866,N_43573);
or U44008 (N_44008,N_43632,N_43514);
nand U44009 (N_44009,N_43702,N_43623);
and U44010 (N_44010,N_43807,N_43772);
nand U44011 (N_44011,N_43579,N_43595);
and U44012 (N_44012,N_43751,N_43957);
xnor U44013 (N_44013,N_43987,N_43540);
and U44014 (N_44014,N_43504,N_43793);
nor U44015 (N_44015,N_43530,N_43737);
nor U44016 (N_44016,N_43534,N_43933);
nor U44017 (N_44017,N_43745,N_43691);
or U44018 (N_44018,N_43763,N_43712);
and U44019 (N_44019,N_43658,N_43792);
xnor U44020 (N_44020,N_43756,N_43606);
or U44021 (N_44021,N_43889,N_43580);
nor U44022 (N_44022,N_43668,N_43518);
or U44023 (N_44023,N_43929,N_43940);
xor U44024 (N_44024,N_43713,N_43890);
or U44025 (N_44025,N_43877,N_43551);
xnor U44026 (N_44026,N_43704,N_43636);
and U44027 (N_44027,N_43934,N_43932);
and U44028 (N_44028,N_43536,N_43562);
or U44029 (N_44029,N_43715,N_43999);
nor U44030 (N_44030,N_43685,N_43984);
xnor U44031 (N_44031,N_43621,N_43502);
nand U44032 (N_44032,N_43741,N_43589);
or U44033 (N_44033,N_43769,N_43523);
xor U44034 (N_44034,N_43863,N_43601);
xnor U44035 (N_44035,N_43787,N_43799);
nand U44036 (N_44036,N_43546,N_43868);
or U44037 (N_44037,N_43732,N_43927);
xor U44038 (N_44038,N_43622,N_43810);
nand U44039 (N_44039,N_43909,N_43812);
nand U44040 (N_44040,N_43572,N_43679);
nand U44041 (N_44041,N_43872,N_43645);
xor U44042 (N_44042,N_43914,N_43571);
xnor U44043 (N_44043,N_43823,N_43662);
or U44044 (N_44044,N_43758,N_43779);
nand U44045 (N_44045,N_43564,N_43528);
nor U44046 (N_44046,N_43790,N_43587);
nand U44047 (N_44047,N_43874,N_43838);
and U44048 (N_44048,N_43628,N_43777);
and U44049 (N_44049,N_43761,N_43603);
and U44050 (N_44050,N_43973,N_43541);
nand U44051 (N_44051,N_43674,N_43716);
or U44052 (N_44052,N_43706,N_43882);
and U44053 (N_44053,N_43859,N_43768);
and U44054 (N_44054,N_43633,N_43726);
nor U44055 (N_44055,N_43646,N_43510);
and U44056 (N_44056,N_43785,N_43576);
nand U44057 (N_44057,N_43888,N_43887);
xnor U44058 (N_44058,N_43854,N_43620);
and U44059 (N_44059,N_43550,N_43886);
and U44060 (N_44060,N_43958,N_43813);
and U44061 (N_44061,N_43804,N_43519);
nor U44062 (N_44062,N_43513,N_43870);
and U44063 (N_44063,N_43982,N_43588);
and U44064 (N_44064,N_43873,N_43664);
and U44065 (N_44065,N_43694,N_43986);
nor U44066 (N_44066,N_43656,N_43781);
and U44067 (N_44067,N_43944,N_43764);
and U44068 (N_44068,N_43831,N_43931);
or U44069 (N_44069,N_43778,N_43654);
xnor U44070 (N_44070,N_43962,N_43738);
xor U44071 (N_44071,N_43964,N_43730);
or U44072 (N_44072,N_43525,N_43891);
nor U44073 (N_44073,N_43667,N_43979);
nor U44074 (N_44074,N_43900,N_43832);
and U44075 (N_44075,N_43757,N_43577);
or U44076 (N_44076,N_43695,N_43553);
or U44077 (N_44077,N_43683,N_43729);
or U44078 (N_44078,N_43592,N_43836);
nor U44079 (N_44079,N_43630,N_43742);
or U44080 (N_44080,N_43844,N_43727);
nor U44081 (N_44081,N_43817,N_43599);
nor U44082 (N_44082,N_43517,N_43901);
xnor U44083 (N_44083,N_43545,N_43903);
and U44084 (N_44084,N_43642,N_43770);
or U44085 (N_44085,N_43723,N_43910);
nand U44086 (N_44086,N_43895,N_43670);
and U44087 (N_44087,N_43912,N_43584);
or U44088 (N_44088,N_43839,N_43833);
xnor U44089 (N_44089,N_43625,N_43512);
nor U44090 (N_44090,N_43818,N_43561);
nor U44091 (N_44091,N_43585,N_43981);
nand U44092 (N_44092,N_43894,N_43916);
nor U44093 (N_44093,N_43602,N_43594);
and U44094 (N_44094,N_43754,N_43581);
xor U44095 (N_44095,N_43722,N_43809);
nor U44096 (N_44096,N_43876,N_43746);
xor U44097 (N_44097,N_43527,N_43521);
nor U44098 (N_44098,N_43791,N_43995);
or U44099 (N_44099,N_43924,N_43923);
or U44100 (N_44100,N_43753,N_43687);
nor U44101 (N_44101,N_43555,N_43678);
nor U44102 (N_44102,N_43568,N_43675);
and U44103 (N_44103,N_43963,N_43985);
nor U44104 (N_44104,N_43867,N_43542);
xor U44105 (N_44105,N_43801,N_43616);
or U44106 (N_44106,N_43776,N_43820);
or U44107 (N_44107,N_43744,N_43762);
nand U44108 (N_44108,N_43938,N_43939);
and U44109 (N_44109,N_43897,N_43676);
xor U44110 (N_44110,N_43841,N_43827);
nor U44111 (N_44111,N_43864,N_43700);
xor U44112 (N_44112,N_43590,N_43953);
or U44113 (N_44113,N_43743,N_43578);
xor U44114 (N_44114,N_43607,N_43794);
xnor U44115 (N_44115,N_43860,N_43816);
or U44116 (N_44116,N_43935,N_43899);
xor U44117 (N_44117,N_43826,N_43515);
or U44118 (N_44118,N_43666,N_43651);
nand U44119 (N_44119,N_43965,N_43819);
nor U44120 (N_44120,N_43803,N_43878);
or U44121 (N_44121,N_43618,N_43795);
or U44122 (N_44122,N_43611,N_43949);
and U44123 (N_44123,N_43608,N_43842);
nor U44124 (N_44124,N_43915,N_43750);
nor U44125 (N_44125,N_43524,N_43988);
nand U44126 (N_44126,N_43857,N_43526);
nand U44127 (N_44127,N_43634,N_43974);
and U44128 (N_44128,N_43908,N_43805);
and U44129 (N_44129,N_43834,N_43991);
and U44130 (N_44130,N_43672,N_43681);
or U44131 (N_44131,N_43548,N_43697);
or U44132 (N_44132,N_43821,N_43640);
or U44133 (N_44133,N_43798,N_43806);
nand U44134 (N_44134,N_43539,N_43789);
nor U44135 (N_44135,N_43814,N_43843);
or U44136 (N_44136,N_43919,N_43677);
nor U44137 (N_44137,N_43647,N_43797);
or U44138 (N_44138,N_43936,N_43922);
and U44139 (N_44139,N_43708,N_43612);
nor U44140 (N_44140,N_43861,N_43771);
and U44141 (N_44141,N_43639,N_43760);
xor U44142 (N_44142,N_43869,N_43747);
or U44143 (N_44143,N_43846,N_43707);
nor U44144 (N_44144,N_43714,N_43709);
and U44145 (N_44145,N_43977,N_43533);
and U44146 (N_44146,N_43906,N_43937);
nand U44147 (N_44147,N_43688,N_43657);
or U44148 (N_44148,N_43720,N_43537);
nor U44149 (N_44149,N_43976,N_43560);
nor U44150 (N_44150,N_43575,N_43946);
or U44151 (N_44151,N_43983,N_43845);
or U44152 (N_44152,N_43849,N_43740);
xor U44153 (N_44153,N_43928,N_43883);
xnor U44154 (N_44154,N_43552,N_43516);
or U44155 (N_44155,N_43699,N_43669);
nor U44156 (N_44156,N_43613,N_43693);
or U44157 (N_44157,N_43808,N_43556);
nor U44158 (N_44158,N_43784,N_43649);
xor U44159 (N_44159,N_43952,N_43629);
xnor U44160 (N_44160,N_43884,N_43898);
or U44161 (N_44161,N_43733,N_43994);
nor U44162 (N_44162,N_43692,N_43724);
and U44163 (N_44163,N_43701,N_43815);
nand U44164 (N_44164,N_43862,N_43505);
xor U44165 (N_44165,N_43975,N_43731);
or U44166 (N_44166,N_43850,N_43925);
or U44167 (N_44167,N_43926,N_43917);
xnor U44168 (N_44168,N_43941,N_43591);
nor U44169 (N_44169,N_43682,N_43644);
xor U44170 (N_44170,N_43538,N_43696);
or U44171 (N_44171,N_43739,N_43661);
nand U44172 (N_44172,N_43705,N_43943);
nand U44173 (N_44173,N_43788,N_43503);
nand U44174 (N_44174,N_43721,N_43875);
xnor U44175 (N_44175,N_43858,N_43617);
or U44176 (N_44176,N_43627,N_43566);
nor U44177 (N_44177,N_43960,N_43852);
nor U44178 (N_44178,N_43650,N_43544);
nand U44179 (N_44179,N_43643,N_43948);
nor U44180 (N_44180,N_43735,N_43614);
or U44181 (N_44181,N_43970,N_43529);
xnor U44182 (N_44182,N_43911,N_43824);
xor U44183 (N_44183,N_43811,N_43961);
nand U44184 (N_44184,N_43947,N_43596);
xnor U44185 (N_44185,N_43848,N_43686);
xnor U44186 (N_44186,N_43881,N_43921);
or U44187 (N_44187,N_43593,N_43969);
or U44188 (N_44188,N_43734,N_43635);
xor U44189 (N_44189,N_43671,N_43583);
nor U44190 (N_44190,N_43655,N_43703);
nor U44191 (N_44191,N_43835,N_43967);
or U44192 (N_44192,N_43638,N_43736);
nand U44193 (N_44193,N_43641,N_43766);
nor U44194 (N_44194,N_43802,N_43786);
or U44195 (N_44195,N_43885,N_43615);
nor U44196 (N_44196,N_43959,N_43610);
and U44197 (N_44197,N_43980,N_43879);
or U44198 (N_44198,N_43631,N_43759);
and U44199 (N_44199,N_43871,N_43569);
and U44200 (N_44200,N_43506,N_43501);
nand U44201 (N_44201,N_43918,N_43950);
nand U44202 (N_44202,N_43567,N_43896);
xor U44203 (N_44203,N_43893,N_43558);
nor U44204 (N_44204,N_43710,N_43565);
and U44205 (N_44205,N_43626,N_43509);
or U44206 (N_44206,N_43563,N_43997);
or U44207 (N_44207,N_43942,N_43880);
nand U44208 (N_44208,N_43972,N_43549);
nand U44209 (N_44209,N_43690,N_43996);
nor U44210 (N_44210,N_43554,N_43775);
xor U44211 (N_44211,N_43847,N_43765);
and U44212 (N_44212,N_43956,N_43684);
xnor U44213 (N_44213,N_43653,N_43907);
nor U44214 (N_44214,N_43825,N_43582);
nor U44215 (N_44215,N_43624,N_43535);
xor U44216 (N_44216,N_43717,N_43855);
and U44217 (N_44217,N_43992,N_43511);
nor U44218 (N_44218,N_43892,N_43913);
nand U44219 (N_44219,N_43990,N_43605);
nand U44220 (N_44220,N_43853,N_43652);
xnor U44221 (N_44221,N_43800,N_43725);
xnor U44222 (N_44222,N_43774,N_43507);
nor U44223 (N_44223,N_43830,N_43570);
nand U44224 (N_44224,N_43531,N_43955);
and U44225 (N_44225,N_43728,N_43773);
xnor U44226 (N_44226,N_43719,N_43648);
nor U44227 (N_44227,N_43782,N_43598);
and U44228 (N_44228,N_43829,N_43989);
and U44229 (N_44229,N_43522,N_43557);
or U44230 (N_44230,N_43547,N_43905);
nand U44231 (N_44231,N_43597,N_43822);
nand U44232 (N_44232,N_43663,N_43968);
xor U44233 (N_44233,N_43586,N_43752);
nand U44234 (N_44234,N_43828,N_43543);
and U44235 (N_44235,N_43559,N_43718);
or U44236 (N_44236,N_43619,N_43673);
nor U44237 (N_44237,N_43920,N_43680);
or U44238 (N_44238,N_43904,N_43604);
nor U44239 (N_44239,N_43637,N_43698);
xor U44240 (N_44240,N_43665,N_43966);
nor U44241 (N_44241,N_43865,N_43659);
xor U44242 (N_44242,N_43971,N_43796);
xor U44243 (N_44243,N_43767,N_43930);
nor U44244 (N_44244,N_43600,N_43993);
xnor U44245 (N_44245,N_43978,N_43609);
and U44246 (N_44246,N_43689,N_43951);
xor U44247 (N_44247,N_43500,N_43711);
and U44248 (N_44248,N_43520,N_43660);
and U44249 (N_44249,N_43851,N_43783);
and U44250 (N_44250,N_43610,N_43941);
and U44251 (N_44251,N_43501,N_43751);
or U44252 (N_44252,N_43532,N_43769);
or U44253 (N_44253,N_43920,N_43508);
or U44254 (N_44254,N_43809,N_43623);
nand U44255 (N_44255,N_43942,N_43720);
and U44256 (N_44256,N_43677,N_43988);
and U44257 (N_44257,N_43861,N_43908);
and U44258 (N_44258,N_43740,N_43576);
nand U44259 (N_44259,N_43710,N_43991);
and U44260 (N_44260,N_43528,N_43947);
or U44261 (N_44261,N_43848,N_43520);
xor U44262 (N_44262,N_43592,N_43889);
xor U44263 (N_44263,N_43771,N_43993);
and U44264 (N_44264,N_43604,N_43907);
nand U44265 (N_44265,N_43726,N_43512);
nor U44266 (N_44266,N_43636,N_43856);
nor U44267 (N_44267,N_43754,N_43719);
and U44268 (N_44268,N_43751,N_43800);
xor U44269 (N_44269,N_43738,N_43716);
xnor U44270 (N_44270,N_43684,N_43747);
and U44271 (N_44271,N_43617,N_43825);
nand U44272 (N_44272,N_43987,N_43858);
or U44273 (N_44273,N_43653,N_43668);
nand U44274 (N_44274,N_43935,N_43730);
or U44275 (N_44275,N_43664,N_43575);
nand U44276 (N_44276,N_43939,N_43620);
xnor U44277 (N_44277,N_43730,N_43840);
nand U44278 (N_44278,N_43549,N_43867);
and U44279 (N_44279,N_43571,N_43961);
nand U44280 (N_44280,N_43657,N_43668);
nand U44281 (N_44281,N_43618,N_43889);
and U44282 (N_44282,N_43990,N_43877);
or U44283 (N_44283,N_43873,N_43855);
and U44284 (N_44284,N_43816,N_43739);
xnor U44285 (N_44285,N_43523,N_43721);
nand U44286 (N_44286,N_43531,N_43729);
or U44287 (N_44287,N_43502,N_43583);
nand U44288 (N_44288,N_43917,N_43595);
nor U44289 (N_44289,N_43683,N_43718);
nor U44290 (N_44290,N_43680,N_43612);
or U44291 (N_44291,N_43910,N_43630);
nand U44292 (N_44292,N_43686,N_43824);
nor U44293 (N_44293,N_43699,N_43546);
nand U44294 (N_44294,N_43533,N_43973);
nand U44295 (N_44295,N_43653,N_43981);
xnor U44296 (N_44296,N_43981,N_43723);
nand U44297 (N_44297,N_43591,N_43912);
or U44298 (N_44298,N_43840,N_43849);
or U44299 (N_44299,N_43916,N_43653);
xnor U44300 (N_44300,N_43839,N_43756);
or U44301 (N_44301,N_43779,N_43919);
nor U44302 (N_44302,N_43790,N_43729);
xor U44303 (N_44303,N_43601,N_43643);
and U44304 (N_44304,N_43666,N_43935);
nor U44305 (N_44305,N_43761,N_43620);
and U44306 (N_44306,N_43572,N_43734);
xnor U44307 (N_44307,N_43696,N_43933);
nor U44308 (N_44308,N_43750,N_43560);
xor U44309 (N_44309,N_43863,N_43976);
xnor U44310 (N_44310,N_43651,N_43770);
or U44311 (N_44311,N_43710,N_43916);
nand U44312 (N_44312,N_43868,N_43743);
and U44313 (N_44313,N_43770,N_43690);
nor U44314 (N_44314,N_43571,N_43670);
nor U44315 (N_44315,N_43739,N_43872);
xor U44316 (N_44316,N_43573,N_43847);
nand U44317 (N_44317,N_43786,N_43992);
nor U44318 (N_44318,N_43502,N_43688);
nor U44319 (N_44319,N_43843,N_43667);
or U44320 (N_44320,N_43869,N_43675);
and U44321 (N_44321,N_43740,N_43540);
and U44322 (N_44322,N_43697,N_43751);
and U44323 (N_44323,N_43539,N_43945);
xnor U44324 (N_44324,N_43812,N_43612);
nor U44325 (N_44325,N_43740,N_43636);
or U44326 (N_44326,N_43800,N_43776);
nor U44327 (N_44327,N_43948,N_43796);
nor U44328 (N_44328,N_43642,N_43547);
nand U44329 (N_44329,N_43709,N_43746);
and U44330 (N_44330,N_43644,N_43876);
and U44331 (N_44331,N_43700,N_43880);
and U44332 (N_44332,N_43747,N_43983);
and U44333 (N_44333,N_43816,N_43878);
nor U44334 (N_44334,N_43928,N_43774);
nand U44335 (N_44335,N_43639,N_43989);
nand U44336 (N_44336,N_43516,N_43959);
nor U44337 (N_44337,N_43760,N_43567);
nand U44338 (N_44338,N_43528,N_43920);
nand U44339 (N_44339,N_43954,N_43856);
or U44340 (N_44340,N_43750,N_43625);
and U44341 (N_44341,N_43569,N_43729);
and U44342 (N_44342,N_43780,N_43604);
and U44343 (N_44343,N_43900,N_43985);
nand U44344 (N_44344,N_43618,N_43894);
nor U44345 (N_44345,N_43613,N_43548);
nand U44346 (N_44346,N_43706,N_43564);
nor U44347 (N_44347,N_43547,N_43561);
xor U44348 (N_44348,N_43623,N_43650);
and U44349 (N_44349,N_43676,N_43893);
or U44350 (N_44350,N_43793,N_43689);
nor U44351 (N_44351,N_43870,N_43947);
nand U44352 (N_44352,N_43939,N_43649);
or U44353 (N_44353,N_43822,N_43914);
nand U44354 (N_44354,N_43762,N_43786);
xnor U44355 (N_44355,N_43705,N_43596);
xnor U44356 (N_44356,N_43848,N_43992);
nor U44357 (N_44357,N_43826,N_43825);
xor U44358 (N_44358,N_43510,N_43886);
or U44359 (N_44359,N_43503,N_43598);
nand U44360 (N_44360,N_43736,N_43667);
nor U44361 (N_44361,N_43970,N_43772);
and U44362 (N_44362,N_43900,N_43858);
and U44363 (N_44363,N_43832,N_43691);
nor U44364 (N_44364,N_43870,N_43943);
or U44365 (N_44365,N_43700,N_43633);
or U44366 (N_44366,N_43975,N_43506);
nor U44367 (N_44367,N_43720,N_43619);
and U44368 (N_44368,N_43520,N_43662);
nand U44369 (N_44369,N_43640,N_43592);
and U44370 (N_44370,N_43894,N_43973);
xnor U44371 (N_44371,N_43728,N_43877);
or U44372 (N_44372,N_43539,N_43603);
nor U44373 (N_44373,N_43594,N_43995);
or U44374 (N_44374,N_43525,N_43684);
xor U44375 (N_44375,N_43719,N_43502);
or U44376 (N_44376,N_43661,N_43986);
or U44377 (N_44377,N_43798,N_43843);
or U44378 (N_44378,N_43708,N_43853);
xnor U44379 (N_44379,N_43518,N_43560);
nand U44380 (N_44380,N_43798,N_43713);
or U44381 (N_44381,N_43617,N_43932);
nand U44382 (N_44382,N_43526,N_43516);
nand U44383 (N_44383,N_43674,N_43999);
or U44384 (N_44384,N_43846,N_43885);
xnor U44385 (N_44385,N_43569,N_43986);
and U44386 (N_44386,N_43513,N_43726);
and U44387 (N_44387,N_43888,N_43757);
or U44388 (N_44388,N_43882,N_43696);
or U44389 (N_44389,N_43911,N_43596);
nor U44390 (N_44390,N_43560,N_43814);
and U44391 (N_44391,N_43573,N_43639);
nor U44392 (N_44392,N_43986,N_43779);
nor U44393 (N_44393,N_43628,N_43644);
and U44394 (N_44394,N_43773,N_43849);
and U44395 (N_44395,N_43513,N_43652);
nand U44396 (N_44396,N_43866,N_43886);
or U44397 (N_44397,N_43778,N_43885);
and U44398 (N_44398,N_43920,N_43823);
nand U44399 (N_44399,N_43879,N_43808);
nand U44400 (N_44400,N_43835,N_43830);
nand U44401 (N_44401,N_43516,N_43846);
xor U44402 (N_44402,N_43725,N_43924);
xnor U44403 (N_44403,N_43881,N_43886);
and U44404 (N_44404,N_43834,N_43791);
nand U44405 (N_44405,N_43782,N_43545);
or U44406 (N_44406,N_43847,N_43923);
nor U44407 (N_44407,N_43674,N_43933);
nor U44408 (N_44408,N_43643,N_43851);
or U44409 (N_44409,N_43989,N_43873);
xor U44410 (N_44410,N_43682,N_43900);
nand U44411 (N_44411,N_43683,N_43673);
or U44412 (N_44412,N_43514,N_43717);
nand U44413 (N_44413,N_43863,N_43813);
or U44414 (N_44414,N_43966,N_43915);
and U44415 (N_44415,N_43673,N_43952);
xnor U44416 (N_44416,N_43980,N_43777);
nand U44417 (N_44417,N_43764,N_43656);
or U44418 (N_44418,N_43982,N_43570);
or U44419 (N_44419,N_43918,N_43831);
xnor U44420 (N_44420,N_43654,N_43773);
nor U44421 (N_44421,N_43855,N_43621);
and U44422 (N_44422,N_43916,N_43676);
and U44423 (N_44423,N_43698,N_43973);
nor U44424 (N_44424,N_43921,N_43552);
or U44425 (N_44425,N_43800,N_43968);
xor U44426 (N_44426,N_43687,N_43871);
or U44427 (N_44427,N_43703,N_43558);
nor U44428 (N_44428,N_43759,N_43929);
xor U44429 (N_44429,N_43517,N_43620);
nor U44430 (N_44430,N_43654,N_43795);
xor U44431 (N_44431,N_43623,N_43575);
nor U44432 (N_44432,N_43998,N_43912);
or U44433 (N_44433,N_43681,N_43919);
and U44434 (N_44434,N_43588,N_43723);
and U44435 (N_44435,N_43715,N_43902);
xnor U44436 (N_44436,N_43984,N_43739);
or U44437 (N_44437,N_43733,N_43875);
nor U44438 (N_44438,N_43989,N_43512);
nand U44439 (N_44439,N_43811,N_43584);
nand U44440 (N_44440,N_43619,N_43524);
xor U44441 (N_44441,N_43876,N_43735);
and U44442 (N_44442,N_43659,N_43617);
nor U44443 (N_44443,N_43871,N_43890);
xor U44444 (N_44444,N_43875,N_43882);
and U44445 (N_44445,N_43840,N_43764);
nor U44446 (N_44446,N_43685,N_43575);
xnor U44447 (N_44447,N_43540,N_43701);
nand U44448 (N_44448,N_43809,N_43837);
or U44449 (N_44449,N_43877,N_43985);
xnor U44450 (N_44450,N_43712,N_43699);
nor U44451 (N_44451,N_43792,N_43975);
nor U44452 (N_44452,N_43503,N_43526);
xnor U44453 (N_44453,N_43668,N_43539);
and U44454 (N_44454,N_43942,N_43579);
nand U44455 (N_44455,N_43861,N_43787);
xnor U44456 (N_44456,N_43585,N_43685);
or U44457 (N_44457,N_43760,N_43915);
xnor U44458 (N_44458,N_43652,N_43786);
nor U44459 (N_44459,N_43886,N_43641);
or U44460 (N_44460,N_43618,N_43670);
nand U44461 (N_44461,N_43979,N_43908);
nand U44462 (N_44462,N_43823,N_43597);
or U44463 (N_44463,N_43681,N_43935);
nand U44464 (N_44464,N_43903,N_43822);
nand U44465 (N_44465,N_43971,N_43919);
nor U44466 (N_44466,N_43667,N_43900);
and U44467 (N_44467,N_43717,N_43527);
xor U44468 (N_44468,N_43824,N_43576);
xor U44469 (N_44469,N_43512,N_43862);
xnor U44470 (N_44470,N_43901,N_43511);
and U44471 (N_44471,N_43614,N_43935);
or U44472 (N_44472,N_43773,N_43946);
or U44473 (N_44473,N_43631,N_43945);
or U44474 (N_44474,N_43718,N_43658);
and U44475 (N_44475,N_43504,N_43883);
and U44476 (N_44476,N_43642,N_43776);
xnor U44477 (N_44477,N_43732,N_43994);
and U44478 (N_44478,N_43707,N_43918);
xnor U44479 (N_44479,N_43621,N_43566);
xor U44480 (N_44480,N_43897,N_43609);
or U44481 (N_44481,N_43658,N_43695);
or U44482 (N_44482,N_43961,N_43555);
nand U44483 (N_44483,N_43782,N_43503);
or U44484 (N_44484,N_43536,N_43818);
nand U44485 (N_44485,N_43737,N_43723);
nor U44486 (N_44486,N_43845,N_43813);
nand U44487 (N_44487,N_43551,N_43575);
or U44488 (N_44488,N_43825,N_43683);
and U44489 (N_44489,N_43943,N_43930);
nand U44490 (N_44490,N_43896,N_43770);
nand U44491 (N_44491,N_43849,N_43505);
and U44492 (N_44492,N_43651,N_43622);
and U44493 (N_44493,N_43684,N_43963);
or U44494 (N_44494,N_43849,N_43823);
nor U44495 (N_44495,N_43550,N_43861);
nand U44496 (N_44496,N_43623,N_43715);
or U44497 (N_44497,N_43708,N_43553);
or U44498 (N_44498,N_43763,N_43607);
xor U44499 (N_44499,N_43573,N_43533);
nor U44500 (N_44500,N_44337,N_44249);
or U44501 (N_44501,N_44365,N_44098);
nand U44502 (N_44502,N_44226,N_44280);
xnor U44503 (N_44503,N_44107,N_44278);
and U44504 (N_44504,N_44385,N_44379);
or U44505 (N_44505,N_44061,N_44206);
nor U44506 (N_44506,N_44053,N_44037);
nor U44507 (N_44507,N_44482,N_44316);
nand U44508 (N_44508,N_44080,N_44058);
nand U44509 (N_44509,N_44052,N_44245);
or U44510 (N_44510,N_44306,N_44148);
nor U44511 (N_44511,N_44464,N_44471);
nor U44512 (N_44512,N_44346,N_44156);
or U44513 (N_44513,N_44152,N_44212);
or U44514 (N_44514,N_44041,N_44421);
and U44515 (N_44515,N_44048,N_44275);
or U44516 (N_44516,N_44017,N_44162);
nor U44517 (N_44517,N_44133,N_44386);
nand U44518 (N_44518,N_44493,N_44217);
nand U44519 (N_44519,N_44260,N_44085);
or U44520 (N_44520,N_44091,N_44353);
xor U44521 (N_44521,N_44042,N_44220);
nor U44522 (N_44522,N_44197,N_44189);
nand U44523 (N_44523,N_44426,N_44372);
nand U44524 (N_44524,N_44185,N_44022);
nor U44525 (N_44525,N_44020,N_44031);
and U44526 (N_44526,N_44259,N_44413);
and U44527 (N_44527,N_44466,N_44113);
xor U44528 (N_44528,N_44474,N_44446);
and U44529 (N_44529,N_44099,N_44011);
and U44530 (N_44530,N_44263,N_44066);
or U44531 (N_44531,N_44139,N_44300);
nand U44532 (N_44532,N_44265,N_44062);
or U44533 (N_44533,N_44431,N_44382);
nand U44534 (N_44534,N_44253,N_44005);
nand U44535 (N_44535,N_44293,N_44318);
xor U44536 (N_44536,N_44046,N_44384);
nor U44537 (N_44537,N_44458,N_44092);
nand U44538 (N_44538,N_44402,N_44355);
or U44539 (N_44539,N_44331,N_44486);
or U44540 (N_44540,N_44014,N_44160);
and U44541 (N_44541,N_44344,N_44254);
and U44542 (N_44542,N_44064,N_44301);
nor U44543 (N_44543,N_44257,N_44078);
nor U44544 (N_44544,N_44494,N_44242);
nor U44545 (N_44545,N_44439,N_44045);
and U44546 (N_44546,N_44327,N_44227);
nand U44547 (N_44547,N_44174,N_44171);
or U44548 (N_44548,N_44200,N_44103);
nand U44549 (N_44549,N_44068,N_44490);
nand U44550 (N_44550,N_44038,N_44118);
or U44551 (N_44551,N_44456,N_44338);
nor U44552 (N_44552,N_44207,N_44349);
xnor U44553 (N_44553,N_44213,N_44360);
xor U44554 (N_44554,N_44291,N_44304);
xnor U44555 (N_44555,N_44181,N_44416);
nand U44556 (N_44556,N_44295,N_44427);
xor U44557 (N_44557,N_44154,N_44069);
nor U44558 (N_44558,N_44376,N_44480);
nor U44559 (N_44559,N_44012,N_44381);
and U44560 (N_44560,N_44237,N_44288);
nand U44561 (N_44561,N_44325,N_44004);
nand U44562 (N_44562,N_44309,N_44423);
or U44563 (N_44563,N_44333,N_44282);
and U44564 (N_44564,N_44027,N_44043);
nor U44565 (N_44565,N_44371,N_44025);
nand U44566 (N_44566,N_44202,N_44044);
nand U44567 (N_44567,N_44463,N_44015);
nor U44568 (N_44568,N_44120,N_44175);
nor U44569 (N_44569,N_44100,N_44215);
nand U44570 (N_44570,N_44125,N_44452);
nor U44571 (N_44571,N_44460,N_44039);
and U44572 (N_44572,N_44296,N_44223);
nor U44573 (N_44573,N_44326,N_44169);
or U44574 (N_44574,N_44201,N_44425);
or U44575 (N_44575,N_44158,N_44131);
nor U44576 (N_44576,N_44082,N_44430);
or U44577 (N_44577,N_44285,N_44214);
nor U44578 (N_44578,N_44434,N_44164);
xnor U44579 (N_44579,N_44467,N_44136);
and U44580 (N_44580,N_44095,N_44356);
xnor U44581 (N_44581,N_44147,N_44188);
nor U44582 (N_44582,N_44040,N_44117);
nor U44583 (N_44583,N_44369,N_44496);
nand U44584 (N_44584,N_44418,N_44252);
xor U44585 (N_44585,N_44395,N_44483);
nor U44586 (N_44586,N_44266,N_44334);
or U44587 (N_44587,N_44396,N_44187);
nor U44588 (N_44588,N_44122,N_44047);
xnor U44589 (N_44589,N_44248,N_44086);
xor U44590 (N_44590,N_44150,N_44083);
or U44591 (N_44591,N_44216,N_44328);
and U44592 (N_44592,N_44271,N_44420);
and U44593 (N_44593,N_44432,N_44303);
xnor U44594 (N_44594,N_44143,N_44350);
nand U44595 (N_44595,N_44116,N_44283);
nor U44596 (N_44596,N_44030,N_44246);
xnor U44597 (N_44597,N_44443,N_44424);
nand U44598 (N_44598,N_44023,N_44234);
nor U44599 (N_44599,N_44233,N_44361);
or U44600 (N_44600,N_44305,N_44221);
nor U44601 (N_44601,N_44009,N_44407);
or U44602 (N_44602,N_44137,N_44232);
xnor U44603 (N_44603,N_44499,N_44114);
xnor U44604 (N_44604,N_44429,N_44236);
nor U44605 (N_44605,N_44315,N_44459);
nand U44606 (N_44606,N_44157,N_44054);
xnor U44607 (N_44607,N_44021,N_44184);
nand U44608 (N_44608,N_44389,N_44241);
and U44609 (N_44609,N_44281,N_44461);
nand U44610 (N_44610,N_44194,N_44388);
nand U44611 (N_44611,N_44279,N_44130);
nand U44612 (N_44612,N_44149,N_44308);
or U44613 (N_44613,N_44168,N_44495);
nand U44614 (N_44614,N_44475,N_44341);
xnor U44615 (N_44615,N_44076,N_44205);
nand U44616 (N_44616,N_44127,N_44404);
nand U44617 (N_44617,N_44172,N_44230);
or U44618 (N_44618,N_44394,N_44177);
nand U44619 (N_44619,N_44477,N_44112);
nand U44620 (N_44620,N_44159,N_44209);
or U44621 (N_44621,N_44391,N_44075);
or U44622 (N_44622,N_44240,N_44183);
nand U44623 (N_44623,N_44138,N_44312);
or U44624 (N_44624,N_44251,N_44294);
nand U44625 (N_44625,N_44492,N_44128);
nor U44626 (N_44626,N_44343,N_44287);
xor U44627 (N_44627,N_44319,N_44250);
nand U44628 (N_44628,N_44104,N_44008);
nand U44629 (N_44629,N_44050,N_44405);
nor U44630 (N_44630,N_44310,N_44060);
xor U44631 (N_44631,N_44269,N_44146);
xnor U44632 (N_44632,N_44419,N_44247);
or U44633 (N_44633,N_44203,N_44115);
nand U44634 (N_44634,N_44070,N_44123);
or U44635 (N_44635,N_44051,N_44244);
nand U44636 (N_44636,N_44406,N_44028);
and U44637 (N_44637,N_44298,N_44093);
xnor U44638 (N_44638,N_44445,N_44457);
nor U44639 (N_44639,N_44163,N_44497);
xor U44640 (N_44640,N_44176,N_44373);
or U44641 (N_44641,N_44032,N_44358);
nor U44642 (N_44642,N_44166,N_44448);
xor U44643 (N_44643,N_44270,N_44442);
xor U44644 (N_44644,N_44342,N_44010);
xor U44645 (N_44645,N_44357,N_44330);
xnor U44646 (N_44646,N_44073,N_44397);
or U44647 (N_44647,N_44468,N_44314);
nand U44648 (N_44648,N_44449,N_44084);
or U44649 (N_44649,N_44210,N_44436);
and U44650 (N_44650,N_44109,N_44204);
nor U44651 (N_44651,N_44057,N_44108);
nor U44652 (N_44652,N_44335,N_44016);
and U44653 (N_44653,N_44299,N_44392);
or U44654 (N_44654,N_44491,N_44261);
nor U44655 (N_44655,N_44322,N_44380);
and U44656 (N_44656,N_44339,N_44074);
nor U44657 (N_44657,N_44367,N_44336);
and U44658 (N_44658,N_44498,N_44178);
xnor U44659 (N_44659,N_44255,N_44155);
xor U44660 (N_44660,N_44311,N_44262);
xor U44661 (N_44661,N_44412,N_44489);
xnor U44662 (N_44662,N_44323,N_44135);
xnor U44663 (N_44663,N_44121,N_44428);
or U44664 (N_44664,N_44354,N_44231);
xnor U44665 (N_44665,N_44003,N_44228);
nor U44666 (N_44666,N_44090,N_44191);
nand U44667 (N_44667,N_44472,N_44444);
nand U44668 (N_44668,N_44351,N_44173);
xnor U44669 (N_44669,N_44000,N_44476);
nor U44670 (N_44670,N_44447,N_44218);
xnor U44671 (N_44671,N_44065,N_44151);
nand U44672 (N_44672,N_44347,N_44059);
and U44673 (N_44673,N_44340,N_44071);
or U44674 (N_44674,N_44454,N_44018);
and U44675 (N_44675,N_44313,N_44393);
xor U44676 (N_44676,N_44195,N_44320);
nor U44677 (N_44677,N_44414,N_44473);
or U44678 (N_44678,N_44140,N_44063);
nand U44679 (N_44679,N_44094,N_44119);
xnor U44680 (N_44680,N_44019,N_44208);
xor U44681 (N_44681,N_44433,N_44081);
nand U44682 (N_44682,N_44134,N_44190);
nand U44683 (N_44683,N_44167,N_44199);
or U44684 (N_44684,N_44161,N_44106);
or U44685 (N_44685,N_44363,N_44451);
and U44686 (N_44686,N_44276,N_44036);
and U44687 (N_44687,N_44193,N_44101);
or U44688 (N_44688,N_44441,N_44111);
and U44689 (N_44689,N_44219,N_44096);
nor U44690 (N_44690,N_44097,N_44180);
nor U44691 (N_44691,N_44274,N_44435);
and U44692 (N_44692,N_44007,N_44034);
and U44693 (N_44693,N_44469,N_44165);
nand U44694 (N_44694,N_44006,N_44470);
xor U44695 (N_44695,N_44235,N_44079);
nor U44696 (N_44696,N_44198,N_44364);
or U44697 (N_44697,N_44284,N_44465);
xnor U44698 (N_44698,N_44307,N_44345);
or U44699 (N_44699,N_44399,N_44484);
xor U44700 (N_44700,N_44029,N_44398);
or U44701 (N_44701,N_44362,N_44411);
or U44702 (N_44702,N_44238,N_44359);
xor U44703 (N_44703,N_44400,N_44132);
nor U44704 (N_44704,N_44481,N_44087);
nand U44705 (N_44705,N_44348,N_44289);
and U44706 (N_44706,N_44478,N_44222);
nor U44707 (N_44707,N_44056,N_44403);
xnor U44708 (N_44708,N_44273,N_44239);
xnor U44709 (N_44709,N_44378,N_44462);
and U44710 (N_44710,N_44033,N_44024);
nor U44711 (N_44711,N_44290,N_44264);
nor U44712 (N_44712,N_44182,N_44243);
nand U44713 (N_44713,N_44002,N_44479);
nand U44714 (N_44714,N_44352,N_44089);
nor U44715 (N_44715,N_44292,N_44297);
nand U44716 (N_44716,N_44153,N_44437);
or U44717 (N_44717,N_44453,N_44409);
nand U44718 (N_44718,N_44317,N_44390);
nand U44719 (N_44719,N_44026,N_44408);
or U44720 (N_44720,N_44410,N_44440);
or U44721 (N_44721,N_44170,N_44383);
nand U44722 (N_44722,N_44110,N_44258);
and U44723 (N_44723,N_44401,N_44387);
and U44724 (N_44724,N_44067,N_44277);
nand U44725 (N_44725,N_44450,N_44001);
and U44726 (N_44726,N_44225,N_44267);
nor U44727 (N_44727,N_44329,N_44105);
nand U44728 (N_44728,N_44229,N_44144);
xor U44729 (N_44729,N_44302,N_44088);
xor U44730 (N_44730,N_44417,N_44332);
nand U44731 (N_44731,N_44377,N_44422);
or U44732 (N_44732,N_44374,N_44455);
or U44733 (N_44733,N_44077,N_44488);
nand U44734 (N_44734,N_44256,N_44370);
nor U44735 (N_44735,N_44013,N_44272);
nor U44736 (N_44736,N_44286,N_44485);
xnor U44737 (N_44737,N_44129,N_44196);
or U44738 (N_44738,N_44268,N_44035);
and U44739 (N_44739,N_44072,N_44211);
xnor U44740 (N_44740,N_44366,N_44438);
nor U44741 (N_44741,N_44415,N_44324);
and U44742 (N_44742,N_44192,N_44102);
nor U44743 (N_44743,N_44141,N_44186);
and U44744 (N_44744,N_44126,N_44375);
xor U44745 (N_44745,N_44368,N_44321);
nor U44746 (N_44746,N_44055,N_44049);
or U44747 (N_44747,N_44487,N_44224);
nor U44748 (N_44748,N_44145,N_44124);
xor U44749 (N_44749,N_44179,N_44142);
xor U44750 (N_44750,N_44404,N_44419);
nand U44751 (N_44751,N_44065,N_44154);
nand U44752 (N_44752,N_44215,N_44312);
or U44753 (N_44753,N_44414,N_44111);
xor U44754 (N_44754,N_44104,N_44235);
nor U44755 (N_44755,N_44273,N_44201);
or U44756 (N_44756,N_44024,N_44282);
and U44757 (N_44757,N_44378,N_44474);
nor U44758 (N_44758,N_44270,N_44175);
nor U44759 (N_44759,N_44196,N_44279);
and U44760 (N_44760,N_44123,N_44168);
nor U44761 (N_44761,N_44304,N_44363);
nor U44762 (N_44762,N_44360,N_44203);
nor U44763 (N_44763,N_44497,N_44275);
nand U44764 (N_44764,N_44270,N_44259);
or U44765 (N_44765,N_44412,N_44382);
nor U44766 (N_44766,N_44066,N_44387);
nor U44767 (N_44767,N_44443,N_44318);
nand U44768 (N_44768,N_44244,N_44194);
and U44769 (N_44769,N_44404,N_44194);
xor U44770 (N_44770,N_44106,N_44368);
nor U44771 (N_44771,N_44112,N_44115);
nor U44772 (N_44772,N_44044,N_44078);
nand U44773 (N_44773,N_44151,N_44296);
and U44774 (N_44774,N_44140,N_44252);
or U44775 (N_44775,N_44269,N_44469);
or U44776 (N_44776,N_44211,N_44249);
nor U44777 (N_44777,N_44074,N_44210);
nor U44778 (N_44778,N_44202,N_44470);
nand U44779 (N_44779,N_44011,N_44021);
or U44780 (N_44780,N_44454,N_44001);
xnor U44781 (N_44781,N_44297,N_44122);
nand U44782 (N_44782,N_44417,N_44151);
or U44783 (N_44783,N_44056,N_44396);
and U44784 (N_44784,N_44197,N_44272);
nand U44785 (N_44785,N_44475,N_44444);
nor U44786 (N_44786,N_44247,N_44167);
nand U44787 (N_44787,N_44344,N_44011);
and U44788 (N_44788,N_44406,N_44310);
nor U44789 (N_44789,N_44496,N_44126);
xnor U44790 (N_44790,N_44025,N_44289);
and U44791 (N_44791,N_44315,N_44464);
and U44792 (N_44792,N_44471,N_44194);
or U44793 (N_44793,N_44422,N_44484);
nand U44794 (N_44794,N_44346,N_44113);
nand U44795 (N_44795,N_44378,N_44026);
or U44796 (N_44796,N_44296,N_44154);
or U44797 (N_44797,N_44103,N_44028);
nor U44798 (N_44798,N_44085,N_44467);
nand U44799 (N_44799,N_44466,N_44151);
and U44800 (N_44800,N_44259,N_44351);
or U44801 (N_44801,N_44150,N_44002);
xnor U44802 (N_44802,N_44267,N_44026);
nor U44803 (N_44803,N_44219,N_44130);
or U44804 (N_44804,N_44405,N_44406);
xor U44805 (N_44805,N_44031,N_44479);
and U44806 (N_44806,N_44144,N_44294);
and U44807 (N_44807,N_44071,N_44450);
nor U44808 (N_44808,N_44056,N_44238);
or U44809 (N_44809,N_44241,N_44289);
xnor U44810 (N_44810,N_44013,N_44107);
nor U44811 (N_44811,N_44056,N_44180);
or U44812 (N_44812,N_44038,N_44287);
or U44813 (N_44813,N_44135,N_44280);
nor U44814 (N_44814,N_44106,N_44073);
or U44815 (N_44815,N_44485,N_44000);
and U44816 (N_44816,N_44106,N_44319);
nand U44817 (N_44817,N_44178,N_44200);
nand U44818 (N_44818,N_44008,N_44096);
and U44819 (N_44819,N_44250,N_44437);
and U44820 (N_44820,N_44336,N_44196);
and U44821 (N_44821,N_44141,N_44416);
xor U44822 (N_44822,N_44492,N_44273);
or U44823 (N_44823,N_44337,N_44457);
nand U44824 (N_44824,N_44489,N_44034);
or U44825 (N_44825,N_44335,N_44472);
nor U44826 (N_44826,N_44360,N_44034);
nor U44827 (N_44827,N_44245,N_44240);
xor U44828 (N_44828,N_44056,N_44485);
nand U44829 (N_44829,N_44362,N_44495);
and U44830 (N_44830,N_44301,N_44153);
nor U44831 (N_44831,N_44426,N_44024);
and U44832 (N_44832,N_44435,N_44010);
nand U44833 (N_44833,N_44246,N_44486);
or U44834 (N_44834,N_44094,N_44471);
and U44835 (N_44835,N_44008,N_44207);
and U44836 (N_44836,N_44083,N_44102);
or U44837 (N_44837,N_44225,N_44443);
xor U44838 (N_44838,N_44476,N_44475);
and U44839 (N_44839,N_44319,N_44025);
nand U44840 (N_44840,N_44065,N_44260);
and U44841 (N_44841,N_44400,N_44009);
xor U44842 (N_44842,N_44311,N_44025);
and U44843 (N_44843,N_44357,N_44106);
nor U44844 (N_44844,N_44361,N_44092);
and U44845 (N_44845,N_44224,N_44185);
nand U44846 (N_44846,N_44015,N_44322);
or U44847 (N_44847,N_44092,N_44295);
nor U44848 (N_44848,N_44028,N_44055);
and U44849 (N_44849,N_44174,N_44478);
nor U44850 (N_44850,N_44006,N_44393);
nand U44851 (N_44851,N_44449,N_44269);
xor U44852 (N_44852,N_44457,N_44091);
nand U44853 (N_44853,N_44201,N_44115);
xor U44854 (N_44854,N_44252,N_44435);
xor U44855 (N_44855,N_44279,N_44355);
or U44856 (N_44856,N_44289,N_44362);
nor U44857 (N_44857,N_44289,N_44173);
nor U44858 (N_44858,N_44050,N_44335);
xor U44859 (N_44859,N_44286,N_44279);
and U44860 (N_44860,N_44370,N_44109);
nor U44861 (N_44861,N_44224,N_44275);
and U44862 (N_44862,N_44408,N_44212);
nor U44863 (N_44863,N_44351,N_44156);
or U44864 (N_44864,N_44281,N_44478);
xor U44865 (N_44865,N_44227,N_44120);
and U44866 (N_44866,N_44316,N_44129);
nor U44867 (N_44867,N_44179,N_44460);
nor U44868 (N_44868,N_44287,N_44291);
and U44869 (N_44869,N_44265,N_44187);
or U44870 (N_44870,N_44081,N_44189);
nor U44871 (N_44871,N_44060,N_44340);
or U44872 (N_44872,N_44386,N_44128);
and U44873 (N_44873,N_44243,N_44455);
or U44874 (N_44874,N_44250,N_44290);
xnor U44875 (N_44875,N_44125,N_44402);
or U44876 (N_44876,N_44465,N_44061);
and U44877 (N_44877,N_44172,N_44311);
xor U44878 (N_44878,N_44286,N_44139);
or U44879 (N_44879,N_44469,N_44120);
xor U44880 (N_44880,N_44473,N_44211);
nand U44881 (N_44881,N_44357,N_44236);
or U44882 (N_44882,N_44025,N_44003);
or U44883 (N_44883,N_44293,N_44084);
or U44884 (N_44884,N_44358,N_44402);
and U44885 (N_44885,N_44183,N_44304);
or U44886 (N_44886,N_44478,N_44349);
and U44887 (N_44887,N_44266,N_44378);
and U44888 (N_44888,N_44009,N_44245);
nor U44889 (N_44889,N_44458,N_44036);
and U44890 (N_44890,N_44453,N_44031);
nand U44891 (N_44891,N_44334,N_44438);
nor U44892 (N_44892,N_44413,N_44085);
nor U44893 (N_44893,N_44020,N_44336);
or U44894 (N_44894,N_44464,N_44198);
nor U44895 (N_44895,N_44112,N_44113);
or U44896 (N_44896,N_44141,N_44443);
nand U44897 (N_44897,N_44152,N_44156);
xor U44898 (N_44898,N_44172,N_44063);
or U44899 (N_44899,N_44044,N_44395);
nor U44900 (N_44900,N_44263,N_44178);
nor U44901 (N_44901,N_44061,N_44113);
or U44902 (N_44902,N_44092,N_44056);
and U44903 (N_44903,N_44405,N_44350);
and U44904 (N_44904,N_44106,N_44030);
or U44905 (N_44905,N_44249,N_44339);
nand U44906 (N_44906,N_44087,N_44312);
xor U44907 (N_44907,N_44466,N_44031);
or U44908 (N_44908,N_44350,N_44339);
nor U44909 (N_44909,N_44282,N_44231);
or U44910 (N_44910,N_44367,N_44386);
and U44911 (N_44911,N_44106,N_44186);
xnor U44912 (N_44912,N_44353,N_44063);
xnor U44913 (N_44913,N_44381,N_44344);
and U44914 (N_44914,N_44336,N_44134);
or U44915 (N_44915,N_44434,N_44445);
and U44916 (N_44916,N_44069,N_44265);
or U44917 (N_44917,N_44289,N_44073);
nand U44918 (N_44918,N_44276,N_44450);
and U44919 (N_44919,N_44259,N_44403);
nand U44920 (N_44920,N_44254,N_44177);
xnor U44921 (N_44921,N_44085,N_44016);
or U44922 (N_44922,N_44222,N_44262);
xnor U44923 (N_44923,N_44297,N_44188);
or U44924 (N_44924,N_44364,N_44246);
and U44925 (N_44925,N_44494,N_44190);
nor U44926 (N_44926,N_44130,N_44306);
or U44927 (N_44927,N_44272,N_44222);
nand U44928 (N_44928,N_44007,N_44202);
nor U44929 (N_44929,N_44065,N_44411);
xor U44930 (N_44930,N_44126,N_44176);
xor U44931 (N_44931,N_44441,N_44039);
nand U44932 (N_44932,N_44090,N_44274);
or U44933 (N_44933,N_44279,N_44184);
nand U44934 (N_44934,N_44206,N_44242);
and U44935 (N_44935,N_44156,N_44497);
or U44936 (N_44936,N_44179,N_44144);
xor U44937 (N_44937,N_44204,N_44077);
nand U44938 (N_44938,N_44465,N_44421);
and U44939 (N_44939,N_44494,N_44363);
and U44940 (N_44940,N_44382,N_44387);
nand U44941 (N_44941,N_44330,N_44134);
nand U44942 (N_44942,N_44194,N_44494);
xnor U44943 (N_44943,N_44468,N_44384);
nor U44944 (N_44944,N_44435,N_44256);
nor U44945 (N_44945,N_44478,N_44154);
or U44946 (N_44946,N_44009,N_44210);
nand U44947 (N_44947,N_44167,N_44195);
xor U44948 (N_44948,N_44352,N_44454);
or U44949 (N_44949,N_44281,N_44087);
and U44950 (N_44950,N_44333,N_44342);
and U44951 (N_44951,N_44461,N_44268);
nand U44952 (N_44952,N_44317,N_44449);
and U44953 (N_44953,N_44056,N_44199);
nand U44954 (N_44954,N_44087,N_44129);
and U44955 (N_44955,N_44391,N_44322);
xnor U44956 (N_44956,N_44241,N_44346);
or U44957 (N_44957,N_44433,N_44056);
nand U44958 (N_44958,N_44441,N_44098);
xor U44959 (N_44959,N_44264,N_44128);
nor U44960 (N_44960,N_44015,N_44411);
nand U44961 (N_44961,N_44382,N_44490);
xor U44962 (N_44962,N_44065,N_44003);
nor U44963 (N_44963,N_44000,N_44045);
nor U44964 (N_44964,N_44289,N_44240);
or U44965 (N_44965,N_44041,N_44143);
xnor U44966 (N_44966,N_44120,N_44105);
nand U44967 (N_44967,N_44089,N_44329);
and U44968 (N_44968,N_44392,N_44008);
and U44969 (N_44969,N_44059,N_44438);
and U44970 (N_44970,N_44142,N_44383);
and U44971 (N_44971,N_44005,N_44242);
and U44972 (N_44972,N_44431,N_44188);
xnor U44973 (N_44973,N_44098,N_44118);
nand U44974 (N_44974,N_44138,N_44248);
and U44975 (N_44975,N_44252,N_44061);
nor U44976 (N_44976,N_44009,N_44051);
nand U44977 (N_44977,N_44486,N_44073);
nor U44978 (N_44978,N_44000,N_44413);
and U44979 (N_44979,N_44017,N_44147);
nor U44980 (N_44980,N_44192,N_44141);
nand U44981 (N_44981,N_44064,N_44460);
or U44982 (N_44982,N_44352,N_44255);
xor U44983 (N_44983,N_44143,N_44428);
xnor U44984 (N_44984,N_44430,N_44066);
and U44985 (N_44985,N_44303,N_44230);
nor U44986 (N_44986,N_44171,N_44268);
and U44987 (N_44987,N_44313,N_44096);
nor U44988 (N_44988,N_44483,N_44488);
and U44989 (N_44989,N_44184,N_44305);
nor U44990 (N_44990,N_44336,N_44460);
and U44991 (N_44991,N_44330,N_44130);
xor U44992 (N_44992,N_44361,N_44026);
nand U44993 (N_44993,N_44490,N_44396);
or U44994 (N_44994,N_44397,N_44253);
nand U44995 (N_44995,N_44374,N_44013);
and U44996 (N_44996,N_44246,N_44019);
nand U44997 (N_44997,N_44091,N_44361);
xnor U44998 (N_44998,N_44321,N_44405);
nor U44999 (N_44999,N_44162,N_44257);
nand U45000 (N_45000,N_44997,N_44953);
or U45001 (N_45001,N_44947,N_44633);
xor U45002 (N_45002,N_44583,N_44928);
nor U45003 (N_45003,N_44627,N_44555);
and U45004 (N_45004,N_44617,N_44973);
nor U45005 (N_45005,N_44670,N_44554);
xnor U45006 (N_45006,N_44578,N_44610);
xor U45007 (N_45007,N_44825,N_44762);
and U45008 (N_45008,N_44969,N_44993);
nand U45009 (N_45009,N_44685,N_44647);
nor U45010 (N_45010,N_44986,N_44641);
xnor U45011 (N_45011,N_44951,N_44924);
xor U45012 (N_45012,N_44939,N_44576);
nand U45013 (N_45013,N_44923,N_44797);
xnor U45014 (N_45014,N_44669,N_44955);
nor U45015 (N_45015,N_44861,N_44862);
or U45016 (N_45016,N_44908,N_44764);
and U45017 (N_45017,N_44952,N_44736);
or U45018 (N_45018,N_44571,N_44638);
nand U45019 (N_45019,N_44719,N_44655);
or U45020 (N_45020,N_44567,N_44806);
or U45021 (N_45021,N_44910,N_44788);
and U45022 (N_45022,N_44602,N_44905);
xor U45023 (N_45023,N_44916,N_44799);
nand U45024 (N_45024,N_44894,N_44998);
and U45025 (N_45025,N_44849,N_44711);
xnor U45026 (N_45026,N_44657,N_44569);
xnor U45027 (N_45027,N_44625,N_44970);
nand U45028 (N_45028,N_44982,N_44903);
nand U45029 (N_45029,N_44748,N_44687);
nor U45030 (N_45030,N_44580,N_44968);
and U45031 (N_45031,N_44902,N_44613);
xnor U45032 (N_45032,N_44850,N_44798);
and U45033 (N_45033,N_44689,N_44786);
and U45034 (N_45034,N_44785,N_44620);
nand U45035 (N_45035,N_44559,N_44887);
nor U45036 (N_45036,N_44726,N_44747);
nor U45037 (N_45037,N_44686,N_44954);
nor U45038 (N_45038,N_44611,N_44824);
or U45039 (N_45039,N_44672,N_44846);
nand U45040 (N_45040,N_44512,N_44929);
nor U45041 (N_45041,N_44558,N_44911);
or U45042 (N_45042,N_44722,N_44515);
or U45043 (N_45043,N_44691,N_44503);
nor U45044 (N_45044,N_44796,N_44618);
xor U45045 (N_45045,N_44933,N_44832);
nor U45046 (N_45046,N_44581,N_44541);
nand U45047 (N_45047,N_44684,N_44716);
nand U45048 (N_45048,N_44906,N_44873);
xor U45049 (N_45049,N_44584,N_44907);
or U45050 (N_45050,N_44866,N_44771);
and U45051 (N_45051,N_44813,N_44889);
nor U45052 (N_45052,N_44508,N_44755);
xor U45053 (N_45053,N_44504,N_44536);
or U45054 (N_45054,N_44869,N_44946);
nor U45055 (N_45055,N_44974,N_44848);
and U45056 (N_45056,N_44802,N_44934);
or U45057 (N_45057,N_44978,N_44704);
or U45058 (N_45058,N_44858,N_44718);
and U45059 (N_45059,N_44740,N_44847);
or U45060 (N_45060,N_44592,N_44927);
and U45061 (N_45061,N_44589,N_44826);
xnor U45062 (N_45062,N_44792,N_44821);
xor U45063 (N_45063,N_44741,N_44958);
or U45064 (N_45064,N_44888,N_44572);
nor U45065 (N_45065,N_44823,N_44738);
xnor U45066 (N_45066,N_44770,N_44604);
and U45067 (N_45067,N_44853,N_44668);
nand U45068 (N_45068,N_44537,N_44895);
xor U45069 (N_45069,N_44854,N_44658);
xor U45070 (N_45070,N_44517,N_44678);
xnor U45071 (N_45071,N_44553,N_44695);
and U45072 (N_45072,N_44865,N_44674);
nand U45073 (N_45073,N_44676,N_44960);
and U45074 (N_45074,N_44949,N_44944);
nand U45075 (N_45075,N_44587,N_44544);
nand U45076 (N_45076,N_44760,N_44656);
nand U45077 (N_45077,N_44876,N_44995);
nor U45078 (N_45078,N_44639,N_44819);
and U45079 (N_45079,N_44715,N_44937);
or U45080 (N_45080,N_44809,N_44883);
and U45081 (N_45081,N_44502,N_44751);
nor U45082 (N_45082,N_44519,N_44521);
and U45083 (N_45083,N_44506,N_44675);
and U45084 (N_45084,N_44935,N_44745);
or U45085 (N_45085,N_44662,N_44977);
nor U45086 (N_45086,N_44758,N_44752);
nand U45087 (N_45087,N_44708,N_44829);
or U45088 (N_45088,N_44963,N_44734);
nand U45089 (N_45089,N_44983,N_44549);
nor U45090 (N_45090,N_44609,N_44667);
xnor U45091 (N_45091,N_44932,N_44579);
or U45092 (N_45092,N_44817,N_44940);
nand U45093 (N_45093,N_44612,N_44661);
and U45094 (N_45094,N_44931,N_44863);
or U45095 (N_45095,N_44828,N_44867);
nand U45096 (N_45096,N_44507,N_44696);
nand U45097 (N_45097,N_44531,N_44720);
and U45098 (N_45098,N_44652,N_44759);
nand U45099 (N_45099,N_44733,N_44831);
xnor U45100 (N_45100,N_44874,N_44925);
xor U45101 (N_45101,N_44956,N_44976);
xnor U45102 (N_45102,N_44631,N_44841);
xnor U45103 (N_45103,N_44980,N_44897);
nand U45104 (N_45104,N_44582,N_44648);
and U45105 (N_45105,N_44607,N_44624);
or U45106 (N_45106,N_44717,N_44896);
or U45107 (N_45107,N_44833,N_44591);
nor U45108 (N_45108,N_44945,N_44560);
and U45109 (N_45109,N_44965,N_44516);
nor U45110 (N_45110,N_44653,N_44810);
nor U45111 (N_45111,N_44706,N_44855);
nand U45112 (N_45112,N_44816,N_44769);
or U45113 (N_45113,N_44514,N_44710);
nor U45114 (N_45114,N_44520,N_44904);
nand U45115 (N_45115,N_44709,N_44790);
xnor U45116 (N_45116,N_44938,N_44860);
xor U45117 (N_45117,N_44509,N_44763);
xnor U45118 (N_45118,N_44577,N_44900);
nor U45119 (N_45119,N_44681,N_44535);
or U45120 (N_45120,N_44981,N_44749);
xnor U45121 (N_45121,N_44814,N_44574);
and U45122 (N_45122,N_44804,N_44562);
and U45123 (N_45123,N_44619,N_44961);
xor U45124 (N_45124,N_44742,N_44550);
or U45125 (N_45125,N_44871,N_44753);
nand U45126 (N_45126,N_44842,N_44513);
or U45127 (N_45127,N_44556,N_44922);
or U45128 (N_45128,N_44728,N_44529);
and U45129 (N_45129,N_44626,N_44999);
xnor U45130 (N_45130,N_44856,N_44530);
and U45131 (N_45131,N_44975,N_44875);
and U45132 (N_45132,N_44926,N_44533);
xnor U45133 (N_45133,N_44901,N_44979);
or U45134 (N_45134,N_44596,N_44701);
xnor U45135 (N_45135,N_44818,N_44527);
nand U45136 (N_45136,N_44528,N_44878);
or U45137 (N_45137,N_44663,N_44700);
and U45138 (N_45138,N_44651,N_44987);
nor U45139 (N_45139,N_44996,N_44721);
nor U45140 (N_45140,N_44899,N_44845);
nand U45141 (N_45141,N_44789,N_44586);
xor U45142 (N_45142,N_44714,N_44561);
xor U45143 (N_45143,N_44957,N_44914);
and U45144 (N_45144,N_44646,N_44615);
and U45145 (N_45145,N_44984,N_44693);
nor U45146 (N_45146,N_44761,N_44882);
and U45147 (N_45147,N_44784,N_44640);
nand U45148 (N_45148,N_44551,N_44967);
nor U45149 (N_45149,N_44827,N_44568);
xnor U45150 (N_45150,N_44563,N_44660);
or U45151 (N_45151,N_44851,N_44893);
and U45152 (N_45152,N_44565,N_44737);
or U45153 (N_45153,N_44622,N_44526);
nor U45154 (N_45154,N_44872,N_44781);
or U45155 (N_45155,N_44636,N_44666);
or U45156 (N_45156,N_44540,N_44608);
nor U45157 (N_45157,N_44634,N_44705);
xnor U45158 (N_45158,N_44621,N_44650);
nor U45159 (N_45159,N_44881,N_44870);
or U45160 (N_45160,N_44912,N_44884);
and U45161 (N_45161,N_44917,N_44595);
nor U45162 (N_45162,N_44523,N_44898);
nor U45163 (N_45163,N_44776,N_44557);
or U45164 (N_45164,N_44918,N_44552);
nand U45165 (N_45165,N_44642,N_44864);
and U45166 (N_45166,N_44564,N_44852);
or U45167 (N_45167,N_44546,N_44843);
nor U45168 (N_45168,N_44600,N_44962);
or U45169 (N_45169,N_44750,N_44692);
or U45170 (N_45170,N_44746,N_44774);
and U45171 (N_45171,N_44773,N_44594);
xor U45172 (N_45172,N_44886,N_44707);
nor U45173 (N_45173,N_44812,N_44915);
nor U45174 (N_45174,N_44808,N_44534);
or U45175 (N_45175,N_44644,N_44511);
and U45176 (N_45176,N_44623,N_44683);
and U45177 (N_45177,N_44545,N_44877);
and U45178 (N_45178,N_44522,N_44988);
nor U45179 (N_45179,N_44913,N_44834);
nand U45180 (N_45180,N_44801,N_44679);
and U45181 (N_45181,N_44820,N_44724);
xor U45182 (N_45182,N_44767,N_44635);
nand U45183 (N_45183,N_44765,N_44501);
or U45184 (N_45184,N_44673,N_44959);
nand U45185 (N_45185,N_44505,N_44713);
xor U45186 (N_45186,N_44548,N_44880);
nor U45187 (N_45187,N_44598,N_44702);
nor U45188 (N_45188,N_44815,N_44891);
or U45189 (N_45189,N_44989,N_44838);
xor U45190 (N_45190,N_44787,N_44654);
and U45191 (N_45191,N_44778,N_44892);
xor U45192 (N_45192,N_44777,N_44920);
nand U45193 (N_45193,N_44588,N_44605);
and U45194 (N_45194,N_44991,N_44699);
or U45195 (N_45195,N_44739,N_44964);
and U45196 (N_45196,N_44775,N_44575);
nand U45197 (N_45197,N_44542,N_44921);
nor U45198 (N_45198,N_44659,N_44682);
and U45199 (N_45199,N_44630,N_44766);
nand U45200 (N_45200,N_44723,N_44791);
xnor U45201 (N_45201,N_44570,N_44538);
xnor U45202 (N_45202,N_44942,N_44990);
and U45203 (N_45203,N_44840,N_44677);
xor U45204 (N_45204,N_44800,N_44698);
nand U45205 (N_45205,N_44950,N_44839);
xor U45206 (N_45206,N_44606,N_44772);
and U45207 (N_45207,N_44879,N_44930);
nor U45208 (N_45208,N_44868,N_44779);
nand U45209 (N_45209,N_44744,N_44835);
xor U45210 (N_45210,N_44730,N_44703);
xor U45211 (N_45211,N_44671,N_44783);
and U45212 (N_45212,N_44628,N_44972);
xor U45213 (N_45213,N_44518,N_44525);
xnor U45214 (N_45214,N_44500,N_44601);
and U45215 (N_45215,N_44857,N_44941);
xor U45216 (N_45216,N_44756,N_44597);
or U45217 (N_45217,N_44593,N_44768);
and U45218 (N_45218,N_44948,N_44690);
and U45219 (N_45219,N_44795,N_44732);
nand U45220 (N_45220,N_44590,N_44782);
nor U45221 (N_45221,N_44807,N_44532);
or U45222 (N_45222,N_44510,N_44725);
nor U45223 (N_45223,N_44712,N_44697);
xor U45224 (N_45224,N_44794,N_44909);
or U45225 (N_45225,N_44637,N_44919);
xnor U45226 (N_45226,N_44688,N_44837);
or U45227 (N_45227,N_44743,N_44727);
xnor U45228 (N_45228,N_44943,N_44992);
nor U45229 (N_45229,N_44585,N_44645);
or U45230 (N_45230,N_44844,N_44649);
xor U45231 (N_45231,N_44539,N_44822);
nor U45232 (N_45232,N_44664,N_44694);
nand U45233 (N_45233,N_44616,N_44524);
nand U45234 (N_45234,N_44543,N_44731);
and U45235 (N_45235,N_44859,N_44603);
or U45236 (N_45236,N_44971,N_44780);
or U45237 (N_45237,N_44985,N_44566);
and U45238 (N_45238,N_44757,N_44994);
xnor U45239 (N_45239,N_44966,N_44614);
and U45240 (N_45240,N_44793,N_44632);
or U45241 (N_45241,N_44629,N_44665);
nor U45242 (N_45242,N_44735,N_44643);
or U45243 (N_45243,N_44836,N_44936);
and U45244 (N_45244,N_44573,N_44885);
nand U45245 (N_45245,N_44803,N_44680);
and U45246 (N_45246,N_44547,N_44811);
nor U45247 (N_45247,N_44729,N_44599);
or U45248 (N_45248,N_44805,N_44890);
or U45249 (N_45249,N_44754,N_44830);
nand U45250 (N_45250,N_44611,N_44692);
nand U45251 (N_45251,N_44959,N_44831);
xor U45252 (N_45252,N_44520,N_44984);
xnor U45253 (N_45253,N_44633,N_44981);
or U45254 (N_45254,N_44744,N_44960);
xnor U45255 (N_45255,N_44939,N_44943);
or U45256 (N_45256,N_44992,N_44916);
and U45257 (N_45257,N_44525,N_44942);
xor U45258 (N_45258,N_44855,N_44737);
nand U45259 (N_45259,N_44924,N_44827);
nand U45260 (N_45260,N_44549,N_44748);
xor U45261 (N_45261,N_44529,N_44967);
or U45262 (N_45262,N_44660,N_44794);
xnor U45263 (N_45263,N_44552,N_44888);
or U45264 (N_45264,N_44661,N_44901);
nor U45265 (N_45265,N_44652,N_44726);
or U45266 (N_45266,N_44944,N_44535);
or U45267 (N_45267,N_44948,N_44613);
nand U45268 (N_45268,N_44584,N_44558);
xnor U45269 (N_45269,N_44679,N_44518);
nand U45270 (N_45270,N_44910,N_44551);
nand U45271 (N_45271,N_44736,N_44558);
or U45272 (N_45272,N_44573,N_44567);
nor U45273 (N_45273,N_44922,N_44879);
and U45274 (N_45274,N_44557,N_44977);
or U45275 (N_45275,N_44548,N_44643);
nor U45276 (N_45276,N_44712,N_44831);
nor U45277 (N_45277,N_44848,N_44594);
or U45278 (N_45278,N_44926,N_44816);
nand U45279 (N_45279,N_44749,N_44845);
nand U45280 (N_45280,N_44688,N_44965);
and U45281 (N_45281,N_44901,N_44557);
nor U45282 (N_45282,N_44805,N_44977);
xnor U45283 (N_45283,N_44840,N_44589);
and U45284 (N_45284,N_44896,N_44969);
and U45285 (N_45285,N_44962,N_44545);
nor U45286 (N_45286,N_44957,N_44906);
and U45287 (N_45287,N_44961,N_44848);
or U45288 (N_45288,N_44727,N_44678);
nor U45289 (N_45289,N_44777,N_44736);
and U45290 (N_45290,N_44632,N_44682);
nor U45291 (N_45291,N_44942,N_44930);
xnor U45292 (N_45292,N_44978,N_44699);
xor U45293 (N_45293,N_44739,N_44884);
and U45294 (N_45294,N_44958,N_44821);
nor U45295 (N_45295,N_44801,N_44579);
and U45296 (N_45296,N_44864,N_44712);
or U45297 (N_45297,N_44921,N_44824);
or U45298 (N_45298,N_44791,N_44656);
nor U45299 (N_45299,N_44771,N_44792);
and U45300 (N_45300,N_44633,N_44779);
or U45301 (N_45301,N_44581,N_44949);
nor U45302 (N_45302,N_44689,N_44807);
nor U45303 (N_45303,N_44907,N_44951);
nand U45304 (N_45304,N_44702,N_44721);
xnor U45305 (N_45305,N_44838,N_44796);
nand U45306 (N_45306,N_44780,N_44720);
and U45307 (N_45307,N_44552,N_44526);
xnor U45308 (N_45308,N_44696,N_44840);
or U45309 (N_45309,N_44905,N_44538);
or U45310 (N_45310,N_44579,N_44635);
and U45311 (N_45311,N_44752,N_44841);
and U45312 (N_45312,N_44853,N_44518);
nor U45313 (N_45313,N_44792,N_44518);
or U45314 (N_45314,N_44565,N_44971);
nor U45315 (N_45315,N_44756,N_44856);
or U45316 (N_45316,N_44703,N_44741);
or U45317 (N_45317,N_44529,N_44686);
nand U45318 (N_45318,N_44649,N_44785);
or U45319 (N_45319,N_44535,N_44542);
and U45320 (N_45320,N_44901,N_44853);
xor U45321 (N_45321,N_44859,N_44849);
nor U45322 (N_45322,N_44644,N_44609);
xnor U45323 (N_45323,N_44583,N_44987);
or U45324 (N_45324,N_44527,N_44679);
xor U45325 (N_45325,N_44533,N_44557);
and U45326 (N_45326,N_44685,N_44748);
nor U45327 (N_45327,N_44604,N_44601);
nor U45328 (N_45328,N_44643,N_44880);
and U45329 (N_45329,N_44785,N_44689);
nor U45330 (N_45330,N_44519,N_44659);
nor U45331 (N_45331,N_44798,N_44871);
xnor U45332 (N_45332,N_44809,N_44941);
xnor U45333 (N_45333,N_44511,N_44809);
or U45334 (N_45334,N_44690,N_44501);
or U45335 (N_45335,N_44624,N_44506);
xnor U45336 (N_45336,N_44906,N_44544);
nand U45337 (N_45337,N_44752,N_44524);
nand U45338 (N_45338,N_44518,N_44534);
and U45339 (N_45339,N_44854,N_44604);
or U45340 (N_45340,N_44832,N_44862);
and U45341 (N_45341,N_44582,N_44679);
nand U45342 (N_45342,N_44702,N_44943);
xnor U45343 (N_45343,N_44667,N_44787);
and U45344 (N_45344,N_44620,N_44743);
or U45345 (N_45345,N_44586,N_44955);
xor U45346 (N_45346,N_44847,N_44900);
or U45347 (N_45347,N_44547,N_44839);
xnor U45348 (N_45348,N_44538,N_44812);
nor U45349 (N_45349,N_44611,N_44988);
or U45350 (N_45350,N_44514,N_44833);
nor U45351 (N_45351,N_44796,N_44839);
nand U45352 (N_45352,N_44781,N_44539);
nor U45353 (N_45353,N_44604,N_44707);
and U45354 (N_45354,N_44694,N_44767);
xnor U45355 (N_45355,N_44522,N_44511);
and U45356 (N_45356,N_44621,N_44652);
nor U45357 (N_45357,N_44530,N_44613);
nor U45358 (N_45358,N_44922,N_44667);
and U45359 (N_45359,N_44803,N_44776);
nor U45360 (N_45360,N_44872,N_44802);
and U45361 (N_45361,N_44731,N_44771);
xor U45362 (N_45362,N_44666,N_44997);
nor U45363 (N_45363,N_44871,N_44735);
nand U45364 (N_45364,N_44887,N_44888);
or U45365 (N_45365,N_44534,N_44556);
nor U45366 (N_45366,N_44593,N_44926);
or U45367 (N_45367,N_44847,N_44914);
nor U45368 (N_45368,N_44544,N_44777);
xnor U45369 (N_45369,N_44897,N_44986);
nor U45370 (N_45370,N_44520,N_44841);
nor U45371 (N_45371,N_44813,N_44831);
and U45372 (N_45372,N_44947,N_44527);
xnor U45373 (N_45373,N_44536,N_44768);
or U45374 (N_45374,N_44892,N_44968);
and U45375 (N_45375,N_44508,N_44567);
nor U45376 (N_45376,N_44893,N_44736);
and U45377 (N_45377,N_44849,N_44887);
and U45378 (N_45378,N_44945,N_44789);
nor U45379 (N_45379,N_44538,N_44598);
nand U45380 (N_45380,N_44572,N_44788);
and U45381 (N_45381,N_44799,N_44503);
xnor U45382 (N_45382,N_44900,N_44649);
xor U45383 (N_45383,N_44824,N_44985);
nand U45384 (N_45384,N_44623,N_44501);
and U45385 (N_45385,N_44572,N_44979);
nand U45386 (N_45386,N_44964,N_44727);
and U45387 (N_45387,N_44882,N_44573);
or U45388 (N_45388,N_44616,N_44767);
nor U45389 (N_45389,N_44529,N_44553);
nor U45390 (N_45390,N_44762,N_44558);
or U45391 (N_45391,N_44916,N_44926);
or U45392 (N_45392,N_44743,N_44637);
or U45393 (N_45393,N_44533,N_44599);
nor U45394 (N_45394,N_44856,N_44947);
and U45395 (N_45395,N_44623,N_44700);
or U45396 (N_45396,N_44579,N_44849);
xnor U45397 (N_45397,N_44720,N_44550);
or U45398 (N_45398,N_44690,N_44598);
or U45399 (N_45399,N_44733,N_44646);
nand U45400 (N_45400,N_44879,N_44697);
nand U45401 (N_45401,N_44880,N_44514);
nand U45402 (N_45402,N_44907,N_44668);
nand U45403 (N_45403,N_44664,N_44724);
xor U45404 (N_45404,N_44966,N_44503);
nand U45405 (N_45405,N_44840,N_44572);
nor U45406 (N_45406,N_44780,N_44744);
nor U45407 (N_45407,N_44984,N_44775);
nor U45408 (N_45408,N_44897,N_44720);
and U45409 (N_45409,N_44972,N_44990);
and U45410 (N_45410,N_44510,N_44536);
and U45411 (N_45411,N_44804,N_44531);
nand U45412 (N_45412,N_44772,N_44757);
nand U45413 (N_45413,N_44781,N_44915);
nor U45414 (N_45414,N_44902,N_44541);
or U45415 (N_45415,N_44507,N_44539);
xor U45416 (N_45416,N_44838,N_44786);
or U45417 (N_45417,N_44627,N_44544);
nor U45418 (N_45418,N_44761,N_44743);
nand U45419 (N_45419,N_44819,N_44793);
xnor U45420 (N_45420,N_44729,N_44606);
and U45421 (N_45421,N_44721,N_44598);
or U45422 (N_45422,N_44866,N_44939);
nor U45423 (N_45423,N_44914,N_44536);
or U45424 (N_45424,N_44676,N_44983);
and U45425 (N_45425,N_44772,N_44529);
and U45426 (N_45426,N_44524,N_44823);
nand U45427 (N_45427,N_44632,N_44713);
nand U45428 (N_45428,N_44663,N_44540);
nand U45429 (N_45429,N_44518,N_44723);
xor U45430 (N_45430,N_44938,N_44903);
xnor U45431 (N_45431,N_44775,N_44751);
nand U45432 (N_45432,N_44822,N_44567);
and U45433 (N_45433,N_44931,N_44656);
nand U45434 (N_45434,N_44742,N_44885);
or U45435 (N_45435,N_44666,N_44503);
nor U45436 (N_45436,N_44679,N_44770);
or U45437 (N_45437,N_44839,N_44746);
and U45438 (N_45438,N_44525,N_44779);
nand U45439 (N_45439,N_44722,N_44901);
xor U45440 (N_45440,N_44595,N_44587);
nor U45441 (N_45441,N_44851,N_44705);
or U45442 (N_45442,N_44722,N_44680);
or U45443 (N_45443,N_44930,N_44839);
or U45444 (N_45444,N_44946,N_44569);
nor U45445 (N_45445,N_44939,N_44824);
xnor U45446 (N_45446,N_44532,N_44783);
nor U45447 (N_45447,N_44715,N_44891);
xor U45448 (N_45448,N_44754,N_44647);
nor U45449 (N_45449,N_44977,N_44904);
and U45450 (N_45450,N_44664,N_44589);
and U45451 (N_45451,N_44543,N_44642);
xnor U45452 (N_45452,N_44561,N_44621);
nor U45453 (N_45453,N_44544,N_44909);
nand U45454 (N_45454,N_44974,N_44912);
or U45455 (N_45455,N_44940,N_44579);
nand U45456 (N_45456,N_44995,N_44783);
nor U45457 (N_45457,N_44948,N_44711);
and U45458 (N_45458,N_44663,N_44876);
xor U45459 (N_45459,N_44716,N_44913);
xnor U45460 (N_45460,N_44826,N_44735);
or U45461 (N_45461,N_44786,N_44626);
and U45462 (N_45462,N_44524,N_44526);
or U45463 (N_45463,N_44874,N_44647);
nor U45464 (N_45464,N_44587,N_44549);
nor U45465 (N_45465,N_44839,N_44853);
or U45466 (N_45466,N_44935,N_44582);
and U45467 (N_45467,N_44539,N_44806);
nand U45468 (N_45468,N_44783,N_44788);
nand U45469 (N_45469,N_44955,N_44884);
nand U45470 (N_45470,N_44901,N_44841);
xnor U45471 (N_45471,N_44611,N_44558);
xnor U45472 (N_45472,N_44748,N_44857);
or U45473 (N_45473,N_44594,N_44655);
nand U45474 (N_45474,N_44936,N_44975);
nand U45475 (N_45475,N_44599,N_44624);
and U45476 (N_45476,N_44671,N_44607);
nor U45477 (N_45477,N_44541,N_44664);
nor U45478 (N_45478,N_44823,N_44968);
or U45479 (N_45479,N_44511,N_44588);
and U45480 (N_45480,N_44787,N_44917);
xor U45481 (N_45481,N_44654,N_44503);
or U45482 (N_45482,N_44803,N_44878);
or U45483 (N_45483,N_44843,N_44841);
xor U45484 (N_45484,N_44713,N_44688);
nor U45485 (N_45485,N_44581,N_44643);
and U45486 (N_45486,N_44846,N_44882);
xor U45487 (N_45487,N_44861,N_44585);
xnor U45488 (N_45488,N_44955,N_44616);
nor U45489 (N_45489,N_44962,N_44924);
xor U45490 (N_45490,N_44548,N_44797);
nor U45491 (N_45491,N_44698,N_44879);
nor U45492 (N_45492,N_44688,N_44896);
or U45493 (N_45493,N_44700,N_44555);
nor U45494 (N_45494,N_44892,N_44644);
nor U45495 (N_45495,N_44612,N_44927);
nor U45496 (N_45496,N_44723,N_44640);
nor U45497 (N_45497,N_44903,N_44966);
nand U45498 (N_45498,N_44663,N_44867);
nor U45499 (N_45499,N_44939,N_44698);
and U45500 (N_45500,N_45225,N_45084);
nor U45501 (N_45501,N_45138,N_45258);
and U45502 (N_45502,N_45127,N_45000);
xor U45503 (N_45503,N_45024,N_45367);
nor U45504 (N_45504,N_45406,N_45214);
and U45505 (N_45505,N_45354,N_45451);
nand U45506 (N_45506,N_45385,N_45414);
and U45507 (N_45507,N_45066,N_45231);
nor U45508 (N_45508,N_45110,N_45409);
nand U45509 (N_45509,N_45198,N_45265);
or U45510 (N_45510,N_45255,N_45310);
and U45511 (N_45511,N_45461,N_45186);
and U45512 (N_45512,N_45471,N_45152);
xnor U45513 (N_45513,N_45318,N_45087);
nand U45514 (N_45514,N_45140,N_45288);
nand U45515 (N_45515,N_45311,N_45041);
nand U45516 (N_45516,N_45182,N_45382);
nor U45517 (N_45517,N_45336,N_45272);
nor U45518 (N_45518,N_45349,N_45492);
nor U45519 (N_45519,N_45365,N_45067);
xnor U45520 (N_45520,N_45165,N_45008);
nor U45521 (N_45521,N_45172,N_45257);
and U45522 (N_45522,N_45259,N_45203);
nand U45523 (N_45523,N_45249,N_45074);
and U45524 (N_45524,N_45237,N_45175);
nor U45525 (N_45525,N_45150,N_45449);
nand U45526 (N_45526,N_45162,N_45435);
or U45527 (N_45527,N_45369,N_45429);
nand U45528 (N_45528,N_45490,N_45081);
and U45529 (N_45529,N_45443,N_45357);
nand U45530 (N_45530,N_45340,N_45242);
nand U45531 (N_45531,N_45358,N_45082);
nand U45532 (N_45532,N_45380,N_45489);
nor U45533 (N_45533,N_45496,N_45252);
xor U45534 (N_45534,N_45405,N_45122);
and U45535 (N_45535,N_45463,N_45497);
nor U45536 (N_45536,N_45038,N_45469);
nor U45537 (N_45537,N_45168,N_45401);
or U45538 (N_45538,N_45109,N_45283);
nor U45539 (N_45539,N_45313,N_45196);
nor U45540 (N_45540,N_45126,N_45077);
or U45541 (N_45541,N_45171,N_45476);
nor U45542 (N_45542,N_45091,N_45247);
nor U45543 (N_45543,N_45013,N_45356);
nor U45544 (N_45544,N_45454,N_45246);
and U45545 (N_45545,N_45072,N_45188);
xnor U45546 (N_45546,N_45190,N_45302);
or U45547 (N_45547,N_45345,N_45238);
xnor U45548 (N_45548,N_45235,N_45053);
nor U45549 (N_45549,N_45210,N_45393);
nand U45550 (N_45550,N_45204,N_45460);
and U45551 (N_45551,N_45381,N_45398);
and U45552 (N_45552,N_45085,N_45342);
nor U45553 (N_45553,N_45105,N_45289);
or U45554 (N_45554,N_45433,N_45417);
and U45555 (N_45555,N_45287,N_45125);
nand U45556 (N_45556,N_45071,N_45120);
nor U45557 (N_45557,N_45177,N_45148);
xnor U45558 (N_45558,N_45379,N_45130);
nand U45559 (N_45559,N_45498,N_45200);
nor U45560 (N_45560,N_45319,N_45368);
xnor U45561 (N_45561,N_45467,N_45108);
xor U45562 (N_45562,N_45309,N_45431);
xor U45563 (N_45563,N_45346,N_45480);
or U45564 (N_45564,N_45452,N_45026);
and U45565 (N_45565,N_45223,N_45332);
or U45566 (N_45566,N_45132,N_45457);
nor U45567 (N_45567,N_45014,N_45093);
or U45568 (N_45568,N_45201,N_45388);
xor U45569 (N_45569,N_45377,N_45320);
and U45570 (N_45570,N_45392,N_45475);
and U45571 (N_45571,N_45391,N_45327);
or U45572 (N_45572,N_45215,N_45364);
and U45573 (N_45573,N_45039,N_45439);
or U45574 (N_45574,N_45396,N_45415);
and U45575 (N_45575,N_45173,N_45139);
or U45576 (N_45576,N_45195,N_45058);
and U45577 (N_45577,N_45297,N_45294);
xor U45578 (N_45578,N_45154,N_45446);
xnor U45579 (N_45579,N_45285,N_45260);
nand U45580 (N_45580,N_45207,N_45020);
or U45581 (N_45581,N_45179,N_45301);
xnor U45582 (N_45582,N_45424,N_45456);
or U45583 (N_45583,N_45135,N_45012);
or U45584 (N_45584,N_45021,N_45176);
and U45585 (N_45585,N_45104,N_45221);
nor U45586 (N_45586,N_45194,N_45158);
and U45587 (N_45587,N_45394,N_45334);
or U45588 (N_45588,N_45161,N_45212);
and U45589 (N_45589,N_45033,N_45184);
and U45590 (N_45590,N_45046,N_45052);
nor U45591 (N_45591,N_45268,N_45006);
nand U45592 (N_45592,N_45253,N_45236);
nand U45593 (N_45593,N_45011,N_45141);
nand U45594 (N_45594,N_45389,N_45015);
xor U45595 (N_45595,N_45434,N_45050);
nand U45596 (N_45596,N_45404,N_45432);
or U45597 (N_45597,N_45232,N_45286);
or U45598 (N_45598,N_45488,N_45244);
and U45599 (N_45599,N_45436,N_45151);
nor U45600 (N_45600,N_45211,N_45222);
nor U45601 (N_45601,N_45267,N_45384);
xnor U45602 (N_45602,N_45484,N_45220);
and U45603 (N_45603,N_45002,N_45437);
nand U45604 (N_45604,N_45464,N_45295);
nand U45605 (N_45605,N_45022,N_45217);
nand U45606 (N_45606,N_45465,N_45183);
nand U45607 (N_45607,N_45343,N_45192);
nand U45608 (N_45608,N_45224,N_45123);
nand U45609 (N_45609,N_45322,N_45054);
and U45610 (N_45610,N_45450,N_45241);
or U45611 (N_45611,N_45118,N_45291);
xnor U45612 (N_45612,N_45423,N_45086);
or U45613 (N_45613,N_45339,N_45124);
nand U45614 (N_45614,N_45070,N_45315);
nor U45615 (N_45615,N_45083,N_45073);
xor U45616 (N_45616,N_45029,N_45305);
nor U45617 (N_45617,N_45037,N_45106);
nor U45618 (N_45618,N_45282,N_45479);
nand U45619 (N_45619,N_45097,N_45303);
xnor U45620 (N_45620,N_45193,N_45482);
and U45621 (N_45621,N_45240,N_45185);
xor U45622 (N_45622,N_45308,N_45411);
xor U45623 (N_45623,N_45229,N_45049);
and U45624 (N_45624,N_45261,N_45060);
nand U45625 (N_45625,N_45474,N_45116);
nand U45626 (N_45626,N_45218,N_45191);
or U45627 (N_45627,N_45157,N_45057);
or U45628 (N_45628,N_45298,N_45239);
and U45629 (N_45629,N_45051,N_45254);
and U45630 (N_45630,N_45062,N_45216);
or U45631 (N_45631,N_45266,N_45293);
xor U45632 (N_45632,N_45316,N_45090);
and U45633 (N_45633,N_45202,N_45228);
xnor U45634 (N_45634,N_45321,N_45048);
xnor U45635 (N_45635,N_45065,N_45243);
and U45636 (N_45636,N_45344,N_45269);
xnor U45637 (N_45637,N_45166,N_45263);
or U45638 (N_45638,N_45399,N_45400);
and U45639 (N_45639,N_45099,N_45167);
nand U45640 (N_45640,N_45477,N_45440);
nor U45641 (N_45641,N_45256,N_45080);
or U45642 (N_45642,N_45300,N_45307);
xor U45643 (N_45643,N_45442,N_45281);
nand U45644 (N_45644,N_45422,N_45353);
nand U45645 (N_45645,N_45360,N_45181);
nor U45646 (N_45646,N_45412,N_45472);
xnor U45647 (N_45647,N_45009,N_45444);
xnor U45648 (N_45648,N_45028,N_45290);
nand U45649 (N_45649,N_45075,N_45438);
nor U45650 (N_45650,N_45078,N_45010);
xnor U45651 (N_45651,N_45373,N_45147);
or U45652 (N_45652,N_45324,N_45164);
nand U45653 (N_45653,N_45351,N_45121);
xnor U45654 (N_45654,N_45416,N_45032);
or U45655 (N_45655,N_45375,N_45441);
nand U45656 (N_45656,N_45248,N_45170);
nand U45657 (N_45657,N_45495,N_45363);
nor U45658 (N_45658,N_45137,N_45453);
xnor U45659 (N_45659,N_45459,N_45299);
nand U45660 (N_45660,N_45296,N_45059);
or U45661 (N_45661,N_45227,N_45410);
nand U45662 (N_45662,N_45473,N_45421);
or U45663 (N_45663,N_45328,N_45102);
or U45664 (N_45664,N_45047,N_45352);
and U45665 (N_45665,N_45447,N_45025);
xnor U45666 (N_45666,N_45205,N_45136);
or U45667 (N_45667,N_45234,N_45430);
nor U45668 (N_45668,N_45361,N_45337);
xnor U45669 (N_45669,N_45355,N_45483);
or U45670 (N_45670,N_45485,N_45378);
xnor U45671 (N_45671,N_45330,N_45003);
xor U45672 (N_45672,N_45304,N_45277);
nor U45673 (N_45673,N_45403,N_45470);
or U45674 (N_45674,N_45493,N_45383);
nand U45675 (N_45675,N_45180,N_45233);
nor U45676 (N_45676,N_45030,N_45329);
or U45677 (N_45677,N_45146,N_45499);
or U45678 (N_45678,N_45209,N_45023);
nor U45679 (N_45679,N_45100,N_45208);
and U45680 (N_45680,N_45478,N_45107);
and U45681 (N_45681,N_45276,N_45306);
xnor U45682 (N_45682,N_45371,N_45331);
nand U45683 (N_45683,N_45055,N_45370);
or U45684 (N_45684,N_45134,N_45487);
nor U45685 (N_45685,N_45387,N_45076);
and U45686 (N_45686,N_45112,N_45213);
or U45687 (N_45687,N_45395,N_45386);
or U45688 (N_45688,N_45230,N_45335);
or U45689 (N_45689,N_45448,N_45016);
or U45690 (N_45690,N_45156,N_45131);
or U45691 (N_45691,N_45468,N_45455);
or U45692 (N_45692,N_45044,N_45056);
nand U45693 (N_45693,N_45144,N_45366);
xor U45694 (N_45694,N_45187,N_45402);
nand U45695 (N_45695,N_45333,N_45007);
xor U45696 (N_45696,N_45348,N_45197);
xnor U45697 (N_45697,N_45462,N_45278);
nand U45698 (N_45698,N_45117,N_45103);
or U45699 (N_45699,N_45017,N_45206);
nand U45700 (N_45700,N_45408,N_45163);
nand U45701 (N_45701,N_45036,N_45251);
nand U45702 (N_45702,N_45491,N_45043);
xor U45703 (N_45703,N_45273,N_45095);
nand U45704 (N_45704,N_45279,N_45005);
or U45705 (N_45705,N_45292,N_45145);
xnor U45706 (N_45706,N_45133,N_45226);
or U45707 (N_45707,N_45111,N_45199);
xor U45708 (N_45708,N_45034,N_45088);
nor U45709 (N_45709,N_45338,N_45169);
or U45710 (N_45710,N_45326,N_45250);
or U45711 (N_45711,N_45096,N_45129);
or U45712 (N_45712,N_45280,N_45418);
and U45713 (N_45713,N_45481,N_45425);
and U45714 (N_45714,N_45153,N_45486);
nor U45715 (N_45715,N_45128,N_45270);
and U45716 (N_45716,N_45061,N_45042);
nor U45717 (N_45717,N_45027,N_45245);
or U45718 (N_45718,N_45031,N_45427);
and U45719 (N_45719,N_45069,N_45045);
xor U45720 (N_45720,N_45219,N_45359);
nand U45721 (N_45721,N_45018,N_45428);
and U45722 (N_45722,N_45374,N_45362);
nand U45723 (N_45723,N_45445,N_45143);
or U45724 (N_45724,N_45092,N_45159);
and U45725 (N_45725,N_45079,N_45174);
nor U45726 (N_45726,N_45040,N_45064);
or U45727 (N_45727,N_45063,N_45407);
or U45728 (N_45728,N_45390,N_45019);
and U45729 (N_45729,N_45262,N_45397);
or U45730 (N_45730,N_45274,N_45275);
nor U45731 (N_45731,N_45035,N_45068);
and U45732 (N_45732,N_45323,N_45325);
and U45733 (N_45733,N_45094,N_45004);
xor U45734 (N_45734,N_45271,N_45142);
and U45735 (N_45735,N_45372,N_45113);
xor U45736 (N_45736,N_45114,N_45264);
nor U45737 (N_45737,N_45312,N_45101);
and U45738 (N_45738,N_45149,N_45098);
or U45739 (N_45739,N_45458,N_45466);
nor U45740 (N_45740,N_45347,N_45089);
or U45741 (N_45741,N_45376,N_45284);
nand U45742 (N_45742,N_45350,N_45420);
or U45743 (N_45743,N_45413,N_45341);
nand U45744 (N_45744,N_45178,N_45160);
and U45745 (N_45745,N_45155,N_45115);
nand U45746 (N_45746,N_45001,N_45426);
nand U45747 (N_45747,N_45314,N_45419);
nor U45748 (N_45748,N_45119,N_45494);
nand U45749 (N_45749,N_45317,N_45189);
nor U45750 (N_45750,N_45025,N_45390);
or U45751 (N_45751,N_45283,N_45060);
nor U45752 (N_45752,N_45192,N_45078);
nor U45753 (N_45753,N_45272,N_45260);
nor U45754 (N_45754,N_45317,N_45241);
or U45755 (N_45755,N_45081,N_45092);
xnor U45756 (N_45756,N_45383,N_45291);
nand U45757 (N_45757,N_45348,N_45239);
xnor U45758 (N_45758,N_45288,N_45352);
or U45759 (N_45759,N_45366,N_45395);
or U45760 (N_45760,N_45242,N_45197);
xor U45761 (N_45761,N_45316,N_45457);
xnor U45762 (N_45762,N_45088,N_45208);
xor U45763 (N_45763,N_45011,N_45250);
and U45764 (N_45764,N_45017,N_45078);
nand U45765 (N_45765,N_45016,N_45131);
nor U45766 (N_45766,N_45337,N_45050);
and U45767 (N_45767,N_45046,N_45114);
and U45768 (N_45768,N_45402,N_45081);
nand U45769 (N_45769,N_45317,N_45338);
nand U45770 (N_45770,N_45288,N_45273);
and U45771 (N_45771,N_45441,N_45005);
xnor U45772 (N_45772,N_45113,N_45285);
nor U45773 (N_45773,N_45150,N_45233);
xnor U45774 (N_45774,N_45302,N_45444);
and U45775 (N_45775,N_45397,N_45494);
or U45776 (N_45776,N_45019,N_45306);
nor U45777 (N_45777,N_45362,N_45396);
and U45778 (N_45778,N_45279,N_45168);
xnor U45779 (N_45779,N_45106,N_45044);
xnor U45780 (N_45780,N_45225,N_45046);
and U45781 (N_45781,N_45237,N_45234);
and U45782 (N_45782,N_45128,N_45139);
xor U45783 (N_45783,N_45294,N_45176);
xnor U45784 (N_45784,N_45448,N_45286);
nor U45785 (N_45785,N_45386,N_45058);
nor U45786 (N_45786,N_45336,N_45226);
xor U45787 (N_45787,N_45071,N_45299);
xor U45788 (N_45788,N_45383,N_45410);
nor U45789 (N_45789,N_45004,N_45393);
or U45790 (N_45790,N_45251,N_45243);
xor U45791 (N_45791,N_45453,N_45310);
nand U45792 (N_45792,N_45321,N_45281);
or U45793 (N_45793,N_45423,N_45391);
nand U45794 (N_45794,N_45211,N_45183);
nand U45795 (N_45795,N_45433,N_45309);
or U45796 (N_45796,N_45228,N_45472);
nor U45797 (N_45797,N_45103,N_45374);
nor U45798 (N_45798,N_45071,N_45344);
and U45799 (N_45799,N_45219,N_45336);
and U45800 (N_45800,N_45152,N_45319);
and U45801 (N_45801,N_45209,N_45470);
and U45802 (N_45802,N_45416,N_45239);
nand U45803 (N_45803,N_45041,N_45300);
xnor U45804 (N_45804,N_45362,N_45223);
xnor U45805 (N_45805,N_45218,N_45085);
and U45806 (N_45806,N_45390,N_45091);
and U45807 (N_45807,N_45300,N_45208);
xnor U45808 (N_45808,N_45259,N_45019);
nand U45809 (N_45809,N_45217,N_45394);
nor U45810 (N_45810,N_45169,N_45127);
or U45811 (N_45811,N_45286,N_45354);
or U45812 (N_45812,N_45297,N_45012);
and U45813 (N_45813,N_45477,N_45076);
or U45814 (N_45814,N_45079,N_45228);
and U45815 (N_45815,N_45430,N_45034);
and U45816 (N_45816,N_45336,N_45263);
or U45817 (N_45817,N_45362,N_45105);
or U45818 (N_45818,N_45295,N_45000);
or U45819 (N_45819,N_45405,N_45040);
nand U45820 (N_45820,N_45127,N_45253);
nand U45821 (N_45821,N_45205,N_45381);
xnor U45822 (N_45822,N_45425,N_45164);
or U45823 (N_45823,N_45101,N_45195);
nand U45824 (N_45824,N_45152,N_45331);
nor U45825 (N_45825,N_45342,N_45236);
or U45826 (N_45826,N_45292,N_45147);
nor U45827 (N_45827,N_45422,N_45315);
xor U45828 (N_45828,N_45076,N_45470);
or U45829 (N_45829,N_45495,N_45055);
and U45830 (N_45830,N_45380,N_45494);
nor U45831 (N_45831,N_45395,N_45456);
xor U45832 (N_45832,N_45284,N_45193);
or U45833 (N_45833,N_45392,N_45328);
nand U45834 (N_45834,N_45440,N_45166);
and U45835 (N_45835,N_45188,N_45044);
nor U45836 (N_45836,N_45089,N_45290);
nand U45837 (N_45837,N_45114,N_45094);
nor U45838 (N_45838,N_45194,N_45473);
or U45839 (N_45839,N_45002,N_45386);
or U45840 (N_45840,N_45298,N_45330);
and U45841 (N_45841,N_45010,N_45303);
xnor U45842 (N_45842,N_45064,N_45340);
nor U45843 (N_45843,N_45303,N_45337);
xor U45844 (N_45844,N_45218,N_45110);
or U45845 (N_45845,N_45439,N_45418);
and U45846 (N_45846,N_45158,N_45411);
nand U45847 (N_45847,N_45191,N_45334);
or U45848 (N_45848,N_45196,N_45224);
xnor U45849 (N_45849,N_45018,N_45170);
or U45850 (N_45850,N_45475,N_45344);
xor U45851 (N_45851,N_45150,N_45230);
nor U45852 (N_45852,N_45085,N_45095);
or U45853 (N_45853,N_45164,N_45189);
and U45854 (N_45854,N_45363,N_45286);
or U45855 (N_45855,N_45273,N_45036);
nand U45856 (N_45856,N_45338,N_45303);
nand U45857 (N_45857,N_45157,N_45340);
and U45858 (N_45858,N_45115,N_45350);
nand U45859 (N_45859,N_45087,N_45071);
or U45860 (N_45860,N_45216,N_45366);
nor U45861 (N_45861,N_45015,N_45450);
nand U45862 (N_45862,N_45306,N_45437);
nor U45863 (N_45863,N_45000,N_45407);
nor U45864 (N_45864,N_45183,N_45303);
nor U45865 (N_45865,N_45243,N_45137);
nor U45866 (N_45866,N_45319,N_45313);
or U45867 (N_45867,N_45415,N_45103);
or U45868 (N_45868,N_45490,N_45410);
xnor U45869 (N_45869,N_45324,N_45418);
xnor U45870 (N_45870,N_45180,N_45171);
and U45871 (N_45871,N_45203,N_45349);
nor U45872 (N_45872,N_45384,N_45339);
xor U45873 (N_45873,N_45328,N_45455);
nor U45874 (N_45874,N_45329,N_45477);
or U45875 (N_45875,N_45266,N_45243);
or U45876 (N_45876,N_45223,N_45303);
and U45877 (N_45877,N_45187,N_45078);
nor U45878 (N_45878,N_45141,N_45020);
nand U45879 (N_45879,N_45470,N_45277);
nor U45880 (N_45880,N_45485,N_45090);
or U45881 (N_45881,N_45245,N_45208);
nand U45882 (N_45882,N_45086,N_45089);
or U45883 (N_45883,N_45401,N_45001);
nand U45884 (N_45884,N_45269,N_45347);
or U45885 (N_45885,N_45171,N_45078);
xnor U45886 (N_45886,N_45251,N_45268);
nor U45887 (N_45887,N_45130,N_45467);
nand U45888 (N_45888,N_45260,N_45047);
nand U45889 (N_45889,N_45176,N_45262);
nor U45890 (N_45890,N_45397,N_45498);
xor U45891 (N_45891,N_45303,N_45032);
or U45892 (N_45892,N_45084,N_45061);
or U45893 (N_45893,N_45223,N_45334);
and U45894 (N_45894,N_45091,N_45057);
or U45895 (N_45895,N_45469,N_45078);
xor U45896 (N_45896,N_45499,N_45184);
and U45897 (N_45897,N_45220,N_45424);
and U45898 (N_45898,N_45295,N_45357);
or U45899 (N_45899,N_45357,N_45060);
and U45900 (N_45900,N_45279,N_45098);
or U45901 (N_45901,N_45234,N_45301);
nor U45902 (N_45902,N_45305,N_45429);
and U45903 (N_45903,N_45194,N_45081);
and U45904 (N_45904,N_45331,N_45230);
or U45905 (N_45905,N_45211,N_45234);
xnor U45906 (N_45906,N_45148,N_45111);
xnor U45907 (N_45907,N_45201,N_45295);
xnor U45908 (N_45908,N_45181,N_45115);
or U45909 (N_45909,N_45391,N_45072);
and U45910 (N_45910,N_45478,N_45041);
nand U45911 (N_45911,N_45422,N_45383);
and U45912 (N_45912,N_45367,N_45201);
and U45913 (N_45913,N_45417,N_45242);
or U45914 (N_45914,N_45020,N_45321);
xnor U45915 (N_45915,N_45104,N_45082);
nand U45916 (N_45916,N_45232,N_45467);
xor U45917 (N_45917,N_45320,N_45252);
nand U45918 (N_45918,N_45155,N_45170);
or U45919 (N_45919,N_45212,N_45439);
and U45920 (N_45920,N_45024,N_45130);
xor U45921 (N_45921,N_45194,N_45333);
nand U45922 (N_45922,N_45393,N_45408);
nand U45923 (N_45923,N_45263,N_45315);
xnor U45924 (N_45924,N_45327,N_45409);
nor U45925 (N_45925,N_45012,N_45203);
and U45926 (N_45926,N_45229,N_45370);
nand U45927 (N_45927,N_45091,N_45055);
nand U45928 (N_45928,N_45184,N_45372);
nand U45929 (N_45929,N_45153,N_45052);
xor U45930 (N_45930,N_45380,N_45362);
or U45931 (N_45931,N_45148,N_45311);
and U45932 (N_45932,N_45441,N_45361);
or U45933 (N_45933,N_45034,N_45053);
nor U45934 (N_45934,N_45085,N_45488);
or U45935 (N_45935,N_45083,N_45001);
or U45936 (N_45936,N_45291,N_45130);
nor U45937 (N_45937,N_45380,N_45089);
or U45938 (N_45938,N_45433,N_45095);
nor U45939 (N_45939,N_45329,N_45057);
or U45940 (N_45940,N_45337,N_45043);
or U45941 (N_45941,N_45322,N_45215);
or U45942 (N_45942,N_45043,N_45436);
or U45943 (N_45943,N_45279,N_45127);
and U45944 (N_45944,N_45457,N_45372);
and U45945 (N_45945,N_45158,N_45187);
nor U45946 (N_45946,N_45065,N_45335);
nor U45947 (N_45947,N_45179,N_45012);
xnor U45948 (N_45948,N_45213,N_45368);
xnor U45949 (N_45949,N_45383,N_45034);
or U45950 (N_45950,N_45276,N_45030);
or U45951 (N_45951,N_45238,N_45413);
nand U45952 (N_45952,N_45280,N_45255);
nand U45953 (N_45953,N_45066,N_45460);
nand U45954 (N_45954,N_45362,N_45388);
xor U45955 (N_45955,N_45120,N_45057);
and U45956 (N_45956,N_45367,N_45373);
nor U45957 (N_45957,N_45456,N_45351);
nand U45958 (N_45958,N_45095,N_45043);
nand U45959 (N_45959,N_45293,N_45203);
nor U45960 (N_45960,N_45350,N_45326);
nand U45961 (N_45961,N_45121,N_45141);
xor U45962 (N_45962,N_45260,N_45296);
and U45963 (N_45963,N_45328,N_45055);
nand U45964 (N_45964,N_45381,N_45025);
nor U45965 (N_45965,N_45274,N_45224);
xor U45966 (N_45966,N_45161,N_45189);
nand U45967 (N_45967,N_45168,N_45114);
and U45968 (N_45968,N_45261,N_45025);
nor U45969 (N_45969,N_45159,N_45356);
or U45970 (N_45970,N_45466,N_45454);
nor U45971 (N_45971,N_45474,N_45081);
and U45972 (N_45972,N_45180,N_45358);
and U45973 (N_45973,N_45482,N_45249);
xor U45974 (N_45974,N_45384,N_45139);
or U45975 (N_45975,N_45325,N_45174);
and U45976 (N_45976,N_45405,N_45066);
nor U45977 (N_45977,N_45393,N_45337);
xnor U45978 (N_45978,N_45433,N_45219);
and U45979 (N_45979,N_45245,N_45248);
nor U45980 (N_45980,N_45254,N_45053);
nor U45981 (N_45981,N_45199,N_45008);
and U45982 (N_45982,N_45062,N_45394);
nor U45983 (N_45983,N_45366,N_45043);
and U45984 (N_45984,N_45258,N_45119);
nand U45985 (N_45985,N_45079,N_45493);
or U45986 (N_45986,N_45402,N_45279);
and U45987 (N_45987,N_45472,N_45259);
nor U45988 (N_45988,N_45379,N_45195);
or U45989 (N_45989,N_45408,N_45334);
xnor U45990 (N_45990,N_45381,N_45095);
and U45991 (N_45991,N_45328,N_45292);
xnor U45992 (N_45992,N_45039,N_45249);
and U45993 (N_45993,N_45419,N_45010);
xnor U45994 (N_45994,N_45359,N_45020);
or U45995 (N_45995,N_45456,N_45401);
xor U45996 (N_45996,N_45032,N_45112);
nand U45997 (N_45997,N_45257,N_45335);
and U45998 (N_45998,N_45342,N_45282);
nor U45999 (N_45999,N_45040,N_45045);
nand U46000 (N_46000,N_45865,N_45864);
nand U46001 (N_46001,N_45694,N_45666);
nor U46002 (N_46002,N_45586,N_45718);
or U46003 (N_46003,N_45761,N_45944);
and U46004 (N_46004,N_45716,N_45857);
xor U46005 (N_46005,N_45844,N_45560);
nand U46006 (N_46006,N_45536,N_45533);
and U46007 (N_46007,N_45519,N_45849);
or U46008 (N_46008,N_45960,N_45820);
xnor U46009 (N_46009,N_45649,N_45840);
nor U46010 (N_46010,N_45851,N_45791);
nor U46011 (N_46011,N_45850,N_45969);
or U46012 (N_46012,N_45826,N_45937);
or U46013 (N_46013,N_45633,N_45725);
nand U46014 (N_46014,N_45641,N_45590);
or U46015 (N_46015,N_45870,N_45819);
nand U46016 (N_46016,N_45654,N_45663);
or U46017 (N_46017,N_45572,N_45787);
nor U46018 (N_46018,N_45839,N_45735);
or U46019 (N_46019,N_45523,N_45550);
or U46020 (N_46020,N_45594,N_45794);
nand U46021 (N_46021,N_45945,N_45585);
and U46022 (N_46022,N_45778,N_45928);
nor U46023 (N_46023,N_45658,N_45577);
xnor U46024 (N_46024,N_45605,N_45738);
and U46025 (N_46025,N_45908,N_45650);
and U46026 (N_46026,N_45852,N_45990);
nand U46027 (N_46027,N_45797,N_45599);
nor U46028 (N_46028,N_45513,N_45744);
xnor U46029 (N_46029,N_45903,N_45770);
nand U46030 (N_46030,N_45991,N_45972);
nand U46031 (N_46031,N_45784,N_45900);
nand U46032 (N_46032,N_45950,N_45809);
and U46033 (N_46033,N_45561,N_45780);
nand U46034 (N_46034,N_45880,N_45795);
and U46035 (N_46035,N_45758,N_45509);
nand U46036 (N_46036,N_45668,N_45992);
xnor U46037 (N_46037,N_45606,N_45506);
nand U46038 (N_46038,N_45899,N_45811);
xor U46039 (N_46039,N_45996,N_45901);
xnor U46040 (N_46040,N_45861,N_45800);
or U46041 (N_46041,N_45918,N_45907);
nand U46042 (N_46042,N_45567,N_45734);
nand U46043 (N_46043,N_45845,N_45843);
or U46044 (N_46044,N_45573,N_45740);
nand U46045 (N_46045,N_45537,N_45952);
or U46046 (N_46046,N_45552,N_45763);
and U46047 (N_46047,N_45722,N_45648);
and U46048 (N_46048,N_45837,N_45730);
xnor U46049 (N_46049,N_45967,N_45879);
nand U46050 (N_46050,N_45833,N_45707);
xor U46051 (N_46051,N_45919,N_45984);
nand U46052 (N_46052,N_45531,N_45579);
xnor U46053 (N_46053,N_45555,N_45538);
xnor U46054 (N_46054,N_45557,N_45569);
xor U46055 (N_46055,N_45587,N_45875);
nand U46056 (N_46056,N_45604,N_45965);
and U46057 (N_46057,N_45540,N_45951);
xnor U46058 (N_46058,N_45546,N_45739);
xor U46059 (N_46059,N_45912,N_45817);
and U46060 (N_46060,N_45511,N_45822);
and U46061 (N_46061,N_45661,N_45553);
nor U46062 (N_46062,N_45893,N_45674);
and U46063 (N_46063,N_45691,N_45554);
and U46064 (N_46064,N_45924,N_45612);
or U46065 (N_46065,N_45772,N_45601);
xor U46066 (N_46066,N_45670,N_45510);
xnor U46067 (N_46067,N_45551,N_45799);
or U46068 (N_46068,N_45611,N_45878);
nor U46069 (N_46069,N_45673,N_45888);
nor U46070 (N_46070,N_45802,N_45524);
xor U46071 (N_46071,N_45986,N_45930);
and U46072 (N_46072,N_45793,N_45710);
and U46073 (N_46073,N_45836,N_45922);
nand U46074 (N_46074,N_45637,N_45999);
nor U46075 (N_46075,N_45915,N_45970);
and U46076 (N_46076,N_45618,N_45501);
or U46077 (N_46077,N_45774,N_45543);
nand U46078 (N_46078,N_45946,N_45568);
xnor U46079 (N_46079,N_45743,N_45589);
and U46080 (N_46080,N_45804,N_45995);
or U46081 (N_46081,N_45783,N_45655);
nor U46082 (N_46082,N_45731,N_45651);
nor U46083 (N_46083,N_45993,N_45838);
and U46084 (N_46084,N_45685,N_45887);
nor U46085 (N_46085,N_45798,N_45860);
or U46086 (N_46086,N_45942,N_45953);
and U46087 (N_46087,N_45853,N_45627);
xnor U46088 (N_46088,N_45571,N_45613);
or U46089 (N_46089,N_45520,N_45976);
nor U46090 (N_46090,N_45977,N_45749);
or U46091 (N_46091,N_45677,N_45834);
and U46092 (N_46092,N_45933,N_45830);
and U46093 (N_46093,N_45527,N_45898);
or U46094 (N_46094,N_45535,N_45994);
xnor U46095 (N_46095,N_45884,N_45848);
nor U46096 (N_46096,N_45588,N_45913);
and U46097 (N_46097,N_45626,N_45748);
xor U46098 (N_46098,N_45726,N_45812);
nor U46099 (N_46099,N_45701,N_45502);
nor U46100 (N_46100,N_45940,N_45989);
or U46101 (N_46101,N_45805,N_45667);
nand U46102 (N_46102,N_45751,N_45835);
nand U46103 (N_46103,N_45746,N_45790);
nor U46104 (N_46104,N_45635,N_45644);
xor U46105 (N_46105,N_45782,N_45760);
nor U46106 (N_46106,N_45825,N_45556);
or U46107 (N_46107,N_45925,N_45679);
or U46108 (N_46108,N_45862,N_45563);
or U46109 (N_46109,N_45905,N_45762);
nor U46110 (N_46110,N_45602,N_45607);
xor U46111 (N_46111,N_45621,N_45712);
nand U46112 (N_46112,N_45534,N_45959);
xnor U46113 (N_46113,N_45764,N_45926);
and U46114 (N_46114,N_45801,N_45842);
and U46115 (N_46115,N_45855,N_45831);
or U46116 (N_46116,N_45623,N_45957);
and U46117 (N_46117,N_45750,N_45985);
xnor U46118 (N_46118,N_45669,N_45688);
nand U46119 (N_46119,N_45935,N_45939);
or U46120 (N_46120,N_45700,N_45958);
nand U46121 (N_46121,N_45962,N_45954);
nor U46122 (N_46122,N_45732,N_45629);
nor U46123 (N_46123,N_45756,N_45948);
or U46124 (N_46124,N_45652,N_45828);
or U46125 (N_46125,N_45771,N_45631);
or U46126 (N_46126,N_45876,N_45708);
nand U46127 (N_46127,N_45891,N_45628);
and U46128 (N_46128,N_45600,N_45630);
or U46129 (N_46129,N_45622,N_45671);
or U46130 (N_46130,N_45776,N_45974);
nor U46131 (N_46131,N_45767,N_45578);
nand U46132 (N_46132,N_45582,N_45896);
and U46133 (N_46133,N_45659,N_45971);
or U46134 (N_46134,N_45709,N_45807);
xnor U46135 (N_46135,N_45541,N_45608);
xnor U46136 (N_46136,N_45752,N_45617);
or U46137 (N_46137,N_45856,N_45777);
xnor U46138 (N_46138,N_45868,N_45619);
and U46139 (N_46139,N_45681,N_45769);
nor U46140 (N_46140,N_45676,N_45934);
nand U46141 (N_46141,N_45713,N_45909);
and U46142 (N_46142,N_45757,N_45522);
nand U46143 (N_46143,N_45684,N_45727);
and U46144 (N_46144,N_45980,N_45558);
or U46145 (N_46145,N_45662,N_45955);
nand U46146 (N_46146,N_45664,N_45936);
nand U46147 (N_46147,N_45824,N_45785);
xnor U46148 (N_46148,N_45987,N_45645);
nand U46149 (N_46149,N_45847,N_45624);
or U46150 (N_46150,N_45647,N_45705);
and U46151 (N_46151,N_45720,N_45711);
nor U46152 (N_46152,N_45904,N_45689);
or U46153 (N_46153,N_45640,N_45877);
or U46154 (N_46154,N_45983,N_45963);
nand U46155 (N_46155,N_45885,N_45503);
nand U46156 (N_46156,N_45789,N_45759);
nand U46157 (N_46157,N_45997,N_45754);
and U46158 (N_46158,N_45547,N_45968);
nor U46159 (N_46159,N_45584,N_45598);
and U46160 (N_46160,N_45724,N_45636);
xnor U46161 (N_46161,N_45530,N_45686);
nand U46162 (N_46162,N_45981,N_45766);
or U46163 (N_46163,N_45656,N_45657);
xor U46164 (N_46164,N_45895,N_45927);
and U46165 (N_46165,N_45975,N_45719);
nand U46166 (N_46166,N_45693,N_45902);
xnor U46167 (N_46167,N_45779,N_45715);
xnor U46168 (N_46168,N_45765,N_45806);
xnor U46169 (N_46169,N_45564,N_45961);
or U46170 (N_46170,N_45886,N_45525);
xor U46171 (N_46171,N_45890,N_45717);
nand U46172 (N_46172,N_45603,N_45544);
nand U46173 (N_46173,N_45583,N_45949);
or U46174 (N_46174,N_45755,N_45858);
and U46175 (N_46175,N_45747,N_45516);
nor U46176 (N_46176,N_45575,N_45881);
and U46177 (N_46177,N_45803,N_45721);
and U46178 (N_46178,N_45775,N_45625);
and U46179 (N_46179,N_45595,N_45808);
xnor U46180 (N_46180,N_45643,N_45871);
or U46181 (N_46181,N_45742,N_45518);
xnor U46182 (N_46182,N_45515,N_45894);
and U46183 (N_46183,N_45580,N_45690);
and U46184 (N_46184,N_45592,N_45532);
or U46185 (N_46185,N_45781,N_45931);
nor U46186 (N_46186,N_45597,N_45832);
nor U46187 (N_46187,N_45660,N_45788);
and U46188 (N_46188,N_45545,N_45883);
or U46189 (N_46189,N_45702,N_45609);
nor U46190 (N_46190,N_45872,N_45892);
nand U46191 (N_46191,N_45815,N_45615);
nor U46192 (N_46192,N_45736,N_45910);
and U46193 (N_46193,N_45526,N_45576);
xnor U46194 (N_46194,N_45796,N_45818);
nor U46195 (N_46195,N_45562,N_45982);
xor U46196 (N_46196,N_45638,N_45911);
or U46197 (N_46197,N_45504,N_45917);
nor U46198 (N_46198,N_45508,N_45929);
nand U46199 (N_46199,N_45680,N_45528);
nor U46200 (N_46200,N_45753,N_45682);
and U46201 (N_46201,N_45813,N_45773);
or U46202 (N_46202,N_45559,N_45823);
xnor U46203 (N_46203,N_45706,N_45768);
xnor U46204 (N_46204,N_45548,N_45687);
and U46205 (N_46205,N_45646,N_45675);
nor U46206 (N_46206,N_45697,N_45846);
or U46207 (N_46207,N_45699,N_45723);
xnor U46208 (N_46208,N_45932,N_45867);
and U46209 (N_46209,N_45733,N_45632);
or U46210 (N_46210,N_45616,N_45916);
and U46211 (N_46211,N_45507,N_45639);
nor U46212 (N_46212,N_45897,N_45874);
or U46213 (N_46213,N_45728,N_45610);
or U46214 (N_46214,N_45542,N_45683);
xor U46215 (N_46215,N_45882,N_45914);
or U46216 (N_46216,N_45570,N_45653);
nor U46217 (N_46217,N_45696,N_45745);
nand U46218 (N_46218,N_45810,N_45786);
nand U46219 (N_46219,N_45678,N_45923);
nor U46220 (N_46220,N_45737,N_45873);
xor U46221 (N_46221,N_45591,N_45614);
or U46222 (N_46222,N_45729,N_45956);
nand U46223 (N_46223,N_45978,N_45964);
nand U46224 (N_46224,N_45889,N_45988);
nand U46225 (N_46225,N_45906,N_45549);
or U46226 (N_46226,N_45943,N_45500);
nor U46227 (N_46227,N_45539,N_45947);
xor U46228 (N_46228,N_45596,N_45869);
or U46229 (N_46229,N_45998,N_45938);
or U46230 (N_46230,N_45841,N_45816);
nor U46231 (N_46231,N_45517,N_45941);
xor U46232 (N_46232,N_45704,N_45966);
or U46233 (N_46233,N_45566,N_45829);
or U46234 (N_46234,N_45695,N_45593);
nor U46235 (N_46235,N_45692,N_45514);
xnor U46236 (N_46236,N_45505,N_45620);
xnor U46237 (N_46237,N_45921,N_45565);
xor U46238 (N_46238,N_45854,N_45512);
xnor U46239 (N_46239,N_45634,N_45863);
or U46240 (N_46240,N_45672,N_45665);
or U46241 (N_46241,N_45792,N_45521);
nor U46242 (N_46242,N_45703,N_45973);
or U46243 (N_46243,N_45741,N_45920);
or U46244 (N_46244,N_45866,N_45642);
xor U46245 (N_46245,N_45581,N_45714);
nor U46246 (N_46246,N_45979,N_45827);
and U46247 (N_46247,N_45814,N_45698);
nor U46248 (N_46248,N_45821,N_45859);
xnor U46249 (N_46249,N_45529,N_45574);
nand U46250 (N_46250,N_45717,N_45854);
and U46251 (N_46251,N_45687,N_45696);
xor U46252 (N_46252,N_45872,N_45657);
and U46253 (N_46253,N_45635,N_45720);
xor U46254 (N_46254,N_45813,N_45780);
nand U46255 (N_46255,N_45663,N_45664);
xnor U46256 (N_46256,N_45789,N_45772);
nor U46257 (N_46257,N_45715,N_45868);
or U46258 (N_46258,N_45983,N_45969);
and U46259 (N_46259,N_45716,N_45617);
xnor U46260 (N_46260,N_45683,N_45754);
nand U46261 (N_46261,N_45886,N_45600);
nand U46262 (N_46262,N_45686,N_45670);
nand U46263 (N_46263,N_45648,N_45893);
nor U46264 (N_46264,N_45650,N_45534);
nor U46265 (N_46265,N_45856,N_45828);
and U46266 (N_46266,N_45567,N_45851);
nor U46267 (N_46267,N_45644,N_45827);
nand U46268 (N_46268,N_45731,N_45594);
nand U46269 (N_46269,N_45704,N_45525);
nor U46270 (N_46270,N_45858,N_45642);
nor U46271 (N_46271,N_45989,N_45704);
nor U46272 (N_46272,N_45856,N_45867);
xor U46273 (N_46273,N_45656,N_45964);
xor U46274 (N_46274,N_45527,N_45813);
and U46275 (N_46275,N_45690,N_45812);
nor U46276 (N_46276,N_45648,N_45688);
nor U46277 (N_46277,N_45789,N_45509);
xor U46278 (N_46278,N_45728,N_45733);
nand U46279 (N_46279,N_45559,N_45539);
nor U46280 (N_46280,N_45923,N_45502);
or U46281 (N_46281,N_45523,N_45572);
or U46282 (N_46282,N_45553,N_45591);
xnor U46283 (N_46283,N_45823,N_45548);
nor U46284 (N_46284,N_45529,N_45843);
nand U46285 (N_46285,N_45891,N_45847);
and U46286 (N_46286,N_45567,N_45754);
nand U46287 (N_46287,N_45873,N_45755);
and U46288 (N_46288,N_45545,N_45532);
nand U46289 (N_46289,N_45863,N_45844);
xnor U46290 (N_46290,N_45722,N_45630);
and U46291 (N_46291,N_45723,N_45667);
nand U46292 (N_46292,N_45750,N_45872);
or U46293 (N_46293,N_45946,N_45897);
and U46294 (N_46294,N_45859,N_45548);
xor U46295 (N_46295,N_45785,N_45526);
nand U46296 (N_46296,N_45611,N_45882);
nor U46297 (N_46297,N_45766,N_45630);
nand U46298 (N_46298,N_45783,N_45757);
or U46299 (N_46299,N_45538,N_45826);
nor U46300 (N_46300,N_45952,N_45741);
nor U46301 (N_46301,N_45718,N_45931);
or U46302 (N_46302,N_45654,N_45676);
nand U46303 (N_46303,N_45858,N_45927);
and U46304 (N_46304,N_45547,N_45875);
and U46305 (N_46305,N_45823,N_45809);
nor U46306 (N_46306,N_45905,N_45679);
nor U46307 (N_46307,N_45798,N_45868);
and U46308 (N_46308,N_45770,N_45781);
or U46309 (N_46309,N_45686,N_45760);
nand U46310 (N_46310,N_45786,N_45672);
xnor U46311 (N_46311,N_45641,N_45562);
nor U46312 (N_46312,N_45860,N_45773);
nor U46313 (N_46313,N_45527,N_45731);
or U46314 (N_46314,N_45515,N_45547);
nand U46315 (N_46315,N_45855,N_45664);
or U46316 (N_46316,N_45766,N_45923);
and U46317 (N_46317,N_45685,N_45652);
or U46318 (N_46318,N_45734,N_45933);
xnor U46319 (N_46319,N_45748,N_45826);
nand U46320 (N_46320,N_45666,N_45884);
xor U46321 (N_46321,N_45889,N_45684);
nor U46322 (N_46322,N_45592,N_45777);
xor U46323 (N_46323,N_45511,N_45712);
xnor U46324 (N_46324,N_45574,N_45819);
xnor U46325 (N_46325,N_45894,N_45510);
or U46326 (N_46326,N_45691,N_45544);
or U46327 (N_46327,N_45644,N_45602);
nand U46328 (N_46328,N_45722,N_45803);
xnor U46329 (N_46329,N_45558,N_45718);
nand U46330 (N_46330,N_45539,N_45719);
nand U46331 (N_46331,N_45877,N_45573);
or U46332 (N_46332,N_45748,N_45554);
nand U46333 (N_46333,N_45850,N_45844);
nand U46334 (N_46334,N_45677,N_45752);
nor U46335 (N_46335,N_45617,N_45806);
nand U46336 (N_46336,N_45980,N_45632);
xnor U46337 (N_46337,N_45612,N_45770);
or U46338 (N_46338,N_45507,N_45809);
xnor U46339 (N_46339,N_45968,N_45702);
nand U46340 (N_46340,N_45701,N_45843);
nor U46341 (N_46341,N_45944,N_45956);
nand U46342 (N_46342,N_45976,N_45958);
and U46343 (N_46343,N_45954,N_45790);
xor U46344 (N_46344,N_45766,N_45700);
and U46345 (N_46345,N_45946,N_45704);
nand U46346 (N_46346,N_45654,N_45791);
and U46347 (N_46347,N_45639,N_45973);
and U46348 (N_46348,N_45621,N_45567);
xor U46349 (N_46349,N_45812,N_45710);
or U46350 (N_46350,N_45912,N_45539);
and U46351 (N_46351,N_45679,N_45667);
nand U46352 (N_46352,N_45863,N_45965);
or U46353 (N_46353,N_45638,N_45696);
nand U46354 (N_46354,N_45566,N_45890);
nand U46355 (N_46355,N_45695,N_45641);
nor U46356 (N_46356,N_45556,N_45798);
nor U46357 (N_46357,N_45813,N_45760);
nor U46358 (N_46358,N_45567,N_45684);
and U46359 (N_46359,N_45504,N_45563);
xor U46360 (N_46360,N_45627,N_45731);
and U46361 (N_46361,N_45791,N_45870);
nor U46362 (N_46362,N_45746,N_45706);
or U46363 (N_46363,N_45839,N_45612);
or U46364 (N_46364,N_45542,N_45629);
and U46365 (N_46365,N_45629,N_45706);
nand U46366 (N_46366,N_45664,N_45602);
nand U46367 (N_46367,N_45648,N_45854);
nor U46368 (N_46368,N_45745,N_45679);
or U46369 (N_46369,N_45940,N_45890);
nand U46370 (N_46370,N_45927,N_45691);
or U46371 (N_46371,N_45997,N_45704);
nor U46372 (N_46372,N_45545,N_45860);
xnor U46373 (N_46373,N_45600,N_45861);
nor U46374 (N_46374,N_45970,N_45743);
nor U46375 (N_46375,N_45668,N_45930);
nor U46376 (N_46376,N_45632,N_45580);
xnor U46377 (N_46377,N_45820,N_45524);
or U46378 (N_46378,N_45553,N_45572);
and U46379 (N_46379,N_45652,N_45671);
nand U46380 (N_46380,N_45705,N_45798);
xnor U46381 (N_46381,N_45939,N_45814);
xor U46382 (N_46382,N_45602,N_45974);
nand U46383 (N_46383,N_45677,N_45756);
and U46384 (N_46384,N_45716,N_45640);
xor U46385 (N_46385,N_45909,N_45915);
nand U46386 (N_46386,N_45903,N_45571);
and U46387 (N_46387,N_45501,N_45945);
nand U46388 (N_46388,N_45698,N_45518);
nand U46389 (N_46389,N_45666,N_45990);
xor U46390 (N_46390,N_45655,N_45940);
xor U46391 (N_46391,N_45698,N_45955);
xor U46392 (N_46392,N_45900,N_45724);
and U46393 (N_46393,N_45748,N_45906);
nor U46394 (N_46394,N_45887,N_45504);
or U46395 (N_46395,N_45913,N_45690);
nor U46396 (N_46396,N_45506,N_45602);
or U46397 (N_46397,N_45745,N_45639);
nor U46398 (N_46398,N_45521,N_45986);
xor U46399 (N_46399,N_45519,N_45922);
and U46400 (N_46400,N_45719,N_45948);
nand U46401 (N_46401,N_45896,N_45885);
nor U46402 (N_46402,N_45746,N_45521);
or U46403 (N_46403,N_45688,N_45760);
or U46404 (N_46404,N_45755,N_45733);
xor U46405 (N_46405,N_45725,N_45953);
or U46406 (N_46406,N_45626,N_45714);
xnor U46407 (N_46407,N_45667,N_45863);
nand U46408 (N_46408,N_45865,N_45737);
and U46409 (N_46409,N_45967,N_45669);
nor U46410 (N_46410,N_45873,N_45866);
or U46411 (N_46411,N_45790,N_45921);
or U46412 (N_46412,N_45610,N_45784);
nor U46413 (N_46413,N_45738,N_45551);
nand U46414 (N_46414,N_45787,N_45692);
and U46415 (N_46415,N_45594,N_45977);
nor U46416 (N_46416,N_45570,N_45878);
or U46417 (N_46417,N_45506,N_45537);
nand U46418 (N_46418,N_45586,N_45637);
xor U46419 (N_46419,N_45867,N_45780);
and U46420 (N_46420,N_45612,N_45677);
and U46421 (N_46421,N_45876,N_45889);
nor U46422 (N_46422,N_45964,N_45905);
nand U46423 (N_46423,N_45561,N_45619);
or U46424 (N_46424,N_45675,N_45752);
or U46425 (N_46425,N_45995,N_45731);
xor U46426 (N_46426,N_45792,N_45894);
and U46427 (N_46427,N_45718,N_45673);
nor U46428 (N_46428,N_45694,N_45652);
xor U46429 (N_46429,N_45926,N_45685);
and U46430 (N_46430,N_45696,N_45864);
or U46431 (N_46431,N_45729,N_45997);
nor U46432 (N_46432,N_45565,N_45800);
and U46433 (N_46433,N_45892,N_45524);
and U46434 (N_46434,N_45947,N_45730);
nand U46435 (N_46435,N_45539,N_45875);
nand U46436 (N_46436,N_45699,N_45525);
xor U46437 (N_46437,N_45874,N_45719);
nand U46438 (N_46438,N_45791,N_45533);
nor U46439 (N_46439,N_45931,N_45640);
or U46440 (N_46440,N_45845,N_45616);
nor U46441 (N_46441,N_45504,N_45704);
or U46442 (N_46442,N_45734,N_45594);
and U46443 (N_46443,N_45927,N_45870);
and U46444 (N_46444,N_45613,N_45729);
and U46445 (N_46445,N_45746,N_45600);
xnor U46446 (N_46446,N_45566,N_45962);
and U46447 (N_46447,N_45564,N_45884);
or U46448 (N_46448,N_45557,N_45516);
nand U46449 (N_46449,N_45785,N_45644);
nor U46450 (N_46450,N_45799,N_45985);
xor U46451 (N_46451,N_45842,N_45886);
nor U46452 (N_46452,N_45500,N_45982);
nor U46453 (N_46453,N_45512,N_45748);
nand U46454 (N_46454,N_45873,N_45910);
nand U46455 (N_46455,N_45680,N_45769);
or U46456 (N_46456,N_45730,N_45713);
xnor U46457 (N_46457,N_45712,N_45579);
nand U46458 (N_46458,N_45634,N_45797);
and U46459 (N_46459,N_45847,N_45835);
and U46460 (N_46460,N_45637,N_45691);
and U46461 (N_46461,N_45813,N_45832);
and U46462 (N_46462,N_45633,N_45761);
nor U46463 (N_46463,N_45716,N_45905);
and U46464 (N_46464,N_45956,N_45918);
nor U46465 (N_46465,N_45919,N_45724);
nor U46466 (N_46466,N_45825,N_45848);
or U46467 (N_46467,N_45702,N_45835);
nand U46468 (N_46468,N_45572,N_45845);
nor U46469 (N_46469,N_45765,N_45590);
nand U46470 (N_46470,N_45625,N_45771);
xnor U46471 (N_46471,N_45746,N_45823);
nor U46472 (N_46472,N_45580,N_45978);
or U46473 (N_46473,N_45734,N_45582);
nor U46474 (N_46474,N_45987,N_45691);
nand U46475 (N_46475,N_45910,N_45875);
or U46476 (N_46476,N_45931,N_45989);
xnor U46477 (N_46477,N_45945,N_45786);
or U46478 (N_46478,N_45609,N_45946);
and U46479 (N_46479,N_45576,N_45675);
or U46480 (N_46480,N_45701,N_45707);
nand U46481 (N_46481,N_45569,N_45885);
xor U46482 (N_46482,N_45829,N_45727);
and U46483 (N_46483,N_45728,N_45905);
xnor U46484 (N_46484,N_45876,N_45651);
or U46485 (N_46485,N_45560,N_45803);
or U46486 (N_46486,N_45908,N_45611);
nand U46487 (N_46487,N_45723,N_45965);
and U46488 (N_46488,N_45972,N_45831);
xnor U46489 (N_46489,N_45579,N_45707);
nor U46490 (N_46490,N_45938,N_45590);
xor U46491 (N_46491,N_45610,N_45997);
and U46492 (N_46492,N_45608,N_45762);
xnor U46493 (N_46493,N_45781,N_45663);
xnor U46494 (N_46494,N_45545,N_45887);
nand U46495 (N_46495,N_45642,N_45954);
and U46496 (N_46496,N_45669,N_45730);
nor U46497 (N_46497,N_45965,N_45984);
nor U46498 (N_46498,N_45620,N_45699);
and U46499 (N_46499,N_45573,N_45804);
nand U46500 (N_46500,N_46149,N_46473);
and U46501 (N_46501,N_46287,N_46437);
and U46502 (N_46502,N_46140,N_46071);
nand U46503 (N_46503,N_46023,N_46286);
xor U46504 (N_46504,N_46277,N_46192);
or U46505 (N_46505,N_46491,N_46032);
xor U46506 (N_46506,N_46103,N_46144);
nand U46507 (N_46507,N_46041,N_46090);
or U46508 (N_46508,N_46462,N_46400);
xor U46509 (N_46509,N_46415,N_46470);
nand U46510 (N_46510,N_46375,N_46463);
nand U46511 (N_46511,N_46214,N_46012);
nor U46512 (N_46512,N_46238,N_46379);
xor U46513 (N_46513,N_46497,N_46332);
nand U46514 (N_46514,N_46361,N_46031);
and U46515 (N_46515,N_46457,N_46407);
nand U46516 (N_46516,N_46424,N_46029);
nand U46517 (N_46517,N_46215,N_46194);
or U46518 (N_46518,N_46322,N_46363);
or U46519 (N_46519,N_46205,N_46364);
or U46520 (N_46520,N_46381,N_46256);
xor U46521 (N_46521,N_46005,N_46037);
nor U46522 (N_46522,N_46383,N_46271);
or U46523 (N_46523,N_46047,N_46116);
or U46524 (N_46524,N_46213,N_46311);
xnor U46525 (N_46525,N_46008,N_46137);
and U46526 (N_46526,N_46474,N_46303);
nand U46527 (N_46527,N_46265,N_46461);
and U46528 (N_46528,N_46024,N_46380);
or U46529 (N_46529,N_46232,N_46203);
and U46530 (N_46530,N_46298,N_46489);
nand U46531 (N_46531,N_46221,N_46083);
nand U46532 (N_46532,N_46114,N_46122);
nand U46533 (N_46533,N_46184,N_46081);
nor U46534 (N_46534,N_46016,N_46366);
and U46535 (N_46535,N_46398,N_46110);
nand U46536 (N_46536,N_46410,N_46347);
and U46537 (N_46537,N_46336,N_46312);
xnor U46538 (N_46538,N_46316,N_46393);
xnor U46539 (N_46539,N_46181,N_46360);
nor U46540 (N_46540,N_46422,N_46257);
and U46541 (N_46541,N_46058,N_46178);
xor U46542 (N_46542,N_46091,N_46406);
and U46543 (N_46543,N_46488,N_46163);
nand U46544 (N_46544,N_46076,N_46451);
xnor U46545 (N_46545,N_46241,N_46426);
or U46546 (N_46546,N_46469,N_46051);
and U46547 (N_46547,N_46447,N_46048);
nand U46548 (N_46548,N_46177,N_46479);
or U46549 (N_46549,N_46189,N_46401);
and U46550 (N_46550,N_46260,N_46471);
nand U46551 (N_46551,N_46409,N_46352);
xnor U46552 (N_46552,N_46066,N_46267);
and U46553 (N_46553,N_46057,N_46227);
nor U46554 (N_46554,N_46362,N_46456);
or U46555 (N_46555,N_46446,N_46033);
xor U46556 (N_46556,N_46390,N_46295);
xor U46557 (N_46557,N_46340,N_46281);
xnor U46558 (N_46558,N_46039,N_46236);
nand U46559 (N_46559,N_46392,N_46134);
nand U46560 (N_46560,N_46145,N_46301);
nor U46561 (N_46561,N_46204,N_46297);
nand U46562 (N_46562,N_46154,N_46142);
nor U46563 (N_46563,N_46234,N_46218);
and U46564 (N_46564,N_46208,N_46111);
or U46565 (N_46565,N_46018,N_46272);
nor U46566 (N_46566,N_46370,N_46198);
nand U46567 (N_46567,N_46388,N_46419);
nor U46568 (N_46568,N_46460,N_46143);
and U46569 (N_46569,N_46342,N_46280);
and U46570 (N_46570,N_46093,N_46268);
or U46571 (N_46571,N_46269,N_46499);
nand U46572 (N_46572,N_46433,N_46112);
xnor U46573 (N_46573,N_46458,N_46070);
nand U46574 (N_46574,N_46243,N_46180);
or U46575 (N_46575,N_46317,N_46060);
nand U46576 (N_46576,N_46250,N_46262);
nand U46577 (N_46577,N_46167,N_46124);
or U46578 (N_46578,N_46273,N_46357);
nand U46579 (N_46579,N_46050,N_46129);
xnor U46580 (N_46580,N_46490,N_46325);
xor U46581 (N_46581,N_46020,N_46373);
nand U46582 (N_46582,N_46484,N_46173);
nand U46583 (N_46583,N_46067,N_46284);
or U46584 (N_46584,N_46450,N_46323);
and U46585 (N_46585,N_46464,N_46334);
xnor U46586 (N_46586,N_46305,N_46126);
xor U46587 (N_46587,N_46132,N_46085);
or U46588 (N_46588,N_46389,N_46444);
and U46589 (N_46589,N_46061,N_46367);
nand U46590 (N_46590,N_46319,N_46349);
nor U46591 (N_46591,N_46130,N_46086);
nor U46592 (N_46592,N_46369,N_46026);
nand U46593 (N_46593,N_46010,N_46141);
xnor U46594 (N_46594,N_46127,N_46007);
and U46595 (N_46595,N_46448,N_46442);
or U46596 (N_46596,N_46465,N_46397);
nor U46597 (N_46597,N_46359,N_46219);
xnor U46598 (N_46598,N_46413,N_46339);
xor U46599 (N_46599,N_46171,N_46253);
nand U46600 (N_46600,N_46368,N_46493);
nand U46601 (N_46601,N_46139,N_46434);
and U46602 (N_46602,N_46344,N_46074);
or U46603 (N_46603,N_46087,N_46259);
or U46604 (N_46604,N_46231,N_46102);
or U46605 (N_46605,N_46396,N_46237);
nor U46606 (N_46606,N_46147,N_46372);
and U46607 (N_46607,N_46411,N_46377);
or U46608 (N_46608,N_46046,N_46402);
or U46609 (N_46609,N_46306,N_46172);
or U46610 (N_46610,N_46498,N_46261);
xnor U46611 (N_46611,N_46240,N_46414);
xnor U46612 (N_46612,N_46439,N_46248);
xnor U46613 (N_46613,N_46329,N_46350);
xor U46614 (N_46614,N_46391,N_46109);
and U46615 (N_46615,N_46436,N_46107);
nand U46616 (N_46616,N_46356,N_46435);
nand U46617 (N_46617,N_46251,N_46068);
and U46618 (N_46618,N_46151,N_46254);
or U46619 (N_46619,N_46176,N_46244);
nand U46620 (N_46620,N_46408,N_46331);
xor U46621 (N_46621,N_46345,N_46494);
xnor U46622 (N_46622,N_46003,N_46064);
xor U46623 (N_46623,N_46378,N_46072);
nor U46624 (N_46624,N_46202,N_46292);
or U46625 (N_46625,N_46477,N_46476);
and U46626 (N_46626,N_46220,N_46001);
xor U46627 (N_46627,N_46043,N_46291);
nand U46628 (N_46628,N_46233,N_46376);
xnor U46629 (N_46629,N_46210,N_46123);
nand U46630 (N_46630,N_46247,N_46193);
and U46631 (N_46631,N_46054,N_46338);
and U46632 (N_46632,N_46166,N_46092);
or U46633 (N_46633,N_46496,N_46153);
or U46634 (N_46634,N_46159,N_46084);
nand U46635 (N_46635,N_46483,N_46217);
and U46636 (N_46636,N_46453,N_46096);
and U46637 (N_46637,N_46445,N_46190);
nor U46638 (N_46638,N_46274,N_46438);
nor U46639 (N_46639,N_46335,N_46307);
nor U46640 (N_46640,N_46098,N_46075);
and U46641 (N_46641,N_46175,N_46384);
nor U46642 (N_46642,N_46069,N_46044);
nand U46643 (N_46643,N_46455,N_46387);
nand U46644 (N_46644,N_46431,N_46355);
nand U46645 (N_46645,N_46206,N_46080);
xnor U46646 (N_46646,N_46374,N_46150);
nand U46647 (N_46647,N_46089,N_46017);
nand U46648 (N_46648,N_46118,N_46136);
nor U46649 (N_46649,N_46152,N_46191);
nor U46650 (N_46650,N_46160,N_46099);
and U46651 (N_46651,N_46412,N_46027);
nand U46652 (N_46652,N_46117,N_46314);
nand U46653 (N_46653,N_46354,N_46289);
xnor U46654 (N_46654,N_46276,N_46346);
nand U46655 (N_46655,N_46014,N_46252);
and U46656 (N_46656,N_46418,N_46207);
xnor U46657 (N_46657,N_46042,N_46337);
xor U46658 (N_46658,N_46482,N_46417);
xor U46659 (N_46659,N_46258,N_46293);
or U46660 (N_46660,N_46230,N_46266);
or U46661 (N_46661,N_46187,N_46224);
and U46662 (N_46662,N_46146,N_46164);
nor U46663 (N_46663,N_46326,N_46330);
nand U46664 (N_46664,N_46310,N_46475);
or U46665 (N_46665,N_46290,N_46053);
and U46666 (N_46666,N_46157,N_46030);
nand U46667 (N_46667,N_46282,N_46135);
or U46668 (N_46668,N_46382,N_46056);
and U46669 (N_46669,N_46327,N_46495);
and U46670 (N_46670,N_46432,N_46263);
xnor U46671 (N_46671,N_46034,N_46430);
or U46672 (N_46672,N_46300,N_46480);
nand U46673 (N_46673,N_46104,N_46079);
nor U46674 (N_46674,N_46222,N_46094);
xor U46675 (N_46675,N_46052,N_46025);
xor U46676 (N_46676,N_46201,N_46425);
nor U46677 (N_46677,N_46420,N_46158);
nand U46678 (N_46678,N_46371,N_46000);
xnor U46679 (N_46679,N_46385,N_46040);
and U46680 (N_46680,N_46321,N_46299);
nand U46681 (N_46681,N_46013,N_46004);
nor U46682 (N_46682,N_46162,N_46120);
or U46683 (N_46683,N_46270,N_46125);
and U46684 (N_46684,N_46174,N_46492);
nand U46685 (N_46685,N_46097,N_46416);
and U46686 (N_46686,N_46228,N_46128);
and U46687 (N_46687,N_46341,N_46468);
nor U46688 (N_46688,N_46138,N_46195);
nor U46689 (N_46689,N_46285,N_46440);
or U46690 (N_46690,N_46036,N_46421);
nor U46691 (N_46691,N_46186,N_46015);
xor U46692 (N_46692,N_46199,N_46200);
xnor U46693 (N_46693,N_46182,N_46133);
xor U46694 (N_46694,N_46188,N_46035);
or U46695 (N_46695,N_46478,N_46324);
xor U46696 (N_46696,N_46209,N_46165);
nand U46697 (N_46697,N_46454,N_46423);
and U46698 (N_46698,N_46155,N_46427);
nand U46699 (N_46699,N_46358,N_46055);
xor U46700 (N_46700,N_46038,N_46021);
or U46701 (N_46701,N_46100,N_46296);
and U46702 (N_46702,N_46333,N_46131);
or U46703 (N_46703,N_46119,N_46028);
or U46704 (N_46704,N_46313,N_46386);
nand U46705 (N_46705,N_46169,N_46156);
nor U46706 (N_46706,N_46487,N_46077);
and U46707 (N_46707,N_46179,N_46328);
and U46708 (N_46708,N_46467,N_46062);
nor U46709 (N_46709,N_46148,N_46403);
nor U46710 (N_46710,N_46108,N_46459);
or U46711 (N_46711,N_46429,N_46065);
nor U46712 (N_46712,N_46019,N_46170);
nand U46713 (N_46713,N_46002,N_46315);
and U46714 (N_46714,N_46318,N_46404);
or U46715 (N_46715,N_46365,N_46353);
xnor U46716 (N_46716,N_46168,N_46229);
or U46717 (N_46717,N_46045,N_46095);
nand U46718 (N_46718,N_46278,N_46308);
or U46719 (N_46719,N_46405,N_46009);
or U46720 (N_46720,N_46082,N_46394);
nand U46721 (N_46721,N_46049,N_46283);
nand U46722 (N_46722,N_46105,N_46216);
xor U46723 (N_46723,N_46279,N_46226);
nand U46724 (N_46724,N_46275,N_46245);
xor U46725 (N_46725,N_46294,N_46212);
nand U46726 (N_46726,N_46255,N_46288);
or U46727 (N_46727,N_46343,N_46428);
nor U46728 (N_46728,N_46101,N_46239);
or U46729 (N_46729,N_46242,N_46223);
nand U46730 (N_46730,N_46106,N_46351);
and U46731 (N_46731,N_46196,N_46481);
xor U46732 (N_46732,N_46115,N_46264);
and U46733 (N_46733,N_46249,N_46235);
nor U46734 (N_46734,N_46183,N_46161);
nor U46735 (N_46735,N_46466,N_46399);
nor U46736 (N_46736,N_46320,N_46011);
or U46737 (N_46737,N_46211,N_46449);
nor U46738 (N_46738,N_46309,N_46485);
xnor U46739 (N_46739,N_46063,N_46059);
nor U46740 (N_46740,N_46246,N_46486);
nor U46741 (N_46741,N_46006,N_46078);
nand U46742 (N_46742,N_46395,N_46348);
nand U46743 (N_46743,N_46472,N_46073);
and U46744 (N_46744,N_46185,N_46441);
and U46745 (N_46745,N_46452,N_46022);
nand U46746 (N_46746,N_46225,N_46302);
nand U46747 (N_46747,N_46088,N_46304);
or U46748 (N_46748,N_46113,N_46443);
nand U46749 (N_46749,N_46121,N_46197);
or U46750 (N_46750,N_46101,N_46387);
nand U46751 (N_46751,N_46075,N_46392);
and U46752 (N_46752,N_46027,N_46006);
or U46753 (N_46753,N_46256,N_46124);
nand U46754 (N_46754,N_46410,N_46069);
nor U46755 (N_46755,N_46069,N_46462);
nor U46756 (N_46756,N_46366,N_46359);
nand U46757 (N_46757,N_46179,N_46308);
and U46758 (N_46758,N_46453,N_46072);
nand U46759 (N_46759,N_46020,N_46028);
or U46760 (N_46760,N_46259,N_46188);
nor U46761 (N_46761,N_46420,N_46173);
nor U46762 (N_46762,N_46434,N_46219);
or U46763 (N_46763,N_46137,N_46234);
xor U46764 (N_46764,N_46132,N_46004);
nor U46765 (N_46765,N_46205,N_46410);
and U46766 (N_46766,N_46405,N_46052);
or U46767 (N_46767,N_46343,N_46478);
nor U46768 (N_46768,N_46323,N_46011);
nor U46769 (N_46769,N_46413,N_46477);
nand U46770 (N_46770,N_46403,N_46109);
xnor U46771 (N_46771,N_46447,N_46109);
or U46772 (N_46772,N_46320,N_46003);
xnor U46773 (N_46773,N_46404,N_46359);
nor U46774 (N_46774,N_46222,N_46297);
or U46775 (N_46775,N_46304,N_46071);
or U46776 (N_46776,N_46235,N_46495);
or U46777 (N_46777,N_46271,N_46379);
nand U46778 (N_46778,N_46124,N_46376);
xnor U46779 (N_46779,N_46380,N_46177);
xnor U46780 (N_46780,N_46348,N_46407);
or U46781 (N_46781,N_46105,N_46025);
nand U46782 (N_46782,N_46168,N_46019);
nand U46783 (N_46783,N_46255,N_46055);
xor U46784 (N_46784,N_46156,N_46455);
or U46785 (N_46785,N_46010,N_46388);
and U46786 (N_46786,N_46103,N_46009);
and U46787 (N_46787,N_46301,N_46047);
and U46788 (N_46788,N_46113,N_46404);
or U46789 (N_46789,N_46152,N_46197);
or U46790 (N_46790,N_46012,N_46455);
nor U46791 (N_46791,N_46061,N_46452);
nand U46792 (N_46792,N_46407,N_46405);
or U46793 (N_46793,N_46275,N_46427);
xor U46794 (N_46794,N_46100,N_46499);
xor U46795 (N_46795,N_46096,N_46308);
nor U46796 (N_46796,N_46138,N_46499);
xor U46797 (N_46797,N_46270,N_46015);
nand U46798 (N_46798,N_46054,N_46198);
xor U46799 (N_46799,N_46121,N_46389);
xnor U46800 (N_46800,N_46186,N_46056);
nand U46801 (N_46801,N_46224,N_46394);
nor U46802 (N_46802,N_46460,N_46230);
and U46803 (N_46803,N_46096,N_46215);
nor U46804 (N_46804,N_46319,N_46217);
nand U46805 (N_46805,N_46440,N_46389);
and U46806 (N_46806,N_46034,N_46314);
xnor U46807 (N_46807,N_46400,N_46309);
nand U46808 (N_46808,N_46228,N_46313);
nand U46809 (N_46809,N_46027,N_46214);
and U46810 (N_46810,N_46453,N_46225);
and U46811 (N_46811,N_46348,N_46356);
and U46812 (N_46812,N_46218,N_46193);
nand U46813 (N_46813,N_46418,N_46192);
and U46814 (N_46814,N_46353,N_46116);
nor U46815 (N_46815,N_46174,N_46496);
xnor U46816 (N_46816,N_46107,N_46473);
or U46817 (N_46817,N_46237,N_46418);
xnor U46818 (N_46818,N_46302,N_46278);
xnor U46819 (N_46819,N_46272,N_46020);
nor U46820 (N_46820,N_46233,N_46498);
nand U46821 (N_46821,N_46000,N_46189);
or U46822 (N_46822,N_46196,N_46453);
or U46823 (N_46823,N_46295,N_46149);
xnor U46824 (N_46824,N_46426,N_46450);
xor U46825 (N_46825,N_46133,N_46304);
xor U46826 (N_46826,N_46210,N_46088);
nor U46827 (N_46827,N_46375,N_46071);
nand U46828 (N_46828,N_46071,N_46012);
xnor U46829 (N_46829,N_46192,N_46311);
and U46830 (N_46830,N_46048,N_46297);
and U46831 (N_46831,N_46166,N_46366);
and U46832 (N_46832,N_46216,N_46027);
nand U46833 (N_46833,N_46241,N_46167);
xnor U46834 (N_46834,N_46443,N_46350);
or U46835 (N_46835,N_46006,N_46335);
nor U46836 (N_46836,N_46449,N_46024);
xor U46837 (N_46837,N_46356,N_46189);
nand U46838 (N_46838,N_46061,N_46417);
xor U46839 (N_46839,N_46164,N_46258);
nor U46840 (N_46840,N_46410,N_46046);
or U46841 (N_46841,N_46265,N_46356);
and U46842 (N_46842,N_46491,N_46384);
nand U46843 (N_46843,N_46040,N_46490);
nor U46844 (N_46844,N_46253,N_46234);
or U46845 (N_46845,N_46429,N_46381);
nor U46846 (N_46846,N_46430,N_46334);
or U46847 (N_46847,N_46124,N_46189);
nand U46848 (N_46848,N_46379,N_46106);
and U46849 (N_46849,N_46355,N_46277);
or U46850 (N_46850,N_46264,N_46141);
and U46851 (N_46851,N_46360,N_46452);
nand U46852 (N_46852,N_46131,N_46197);
xor U46853 (N_46853,N_46311,N_46416);
nand U46854 (N_46854,N_46479,N_46324);
xor U46855 (N_46855,N_46188,N_46449);
or U46856 (N_46856,N_46232,N_46428);
or U46857 (N_46857,N_46297,N_46076);
and U46858 (N_46858,N_46448,N_46476);
or U46859 (N_46859,N_46224,N_46167);
or U46860 (N_46860,N_46488,N_46155);
and U46861 (N_46861,N_46116,N_46338);
or U46862 (N_46862,N_46125,N_46341);
nand U46863 (N_46863,N_46039,N_46442);
nor U46864 (N_46864,N_46391,N_46142);
and U46865 (N_46865,N_46411,N_46128);
nand U46866 (N_46866,N_46048,N_46287);
xor U46867 (N_46867,N_46437,N_46181);
nor U46868 (N_46868,N_46136,N_46437);
nor U46869 (N_46869,N_46416,N_46295);
or U46870 (N_46870,N_46245,N_46026);
or U46871 (N_46871,N_46412,N_46052);
or U46872 (N_46872,N_46331,N_46263);
and U46873 (N_46873,N_46121,N_46117);
or U46874 (N_46874,N_46128,N_46032);
nand U46875 (N_46875,N_46106,N_46171);
or U46876 (N_46876,N_46149,N_46021);
or U46877 (N_46877,N_46261,N_46004);
or U46878 (N_46878,N_46354,N_46200);
and U46879 (N_46879,N_46106,N_46490);
xnor U46880 (N_46880,N_46371,N_46428);
nand U46881 (N_46881,N_46237,N_46273);
nor U46882 (N_46882,N_46442,N_46166);
nor U46883 (N_46883,N_46359,N_46346);
nor U46884 (N_46884,N_46409,N_46289);
and U46885 (N_46885,N_46280,N_46111);
nor U46886 (N_46886,N_46002,N_46401);
nor U46887 (N_46887,N_46157,N_46266);
nand U46888 (N_46888,N_46253,N_46369);
and U46889 (N_46889,N_46034,N_46291);
nand U46890 (N_46890,N_46088,N_46004);
nor U46891 (N_46891,N_46247,N_46015);
xnor U46892 (N_46892,N_46207,N_46299);
xnor U46893 (N_46893,N_46019,N_46422);
nor U46894 (N_46894,N_46411,N_46442);
or U46895 (N_46895,N_46115,N_46127);
and U46896 (N_46896,N_46047,N_46239);
or U46897 (N_46897,N_46280,N_46269);
or U46898 (N_46898,N_46018,N_46261);
nor U46899 (N_46899,N_46068,N_46430);
nand U46900 (N_46900,N_46179,N_46288);
xnor U46901 (N_46901,N_46391,N_46464);
or U46902 (N_46902,N_46411,N_46253);
nand U46903 (N_46903,N_46405,N_46161);
and U46904 (N_46904,N_46168,N_46001);
or U46905 (N_46905,N_46334,N_46009);
nand U46906 (N_46906,N_46190,N_46433);
nor U46907 (N_46907,N_46223,N_46339);
and U46908 (N_46908,N_46185,N_46258);
or U46909 (N_46909,N_46289,N_46197);
nor U46910 (N_46910,N_46112,N_46279);
nor U46911 (N_46911,N_46121,N_46105);
or U46912 (N_46912,N_46078,N_46051);
xor U46913 (N_46913,N_46339,N_46009);
nand U46914 (N_46914,N_46309,N_46464);
nand U46915 (N_46915,N_46233,N_46074);
and U46916 (N_46916,N_46479,N_46451);
nor U46917 (N_46917,N_46271,N_46441);
or U46918 (N_46918,N_46489,N_46413);
and U46919 (N_46919,N_46170,N_46244);
and U46920 (N_46920,N_46377,N_46446);
nor U46921 (N_46921,N_46347,N_46254);
or U46922 (N_46922,N_46429,N_46173);
nand U46923 (N_46923,N_46231,N_46495);
and U46924 (N_46924,N_46183,N_46187);
nor U46925 (N_46925,N_46356,N_46331);
and U46926 (N_46926,N_46133,N_46121);
nor U46927 (N_46927,N_46485,N_46130);
and U46928 (N_46928,N_46229,N_46075);
nor U46929 (N_46929,N_46314,N_46289);
or U46930 (N_46930,N_46191,N_46397);
nand U46931 (N_46931,N_46109,N_46382);
nor U46932 (N_46932,N_46402,N_46193);
nor U46933 (N_46933,N_46085,N_46093);
nand U46934 (N_46934,N_46402,N_46435);
nand U46935 (N_46935,N_46012,N_46361);
or U46936 (N_46936,N_46349,N_46100);
or U46937 (N_46937,N_46425,N_46154);
or U46938 (N_46938,N_46482,N_46393);
and U46939 (N_46939,N_46458,N_46114);
nor U46940 (N_46940,N_46326,N_46081);
nor U46941 (N_46941,N_46004,N_46089);
nor U46942 (N_46942,N_46102,N_46386);
nor U46943 (N_46943,N_46123,N_46449);
nand U46944 (N_46944,N_46205,N_46407);
xnor U46945 (N_46945,N_46317,N_46407);
xnor U46946 (N_46946,N_46061,N_46344);
xnor U46947 (N_46947,N_46095,N_46245);
and U46948 (N_46948,N_46074,N_46105);
nand U46949 (N_46949,N_46364,N_46152);
xor U46950 (N_46950,N_46099,N_46198);
xnor U46951 (N_46951,N_46054,N_46127);
and U46952 (N_46952,N_46192,N_46322);
nand U46953 (N_46953,N_46378,N_46394);
nor U46954 (N_46954,N_46016,N_46368);
xnor U46955 (N_46955,N_46326,N_46333);
nand U46956 (N_46956,N_46194,N_46292);
nor U46957 (N_46957,N_46470,N_46268);
nor U46958 (N_46958,N_46349,N_46175);
nand U46959 (N_46959,N_46453,N_46274);
or U46960 (N_46960,N_46217,N_46445);
nor U46961 (N_46961,N_46243,N_46205);
nor U46962 (N_46962,N_46269,N_46425);
nand U46963 (N_46963,N_46037,N_46014);
and U46964 (N_46964,N_46414,N_46073);
or U46965 (N_46965,N_46308,N_46145);
nand U46966 (N_46966,N_46097,N_46028);
and U46967 (N_46967,N_46222,N_46025);
xor U46968 (N_46968,N_46100,N_46186);
or U46969 (N_46969,N_46301,N_46374);
xnor U46970 (N_46970,N_46479,N_46003);
and U46971 (N_46971,N_46202,N_46354);
xnor U46972 (N_46972,N_46014,N_46234);
nand U46973 (N_46973,N_46338,N_46115);
xor U46974 (N_46974,N_46454,N_46434);
nand U46975 (N_46975,N_46102,N_46262);
or U46976 (N_46976,N_46054,N_46479);
or U46977 (N_46977,N_46079,N_46230);
xnor U46978 (N_46978,N_46329,N_46098);
nand U46979 (N_46979,N_46083,N_46089);
and U46980 (N_46980,N_46142,N_46147);
nor U46981 (N_46981,N_46471,N_46484);
or U46982 (N_46982,N_46350,N_46148);
nand U46983 (N_46983,N_46045,N_46055);
and U46984 (N_46984,N_46481,N_46151);
nand U46985 (N_46985,N_46403,N_46402);
or U46986 (N_46986,N_46396,N_46385);
xor U46987 (N_46987,N_46268,N_46486);
and U46988 (N_46988,N_46150,N_46258);
or U46989 (N_46989,N_46452,N_46384);
nand U46990 (N_46990,N_46155,N_46390);
and U46991 (N_46991,N_46363,N_46240);
nor U46992 (N_46992,N_46270,N_46353);
xor U46993 (N_46993,N_46452,N_46252);
and U46994 (N_46994,N_46464,N_46112);
xor U46995 (N_46995,N_46134,N_46376);
and U46996 (N_46996,N_46249,N_46370);
or U46997 (N_46997,N_46128,N_46043);
nor U46998 (N_46998,N_46030,N_46411);
xor U46999 (N_46999,N_46259,N_46313);
nand U47000 (N_47000,N_46667,N_46818);
nor U47001 (N_47001,N_46586,N_46599);
and U47002 (N_47002,N_46585,N_46921);
and U47003 (N_47003,N_46775,N_46502);
or U47004 (N_47004,N_46985,N_46773);
nand U47005 (N_47005,N_46992,N_46843);
and U47006 (N_47006,N_46969,N_46834);
xor U47007 (N_47007,N_46870,N_46763);
xor U47008 (N_47008,N_46690,N_46875);
and U47009 (N_47009,N_46766,N_46751);
nor U47010 (N_47010,N_46906,N_46953);
or U47011 (N_47011,N_46967,N_46642);
nor U47012 (N_47012,N_46598,N_46643);
and U47013 (N_47013,N_46744,N_46680);
and U47014 (N_47014,N_46511,N_46539);
nand U47015 (N_47015,N_46804,N_46943);
and U47016 (N_47016,N_46646,N_46639);
or U47017 (N_47017,N_46644,N_46855);
xor U47018 (N_47018,N_46674,N_46576);
and U47019 (N_47019,N_46512,N_46662);
nand U47020 (N_47020,N_46507,N_46964);
nor U47021 (N_47021,N_46799,N_46900);
or U47022 (N_47022,N_46946,N_46737);
and U47023 (N_47023,N_46790,N_46853);
nand U47024 (N_47024,N_46968,N_46919);
nor U47025 (N_47025,N_46890,N_46983);
nand U47026 (N_47026,N_46738,N_46877);
and U47027 (N_47027,N_46679,N_46572);
xnor U47028 (N_47028,N_46669,N_46987);
xnor U47029 (N_47029,N_46889,N_46725);
xor U47030 (N_47030,N_46620,N_46527);
nand U47031 (N_47031,N_46811,N_46610);
and U47032 (N_47032,N_46709,N_46924);
or U47033 (N_47033,N_46684,N_46581);
and U47034 (N_47034,N_46794,N_46791);
xor U47035 (N_47035,N_46508,N_46869);
or U47036 (N_47036,N_46827,N_46768);
or U47037 (N_47037,N_46503,N_46606);
nand U47038 (N_47038,N_46863,N_46991);
or U47039 (N_47039,N_46640,N_46857);
nand U47040 (N_47040,N_46626,N_46904);
nor U47041 (N_47041,N_46721,N_46526);
nor U47042 (N_47042,N_46665,N_46808);
or U47043 (N_47043,N_46696,N_46578);
nor U47044 (N_47044,N_46510,N_46828);
and U47045 (N_47045,N_46830,N_46530);
and U47046 (N_47046,N_46745,N_46687);
and U47047 (N_47047,N_46936,N_46755);
nor U47048 (N_47048,N_46541,N_46705);
and U47049 (N_47049,N_46899,N_46786);
and U47050 (N_47050,N_46901,N_46603);
and U47051 (N_47051,N_46734,N_46742);
nor U47052 (N_47052,N_46522,N_46501);
or U47053 (N_47053,N_46693,N_46762);
or U47054 (N_47054,N_46575,N_46944);
or U47055 (N_47055,N_46874,N_46926);
nand U47056 (N_47056,N_46951,N_46880);
nor U47057 (N_47057,N_46698,N_46653);
xnor U47058 (N_47058,N_46878,N_46938);
or U47059 (N_47059,N_46883,N_46868);
nand U47060 (N_47060,N_46905,N_46701);
nand U47061 (N_47061,N_46947,N_46935);
or U47062 (N_47062,N_46810,N_46723);
nand U47063 (N_47063,N_46892,N_46859);
and U47064 (N_47064,N_46956,N_46556);
nand U47065 (N_47065,N_46689,N_46547);
nand U47066 (N_47066,N_46776,N_46706);
xnor U47067 (N_47067,N_46993,N_46633);
and U47068 (N_47068,N_46712,N_46719);
or U47069 (N_47069,N_46702,N_46990);
and U47070 (N_47070,N_46845,N_46873);
or U47071 (N_47071,N_46931,N_46858);
nor U47072 (N_47072,N_46849,N_46523);
nor U47073 (N_47073,N_46722,N_46909);
xor U47074 (N_47074,N_46675,N_46937);
nand U47075 (N_47075,N_46865,N_46817);
nand U47076 (N_47076,N_46695,N_46761);
or U47077 (N_47077,N_46846,N_46566);
nand U47078 (N_47078,N_46941,N_46772);
and U47079 (N_47079,N_46895,N_46717);
and U47080 (N_47080,N_46715,N_46797);
and U47081 (N_47081,N_46513,N_46713);
xnor U47082 (N_47082,N_46589,N_46559);
and U47083 (N_47083,N_46622,N_46929);
nand U47084 (N_47084,N_46882,N_46793);
nor U47085 (N_47085,N_46978,N_46739);
and U47086 (N_47086,N_46542,N_46861);
nor U47087 (N_47087,N_46822,N_46902);
xnor U47088 (N_47088,N_46917,N_46749);
xnor U47089 (N_47089,N_46995,N_46914);
and U47090 (N_47090,N_46879,N_46652);
nor U47091 (N_47091,N_46650,N_46664);
nand U47092 (N_47092,N_46688,N_46597);
or U47093 (N_47093,N_46796,N_46996);
and U47094 (N_47094,N_46711,N_46989);
xnor U47095 (N_47095,N_46960,N_46984);
nor U47096 (N_47096,N_46618,N_46694);
or U47097 (N_47097,N_46886,N_46505);
and U47098 (N_47098,N_46979,N_46959);
xnor U47099 (N_47099,N_46641,N_46515);
and U47100 (N_47100,N_46638,N_46560);
and U47101 (N_47101,N_46631,N_46747);
and U47102 (N_47102,N_46840,N_46866);
and U47103 (N_47103,N_46893,N_46668);
nand U47104 (N_47104,N_46833,N_46700);
or U47105 (N_47105,N_46608,N_46624);
nand U47106 (N_47106,N_46757,N_46837);
xor U47107 (N_47107,N_46660,N_46795);
or U47108 (N_47108,N_46927,N_46699);
nor U47109 (N_47109,N_46881,N_46970);
nand U47110 (N_47110,N_46732,N_46820);
nor U47111 (N_47111,N_46814,N_46545);
nor U47112 (N_47112,N_46821,N_46832);
nand U47113 (N_47113,N_46649,N_46752);
xor U47114 (N_47114,N_46982,N_46816);
nand U47115 (N_47115,N_46678,N_46933);
and U47116 (N_47116,N_46587,N_46677);
or U47117 (N_47117,N_46916,N_46600);
or U47118 (N_47118,N_46731,N_46850);
nor U47119 (N_47119,N_46656,N_46577);
nand U47120 (N_47120,N_46518,N_46525);
nor U47121 (N_47121,N_46555,N_46798);
xnor U47122 (N_47122,N_46623,N_46676);
xnor U47123 (N_47123,N_46976,N_46912);
nor U47124 (N_47124,N_46546,N_46609);
or U47125 (N_47125,N_46844,N_46614);
nand U47126 (N_47126,N_46683,N_46841);
and U47127 (N_47127,N_46686,N_46565);
and U47128 (N_47128,N_46852,N_46704);
and U47129 (N_47129,N_46788,N_46862);
and U47130 (N_47130,N_46682,N_46787);
nor U47131 (N_47131,N_46955,N_46531);
and U47132 (N_47132,N_46888,N_46672);
or U47133 (N_47133,N_46898,N_46860);
and U47134 (N_47134,N_46645,N_46663);
or U47135 (N_47135,N_46519,N_46973);
nand U47136 (N_47136,N_46703,N_46544);
and U47137 (N_47137,N_46537,N_46911);
xor U47138 (N_47138,N_46602,N_46753);
xnor U47139 (N_47139,N_46651,N_46500);
nand U47140 (N_47140,N_46908,N_46948);
nor U47141 (N_47141,N_46759,N_46961);
and U47142 (N_47142,N_46553,N_46552);
nand U47143 (N_47143,N_46764,N_46897);
nor U47144 (N_47144,N_46940,N_46743);
nor U47145 (N_47145,N_46774,N_46517);
xnor U47146 (N_47146,N_46750,N_46819);
nor U47147 (N_47147,N_46516,N_46885);
or U47148 (N_47148,N_46997,N_46634);
and U47149 (N_47149,N_46627,N_46681);
nand U47150 (N_47150,N_46864,N_46907);
nand U47151 (N_47151,N_46685,N_46671);
and U47152 (N_47152,N_46872,N_46661);
nor U47153 (N_47153,N_46708,N_46925);
nor U47154 (N_47154,N_46584,N_46760);
or U47155 (N_47155,N_46957,N_46839);
nor U47156 (N_47156,N_46632,N_46966);
or U47157 (N_47157,N_46746,N_46616);
nand U47158 (N_47158,N_46601,N_46777);
or U47159 (N_47159,N_46724,N_46758);
nand U47160 (N_47160,N_46812,N_46806);
and U47161 (N_47161,N_46570,N_46654);
and U47162 (N_47162,N_46548,N_46971);
nor U47163 (N_47163,N_46952,N_46736);
or U47164 (N_47164,N_46965,N_46949);
nor U47165 (N_47165,N_46692,N_46670);
or U47166 (N_47166,N_46856,N_46784);
xnor U47167 (N_47167,N_46536,N_46592);
nand U47168 (N_47168,N_46612,N_46563);
nand U47169 (N_47169,N_46781,N_46574);
nand U47170 (N_47170,N_46615,N_46756);
nor U47171 (N_47171,N_46807,N_46792);
xnor U47172 (N_47172,N_46923,N_46915);
or U47173 (N_47173,N_46504,N_46520);
or U47174 (N_47174,N_46625,N_46826);
and U47175 (N_47175,N_46876,N_46999);
or U47176 (N_47176,N_46932,N_46802);
nand U47177 (N_47177,N_46735,N_46564);
and U47178 (N_47178,N_46655,N_46697);
and U47179 (N_47179,N_46887,N_46836);
nor U47180 (N_47180,N_46729,N_46958);
or U47181 (N_47181,N_46803,N_46783);
nand U47182 (N_47182,N_46628,N_46588);
xor U47183 (N_47183,N_46621,N_46558);
nor U47184 (N_47184,N_46557,N_46707);
nand U47185 (N_47185,N_46580,N_46673);
xor U47186 (N_47186,N_46934,N_46813);
and U47187 (N_47187,N_46854,N_46535);
xnor U47188 (N_47188,N_46521,N_46613);
nand U47189 (N_47189,N_46720,N_46963);
xor U47190 (N_47190,N_46789,N_46824);
or U47191 (N_47191,N_46590,N_46630);
nand U47192 (N_47192,N_46962,N_46851);
and U47193 (N_47193,N_46842,N_46569);
or U47194 (N_47194,N_46972,N_46939);
nand U47195 (N_47195,N_46691,N_46551);
nand U47196 (N_47196,N_46910,N_46740);
and U47197 (N_47197,N_46771,N_46727);
xor U47198 (N_47198,N_46835,N_46884);
and U47199 (N_47199,N_46894,N_46891);
nand U47200 (N_47200,N_46604,N_46617);
nor U47201 (N_47201,N_46954,N_46658);
nand U47202 (N_47202,N_46831,N_46710);
nand U47203 (N_47203,N_46847,N_46533);
nor U47204 (N_47204,N_46648,N_46550);
xor U47205 (N_47205,N_46805,N_46778);
xnor U47206 (N_47206,N_46896,N_46605);
and U47207 (N_47207,N_46619,N_46611);
or U47208 (N_47208,N_46568,N_46540);
and U47209 (N_47209,N_46593,N_46524);
xnor U47210 (N_47210,N_46629,N_46657);
nor U47211 (N_47211,N_46986,N_46918);
or U47212 (N_47212,N_46591,N_46977);
or U47213 (N_47213,N_46922,N_46636);
xnor U47214 (N_47214,N_46748,N_46903);
xor U47215 (N_47215,N_46514,N_46928);
nor U47216 (N_47216,N_46782,N_46543);
nand U47217 (N_47217,N_46561,N_46779);
nand U47218 (N_47218,N_46998,N_46838);
and U47219 (N_47219,N_46871,N_46981);
nor U47220 (N_47220,N_46988,N_46980);
and U47221 (N_47221,N_46741,N_46809);
and U47222 (N_47222,N_46974,N_46538);
xnor U47223 (N_47223,N_46765,N_46770);
nand U47224 (N_47224,N_46714,N_46637);
nand U47225 (N_47225,N_46607,N_46801);
xor U47226 (N_47226,N_46594,N_46567);
xnor U47227 (N_47227,N_46945,N_46529);
or U47228 (N_47228,N_46554,N_46635);
or U47229 (N_47229,N_46848,N_46728);
xor U47230 (N_47230,N_46579,N_46754);
xor U47231 (N_47231,N_46930,N_46920);
or U47232 (N_47232,N_46942,N_46730);
and U47233 (N_47233,N_46780,N_46647);
or U47234 (N_47234,N_46562,N_46583);
xnor U47235 (N_47235,N_46596,N_46829);
xnor U47236 (N_47236,N_46785,N_46825);
or U47237 (N_47237,N_46528,N_46815);
xor U47238 (N_47238,N_46994,N_46716);
and U47239 (N_47239,N_46769,N_46823);
nand U47240 (N_47240,N_46509,N_46867);
nor U47241 (N_47241,N_46718,N_46532);
nor U47242 (N_47242,N_46573,N_46733);
xnor U47243 (N_47243,N_46595,N_46666);
nand U47244 (N_47244,N_46726,N_46913);
xnor U47245 (N_47245,N_46800,N_46975);
nor U47246 (N_47246,N_46534,N_46950);
xnor U47247 (N_47247,N_46582,N_46549);
nand U47248 (N_47248,N_46506,N_46767);
nand U47249 (N_47249,N_46571,N_46659);
nand U47250 (N_47250,N_46927,N_46977);
or U47251 (N_47251,N_46840,N_46514);
or U47252 (N_47252,N_46953,N_46698);
and U47253 (N_47253,N_46507,N_46549);
xor U47254 (N_47254,N_46565,N_46532);
xnor U47255 (N_47255,N_46526,N_46792);
nor U47256 (N_47256,N_46672,N_46807);
and U47257 (N_47257,N_46774,N_46756);
or U47258 (N_47258,N_46981,N_46992);
nand U47259 (N_47259,N_46903,N_46701);
and U47260 (N_47260,N_46747,N_46717);
or U47261 (N_47261,N_46854,N_46985);
or U47262 (N_47262,N_46816,N_46877);
nand U47263 (N_47263,N_46580,N_46657);
nor U47264 (N_47264,N_46765,N_46971);
nor U47265 (N_47265,N_46851,N_46655);
nor U47266 (N_47266,N_46521,N_46638);
nor U47267 (N_47267,N_46578,N_46626);
and U47268 (N_47268,N_46795,N_46644);
nand U47269 (N_47269,N_46835,N_46975);
nand U47270 (N_47270,N_46544,N_46964);
nand U47271 (N_47271,N_46595,N_46653);
nor U47272 (N_47272,N_46530,N_46619);
xnor U47273 (N_47273,N_46753,N_46601);
or U47274 (N_47274,N_46879,N_46782);
and U47275 (N_47275,N_46684,N_46953);
nor U47276 (N_47276,N_46843,N_46747);
nand U47277 (N_47277,N_46919,N_46728);
nand U47278 (N_47278,N_46799,N_46758);
or U47279 (N_47279,N_46684,N_46984);
nand U47280 (N_47280,N_46945,N_46911);
xnor U47281 (N_47281,N_46932,N_46759);
or U47282 (N_47282,N_46978,N_46641);
and U47283 (N_47283,N_46523,N_46589);
nor U47284 (N_47284,N_46719,N_46627);
nor U47285 (N_47285,N_46950,N_46597);
nor U47286 (N_47286,N_46646,N_46609);
and U47287 (N_47287,N_46681,N_46647);
or U47288 (N_47288,N_46777,N_46523);
nor U47289 (N_47289,N_46707,N_46978);
xnor U47290 (N_47290,N_46604,N_46500);
nor U47291 (N_47291,N_46926,N_46596);
or U47292 (N_47292,N_46653,N_46849);
and U47293 (N_47293,N_46622,N_46519);
and U47294 (N_47294,N_46526,N_46672);
and U47295 (N_47295,N_46749,N_46632);
xnor U47296 (N_47296,N_46562,N_46845);
nor U47297 (N_47297,N_46713,N_46569);
nand U47298 (N_47298,N_46925,N_46573);
nor U47299 (N_47299,N_46704,N_46605);
nor U47300 (N_47300,N_46915,N_46714);
nand U47301 (N_47301,N_46728,N_46591);
xor U47302 (N_47302,N_46861,N_46956);
nor U47303 (N_47303,N_46730,N_46533);
or U47304 (N_47304,N_46856,N_46916);
or U47305 (N_47305,N_46951,N_46583);
xor U47306 (N_47306,N_46697,N_46877);
xor U47307 (N_47307,N_46962,N_46889);
nor U47308 (N_47308,N_46739,N_46917);
and U47309 (N_47309,N_46959,N_46944);
xor U47310 (N_47310,N_46729,N_46748);
or U47311 (N_47311,N_46736,N_46903);
and U47312 (N_47312,N_46626,N_46833);
nor U47313 (N_47313,N_46550,N_46775);
or U47314 (N_47314,N_46534,N_46750);
or U47315 (N_47315,N_46512,N_46766);
nand U47316 (N_47316,N_46806,N_46784);
or U47317 (N_47317,N_46738,N_46653);
xor U47318 (N_47318,N_46827,N_46599);
and U47319 (N_47319,N_46617,N_46705);
and U47320 (N_47320,N_46515,N_46933);
and U47321 (N_47321,N_46550,N_46656);
or U47322 (N_47322,N_46565,N_46994);
nor U47323 (N_47323,N_46638,N_46831);
and U47324 (N_47324,N_46992,N_46849);
or U47325 (N_47325,N_46961,N_46691);
and U47326 (N_47326,N_46890,N_46529);
and U47327 (N_47327,N_46832,N_46838);
and U47328 (N_47328,N_46848,N_46900);
or U47329 (N_47329,N_46952,N_46748);
or U47330 (N_47330,N_46693,N_46665);
xor U47331 (N_47331,N_46926,N_46839);
or U47332 (N_47332,N_46512,N_46840);
or U47333 (N_47333,N_46617,N_46615);
and U47334 (N_47334,N_46982,N_46645);
or U47335 (N_47335,N_46691,N_46771);
nor U47336 (N_47336,N_46625,N_46664);
nor U47337 (N_47337,N_46944,N_46698);
nor U47338 (N_47338,N_46794,N_46801);
xnor U47339 (N_47339,N_46613,N_46792);
nor U47340 (N_47340,N_46635,N_46773);
xor U47341 (N_47341,N_46737,N_46967);
nand U47342 (N_47342,N_46904,N_46987);
and U47343 (N_47343,N_46595,N_46737);
nor U47344 (N_47344,N_46751,N_46698);
xor U47345 (N_47345,N_46891,N_46890);
and U47346 (N_47346,N_46987,N_46716);
nor U47347 (N_47347,N_46964,N_46638);
or U47348 (N_47348,N_46614,N_46966);
and U47349 (N_47349,N_46921,N_46792);
nand U47350 (N_47350,N_46784,N_46588);
nor U47351 (N_47351,N_46562,N_46714);
nand U47352 (N_47352,N_46891,N_46615);
and U47353 (N_47353,N_46584,N_46504);
nand U47354 (N_47354,N_46609,N_46749);
or U47355 (N_47355,N_46901,N_46816);
nand U47356 (N_47356,N_46827,N_46794);
nor U47357 (N_47357,N_46759,N_46663);
nand U47358 (N_47358,N_46591,N_46527);
xnor U47359 (N_47359,N_46907,N_46500);
nor U47360 (N_47360,N_46779,N_46862);
and U47361 (N_47361,N_46869,N_46927);
nor U47362 (N_47362,N_46521,N_46515);
or U47363 (N_47363,N_46654,N_46673);
or U47364 (N_47364,N_46558,N_46683);
nor U47365 (N_47365,N_46685,N_46716);
xor U47366 (N_47366,N_46749,N_46715);
nand U47367 (N_47367,N_46520,N_46900);
xnor U47368 (N_47368,N_46853,N_46924);
xor U47369 (N_47369,N_46857,N_46585);
or U47370 (N_47370,N_46911,N_46704);
nand U47371 (N_47371,N_46623,N_46772);
or U47372 (N_47372,N_46830,N_46996);
and U47373 (N_47373,N_46839,N_46694);
xnor U47374 (N_47374,N_46657,N_46805);
or U47375 (N_47375,N_46755,N_46686);
nor U47376 (N_47376,N_46523,N_46678);
and U47377 (N_47377,N_46538,N_46809);
xnor U47378 (N_47378,N_46922,N_46529);
and U47379 (N_47379,N_46889,N_46903);
xnor U47380 (N_47380,N_46647,N_46700);
and U47381 (N_47381,N_46992,N_46502);
nand U47382 (N_47382,N_46801,N_46637);
or U47383 (N_47383,N_46972,N_46599);
xor U47384 (N_47384,N_46735,N_46755);
or U47385 (N_47385,N_46916,N_46662);
and U47386 (N_47386,N_46605,N_46905);
nor U47387 (N_47387,N_46690,N_46646);
nor U47388 (N_47388,N_46536,N_46691);
xor U47389 (N_47389,N_46859,N_46692);
xor U47390 (N_47390,N_46793,N_46825);
nand U47391 (N_47391,N_46634,N_46573);
and U47392 (N_47392,N_46657,N_46614);
nand U47393 (N_47393,N_46685,N_46818);
nor U47394 (N_47394,N_46780,N_46627);
nand U47395 (N_47395,N_46827,N_46979);
or U47396 (N_47396,N_46793,N_46839);
nand U47397 (N_47397,N_46595,N_46734);
xnor U47398 (N_47398,N_46759,N_46805);
nor U47399 (N_47399,N_46541,N_46647);
nor U47400 (N_47400,N_46536,N_46544);
xnor U47401 (N_47401,N_46812,N_46745);
or U47402 (N_47402,N_46768,N_46666);
nor U47403 (N_47403,N_46956,N_46578);
nand U47404 (N_47404,N_46592,N_46983);
or U47405 (N_47405,N_46927,N_46503);
and U47406 (N_47406,N_46876,N_46890);
nand U47407 (N_47407,N_46998,N_46763);
nand U47408 (N_47408,N_46783,N_46721);
nor U47409 (N_47409,N_46882,N_46795);
nor U47410 (N_47410,N_46647,N_46512);
nor U47411 (N_47411,N_46583,N_46804);
nor U47412 (N_47412,N_46797,N_46887);
nand U47413 (N_47413,N_46921,N_46687);
or U47414 (N_47414,N_46618,N_46926);
or U47415 (N_47415,N_46843,N_46738);
xnor U47416 (N_47416,N_46901,N_46584);
and U47417 (N_47417,N_46697,N_46695);
nor U47418 (N_47418,N_46935,N_46929);
nand U47419 (N_47419,N_46570,N_46567);
nor U47420 (N_47420,N_46599,N_46886);
nor U47421 (N_47421,N_46511,N_46831);
xor U47422 (N_47422,N_46673,N_46696);
nand U47423 (N_47423,N_46875,N_46545);
or U47424 (N_47424,N_46689,N_46803);
nand U47425 (N_47425,N_46636,N_46677);
nand U47426 (N_47426,N_46542,N_46739);
xnor U47427 (N_47427,N_46636,N_46535);
nor U47428 (N_47428,N_46998,N_46902);
nand U47429 (N_47429,N_46916,N_46771);
or U47430 (N_47430,N_46963,N_46941);
nor U47431 (N_47431,N_46790,N_46919);
and U47432 (N_47432,N_46612,N_46674);
nor U47433 (N_47433,N_46926,N_46551);
nor U47434 (N_47434,N_46707,N_46942);
nand U47435 (N_47435,N_46758,N_46631);
and U47436 (N_47436,N_46849,N_46777);
nor U47437 (N_47437,N_46893,N_46538);
and U47438 (N_47438,N_46723,N_46511);
and U47439 (N_47439,N_46643,N_46774);
or U47440 (N_47440,N_46897,N_46549);
nand U47441 (N_47441,N_46766,N_46678);
or U47442 (N_47442,N_46906,N_46624);
xnor U47443 (N_47443,N_46622,N_46712);
nor U47444 (N_47444,N_46867,N_46857);
or U47445 (N_47445,N_46851,N_46951);
nor U47446 (N_47446,N_46758,N_46625);
or U47447 (N_47447,N_46869,N_46767);
nor U47448 (N_47448,N_46727,N_46556);
or U47449 (N_47449,N_46743,N_46790);
nand U47450 (N_47450,N_46668,N_46707);
and U47451 (N_47451,N_46516,N_46556);
xnor U47452 (N_47452,N_46872,N_46607);
or U47453 (N_47453,N_46902,N_46698);
or U47454 (N_47454,N_46614,N_46520);
nand U47455 (N_47455,N_46803,N_46811);
or U47456 (N_47456,N_46725,N_46520);
nand U47457 (N_47457,N_46784,N_46611);
xnor U47458 (N_47458,N_46837,N_46632);
or U47459 (N_47459,N_46764,N_46573);
nor U47460 (N_47460,N_46529,N_46990);
nor U47461 (N_47461,N_46606,N_46790);
and U47462 (N_47462,N_46708,N_46835);
nor U47463 (N_47463,N_46593,N_46709);
xor U47464 (N_47464,N_46543,N_46875);
or U47465 (N_47465,N_46555,N_46596);
and U47466 (N_47466,N_46791,N_46608);
and U47467 (N_47467,N_46576,N_46967);
xnor U47468 (N_47468,N_46970,N_46710);
and U47469 (N_47469,N_46981,N_46679);
and U47470 (N_47470,N_46955,N_46681);
xnor U47471 (N_47471,N_46787,N_46560);
nand U47472 (N_47472,N_46964,N_46671);
nand U47473 (N_47473,N_46827,N_46822);
xnor U47474 (N_47474,N_46875,N_46801);
nand U47475 (N_47475,N_46745,N_46688);
nor U47476 (N_47476,N_46737,N_46887);
nand U47477 (N_47477,N_46578,N_46661);
or U47478 (N_47478,N_46952,N_46719);
and U47479 (N_47479,N_46692,N_46866);
or U47480 (N_47480,N_46692,N_46643);
xor U47481 (N_47481,N_46612,N_46532);
nand U47482 (N_47482,N_46755,N_46913);
and U47483 (N_47483,N_46619,N_46967);
xor U47484 (N_47484,N_46543,N_46704);
or U47485 (N_47485,N_46627,N_46561);
nor U47486 (N_47486,N_46608,N_46893);
or U47487 (N_47487,N_46624,N_46692);
and U47488 (N_47488,N_46640,N_46513);
nand U47489 (N_47489,N_46570,N_46802);
nor U47490 (N_47490,N_46776,N_46993);
and U47491 (N_47491,N_46596,N_46589);
nor U47492 (N_47492,N_46963,N_46596);
xnor U47493 (N_47493,N_46930,N_46988);
nand U47494 (N_47494,N_46694,N_46905);
or U47495 (N_47495,N_46536,N_46950);
xnor U47496 (N_47496,N_46843,N_46857);
or U47497 (N_47497,N_46548,N_46561);
and U47498 (N_47498,N_46595,N_46920);
nand U47499 (N_47499,N_46548,N_46786);
or U47500 (N_47500,N_47039,N_47125);
or U47501 (N_47501,N_47095,N_47460);
and U47502 (N_47502,N_47214,N_47316);
and U47503 (N_47503,N_47185,N_47149);
xor U47504 (N_47504,N_47428,N_47348);
nand U47505 (N_47505,N_47181,N_47263);
and U47506 (N_47506,N_47400,N_47497);
nand U47507 (N_47507,N_47123,N_47220);
nor U47508 (N_47508,N_47137,N_47006);
xnor U47509 (N_47509,N_47332,N_47398);
or U47510 (N_47510,N_47441,N_47446);
and U47511 (N_47511,N_47242,N_47094);
and U47512 (N_47512,N_47075,N_47250);
nor U47513 (N_47513,N_47043,N_47223);
nand U47514 (N_47514,N_47403,N_47231);
xnor U47515 (N_47515,N_47319,N_47432);
and U47516 (N_47516,N_47292,N_47443);
nand U47517 (N_47517,N_47329,N_47227);
and U47518 (N_47518,N_47254,N_47297);
and U47519 (N_47519,N_47208,N_47176);
or U47520 (N_47520,N_47007,N_47311);
or U47521 (N_47521,N_47114,N_47093);
xor U47522 (N_47522,N_47005,N_47057);
nand U47523 (N_47523,N_47483,N_47140);
nor U47524 (N_47524,N_47285,N_47042);
nor U47525 (N_47525,N_47045,N_47028);
or U47526 (N_47526,N_47378,N_47030);
and U47527 (N_47527,N_47325,N_47321);
xor U47528 (N_47528,N_47022,N_47182);
nand U47529 (N_47529,N_47178,N_47277);
or U47530 (N_47530,N_47296,N_47097);
or U47531 (N_47531,N_47156,N_47146);
nor U47532 (N_47532,N_47308,N_47420);
nor U47533 (N_47533,N_47422,N_47035);
nor U47534 (N_47534,N_47279,N_47433);
xor U47535 (N_47535,N_47496,N_47239);
and U47536 (N_47536,N_47038,N_47134);
nand U47537 (N_47537,N_47475,N_47405);
nand U47538 (N_47538,N_47417,N_47455);
nand U47539 (N_47539,N_47143,N_47047);
or U47540 (N_47540,N_47101,N_47334);
xor U47541 (N_47541,N_47286,N_47488);
and U47542 (N_47542,N_47431,N_47027);
nor U47543 (N_47543,N_47023,N_47133);
nand U47544 (N_47544,N_47380,N_47485);
nand U47545 (N_47545,N_47365,N_47258);
nand U47546 (N_47546,N_47491,N_47328);
nand U47547 (N_47547,N_47304,N_47190);
nand U47548 (N_47548,N_47440,N_47291);
nand U47549 (N_47549,N_47333,N_47418);
nand U47550 (N_47550,N_47415,N_47111);
xnor U47551 (N_47551,N_47335,N_47071);
and U47552 (N_47552,N_47152,N_47031);
xnor U47553 (N_47553,N_47289,N_47262);
and U47554 (N_47554,N_47069,N_47487);
and U47555 (N_47555,N_47476,N_47421);
xnor U47556 (N_47556,N_47369,N_47426);
nor U47557 (N_47557,N_47486,N_47495);
or U47558 (N_47558,N_47351,N_47465);
or U47559 (N_47559,N_47135,N_47276);
xor U47560 (N_47560,N_47040,N_47237);
nor U47561 (N_47561,N_47126,N_47272);
nand U47562 (N_47562,N_47230,N_47419);
xor U47563 (N_47563,N_47013,N_47144);
nand U47564 (N_47564,N_47068,N_47303);
and U47565 (N_47565,N_47383,N_47046);
and U47566 (N_47566,N_47171,N_47194);
nand U47567 (N_47567,N_47079,N_47367);
or U47568 (N_47568,N_47092,N_47467);
xor U47569 (N_47569,N_47294,N_47412);
xnor U47570 (N_47570,N_47067,N_47162);
nor U47571 (N_47571,N_47241,N_47240);
and U47572 (N_47572,N_47142,N_47281);
nor U47573 (N_47573,N_47016,N_47169);
and U47574 (N_47574,N_47025,N_47179);
xor U47575 (N_47575,N_47138,N_47130);
or U47576 (N_47576,N_47116,N_47245);
nor U47577 (N_47577,N_47127,N_47273);
nand U47578 (N_47578,N_47484,N_47059);
and U47579 (N_47579,N_47355,N_47078);
or U47580 (N_47580,N_47119,N_47124);
nor U47581 (N_47581,N_47393,N_47256);
nor U47582 (N_47582,N_47280,N_47425);
nand U47583 (N_47583,N_47345,N_47228);
and U47584 (N_47584,N_47474,N_47158);
nor U47585 (N_47585,N_47009,N_47100);
nor U47586 (N_47586,N_47155,N_47370);
nor U47587 (N_47587,N_47340,N_47064);
nand U47588 (N_47588,N_47339,N_47048);
xnor U47589 (N_47589,N_47165,N_47480);
or U47590 (N_47590,N_47438,N_47459);
xnor U47591 (N_47591,N_47331,N_47018);
or U47592 (N_47592,N_47344,N_47139);
or U47593 (N_47593,N_47478,N_47060);
nand U47594 (N_47594,N_47056,N_47051);
nor U47595 (N_47595,N_47395,N_47014);
and U47596 (N_47596,N_47357,N_47387);
nand U47597 (N_47597,N_47347,N_47390);
and U47598 (N_47598,N_47498,N_47342);
nand U47599 (N_47599,N_47210,N_47066);
nand U47600 (N_47600,N_47129,N_47427);
nand U47601 (N_47601,N_47320,N_47274);
nand U47602 (N_47602,N_47336,N_47188);
and U47603 (N_47603,N_47184,N_47055);
xnor U47604 (N_47604,N_47375,N_47206);
or U47605 (N_47605,N_47349,N_47472);
xor U47606 (N_47606,N_47350,N_47269);
xnor U47607 (N_47607,N_47310,N_47298);
nor U47608 (N_47608,N_47106,N_47121);
xor U47609 (N_47609,N_47207,N_47074);
and U47610 (N_47610,N_47011,N_47456);
or U47611 (N_47611,N_47032,N_47430);
or U47612 (N_47612,N_47166,N_47037);
or U47613 (N_47613,N_47371,N_47110);
nand U47614 (N_47614,N_47406,N_47172);
and U47615 (N_47615,N_47163,N_47482);
or U47616 (N_47616,N_47209,N_47015);
nand U47617 (N_47617,N_47204,N_47236);
nor U47618 (N_47618,N_47361,N_47282);
nand U47619 (N_47619,N_47225,N_47213);
and U47620 (N_47620,N_47265,N_47235);
nor U47621 (N_47621,N_47243,N_47299);
nand U47622 (N_47622,N_47479,N_47004);
or U47623 (N_47623,N_47413,N_47324);
nand U47624 (N_47624,N_47392,N_47359);
xnor U47625 (N_47625,N_47452,N_47362);
nor U47626 (N_47626,N_47318,N_47122);
nand U47627 (N_47627,N_47466,N_47330);
nand U47628 (N_47628,N_47312,N_47346);
xor U47629 (N_47629,N_47315,N_47211);
or U47630 (N_47630,N_47453,N_47275);
and U47631 (N_47631,N_47192,N_47128);
nor U47632 (N_47632,N_47065,N_47408);
nor U47633 (N_47633,N_47195,N_47113);
nor U47634 (N_47634,N_47458,N_47463);
or U47635 (N_47635,N_47451,N_47096);
and U47636 (N_47636,N_47434,N_47222);
and U47637 (N_47637,N_47360,N_47202);
nor U47638 (N_47638,N_47382,N_47411);
xor U47639 (N_47639,N_47401,N_47264);
and U47640 (N_47640,N_47353,N_47221);
nor U47641 (N_47641,N_47464,N_47232);
nor U47642 (N_47642,N_47376,N_47468);
xnor U47643 (N_47643,N_47091,N_47020);
and U47644 (N_47644,N_47164,N_47087);
nand U47645 (N_47645,N_47073,N_47153);
and U47646 (N_47646,N_47154,N_47049);
nor U47647 (N_47647,N_47193,N_47098);
nor U47648 (N_47648,N_47255,N_47454);
or U47649 (N_47649,N_47061,N_47224);
nor U47650 (N_47650,N_47302,N_47167);
or U47651 (N_47651,N_47120,N_47248);
nor U47652 (N_47652,N_47008,N_47283);
nor U47653 (N_47653,N_47019,N_47034);
and U47654 (N_47654,N_47323,N_47307);
nand U47655 (N_47655,N_47216,N_47381);
nor U47656 (N_47656,N_47377,N_47186);
or U47657 (N_47657,N_47259,N_47215);
or U47658 (N_47658,N_47112,N_47388);
xor U47659 (N_47659,N_47327,N_47352);
and U47660 (N_47660,N_47470,N_47471);
and U47661 (N_47661,N_47338,N_47033);
and U47662 (N_47662,N_47189,N_47099);
nand U47663 (N_47663,N_47226,N_47147);
and U47664 (N_47664,N_47212,N_47402);
nor U47665 (N_47665,N_47436,N_47477);
or U47666 (N_47666,N_47450,N_47145);
or U47667 (N_47667,N_47300,N_47151);
nand U47668 (N_47668,N_47131,N_47414);
xor U47669 (N_47669,N_47322,N_47379);
or U47670 (N_47670,N_47109,N_47218);
nand U47671 (N_47671,N_47284,N_47253);
xor U47672 (N_47672,N_47257,N_47293);
xnor U47673 (N_47673,N_47159,N_47423);
nor U47674 (N_47674,N_47054,N_47077);
nand U47675 (N_47675,N_47437,N_47197);
xor U47676 (N_47676,N_47170,N_47180);
nor U47677 (N_47677,N_47058,N_47010);
xnor U47678 (N_47678,N_47052,N_47448);
or U47679 (N_47679,N_47088,N_47244);
nor U47680 (N_47680,N_47001,N_47337);
and U47681 (N_47681,N_47187,N_47251);
and U47682 (N_47682,N_47288,N_47374);
nand U47683 (N_47683,N_47386,N_47409);
or U47684 (N_47684,N_47341,N_47416);
nand U47685 (N_47685,N_47117,N_47410);
nand U47686 (N_47686,N_47229,N_47270);
xnor U47687 (N_47687,N_47175,N_47354);
nand U47688 (N_47688,N_47000,N_47404);
xnor U47689 (N_47689,N_47385,N_47083);
xor U47690 (N_47690,N_47309,N_47490);
nor U47691 (N_47691,N_47026,N_47118);
nor U47692 (N_47692,N_47160,N_47107);
nand U47693 (N_47693,N_47072,N_47183);
xnor U47694 (N_47694,N_47287,N_47198);
nor U47695 (N_47695,N_47234,N_47203);
nand U47696 (N_47696,N_47247,N_47391);
or U47697 (N_47697,N_47306,N_47090);
and U47698 (N_47698,N_47373,N_47021);
or U47699 (N_47699,N_47044,N_47396);
and U47700 (N_47700,N_47317,N_47080);
and U47701 (N_47701,N_47070,N_47394);
xnor U47702 (N_47702,N_47063,N_47260);
nor U47703 (N_47703,N_47002,N_47429);
nand U47704 (N_47704,N_47492,N_47389);
xnor U47705 (N_47705,N_47267,N_47363);
xor U47706 (N_47706,N_47278,N_47366);
xor U47707 (N_47707,N_47108,N_47136);
nand U47708 (N_47708,N_47177,N_47238);
or U47709 (N_47709,N_47196,N_47115);
xor U47710 (N_47710,N_47089,N_47449);
nor U47711 (N_47711,N_47062,N_47364);
or U47712 (N_47712,N_47301,N_47104);
nand U47713 (N_47713,N_47105,N_47174);
nor U47714 (N_47714,N_47295,N_47086);
or U47715 (N_47715,N_47199,N_47252);
and U47716 (N_47716,N_47246,N_47102);
nor U47717 (N_47717,N_47012,N_47290);
xor U47718 (N_47718,N_47442,N_47141);
or U47719 (N_47719,N_47368,N_47444);
nor U47720 (N_47720,N_47173,N_47481);
xnor U47721 (N_47721,N_47305,N_47233);
or U47722 (N_47722,N_47445,N_47372);
and U47723 (N_47723,N_47205,N_47003);
nor U47724 (N_47724,N_47219,N_47457);
nor U47725 (N_47725,N_47469,N_47494);
xnor U47726 (N_47726,N_47473,N_47053);
xor U47727 (N_47727,N_47085,N_47461);
nor U47728 (N_47728,N_47168,N_47499);
xor U47729 (N_47729,N_47200,N_47314);
xnor U47730 (N_47730,N_47161,N_47384);
or U47731 (N_47731,N_47082,N_47076);
or U47732 (N_47732,N_47447,N_47266);
or U47733 (N_47733,N_47343,N_47261);
or U47734 (N_47734,N_47217,N_47036);
nand U47735 (N_47735,N_47132,N_47041);
and U47736 (N_47736,N_47081,N_47397);
or U47737 (N_47737,N_47050,N_47489);
or U47738 (N_47738,N_47268,N_47493);
nand U47739 (N_47739,N_47148,N_47084);
xnor U47740 (N_47740,N_47249,N_47271);
or U47741 (N_47741,N_47326,N_47399);
nand U47742 (N_47742,N_47191,N_47462);
nand U47743 (N_47743,N_47439,N_47356);
nor U47744 (N_47744,N_47029,N_47201);
xor U47745 (N_47745,N_47150,N_47157);
or U47746 (N_47746,N_47313,N_47435);
nand U47747 (N_47747,N_47358,N_47024);
or U47748 (N_47748,N_47424,N_47407);
or U47749 (N_47749,N_47017,N_47103);
and U47750 (N_47750,N_47324,N_47109);
and U47751 (N_47751,N_47038,N_47493);
nand U47752 (N_47752,N_47082,N_47241);
xnor U47753 (N_47753,N_47123,N_47318);
xor U47754 (N_47754,N_47394,N_47483);
or U47755 (N_47755,N_47399,N_47288);
xor U47756 (N_47756,N_47234,N_47242);
nand U47757 (N_47757,N_47302,N_47241);
xnor U47758 (N_47758,N_47051,N_47190);
xnor U47759 (N_47759,N_47152,N_47390);
nand U47760 (N_47760,N_47080,N_47029);
or U47761 (N_47761,N_47236,N_47073);
or U47762 (N_47762,N_47065,N_47434);
or U47763 (N_47763,N_47385,N_47016);
nand U47764 (N_47764,N_47399,N_47431);
nor U47765 (N_47765,N_47310,N_47061);
and U47766 (N_47766,N_47087,N_47374);
nand U47767 (N_47767,N_47290,N_47317);
or U47768 (N_47768,N_47258,N_47059);
xor U47769 (N_47769,N_47376,N_47211);
and U47770 (N_47770,N_47005,N_47104);
xor U47771 (N_47771,N_47493,N_47186);
xnor U47772 (N_47772,N_47193,N_47348);
and U47773 (N_47773,N_47220,N_47085);
nand U47774 (N_47774,N_47398,N_47354);
nor U47775 (N_47775,N_47354,N_47261);
xnor U47776 (N_47776,N_47410,N_47019);
or U47777 (N_47777,N_47382,N_47273);
nand U47778 (N_47778,N_47056,N_47461);
or U47779 (N_47779,N_47357,N_47437);
nand U47780 (N_47780,N_47081,N_47070);
and U47781 (N_47781,N_47289,N_47053);
or U47782 (N_47782,N_47152,N_47105);
and U47783 (N_47783,N_47488,N_47372);
nor U47784 (N_47784,N_47160,N_47121);
or U47785 (N_47785,N_47211,N_47071);
or U47786 (N_47786,N_47359,N_47327);
and U47787 (N_47787,N_47066,N_47280);
xor U47788 (N_47788,N_47343,N_47268);
nor U47789 (N_47789,N_47218,N_47075);
nor U47790 (N_47790,N_47415,N_47356);
or U47791 (N_47791,N_47106,N_47394);
nor U47792 (N_47792,N_47131,N_47007);
nor U47793 (N_47793,N_47056,N_47273);
and U47794 (N_47794,N_47037,N_47194);
and U47795 (N_47795,N_47189,N_47180);
or U47796 (N_47796,N_47092,N_47133);
or U47797 (N_47797,N_47136,N_47490);
and U47798 (N_47798,N_47273,N_47360);
or U47799 (N_47799,N_47452,N_47093);
nand U47800 (N_47800,N_47391,N_47283);
xnor U47801 (N_47801,N_47065,N_47347);
nor U47802 (N_47802,N_47212,N_47171);
xor U47803 (N_47803,N_47147,N_47266);
nor U47804 (N_47804,N_47009,N_47235);
or U47805 (N_47805,N_47255,N_47384);
nor U47806 (N_47806,N_47109,N_47427);
xor U47807 (N_47807,N_47412,N_47480);
nor U47808 (N_47808,N_47274,N_47446);
nand U47809 (N_47809,N_47202,N_47117);
or U47810 (N_47810,N_47480,N_47300);
or U47811 (N_47811,N_47265,N_47396);
or U47812 (N_47812,N_47153,N_47177);
or U47813 (N_47813,N_47234,N_47083);
nand U47814 (N_47814,N_47440,N_47003);
nand U47815 (N_47815,N_47009,N_47438);
nor U47816 (N_47816,N_47280,N_47256);
nand U47817 (N_47817,N_47449,N_47360);
xor U47818 (N_47818,N_47451,N_47018);
nor U47819 (N_47819,N_47163,N_47318);
xnor U47820 (N_47820,N_47296,N_47047);
nand U47821 (N_47821,N_47499,N_47152);
nor U47822 (N_47822,N_47084,N_47176);
or U47823 (N_47823,N_47130,N_47293);
nor U47824 (N_47824,N_47107,N_47037);
or U47825 (N_47825,N_47033,N_47455);
and U47826 (N_47826,N_47193,N_47416);
and U47827 (N_47827,N_47126,N_47452);
and U47828 (N_47828,N_47493,N_47338);
and U47829 (N_47829,N_47143,N_47246);
or U47830 (N_47830,N_47011,N_47282);
or U47831 (N_47831,N_47494,N_47159);
nor U47832 (N_47832,N_47410,N_47196);
or U47833 (N_47833,N_47318,N_47478);
nor U47834 (N_47834,N_47359,N_47273);
nor U47835 (N_47835,N_47094,N_47080);
nor U47836 (N_47836,N_47045,N_47285);
or U47837 (N_47837,N_47376,N_47499);
nor U47838 (N_47838,N_47239,N_47082);
xor U47839 (N_47839,N_47084,N_47272);
xor U47840 (N_47840,N_47209,N_47366);
and U47841 (N_47841,N_47395,N_47495);
nor U47842 (N_47842,N_47221,N_47340);
or U47843 (N_47843,N_47088,N_47188);
nand U47844 (N_47844,N_47046,N_47321);
nand U47845 (N_47845,N_47379,N_47324);
nand U47846 (N_47846,N_47346,N_47410);
and U47847 (N_47847,N_47369,N_47247);
and U47848 (N_47848,N_47373,N_47326);
nand U47849 (N_47849,N_47024,N_47473);
or U47850 (N_47850,N_47424,N_47402);
and U47851 (N_47851,N_47169,N_47063);
xnor U47852 (N_47852,N_47177,N_47372);
xnor U47853 (N_47853,N_47206,N_47476);
xnor U47854 (N_47854,N_47033,N_47213);
xor U47855 (N_47855,N_47216,N_47130);
xor U47856 (N_47856,N_47180,N_47093);
nor U47857 (N_47857,N_47267,N_47244);
and U47858 (N_47858,N_47492,N_47226);
and U47859 (N_47859,N_47062,N_47262);
nor U47860 (N_47860,N_47338,N_47306);
nand U47861 (N_47861,N_47322,N_47002);
nand U47862 (N_47862,N_47326,N_47032);
xnor U47863 (N_47863,N_47457,N_47410);
xnor U47864 (N_47864,N_47172,N_47307);
nor U47865 (N_47865,N_47447,N_47386);
and U47866 (N_47866,N_47071,N_47234);
nand U47867 (N_47867,N_47397,N_47020);
nor U47868 (N_47868,N_47026,N_47442);
or U47869 (N_47869,N_47354,N_47121);
nor U47870 (N_47870,N_47338,N_47427);
xor U47871 (N_47871,N_47016,N_47302);
xor U47872 (N_47872,N_47125,N_47021);
nand U47873 (N_47873,N_47400,N_47323);
or U47874 (N_47874,N_47351,N_47334);
and U47875 (N_47875,N_47077,N_47124);
nand U47876 (N_47876,N_47447,N_47287);
xor U47877 (N_47877,N_47038,N_47451);
nor U47878 (N_47878,N_47297,N_47462);
xnor U47879 (N_47879,N_47181,N_47402);
or U47880 (N_47880,N_47300,N_47311);
xnor U47881 (N_47881,N_47455,N_47460);
nand U47882 (N_47882,N_47062,N_47311);
and U47883 (N_47883,N_47190,N_47242);
nand U47884 (N_47884,N_47270,N_47126);
and U47885 (N_47885,N_47342,N_47080);
nor U47886 (N_47886,N_47269,N_47005);
xor U47887 (N_47887,N_47441,N_47122);
and U47888 (N_47888,N_47449,N_47343);
or U47889 (N_47889,N_47218,N_47216);
and U47890 (N_47890,N_47031,N_47098);
nand U47891 (N_47891,N_47209,N_47357);
or U47892 (N_47892,N_47410,N_47414);
and U47893 (N_47893,N_47060,N_47461);
or U47894 (N_47894,N_47325,N_47320);
xnor U47895 (N_47895,N_47001,N_47439);
nand U47896 (N_47896,N_47230,N_47373);
nor U47897 (N_47897,N_47236,N_47347);
xnor U47898 (N_47898,N_47405,N_47082);
nand U47899 (N_47899,N_47067,N_47456);
nor U47900 (N_47900,N_47457,N_47498);
and U47901 (N_47901,N_47080,N_47047);
or U47902 (N_47902,N_47473,N_47417);
xnor U47903 (N_47903,N_47041,N_47112);
nor U47904 (N_47904,N_47180,N_47032);
nand U47905 (N_47905,N_47492,N_47336);
and U47906 (N_47906,N_47123,N_47282);
nor U47907 (N_47907,N_47457,N_47069);
or U47908 (N_47908,N_47367,N_47174);
xnor U47909 (N_47909,N_47373,N_47263);
xor U47910 (N_47910,N_47323,N_47273);
nand U47911 (N_47911,N_47234,N_47466);
nand U47912 (N_47912,N_47426,N_47186);
nand U47913 (N_47913,N_47390,N_47175);
nand U47914 (N_47914,N_47015,N_47343);
nor U47915 (N_47915,N_47223,N_47061);
and U47916 (N_47916,N_47081,N_47021);
nand U47917 (N_47917,N_47368,N_47291);
nor U47918 (N_47918,N_47071,N_47355);
nand U47919 (N_47919,N_47263,N_47139);
nor U47920 (N_47920,N_47467,N_47442);
nand U47921 (N_47921,N_47442,N_47131);
nand U47922 (N_47922,N_47118,N_47299);
nor U47923 (N_47923,N_47109,N_47446);
nor U47924 (N_47924,N_47478,N_47225);
and U47925 (N_47925,N_47482,N_47052);
and U47926 (N_47926,N_47177,N_47313);
and U47927 (N_47927,N_47295,N_47447);
or U47928 (N_47928,N_47270,N_47004);
and U47929 (N_47929,N_47423,N_47002);
nor U47930 (N_47930,N_47177,N_47409);
nor U47931 (N_47931,N_47468,N_47388);
xnor U47932 (N_47932,N_47128,N_47431);
nand U47933 (N_47933,N_47077,N_47070);
nor U47934 (N_47934,N_47335,N_47112);
xnor U47935 (N_47935,N_47169,N_47162);
xnor U47936 (N_47936,N_47100,N_47395);
and U47937 (N_47937,N_47203,N_47441);
xor U47938 (N_47938,N_47085,N_47073);
and U47939 (N_47939,N_47402,N_47290);
nor U47940 (N_47940,N_47065,N_47281);
xor U47941 (N_47941,N_47294,N_47130);
nand U47942 (N_47942,N_47233,N_47412);
xnor U47943 (N_47943,N_47471,N_47032);
nand U47944 (N_47944,N_47221,N_47399);
xor U47945 (N_47945,N_47184,N_47113);
xor U47946 (N_47946,N_47397,N_47364);
or U47947 (N_47947,N_47315,N_47002);
nor U47948 (N_47948,N_47375,N_47499);
nand U47949 (N_47949,N_47051,N_47441);
and U47950 (N_47950,N_47043,N_47234);
and U47951 (N_47951,N_47143,N_47445);
nand U47952 (N_47952,N_47006,N_47027);
xor U47953 (N_47953,N_47051,N_47422);
or U47954 (N_47954,N_47426,N_47139);
nor U47955 (N_47955,N_47313,N_47209);
or U47956 (N_47956,N_47154,N_47425);
xor U47957 (N_47957,N_47095,N_47442);
or U47958 (N_47958,N_47101,N_47149);
nor U47959 (N_47959,N_47233,N_47124);
or U47960 (N_47960,N_47196,N_47304);
and U47961 (N_47961,N_47058,N_47146);
or U47962 (N_47962,N_47315,N_47231);
nor U47963 (N_47963,N_47205,N_47335);
xnor U47964 (N_47964,N_47247,N_47418);
nand U47965 (N_47965,N_47129,N_47058);
and U47966 (N_47966,N_47160,N_47109);
or U47967 (N_47967,N_47192,N_47273);
and U47968 (N_47968,N_47019,N_47336);
xnor U47969 (N_47969,N_47163,N_47331);
and U47970 (N_47970,N_47192,N_47392);
nor U47971 (N_47971,N_47400,N_47397);
nor U47972 (N_47972,N_47163,N_47188);
nor U47973 (N_47973,N_47278,N_47348);
nor U47974 (N_47974,N_47293,N_47164);
xnor U47975 (N_47975,N_47049,N_47252);
nor U47976 (N_47976,N_47331,N_47219);
nor U47977 (N_47977,N_47394,N_47143);
xnor U47978 (N_47978,N_47277,N_47069);
nand U47979 (N_47979,N_47199,N_47024);
nor U47980 (N_47980,N_47273,N_47352);
nand U47981 (N_47981,N_47360,N_47280);
nand U47982 (N_47982,N_47415,N_47399);
nor U47983 (N_47983,N_47280,N_47016);
nand U47984 (N_47984,N_47035,N_47276);
nor U47985 (N_47985,N_47300,N_47032);
nor U47986 (N_47986,N_47464,N_47316);
and U47987 (N_47987,N_47149,N_47337);
nor U47988 (N_47988,N_47082,N_47450);
and U47989 (N_47989,N_47377,N_47015);
xnor U47990 (N_47990,N_47173,N_47125);
nor U47991 (N_47991,N_47182,N_47491);
nor U47992 (N_47992,N_47343,N_47085);
and U47993 (N_47993,N_47004,N_47109);
nor U47994 (N_47994,N_47181,N_47086);
and U47995 (N_47995,N_47373,N_47412);
and U47996 (N_47996,N_47365,N_47267);
or U47997 (N_47997,N_47355,N_47419);
and U47998 (N_47998,N_47453,N_47455);
or U47999 (N_47999,N_47269,N_47192);
and U48000 (N_48000,N_47867,N_47777);
xnor U48001 (N_48001,N_47728,N_47774);
and U48002 (N_48002,N_47831,N_47905);
and U48003 (N_48003,N_47588,N_47579);
or U48004 (N_48004,N_47821,N_47711);
nand U48005 (N_48005,N_47845,N_47619);
nand U48006 (N_48006,N_47833,N_47855);
nor U48007 (N_48007,N_47808,N_47775);
nor U48008 (N_48008,N_47875,N_47734);
nand U48009 (N_48009,N_47856,N_47758);
nor U48010 (N_48010,N_47853,N_47832);
or U48011 (N_48011,N_47769,N_47542);
or U48012 (N_48012,N_47989,N_47556);
nor U48013 (N_48013,N_47710,N_47953);
nand U48014 (N_48014,N_47822,N_47538);
xor U48015 (N_48015,N_47693,N_47763);
nand U48016 (N_48016,N_47918,N_47784);
and U48017 (N_48017,N_47799,N_47912);
and U48018 (N_48018,N_47985,N_47692);
nand U48019 (N_48019,N_47502,N_47826);
nor U48020 (N_48020,N_47680,N_47825);
or U48021 (N_48021,N_47932,N_47741);
or U48022 (N_48022,N_47585,N_47590);
and U48023 (N_48023,N_47827,N_47682);
nor U48024 (N_48024,N_47917,N_47852);
nand U48025 (N_48025,N_47963,N_47886);
nand U48026 (N_48026,N_47697,N_47877);
and U48027 (N_48027,N_47636,N_47801);
xor U48028 (N_48028,N_47678,N_47614);
or U48029 (N_48029,N_47771,N_47861);
or U48030 (N_48030,N_47521,N_47851);
and U48031 (N_48031,N_47767,N_47530);
or U48032 (N_48032,N_47837,N_47787);
and U48033 (N_48033,N_47923,N_47978);
nor U48034 (N_48034,N_47737,N_47653);
nor U48035 (N_48035,N_47570,N_47804);
or U48036 (N_48036,N_47543,N_47935);
nor U48037 (N_48037,N_47535,N_47577);
nor U48038 (N_48038,N_47926,N_47715);
nor U48039 (N_48039,N_47562,N_47965);
or U48040 (N_48040,N_47526,N_47914);
and U48041 (N_48041,N_47657,N_47672);
nor U48042 (N_48042,N_47744,N_47794);
nand U48043 (N_48043,N_47760,N_47576);
or U48044 (N_48044,N_47980,N_47990);
nand U48045 (N_48045,N_47584,N_47747);
nand U48046 (N_48046,N_47587,N_47733);
nor U48047 (N_48047,N_47607,N_47709);
nor U48048 (N_48048,N_47949,N_47836);
or U48049 (N_48049,N_47817,N_47726);
nand U48050 (N_48050,N_47762,N_47934);
nand U48051 (N_48051,N_47950,N_47879);
nor U48052 (N_48052,N_47811,N_47776);
or U48053 (N_48053,N_47639,N_47532);
xor U48054 (N_48054,N_47671,N_47999);
nor U48055 (N_48055,N_47522,N_47509);
xnor U48056 (N_48056,N_47644,N_47798);
and U48057 (N_48057,N_47838,N_47878);
or U48058 (N_48058,N_47649,N_47527);
nand U48059 (N_48059,N_47730,N_47885);
or U48060 (N_48060,N_47544,N_47610);
xnor U48061 (N_48061,N_47900,N_47754);
and U48062 (N_48062,N_47647,N_47673);
xnor U48063 (N_48063,N_47541,N_47551);
and U48064 (N_48064,N_47898,N_47891);
nor U48065 (N_48065,N_47604,N_47514);
xnor U48066 (N_48066,N_47596,N_47864);
xnor U48067 (N_48067,N_47515,N_47951);
nand U48068 (N_48068,N_47840,N_47890);
xnor U48069 (N_48069,N_47727,N_47640);
xor U48070 (N_48070,N_47669,N_47518);
xor U48071 (N_48071,N_47651,N_47547);
nor U48072 (N_48072,N_47531,N_47700);
and U48073 (N_48073,N_47504,N_47723);
xor U48074 (N_48074,N_47979,N_47524);
nand U48075 (N_48075,N_47929,N_47847);
or U48076 (N_48076,N_47966,N_47901);
nand U48077 (N_48077,N_47937,N_47605);
or U48078 (N_48078,N_47871,N_47615);
nand U48079 (N_48079,N_47944,N_47906);
and U48080 (N_48080,N_47717,N_47971);
xnor U48081 (N_48081,N_47635,N_47920);
nand U48082 (N_48082,N_47996,N_47788);
nand U48083 (N_48083,N_47998,N_47571);
nand U48084 (N_48084,N_47735,N_47621);
or U48085 (N_48085,N_47789,N_47660);
nor U48086 (N_48086,N_47563,N_47907);
xor U48087 (N_48087,N_47601,N_47959);
nand U48088 (N_48088,N_47573,N_47948);
nand U48089 (N_48089,N_47703,N_47882);
and U48090 (N_48090,N_47930,N_47820);
nand U48091 (N_48091,N_47519,N_47681);
and U48092 (N_48092,N_47553,N_47969);
or U48093 (N_48093,N_47779,N_47706);
and U48094 (N_48094,N_47782,N_47738);
xor U48095 (N_48095,N_47513,N_47714);
nor U48096 (N_48096,N_47752,N_47940);
nor U48097 (N_48097,N_47548,N_47961);
and U48098 (N_48098,N_47984,N_47893);
nor U48099 (N_48099,N_47628,N_47835);
or U48100 (N_48100,N_47667,N_47987);
and U48101 (N_48101,N_47765,N_47954);
xor U48102 (N_48102,N_47997,N_47525);
nand U48103 (N_48103,N_47819,N_47583);
xnor U48104 (N_48104,N_47761,N_47575);
nand U48105 (N_48105,N_47627,N_47591);
or U48106 (N_48106,N_47574,N_47818);
or U48107 (N_48107,N_47824,N_47793);
nand U48108 (N_48108,N_47510,N_47537);
nand U48109 (N_48109,N_47668,N_47582);
nand U48110 (N_48110,N_47505,N_47638);
or U48111 (N_48111,N_47724,N_47815);
nor U48112 (N_48112,N_47523,N_47564);
or U48113 (N_48113,N_47993,N_47659);
nand U48114 (N_48114,N_47873,N_47859);
xor U48115 (N_48115,N_47546,N_47982);
or U48116 (N_48116,N_47972,N_47592);
nor U48117 (N_48117,N_47842,N_47874);
nand U48118 (N_48118,N_47858,N_47609);
nor U48119 (N_48119,N_47854,N_47862);
nor U48120 (N_48120,N_47641,N_47528);
or U48121 (N_48121,N_47828,N_47910);
nor U48122 (N_48122,N_47816,N_47568);
or U48123 (N_48123,N_47974,N_47599);
or U48124 (N_48124,N_47554,N_47536);
nand U48125 (N_48125,N_47566,N_47909);
nand U48126 (N_48126,N_47705,N_47748);
and U48127 (N_48127,N_47589,N_47964);
and U48128 (N_48128,N_47889,N_47939);
or U48129 (N_48129,N_47740,N_47608);
nand U48130 (N_48130,N_47642,N_47720);
nor U48131 (N_48131,N_47970,N_47557);
nand U48132 (N_48132,N_47973,N_47507);
nand U48133 (N_48133,N_47880,N_47648);
and U48134 (N_48134,N_47606,N_47662);
and U48135 (N_48135,N_47823,N_47806);
and U48136 (N_48136,N_47688,N_47931);
xor U48137 (N_48137,N_47704,N_47634);
or U48138 (N_48138,N_47674,N_47839);
xor U48139 (N_48139,N_47743,N_47629);
or U48140 (N_48140,N_47666,N_47729);
nor U48141 (N_48141,N_47722,N_47701);
and U48142 (N_48142,N_47834,N_47511);
and U48143 (N_48143,N_47921,N_47795);
nand U48144 (N_48144,N_47578,N_47742);
nor U48145 (N_48145,N_47529,N_47908);
and U48146 (N_48146,N_47655,N_47708);
and U48147 (N_48147,N_47707,N_47679);
or U48148 (N_48148,N_47683,N_47611);
or U48149 (N_48149,N_47872,N_47942);
nand U48150 (N_48150,N_47612,N_47753);
and U48151 (N_48151,N_47983,N_47665);
xnor U48152 (N_48152,N_47933,N_47516);
nor U48153 (N_48153,N_47580,N_47731);
and U48154 (N_48154,N_47721,N_47746);
nor U48155 (N_48155,N_47791,N_47618);
xor U48156 (N_48156,N_47603,N_47550);
xnor U48157 (N_48157,N_47768,N_47786);
or U48158 (N_48158,N_47915,N_47805);
xor U48159 (N_48159,N_47843,N_47925);
or U48160 (N_48160,N_47764,N_47988);
xnor U48161 (N_48161,N_47713,N_47637);
nor U48162 (N_48162,N_47630,N_47560);
nor U48163 (N_48163,N_47597,N_47892);
and U48164 (N_48164,N_47687,N_47781);
or U48165 (N_48165,N_47745,N_47677);
and U48166 (N_48166,N_47991,N_47616);
xnor U48167 (N_48167,N_47620,N_47897);
nand U48168 (N_48168,N_47622,N_47904);
and U48169 (N_48169,N_47569,N_47780);
nor U48170 (N_48170,N_47626,N_47870);
nand U48171 (N_48171,N_47957,N_47809);
and U48172 (N_48172,N_47895,N_47902);
and U48173 (N_48173,N_47947,N_47958);
nor U48174 (N_48174,N_47623,N_47883);
and U48175 (N_48175,N_47807,N_47863);
xnor U48176 (N_48176,N_47664,N_47981);
nor U48177 (N_48177,N_47975,N_47501);
or U48178 (N_48178,N_47756,N_47749);
xor U48179 (N_48179,N_47732,N_47695);
and U48180 (N_48180,N_47814,N_47995);
nor U48181 (N_48181,N_47773,N_47739);
or U48182 (N_48182,N_47602,N_47846);
xnor U48183 (N_48183,N_47690,N_47955);
and U48184 (N_48184,N_47689,N_47506);
nand U48185 (N_48185,N_47830,N_47927);
and U48186 (N_48186,N_47860,N_47894);
nor U48187 (N_48187,N_47539,N_47876);
nand U48188 (N_48188,N_47943,N_47881);
nor U48189 (N_48189,N_47797,N_47684);
and U48190 (N_48190,N_47661,N_47725);
or U48191 (N_48191,N_47884,N_47887);
or U48192 (N_48192,N_47792,N_47656);
and U48193 (N_48193,N_47699,N_47850);
nand U48194 (N_48194,N_47572,N_47559);
and U48195 (N_48195,N_47631,N_47652);
or U48196 (N_48196,N_47960,N_47718);
nand U48197 (N_48197,N_47552,N_47702);
or U48198 (N_48198,N_47755,N_47658);
xnor U48199 (N_48199,N_47540,N_47936);
xnor U48200 (N_48200,N_47857,N_47586);
or U48201 (N_48201,N_47848,N_47924);
and U48202 (N_48202,N_47561,N_47645);
nor U48203 (N_48203,N_47813,N_47962);
and U48204 (N_48204,N_47508,N_47675);
nand U48205 (N_48205,N_47500,N_47685);
or U48206 (N_48206,N_47654,N_47829);
nand U48207 (N_48207,N_47759,N_47952);
nand U48208 (N_48208,N_47844,N_47751);
and U48209 (N_48209,N_47650,N_47946);
nor U48210 (N_48210,N_47549,N_47785);
xor U48211 (N_48211,N_47869,N_47913);
and U48212 (N_48212,N_47896,N_47766);
nor U48213 (N_48213,N_47812,N_47632);
xnor U48214 (N_48214,N_47956,N_47919);
or U48215 (N_48215,N_47941,N_47694);
nand U48216 (N_48216,N_47750,N_47772);
nor U48217 (N_48217,N_47691,N_47803);
xor U48218 (N_48218,N_47800,N_47967);
nand U48219 (N_48219,N_47643,N_47986);
nor U48220 (N_48220,N_47992,N_47533);
nand U48221 (N_48221,N_47617,N_47790);
or U48222 (N_48222,N_47770,N_47646);
xnor U48223 (N_48223,N_47778,N_47676);
nand U48224 (N_48224,N_47938,N_47968);
nor U48225 (N_48225,N_47670,N_47976);
or U48226 (N_48226,N_47911,N_47868);
nand U48227 (N_48227,N_47916,N_47595);
nor U48228 (N_48228,N_47593,N_47565);
and U48229 (N_48229,N_47633,N_47712);
xor U48230 (N_48230,N_47866,N_47567);
xor U48231 (N_48231,N_47849,N_47810);
and U48232 (N_48232,N_47686,N_47625);
or U48233 (N_48233,N_47757,N_47512);
xor U48234 (N_48234,N_47520,N_47928);
nor U48235 (N_48235,N_47716,N_47696);
xor U48236 (N_48236,N_47977,N_47736);
xnor U48237 (N_48237,N_47598,N_47613);
and U48238 (N_48238,N_47581,N_47899);
and U48239 (N_48239,N_47841,N_47624);
nand U48240 (N_48240,N_47802,N_47594);
xor U48241 (N_48241,N_47945,N_47503);
nor U48242 (N_48242,N_47865,N_47698);
nor U48243 (N_48243,N_47555,N_47888);
nand U48244 (N_48244,N_47663,N_47922);
xnor U48245 (N_48245,N_47783,N_47994);
xnor U48246 (N_48246,N_47600,N_47719);
xnor U48247 (N_48247,N_47534,N_47545);
or U48248 (N_48248,N_47903,N_47558);
xnor U48249 (N_48249,N_47796,N_47517);
xnor U48250 (N_48250,N_47943,N_47598);
nand U48251 (N_48251,N_47595,N_47939);
or U48252 (N_48252,N_47715,N_47780);
nor U48253 (N_48253,N_47809,N_47663);
nor U48254 (N_48254,N_47529,N_47673);
nand U48255 (N_48255,N_47694,N_47825);
and U48256 (N_48256,N_47766,N_47618);
xnor U48257 (N_48257,N_47583,N_47848);
nand U48258 (N_48258,N_47993,N_47923);
or U48259 (N_48259,N_47568,N_47917);
and U48260 (N_48260,N_47630,N_47844);
and U48261 (N_48261,N_47984,N_47913);
nor U48262 (N_48262,N_47913,N_47516);
nor U48263 (N_48263,N_47533,N_47984);
or U48264 (N_48264,N_47934,N_47727);
nand U48265 (N_48265,N_47848,N_47605);
and U48266 (N_48266,N_47576,N_47620);
nor U48267 (N_48267,N_47639,N_47749);
nand U48268 (N_48268,N_47793,N_47894);
nor U48269 (N_48269,N_47879,N_47563);
nand U48270 (N_48270,N_47732,N_47700);
xnor U48271 (N_48271,N_47741,N_47935);
nor U48272 (N_48272,N_47518,N_47645);
nor U48273 (N_48273,N_47833,N_47735);
xor U48274 (N_48274,N_47876,N_47768);
nand U48275 (N_48275,N_47965,N_47718);
or U48276 (N_48276,N_47877,N_47807);
or U48277 (N_48277,N_47570,N_47822);
xor U48278 (N_48278,N_47818,N_47742);
or U48279 (N_48279,N_47663,N_47996);
nand U48280 (N_48280,N_47803,N_47552);
xor U48281 (N_48281,N_47746,N_47639);
xnor U48282 (N_48282,N_47881,N_47982);
and U48283 (N_48283,N_47791,N_47657);
or U48284 (N_48284,N_47608,N_47734);
nand U48285 (N_48285,N_47550,N_47888);
nand U48286 (N_48286,N_47883,N_47532);
xor U48287 (N_48287,N_47569,N_47998);
nand U48288 (N_48288,N_47787,N_47645);
nor U48289 (N_48289,N_47863,N_47984);
nand U48290 (N_48290,N_47966,N_47575);
and U48291 (N_48291,N_47720,N_47690);
nand U48292 (N_48292,N_47525,N_47606);
nand U48293 (N_48293,N_47586,N_47992);
nor U48294 (N_48294,N_47836,N_47782);
and U48295 (N_48295,N_47639,N_47689);
nor U48296 (N_48296,N_47519,N_47811);
or U48297 (N_48297,N_47629,N_47795);
nor U48298 (N_48298,N_47679,N_47681);
nand U48299 (N_48299,N_47705,N_47995);
nand U48300 (N_48300,N_47689,N_47895);
nand U48301 (N_48301,N_47813,N_47563);
and U48302 (N_48302,N_47856,N_47740);
nor U48303 (N_48303,N_47929,N_47500);
and U48304 (N_48304,N_47978,N_47946);
and U48305 (N_48305,N_47744,N_47667);
nand U48306 (N_48306,N_47630,N_47815);
and U48307 (N_48307,N_47889,N_47759);
and U48308 (N_48308,N_47618,N_47990);
or U48309 (N_48309,N_47908,N_47665);
and U48310 (N_48310,N_47951,N_47808);
or U48311 (N_48311,N_47986,N_47895);
nor U48312 (N_48312,N_47770,N_47647);
and U48313 (N_48313,N_47811,N_47501);
and U48314 (N_48314,N_47681,N_47773);
nor U48315 (N_48315,N_47838,N_47975);
nand U48316 (N_48316,N_47684,N_47533);
nor U48317 (N_48317,N_47862,N_47960);
nand U48318 (N_48318,N_47680,N_47585);
and U48319 (N_48319,N_47964,N_47750);
nor U48320 (N_48320,N_47822,N_47834);
nand U48321 (N_48321,N_47771,N_47967);
nand U48322 (N_48322,N_47525,N_47771);
nor U48323 (N_48323,N_47960,N_47691);
nand U48324 (N_48324,N_47560,N_47975);
nand U48325 (N_48325,N_47893,N_47530);
nor U48326 (N_48326,N_47897,N_47526);
nor U48327 (N_48327,N_47569,N_47534);
or U48328 (N_48328,N_47798,N_47948);
nand U48329 (N_48329,N_47914,N_47577);
and U48330 (N_48330,N_47550,N_47583);
xor U48331 (N_48331,N_47517,N_47798);
nor U48332 (N_48332,N_47997,N_47521);
nand U48333 (N_48333,N_47734,N_47841);
or U48334 (N_48334,N_47532,N_47578);
and U48335 (N_48335,N_47783,N_47989);
or U48336 (N_48336,N_47686,N_47674);
nor U48337 (N_48337,N_47629,N_47974);
and U48338 (N_48338,N_47633,N_47760);
nor U48339 (N_48339,N_47711,N_47960);
and U48340 (N_48340,N_47835,N_47857);
xor U48341 (N_48341,N_47722,N_47811);
xor U48342 (N_48342,N_47603,N_47728);
or U48343 (N_48343,N_47787,N_47655);
nand U48344 (N_48344,N_47784,N_47753);
and U48345 (N_48345,N_47850,N_47650);
nand U48346 (N_48346,N_47824,N_47937);
or U48347 (N_48347,N_47908,N_47766);
xnor U48348 (N_48348,N_47545,N_47542);
nor U48349 (N_48349,N_47892,N_47612);
nand U48350 (N_48350,N_47903,N_47908);
xnor U48351 (N_48351,N_47991,N_47822);
and U48352 (N_48352,N_47876,N_47549);
nand U48353 (N_48353,N_47747,N_47549);
and U48354 (N_48354,N_47506,N_47789);
xnor U48355 (N_48355,N_47682,N_47809);
nor U48356 (N_48356,N_47585,N_47732);
xor U48357 (N_48357,N_47673,N_47653);
or U48358 (N_48358,N_47789,N_47594);
and U48359 (N_48359,N_47791,N_47752);
and U48360 (N_48360,N_47842,N_47766);
or U48361 (N_48361,N_47541,N_47795);
nor U48362 (N_48362,N_47998,N_47819);
or U48363 (N_48363,N_47869,N_47689);
nor U48364 (N_48364,N_47724,N_47890);
and U48365 (N_48365,N_47979,N_47685);
and U48366 (N_48366,N_47824,N_47810);
and U48367 (N_48367,N_47596,N_47886);
xnor U48368 (N_48368,N_47710,N_47674);
nor U48369 (N_48369,N_47509,N_47709);
and U48370 (N_48370,N_47522,N_47978);
nand U48371 (N_48371,N_47826,N_47718);
nor U48372 (N_48372,N_47654,N_47614);
nand U48373 (N_48373,N_47789,N_47518);
or U48374 (N_48374,N_47718,N_47795);
nor U48375 (N_48375,N_47816,N_47615);
nand U48376 (N_48376,N_47501,N_47884);
and U48377 (N_48377,N_47697,N_47740);
or U48378 (N_48378,N_47613,N_47589);
xnor U48379 (N_48379,N_47547,N_47921);
nor U48380 (N_48380,N_47889,N_47814);
nand U48381 (N_48381,N_47637,N_47670);
xor U48382 (N_48382,N_47786,N_47562);
or U48383 (N_48383,N_47837,N_47823);
xnor U48384 (N_48384,N_47502,N_47655);
nor U48385 (N_48385,N_47983,N_47922);
nor U48386 (N_48386,N_47793,N_47572);
nand U48387 (N_48387,N_47924,N_47866);
or U48388 (N_48388,N_47744,N_47668);
or U48389 (N_48389,N_47833,N_47545);
or U48390 (N_48390,N_47583,N_47785);
or U48391 (N_48391,N_47919,N_47748);
nor U48392 (N_48392,N_47623,N_47863);
nand U48393 (N_48393,N_47996,N_47988);
and U48394 (N_48394,N_47562,N_47824);
or U48395 (N_48395,N_47956,N_47979);
nand U48396 (N_48396,N_47811,N_47902);
or U48397 (N_48397,N_47810,N_47608);
or U48398 (N_48398,N_47694,N_47713);
nand U48399 (N_48399,N_47644,N_47506);
nand U48400 (N_48400,N_47963,N_47808);
nand U48401 (N_48401,N_47936,N_47839);
xor U48402 (N_48402,N_47513,N_47971);
nor U48403 (N_48403,N_47566,N_47978);
or U48404 (N_48404,N_47729,N_47672);
or U48405 (N_48405,N_47552,N_47695);
and U48406 (N_48406,N_47817,N_47905);
nor U48407 (N_48407,N_47594,N_47645);
or U48408 (N_48408,N_47526,N_47862);
nand U48409 (N_48409,N_47733,N_47584);
or U48410 (N_48410,N_47785,N_47888);
or U48411 (N_48411,N_47774,N_47711);
nand U48412 (N_48412,N_47878,N_47971);
nand U48413 (N_48413,N_47980,N_47812);
xor U48414 (N_48414,N_47543,N_47898);
or U48415 (N_48415,N_47529,N_47812);
nor U48416 (N_48416,N_47703,N_47608);
nand U48417 (N_48417,N_47556,N_47831);
xor U48418 (N_48418,N_47878,N_47564);
or U48419 (N_48419,N_47560,N_47787);
nand U48420 (N_48420,N_47737,N_47561);
nor U48421 (N_48421,N_47691,N_47677);
nand U48422 (N_48422,N_47704,N_47964);
or U48423 (N_48423,N_47604,N_47851);
nor U48424 (N_48424,N_47688,N_47592);
xor U48425 (N_48425,N_47580,N_47794);
or U48426 (N_48426,N_47965,N_47855);
or U48427 (N_48427,N_47795,N_47542);
nor U48428 (N_48428,N_47726,N_47742);
or U48429 (N_48429,N_47619,N_47789);
or U48430 (N_48430,N_47981,N_47749);
nand U48431 (N_48431,N_47896,N_47794);
nand U48432 (N_48432,N_47577,N_47648);
xnor U48433 (N_48433,N_47628,N_47593);
nand U48434 (N_48434,N_47521,N_47837);
xnor U48435 (N_48435,N_47703,N_47974);
nor U48436 (N_48436,N_47545,N_47979);
or U48437 (N_48437,N_47579,N_47710);
nand U48438 (N_48438,N_47684,N_47570);
nand U48439 (N_48439,N_47699,N_47841);
nor U48440 (N_48440,N_47956,N_47543);
xnor U48441 (N_48441,N_47564,N_47795);
nand U48442 (N_48442,N_47897,N_47908);
nor U48443 (N_48443,N_47871,N_47792);
xor U48444 (N_48444,N_47611,N_47666);
xnor U48445 (N_48445,N_47771,N_47528);
nand U48446 (N_48446,N_47815,N_47645);
xor U48447 (N_48447,N_47661,N_47913);
nand U48448 (N_48448,N_47931,N_47669);
or U48449 (N_48449,N_47752,N_47603);
or U48450 (N_48450,N_47762,N_47662);
nand U48451 (N_48451,N_47896,N_47936);
xnor U48452 (N_48452,N_47992,N_47539);
xor U48453 (N_48453,N_47626,N_47526);
and U48454 (N_48454,N_47785,N_47753);
nand U48455 (N_48455,N_47696,N_47965);
or U48456 (N_48456,N_47611,N_47774);
and U48457 (N_48457,N_47752,N_47958);
nor U48458 (N_48458,N_47658,N_47821);
or U48459 (N_48459,N_47947,N_47990);
xor U48460 (N_48460,N_47936,N_47772);
nand U48461 (N_48461,N_47593,N_47606);
nand U48462 (N_48462,N_47922,N_47793);
or U48463 (N_48463,N_47813,N_47914);
nor U48464 (N_48464,N_47535,N_47634);
or U48465 (N_48465,N_47557,N_47931);
nor U48466 (N_48466,N_47841,N_47886);
or U48467 (N_48467,N_47514,N_47528);
nor U48468 (N_48468,N_47913,N_47589);
nor U48469 (N_48469,N_47887,N_47650);
or U48470 (N_48470,N_47826,N_47789);
or U48471 (N_48471,N_47666,N_47755);
nor U48472 (N_48472,N_47923,N_47891);
nand U48473 (N_48473,N_47937,N_47799);
nor U48474 (N_48474,N_47633,N_47673);
and U48475 (N_48475,N_47766,N_47637);
nand U48476 (N_48476,N_47825,N_47805);
nand U48477 (N_48477,N_47531,N_47567);
nand U48478 (N_48478,N_47582,N_47993);
xor U48479 (N_48479,N_47871,N_47996);
nor U48480 (N_48480,N_47948,N_47892);
nand U48481 (N_48481,N_47517,N_47548);
and U48482 (N_48482,N_47758,N_47903);
nor U48483 (N_48483,N_47938,N_47916);
or U48484 (N_48484,N_47702,N_47622);
or U48485 (N_48485,N_47617,N_47531);
nand U48486 (N_48486,N_47532,N_47754);
nor U48487 (N_48487,N_47960,N_47662);
or U48488 (N_48488,N_47836,N_47700);
nor U48489 (N_48489,N_47511,N_47542);
nor U48490 (N_48490,N_47680,N_47560);
xor U48491 (N_48491,N_47656,N_47764);
nand U48492 (N_48492,N_47610,N_47962);
or U48493 (N_48493,N_47772,N_47665);
or U48494 (N_48494,N_47929,N_47850);
nor U48495 (N_48495,N_47770,N_47778);
xor U48496 (N_48496,N_47954,N_47782);
and U48497 (N_48497,N_47954,N_47710);
or U48498 (N_48498,N_47691,N_47841);
nand U48499 (N_48499,N_47980,N_47902);
or U48500 (N_48500,N_48032,N_48405);
or U48501 (N_48501,N_48464,N_48013);
nand U48502 (N_48502,N_48471,N_48340);
nand U48503 (N_48503,N_48285,N_48179);
nor U48504 (N_48504,N_48237,N_48304);
xnor U48505 (N_48505,N_48201,N_48117);
and U48506 (N_48506,N_48165,N_48494);
nand U48507 (N_48507,N_48424,N_48188);
nor U48508 (N_48508,N_48328,N_48491);
xnor U48509 (N_48509,N_48426,N_48219);
and U48510 (N_48510,N_48394,N_48287);
and U48511 (N_48511,N_48213,N_48008);
or U48512 (N_48512,N_48159,N_48296);
or U48513 (N_48513,N_48356,N_48072);
nand U48514 (N_48514,N_48268,N_48468);
xor U48515 (N_48515,N_48455,N_48336);
and U48516 (N_48516,N_48205,N_48136);
xor U48517 (N_48517,N_48300,N_48099);
xor U48518 (N_48518,N_48087,N_48191);
nand U48519 (N_48519,N_48396,N_48104);
nor U48520 (N_48520,N_48027,N_48453);
nand U48521 (N_48521,N_48315,N_48368);
xnor U48522 (N_48522,N_48390,N_48395);
nor U48523 (N_48523,N_48193,N_48005);
nand U48524 (N_48524,N_48323,N_48123);
xor U48525 (N_48525,N_48486,N_48383);
and U48526 (N_48526,N_48298,N_48399);
and U48527 (N_48527,N_48065,N_48366);
nand U48528 (N_48528,N_48319,N_48031);
and U48529 (N_48529,N_48427,N_48387);
and U48530 (N_48530,N_48046,N_48433);
and U48531 (N_48531,N_48158,N_48373);
xor U48532 (N_48532,N_48009,N_48348);
and U48533 (N_48533,N_48052,N_48311);
xnor U48534 (N_48534,N_48037,N_48370);
nand U48535 (N_48535,N_48185,N_48406);
nor U48536 (N_48536,N_48422,N_48187);
nor U48537 (N_48537,N_48275,N_48217);
xnor U48538 (N_48538,N_48262,N_48174);
xnor U48539 (N_48539,N_48404,N_48069);
and U48540 (N_48540,N_48246,N_48408);
and U48541 (N_48541,N_48225,N_48147);
or U48542 (N_48542,N_48282,N_48414);
nand U48543 (N_48543,N_48049,N_48290);
or U48544 (N_48544,N_48301,N_48145);
xnor U48545 (N_48545,N_48128,N_48445);
or U48546 (N_48546,N_48017,N_48164);
xnor U48547 (N_48547,N_48271,N_48428);
and U48548 (N_48548,N_48284,N_48143);
and U48549 (N_48549,N_48144,N_48379);
and U48550 (N_48550,N_48011,N_48086);
xnor U48551 (N_48551,N_48446,N_48261);
nand U48552 (N_48552,N_48239,N_48059);
nand U48553 (N_48553,N_48258,N_48444);
nand U48554 (N_48554,N_48350,N_48389);
and U48555 (N_48555,N_48153,N_48060);
nand U48556 (N_48556,N_48007,N_48110);
and U48557 (N_48557,N_48068,N_48266);
nor U48558 (N_48558,N_48384,N_48121);
nor U48559 (N_48559,N_48369,N_48091);
nor U48560 (N_48560,N_48294,N_48251);
nor U48561 (N_48561,N_48126,N_48056);
or U48562 (N_48562,N_48160,N_48197);
and U48563 (N_48563,N_48460,N_48139);
and U48564 (N_48564,N_48089,N_48302);
and U48565 (N_48565,N_48498,N_48034);
and U48566 (N_48566,N_48088,N_48295);
xor U48567 (N_48567,N_48211,N_48398);
and U48568 (N_48568,N_48478,N_48359);
xnor U48569 (N_48569,N_48434,N_48083);
xor U48570 (N_48570,N_48475,N_48331);
or U48571 (N_48571,N_48283,N_48012);
nand U48572 (N_48572,N_48452,N_48157);
or U48573 (N_48573,N_48047,N_48463);
and U48574 (N_48574,N_48499,N_48403);
nand U48575 (N_48575,N_48353,N_48004);
nand U48576 (N_48576,N_48106,N_48272);
nor U48577 (N_48577,N_48002,N_48163);
and U48578 (N_48578,N_48410,N_48364);
nor U48579 (N_48579,N_48097,N_48352);
xor U48580 (N_48580,N_48076,N_48462);
nand U48581 (N_48581,N_48092,N_48289);
xnor U48582 (N_48582,N_48469,N_48199);
or U48583 (N_48583,N_48149,N_48345);
nor U48584 (N_48584,N_48150,N_48280);
or U48585 (N_48585,N_48200,N_48074);
or U48586 (N_48586,N_48210,N_48124);
nand U48587 (N_48587,N_48137,N_48443);
xor U48588 (N_48588,N_48112,N_48357);
and U48589 (N_48589,N_48098,N_48391);
or U48590 (N_48590,N_48080,N_48477);
xor U48591 (N_48591,N_48223,N_48079);
nor U48592 (N_48592,N_48381,N_48448);
nand U48593 (N_48593,N_48053,N_48155);
nor U48594 (N_48594,N_48423,N_48024);
nor U48595 (N_48595,N_48335,N_48479);
nor U48596 (N_48596,N_48413,N_48156);
or U48597 (N_48597,N_48279,N_48457);
and U48598 (N_48598,N_48485,N_48317);
xor U48599 (N_48599,N_48062,N_48209);
or U48600 (N_48600,N_48073,N_48376);
and U48601 (N_48601,N_48194,N_48162);
xor U48602 (N_48602,N_48385,N_48299);
nor U48603 (N_48603,N_48343,N_48168);
or U48604 (N_48604,N_48016,N_48267);
nand U48605 (N_48605,N_48313,N_48361);
and U48606 (N_48606,N_48467,N_48257);
xor U48607 (N_48607,N_48135,N_48130);
nor U48608 (N_48608,N_48263,N_48248);
nand U48609 (N_48609,N_48397,N_48242);
nor U48610 (N_48610,N_48273,N_48349);
xnor U48611 (N_48611,N_48245,N_48231);
and U48612 (N_48612,N_48182,N_48419);
and U48613 (N_48613,N_48264,N_48167);
or U48614 (N_48614,N_48067,N_48456);
nor U48615 (N_48615,N_48429,N_48442);
xor U48616 (N_48616,N_48438,N_48222);
or U48617 (N_48617,N_48186,N_48189);
and U48618 (N_48618,N_48496,N_48006);
or U48619 (N_48619,N_48041,N_48244);
and U48620 (N_48620,N_48255,N_48288);
or U48621 (N_48621,N_48202,N_48240);
xnor U48622 (N_48622,N_48487,N_48044);
or U48623 (N_48623,N_48458,N_48449);
and U48624 (N_48624,N_48447,N_48019);
nand U48625 (N_48625,N_48082,N_48171);
xor U48626 (N_48626,N_48105,N_48281);
xnor U48627 (N_48627,N_48161,N_48127);
xor U48628 (N_48628,N_48293,N_48178);
nor U48629 (N_48629,N_48192,N_48380);
nor U48630 (N_48630,N_48101,N_48474);
xnor U48631 (N_48631,N_48259,N_48030);
nand U48632 (N_48632,N_48324,N_48085);
xor U48633 (N_48633,N_48071,N_48152);
nand U48634 (N_48634,N_48431,N_48206);
nor U48635 (N_48635,N_48409,N_48420);
xnor U48636 (N_48636,N_48039,N_48221);
and U48637 (N_48637,N_48354,N_48040);
and U48638 (N_48638,N_48115,N_48325);
or U48639 (N_48639,N_48208,N_48363);
and U48640 (N_48640,N_48400,N_48138);
nor U48641 (N_48641,N_48274,N_48081);
or U48642 (N_48642,N_48392,N_48236);
nand U48643 (N_48643,N_48297,N_48465);
and U48644 (N_48644,N_48234,N_48094);
nor U48645 (N_48645,N_48113,N_48175);
or U48646 (N_48646,N_48358,N_48227);
xor U48647 (N_48647,N_48412,N_48181);
nand U48648 (N_48648,N_48365,N_48241);
nor U48649 (N_48649,N_48061,N_48411);
xnor U48650 (N_48650,N_48393,N_48107);
xnor U48651 (N_48651,N_48440,N_48022);
xor U48652 (N_48652,N_48309,N_48307);
or U48653 (N_48653,N_48064,N_48450);
or U48654 (N_48654,N_48020,N_48042);
nor U48655 (N_48655,N_48235,N_48292);
and U48656 (N_48656,N_48341,N_48054);
and U48657 (N_48657,N_48125,N_48483);
xnor U48658 (N_48658,N_48382,N_48035);
nand U48659 (N_48659,N_48220,N_48131);
or U48660 (N_48660,N_48430,N_48184);
nor U48661 (N_48661,N_48493,N_48332);
and U48662 (N_48662,N_48407,N_48377);
nand U48663 (N_48663,N_48484,N_48025);
and U48664 (N_48664,N_48371,N_48269);
nor U48665 (N_48665,N_48001,N_48432);
nand U48666 (N_48666,N_48229,N_48333);
nor U48667 (N_48667,N_48495,N_48003);
nand U48668 (N_48668,N_48111,N_48388);
or U48669 (N_48669,N_48488,N_48439);
or U48670 (N_48670,N_48226,N_48166);
xnor U48671 (N_48671,N_48416,N_48015);
and U48672 (N_48672,N_48134,N_48492);
nand U48673 (N_48673,N_48095,N_48109);
nand U48674 (N_48674,N_48203,N_48466);
and U48675 (N_48675,N_48114,N_48250);
and U48676 (N_48676,N_48055,N_48421);
and U48677 (N_48677,N_48334,N_48063);
nand U48678 (N_48678,N_48146,N_48118);
xnor U48679 (N_48679,N_48310,N_48473);
and U48680 (N_48680,N_48344,N_48362);
nand U48681 (N_48681,N_48119,N_48230);
nand U48682 (N_48682,N_48314,N_48051);
nor U48683 (N_48683,N_48253,N_48129);
xor U48684 (N_48684,N_48215,N_48048);
xnor U48685 (N_48685,N_48330,N_48077);
nand U48686 (N_48686,N_48254,N_48151);
nor U48687 (N_48687,N_48102,N_48472);
or U48688 (N_48688,N_48096,N_48000);
nand U48689 (N_48689,N_48322,N_48351);
and U48690 (N_48690,N_48238,N_48026);
and U48691 (N_48691,N_48276,N_48260);
nor U48692 (N_48692,N_48023,N_48122);
and U48693 (N_48693,N_48176,N_48436);
and U48694 (N_48694,N_48372,N_48338);
and U48695 (N_48695,N_48228,N_48247);
nand U48696 (N_48696,N_48342,N_48378);
xor U48697 (N_48697,N_48021,N_48497);
nand U48698 (N_48698,N_48033,N_48133);
nor U48699 (N_48699,N_48265,N_48093);
xnor U48700 (N_48700,N_48320,N_48252);
nor U48701 (N_48701,N_48489,N_48141);
xor U48702 (N_48702,N_48036,N_48103);
nand U48703 (N_48703,N_48454,N_48018);
or U48704 (N_48704,N_48190,N_48154);
xor U48705 (N_48705,N_48216,N_48401);
xnor U48706 (N_48706,N_48437,N_48169);
and U48707 (N_48707,N_48078,N_48195);
xnor U48708 (N_48708,N_48337,N_48090);
xor U48709 (N_48709,N_48318,N_48476);
xnor U48710 (N_48710,N_48441,N_48305);
nor U48711 (N_48711,N_48347,N_48170);
or U48712 (N_48712,N_48417,N_48142);
and U48713 (N_48713,N_48470,N_48029);
xor U48714 (N_48714,N_48327,N_48256);
nand U48715 (N_48715,N_48243,N_48367);
or U48716 (N_48716,N_48291,N_48207);
nor U48717 (N_48717,N_48196,N_48116);
and U48718 (N_48718,N_48312,N_48329);
or U48719 (N_48719,N_48066,N_48058);
nor U48720 (N_48720,N_48132,N_48451);
and U48721 (N_48721,N_48277,N_48084);
and U48722 (N_48722,N_48233,N_48375);
and U48723 (N_48723,N_48270,N_48481);
nand U48724 (N_48724,N_48425,N_48326);
xor U48725 (N_48725,N_48316,N_48461);
nand U48726 (N_48726,N_48218,N_48180);
nor U48727 (N_48727,N_48435,N_48415);
nand U48728 (N_48728,N_48212,N_48308);
xnor U48729 (N_48729,N_48490,N_48303);
or U48730 (N_48730,N_48321,N_48172);
xor U48731 (N_48731,N_48482,N_48214);
xor U48732 (N_48732,N_48232,N_48386);
or U48733 (N_48733,N_48140,N_48183);
nand U48734 (N_48734,N_48374,N_48339);
nand U48735 (N_48735,N_48120,N_48418);
or U48736 (N_48736,N_48360,N_48402);
or U48737 (N_48737,N_48224,N_48249);
xor U48738 (N_48738,N_48278,N_48346);
and U48739 (N_48739,N_48306,N_48045);
or U48740 (N_48740,N_48286,N_48043);
or U48741 (N_48741,N_48355,N_48075);
nand U48742 (N_48742,N_48173,N_48010);
nor U48743 (N_48743,N_48038,N_48459);
nand U48744 (N_48744,N_48057,N_48050);
nand U48745 (N_48745,N_48480,N_48198);
nand U48746 (N_48746,N_48148,N_48177);
xor U48747 (N_48747,N_48070,N_48100);
xnor U48748 (N_48748,N_48204,N_48108);
or U48749 (N_48749,N_48028,N_48014);
and U48750 (N_48750,N_48138,N_48491);
and U48751 (N_48751,N_48452,N_48040);
xor U48752 (N_48752,N_48368,N_48053);
nand U48753 (N_48753,N_48428,N_48391);
and U48754 (N_48754,N_48083,N_48355);
nand U48755 (N_48755,N_48032,N_48342);
xnor U48756 (N_48756,N_48350,N_48222);
nand U48757 (N_48757,N_48102,N_48446);
nand U48758 (N_48758,N_48085,N_48417);
nor U48759 (N_48759,N_48418,N_48043);
or U48760 (N_48760,N_48463,N_48467);
nand U48761 (N_48761,N_48025,N_48109);
nand U48762 (N_48762,N_48422,N_48005);
nor U48763 (N_48763,N_48352,N_48006);
and U48764 (N_48764,N_48150,N_48419);
and U48765 (N_48765,N_48042,N_48468);
xor U48766 (N_48766,N_48378,N_48259);
nor U48767 (N_48767,N_48022,N_48220);
or U48768 (N_48768,N_48038,N_48242);
or U48769 (N_48769,N_48209,N_48093);
nor U48770 (N_48770,N_48346,N_48418);
nor U48771 (N_48771,N_48426,N_48482);
nor U48772 (N_48772,N_48066,N_48211);
xor U48773 (N_48773,N_48282,N_48370);
nor U48774 (N_48774,N_48327,N_48071);
xor U48775 (N_48775,N_48051,N_48498);
and U48776 (N_48776,N_48481,N_48454);
nand U48777 (N_48777,N_48093,N_48234);
nand U48778 (N_48778,N_48196,N_48113);
nor U48779 (N_48779,N_48470,N_48390);
and U48780 (N_48780,N_48079,N_48074);
xor U48781 (N_48781,N_48128,N_48065);
or U48782 (N_48782,N_48376,N_48218);
or U48783 (N_48783,N_48160,N_48269);
nand U48784 (N_48784,N_48054,N_48416);
or U48785 (N_48785,N_48339,N_48218);
xnor U48786 (N_48786,N_48253,N_48067);
nand U48787 (N_48787,N_48274,N_48196);
nor U48788 (N_48788,N_48220,N_48109);
or U48789 (N_48789,N_48076,N_48421);
nand U48790 (N_48790,N_48126,N_48175);
or U48791 (N_48791,N_48441,N_48121);
xor U48792 (N_48792,N_48328,N_48482);
nor U48793 (N_48793,N_48414,N_48387);
or U48794 (N_48794,N_48027,N_48304);
nor U48795 (N_48795,N_48450,N_48195);
or U48796 (N_48796,N_48382,N_48268);
and U48797 (N_48797,N_48429,N_48195);
or U48798 (N_48798,N_48329,N_48023);
nor U48799 (N_48799,N_48060,N_48044);
and U48800 (N_48800,N_48387,N_48007);
or U48801 (N_48801,N_48271,N_48195);
or U48802 (N_48802,N_48109,N_48114);
xnor U48803 (N_48803,N_48308,N_48144);
or U48804 (N_48804,N_48085,N_48311);
xnor U48805 (N_48805,N_48227,N_48281);
nor U48806 (N_48806,N_48132,N_48186);
or U48807 (N_48807,N_48006,N_48063);
nand U48808 (N_48808,N_48004,N_48197);
nor U48809 (N_48809,N_48186,N_48012);
xnor U48810 (N_48810,N_48302,N_48299);
xor U48811 (N_48811,N_48151,N_48032);
nand U48812 (N_48812,N_48435,N_48011);
xnor U48813 (N_48813,N_48040,N_48099);
xor U48814 (N_48814,N_48375,N_48456);
xnor U48815 (N_48815,N_48103,N_48195);
nand U48816 (N_48816,N_48421,N_48475);
nor U48817 (N_48817,N_48382,N_48425);
nor U48818 (N_48818,N_48373,N_48096);
nand U48819 (N_48819,N_48109,N_48302);
or U48820 (N_48820,N_48288,N_48221);
or U48821 (N_48821,N_48263,N_48481);
or U48822 (N_48822,N_48122,N_48104);
xor U48823 (N_48823,N_48422,N_48333);
xnor U48824 (N_48824,N_48292,N_48152);
or U48825 (N_48825,N_48098,N_48065);
nor U48826 (N_48826,N_48141,N_48198);
nand U48827 (N_48827,N_48239,N_48396);
xor U48828 (N_48828,N_48149,N_48372);
and U48829 (N_48829,N_48325,N_48300);
or U48830 (N_48830,N_48150,N_48480);
and U48831 (N_48831,N_48058,N_48219);
or U48832 (N_48832,N_48038,N_48355);
nand U48833 (N_48833,N_48370,N_48052);
or U48834 (N_48834,N_48154,N_48136);
or U48835 (N_48835,N_48230,N_48027);
nand U48836 (N_48836,N_48368,N_48168);
or U48837 (N_48837,N_48408,N_48068);
nor U48838 (N_48838,N_48158,N_48071);
and U48839 (N_48839,N_48448,N_48405);
or U48840 (N_48840,N_48494,N_48182);
nand U48841 (N_48841,N_48447,N_48329);
or U48842 (N_48842,N_48398,N_48237);
nor U48843 (N_48843,N_48212,N_48039);
or U48844 (N_48844,N_48038,N_48130);
and U48845 (N_48845,N_48329,N_48397);
nand U48846 (N_48846,N_48251,N_48124);
nand U48847 (N_48847,N_48257,N_48057);
nor U48848 (N_48848,N_48417,N_48498);
xor U48849 (N_48849,N_48344,N_48372);
nand U48850 (N_48850,N_48124,N_48491);
xnor U48851 (N_48851,N_48264,N_48029);
nand U48852 (N_48852,N_48493,N_48215);
and U48853 (N_48853,N_48281,N_48082);
nand U48854 (N_48854,N_48464,N_48026);
nor U48855 (N_48855,N_48260,N_48383);
and U48856 (N_48856,N_48275,N_48353);
and U48857 (N_48857,N_48111,N_48155);
nand U48858 (N_48858,N_48195,N_48132);
xor U48859 (N_48859,N_48263,N_48250);
nor U48860 (N_48860,N_48110,N_48098);
or U48861 (N_48861,N_48419,N_48469);
and U48862 (N_48862,N_48203,N_48316);
or U48863 (N_48863,N_48468,N_48397);
xor U48864 (N_48864,N_48091,N_48475);
nand U48865 (N_48865,N_48300,N_48283);
nand U48866 (N_48866,N_48220,N_48445);
nand U48867 (N_48867,N_48395,N_48475);
xor U48868 (N_48868,N_48030,N_48386);
and U48869 (N_48869,N_48221,N_48433);
xor U48870 (N_48870,N_48228,N_48358);
nand U48871 (N_48871,N_48116,N_48168);
or U48872 (N_48872,N_48126,N_48176);
or U48873 (N_48873,N_48314,N_48332);
or U48874 (N_48874,N_48081,N_48101);
and U48875 (N_48875,N_48022,N_48131);
nand U48876 (N_48876,N_48071,N_48175);
nand U48877 (N_48877,N_48066,N_48224);
nand U48878 (N_48878,N_48017,N_48407);
nand U48879 (N_48879,N_48313,N_48288);
xnor U48880 (N_48880,N_48392,N_48159);
and U48881 (N_48881,N_48368,N_48462);
nor U48882 (N_48882,N_48381,N_48408);
or U48883 (N_48883,N_48044,N_48494);
or U48884 (N_48884,N_48144,N_48212);
nand U48885 (N_48885,N_48252,N_48490);
nand U48886 (N_48886,N_48030,N_48424);
nand U48887 (N_48887,N_48270,N_48432);
and U48888 (N_48888,N_48283,N_48424);
or U48889 (N_48889,N_48287,N_48291);
xor U48890 (N_48890,N_48186,N_48035);
nor U48891 (N_48891,N_48446,N_48035);
and U48892 (N_48892,N_48413,N_48385);
nand U48893 (N_48893,N_48191,N_48315);
nor U48894 (N_48894,N_48421,N_48230);
nand U48895 (N_48895,N_48200,N_48320);
nand U48896 (N_48896,N_48314,N_48369);
nand U48897 (N_48897,N_48369,N_48122);
nor U48898 (N_48898,N_48218,N_48406);
and U48899 (N_48899,N_48449,N_48000);
xor U48900 (N_48900,N_48122,N_48314);
or U48901 (N_48901,N_48151,N_48304);
or U48902 (N_48902,N_48126,N_48433);
nor U48903 (N_48903,N_48033,N_48213);
nand U48904 (N_48904,N_48468,N_48076);
xor U48905 (N_48905,N_48040,N_48433);
xnor U48906 (N_48906,N_48317,N_48223);
nand U48907 (N_48907,N_48353,N_48430);
nor U48908 (N_48908,N_48153,N_48303);
and U48909 (N_48909,N_48146,N_48154);
nor U48910 (N_48910,N_48085,N_48496);
and U48911 (N_48911,N_48280,N_48274);
and U48912 (N_48912,N_48298,N_48109);
nand U48913 (N_48913,N_48436,N_48496);
nor U48914 (N_48914,N_48458,N_48037);
or U48915 (N_48915,N_48000,N_48319);
nand U48916 (N_48916,N_48276,N_48068);
or U48917 (N_48917,N_48051,N_48358);
xnor U48918 (N_48918,N_48237,N_48087);
or U48919 (N_48919,N_48374,N_48284);
nor U48920 (N_48920,N_48165,N_48442);
or U48921 (N_48921,N_48268,N_48145);
nor U48922 (N_48922,N_48163,N_48362);
nor U48923 (N_48923,N_48292,N_48084);
or U48924 (N_48924,N_48373,N_48303);
nor U48925 (N_48925,N_48174,N_48423);
nand U48926 (N_48926,N_48357,N_48276);
and U48927 (N_48927,N_48135,N_48202);
xnor U48928 (N_48928,N_48249,N_48197);
nor U48929 (N_48929,N_48268,N_48316);
nor U48930 (N_48930,N_48207,N_48129);
and U48931 (N_48931,N_48461,N_48186);
or U48932 (N_48932,N_48361,N_48427);
nor U48933 (N_48933,N_48198,N_48299);
and U48934 (N_48934,N_48053,N_48458);
xor U48935 (N_48935,N_48155,N_48377);
nand U48936 (N_48936,N_48482,N_48256);
or U48937 (N_48937,N_48218,N_48307);
nand U48938 (N_48938,N_48353,N_48060);
xnor U48939 (N_48939,N_48419,N_48312);
or U48940 (N_48940,N_48329,N_48389);
nor U48941 (N_48941,N_48056,N_48125);
and U48942 (N_48942,N_48445,N_48229);
nand U48943 (N_48943,N_48325,N_48228);
or U48944 (N_48944,N_48265,N_48386);
xor U48945 (N_48945,N_48339,N_48289);
xnor U48946 (N_48946,N_48484,N_48381);
or U48947 (N_48947,N_48480,N_48157);
nand U48948 (N_48948,N_48153,N_48176);
xnor U48949 (N_48949,N_48170,N_48390);
nor U48950 (N_48950,N_48389,N_48049);
and U48951 (N_48951,N_48465,N_48007);
nor U48952 (N_48952,N_48368,N_48105);
nand U48953 (N_48953,N_48041,N_48387);
nor U48954 (N_48954,N_48121,N_48017);
xor U48955 (N_48955,N_48249,N_48303);
and U48956 (N_48956,N_48396,N_48474);
nor U48957 (N_48957,N_48326,N_48238);
nand U48958 (N_48958,N_48137,N_48152);
and U48959 (N_48959,N_48309,N_48353);
and U48960 (N_48960,N_48497,N_48083);
nand U48961 (N_48961,N_48395,N_48011);
or U48962 (N_48962,N_48167,N_48172);
or U48963 (N_48963,N_48149,N_48101);
or U48964 (N_48964,N_48075,N_48181);
nand U48965 (N_48965,N_48402,N_48049);
xnor U48966 (N_48966,N_48094,N_48194);
and U48967 (N_48967,N_48037,N_48418);
and U48968 (N_48968,N_48333,N_48327);
and U48969 (N_48969,N_48182,N_48243);
xor U48970 (N_48970,N_48422,N_48463);
nand U48971 (N_48971,N_48171,N_48099);
or U48972 (N_48972,N_48142,N_48372);
xnor U48973 (N_48973,N_48308,N_48263);
nor U48974 (N_48974,N_48009,N_48062);
xor U48975 (N_48975,N_48431,N_48321);
xnor U48976 (N_48976,N_48345,N_48382);
xnor U48977 (N_48977,N_48156,N_48292);
or U48978 (N_48978,N_48259,N_48275);
nor U48979 (N_48979,N_48442,N_48471);
and U48980 (N_48980,N_48027,N_48335);
xnor U48981 (N_48981,N_48164,N_48492);
or U48982 (N_48982,N_48342,N_48288);
xnor U48983 (N_48983,N_48432,N_48382);
xnor U48984 (N_48984,N_48145,N_48415);
or U48985 (N_48985,N_48284,N_48395);
or U48986 (N_48986,N_48404,N_48075);
nand U48987 (N_48987,N_48422,N_48482);
nor U48988 (N_48988,N_48239,N_48460);
nor U48989 (N_48989,N_48008,N_48486);
xnor U48990 (N_48990,N_48421,N_48449);
and U48991 (N_48991,N_48346,N_48031);
or U48992 (N_48992,N_48133,N_48256);
xnor U48993 (N_48993,N_48082,N_48006);
xor U48994 (N_48994,N_48354,N_48309);
and U48995 (N_48995,N_48079,N_48469);
nand U48996 (N_48996,N_48009,N_48072);
xnor U48997 (N_48997,N_48039,N_48274);
and U48998 (N_48998,N_48226,N_48355);
nand U48999 (N_48999,N_48157,N_48286);
nor U49000 (N_49000,N_48611,N_48994);
and U49001 (N_49001,N_48836,N_48515);
nor U49002 (N_49002,N_48901,N_48630);
nor U49003 (N_49003,N_48988,N_48724);
nand U49004 (N_49004,N_48944,N_48531);
xor U49005 (N_49005,N_48508,N_48550);
nor U49006 (N_49006,N_48799,N_48964);
xor U49007 (N_49007,N_48807,N_48601);
nand U49008 (N_49008,N_48652,N_48654);
or U49009 (N_49009,N_48942,N_48712);
and U49010 (N_49010,N_48998,N_48958);
nand U49011 (N_49011,N_48664,N_48810);
and U49012 (N_49012,N_48589,N_48603);
nand U49013 (N_49013,N_48697,N_48804);
and U49014 (N_49014,N_48681,N_48838);
and U49015 (N_49015,N_48731,N_48564);
nand U49016 (N_49016,N_48881,N_48797);
xor U49017 (N_49017,N_48686,N_48919);
and U49018 (N_49018,N_48955,N_48666);
nor U49019 (N_49019,N_48759,N_48661);
or U49020 (N_49020,N_48997,N_48925);
nand U49021 (N_49021,N_48619,N_48648);
xnor U49022 (N_49022,N_48678,N_48990);
nor U49023 (N_49023,N_48506,N_48667);
or U49024 (N_49024,N_48653,N_48704);
xor U49025 (N_49025,N_48702,N_48597);
nor U49026 (N_49026,N_48920,N_48915);
and U49027 (N_49027,N_48521,N_48628);
nor U49028 (N_49028,N_48764,N_48688);
xor U49029 (N_49029,N_48812,N_48636);
or U49030 (N_49030,N_48736,N_48852);
and U49031 (N_49031,N_48943,N_48763);
nand U49032 (N_49032,N_48670,N_48862);
or U49033 (N_49033,N_48594,N_48840);
nand U49034 (N_49034,N_48673,N_48675);
nor U49035 (N_49035,N_48959,N_48844);
nor U49036 (N_49036,N_48834,N_48888);
and U49037 (N_49037,N_48705,N_48741);
and U49038 (N_49038,N_48856,N_48726);
nor U49039 (N_49039,N_48947,N_48911);
and U49040 (N_49040,N_48534,N_48869);
nor U49041 (N_49041,N_48820,N_48608);
or U49042 (N_49042,N_48974,N_48950);
or U49043 (N_49043,N_48685,N_48918);
xor U49044 (N_49044,N_48742,N_48575);
nand U49045 (N_49045,N_48533,N_48596);
xor U49046 (N_49046,N_48641,N_48809);
and U49047 (N_49047,N_48817,N_48900);
nand U49048 (N_49048,N_48985,N_48937);
or U49049 (N_49049,N_48978,N_48766);
xnor U49050 (N_49050,N_48617,N_48793);
or U49051 (N_49051,N_48903,N_48595);
and U49052 (N_49052,N_48879,N_48584);
xnor U49053 (N_49053,N_48708,N_48863);
or U49054 (N_49054,N_48749,N_48948);
and U49055 (N_49055,N_48612,N_48677);
xnor U49056 (N_49056,N_48757,N_48668);
nor U49057 (N_49057,N_48634,N_48806);
xor U49058 (N_49058,N_48695,N_48605);
or U49059 (N_49059,N_48845,N_48982);
xnor U49060 (N_49060,N_48541,N_48819);
and U49061 (N_49061,N_48962,N_48588);
or U49062 (N_49062,N_48907,N_48660);
or U49063 (N_49063,N_48502,N_48853);
xnor U49064 (N_49064,N_48535,N_48859);
or U49065 (N_49065,N_48893,N_48582);
or U49066 (N_49066,N_48719,N_48934);
nor U49067 (N_49067,N_48583,N_48610);
xnor U49068 (N_49068,N_48837,N_48530);
nand U49069 (N_49069,N_48722,N_48623);
and U49070 (N_49070,N_48665,N_48880);
or U49071 (N_49071,N_48750,N_48684);
xor U49072 (N_49072,N_48885,N_48713);
or U49073 (N_49073,N_48663,N_48791);
or U49074 (N_49074,N_48646,N_48895);
xnor U49075 (N_49075,N_48536,N_48822);
and U49076 (N_49076,N_48910,N_48557);
xor U49077 (N_49077,N_48890,N_48926);
and U49078 (N_49078,N_48577,N_48587);
xnor U49079 (N_49079,N_48669,N_48560);
nor U49080 (N_49080,N_48546,N_48699);
or U49081 (N_49081,N_48821,N_48873);
nand U49082 (N_49082,N_48854,N_48633);
or U49083 (N_49083,N_48540,N_48656);
or U49084 (N_49084,N_48957,N_48929);
and U49085 (N_49085,N_48805,N_48867);
xor U49086 (N_49086,N_48831,N_48671);
xor U49087 (N_49087,N_48659,N_48643);
and U49088 (N_49088,N_48710,N_48874);
nand U49089 (N_49089,N_48725,N_48800);
and U49090 (N_49090,N_48839,N_48606);
or U49091 (N_49091,N_48701,N_48543);
or U49092 (N_49092,N_48861,N_48905);
nand U49093 (N_49093,N_48761,N_48753);
and U49094 (N_49094,N_48518,N_48878);
nor U49095 (N_49095,N_48832,N_48884);
xor U49096 (N_49096,N_48816,N_48877);
nand U49097 (N_49097,N_48609,N_48523);
xnor U49098 (N_49098,N_48931,N_48732);
or U49099 (N_49099,N_48991,N_48938);
xor U49100 (N_49100,N_48917,N_48871);
and U49101 (N_49101,N_48908,N_48566);
nand U49102 (N_49102,N_48813,N_48554);
xnor U49103 (N_49103,N_48751,N_48565);
and U49104 (N_49104,N_48754,N_48969);
nor U49105 (N_49105,N_48516,N_48717);
nand U49106 (N_49106,N_48904,N_48971);
nor U49107 (N_49107,N_48932,N_48616);
and U49108 (N_49108,N_48896,N_48585);
nor U49109 (N_49109,N_48841,N_48857);
nor U49110 (N_49110,N_48922,N_48872);
or U49111 (N_49111,N_48501,N_48735);
or U49112 (N_49112,N_48696,N_48966);
xnor U49113 (N_49113,N_48507,N_48892);
or U49114 (N_49114,N_48760,N_48963);
xor U49115 (N_49115,N_48563,N_48887);
xor U49116 (N_49116,N_48542,N_48614);
or U49117 (N_49117,N_48928,N_48548);
and U49118 (N_49118,N_48823,N_48782);
xnor U49119 (N_49119,N_48647,N_48714);
and U49120 (N_49120,N_48730,N_48644);
xor U49121 (N_49121,N_48989,N_48980);
nand U49122 (N_49122,N_48503,N_48939);
or U49123 (N_49123,N_48622,N_48711);
nor U49124 (N_49124,N_48776,N_48842);
or U49125 (N_49125,N_48627,N_48788);
nor U49126 (N_49126,N_48602,N_48522);
xnor U49127 (N_49127,N_48744,N_48626);
xor U49128 (N_49128,N_48851,N_48586);
nand U49129 (N_49129,N_48555,N_48707);
nand U49130 (N_49130,N_48723,N_48549);
nand U49131 (N_49131,N_48568,N_48970);
nor U49132 (N_49132,N_48818,N_48520);
xor U49133 (N_49133,N_48956,N_48519);
nand U49134 (N_49134,N_48784,N_48933);
nand U49135 (N_49135,N_48829,N_48987);
nand U49136 (N_49136,N_48651,N_48729);
nor U49137 (N_49137,N_48561,N_48815);
nand U49138 (N_49138,N_48796,N_48572);
xnor U49139 (N_49139,N_48936,N_48954);
nand U49140 (N_49140,N_48765,N_48870);
xor U49141 (N_49141,N_48960,N_48983);
and U49142 (N_49142,N_48849,N_48914);
nor U49143 (N_49143,N_48899,N_48514);
or U49144 (N_49144,N_48738,N_48591);
nand U49145 (N_49145,N_48858,N_48783);
or U49146 (N_49146,N_48968,N_48883);
nor U49147 (N_49147,N_48700,N_48683);
xor U49148 (N_49148,N_48930,N_48965);
nand U49149 (N_49149,N_48780,N_48935);
nor U49150 (N_49150,N_48547,N_48527);
and U49151 (N_49151,N_48777,N_48637);
or U49152 (N_49152,N_48803,N_48607);
nand U49153 (N_49153,N_48779,N_48740);
nand U49154 (N_49154,N_48544,N_48642);
xor U49155 (N_49155,N_48635,N_48752);
nand U49156 (N_49156,N_48655,N_48848);
and U49157 (N_49157,N_48762,N_48792);
xor U49158 (N_49158,N_48865,N_48785);
xnor U49159 (N_49159,N_48945,N_48747);
nand U49160 (N_49160,N_48986,N_48539);
xnor U49161 (N_49161,N_48794,N_48946);
nor U49162 (N_49162,N_48676,N_48500);
xor U49163 (N_49163,N_48787,N_48973);
or U49164 (N_49164,N_48625,N_48868);
nor U49165 (N_49165,N_48967,N_48802);
xnor U49166 (N_49166,N_48827,N_48524);
or U49167 (N_49167,N_48882,N_48620);
or U49168 (N_49168,N_48769,N_48748);
or U49169 (N_49169,N_48513,N_48758);
xnor U49170 (N_49170,N_48734,N_48579);
xnor U49171 (N_49171,N_48772,N_48739);
nand U49172 (N_49172,N_48941,N_48672);
xor U49173 (N_49173,N_48505,N_48774);
nand U49174 (N_49174,N_48662,N_48801);
nand U49175 (N_49175,N_48733,N_48613);
nor U49176 (N_49176,N_48771,N_48658);
nor U49177 (N_49177,N_48924,N_48592);
nand U49178 (N_49178,N_48961,N_48756);
or U49179 (N_49179,N_48814,N_48649);
nor U49180 (N_49180,N_48843,N_48570);
or U49181 (N_49181,N_48847,N_48745);
nor U49182 (N_49182,N_48808,N_48721);
nor U49183 (N_49183,N_48770,N_48599);
nand U49184 (N_49184,N_48786,N_48992);
nor U49185 (N_49185,N_48940,N_48909);
nand U49186 (N_49186,N_48835,N_48559);
nand U49187 (N_49187,N_48826,N_48993);
xor U49188 (N_49188,N_48682,N_48687);
xor U49189 (N_49189,N_48569,N_48604);
nand U49190 (N_49190,N_48906,N_48860);
nor U49191 (N_49191,N_48645,N_48889);
and U49192 (N_49192,N_48578,N_48538);
or U49193 (N_49193,N_48529,N_48876);
and U49194 (N_49194,N_48981,N_48545);
and U49195 (N_49195,N_48850,N_48718);
xor U49196 (N_49196,N_48979,N_48828);
or U49197 (N_49197,N_48715,N_48590);
nor U49198 (N_49198,N_48984,N_48698);
nor U49199 (N_49199,N_48833,N_48709);
or U49200 (N_49200,N_48875,N_48855);
and U49201 (N_49201,N_48825,N_48913);
nand U49202 (N_49202,N_48703,N_48621);
nor U49203 (N_49203,N_48511,N_48552);
nor U49204 (N_49204,N_48912,N_48693);
and U49205 (N_49205,N_48746,N_48689);
and U49206 (N_49206,N_48551,N_48571);
and U49207 (N_49207,N_48692,N_48830);
xnor U49208 (N_49208,N_48716,N_48999);
and U49209 (N_49209,N_48789,N_48574);
xor U49210 (N_49210,N_48562,N_48593);
nand U49211 (N_49211,N_48728,N_48640);
nor U49212 (N_49212,N_48706,N_48743);
nand U49213 (N_49213,N_48995,N_48674);
xor U49214 (N_49214,N_48512,N_48949);
nor U49215 (N_49215,N_48615,N_48775);
or U49216 (N_49216,N_48558,N_48894);
or U49217 (N_49217,N_48790,N_48629);
or U49218 (N_49218,N_48866,N_48532);
nor U49219 (N_49219,N_48510,N_48690);
or U49220 (N_49220,N_48755,N_48996);
and U49221 (N_49221,N_48504,N_48638);
nand U49222 (N_49222,N_48691,N_48581);
and U49223 (N_49223,N_48509,N_48916);
nand U49224 (N_49224,N_48650,N_48972);
and U49225 (N_49225,N_48580,N_48598);
nor U49226 (N_49226,N_48891,N_48567);
or U49227 (N_49227,N_48576,N_48727);
nand U49228 (N_49228,N_48526,N_48795);
xor U49229 (N_49229,N_48923,N_48952);
and U49230 (N_49230,N_48525,N_48767);
nor U49231 (N_49231,N_48773,N_48618);
xnor U49232 (N_49232,N_48657,N_48886);
xnor U49233 (N_49233,N_48927,N_48768);
nor U49234 (N_49234,N_48631,N_48573);
or U49235 (N_49235,N_48897,N_48977);
and U49236 (N_49236,N_48632,N_48953);
and U49237 (N_49237,N_48798,N_48556);
nand U49238 (N_49238,N_48537,N_48528);
and U49239 (N_49239,N_48720,N_48517);
xor U49240 (N_49240,N_48921,N_48824);
nand U49241 (N_49241,N_48679,N_48975);
nand U49242 (N_49242,N_48639,N_48624);
xor U49243 (N_49243,N_48902,N_48811);
and U49244 (N_49244,N_48778,N_48680);
or U49245 (N_49245,N_48781,N_48898);
or U49246 (N_49246,N_48951,N_48976);
nand U49247 (N_49247,N_48553,N_48694);
nor U49248 (N_49248,N_48864,N_48737);
or U49249 (N_49249,N_48846,N_48600);
or U49250 (N_49250,N_48741,N_48825);
nor U49251 (N_49251,N_48998,N_48716);
nor U49252 (N_49252,N_48649,N_48981);
nor U49253 (N_49253,N_48524,N_48862);
nor U49254 (N_49254,N_48973,N_48922);
xor U49255 (N_49255,N_48949,N_48553);
nor U49256 (N_49256,N_48779,N_48775);
xor U49257 (N_49257,N_48749,N_48673);
and U49258 (N_49258,N_48882,N_48777);
nor U49259 (N_49259,N_48648,N_48867);
and U49260 (N_49260,N_48884,N_48913);
or U49261 (N_49261,N_48916,N_48776);
and U49262 (N_49262,N_48959,N_48768);
and U49263 (N_49263,N_48719,N_48920);
and U49264 (N_49264,N_48966,N_48984);
nand U49265 (N_49265,N_48725,N_48759);
nor U49266 (N_49266,N_48566,N_48780);
xnor U49267 (N_49267,N_48661,N_48652);
or U49268 (N_49268,N_48886,N_48604);
xnor U49269 (N_49269,N_48651,N_48795);
or U49270 (N_49270,N_48807,N_48685);
or U49271 (N_49271,N_48869,N_48796);
xor U49272 (N_49272,N_48871,N_48676);
xor U49273 (N_49273,N_48883,N_48609);
and U49274 (N_49274,N_48981,N_48988);
xor U49275 (N_49275,N_48713,N_48817);
or U49276 (N_49276,N_48990,N_48873);
xnor U49277 (N_49277,N_48987,N_48839);
or U49278 (N_49278,N_48690,N_48954);
and U49279 (N_49279,N_48696,N_48599);
nand U49280 (N_49280,N_48534,N_48807);
xnor U49281 (N_49281,N_48839,N_48911);
xor U49282 (N_49282,N_48819,N_48747);
nor U49283 (N_49283,N_48788,N_48849);
and U49284 (N_49284,N_48810,N_48788);
nor U49285 (N_49285,N_48895,N_48645);
nor U49286 (N_49286,N_48831,N_48935);
nand U49287 (N_49287,N_48994,N_48685);
xor U49288 (N_49288,N_48880,N_48779);
and U49289 (N_49289,N_48783,N_48536);
or U49290 (N_49290,N_48828,N_48535);
and U49291 (N_49291,N_48963,N_48843);
nand U49292 (N_49292,N_48666,N_48710);
and U49293 (N_49293,N_48615,N_48640);
nand U49294 (N_49294,N_48645,N_48587);
and U49295 (N_49295,N_48731,N_48710);
nor U49296 (N_49296,N_48561,N_48947);
or U49297 (N_49297,N_48535,N_48847);
xor U49298 (N_49298,N_48960,N_48749);
nor U49299 (N_49299,N_48626,N_48779);
and U49300 (N_49300,N_48628,N_48877);
nand U49301 (N_49301,N_48832,N_48743);
xor U49302 (N_49302,N_48969,N_48848);
and U49303 (N_49303,N_48762,N_48679);
nand U49304 (N_49304,N_48823,N_48856);
or U49305 (N_49305,N_48528,N_48513);
and U49306 (N_49306,N_48656,N_48808);
or U49307 (N_49307,N_48865,N_48812);
nand U49308 (N_49308,N_48552,N_48641);
and U49309 (N_49309,N_48771,N_48881);
xor U49310 (N_49310,N_48817,N_48970);
xor U49311 (N_49311,N_48854,N_48614);
or U49312 (N_49312,N_48814,N_48867);
or U49313 (N_49313,N_48991,N_48921);
and U49314 (N_49314,N_48568,N_48914);
xnor U49315 (N_49315,N_48733,N_48804);
nor U49316 (N_49316,N_48591,N_48736);
or U49317 (N_49317,N_48752,N_48986);
nor U49318 (N_49318,N_48620,N_48702);
and U49319 (N_49319,N_48895,N_48816);
nand U49320 (N_49320,N_48924,N_48578);
xnor U49321 (N_49321,N_48934,N_48616);
nor U49322 (N_49322,N_48623,N_48654);
nor U49323 (N_49323,N_48575,N_48603);
nand U49324 (N_49324,N_48897,N_48543);
or U49325 (N_49325,N_48776,N_48682);
nor U49326 (N_49326,N_48544,N_48860);
nand U49327 (N_49327,N_48837,N_48528);
nor U49328 (N_49328,N_48637,N_48968);
nand U49329 (N_49329,N_48779,N_48523);
and U49330 (N_49330,N_48646,N_48887);
or U49331 (N_49331,N_48548,N_48659);
and U49332 (N_49332,N_48928,N_48604);
and U49333 (N_49333,N_48598,N_48968);
nand U49334 (N_49334,N_48798,N_48520);
and U49335 (N_49335,N_48777,N_48929);
or U49336 (N_49336,N_48797,N_48874);
and U49337 (N_49337,N_48659,N_48957);
or U49338 (N_49338,N_48743,N_48858);
nand U49339 (N_49339,N_48532,N_48991);
nor U49340 (N_49340,N_48930,N_48704);
xor U49341 (N_49341,N_48624,N_48562);
xnor U49342 (N_49342,N_48838,N_48564);
xor U49343 (N_49343,N_48512,N_48889);
or U49344 (N_49344,N_48792,N_48843);
or U49345 (N_49345,N_48990,N_48612);
and U49346 (N_49346,N_48595,N_48643);
and U49347 (N_49347,N_48822,N_48626);
nand U49348 (N_49348,N_48807,N_48869);
xnor U49349 (N_49349,N_48957,N_48741);
and U49350 (N_49350,N_48933,N_48591);
or U49351 (N_49351,N_48612,N_48577);
nand U49352 (N_49352,N_48796,N_48646);
and U49353 (N_49353,N_48874,N_48546);
nand U49354 (N_49354,N_48861,N_48891);
nand U49355 (N_49355,N_48940,N_48858);
nor U49356 (N_49356,N_48692,N_48949);
xnor U49357 (N_49357,N_48732,N_48616);
or U49358 (N_49358,N_48593,N_48841);
nor U49359 (N_49359,N_48636,N_48510);
nor U49360 (N_49360,N_48639,N_48679);
nand U49361 (N_49361,N_48982,N_48670);
xnor U49362 (N_49362,N_48710,N_48579);
xor U49363 (N_49363,N_48546,N_48711);
nor U49364 (N_49364,N_48779,N_48716);
xnor U49365 (N_49365,N_48984,N_48757);
and U49366 (N_49366,N_48772,N_48749);
xor U49367 (N_49367,N_48661,N_48862);
nor U49368 (N_49368,N_48758,N_48563);
xnor U49369 (N_49369,N_48789,N_48544);
nor U49370 (N_49370,N_48842,N_48637);
nor U49371 (N_49371,N_48917,N_48831);
xnor U49372 (N_49372,N_48984,N_48866);
and U49373 (N_49373,N_48819,N_48754);
xor U49374 (N_49374,N_48564,N_48535);
and U49375 (N_49375,N_48768,N_48666);
xor U49376 (N_49376,N_48552,N_48933);
nand U49377 (N_49377,N_48934,N_48649);
xor U49378 (N_49378,N_48622,N_48526);
and U49379 (N_49379,N_48835,N_48512);
nor U49380 (N_49380,N_48935,N_48958);
or U49381 (N_49381,N_48911,N_48927);
nand U49382 (N_49382,N_48519,N_48803);
xnor U49383 (N_49383,N_48890,N_48616);
xnor U49384 (N_49384,N_48840,N_48612);
nor U49385 (N_49385,N_48689,N_48822);
nand U49386 (N_49386,N_48931,N_48542);
nand U49387 (N_49387,N_48618,N_48617);
or U49388 (N_49388,N_48705,N_48823);
and U49389 (N_49389,N_48767,N_48621);
nor U49390 (N_49390,N_48643,N_48887);
xnor U49391 (N_49391,N_48510,N_48823);
and U49392 (N_49392,N_48896,N_48622);
nand U49393 (N_49393,N_48574,N_48817);
or U49394 (N_49394,N_48987,N_48891);
nor U49395 (N_49395,N_48755,N_48912);
nand U49396 (N_49396,N_48862,N_48965);
or U49397 (N_49397,N_48677,N_48516);
nand U49398 (N_49398,N_48643,N_48539);
nand U49399 (N_49399,N_48849,N_48839);
nand U49400 (N_49400,N_48722,N_48552);
or U49401 (N_49401,N_48603,N_48582);
nor U49402 (N_49402,N_48576,N_48664);
or U49403 (N_49403,N_48808,N_48720);
nand U49404 (N_49404,N_48659,N_48791);
or U49405 (N_49405,N_48922,N_48896);
and U49406 (N_49406,N_48935,N_48537);
nand U49407 (N_49407,N_48599,N_48564);
and U49408 (N_49408,N_48641,N_48654);
nand U49409 (N_49409,N_48865,N_48671);
nor U49410 (N_49410,N_48818,N_48896);
nor U49411 (N_49411,N_48801,N_48921);
and U49412 (N_49412,N_48834,N_48627);
and U49413 (N_49413,N_48514,N_48864);
nand U49414 (N_49414,N_48733,N_48521);
and U49415 (N_49415,N_48611,N_48768);
or U49416 (N_49416,N_48545,N_48697);
xor U49417 (N_49417,N_48921,N_48988);
nand U49418 (N_49418,N_48957,N_48951);
nor U49419 (N_49419,N_48735,N_48568);
nor U49420 (N_49420,N_48718,N_48948);
or U49421 (N_49421,N_48613,N_48788);
and U49422 (N_49422,N_48587,N_48963);
nand U49423 (N_49423,N_48706,N_48510);
nor U49424 (N_49424,N_48804,N_48819);
xnor U49425 (N_49425,N_48799,N_48996);
xnor U49426 (N_49426,N_48973,N_48717);
nor U49427 (N_49427,N_48900,N_48826);
or U49428 (N_49428,N_48723,N_48976);
or U49429 (N_49429,N_48626,N_48998);
and U49430 (N_49430,N_48971,N_48876);
nor U49431 (N_49431,N_48689,N_48638);
and U49432 (N_49432,N_48692,N_48530);
and U49433 (N_49433,N_48712,N_48868);
nor U49434 (N_49434,N_48849,N_48730);
nand U49435 (N_49435,N_48739,N_48514);
or U49436 (N_49436,N_48564,N_48850);
and U49437 (N_49437,N_48833,N_48844);
xor U49438 (N_49438,N_48738,N_48773);
nor U49439 (N_49439,N_48824,N_48792);
nor U49440 (N_49440,N_48564,N_48763);
xor U49441 (N_49441,N_48979,N_48567);
or U49442 (N_49442,N_48541,N_48813);
or U49443 (N_49443,N_48747,N_48852);
xor U49444 (N_49444,N_48593,N_48738);
or U49445 (N_49445,N_48870,N_48619);
nand U49446 (N_49446,N_48588,N_48790);
nand U49447 (N_49447,N_48798,N_48764);
nand U49448 (N_49448,N_48897,N_48659);
nand U49449 (N_49449,N_48705,N_48764);
xnor U49450 (N_49450,N_48558,N_48857);
nor U49451 (N_49451,N_48866,N_48646);
nor U49452 (N_49452,N_48884,N_48608);
or U49453 (N_49453,N_48862,N_48514);
and U49454 (N_49454,N_48571,N_48615);
xor U49455 (N_49455,N_48959,N_48612);
nand U49456 (N_49456,N_48776,N_48860);
nor U49457 (N_49457,N_48731,N_48942);
and U49458 (N_49458,N_48733,N_48882);
xnor U49459 (N_49459,N_48775,N_48924);
and U49460 (N_49460,N_48732,N_48651);
and U49461 (N_49461,N_48673,N_48795);
and U49462 (N_49462,N_48789,N_48836);
or U49463 (N_49463,N_48694,N_48545);
nor U49464 (N_49464,N_48792,N_48544);
nor U49465 (N_49465,N_48956,N_48743);
xor U49466 (N_49466,N_48694,N_48560);
nand U49467 (N_49467,N_48837,N_48701);
and U49468 (N_49468,N_48638,N_48644);
nand U49469 (N_49469,N_48541,N_48970);
and U49470 (N_49470,N_48629,N_48558);
xnor U49471 (N_49471,N_48512,N_48623);
nand U49472 (N_49472,N_48847,N_48765);
or U49473 (N_49473,N_48864,N_48835);
nand U49474 (N_49474,N_48979,N_48683);
or U49475 (N_49475,N_48789,N_48838);
or U49476 (N_49476,N_48644,N_48784);
or U49477 (N_49477,N_48820,N_48984);
nor U49478 (N_49478,N_48888,N_48581);
and U49479 (N_49479,N_48621,N_48776);
or U49480 (N_49480,N_48796,N_48611);
and U49481 (N_49481,N_48831,N_48903);
nor U49482 (N_49482,N_48687,N_48644);
or U49483 (N_49483,N_48605,N_48744);
nor U49484 (N_49484,N_48881,N_48988);
nand U49485 (N_49485,N_48956,N_48808);
and U49486 (N_49486,N_48743,N_48964);
nor U49487 (N_49487,N_48566,N_48910);
xnor U49488 (N_49488,N_48837,N_48551);
nor U49489 (N_49489,N_48649,N_48568);
nand U49490 (N_49490,N_48558,N_48502);
nand U49491 (N_49491,N_48707,N_48913);
xnor U49492 (N_49492,N_48867,N_48641);
xnor U49493 (N_49493,N_48540,N_48722);
and U49494 (N_49494,N_48861,N_48991);
or U49495 (N_49495,N_48806,N_48598);
nand U49496 (N_49496,N_48791,N_48762);
xnor U49497 (N_49497,N_48643,N_48583);
xor U49498 (N_49498,N_48843,N_48824);
nor U49499 (N_49499,N_48809,N_48763);
nor U49500 (N_49500,N_49107,N_49072);
nor U49501 (N_49501,N_49446,N_49362);
nand U49502 (N_49502,N_49332,N_49337);
or U49503 (N_49503,N_49472,N_49271);
or U49504 (N_49504,N_49244,N_49343);
or U49505 (N_49505,N_49402,N_49160);
and U49506 (N_49506,N_49350,N_49341);
nand U49507 (N_49507,N_49404,N_49322);
nand U49508 (N_49508,N_49193,N_49159);
nor U49509 (N_49509,N_49222,N_49098);
nand U49510 (N_49510,N_49182,N_49038);
or U49511 (N_49511,N_49099,N_49260);
and U49512 (N_49512,N_49073,N_49401);
nor U49513 (N_49513,N_49115,N_49128);
and U49514 (N_49514,N_49228,N_49342);
nand U49515 (N_49515,N_49375,N_49241);
xnor U49516 (N_49516,N_49360,N_49328);
and U49517 (N_49517,N_49023,N_49434);
and U49518 (N_49518,N_49424,N_49289);
and U49519 (N_49519,N_49443,N_49188);
nand U49520 (N_49520,N_49365,N_49378);
and U49521 (N_49521,N_49339,N_49471);
xor U49522 (N_49522,N_49161,N_49207);
nor U49523 (N_49523,N_49213,N_49199);
nor U49524 (N_49524,N_49211,N_49103);
or U49525 (N_49525,N_49309,N_49052);
or U49526 (N_49526,N_49467,N_49022);
nand U49527 (N_49527,N_49284,N_49438);
or U49528 (N_49528,N_49266,N_49409);
nand U49529 (N_49529,N_49297,N_49283);
nor U49530 (N_49530,N_49212,N_49081);
nor U49531 (N_49531,N_49123,N_49089);
or U49532 (N_49532,N_49315,N_49245);
xor U49533 (N_49533,N_49435,N_49408);
nand U49534 (N_49534,N_49361,N_49410);
xnor U49535 (N_49535,N_49096,N_49058);
nor U49536 (N_49536,N_49464,N_49479);
and U49537 (N_49537,N_49458,N_49238);
nor U49538 (N_49538,N_49195,N_49324);
nor U49539 (N_49539,N_49333,N_49302);
nand U49540 (N_49540,N_49033,N_49168);
or U49541 (N_49541,N_49304,N_49247);
and U49542 (N_49542,N_49000,N_49327);
xnor U49543 (N_49543,N_49173,N_49153);
and U49544 (N_49544,N_49232,N_49396);
nor U49545 (N_49545,N_49053,N_49192);
and U49546 (N_49546,N_49412,N_49138);
xor U49547 (N_49547,N_49068,N_49205);
xnor U49548 (N_49548,N_49445,N_49061);
and U49549 (N_49549,N_49394,N_49456);
and U49550 (N_49550,N_49013,N_49063);
and U49551 (N_49551,N_49385,N_49383);
and U49552 (N_49552,N_49219,N_49301);
nand U49553 (N_49553,N_49175,N_49494);
nor U49554 (N_49554,N_49248,N_49169);
nand U49555 (N_49555,N_49012,N_49497);
or U49556 (N_49556,N_49118,N_49320);
nand U49557 (N_49557,N_49144,N_49425);
or U49558 (N_49558,N_49203,N_49393);
or U49559 (N_49559,N_49495,N_49157);
xor U49560 (N_49560,N_49079,N_49119);
nand U49561 (N_49561,N_49489,N_49121);
nor U49562 (N_49562,N_49214,N_49487);
nor U49563 (N_49563,N_49194,N_49481);
xor U49564 (N_49564,N_49427,N_49454);
nand U49565 (N_49565,N_49016,N_49218);
and U49566 (N_49566,N_49368,N_49091);
xor U49567 (N_49567,N_49312,N_49116);
xnor U49568 (N_49568,N_49384,N_49178);
and U49569 (N_49569,N_49136,N_49109);
or U49570 (N_49570,N_49190,N_49496);
nor U49571 (N_49571,N_49331,N_49014);
xor U49572 (N_49572,N_49269,N_49132);
xor U49573 (N_49573,N_49423,N_49381);
xnor U49574 (N_49574,N_49223,N_49449);
nor U49575 (N_49575,N_49416,N_49480);
or U49576 (N_49576,N_49366,N_49330);
and U49577 (N_49577,N_49010,N_49236);
xor U49578 (N_49578,N_49256,N_49251);
nor U49579 (N_49579,N_49032,N_49083);
nand U49580 (N_49580,N_49078,N_49407);
nand U49581 (N_49581,N_49235,N_49198);
xor U49582 (N_49582,N_49286,N_49146);
nand U49583 (N_49583,N_49162,N_49314);
and U49584 (N_49584,N_49059,N_49352);
nand U49585 (N_49585,N_49265,N_49197);
or U49586 (N_49586,N_49444,N_49268);
or U49587 (N_49587,N_49498,N_49370);
nand U49588 (N_49588,N_49104,N_49097);
or U49589 (N_49589,N_49359,N_49143);
xor U49590 (N_49590,N_49376,N_49149);
and U49591 (N_49591,N_49379,N_49036);
and U49592 (N_49592,N_49240,N_49246);
nor U49593 (N_49593,N_49015,N_49221);
xnor U49594 (N_49594,N_49201,N_49448);
nor U49595 (N_49595,N_49447,N_49374);
and U49596 (N_49596,N_49291,N_49024);
nor U49597 (N_49597,N_49007,N_49349);
or U49598 (N_49598,N_49413,N_49432);
xnor U49599 (N_49599,N_49442,N_49461);
or U49600 (N_49600,N_49187,N_49317);
xnor U49601 (N_49601,N_49165,N_49278);
nand U49602 (N_49602,N_49484,N_49272);
nor U49603 (N_49603,N_49049,N_49209);
and U49604 (N_49604,N_49348,N_49156);
nand U49605 (N_49605,N_49029,N_49474);
and U49606 (N_49606,N_49344,N_49074);
or U49607 (N_49607,N_49397,N_49428);
and U49608 (N_49608,N_49263,N_49371);
nand U49609 (N_49609,N_49180,N_49280);
nand U49610 (N_49610,N_49421,N_49418);
nand U49611 (N_49611,N_49369,N_49230);
xnor U49612 (N_49612,N_49492,N_49056);
xor U49613 (N_49613,N_49047,N_49380);
and U49614 (N_49614,N_49057,N_49183);
nand U49615 (N_49615,N_49112,N_49135);
and U49616 (N_49616,N_49430,N_49486);
and U49617 (N_49617,N_49050,N_49101);
xnor U49618 (N_49618,N_49395,N_49100);
xnor U49619 (N_49619,N_49319,N_49224);
or U49620 (N_49620,N_49372,N_49318);
and U49621 (N_49621,N_49028,N_49220);
and U49622 (N_49622,N_49389,N_49436);
nand U49623 (N_49623,N_49499,N_49026);
or U49624 (N_49624,N_49206,N_49133);
nor U49625 (N_49625,N_49329,N_49094);
nor U49626 (N_49626,N_49273,N_49176);
nand U49627 (N_49627,N_49400,N_49483);
or U49628 (N_49628,N_49358,N_49117);
nand U49629 (N_49629,N_49035,N_49229);
or U49630 (N_49630,N_49031,N_49090);
nor U49631 (N_49631,N_49001,N_49452);
xor U49632 (N_49632,N_49282,N_49264);
or U49633 (N_49633,N_49186,N_49255);
and U49634 (N_49634,N_49477,N_49253);
nand U49635 (N_49635,N_49279,N_49155);
nor U49636 (N_49636,N_49170,N_49150);
or U49637 (N_49637,N_49285,N_49124);
or U49638 (N_49638,N_49105,N_49457);
and U49639 (N_49639,N_49310,N_49179);
or U49640 (N_49640,N_49114,N_49335);
nand U49641 (N_49641,N_49391,N_49488);
or U49642 (N_49642,N_49377,N_49305);
nand U49643 (N_49643,N_49345,N_49478);
and U49644 (N_49644,N_49233,N_49463);
and U49645 (N_49645,N_49390,N_49415);
nand U49646 (N_49646,N_49111,N_49152);
and U49647 (N_49647,N_49102,N_49465);
xnor U49648 (N_49648,N_49429,N_49355);
nand U49649 (N_49649,N_49171,N_49051);
nor U49650 (N_49650,N_49411,N_49473);
xor U49651 (N_49651,N_49039,N_49356);
nor U49652 (N_49652,N_49046,N_49225);
or U49653 (N_49653,N_49076,N_49354);
nor U49654 (N_49654,N_49011,N_49267);
xnor U49655 (N_49655,N_49326,N_49237);
xnor U49656 (N_49656,N_49060,N_49130);
nor U49657 (N_49657,N_49226,N_49299);
xor U49658 (N_49658,N_49154,N_49070);
or U49659 (N_49659,N_49249,N_49419);
nor U49660 (N_49660,N_49466,N_49462);
or U49661 (N_49661,N_49387,N_49294);
and U49662 (N_49662,N_49274,N_49093);
and U49663 (N_49663,N_49202,N_49303);
and U49664 (N_49664,N_49367,N_49134);
xor U49665 (N_49665,N_49009,N_49295);
nor U49666 (N_49666,N_49234,N_49306);
nor U49667 (N_49667,N_49002,N_49262);
nand U49668 (N_49668,N_49084,N_49043);
or U49669 (N_49669,N_49086,N_49298);
nand U49670 (N_49670,N_49145,N_49441);
nor U49671 (N_49671,N_49064,N_49040);
and U49672 (N_49672,N_49313,N_49300);
xor U49673 (N_49673,N_49021,N_49125);
xor U49674 (N_49674,N_49087,N_49216);
xor U49675 (N_49675,N_49276,N_49281);
and U49676 (N_49676,N_49200,N_49177);
nand U49677 (N_49677,N_49351,N_49363);
nand U49678 (N_49678,N_49293,N_49215);
and U49679 (N_49679,N_49257,N_49082);
nor U49680 (N_49680,N_49403,N_49185);
and U49681 (N_49681,N_49045,N_49325);
and U49682 (N_49682,N_49414,N_49485);
nor U49683 (N_49683,N_49316,N_49034);
nor U49684 (N_49684,N_49227,N_49288);
nor U49685 (N_49685,N_49077,N_49048);
nor U49686 (N_49686,N_49455,N_49392);
xor U49687 (N_49687,N_49364,N_49174);
nand U49688 (N_49688,N_49044,N_49426);
nand U49689 (N_49689,N_49018,N_49440);
or U49690 (N_49690,N_49431,N_49406);
nand U49691 (N_49691,N_49482,N_49296);
and U49692 (N_49692,N_49321,N_49353);
and U49693 (N_49693,N_49095,N_49191);
nor U49694 (N_49694,N_49042,N_49181);
and U49695 (N_49695,N_49164,N_49490);
nand U49696 (N_49696,N_49250,N_49292);
and U49697 (N_49697,N_49308,N_49261);
nor U49698 (N_49698,N_49270,N_49166);
xor U49699 (N_49699,N_49338,N_49122);
and U49700 (N_49700,N_49126,N_49252);
or U49701 (N_49701,N_49439,N_49451);
nor U49702 (N_49702,N_49141,N_49311);
xor U49703 (N_49703,N_49357,N_49459);
or U49704 (N_49704,N_49258,N_49493);
xnor U49705 (N_49705,N_49460,N_49437);
xor U49706 (N_49706,N_49172,N_49139);
xnor U49707 (N_49707,N_49468,N_49373);
nand U49708 (N_49708,N_49347,N_49037);
nand U49709 (N_49709,N_49275,N_49204);
xnor U49710 (N_49710,N_49336,N_49080);
and U49711 (N_49711,N_49388,N_49067);
or U49712 (N_49712,N_49108,N_49287);
and U49713 (N_49713,N_49417,N_49398);
nand U49714 (N_49714,N_49054,N_49450);
nand U49715 (N_49715,N_49005,N_49140);
and U49716 (N_49716,N_49243,N_49003);
nor U49717 (N_49717,N_49137,N_49231);
and U49718 (N_49718,N_49346,N_49340);
nand U49719 (N_49719,N_49004,N_49113);
nor U49720 (N_49720,N_49131,N_49092);
nand U49721 (N_49721,N_49167,N_49055);
nand U49722 (N_49722,N_49420,N_49163);
nand U49723 (N_49723,N_49158,N_49189);
xnor U49724 (N_49724,N_49062,N_49151);
nand U49725 (N_49725,N_49020,N_49242);
xnor U49726 (N_49726,N_49085,N_49307);
nand U49727 (N_49727,N_49386,N_49142);
and U49728 (N_49728,N_49127,N_49476);
nor U49729 (N_49729,N_49382,N_49071);
nor U49730 (N_49730,N_49041,N_49106);
xnor U49731 (N_49731,N_49066,N_49491);
nand U49732 (N_49732,N_49129,N_49277);
or U49733 (N_49733,N_49323,N_49184);
nand U49734 (N_49734,N_49075,N_49069);
or U49735 (N_49735,N_49008,N_49208);
or U49736 (N_49736,N_49334,N_49469);
and U49737 (N_49737,N_49239,N_49290);
nand U49738 (N_49738,N_49017,N_49110);
nand U49739 (N_49739,N_49217,N_49433);
nor U49740 (N_49740,N_49470,N_49065);
xor U49741 (N_49741,N_49088,N_49210);
or U49742 (N_49742,N_49405,N_49019);
and U49743 (N_49743,N_49399,N_49148);
xor U49744 (N_49744,N_49475,N_49254);
xnor U49745 (N_49745,N_49030,N_49196);
nand U49746 (N_49746,N_49259,N_49147);
xor U49747 (N_49747,N_49025,N_49006);
nor U49748 (N_49748,N_49453,N_49027);
or U49749 (N_49749,N_49422,N_49120);
nand U49750 (N_49750,N_49381,N_49087);
xnor U49751 (N_49751,N_49208,N_49339);
or U49752 (N_49752,N_49346,N_49055);
xor U49753 (N_49753,N_49409,N_49233);
xor U49754 (N_49754,N_49253,N_49462);
nand U49755 (N_49755,N_49122,N_49392);
xor U49756 (N_49756,N_49192,N_49004);
xnor U49757 (N_49757,N_49276,N_49268);
xnor U49758 (N_49758,N_49307,N_49211);
nand U49759 (N_49759,N_49011,N_49033);
nand U49760 (N_49760,N_49147,N_49333);
xor U49761 (N_49761,N_49288,N_49172);
or U49762 (N_49762,N_49239,N_49195);
xor U49763 (N_49763,N_49032,N_49040);
or U49764 (N_49764,N_49265,N_49103);
nor U49765 (N_49765,N_49051,N_49337);
or U49766 (N_49766,N_49471,N_49131);
nand U49767 (N_49767,N_49348,N_49023);
and U49768 (N_49768,N_49381,N_49048);
xor U49769 (N_49769,N_49451,N_49335);
and U49770 (N_49770,N_49240,N_49095);
xor U49771 (N_49771,N_49414,N_49001);
or U49772 (N_49772,N_49328,N_49377);
xnor U49773 (N_49773,N_49443,N_49477);
xnor U49774 (N_49774,N_49028,N_49146);
or U49775 (N_49775,N_49439,N_49052);
nand U49776 (N_49776,N_49190,N_49346);
nor U49777 (N_49777,N_49269,N_49012);
nand U49778 (N_49778,N_49020,N_49414);
nor U49779 (N_49779,N_49429,N_49476);
and U49780 (N_49780,N_49471,N_49159);
or U49781 (N_49781,N_49032,N_49221);
or U49782 (N_49782,N_49135,N_49475);
xor U49783 (N_49783,N_49107,N_49033);
and U49784 (N_49784,N_49437,N_49422);
nand U49785 (N_49785,N_49313,N_49334);
nand U49786 (N_49786,N_49215,N_49452);
and U49787 (N_49787,N_49442,N_49177);
nor U49788 (N_49788,N_49134,N_49162);
and U49789 (N_49789,N_49266,N_49487);
nand U49790 (N_49790,N_49212,N_49450);
xnor U49791 (N_49791,N_49004,N_49136);
or U49792 (N_49792,N_49147,N_49311);
or U49793 (N_49793,N_49109,N_49130);
xnor U49794 (N_49794,N_49389,N_49115);
and U49795 (N_49795,N_49458,N_49164);
nand U49796 (N_49796,N_49289,N_49074);
or U49797 (N_49797,N_49122,N_49450);
nand U49798 (N_49798,N_49467,N_49354);
and U49799 (N_49799,N_49040,N_49403);
xor U49800 (N_49800,N_49480,N_49031);
xor U49801 (N_49801,N_49115,N_49099);
or U49802 (N_49802,N_49457,N_49005);
and U49803 (N_49803,N_49391,N_49115);
and U49804 (N_49804,N_49448,N_49410);
or U49805 (N_49805,N_49064,N_49102);
or U49806 (N_49806,N_49404,N_49021);
or U49807 (N_49807,N_49301,N_49485);
xor U49808 (N_49808,N_49372,N_49294);
xor U49809 (N_49809,N_49359,N_49179);
nand U49810 (N_49810,N_49467,N_49438);
xnor U49811 (N_49811,N_49200,N_49180);
xor U49812 (N_49812,N_49061,N_49163);
nor U49813 (N_49813,N_49020,N_49435);
nand U49814 (N_49814,N_49423,N_49061);
nor U49815 (N_49815,N_49018,N_49344);
and U49816 (N_49816,N_49089,N_49331);
and U49817 (N_49817,N_49321,N_49222);
or U49818 (N_49818,N_49063,N_49135);
or U49819 (N_49819,N_49430,N_49269);
and U49820 (N_49820,N_49397,N_49028);
xnor U49821 (N_49821,N_49289,N_49277);
or U49822 (N_49822,N_49436,N_49482);
nor U49823 (N_49823,N_49156,N_49024);
and U49824 (N_49824,N_49074,N_49181);
xor U49825 (N_49825,N_49299,N_49447);
xor U49826 (N_49826,N_49215,N_49032);
and U49827 (N_49827,N_49203,N_49310);
xnor U49828 (N_49828,N_49429,N_49251);
nor U49829 (N_49829,N_49383,N_49276);
and U49830 (N_49830,N_49052,N_49212);
nor U49831 (N_49831,N_49287,N_49414);
nand U49832 (N_49832,N_49276,N_49279);
nand U49833 (N_49833,N_49370,N_49458);
nor U49834 (N_49834,N_49459,N_49262);
or U49835 (N_49835,N_49326,N_49209);
or U49836 (N_49836,N_49036,N_49201);
or U49837 (N_49837,N_49254,N_49409);
nand U49838 (N_49838,N_49457,N_49332);
or U49839 (N_49839,N_49252,N_49323);
nor U49840 (N_49840,N_49171,N_49036);
nand U49841 (N_49841,N_49146,N_49388);
and U49842 (N_49842,N_49204,N_49017);
and U49843 (N_49843,N_49178,N_49187);
xnor U49844 (N_49844,N_49152,N_49147);
nor U49845 (N_49845,N_49309,N_49289);
or U49846 (N_49846,N_49240,N_49107);
and U49847 (N_49847,N_49010,N_49167);
xnor U49848 (N_49848,N_49402,N_49244);
and U49849 (N_49849,N_49361,N_49023);
or U49850 (N_49850,N_49087,N_49208);
nand U49851 (N_49851,N_49390,N_49103);
or U49852 (N_49852,N_49318,N_49196);
xor U49853 (N_49853,N_49184,N_49320);
and U49854 (N_49854,N_49084,N_49262);
or U49855 (N_49855,N_49061,N_49213);
and U49856 (N_49856,N_49070,N_49419);
or U49857 (N_49857,N_49065,N_49426);
nand U49858 (N_49858,N_49440,N_49146);
nand U49859 (N_49859,N_49031,N_49332);
and U49860 (N_49860,N_49204,N_49240);
and U49861 (N_49861,N_49057,N_49234);
xnor U49862 (N_49862,N_49273,N_49376);
or U49863 (N_49863,N_49461,N_49126);
xor U49864 (N_49864,N_49346,N_49023);
nand U49865 (N_49865,N_49442,N_49043);
and U49866 (N_49866,N_49391,N_49306);
xnor U49867 (N_49867,N_49243,N_49394);
nor U49868 (N_49868,N_49074,N_49333);
and U49869 (N_49869,N_49314,N_49467);
nor U49870 (N_49870,N_49209,N_49382);
or U49871 (N_49871,N_49438,N_49430);
or U49872 (N_49872,N_49145,N_49368);
nand U49873 (N_49873,N_49356,N_49349);
and U49874 (N_49874,N_49267,N_49260);
xnor U49875 (N_49875,N_49347,N_49336);
or U49876 (N_49876,N_49402,N_49430);
nor U49877 (N_49877,N_49106,N_49280);
nor U49878 (N_49878,N_49372,N_49038);
nand U49879 (N_49879,N_49256,N_49159);
nor U49880 (N_49880,N_49056,N_49223);
or U49881 (N_49881,N_49133,N_49417);
or U49882 (N_49882,N_49435,N_49031);
nand U49883 (N_49883,N_49191,N_49325);
xor U49884 (N_49884,N_49371,N_49354);
and U49885 (N_49885,N_49018,N_49102);
nand U49886 (N_49886,N_49267,N_49268);
nor U49887 (N_49887,N_49414,N_49426);
nor U49888 (N_49888,N_49336,N_49391);
xnor U49889 (N_49889,N_49328,N_49104);
or U49890 (N_49890,N_49421,N_49036);
nor U49891 (N_49891,N_49248,N_49322);
nor U49892 (N_49892,N_49404,N_49424);
nor U49893 (N_49893,N_49028,N_49192);
or U49894 (N_49894,N_49462,N_49354);
nand U49895 (N_49895,N_49461,N_49047);
and U49896 (N_49896,N_49439,N_49452);
nor U49897 (N_49897,N_49188,N_49390);
nor U49898 (N_49898,N_49431,N_49044);
nor U49899 (N_49899,N_49238,N_49003);
and U49900 (N_49900,N_49491,N_49137);
nand U49901 (N_49901,N_49133,N_49367);
nand U49902 (N_49902,N_49397,N_49078);
xnor U49903 (N_49903,N_49331,N_49421);
or U49904 (N_49904,N_49002,N_49498);
and U49905 (N_49905,N_49139,N_49356);
nand U49906 (N_49906,N_49013,N_49415);
and U49907 (N_49907,N_49138,N_49235);
or U49908 (N_49908,N_49236,N_49193);
nor U49909 (N_49909,N_49205,N_49458);
nor U49910 (N_49910,N_49159,N_49477);
nand U49911 (N_49911,N_49481,N_49477);
and U49912 (N_49912,N_49233,N_49141);
nor U49913 (N_49913,N_49384,N_49255);
and U49914 (N_49914,N_49054,N_49324);
xnor U49915 (N_49915,N_49094,N_49243);
nand U49916 (N_49916,N_49182,N_49344);
and U49917 (N_49917,N_49356,N_49400);
nor U49918 (N_49918,N_49086,N_49088);
or U49919 (N_49919,N_49478,N_49380);
nor U49920 (N_49920,N_49188,N_49009);
nor U49921 (N_49921,N_49474,N_49430);
and U49922 (N_49922,N_49022,N_49207);
and U49923 (N_49923,N_49366,N_49479);
or U49924 (N_49924,N_49107,N_49116);
nand U49925 (N_49925,N_49341,N_49362);
and U49926 (N_49926,N_49413,N_49341);
and U49927 (N_49927,N_49145,N_49004);
nor U49928 (N_49928,N_49489,N_49041);
nor U49929 (N_49929,N_49016,N_49315);
and U49930 (N_49930,N_49165,N_49369);
nor U49931 (N_49931,N_49439,N_49104);
or U49932 (N_49932,N_49386,N_49138);
nor U49933 (N_49933,N_49458,N_49252);
or U49934 (N_49934,N_49000,N_49022);
nand U49935 (N_49935,N_49325,N_49214);
nor U49936 (N_49936,N_49055,N_49476);
nand U49937 (N_49937,N_49370,N_49285);
nand U49938 (N_49938,N_49304,N_49115);
and U49939 (N_49939,N_49228,N_49335);
or U49940 (N_49940,N_49273,N_49497);
nor U49941 (N_49941,N_49004,N_49414);
and U49942 (N_49942,N_49470,N_49483);
nor U49943 (N_49943,N_49378,N_49184);
nor U49944 (N_49944,N_49073,N_49127);
nand U49945 (N_49945,N_49470,N_49457);
nand U49946 (N_49946,N_49279,N_49031);
and U49947 (N_49947,N_49226,N_49411);
nor U49948 (N_49948,N_49060,N_49241);
or U49949 (N_49949,N_49144,N_49076);
nor U49950 (N_49950,N_49341,N_49130);
nand U49951 (N_49951,N_49248,N_49454);
and U49952 (N_49952,N_49044,N_49158);
and U49953 (N_49953,N_49352,N_49295);
xor U49954 (N_49954,N_49316,N_49081);
nor U49955 (N_49955,N_49188,N_49257);
nand U49956 (N_49956,N_49315,N_49129);
nor U49957 (N_49957,N_49382,N_49296);
and U49958 (N_49958,N_49446,N_49474);
nor U49959 (N_49959,N_49126,N_49009);
nand U49960 (N_49960,N_49419,N_49222);
xor U49961 (N_49961,N_49312,N_49398);
or U49962 (N_49962,N_49315,N_49234);
nor U49963 (N_49963,N_49005,N_49289);
nor U49964 (N_49964,N_49333,N_49005);
nand U49965 (N_49965,N_49400,N_49096);
nor U49966 (N_49966,N_49197,N_49309);
nor U49967 (N_49967,N_49116,N_49090);
nand U49968 (N_49968,N_49497,N_49401);
or U49969 (N_49969,N_49238,N_49267);
xor U49970 (N_49970,N_49142,N_49401);
nor U49971 (N_49971,N_49027,N_49325);
xnor U49972 (N_49972,N_49403,N_49429);
and U49973 (N_49973,N_49033,N_49484);
nand U49974 (N_49974,N_49472,N_49216);
nand U49975 (N_49975,N_49422,N_49225);
xnor U49976 (N_49976,N_49433,N_49011);
or U49977 (N_49977,N_49328,N_49123);
nor U49978 (N_49978,N_49114,N_49135);
xor U49979 (N_49979,N_49188,N_49347);
or U49980 (N_49980,N_49355,N_49091);
nand U49981 (N_49981,N_49080,N_49417);
xnor U49982 (N_49982,N_49101,N_49239);
or U49983 (N_49983,N_49217,N_49248);
nor U49984 (N_49984,N_49105,N_49344);
and U49985 (N_49985,N_49034,N_49383);
nand U49986 (N_49986,N_49030,N_49095);
xnor U49987 (N_49987,N_49412,N_49084);
nor U49988 (N_49988,N_49048,N_49362);
nand U49989 (N_49989,N_49409,N_49305);
or U49990 (N_49990,N_49405,N_49361);
and U49991 (N_49991,N_49172,N_49255);
xor U49992 (N_49992,N_49406,N_49422);
nor U49993 (N_49993,N_49177,N_49425);
nand U49994 (N_49994,N_49187,N_49428);
nor U49995 (N_49995,N_49465,N_49476);
nor U49996 (N_49996,N_49403,N_49478);
xor U49997 (N_49997,N_49038,N_49157);
nor U49998 (N_49998,N_49174,N_49416);
nor U49999 (N_49999,N_49448,N_49269);
nor UO_0 (O_0,N_49975,N_49591);
or UO_1 (O_1,N_49822,N_49914);
and UO_2 (O_2,N_49817,N_49505);
nand UO_3 (O_3,N_49983,N_49789);
or UO_4 (O_4,N_49830,N_49570);
and UO_5 (O_5,N_49917,N_49744);
nor UO_6 (O_6,N_49857,N_49986);
or UO_7 (O_7,N_49939,N_49646);
xnor UO_8 (O_8,N_49850,N_49783);
and UO_9 (O_9,N_49928,N_49978);
nand UO_10 (O_10,N_49916,N_49993);
or UO_11 (O_11,N_49927,N_49812);
nand UO_12 (O_12,N_49934,N_49786);
and UO_13 (O_13,N_49540,N_49660);
nand UO_14 (O_14,N_49543,N_49823);
xor UO_15 (O_15,N_49877,N_49717);
xnor UO_16 (O_16,N_49523,N_49611);
and UO_17 (O_17,N_49856,N_49561);
nand UO_18 (O_18,N_49898,N_49662);
or UO_19 (O_19,N_49728,N_49520);
nand UO_20 (O_20,N_49628,N_49528);
nand UO_21 (O_21,N_49743,N_49692);
nand UO_22 (O_22,N_49977,N_49573);
and UO_23 (O_23,N_49669,N_49959);
xor UO_24 (O_24,N_49569,N_49574);
and UO_25 (O_25,N_49947,N_49992);
nand UO_26 (O_26,N_49674,N_49851);
and UO_27 (O_27,N_49776,N_49995);
nand UO_28 (O_28,N_49658,N_49557);
xnor UO_29 (O_29,N_49698,N_49773);
xnor UO_30 (O_30,N_49513,N_49834);
and UO_31 (O_31,N_49852,N_49586);
nand UO_32 (O_32,N_49533,N_49963);
or UO_33 (O_33,N_49577,N_49893);
and UO_34 (O_34,N_49951,N_49645);
nor UO_35 (O_35,N_49584,N_49826);
nor UO_36 (O_36,N_49648,N_49797);
nand UO_37 (O_37,N_49517,N_49595);
and UO_38 (O_38,N_49861,N_49688);
nor UO_39 (O_39,N_49878,N_49883);
and UO_40 (O_40,N_49887,N_49622);
or UO_41 (O_41,N_49976,N_49661);
and UO_42 (O_42,N_49905,N_49945);
or UO_43 (O_43,N_49757,N_49832);
and UO_44 (O_44,N_49871,N_49514);
and UO_45 (O_45,N_49736,N_49695);
xnor UO_46 (O_46,N_49711,N_49726);
nor UO_47 (O_47,N_49705,N_49718);
or UO_48 (O_48,N_49924,N_49954);
nor UO_49 (O_49,N_49549,N_49998);
nand UO_50 (O_50,N_49770,N_49865);
or UO_51 (O_51,N_49870,N_49920);
xor UO_52 (O_52,N_49957,N_49672);
nand UO_53 (O_53,N_49879,N_49709);
xor UO_54 (O_54,N_49537,N_49946);
or UO_55 (O_55,N_49833,N_49530);
and UO_56 (O_56,N_49876,N_49696);
and UO_57 (O_57,N_49619,N_49962);
nor UO_58 (O_58,N_49522,N_49863);
nand UO_59 (O_59,N_49775,N_49875);
and UO_60 (O_60,N_49506,N_49607);
or UO_61 (O_61,N_49604,N_49548);
and UO_62 (O_62,N_49815,N_49710);
nor UO_63 (O_63,N_49862,N_49587);
nor UO_64 (O_64,N_49578,N_49827);
nor UO_65 (O_65,N_49810,N_49748);
or UO_66 (O_66,N_49637,N_49801);
xnor UO_67 (O_67,N_49635,N_49971);
nor UO_68 (O_68,N_49771,N_49930);
nor UO_69 (O_69,N_49665,N_49596);
and UO_70 (O_70,N_49910,N_49614);
xor UO_71 (O_71,N_49932,N_49787);
and UO_72 (O_72,N_49855,N_49583);
nor UO_73 (O_73,N_49994,N_49511);
or UO_74 (O_74,N_49542,N_49938);
nor UO_75 (O_75,N_49866,N_49845);
and UO_76 (O_76,N_49652,N_49747);
nand UO_77 (O_77,N_49690,N_49746);
xor UO_78 (O_78,N_49982,N_49687);
or UO_79 (O_79,N_49781,N_49782);
nand UO_80 (O_80,N_49539,N_49682);
xor UO_81 (O_81,N_49656,N_49667);
xor UO_82 (O_82,N_49700,N_49760);
or UO_83 (O_83,N_49634,N_49551);
xor UO_84 (O_84,N_49545,N_49860);
nor UO_85 (O_85,N_49740,N_49800);
or UO_86 (O_86,N_49684,N_49599);
nand UO_87 (O_87,N_49921,N_49967);
nor UO_88 (O_88,N_49980,N_49825);
xnor UO_89 (O_89,N_49902,N_49550);
or UO_90 (O_90,N_49880,N_49721);
or UO_91 (O_91,N_49942,N_49673);
and UO_92 (O_92,N_49929,N_49714);
or UO_93 (O_93,N_49849,N_49922);
nor UO_94 (O_94,N_49739,N_49538);
nand UO_95 (O_95,N_49791,N_49702);
xnor UO_96 (O_96,N_49680,N_49794);
nor UO_97 (O_97,N_49593,N_49663);
nor UO_98 (O_98,N_49885,N_49670);
or UO_99 (O_99,N_49693,N_49803);
or UO_100 (O_100,N_49544,N_49753);
and UO_101 (O_101,N_49864,N_49654);
nor UO_102 (O_102,N_49608,N_49919);
nor UO_103 (O_103,N_49949,N_49935);
nand UO_104 (O_104,N_49846,N_49940);
xnor UO_105 (O_105,N_49890,N_49598);
and UO_106 (O_106,N_49759,N_49639);
or UO_107 (O_107,N_49899,N_49808);
and UO_108 (O_108,N_49869,N_49751);
and UO_109 (O_109,N_49948,N_49555);
nor UO_110 (O_110,N_49582,N_49854);
nor UO_111 (O_111,N_49676,N_49891);
or UO_112 (O_112,N_49886,N_49572);
or UO_113 (O_113,N_49612,N_49666);
nand UO_114 (O_114,N_49741,N_49524);
xor UO_115 (O_115,N_49955,N_49507);
or UO_116 (O_116,N_49589,N_49972);
nand UO_117 (O_117,N_49950,N_49772);
or UO_118 (O_118,N_49566,N_49501);
or UO_119 (O_119,N_49853,N_49563);
or UO_120 (O_120,N_49636,N_49937);
or UO_121 (O_121,N_49556,N_49754);
nand UO_122 (O_122,N_49761,N_49819);
nor UO_123 (O_123,N_49686,N_49685);
nor UO_124 (O_124,N_49562,N_49923);
and UO_125 (O_125,N_49559,N_49733);
nand UO_126 (O_126,N_49915,N_49839);
nor UO_127 (O_127,N_49807,N_49504);
and UO_128 (O_128,N_49884,N_49848);
and UO_129 (O_129,N_49926,N_49668);
or UO_130 (O_130,N_49704,N_49991);
nor UO_131 (O_131,N_49756,N_49681);
xor UO_132 (O_132,N_49554,N_49953);
and UO_133 (O_133,N_49906,N_49713);
or UO_134 (O_134,N_49627,N_49931);
and UO_135 (O_135,N_49722,N_49502);
and UO_136 (O_136,N_49897,N_49703);
or UO_137 (O_137,N_49647,N_49943);
nor UO_138 (O_138,N_49859,N_49689);
nand UO_139 (O_139,N_49742,N_49996);
nor UO_140 (O_140,N_49867,N_49966);
and UO_141 (O_141,N_49625,N_49701);
nor UO_142 (O_142,N_49987,N_49521);
or UO_143 (O_143,N_49610,N_49626);
and UO_144 (O_144,N_49729,N_49529);
or UO_145 (O_145,N_49762,N_49694);
nor UO_146 (O_146,N_49969,N_49630);
and UO_147 (O_147,N_49970,N_49552);
nor UO_148 (O_148,N_49990,N_49576);
nand UO_149 (O_149,N_49525,N_49677);
nor UO_150 (O_150,N_49838,N_49961);
or UO_151 (O_151,N_49640,N_49588);
xnor UO_152 (O_152,N_49723,N_49602);
and UO_153 (O_153,N_49553,N_49774);
nor UO_154 (O_154,N_49780,N_49769);
xnor UO_155 (O_155,N_49802,N_49795);
and UO_156 (O_156,N_49605,N_49590);
nor UO_157 (O_157,N_49872,N_49793);
xnor UO_158 (O_158,N_49638,N_49974);
or UO_159 (O_159,N_49631,N_49623);
nand UO_160 (O_160,N_49567,N_49650);
nor UO_161 (O_161,N_49565,N_49904);
and UO_162 (O_162,N_49835,N_49911);
or UO_163 (O_163,N_49571,N_49657);
xnor UO_164 (O_164,N_49601,N_49809);
and UO_165 (O_165,N_49732,N_49824);
xnor UO_166 (O_166,N_49738,N_49936);
nand UO_167 (O_167,N_49843,N_49734);
and UO_168 (O_168,N_49725,N_49651);
or UO_169 (O_169,N_49784,N_49644);
xor UO_170 (O_170,N_49913,N_49706);
nor UO_171 (O_171,N_49617,N_49632);
nor UO_172 (O_172,N_49519,N_49818);
xnor UO_173 (O_173,N_49873,N_49821);
and UO_174 (O_174,N_49568,N_49516);
and UO_175 (O_175,N_49988,N_49820);
and UO_176 (O_176,N_49629,N_49708);
and UO_177 (O_177,N_49785,N_49624);
or UO_178 (O_178,N_49960,N_49527);
nand UO_179 (O_179,N_49958,N_49616);
nor UO_180 (O_180,N_49765,N_49500);
nand UO_181 (O_181,N_49618,N_49678);
nand UO_182 (O_182,N_49560,N_49813);
or UO_183 (O_183,N_49964,N_49758);
and UO_184 (O_184,N_49510,N_49811);
nor UO_185 (O_185,N_49615,N_49541);
nand UO_186 (O_186,N_49564,N_49581);
nor UO_187 (O_187,N_49633,N_49896);
xnor UO_188 (O_188,N_49749,N_49512);
nand UO_189 (O_189,N_49597,N_49844);
or UO_190 (O_190,N_49752,N_49755);
xor UO_191 (O_191,N_49727,N_49925);
nor UO_192 (O_192,N_49641,N_49842);
xnor UO_193 (O_193,N_49737,N_49814);
and UO_194 (O_194,N_49659,N_49888);
xor UO_195 (O_195,N_49881,N_49829);
nor UO_196 (O_196,N_49777,N_49613);
nor UO_197 (O_197,N_49903,N_49792);
or UO_198 (O_198,N_49580,N_49944);
xnor UO_199 (O_199,N_49730,N_49778);
nor UO_200 (O_200,N_49894,N_49536);
nand UO_201 (O_201,N_49837,N_49575);
and UO_202 (O_202,N_49768,N_49874);
nand UO_203 (O_203,N_49509,N_49724);
and UO_204 (O_204,N_49779,N_49828);
or UO_205 (O_205,N_49796,N_49900);
or UO_206 (O_206,N_49620,N_49735);
xor UO_207 (O_207,N_49518,N_49788);
nand UO_208 (O_208,N_49831,N_49767);
xor UO_209 (O_209,N_49526,N_49600);
or UO_210 (O_210,N_49892,N_49981);
xnor UO_211 (O_211,N_49683,N_49719);
nor UO_212 (O_212,N_49503,N_49655);
nand UO_213 (O_213,N_49933,N_49508);
or UO_214 (O_214,N_49908,N_49606);
nor UO_215 (O_215,N_49547,N_49965);
nand UO_216 (O_216,N_49889,N_49649);
nor UO_217 (O_217,N_49806,N_49816);
xor UO_218 (O_218,N_49868,N_49973);
nand UO_219 (O_219,N_49558,N_49592);
xnor UO_220 (O_220,N_49609,N_49840);
nand UO_221 (O_221,N_49941,N_49997);
xor UO_222 (O_222,N_49679,N_49621);
and UO_223 (O_223,N_49841,N_49643);
nor UO_224 (O_224,N_49642,N_49901);
nand UO_225 (O_225,N_49790,N_49999);
nor UO_226 (O_226,N_49798,N_49546);
nand UO_227 (O_227,N_49715,N_49952);
nor UO_228 (O_228,N_49763,N_49653);
and UO_229 (O_229,N_49984,N_49675);
nor UO_230 (O_230,N_49799,N_49912);
xnor UO_231 (O_231,N_49671,N_49989);
nand UO_232 (O_232,N_49594,N_49979);
nor UO_233 (O_233,N_49907,N_49716);
nor UO_234 (O_234,N_49532,N_49720);
nor UO_235 (O_235,N_49731,N_49534);
nand UO_236 (O_236,N_49531,N_49858);
nand UO_237 (O_237,N_49579,N_49766);
nor UO_238 (O_238,N_49707,N_49535);
xor UO_239 (O_239,N_49764,N_49712);
nor UO_240 (O_240,N_49847,N_49745);
or UO_241 (O_241,N_49895,N_49882);
nand UO_242 (O_242,N_49585,N_49750);
nand UO_243 (O_243,N_49699,N_49836);
or UO_244 (O_244,N_49804,N_49985);
nor UO_245 (O_245,N_49515,N_49956);
nor UO_246 (O_246,N_49909,N_49805);
xor UO_247 (O_247,N_49691,N_49664);
nor UO_248 (O_248,N_49918,N_49697);
and UO_249 (O_249,N_49968,N_49603);
and UO_250 (O_250,N_49592,N_49510);
xor UO_251 (O_251,N_49530,N_49519);
or UO_252 (O_252,N_49716,N_49919);
nor UO_253 (O_253,N_49654,N_49814);
or UO_254 (O_254,N_49973,N_49705);
nand UO_255 (O_255,N_49579,N_49563);
and UO_256 (O_256,N_49742,N_49812);
nor UO_257 (O_257,N_49570,N_49773);
nand UO_258 (O_258,N_49852,N_49777);
nor UO_259 (O_259,N_49923,N_49540);
and UO_260 (O_260,N_49808,N_49775);
xor UO_261 (O_261,N_49893,N_49761);
nand UO_262 (O_262,N_49738,N_49981);
or UO_263 (O_263,N_49898,N_49857);
xnor UO_264 (O_264,N_49598,N_49702);
nor UO_265 (O_265,N_49779,N_49936);
nand UO_266 (O_266,N_49847,N_49819);
nand UO_267 (O_267,N_49547,N_49759);
or UO_268 (O_268,N_49687,N_49775);
and UO_269 (O_269,N_49636,N_49556);
nand UO_270 (O_270,N_49639,N_49884);
nand UO_271 (O_271,N_49565,N_49803);
xor UO_272 (O_272,N_49732,N_49613);
or UO_273 (O_273,N_49845,N_49611);
and UO_274 (O_274,N_49925,N_49943);
and UO_275 (O_275,N_49880,N_49960);
or UO_276 (O_276,N_49602,N_49840);
nor UO_277 (O_277,N_49937,N_49677);
and UO_278 (O_278,N_49960,N_49794);
xor UO_279 (O_279,N_49577,N_49891);
nor UO_280 (O_280,N_49616,N_49695);
or UO_281 (O_281,N_49798,N_49882);
and UO_282 (O_282,N_49529,N_49553);
nand UO_283 (O_283,N_49565,N_49520);
nand UO_284 (O_284,N_49987,N_49718);
and UO_285 (O_285,N_49744,N_49764);
xor UO_286 (O_286,N_49745,N_49700);
xor UO_287 (O_287,N_49823,N_49552);
and UO_288 (O_288,N_49721,N_49795);
and UO_289 (O_289,N_49758,N_49947);
nand UO_290 (O_290,N_49746,N_49798);
nor UO_291 (O_291,N_49879,N_49966);
or UO_292 (O_292,N_49949,N_49979);
nor UO_293 (O_293,N_49992,N_49900);
or UO_294 (O_294,N_49511,N_49559);
nand UO_295 (O_295,N_49805,N_49912);
and UO_296 (O_296,N_49739,N_49506);
xor UO_297 (O_297,N_49910,N_49779);
and UO_298 (O_298,N_49722,N_49950);
nand UO_299 (O_299,N_49805,N_49713);
nor UO_300 (O_300,N_49730,N_49787);
nor UO_301 (O_301,N_49847,N_49727);
nand UO_302 (O_302,N_49982,N_49712);
nand UO_303 (O_303,N_49648,N_49574);
nand UO_304 (O_304,N_49656,N_49891);
or UO_305 (O_305,N_49901,N_49817);
nor UO_306 (O_306,N_49748,N_49535);
nand UO_307 (O_307,N_49766,N_49591);
nor UO_308 (O_308,N_49768,N_49717);
or UO_309 (O_309,N_49705,N_49896);
and UO_310 (O_310,N_49560,N_49924);
and UO_311 (O_311,N_49783,N_49683);
nand UO_312 (O_312,N_49902,N_49812);
xnor UO_313 (O_313,N_49718,N_49619);
or UO_314 (O_314,N_49559,N_49504);
xor UO_315 (O_315,N_49815,N_49888);
xor UO_316 (O_316,N_49968,N_49895);
xnor UO_317 (O_317,N_49762,N_49505);
nand UO_318 (O_318,N_49770,N_49741);
nor UO_319 (O_319,N_49725,N_49845);
or UO_320 (O_320,N_49873,N_49825);
nand UO_321 (O_321,N_49939,N_49508);
and UO_322 (O_322,N_49993,N_49657);
nor UO_323 (O_323,N_49928,N_49777);
nand UO_324 (O_324,N_49753,N_49674);
xor UO_325 (O_325,N_49943,N_49926);
and UO_326 (O_326,N_49999,N_49825);
or UO_327 (O_327,N_49612,N_49538);
or UO_328 (O_328,N_49961,N_49558);
nand UO_329 (O_329,N_49876,N_49726);
or UO_330 (O_330,N_49808,N_49693);
nand UO_331 (O_331,N_49800,N_49642);
and UO_332 (O_332,N_49574,N_49897);
xor UO_333 (O_333,N_49709,N_49871);
and UO_334 (O_334,N_49615,N_49931);
and UO_335 (O_335,N_49822,N_49763);
nor UO_336 (O_336,N_49551,N_49712);
nand UO_337 (O_337,N_49999,N_49559);
and UO_338 (O_338,N_49779,N_49746);
xor UO_339 (O_339,N_49752,N_49565);
nand UO_340 (O_340,N_49582,N_49639);
or UO_341 (O_341,N_49664,N_49895);
and UO_342 (O_342,N_49827,N_49705);
nand UO_343 (O_343,N_49821,N_49906);
and UO_344 (O_344,N_49687,N_49851);
or UO_345 (O_345,N_49794,N_49822);
and UO_346 (O_346,N_49988,N_49951);
and UO_347 (O_347,N_49564,N_49828);
xnor UO_348 (O_348,N_49737,N_49771);
and UO_349 (O_349,N_49897,N_49820);
xnor UO_350 (O_350,N_49993,N_49775);
nor UO_351 (O_351,N_49781,N_49507);
and UO_352 (O_352,N_49702,N_49797);
and UO_353 (O_353,N_49762,N_49542);
or UO_354 (O_354,N_49738,N_49835);
nor UO_355 (O_355,N_49950,N_49898);
xnor UO_356 (O_356,N_49574,N_49768);
and UO_357 (O_357,N_49727,N_49872);
xor UO_358 (O_358,N_49774,N_49714);
nand UO_359 (O_359,N_49641,N_49642);
and UO_360 (O_360,N_49623,N_49979);
and UO_361 (O_361,N_49762,N_49743);
xor UO_362 (O_362,N_49887,N_49572);
or UO_363 (O_363,N_49941,N_49903);
nand UO_364 (O_364,N_49640,N_49770);
and UO_365 (O_365,N_49905,N_49951);
nor UO_366 (O_366,N_49775,N_49928);
nor UO_367 (O_367,N_49589,N_49928);
or UO_368 (O_368,N_49699,N_49594);
or UO_369 (O_369,N_49723,N_49931);
and UO_370 (O_370,N_49617,N_49711);
xor UO_371 (O_371,N_49652,N_49673);
or UO_372 (O_372,N_49975,N_49945);
xnor UO_373 (O_373,N_49733,N_49771);
or UO_374 (O_374,N_49983,N_49518);
and UO_375 (O_375,N_49589,N_49973);
and UO_376 (O_376,N_49989,N_49818);
nand UO_377 (O_377,N_49543,N_49579);
or UO_378 (O_378,N_49951,N_49902);
nor UO_379 (O_379,N_49847,N_49569);
and UO_380 (O_380,N_49865,N_49762);
nand UO_381 (O_381,N_49776,N_49913);
and UO_382 (O_382,N_49582,N_49684);
and UO_383 (O_383,N_49748,N_49819);
or UO_384 (O_384,N_49900,N_49762);
xor UO_385 (O_385,N_49584,N_49765);
xnor UO_386 (O_386,N_49753,N_49927);
xor UO_387 (O_387,N_49902,N_49888);
xor UO_388 (O_388,N_49886,N_49953);
xnor UO_389 (O_389,N_49676,N_49651);
nand UO_390 (O_390,N_49515,N_49771);
xor UO_391 (O_391,N_49920,N_49981);
nand UO_392 (O_392,N_49588,N_49728);
nor UO_393 (O_393,N_49689,N_49796);
and UO_394 (O_394,N_49609,N_49524);
and UO_395 (O_395,N_49867,N_49573);
xnor UO_396 (O_396,N_49863,N_49965);
nor UO_397 (O_397,N_49982,N_49502);
nor UO_398 (O_398,N_49696,N_49871);
or UO_399 (O_399,N_49599,N_49737);
or UO_400 (O_400,N_49877,N_49555);
nand UO_401 (O_401,N_49790,N_49824);
nand UO_402 (O_402,N_49709,N_49979);
xnor UO_403 (O_403,N_49754,N_49557);
xnor UO_404 (O_404,N_49841,N_49741);
or UO_405 (O_405,N_49812,N_49974);
and UO_406 (O_406,N_49872,N_49958);
and UO_407 (O_407,N_49641,N_49518);
or UO_408 (O_408,N_49764,N_49823);
nor UO_409 (O_409,N_49544,N_49520);
nand UO_410 (O_410,N_49724,N_49691);
nor UO_411 (O_411,N_49654,N_49659);
or UO_412 (O_412,N_49648,N_49719);
xnor UO_413 (O_413,N_49531,N_49907);
and UO_414 (O_414,N_49820,N_49544);
or UO_415 (O_415,N_49596,N_49780);
or UO_416 (O_416,N_49570,N_49514);
and UO_417 (O_417,N_49878,N_49963);
nor UO_418 (O_418,N_49610,N_49853);
or UO_419 (O_419,N_49855,N_49613);
xnor UO_420 (O_420,N_49510,N_49501);
nand UO_421 (O_421,N_49631,N_49859);
and UO_422 (O_422,N_49831,N_49684);
xnor UO_423 (O_423,N_49665,N_49963);
nand UO_424 (O_424,N_49606,N_49511);
nor UO_425 (O_425,N_49547,N_49691);
or UO_426 (O_426,N_49935,N_49827);
and UO_427 (O_427,N_49982,N_49947);
nor UO_428 (O_428,N_49753,N_49779);
nand UO_429 (O_429,N_49969,N_49571);
and UO_430 (O_430,N_49647,N_49967);
nor UO_431 (O_431,N_49904,N_49569);
nor UO_432 (O_432,N_49872,N_49986);
or UO_433 (O_433,N_49654,N_49771);
nand UO_434 (O_434,N_49742,N_49574);
xnor UO_435 (O_435,N_49544,N_49981);
nor UO_436 (O_436,N_49790,N_49571);
nor UO_437 (O_437,N_49562,N_49708);
xnor UO_438 (O_438,N_49606,N_49987);
nor UO_439 (O_439,N_49832,N_49612);
nand UO_440 (O_440,N_49791,N_49953);
and UO_441 (O_441,N_49765,N_49968);
nand UO_442 (O_442,N_49572,N_49718);
nor UO_443 (O_443,N_49947,N_49659);
or UO_444 (O_444,N_49672,N_49576);
or UO_445 (O_445,N_49756,N_49933);
nor UO_446 (O_446,N_49739,N_49607);
nand UO_447 (O_447,N_49840,N_49985);
xor UO_448 (O_448,N_49560,N_49875);
nor UO_449 (O_449,N_49976,N_49787);
and UO_450 (O_450,N_49878,N_49532);
nor UO_451 (O_451,N_49503,N_49923);
or UO_452 (O_452,N_49533,N_49686);
and UO_453 (O_453,N_49609,N_49941);
nor UO_454 (O_454,N_49573,N_49564);
xnor UO_455 (O_455,N_49576,N_49742);
and UO_456 (O_456,N_49919,N_49515);
nand UO_457 (O_457,N_49535,N_49607);
nor UO_458 (O_458,N_49783,N_49922);
nor UO_459 (O_459,N_49598,N_49905);
nor UO_460 (O_460,N_49701,N_49769);
nor UO_461 (O_461,N_49875,N_49801);
and UO_462 (O_462,N_49635,N_49912);
and UO_463 (O_463,N_49879,N_49524);
and UO_464 (O_464,N_49584,N_49961);
nor UO_465 (O_465,N_49601,N_49976);
nand UO_466 (O_466,N_49934,N_49663);
nand UO_467 (O_467,N_49626,N_49636);
nand UO_468 (O_468,N_49763,N_49940);
nor UO_469 (O_469,N_49984,N_49923);
nand UO_470 (O_470,N_49781,N_49549);
nor UO_471 (O_471,N_49524,N_49695);
nor UO_472 (O_472,N_49960,N_49999);
nor UO_473 (O_473,N_49718,N_49679);
or UO_474 (O_474,N_49531,N_49734);
nand UO_475 (O_475,N_49751,N_49924);
and UO_476 (O_476,N_49657,N_49997);
xnor UO_477 (O_477,N_49654,N_49696);
nor UO_478 (O_478,N_49785,N_49518);
and UO_479 (O_479,N_49666,N_49892);
nor UO_480 (O_480,N_49728,N_49879);
and UO_481 (O_481,N_49934,N_49710);
and UO_482 (O_482,N_49648,N_49807);
xor UO_483 (O_483,N_49752,N_49503);
or UO_484 (O_484,N_49564,N_49819);
and UO_485 (O_485,N_49613,N_49949);
and UO_486 (O_486,N_49802,N_49798);
and UO_487 (O_487,N_49696,N_49593);
and UO_488 (O_488,N_49846,N_49736);
xnor UO_489 (O_489,N_49773,N_49811);
or UO_490 (O_490,N_49787,N_49719);
or UO_491 (O_491,N_49507,N_49812);
nand UO_492 (O_492,N_49850,N_49908);
nand UO_493 (O_493,N_49891,N_49636);
and UO_494 (O_494,N_49756,N_49682);
xnor UO_495 (O_495,N_49797,N_49745);
xnor UO_496 (O_496,N_49793,N_49855);
xnor UO_497 (O_497,N_49623,N_49792);
and UO_498 (O_498,N_49859,N_49699);
xnor UO_499 (O_499,N_49958,N_49517);
nor UO_500 (O_500,N_49852,N_49727);
and UO_501 (O_501,N_49743,N_49776);
nand UO_502 (O_502,N_49815,N_49684);
and UO_503 (O_503,N_49869,N_49661);
nand UO_504 (O_504,N_49658,N_49706);
or UO_505 (O_505,N_49622,N_49546);
nor UO_506 (O_506,N_49884,N_49648);
and UO_507 (O_507,N_49825,N_49524);
nor UO_508 (O_508,N_49854,N_49866);
or UO_509 (O_509,N_49645,N_49607);
and UO_510 (O_510,N_49789,N_49730);
xnor UO_511 (O_511,N_49774,N_49528);
nand UO_512 (O_512,N_49702,N_49759);
and UO_513 (O_513,N_49754,N_49546);
nand UO_514 (O_514,N_49852,N_49561);
nor UO_515 (O_515,N_49534,N_49901);
nand UO_516 (O_516,N_49842,N_49937);
nand UO_517 (O_517,N_49811,N_49861);
or UO_518 (O_518,N_49627,N_49706);
nand UO_519 (O_519,N_49501,N_49551);
nand UO_520 (O_520,N_49975,N_49925);
and UO_521 (O_521,N_49693,N_49759);
or UO_522 (O_522,N_49520,N_49514);
or UO_523 (O_523,N_49929,N_49986);
xor UO_524 (O_524,N_49861,N_49611);
nor UO_525 (O_525,N_49771,N_49836);
nand UO_526 (O_526,N_49770,N_49912);
xnor UO_527 (O_527,N_49976,N_49687);
or UO_528 (O_528,N_49832,N_49587);
xor UO_529 (O_529,N_49551,N_49598);
nand UO_530 (O_530,N_49678,N_49627);
nor UO_531 (O_531,N_49598,N_49974);
nor UO_532 (O_532,N_49703,N_49901);
nand UO_533 (O_533,N_49556,N_49557);
or UO_534 (O_534,N_49654,N_49705);
xor UO_535 (O_535,N_49580,N_49711);
nand UO_536 (O_536,N_49536,N_49971);
xor UO_537 (O_537,N_49967,N_49794);
nand UO_538 (O_538,N_49592,N_49847);
or UO_539 (O_539,N_49546,N_49603);
nor UO_540 (O_540,N_49946,N_49924);
and UO_541 (O_541,N_49880,N_49722);
nand UO_542 (O_542,N_49895,N_49928);
nand UO_543 (O_543,N_49707,N_49995);
xnor UO_544 (O_544,N_49671,N_49814);
nand UO_545 (O_545,N_49871,N_49929);
nand UO_546 (O_546,N_49626,N_49876);
nor UO_547 (O_547,N_49541,N_49614);
or UO_548 (O_548,N_49772,N_49790);
nor UO_549 (O_549,N_49550,N_49690);
nor UO_550 (O_550,N_49506,N_49759);
xor UO_551 (O_551,N_49855,N_49977);
xor UO_552 (O_552,N_49604,N_49609);
and UO_553 (O_553,N_49939,N_49858);
nand UO_554 (O_554,N_49770,N_49857);
or UO_555 (O_555,N_49606,N_49521);
or UO_556 (O_556,N_49567,N_49969);
xor UO_557 (O_557,N_49813,N_49653);
and UO_558 (O_558,N_49703,N_49669);
nand UO_559 (O_559,N_49746,N_49544);
nor UO_560 (O_560,N_49992,N_49588);
or UO_561 (O_561,N_49844,N_49888);
and UO_562 (O_562,N_49821,N_49667);
nand UO_563 (O_563,N_49568,N_49929);
and UO_564 (O_564,N_49703,N_49967);
and UO_565 (O_565,N_49831,N_49591);
nand UO_566 (O_566,N_49673,N_49771);
xnor UO_567 (O_567,N_49824,N_49695);
and UO_568 (O_568,N_49737,N_49703);
nand UO_569 (O_569,N_49501,N_49547);
nand UO_570 (O_570,N_49681,N_49665);
or UO_571 (O_571,N_49642,N_49566);
and UO_572 (O_572,N_49888,N_49954);
xor UO_573 (O_573,N_49918,N_49865);
nor UO_574 (O_574,N_49717,N_49719);
and UO_575 (O_575,N_49534,N_49950);
xnor UO_576 (O_576,N_49562,N_49774);
xor UO_577 (O_577,N_49887,N_49509);
nor UO_578 (O_578,N_49969,N_49723);
or UO_579 (O_579,N_49527,N_49590);
nor UO_580 (O_580,N_49794,N_49658);
and UO_581 (O_581,N_49538,N_49736);
and UO_582 (O_582,N_49735,N_49924);
nand UO_583 (O_583,N_49699,N_49981);
nand UO_584 (O_584,N_49726,N_49698);
or UO_585 (O_585,N_49643,N_49649);
xor UO_586 (O_586,N_49909,N_49509);
or UO_587 (O_587,N_49601,N_49987);
and UO_588 (O_588,N_49532,N_49773);
xor UO_589 (O_589,N_49996,N_49660);
nor UO_590 (O_590,N_49991,N_49515);
xnor UO_591 (O_591,N_49504,N_49583);
nor UO_592 (O_592,N_49987,N_49921);
and UO_593 (O_593,N_49626,N_49593);
nand UO_594 (O_594,N_49639,N_49564);
xor UO_595 (O_595,N_49796,N_49673);
nor UO_596 (O_596,N_49598,N_49637);
nor UO_597 (O_597,N_49595,N_49774);
xor UO_598 (O_598,N_49688,N_49920);
nor UO_599 (O_599,N_49770,N_49727);
or UO_600 (O_600,N_49630,N_49761);
nor UO_601 (O_601,N_49992,N_49762);
or UO_602 (O_602,N_49659,N_49691);
nand UO_603 (O_603,N_49582,N_49520);
and UO_604 (O_604,N_49854,N_49938);
nor UO_605 (O_605,N_49698,N_49858);
and UO_606 (O_606,N_49628,N_49930);
and UO_607 (O_607,N_49931,N_49559);
xor UO_608 (O_608,N_49621,N_49531);
nor UO_609 (O_609,N_49723,N_49915);
and UO_610 (O_610,N_49924,N_49531);
and UO_611 (O_611,N_49919,N_49743);
xnor UO_612 (O_612,N_49850,N_49874);
and UO_613 (O_613,N_49814,N_49891);
nor UO_614 (O_614,N_49815,N_49539);
and UO_615 (O_615,N_49519,N_49892);
nor UO_616 (O_616,N_49590,N_49687);
and UO_617 (O_617,N_49959,N_49526);
xor UO_618 (O_618,N_49627,N_49694);
and UO_619 (O_619,N_49980,N_49550);
nand UO_620 (O_620,N_49801,N_49771);
nor UO_621 (O_621,N_49804,N_49795);
nor UO_622 (O_622,N_49745,N_49972);
nand UO_623 (O_623,N_49890,N_49690);
xor UO_624 (O_624,N_49674,N_49783);
nand UO_625 (O_625,N_49858,N_49516);
xor UO_626 (O_626,N_49736,N_49928);
and UO_627 (O_627,N_49521,N_49608);
or UO_628 (O_628,N_49587,N_49603);
nor UO_629 (O_629,N_49509,N_49707);
xnor UO_630 (O_630,N_49516,N_49725);
and UO_631 (O_631,N_49665,N_49504);
or UO_632 (O_632,N_49976,N_49673);
nand UO_633 (O_633,N_49712,N_49923);
and UO_634 (O_634,N_49758,N_49989);
xor UO_635 (O_635,N_49635,N_49957);
xor UO_636 (O_636,N_49568,N_49519);
xnor UO_637 (O_637,N_49908,N_49924);
or UO_638 (O_638,N_49591,N_49869);
xor UO_639 (O_639,N_49629,N_49917);
xor UO_640 (O_640,N_49704,N_49547);
and UO_641 (O_641,N_49877,N_49553);
or UO_642 (O_642,N_49583,N_49867);
or UO_643 (O_643,N_49647,N_49766);
nand UO_644 (O_644,N_49776,N_49542);
xnor UO_645 (O_645,N_49539,N_49841);
and UO_646 (O_646,N_49677,N_49522);
and UO_647 (O_647,N_49628,N_49656);
nor UO_648 (O_648,N_49876,N_49563);
nand UO_649 (O_649,N_49840,N_49686);
and UO_650 (O_650,N_49543,N_49512);
nand UO_651 (O_651,N_49959,N_49924);
and UO_652 (O_652,N_49901,N_49785);
and UO_653 (O_653,N_49741,N_49613);
nor UO_654 (O_654,N_49607,N_49748);
xor UO_655 (O_655,N_49990,N_49828);
nor UO_656 (O_656,N_49671,N_49652);
or UO_657 (O_657,N_49573,N_49591);
nor UO_658 (O_658,N_49550,N_49571);
and UO_659 (O_659,N_49808,N_49592);
xor UO_660 (O_660,N_49626,N_49695);
or UO_661 (O_661,N_49846,N_49893);
xor UO_662 (O_662,N_49949,N_49989);
nor UO_663 (O_663,N_49830,N_49693);
or UO_664 (O_664,N_49908,N_49660);
nor UO_665 (O_665,N_49776,N_49937);
nor UO_666 (O_666,N_49599,N_49751);
nand UO_667 (O_667,N_49743,N_49535);
nand UO_668 (O_668,N_49625,N_49809);
and UO_669 (O_669,N_49552,N_49822);
xnor UO_670 (O_670,N_49556,N_49937);
and UO_671 (O_671,N_49802,N_49720);
or UO_672 (O_672,N_49786,N_49859);
xor UO_673 (O_673,N_49525,N_49980);
xnor UO_674 (O_674,N_49638,N_49644);
nor UO_675 (O_675,N_49634,N_49825);
and UO_676 (O_676,N_49524,N_49536);
xor UO_677 (O_677,N_49500,N_49632);
or UO_678 (O_678,N_49507,N_49601);
nor UO_679 (O_679,N_49758,N_49615);
nor UO_680 (O_680,N_49848,N_49724);
xor UO_681 (O_681,N_49747,N_49842);
or UO_682 (O_682,N_49629,N_49847);
nand UO_683 (O_683,N_49529,N_49850);
nor UO_684 (O_684,N_49974,N_49678);
nor UO_685 (O_685,N_49515,N_49714);
nand UO_686 (O_686,N_49623,N_49660);
and UO_687 (O_687,N_49754,N_49867);
nand UO_688 (O_688,N_49905,N_49953);
xor UO_689 (O_689,N_49616,N_49841);
nand UO_690 (O_690,N_49651,N_49652);
nand UO_691 (O_691,N_49802,N_49977);
nand UO_692 (O_692,N_49863,N_49738);
or UO_693 (O_693,N_49755,N_49996);
and UO_694 (O_694,N_49681,N_49590);
nor UO_695 (O_695,N_49675,N_49946);
or UO_696 (O_696,N_49516,N_49845);
nand UO_697 (O_697,N_49906,N_49847);
and UO_698 (O_698,N_49863,N_49699);
xor UO_699 (O_699,N_49651,N_49800);
and UO_700 (O_700,N_49617,N_49894);
nor UO_701 (O_701,N_49959,N_49731);
xnor UO_702 (O_702,N_49938,N_49915);
xor UO_703 (O_703,N_49695,N_49669);
xnor UO_704 (O_704,N_49927,N_49886);
or UO_705 (O_705,N_49682,N_49827);
xor UO_706 (O_706,N_49924,N_49535);
and UO_707 (O_707,N_49808,N_49666);
xnor UO_708 (O_708,N_49637,N_49953);
and UO_709 (O_709,N_49605,N_49849);
and UO_710 (O_710,N_49867,N_49981);
or UO_711 (O_711,N_49503,N_49972);
nor UO_712 (O_712,N_49530,N_49655);
and UO_713 (O_713,N_49637,N_49866);
or UO_714 (O_714,N_49950,N_49789);
or UO_715 (O_715,N_49836,N_49573);
nor UO_716 (O_716,N_49877,N_49803);
or UO_717 (O_717,N_49978,N_49753);
or UO_718 (O_718,N_49750,N_49575);
nor UO_719 (O_719,N_49779,N_49522);
xnor UO_720 (O_720,N_49987,N_49663);
nor UO_721 (O_721,N_49683,N_49715);
or UO_722 (O_722,N_49692,N_49572);
or UO_723 (O_723,N_49948,N_49644);
nand UO_724 (O_724,N_49784,N_49995);
or UO_725 (O_725,N_49804,N_49569);
or UO_726 (O_726,N_49577,N_49896);
nand UO_727 (O_727,N_49880,N_49693);
nand UO_728 (O_728,N_49739,N_49546);
xnor UO_729 (O_729,N_49893,N_49781);
and UO_730 (O_730,N_49788,N_49651);
nand UO_731 (O_731,N_49952,N_49613);
nor UO_732 (O_732,N_49700,N_49784);
xnor UO_733 (O_733,N_49839,N_49921);
nor UO_734 (O_734,N_49741,N_49855);
xor UO_735 (O_735,N_49904,N_49908);
xnor UO_736 (O_736,N_49556,N_49647);
and UO_737 (O_737,N_49830,N_49804);
and UO_738 (O_738,N_49505,N_49831);
nor UO_739 (O_739,N_49824,N_49686);
and UO_740 (O_740,N_49941,N_49782);
and UO_741 (O_741,N_49576,N_49838);
nand UO_742 (O_742,N_49800,N_49581);
nand UO_743 (O_743,N_49731,N_49945);
nand UO_744 (O_744,N_49631,N_49896);
nand UO_745 (O_745,N_49987,N_49561);
and UO_746 (O_746,N_49745,N_49941);
or UO_747 (O_747,N_49779,N_49512);
xor UO_748 (O_748,N_49728,N_49731);
nand UO_749 (O_749,N_49561,N_49602);
or UO_750 (O_750,N_49549,N_49825);
xnor UO_751 (O_751,N_49831,N_49578);
nor UO_752 (O_752,N_49762,N_49705);
nand UO_753 (O_753,N_49811,N_49930);
nand UO_754 (O_754,N_49927,N_49863);
nor UO_755 (O_755,N_49604,N_49933);
and UO_756 (O_756,N_49522,N_49902);
and UO_757 (O_757,N_49678,N_49761);
nor UO_758 (O_758,N_49525,N_49575);
nor UO_759 (O_759,N_49899,N_49728);
or UO_760 (O_760,N_49904,N_49850);
and UO_761 (O_761,N_49926,N_49844);
xor UO_762 (O_762,N_49742,N_49615);
nand UO_763 (O_763,N_49941,N_49804);
nand UO_764 (O_764,N_49793,N_49890);
nand UO_765 (O_765,N_49613,N_49672);
nor UO_766 (O_766,N_49552,N_49598);
nand UO_767 (O_767,N_49964,N_49546);
or UO_768 (O_768,N_49984,N_49660);
nor UO_769 (O_769,N_49932,N_49513);
and UO_770 (O_770,N_49597,N_49619);
or UO_771 (O_771,N_49526,N_49621);
nand UO_772 (O_772,N_49976,N_49995);
nor UO_773 (O_773,N_49905,N_49502);
or UO_774 (O_774,N_49895,N_49756);
nand UO_775 (O_775,N_49934,N_49841);
nor UO_776 (O_776,N_49820,N_49528);
nand UO_777 (O_777,N_49521,N_49565);
and UO_778 (O_778,N_49905,N_49931);
nand UO_779 (O_779,N_49639,N_49665);
nand UO_780 (O_780,N_49721,N_49981);
and UO_781 (O_781,N_49521,N_49906);
and UO_782 (O_782,N_49569,N_49837);
and UO_783 (O_783,N_49862,N_49776);
nand UO_784 (O_784,N_49938,N_49602);
or UO_785 (O_785,N_49514,N_49511);
nand UO_786 (O_786,N_49919,N_49871);
nor UO_787 (O_787,N_49682,N_49764);
nand UO_788 (O_788,N_49860,N_49929);
nand UO_789 (O_789,N_49890,N_49957);
nand UO_790 (O_790,N_49994,N_49737);
xnor UO_791 (O_791,N_49631,N_49988);
and UO_792 (O_792,N_49917,N_49802);
xnor UO_793 (O_793,N_49622,N_49989);
nand UO_794 (O_794,N_49847,N_49859);
nor UO_795 (O_795,N_49697,N_49555);
nand UO_796 (O_796,N_49984,N_49911);
nor UO_797 (O_797,N_49907,N_49814);
nand UO_798 (O_798,N_49695,N_49632);
nor UO_799 (O_799,N_49979,N_49927);
nand UO_800 (O_800,N_49988,N_49558);
nor UO_801 (O_801,N_49508,N_49555);
and UO_802 (O_802,N_49522,N_49783);
and UO_803 (O_803,N_49634,N_49901);
nor UO_804 (O_804,N_49814,N_49559);
xor UO_805 (O_805,N_49515,N_49980);
or UO_806 (O_806,N_49625,N_49977);
xor UO_807 (O_807,N_49915,N_49569);
and UO_808 (O_808,N_49578,N_49811);
or UO_809 (O_809,N_49662,N_49518);
nor UO_810 (O_810,N_49888,N_49727);
nand UO_811 (O_811,N_49719,N_49732);
and UO_812 (O_812,N_49895,N_49531);
or UO_813 (O_813,N_49758,N_49757);
or UO_814 (O_814,N_49549,N_49907);
xor UO_815 (O_815,N_49515,N_49989);
nand UO_816 (O_816,N_49764,N_49769);
nor UO_817 (O_817,N_49719,N_49593);
nor UO_818 (O_818,N_49575,N_49943);
xnor UO_819 (O_819,N_49893,N_49537);
nand UO_820 (O_820,N_49639,N_49958);
and UO_821 (O_821,N_49799,N_49560);
or UO_822 (O_822,N_49724,N_49557);
nor UO_823 (O_823,N_49836,N_49748);
nand UO_824 (O_824,N_49580,N_49913);
and UO_825 (O_825,N_49755,N_49761);
and UO_826 (O_826,N_49886,N_49908);
and UO_827 (O_827,N_49708,N_49829);
and UO_828 (O_828,N_49691,N_49816);
and UO_829 (O_829,N_49640,N_49566);
xor UO_830 (O_830,N_49872,N_49980);
xor UO_831 (O_831,N_49857,N_49518);
and UO_832 (O_832,N_49705,N_49871);
xnor UO_833 (O_833,N_49810,N_49888);
and UO_834 (O_834,N_49804,N_49933);
xor UO_835 (O_835,N_49626,N_49608);
xor UO_836 (O_836,N_49931,N_49997);
and UO_837 (O_837,N_49955,N_49654);
and UO_838 (O_838,N_49558,N_49791);
nand UO_839 (O_839,N_49764,N_49527);
nand UO_840 (O_840,N_49980,N_49762);
nand UO_841 (O_841,N_49824,N_49643);
and UO_842 (O_842,N_49837,N_49941);
and UO_843 (O_843,N_49572,N_49688);
nor UO_844 (O_844,N_49858,N_49500);
xnor UO_845 (O_845,N_49531,N_49911);
or UO_846 (O_846,N_49950,N_49512);
nor UO_847 (O_847,N_49609,N_49697);
nor UO_848 (O_848,N_49777,N_49507);
nand UO_849 (O_849,N_49960,N_49553);
nor UO_850 (O_850,N_49814,N_49552);
nand UO_851 (O_851,N_49805,N_49850);
nor UO_852 (O_852,N_49614,N_49886);
and UO_853 (O_853,N_49943,N_49572);
and UO_854 (O_854,N_49929,N_49792);
nor UO_855 (O_855,N_49562,N_49535);
nand UO_856 (O_856,N_49502,N_49561);
and UO_857 (O_857,N_49905,N_49691);
nor UO_858 (O_858,N_49872,N_49808);
xor UO_859 (O_859,N_49972,N_49907);
xnor UO_860 (O_860,N_49860,N_49715);
nor UO_861 (O_861,N_49564,N_49700);
nor UO_862 (O_862,N_49542,N_49818);
xnor UO_863 (O_863,N_49707,N_49533);
and UO_864 (O_864,N_49791,N_49993);
xnor UO_865 (O_865,N_49534,N_49566);
and UO_866 (O_866,N_49893,N_49804);
and UO_867 (O_867,N_49845,N_49984);
nor UO_868 (O_868,N_49723,N_49870);
and UO_869 (O_869,N_49975,N_49835);
or UO_870 (O_870,N_49627,N_49548);
nor UO_871 (O_871,N_49921,N_49676);
and UO_872 (O_872,N_49943,N_49611);
nand UO_873 (O_873,N_49762,N_49758);
nand UO_874 (O_874,N_49659,N_49583);
or UO_875 (O_875,N_49777,N_49720);
and UO_876 (O_876,N_49985,N_49989);
xor UO_877 (O_877,N_49575,N_49910);
xor UO_878 (O_878,N_49990,N_49668);
nor UO_879 (O_879,N_49869,N_49938);
xor UO_880 (O_880,N_49703,N_49826);
nor UO_881 (O_881,N_49775,N_49700);
nor UO_882 (O_882,N_49501,N_49638);
xor UO_883 (O_883,N_49794,N_49829);
or UO_884 (O_884,N_49519,N_49701);
xnor UO_885 (O_885,N_49730,N_49753);
xor UO_886 (O_886,N_49540,N_49972);
nor UO_887 (O_887,N_49688,N_49817);
nor UO_888 (O_888,N_49705,N_49932);
or UO_889 (O_889,N_49668,N_49601);
xnor UO_890 (O_890,N_49571,N_49798);
or UO_891 (O_891,N_49548,N_49590);
nor UO_892 (O_892,N_49635,N_49972);
nor UO_893 (O_893,N_49868,N_49977);
nor UO_894 (O_894,N_49987,N_49630);
xor UO_895 (O_895,N_49637,N_49975);
xor UO_896 (O_896,N_49821,N_49560);
nand UO_897 (O_897,N_49843,N_49585);
and UO_898 (O_898,N_49798,N_49799);
nor UO_899 (O_899,N_49664,N_49610);
nor UO_900 (O_900,N_49889,N_49987);
and UO_901 (O_901,N_49841,N_49963);
and UO_902 (O_902,N_49515,N_49542);
xor UO_903 (O_903,N_49546,N_49618);
nor UO_904 (O_904,N_49611,N_49828);
nor UO_905 (O_905,N_49592,N_49730);
or UO_906 (O_906,N_49646,N_49749);
or UO_907 (O_907,N_49515,N_49888);
nand UO_908 (O_908,N_49596,N_49786);
xor UO_909 (O_909,N_49501,N_49997);
xor UO_910 (O_910,N_49857,N_49985);
or UO_911 (O_911,N_49783,N_49939);
and UO_912 (O_912,N_49749,N_49795);
xnor UO_913 (O_913,N_49687,N_49841);
nand UO_914 (O_914,N_49579,N_49933);
nand UO_915 (O_915,N_49552,N_49926);
and UO_916 (O_916,N_49930,N_49777);
and UO_917 (O_917,N_49928,N_49588);
or UO_918 (O_918,N_49602,N_49539);
or UO_919 (O_919,N_49764,N_49807);
nand UO_920 (O_920,N_49968,N_49798);
or UO_921 (O_921,N_49825,N_49991);
nand UO_922 (O_922,N_49640,N_49561);
xor UO_923 (O_923,N_49808,N_49593);
nand UO_924 (O_924,N_49766,N_49605);
or UO_925 (O_925,N_49645,N_49685);
nand UO_926 (O_926,N_49527,N_49537);
nor UO_927 (O_927,N_49549,N_49727);
nand UO_928 (O_928,N_49885,N_49951);
nand UO_929 (O_929,N_49839,N_49581);
nand UO_930 (O_930,N_49755,N_49572);
nor UO_931 (O_931,N_49825,N_49835);
and UO_932 (O_932,N_49505,N_49747);
nand UO_933 (O_933,N_49510,N_49675);
and UO_934 (O_934,N_49656,N_49646);
nand UO_935 (O_935,N_49674,N_49624);
or UO_936 (O_936,N_49632,N_49736);
and UO_937 (O_937,N_49752,N_49703);
xnor UO_938 (O_938,N_49686,N_49889);
nand UO_939 (O_939,N_49716,N_49705);
nor UO_940 (O_940,N_49720,N_49892);
xor UO_941 (O_941,N_49726,N_49626);
and UO_942 (O_942,N_49909,N_49903);
xnor UO_943 (O_943,N_49973,N_49928);
or UO_944 (O_944,N_49731,N_49874);
and UO_945 (O_945,N_49983,N_49555);
or UO_946 (O_946,N_49969,N_49684);
nand UO_947 (O_947,N_49550,N_49637);
nor UO_948 (O_948,N_49682,N_49725);
nand UO_949 (O_949,N_49849,N_49566);
nand UO_950 (O_950,N_49929,N_49737);
and UO_951 (O_951,N_49518,N_49549);
nor UO_952 (O_952,N_49916,N_49626);
nand UO_953 (O_953,N_49964,N_49821);
xnor UO_954 (O_954,N_49924,N_49765);
xnor UO_955 (O_955,N_49579,N_49557);
or UO_956 (O_956,N_49784,N_49685);
and UO_957 (O_957,N_49571,N_49523);
nand UO_958 (O_958,N_49623,N_49522);
nor UO_959 (O_959,N_49508,N_49530);
or UO_960 (O_960,N_49725,N_49686);
nand UO_961 (O_961,N_49627,N_49527);
or UO_962 (O_962,N_49514,N_49812);
xor UO_963 (O_963,N_49669,N_49964);
nand UO_964 (O_964,N_49839,N_49803);
xor UO_965 (O_965,N_49634,N_49800);
xor UO_966 (O_966,N_49564,N_49882);
or UO_967 (O_967,N_49501,N_49962);
and UO_968 (O_968,N_49955,N_49653);
nor UO_969 (O_969,N_49730,N_49679);
xor UO_970 (O_970,N_49872,N_49881);
xnor UO_971 (O_971,N_49760,N_49802);
xor UO_972 (O_972,N_49847,N_49522);
xnor UO_973 (O_973,N_49994,N_49572);
and UO_974 (O_974,N_49813,N_49946);
xor UO_975 (O_975,N_49946,N_49752);
nor UO_976 (O_976,N_49818,N_49657);
and UO_977 (O_977,N_49529,N_49983);
nand UO_978 (O_978,N_49949,N_49761);
and UO_979 (O_979,N_49648,N_49747);
and UO_980 (O_980,N_49871,N_49500);
and UO_981 (O_981,N_49723,N_49734);
or UO_982 (O_982,N_49943,N_49930);
nand UO_983 (O_983,N_49751,N_49951);
or UO_984 (O_984,N_49900,N_49509);
and UO_985 (O_985,N_49898,N_49886);
nand UO_986 (O_986,N_49809,N_49965);
and UO_987 (O_987,N_49634,N_49954);
nand UO_988 (O_988,N_49607,N_49599);
nor UO_989 (O_989,N_49696,N_49793);
and UO_990 (O_990,N_49761,N_49692);
and UO_991 (O_991,N_49732,N_49919);
and UO_992 (O_992,N_49551,N_49655);
nand UO_993 (O_993,N_49882,N_49736);
nand UO_994 (O_994,N_49799,N_49518);
nor UO_995 (O_995,N_49918,N_49610);
nor UO_996 (O_996,N_49943,N_49905);
nand UO_997 (O_997,N_49875,N_49578);
nand UO_998 (O_998,N_49745,N_49964);
nand UO_999 (O_999,N_49602,N_49967);
or UO_1000 (O_1000,N_49898,N_49839);
nor UO_1001 (O_1001,N_49531,N_49620);
xnor UO_1002 (O_1002,N_49672,N_49906);
and UO_1003 (O_1003,N_49760,N_49735);
or UO_1004 (O_1004,N_49725,N_49611);
xor UO_1005 (O_1005,N_49717,N_49545);
and UO_1006 (O_1006,N_49815,N_49696);
xor UO_1007 (O_1007,N_49970,N_49686);
nand UO_1008 (O_1008,N_49524,N_49806);
nor UO_1009 (O_1009,N_49618,N_49579);
xor UO_1010 (O_1010,N_49523,N_49775);
xor UO_1011 (O_1011,N_49737,N_49898);
xnor UO_1012 (O_1012,N_49937,N_49786);
or UO_1013 (O_1013,N_49918,N_49768);
or UO_1014 (O_1014,N_49634,N_49739);
nand UO_1015 (O_1015,N_49982,N_49552);
xor UO_1016 (O_1016,N_49512,N_49544);
and UO_1017 (O_1017,N_49552,N_49914);
and UO_1018 (O_1018,N_49695,N_49845);
or UO_1019 (O_1019,N_49940,N_49535);
nor UO_1020 (O_1020,N_49741,N_49862);
nor UO_1021 (O_1021,N_49950,N_49612);
nor UO_1022 (O_1022,N_49724,N_49564);
xor UO_1023 (O_1023,N_49557,N_49954);
or UO_1024 (O_1024,N_49779,N_49960);
and UO_1025 (O_1025,N_49999,N_49769);
or UO_1026 (O_1026,N_49748,N_49572);
nand UO_1027 (O_1027,N_49685,N_49898);
and UO_1028 (O_1028,N_49508,N_49565);
and UO_1029 (O_1029,N_49735,N_49856);
and UO_1030 (O_1030,N_49552,N_49752);
and UO_1031 (O_1031,N_49852,N_49842);
nand UO_1032 (O_1032,N_49829,N_49874);
and UO_1033 (O_1033,N_49922,N_49525);
or UO_1034 (O_1034,N_49978,N_49897);
xnor UO_1035 (O_1035,N_49892,N_49880);
xor UO_1036 (O_1036,N_49627,N_49782);
nand UO_1037 (O_1037,N_49958,N_49904);
nor UO_1038 (O_1038,N_49880,N_49630);
or UO_1039 (O_1039,N_49527,N_49884);
nor UO_1040 (O_1040,N_49607,N_49711);
nand UO_1041 (O_1041,N_49991,N_49651);
xor UO_1042 (O_1042,N_49663,N_49816);
nor UO_1043 (O_1043,N_49766,N_49800);
and UO_1044 (O_1044,N_49710,N_49634);
nor UO_1045 (O_1045,N_49940,N_49994);
or UO_1046 (O_1046,N_49605,N_49678);
xnor UO_1047 (O_1047,N_49718,N_49749);
xnor UO_1048 (O_1048,N_49563,N_49884);
or UO_1049 (O_1049,N_49731,N_49914);
xnor UO_1050 (O_1050,N_49898,N_49771);
nand UO_1051 (O_1051,N_49617,N_49835);
xor UO_1052 (O_1052,N_49953,N_49719);
and UO_1053 (O_1053,N_49633,N_49682);
nor UO_1054 (O_1054,N_49704,N_49923);
and UO_1055 (O_1055,N_49809,N_49890);
nand UO_1056 (O_1056,N_49982,N_49672);
xor UO_1057 (O_1057,N_49985,N_49758);
and UO_1058 (O_1058,N_49706,N_49539);
or UO_1059 (O_1059,N_49613,N_49726);
or UO_1060 (O_1060,N_49682,N_49875);
xnor UO_1061 (O_1061,N_49814,N_49521);
xnor UO_1062 (O_1062,N_49956,N_49516);
nor UO_1063 (O_1063,N_49536,N_49933);
nor UO_1064 (O_1064,N_49610,N_49784);
nor UO_1065 (O_1065,N_49725,N_49715);
and UO_1066 (O_1066,N_49516,N_49927);
nand UO_1067 (O_1067,N_49915,N_49802);
nand UO_1068 (O_1068,N_49682,N_49848);
and UO_1069 (O_1069,N_49897,N_49843);
or UO_1070 (O_1070,N_49663,N_49758);
and UO_1071 (O_1071,N_49935,N_49693);
and UO_1072 (O_1072,N_49995,N_49629);
or UO_1073 (O_1073,N_49514,N_49853);
nor UO_1074 (O_1074,N_49934,N_49859);
or UO_1075 (O_1075,N_49769,N_49791);
and UO_1076 (O_1076,N_49584,N_49998);
or UO_1077 (O_1077,N_49643,N_49830);
and UO_1078 (O_1078,N_49694,N_49649);
and UO_1079 (O_1079,N_49944,N_49852);
nor UO_1080 (O_1080,N_49992,N_49862);
or UO_1081 (O_1081,N_49834,N_49878);
or UO_1082 (O_1082,N_49599,N_49826);
or UO_1083 (O_1083,N_49793,N_49533);
nor UO_1084 (O_1084,N_49977,N_49732);
nor UO_1085 (O_1085,N_49933,N_49548);
xor UO_1086 (O_1086,N_49640,N_49517);
or UO_1087 (O_1087,N_49594,N_49928);
and UO_1088 (O_1088,N_49735,N_49885);
nand UO_1089 (O_1089,N_49568,N_49560);
or UO_1090 (O_1090,N_49664,N_49965);
or UO_1091 (O_1091,N_49810,N_49669);
or UO_1092 (O_1092,N_49844,N_49523);
nand UO_1093 (O_1093,N_49583,N_49509);
xnor UO_1094 (O_1094,N_49832,N_49930);
nand UO_1095 (O_1095,N_49670,N_49531);
nor UO_1096 (O_1096,N_49971,N_49989);
nand UO_1097 (O_1097,N_49718,N_49881);
nor UO_1098 (O_1098,N_49710,N_49567);
and UO_1099 (O_1099,N_49571,N_49521);
xnor UO_1100 (O_1100,N_49907,N_49585);
nand UO_1101 (O_1101,N_49646,N_49548);
nor UO_1102 (O_1102,N_49517,N_49738);
xnor UO_1103 (O_1103,N_49951,N_49892);
or UO_1104 (O_1104,N_49983,N_49561);
and UO_1105 (O_1105,N_49877,N_49862);
nor UO_1106 (O_1106,N_49582,N_49630);
or UO_1107 (O_1107,N_49964,N_49862);
and UO_1108 (O_1108,N_49713,N_49773);
and UO_1109 (O_1109,N_49694,N_49819);
or UO_1110 (O_1110,N_49527,N_49500);
or UO_1111 (O_1111,N_49869,N_49942);
xor UO_1112 (O_1112,N_49979,N_49805);
nand UO_1113 (O_1113,N_49699,N_49767);
xnor UO_1114 (O_1114,N_49611,N_49548);
nand UO_1115 (O_1115,N_49670,N_49898);
nor UO_1116 (O_1116,N_49779,N_49956);
nor UO_1117 (O_1117,N_49626,N_49517);
nor UO_1118 (O_1118,N_49705,N_49719);
nand UO_1119 (O_1119,N_49935,N_49626);
or UO_1120 (O_1120,N_49733,N_49598);
xnor UO_1121 (O_1121,N_49670,N_49811);
and UO_1122 (O_1122,N_49876,N_49518);
nor UO_1123 (O_1123,N_49719,N_49629);
nor UO_1124 (O_1124,N_49857,N_49902);
xor UO_1125 (O_1125,N_49604,N_49827);
xor UO_1126 (O_1126,N_49865,N_49678);
and UO_1127 (O_1127,N_49649,N_49515);
nor UO_1128 (O_1128,N_49884,N_49836);
and UO_1129 (O_1129,N_49863,N_49620);
or UO_1130 (O_1130,N_49988,N_49592);
and UO_1131 (O_1131,N_49919,N_49722);
or UO_1132 (O_1132,N_49781,N_49694);
xnor UO_1133 (O_1133,N_49787,N_49816);
nor UO_1134 (O_1134,N_49598,N_49910);
and UO_1135 (O_1135,N_49702,N_49957);
nand UO_1136 (O_1136,N_49648,N_49954);
nand UO_1137 (O_1137,N_49799,N_49517);
nor UO_1138 (O_1138,N_49956,N_49959);
nor UO_1139 (O_1139,N_49890,N_49903);
nand UO_1140 (O_1140,N_49727,N_49741);
or UO_1141 (O_1141,N_49704,N_49705);
xor UO_1142 (O_1142,N_49590,N_49684);
xnor UO_1143 (O_1143,N_49611,N_49579);
xnor UO_1144 (O_1144,N_49916,N_49702);
xor UO_1145 (O_1145,N_49651,N_49710);
xor UO_1146 (O_1146,N_49735,N_49557);
nand UO_1147 (O_1147,N_49770,N_49668);
nand UO_1148 (O_1148,N_49928,N_49702);
and UO_1149 (O_1149,N_49599,N_49953);
or UO_1150 (O_1150,N_49551,N_49776);
xor UO_1151 (O_1151,N_49651,N_49625);
nand UO_1152 (O_1152,N_49684,N_49726);
nand UO_1153 (O_1153,N_49615,N_49558);
or UO_1154 (O_1154,N_49864,N_49824);
or UO_1155 (O_1155,N_49648,N_49789);
xnor UO_1156 (O_1156,N_49672,N_49700);
nor UO_1157 (O_1157,N_49740,N_49710);
xor UO_1158 (O_1158,N_49918,N_49744);
nand UO_1159 (O_1159,N_49507,N_49929);
or UO_1160 (O_1160,N_49812,N_49815);
nor UO_1161 (O_1161,N_49741,N_49645);
and UO_1162 (O_1162,N_49696,N_49814);
and UO_1163 (O_1163,N_49775,N_49799);
nor UO_1164 (O_1164,N_49856,N_49973);
nor UO_1165 (O_1165,N_49918,N_49881);
nand UO_1166 (O_1166,N_49663,N_49847);
nor UO_1167 (O_1167,N_49891,N_49668);
nor UO_1168 (O_1168,N_49740,N_49876);
nor UO_1169 (O_1169,N_49545,N_49744);
nand UO_1170 (O_1170,N_49504,N_49721);
xor UO_1171 (O_1171,N_49882,N_49755);
nor UO_1172 (O_1172,N_49926,N_49846);
nor UO_1173 (O_1173,N_49641,N_49830);
nor UO_1174 (O_1174,N_49869,N_49705);
nand UO_1175 (O_1175,N_49798,N_49942);
or UO_1176 (O_1176,N_49689,N_49783);
nor UO_1177 (O_1177,N_49645,N_49691);
xnor UO_1178 (O_1178,N_49529,N_49818);
xor UO_1179 (O_1179,N_49827,N_49597);
nor UO_1180 (O_1180,N_49623,N_49947);
and UO_1181 (O_1181,N_49657,N_49752);
nor UO_1182 (O_1182,N_49674,N_49780);
or UO_1183 (O_1183,N_49993,N_49511);
or UO_1184 (O_1184,N_49671,N_49796);
or UO_1185 (O_1185,N_49654,N_49636);
and UO_1186 (O_1186,N_49518,N_49563);
or UO_1187 (O_1187,N_49636,N_49692);
nor UO_1188 (O_1188,N_49990,N_49883);
nor UO_1189 (O_1189,N_49954,N_49998);
xnor UO_1190 (O_1190,N_49971,N_49624);
nor UO_1191 (O_1191,N_49806,N_49662);
xor UO_1192 (O_1192,N_49507,N_49633);
xnor UO_1193 (O_1193,N_49830,N_49669);
xor UO_1194 (O_1194,N_49849,N_49887);
or UO_1195 (O_1195,N_49588,N_49626);
xor UO_1196 (O_1196,N_49637,N_49962);
or UO_1197 (O_1197,N_49539,N_49554);
or UO_1198 (O_1198,N_49584,N_49967);
xnor UO_1199 (O_1199,N_49645,N_49759);
nor UO_1200 (O_1200,N_49515,N_49792);
nor UO_1201 (O_1201,N_49513,N_49533);
nand UO_1202 (O_1202,N_49786,N_49727);
xor UO_1203 (O_1203,N_49804,N_49687);
nand UO_1204 (O_1204,N_49721,N_49691);
nand UO_1205 (O_1205,N_49596,N_49607);
xor UO_1206 (O_1206,N_49681,N_49758);
or UO_1207 (O_1207,N_49847,N_49740);
nand UO_1208 (O_1208,N_49513,N_49678);
nor UO_1209 (O_1209,N_49505,N_49944);
nand UO_1210 (O_1210,N_49595,N_49953);
nor UO_1211 (O_1211,N_49674,N_49558);
or UO_1212 (O_1212,N_49630,N_49742);
nor UO_1213 (O_1213,N_49538,N_49804);
nand UO_1214 (O_1214,N_49860,N_49908);
nor UO_1215 (O_1215,N_49690,N_49784);
xnor UO_1216 (O_1216,N_49973,N_49948);
nand UO_1217 (O_1217,N_49958,N_49532);
and UO_1218 (O_1218,N_49845,N_49674);
nand UO_1219 (O_1219,N_49660,N_49544);
nor UO_1220 (O_1220,N_49754,N_49998);
nand UO_1221 (O_1221,N_49996,N_49609);
or UO_1222 (O_1222,N_49771,N_49766);
nand UO_1223 (O_1223,N_49700,N_49813);
or UO_1224 (O_1224,N_49909,N_49627);
or UO_1225 (O_1225,N_49852,N_49611);
nor UO_1226 (O_1226,N_49720,N_49693);
or UO_1227 (O_1227,N_49800,N_49861);
nor UO_1228 (O_1228,N_49755,N_49505);
and UO_1229 (O_1229,N_49725,N_49930);
nand UO_1230 (O_1230,N_49932,N_49836);
xnor UO_1231 (O_1231,N_49752,N_49785);
and UO_1232 (O_1232,N_49716,N_49658);
nand UO_1233 (O_1233,N_49730,N_49526);
nor UO_1234 (O_1234,N_49837,N_49808);
and UO_1235 (O_1235,N_49533,N_49622);
nand UO_1236 (O_1236,N_49566,N_49844);
nor UO_1237 (O_1237,N_49910,N_49940);
xor UO_1238 (O_1238,N_49678,N_49623);
and UO_1239 (O_1239,N_49655,N_49544);
nor UO_1240 (O_1240,N_49951,N_49684);
nand UO_1241 (O_1241,N_49888,N_49933);
nand UO_1242 (O_1242,N_49618,N_49768);
and UO_1243 (O_1243,N_49889,N_49605);
and UO_1244 (O_1244,N_49561,N_49617);
and UO_1245 (O_1245,N_49609,N_49858);
or UO_1246 (O_1246,N_49597,N_49826);
nand UO_1247 (O_1247,N_49702,N_49961);
nand UO_1248 (O_1248,N_49662,N_49918);
or UO_1249 (O_1249,N_49729,N_49631);
xor UO_1250 (O_1250,N_49864,N_49779);
nor UO_1251 (O_1251,N_49995,N_49944);
xnor UO_1252 (O_1252,N_49765,N_49694);
or UO_1253 (O_1253,N_49677,N_49794);
or UO_1254 (O_1254,N_49610,N_49689);
nand UO_1255 (O_1255,N_49647,N_49744);
xor UO_1256 (O_1256,N_49827,N_49691);
nor UO_1257 (O_1257,N_49912,N_49777);
or UO_1258 (O_1258,N_49648,N_49772);
xor UO_1259 (O_1259,N_49950,N_49655);
and UO_1260 (O_1260,N_49833,N_49520);
and UO_1261 (O_1261,N_49914,N_49630);
nor UO_1262 (O_1262,N_49833,N_49928);
and UO_1263 (O_1263,N_49605,N_49770);
nor UO_1264 (O_1264,N_49775,N_49521);
and UO_1265 (O_1265,N_49596,N_49816);
xor UO_1266 (O_1266,N_49840,N_49614);
and UO_1267 (O_1267,N_49734,N_49933);
or UO_1268 (O_1268,N_49701,N_49675);
or UO_1269 (O_1269,N_49572,N_49704);
nor UO_1270 (O_1270,N_49688,N_49767);
or UO_1271 (O_1271,N_49549,N_49798);
xor UO_1272 (O_1272,N_49821,N_49991);
xnor UO_1273 (O_1273,N_49863,N_49884);
nor UO_1274 (O_1274,N_49615,N_49863);
nand UO_1275 (O_1275,N_49664,N_49515);
or UO_1276 (O_1276,N_49886,N_49583);
nand UO_1277 (O_1277,N_49818,N_49848);
nor UO_1278 (O_1278,N_49559,N_49954);
nand UO_1279 (O_1279,N_49641,N_49875);
xor UO_1280 (O_1280,N_49584,N_49876);
xor UO_1281 (O_1281,N_49781,N_49908);
or UO_1282 (O_1282,N_49927,N_49549);
nor UO_1283 (O_1283,N_49892,N_49911);
nand UO_1284 (O_1284,N_49645,N_49667);
nor UO_1285 (O_1285,N_49887,N_49523);
and UO_1286 (O_1286,N_49586,N_49677);
nor UO_1287 (O_1287,N_49502,N_49524);
xnor UO_1288 (O_1288,N_49927,N_49700);
xor UO_1289 (O_1289,N_49871,N_49958);
nor UO_1290 (O_1290,N_49863,N_49671);
nand UO_1291 (O_1291,N_49850,N_49646);
xnor UO_1292 (O_1292,N_49675,N_49790);
nor UO_1293 (O_1293,N_49662,N_49965);
nor UO_1294 (O_1294,N_49846,N_49780);
nand UO_1295 (O_1295,N_49650,N_49778);
or UO_1296 (O_1296,N_49799,N_49715);
and UO_1297 (O_1297,N_49675,N_49967);
or UO_1298 (O_1298,N_49861,N_49508);
nand UO_1299 (O_1299,N_49563,N_49633);
nor UO_1300 (O_1300,N_49670,N_49960);
xnor UO_1301 (O_1301,N_49573,N_49618);
nand UO_1302 (O_1302,N_49783,N_49510);
nand UO_1303 (O_1303,N_49715,N_49682);
xnor UO_1304 (O_1304,N_49914,N_49739);
and UO_1305 (O_1305,N_49672,N_49950);
or UO_1306 (O_1306,N_49753,N_49642);
nand UO_1307 (O_1307,N_49802,N_49853);
nand UO_1308 (O_1308,N_49941,N_49799);
nand UO_1309 (O_1309,N_49507,N_49717);
or UO_1310 (O_1310,N_49524,N_49597);
nand UO_1311 (O_1311,N_49662,N_49509);
nor UO_1312 (O_1312,N_49551,N_49775);
xor UO_1313 (O_1313,N_49802,N_49625);
and UO_1314 (O_1314,N_49660,N_49883);
nor UO_1315 (O_1315,N_49788,N_49729);
and UO_1316 (O_1316,N_49936,N_49974);
or UO_1317 (O_1317,N_49603,N_49504);
nor UO_1318 (O_1318,N_49795,N_49912);
or UO_1319 (O_1319,N_49866,N_49877);
and UO_1320 (O_1320,N_49626,N_49507);
xnor UO_1321 (O_1321,N_49946,N_49777);
and UO_1322 (O_1322,N_49733,N_49787);
nand UO_1323 (O_1323,N_49719,N_49678);
or UO_1324 (O_1324,N_49810,N_49692);
or UO_1325 (O_1325,N_49749,N_49881);
and UO_1326 (O_1326,N_49950,N_49531);
nor UO_1327 (O_1327,N_49960,N_49936);
and UO_1328 (O_1328,N_49844,N_49755);
or UO_1329 (O_1329,N_49622,N_49712);
xnor UO_1330 (O_1330,N_49693,N_49749);
and UO_1331 (O_1331,N_49751,N_49985);
nor UO_1332 (O_1332,N_49860,N_49985);
and UO_1333 (O_1333,N_49904,N_49878);
or UO_1334 (O_1334,N_49649,N_49966);
or UO_1335 (O_1335,N_49885,N_49603);
nor UO_1336 (O_1336,N_49613,N_49896);
or UO_1337 (O_1337,N_49664,N_49743);
xor UO_1338 (O_1338,N_49893,N_49614);
nand UO_1339 (O_1339,N_49621,N_49982);
xor UO_1340 (O_1340,N_49808,N_49606);
and UO_1341 (O_1341,N_49594,N_49763);
nand UO_1342 (O_1342,N_49993,N_49781);
or UO_1343 (O_1343,N_49883,N_49649);
or UO_1344 (O_1344,N_49714,N_49775);
nor UO_1345 (O_1345,N_49798,N_49981);
nand UO_1346 (O_1346,N_49511,N_49898);
nand UO_1347 (O_1347,N_49719,N_49980);
nand UO_1348 (O_1348,N_49779,N_49715);
or UO_1349 (O_1349,N_49705,N_49693);
or UO_1350 (O_1350,N_49924,N_49565);
or UO_1351 (O_1351,N_49957,N_49638);
nor UO_1352 (O_1352,N_49893,N_49699);
xnor UO_1353 (O_1353,N_49520,N_49942);
nand UO_1354 (O_1354,N_49786,N_49967);
and UO_1355 (O_1355,N_49945,N_49503);
xnor UO_1356 (O_1356,N_49729,N_49528);
xor UO_1357 (O_1357,N_49977,N_49638);
nor UO_1358 (O_1358,N_49925,N_49553);
nand UO_1359 (O_1359,N_49941,N_49621);
xor UO_1360 (O_1360,N_49740,N_49918);
nand UO_1361 (O_1361,N_49512,N_49566);
nand UO_1362 (O_1362,N_49510,N_49994);
nand UO_1363 (O_1363,N_49825,N_49876);
nor UO_1364 (O_1364,N_49630,N_49530);
xor UO_1365 (O_1365,N_49894,N_49726);
xnor UO_1366 (O_1366,N_49662,N_49540);
xor UO_1367 (O_1367,N_49612,N_49688);
xnor UO_1368 (O_1368,N_49624,N_49610);
and UO_1369 (O_1369,N_49709,N_49812);
nand UO_1370 (O_1370,N_49709,N_49783);
and UO_1371 (O_1371,N_49522,N_49910);
nand UO_1372 (O_1372,N_49525,N_49591);
nand UO_1373 (O_1373,N_49900,N_49951);
nand UO_1374 (O_1374,N_49563,N_49990);
xnor UO_1375 (O_1375,N_49554,N_49797);
and UO_1376 (O_1376,N_49910,N_49948);
nand UO_1377 (O_1377,N_49838,N_49932);
or UO_1378 (O_1378,N_49961,N_49572);
nand UO_1379 (O_1379,N_49994,N_49705);
xnor UO_1380 (O_1380,N_49638,N_49853);
nor UO_1381 (O_1381,N_49807,N_49612);
xor UO_1382 (O_1382,N_49977,N_49644);
xnor UO_1383 (O_1383,N_49902,N_49540);
nand UO_1384 (O_1384,N_49595,N_49917);
nand UO_1385 (O_1385,N_49879,N_49951);
and UO_1386 (O_1386,N_49674,N_49800);
and UO_1387 (O_1387,N_49594,N_49819);
nor UO_1388 (O_1388,N_49750,N_49507);
nand UO_1389 (O_1389,N_49928,N_49730);
nor UO_1390 (O_1390,N_49923,N_49702);
nor UO_1391 (O_1391,N_49724,N_49605);
or UO_1392 (O_1392,N_49821,N_49792);
or UO_1393 (O_1393,N_49739,N_49521);
nand UO_1394 (O_1394,N_49541,N_49657);
nor UO_1395 (O_1395,N_49902,N_49945);
nor UO_1396 (O_1396,N_49647,N_49825);
or UO_1397 (O_1397,N_49835,N_49581);
nor UO_1398 (O_1398,N_49512,N_49977);
nand UO_1399 (O_1399,N_49969,N_49627);
or UO_1400 (O_1400,N_49510,N_49762);
nand UO_1401 (O_1401,N_49642,N_49747);
nor UO_1402 (O_1402,N_49709,N_49989);
nor UO_1403 (O_1403,N_49634,N_49748);
and UO_1404 (O_1404,N_49885,N_49625);
and UO_1405 (O_1405,N_49504,N_49601);
xor UO_1406 (O_1406,N_49556,N_49689);
nor UO_1407 (O_1407,N_49675,N_49963);
nand UO_1408 (O_1408,N_49849,N_49715);
and UO_1409 (O_1409,N_49521,N_49947);
or UO_1410 (O_1410,N_49591,N_49548);
nand UO_1411 (O_1411,N_49610,N_49660);
or UO_1412 (O_1412,N_49698,N_49853);
and UO_1413 (O_1413,N_49982,N_49936);
xnor UO_1414 (O_1414,N_49865,N_49928);
nor UO_1415 (O_1415,N_49598,N_49979);
nand UO_1416 (O_1416,N_49569,N_49957);
and UO_1417 (O_1417,N_49559,N_49831);
xnor UO_1418 (O_1418,N_49585,N_49838);
nand UO_1419 (O_1419,N_49974,N_49806);
xnor UO_1420 (O_1420,N_49683,N_49877);
or UO_1421 (O_1421,N_49745,N_49692);
nor UO_1422 (O_1422,N_49619,N_49860);
nand UO_1423 (O_1423,N_49856,N_49550);
or UO_1424 (O_1424,N_49742,N_49684);
and UO_1425 (O_1425,N_49938,N_49982);
xnor UO_1426 (O_1426,N_49770,N_49644);
and UO_1427 (O_1427,N_49901,N_49720);
or UO_1428 (O_1428,N_49562,N_49669);
xnor UO_1429 (O_1429,N_49511,N_49682);
nand UO_1430 (O_1430,N_49571,N_49772);
xor UO_1431 (O_1431,N_49586,N_49721);
and UO_1432 (O_1432,N_49742,N_49745);
xor UO_1433 (O_1433,N_49944,N_49733);
nand UO_1434 (O_1434,N_49760,N_49961);
or UO_1435 (O_1435,N_49594,N_49851);
nor UO_1436 (O_1436,N_49914,N_49518);
xnor UO_1437 (O_1437,N_49728,N_49781);
nand UO_1438 (O_1438,N_49705,N_49659);
nor UO_1439 (O_1439,N_49961,N_49926);
and UO_1440 (O_1440,N_49697,N_49936);
nand UO_1441 (O_1441,N_49876,N_49552);
or UO_1442 (O_1442,N_49742,N_49899);
nor UO_1443 (O_1443,N_49754,N_49523);
xnor UO_1444 (O_1444,N_49532,N_49607);
xor UO_1445 (O_1445,N_49969,N_49965);
or UO_1446 (O_1446,N_49609,N_49975);
xnor UO_1447 (O_1447,N_49966,N_49631);
nand UO_1448 (O_1448,N_49669,N_49686);
or UO_1449 (O_1449,N_49741,N_49502);
and UO_1450 (O_1450,N_49542,N_49618);
and UO_1451 (O_1451,N_49896,N_49554);
nand UO_1452 (O_1452,N_49910,N_49521);
xor UO_1453 (O_1453,N_49630,N_49731);
nor UO_1454 (O_1454,N_49943,N_49953);
xor UO_1455 (O_1455,N_49887,N_49748);
nor UO_1456 (O_1456,N_49595,N_49667);
nor UO_1457 (O_1457,N_49709,N_49680);
and UO_1458 (O_1458,N_49608,N_49927);
or UO_1459 (O_1459,N_49667,N_49751);
or UO_1460 (O_1460,N_49861,N_49844);
and UO_1461 (O_1461,N_49830,N_49703);
nor UO_1462 (O_1462,N_49725,N_49770);
nand UO_1463 (O_1463,N_49932,N_49590);
nand UO_1464 (O_1464,N_49854,N_49565);
or UO_1465 (O_1465,N_49795,N_49731);
or UO_1466 (O_1466,N_49833,N_49717);
or UO_1467 (O_1467,N_49785,N_49533);
nor UO_1468 (O_1468,N_49981,N_49856);
nand UO_1469 (O_1469,N_49907,N_49761);
nor UO_1470 (O_1470,N_49827,N_49852);
xnor UO_1471 (O_1471,N_49822,N_49965);
nand UO_1472 (O_1472,N_49516,N_49815);
xor UO_1473 (O_1473,N_49728,N_49857);
or UO_1474 (O_1474,N_49953,N_49613);
nor UO_1475 (O_1475,N_49540,N_49532);
xnor UO_1476 (O_1476,N_49838,N_49977);
nand UO_1477 (O_1477,N_49810,N_49512);
and UO_1478 (O_1478,N_49897,N_49887);
nor UO_1479 (O_1479,N_49642,N_49996);
or UO_1480 (O_1480,N_49909,N_49818);
and UO_1481 (O_1481,N_49640,N_49761);
xor UO_1482 (O_1482,N_49742,N_49564);
xor UO_1483 (O_1483,N_49532,N_49620);
nand UO_1484 (O_1484,N_49690,N_49854);
nand UO_1485 (O_1485,N_49603,N_49552);
and UO_1486 (O_1486,N_49922,N_49684);
nor UO_1487 (O_1487,N_49837,N_49746);
nor UO_1488 (O_1488,N_49718,N_49816);
nand UO_1489 (O_1489,N_49710,N_49687);
xor UO_1490 (O_1490,N_49778,N_49591);
xor UO_1491 (O_1491,N_49880,N_49889);
nand UO_1492 (O_1492,N_49644,N_49815);
xnor UO_1493 (O_1493,N_49775,N_49585);
nor UO_1494 (O_1494,N_49725,N_49583);
nor UO_1495 (O_1495,N_49527,N_49542);
nor UO_1496 (O_1496,N_49598,N_49864);
or UO_1497 (O_1497,N_49685,N_49934);
and UO_1498 (O_1498,N_49552,N_49874);
nor UO_1499 (O_1499,N_49868,N_49962);
xor UO_1500 (O_1500,N_49699,N_49946);
nor UO_1501 (O_1501,N_49951,N_49772);
and UO_1502 (O_1502,N_49722,N_49741);
or UO_1503 (O_1503,N_49696,N_49621);
nor UO_1504 (O_1504,N_49871,N_49685);
nand UO_1505 (O_1505,N_49892,N_49920);
nor UO_1506 (O_1506,N_49769,N_49759);
nand UO_1507 (O_1507,N_49501,N_49644);
or UO_1508 (O_1508,N_49693,N_49509);
nor UO_1509 (O_1509,N_49793,N_49737);
or UO_1510 (O_1510,N_49794,N_49877);
and UO_1511 (O_1511,N_49897,N_49992);
nor UO_1512 (O_1512,N_49754,N_49771);
nand UO_1513 (O_1513,N_49595,N_49543);
nor UO_1514 (O_1514,N_49584,N_49519);
nor UO_1515 (O_1515,N_49518,N_49630);
xnor UO_1516 (O_1516,N_49806,N_49642);
or UO_1517 (O_1517,N_49649,N_49579);
nor UO_1518 (O_1518,N_49816,N_49700);
nor UO_1519 (O_1519,N_49768,N_49854);
nand UO_1520 (O_1520,N_49915,N_49614);
nand UO_1521 (O_1521,N_49842,N_49585);
xnor UO_1522 (O_1522,N_49870,N_49703);
xor UO_1523 (O_1523,N_49615,N_49790);
and UO_1524 (O_1524,N_49580,N_49753);
nor UO_1525 (O_1525,N_49733,N_49567);
xor UO_1526 (O_1526,N_49758,N_49993);
and UO_1527 (O_1527,N_49978,N_49566);
and UO_1528 (O_1528,N_49776,N_49644);
or UO_1529 (O_1529,N_49586,N_49909);
xor UO_1530 (O_1530,N_49740,N_49691);
nor UO_1531 (O_1531,N_49955,N_49571);
nand UO_1532 (O_1532,N_49781,N_49602);
nand UO_1533 (O_1533,N_49559,N_49695);
nor UO_1534 (O_1534,N_49613,N_49655);
xnor UO_1535 (O_1535,N_49842,N_49773);
nor UO_1536 (O_1536,N_49898,N_49795);
and UO_1537 (O_1537,N_49724,N_49730);
nand UO_1538 (O_1538,N_49731,N_49828);
or UO_1539 (O_1539,N_49786,N_49938);
xnor UO_1540 (O_1540,N_49707,N_49592);
and UO_1541 (O_1541,N_49740,N_49929);
nor UO_1542 (O_1542,N_49514,N_49636);
nor UO_1543 (O_1543,N_49780,N_49986);
or UO_1544 (O_1544,N_49957,N_49703);
xnor UO_1545 (O_1545,N_49632,N_49613);
nor UO_1546 (O_1546,N_49968,N_49914);
and UO_1547 (O_1547,N_49751,N_49944);
and UO_1548 (O_1548,N_49617,N_49859);
or UO_1549 (O_1549,N_49922,N_49979);
xnor UO_1550 (O_1550,N_49645,N_49899);
and UO_1551 (O_1551,N_49782,N_49564);
nor UO_1552 (O_1552,N_49619,N_49829);
nor UO_1553 (O_1553,N_49640,N_49864);
nand UO_1554 (O_1554,N_49857,N_49912);
nand UO_1555 (O_1555,N_49677,N_49661);
xor UO_1556 (O_1556,N_49759,N_49816);
nor UO_1557 (O_1557,N_49786,N_49682);
and UO_1558 (O_1558,N_49865,N_49814);
xor UO_1559 (O_1559,N_49937,N_49721);
or UO_1560 (O_1560,N_49947,N_49531);
xnor UO_1561 (O_1561,N_49757,N_49854);
xor UO_1562 (O_1562,N_49928,N_49828);
nand UO_1563 (O_1563,N_49799,N_49720);
nor UO_1564 (O_1564,N_49642,N_49762);
xor UO_1565 (O_1565,N_49523,N_49876);
nor UO_1566 (O_1566,N_49617,N_49776);
nand UO_1567 (O_1567,N_49747,N_49708);
and UO_1568 (O_1568,N_49575,N_49532);
xnor UO_1569 (O_1569,N_49813,N_49621);
and UO_1570 (O_1570,N_49602,N_49739);
and UO_1571 (O_1571,N_49521,N_49679);
nor UO_1572 (O_1572,N_49726,N_49992);
xor UO_1573 (O_1573,N_49651,N_49972);
xnor UO_1574 (O_1574,N_49588,N_49748);
nor UO_1575 (O_1575,N_49924,N_49875);
and UO_1576 (O_1576,N_49700,N_49805);
nor UO_1577 (O_1577,N_49829,N_49584);
xor UO_1578 (O_1578,N_49938,N_49880);
nand UO_1579 (O_1579,N_49906,N_49792);
nor UO_1580 (O_1580,N_49906,N_49588);
or UO_1581 (O_1581,N_49763,N_49528);
xor UO_1582 (O_1582,N_49807,N_49741);
xnor UO_1583 (O_1583,N_49591,N_49832);
nand UO_1584 (O_1584,N_49788,N_49702);
nor UO_1585 (O_1585,N_49927,N_49746);
xnor UO_1586 (O_1586,N_49979,N_49692);
xnor UO_1587 (O_1587,N_49643,N_49984);
or UO_1588 (O_1588,N_49859,N_49648);
or UO_1589 (O_1589,N_49718,N_49575);
nand UO_1590 (O_1590,N_49832,N_49537);
or UO_1591 (O_1591,N_49790,N_49574);
xor UO_1592 (O_1592,N_49565,N_49869);
or UO_1593 (O_1593,N_49675,N_49582);
or UO_1594 (O_1594,N_49558,N_49651);
xor UO_1595 (O_1595,N_49707,N_49590);
nand UO_1596 (O_1596,N_49624,N_49537);
nand UO_1597 (O_1597,N_49514,N_49893);
nor UO_1598 (O_1598,N_49622,N_49742);
or UO_1599 (O_1599,N_49587,N_49747);
xor UO_1600 (O_1600,N_49872,N_49953);
or UO_1601 (O_1601,N_49930,N_49765);
xnor UO_1602 (O_1602,N_49896,N_49630);
or UO_1603 (O_1603,N_49634,N_49539);
and UO_1604 (O_1604,N_49912,N_49906);
xor UO_1605 (O_1605,N_49895,N_49878);
nor UO_1606 (O_1606,N_49676,N_49769);
nand UO_1607 (O_1607,N_49592,N_49720);
or UO_1608 (O_1608,N_49926,N_49826);
nor UO_1609 (O_1609,N_49502,N_49849);
nand UO_1610 (O_1610,N_49523,N_49675);
and UO_1611 (O_1611,N_49519,N_49835);
or UO_1612 (O_1612,N_49515,N_49558);
and UO_1613 (O_1613,N_49594,N_49902);
nand UO_1614 (O_1614,N_49846,N_49581);
or UO_1615 (O_1615,N_49933,N_49735);
xnor UO_1616 (O_1616,N_49859,N_49564);
xor UO_1617 (O_1617,N_49772,N_49798);
xnor UO_1618 (O_1618,N_49592,N_49637);
or UO_1619 (O_1619,N_49502,N_49658);
nand UO_1620 (O_1620,N_49705,N_49972);
nand UO_1621 (O_1621,N_49578,N_49889);
nor UO_1622 (O_1622,N_49646,N_49500);
or UO_1623 (O_1623,N_49634,N_49511);
or UO_1624 (O_1624,N_49730,N_49525);
xor UO_1625 (O_1625,N_49695,N_49955);
nor UO_1626 (O_1626,N_49653,N_49926);
and UO_1627 (O_1627,N_49566,N_49961);
nand UO_1628 (O_1628,N_49971,N_49849);
and UO_1629 (O_1629,N_49536,N_49960);
xnor UO_1630 (O_1630,N_49757,N_49789);
xnor UO_1631 (O_1631,N_49776,N_49529);
nor UO_1632 (O_1632,N_49844,N_49856);
and UO_1633 (O_1633,N_49668,N_49916);
and UO_1634 (O_1634,N_49782,N_49864);
xor UO_1635 (O_1635,N_49915,N_49752);
or UO_1636 (O_1636,N_49959,N_49725);
nand UO_1637 (O_1637,N_49537,N_49856);
and UO_1638 (O_1638,N_49659,N_49822);
or UO_1639 (O_1639,N_49794,N_49995);
or UO_1640 (O_1640,N_49614,N_49775);
nand UO_1641 (O_1641,N_49551,N_49533);
xnor UO_1642 (O_1642,N_49851,N_49640);
nand UO_1643 (O_1643,N_49576,N_49874);
xnor UO_1644 (O_1644,N_49880,N_49536);
and UO_1645 (O_1645,N_49570,N_49741);
nand UO_1646 (O_1646,N_49709,N_49818);
or UO_1647 (O_1647,N_49549,N_49569);
or UO_1648 (O_1648,N_49585,N_49763);
or UO_1649 (O_1649,N_49968,N_49910);
or UO_1650 (O_1650,N_49985,N_49577);
nor UO_1651 (O_1651,N_49900,N_49512);
xor UO_1652 (O_1652,N_49760,N_49545);
and UO_1653 (O_1653,N_49747,N_49884);
nor UO_1654 (O_1654,N_49767,N_49830);
nand UO_1655 (O_1655,N_49592,N_49957);
and UO_1656 (O_1656,N_49810,N_49974);
nand UO_1657 (O_1657,N_49579,N_49505);
or UO_1658 (O_1658,N_49992,N_49555);
and UO_1659 (O_1659,N_49584,N_49719);
or UO_1660 (O_1660,N_49691,N_49858);
nand UO_1661 (O_1661,N_49684,N_49917);
xnor UO_1662 (O_1662,N_49909,N_49579);
nor UO_1663 (O_1663,N_49815,N_49784);
nor UO_1664 (O_1664,N_49918,N_49760);
or UO_1665 (O_1665,N_49737,N_49838);
nor UO_1666 (O_1666,N_49725,N_49969);
and UO_1667 (O_1667,N_49779,N_49621);
or UO_1668 (O_1668,N_49720,N_49531);
and UO_1669 (O_1669,N_49891,N_49837);
nor UO_1670 (O_1670,N_49598,N_49739);
and UO_1671 (O_1671,N_49753,N_49946);
or UO_1672 (O_1672,N_49694,N_49663);
nor UO_1673 (O_1673,N_49585,N_49981);
or UO_1674 (O_1674,N_49851,N_49765);
nor UO_1675 (O_1675,N_49953,N_49729);
and UO_1676 (O_1676,N_49946,N_49843);
nor UO_1677 (O_1677,N_49685,N_49533);
and UO_1678 (O_1678,N_49737,N_49739);
and UO_1679 (O_1679,N_49765,N_49937);
or UO_1680 (O_1680,N_49852,N_49600);
nor UO_1681 (O_1681,N_49727,N_49940);
or UO_1682 (O_1682,N_49699,N_49627);
nand UO_1683 (O_1683,N_49599,N_49969);
or UO_1684 (O_1684,N_49539,N_49909);
nor UO_1685 (O_1685,N_49651,N_49508);
nor UO_1686 (O_1686,N_49531,N_49638);
or UO_1687 (O_1687,N_49748,N_49579);
nor UO_1688 (O_1688,N_49788,N_49757);
xnor UO_1689 (O_1689,N_49585,N_49768);
nor UO_1690 (O_1690,N_49788,N_49641);
or UO_1691 (O_1691,N_49583,N_49805);
nand UO_1692 (O_1692,N_49880,N_49739);
nand UO_1693 (O_1693,N_49877,N_49552);
or UO_1694 (O_1694,N_49737,N_49587);
nand UO_1695 (O_1695,N_49510,N_49679);
nor UO_1696 (O_1696,N_49573,N_49785);
nor UO_1697 (O_1697,N_49911,N_49753);
or UO_1698 (O_1698,N_49689,N_49853);
and UO_1699 (O_1699,N_49956,N_49609);
and UO_1700 (O_1700,N_49715,N_49537);
and UO_1701 (O_1701,N_49979,N_49754);
or UO_1702 (O_1702,N_49668,N_49772);
and UO_1703 (O_1703,N_49985,N_49760);
xnor UO_1704 (O_1704,N_49650,N_49501);
nand UO_1705 (O_1705,N_49872,N_49654);
nand UO_1706 (O_1706,N_49659,N_49609);
nor UO_1707 (O_1707,N_49627,N_49533);
nand UO_1708 (O_1708,N_49545,N_49984);
nor UO_1709 (O_1709,N_49877,N_49868);
nand UO_1710 (O_1710,N_49715,N_49834);
and UO_1711 (O_1711,N_49501,N_49504);
nor UO_1712 (O_1712,N_49824,N_49986);
and UO_1713 (O_1713,N_49504,N_49700);
nand UO_1714 (O_1714,N_49765,N_49955);
nand UO_1715 (O_1715,N_49716,N_49709);
nand UO_1716 (O_1716,N_49509,N_49833);
nand UO_1717 (O_1717,N_49681,N_49828);
and UO_1718 (O_1718,N_49867,N_49690);
nand UO_1719 (O_1719,N_49563,N_49743);
and UO_1720 (O_1720,N_49957,N_49945);
nor UO_1721 (O_1721,N_49893,N_49532);
xor UO_1722 (O_1722,N_49941,N_49676);
nand UO_1723 (O_1723,N_49750,N_49656);
or UO_1724 (O_1724,N_49857,N_49826);
nand UO_1725 (O_1725,N_49983,N_49636);
nand UO_1726 (O_1726,N_49771,N_49908);
or UO_1727 (O_1727,N_49871,N_49524);
and UO_1728 (O_1728,N_49925,N_49815);
nand UO_1729 (O_1729,N_49990,N_49764);
nand UO_1730 (O_1730,N_49720,N_49639);
nor UO_1731 (O_1731,N_49633,N_49800);
nor UO_1732 (O_1732,N_49724,N_49743);
nor UO_1733 (O_1733,N_49664,N_49648);
nor UO_1734 (O_1734,N_49706,N_49999);
or UO_1735 (O_1735,N_49522,N_49924);
nor UO_1736 (O_1736,N_49561,N_49945);
and UO_1737 (O_1737,N_49700,N_49537);
and UO_1738 (O_1738,N_49699,N_49756);
or UO_1739 (O_1739,N_49781,N_49648);
or UO_1740 (O_1740,N_49524,N_49894);
nor UO_1741 (O_1741,N_49603,N_49571);
nand UO_1742 (O_1742,N_49838,N_49597);
nand UO_1743 (O_1743,N_49612,N_49509);
nor UO_1744 (O_1744,N_49601,N_49903);
xnor UO_1745 (O_1745,N_49970,N_49743);
nor UO_1746 (O_1746,N_49655,N_49818);
nand UO_1747 (O_1747,N_49756,N_49904);
xnor UO_1748 (O_1748,N_49550,N_49759);
nor UO_1749 (O_1749,N_49635,N_49579);
or UO_1750 (O_1750,N_49663,N_49577);
xor UO_1751 (O_1751,N_49638,N_49990);
nor UO_1752 (O_1752,N_49792,N_49628);
or UO_1753 (O_1753,N_49595,N_49976);
or UO_1754 (O_1754,N_49982,N_49691);
and UO_1755 (O_1755,N_49912,N_49555);
xor UO_1756 (O_1756,N_49920,N_49849);
or UO_1757 (O_1757,N_49937,N_49681);
nand UO_1758 (O_1758,N_49930,N_49822);
nor UO_1759 (O_1759,N_49798,N_49811);
nor UO_1760 (O_1760,N_49742,N_49733);
and UO_1761 (O_1761,N_49771,N_49817);
xnor UO_1762 (O_1762,N_49940,N_49896);
and UO_1763 (O_1763,N_49660,N_49918);
nand UO_1764 (O_1764,N_49759,N_49527);
or UO_1765 (O_1765,N_49629,N_49655);
and UO_1766 (O_1766,N_49653,N_49570);
and UO_1767 (O_1767,N_49652,N_49563);
nand UO_1768 (O_1768,N_49526,N_49690);
nor UO_1769 (O_1769,N_49876,N_49786);
xnor UO_1770 (O_1770,N_49744,N_49594);
nand UO_1771 (O_1771,N_49998,N_49540);
and UO_1772 (O_1772,N_49812,N_49638);
nor UO_1773 (O_1773,N_49735,N_49628);
nand UO_1774 (O_1774,N_49636,N_49777);
xor UO_1775 (O_1775,N_49934,N_49845);
and UO_1776 (O_1776,N_49872,N_49743);
nand UO_1777 (O_1777,N_49531,N_49732);
or UO_1778 (O_1778,N_49900,N_49563);
xnor UO_1779 (O_1779,N_49692,N_49691);
xor UO_1780 (O_1780,N_49883,N_49941);
xor UO_1781 (O_1781,N_49675,N_49912);
and UO_1782 (O_1782,N_49859,N_49547);
nand UO_1783 (O_1783,N_49973,N_49527);
xor UO_1784 (O_1784,N_49878,N_49554);
xor UO_1785 (O_1785,N_49985,N_49502);
and UO_1786 (O_1786,N_49592,N_49513);
and UO_1787 (O_1787,N_49668,N_49606);
or UO_1788 (O_1788,N_49577,N_49750);
nand UO_1789 (O_1789,N_49917,N_49717);
xor UO_1790 (O_1790,N_49919,N_49943);
and UO_1791 (O_1791,N_49875,N_49805);
and UO_1792 (O_1792,N_49884,N_49725);
nor UO_1793 (O_1793,N_49941,N_49734);
nand UO_1794 (O_1794,N_49535,N_49776);
xor UO_1795 (O_1795,N_49647,N_49719);
nand UO_1796 (O_1796,N_49666,N_49738);
nor UO_1797 (O_1797,N_49713,N_49634);
or UO_1798 (O_1798,N_49975,N_49857);
xnor UO_1799 (O_1799,N_49862,N_49652);
nand UO_1800 (O_1800,N_49989,N_49981);
nand UO_1801 (O_1801,N_49693,N_49979);
nand UO_1802 (O_1802,N_49569,N_49621);
xnor UO_1803 (O_1803,N_49660,N_49964);
nor UO_1804 (O_1804,N_49621,N_49770);
or UO_1805 (O_1805,N_49514,N_49559);
and UO_1806 (O_1806,N_49869,N_49887);
or UO_1807 (O_1807,N_49651,N_49630);
nor UO_1808 (O_1808,N_49506,N_49949);
and UO_1809 (O_1809,N_49918,N_49555);
and UO_1810 (O_1810,N_49964,N_49942);
xnor UO_1811 (O_1811,N_49881,N_49796);
nor UO_1812 (O_1812,N_49628,N_49906);
or UO_1813 (O_1813,N_49525,N_49886);
nor UO_1814 (O_1814,N_49876,N_49660);
nand UO_1815 (O_1815,N_49701,N_49819);
xor UO_1816 (O_1816,N_49773,N_49857);
or UO_1817 (O_1817,N_49585,N_49714);
and UO_1818 (O_1818,N_49649,N_49566);
or UO_1819 (O_1819,N_49738,N_49867);
nand UO_1820 (O_1820,N_49616,N_49988);
or UO_1821 (O_1821,N_49633,N_49755);
nor UO_1822 (O_1822,N_49627,N_49657);
xor UO_1823 (O_1823,N_49732,N_49889);
or UO_1824 (O_1824,N_49638,N_49758);
and UO_1825 (O_1825,N_49629,N_49619);
nor UO_1826 (O_1826,N_49740,N_49610);
nand UO_1827 (O_1827,N_49824,N_49737);
nor UO_1828 (O_1828,N_49714,N_49887);
and UO_1829 (O_1829,N_49868,N_49524);
or UO_1830 (O_1830,N_49618,N_49909);
nand UO_1831 (O_1831,N_49866,N_49567);
xor UO_1832 (O_1832,N_49896,N_49642);
xnor UO_1833 (O_1833,N_49849,N_49987);
and UO_1834 (O_1834,N_49767,N_49792);
xnor UO_1835 (O_1835,N_49735,N_49639);
or UO_1836 (O_1836,N_49821,N_49635);
xnor UO_1837 (O_1837,N_49864,N_49649);
nor UO_1838 (O_1838,N_49831,N_49837);
nand UO_1839 (O_1839,N_49915,N_49952);
or UO_1840 (O_1840,N_49541,N_49888);
or UO_1841 (O_1841,N_49565,N_49807);
nor UO_1842 (O_1842,N_49962,N_49798);
nor UO_1843 (O_1843,N_49713,N_49580);
xor UO_1844 (O_1844,N_49793,N_49555);
nor UO_1845 (O_1845,N_49746,N_49638);
or UO_1846 (O_1846,N_49930,N_49983);
and UO_1847 (O_1847,N_49963,N_49748);
nand UO_1848 (O_1848,N_49807,N_49866);
or UO_1849 (O_1849,N_49545,N_49763);
nor UO_1850 (O_1850,N_49993,N_49613);
nand UO_1851 (O_1851,N_49738,N_49817);
xnor UO_1852 (O_1852,N_49673,N_49604);
xor UO_1853 (O_1853,N_49712,N_49914);
xnor UO_1854 (O_1854,N_49819,N_49880);
xnor UO_1855 (O_1855,N_49918,N_49799);
xnor UO_1856 (O_1856,N_49988,N_49971);
or UO_1857 (O_1857,N_49782,N_49915);
and UO_1858 (O_1858,N_49707,N_49872);
or UO_1859 (O_1859,N_49940,N_49783);
nor UO_1860 (O_1860,N_49893,N_49852);
xnor UO_1861 (O_1861,N_49927,N_49656);
nor UO_1862 (O_1862,N_49822,N_49676);
or UO_1863 (O_1863,N_49786,N_49935);
nor UO_1864 (O_1864,N_49956,N_49701);
xor UO_1865 (O_1865,N_49596,N_49734);
xor UO_1866 (O_1866,N_49889,N_49949);
nand UO_1867 (O_1867,N_49757,N_49593);
or UO_1868 (O_1868,N_49748,N_49687);
and UO_1869 (O_1869,N_49718,N_49780);
and UO_1870 (O_1870,N_49982,N_49763);
nor UO_1871 (O_1871,N_49918,N_49806);
or UO_1872 (O_1872,N_49581,N_49981);
nand UO_1873 (O_1873,N_49837,N_49942);
xor UO_1874 (O_1874,N_49937,N_49541);
xnor UO_1875 (O_1875,N_49512,N_49860);
xor UO_1876 (O_1876,N_49742,N_49880);
and UO_1877 (O_1877,N_49845,N_49627);
and UO_1878 (O_1878,N_49757,N_49587);
nor UO_1879 (O_1879,N_49716,N_49944);
nor UO_1880 (O_1880,N_49754,N_49691);
and UO_1881 (O_1881,N_49927,N_49911);
or UO_1882 (O_1882,N_49963,N_49573);
or UO_1883 (O_1883,N_49955,N_49533);
nand UO_1884 (O_1884,N_49538,N_49914);
and UO_1885 (O_1885,N_49930,N_49707);
nand UO_1886 (O_1886,N_49505,N_49510);
xnor UO_1887 (O_1887,N_49899,N_49938);
nor UO_1888 (O_1888,N_49627,N_49614);
and UO_1889 (O_1889,N_49654,N_49615);
xnor UO_1890 (O_1890,N_49655,N_49653);
nand UO_1891 (O_1891,N_49788,N_49900);
xor UO_1892 (O_1892,N_49833,N_49508);
and UO_1893 (O_1893,N_49728,N_49531);
nand UO_1894 (O_1894,N_49583,N_49940);
and UO_1895 (O_1895,N_49566,N_49692);
or UO_1896 (O_1896,N_49640,N_49599);
xnor UO_1897 (O_1897,N_49932,N_49976);
and UO_1898 (O_1898,N_49660,N_49838);
nor UO_1899 (O_1899,N_49548,N_49857);
or UO_1900 (O_1900,N_49572,N_49914);
and UO_1901 (O_1901,N_49792,N_49992);
nand UO_1902 (O_1902,N_49779,N_49841);
nor UO_1903 (O_1903,N_49771,N_49887);
nor UO_1904 (O_1904,N_49630,N_49656);
and UO_1905 (O_1905,N_49535,N_49938);
or UO_1906 (O_1906,N_49875,N_49758);
nor UO_1907 (O_1907,N_49716,N_49667);
nand UO_1908 (O_1908,N_49535,N_49629);
xor UO_1909 (O_1909,N_49995,N_49641);
nand UO_1910 (O_1910,N_49963,N_49834);
or UO_1911 (O_1911,N_49861,N_49933);
or UO_1912 (O_1912,N_49915,N_49676);
xor UO_1913 (O_1913,N_49917,N_49916);
nand UO_1914 (O_1914,N_49892,N_49768);
or UO_1915 (O_1915,N_49779,N_49893);
nand UO_1916 (O_1916,N_49618,N_49550);
nor UO_1917 (O_1917,N_49796,N_49695);
or UO_1918 (O_1918,N_49821,N_49879);
nand UO_1919 (O_1919,N_49538,N_49890);
or UO_1920 (O_1920,N_49836,N_49610);
and UO_1921 (O_1921,N_49527,N_49937);
and UO_1922 (O_1922,N_49914,N_49970);
or UO_1923 (O_1923,N_49935,N_49957);
or UO_1924 (O_1924,N_49924,N_49595);
and UO_1925 (O_1925,N_49875,N_49940);
and UO_1926 (O_1926,N_49511,N_49897);
nand UO_1927 (O_1927,N_49601,N_49701);
and UO_1928 (O_1928,N_49603,N_49788);
and UO_1929 (O_1929,N_49911,N_49586);
nand UO_1930 (O_1930,N_49865,N_49802);
and UO_1931 (O_1931,N_49807,N_49977);
nand UO_1932 (O_1932,N_49502,N_49823);
or UO_1933 (O_1933,N_49780,N_49753);
xnor UO_1934 (O_1934,N_49637,N_49682);
and UO_1935 (O_1935,N_49667,N_49793);
xor UO_1936 (O_1936,N_49654,N_49750);
and UO_1937 (O_1937,N_49580,N_49772);
and UO_1938 (O_1938,N_49834,N_49936);
nand UO_1939 (O_1939,N_49848,N_49718);
and UO_1940 (O_1940,N_49704,N_49608);
nor UO_1941 (O_1941,N_49578,N_49702);
xnor UO_1942 (O_1942,N_49857,N_49617);
and UO_1943 (O_1943,N_49529,N_49536);
nand UO_1944 (O_1944,N_49983,N_49538);
nand UO_1945 (O_1945,N_49966,N_49955);
nor UO_1946 (O_1946,N_49717,N_49649);
and UO_1947 (O_1947,N_49863,N_49759);
xnor UO_1948 (O_1948,N_49657,N_49690);
nand UO_1949 (O_1949,N_49685,N_49739);
and UO_1950 (O_1950,N_49583,N_49634);
and UO_1951 (O_1951,N_49856,N_49664);
and UO_1952 (O_1952,N_49723,N_49742);
and UO_1953 (O_1953,N_49967,N_49604);
nor UO_1954 (O_1954,N_49589,N_49581);
nand UO_1955 (O_1955,N_49955,N_49953);
xnor UO_1956 (O_1956,N_49703,N_49975);
or UO_1957 (O_1957,N_49519,N_49916);
nor UO_1958 (O_1958,N_49551,N_49936);
nor UO_1959 (O_1959,N_49744,N_49657);
nand UO_1960 (O_1960,N_49943,N_49889);
nand UO_1961 (O_1961,N_49573,N_49882);
nand UO_1962 (O_1962,N_49658,N_49989);
nand UO_1963 (O_1963,N_49635,N_49993);
and UO_1964 (O_1964,N_49957,N_49615);
nand UO_1965 (O_1965,N_49542,N_49887);
or UO_1966 (O_1966,N_49564,N_49799);
and UO_1967 (O_1967,N_49625,N_49876);
and UO_1968 (O_1968,N_49759,N_49934);
or UO_1969 (O_1969,N_49966,N_49897);
xor UO_1970 (O_1970,N_49698,N_49505);
nand UO_1971 (O_1971,N_49609,N_49622);
and UO_1972 (O_1972,N_49904,N_49706);
nand UO_1973 (O_1973,N_49691,N_49539);
and UO_1974 (O_1974,N_49500,N_49657);
xor UO_1975 (O_1975,N_49936,N_49839);
xnor UO_1976 (O_1976,N_49761,N_49682);
and UO_1977 (O_1977,N_49658,N_49668);
nand UO_1978 (O_1978,N_49718,N_49586);
nand UO_1979 (O_1979,N_49702,N_49582);
nor UO_1980 (O_1980,N_49939,N_49830);
or UO_1981 (O_1981,N_49786,N_49998);
and UO_1982 (O_1982,N_49623,N_49722);
xor UO_1983 (O_1983,N_49808,N_49866);
xnor UO_1984 (O_1984,N_49686,N_49664);
and UO_1985 (O_1985,N_49621,N_49761);
or UO_1986 (O_1986,N_49730,N_49625);
xor UO_1987 (O_1987,N_49528,N_49606);
nand UO_1988 (O_1988,N_49765,N_49843);
nor UO_1989 (O_1989,N_49879,N_49845);
and UO_1990 (O_1990,N_49857,N_49992);
nand UO_1991 (O_1991,N_49674,N_49615);
xor UO_1992 (O_1992,N_49690,N_49934);
and UO_1993 (O_1993,N_49983,N_49594);
nand UO_1994 (O_1994,N_49916,N_49908);
nand UO_1995 (O_1995,N_49977,N_49821);
and UO_1996 (O_1996,N_49796,N_49652);
or UO_1997 (O_1997,N_49592,N_49797);
xor UO_1998 (O_1998,N_49626,N_49503);
nand UO_1999 (O_1999,N_49838,N_49821);
xnor UO_2000 (O_2000,N_49607,N_49908);
and UO_2001 (O_2001,N_49740,N_49753);
nand UO_2002 (O_2002,N_49818,N_49662);
and UO_2003 (O_2003,N_49942,N_49761);
and UO_2004 (O_2004,N_49912,N_49648);
or UO_2005 (O_2005,N_49521,N_49659);
nor UO_2006 (O_2006,N_49619,N_49613);
and UO_2007 (O_2007,N_49933,N_49937);
or UO_2008 (O_2008,N_49521,N_49902);
nor UO_2009 (O_2009,N_49606,N_49594);
and UO_2010 (O_2010,N_49537,N_49586);
and UO_2011 (O_2011,N_49505,N_49881);
nand UO_2012 (O_2012,N_49820,N_49677);
nor UO_2013 (O_2013,N_49899,N_49605);
nor UO_2014 (O_2014,N_49536,N_49676);
nand UO_2015 (O_2015,N_49642,N_49805);
nor UO_2016 (O_2016,N_49716,N_49536);
nand UO_2017 (O_2017,N_49827,N_49641);
and UO_2018 (O_2018,N_49806,N_49540);
xnor UO_2019 (O_2019,N_49784,N_49715);
nor UO_2020 (O_2020,N_49883,N_49654);
nor UO_2021 (O_2021,N_49594,N_49768);
nand UO_2022 (O_2022,N_49993,N_49919);
and UO_2023 (O_2023,N_49992,N_49634);
xnor UO_2024 (O_2024,N_49981,N_49783);
nand UO_2025 (O_2025,N_49965,N_49955);
xor UO_2026 (O_2026,N_49852,N_49697);
nor UO_2027 (O_2027,N_49648,N_49662);
and UO_2028 (O_2028,N_49972,N_49951);
or UO_2029 (O_2029,N_49504,N_49548);
nor UO_2030 (O_2030,N_49527,N_49513);
nand UO_2031 (O_2031,N_49554,N_49989);
or UO_2032 (O_2032,N_49522,N_49668);
nor UO_2033 (O_2033,N_49611,N_49821);
nor UO_2034 (O_2034,N_49741,N_49856);
nand UO_2035 (O_2035,N_49961,N_49868);
nor UO_2036 (O_2036,N_49981,N_49579);
xnor UO_2037 (O_2037,N_49784,N_49812);
or UO_2038 (O_2038,N_49590,N_49930);
and UO_2039 (O_2039,N_49922,N_49509);
and UO_2040 (O_2040,N_49628,N_49598);
and UO_2041 (O_2041,N_49662,N_49642);
nand UO_2042 (O_2042,N_49798,N_49617);
xor UO_2043 (O_2043,N_49849,N_49786);
nand UO_2044 (O_2044,N_49906,N_49504);
xor UO_2045 (O_2045,N_49853,N_49890);
nor UO_2046 (O_2046,N_49645,N_49780);
nor UO_2047 (O_2047,N_49659,N_49792);
nand UO_2048 (O_2048,N_49873,N_49608);
nor UO_2049 (O_2049,N_49826,N_49521);
nor UO_2050 (O_2050,N_49663,N_49587);
nor UO_2051 (O_2051,N_49872,N_49604);
or UO_2052 (O_2052,N_49500,N_49937);
or UO_2053 (O_2053,N_49509,N_49801);
or UO_2054 (O_2054,N_49750,N_49641);
nor UO_2055 (O_2055,N_49645,N_49673);
nor UO_2056 (O_2056,N_49875,N_49970);
xnor UO_2057 (O_2057,N_49872,N_49685);
xor UO_2058 (O_2058,N_49798,N_49939);
xor UO_2059 (O_2059,N_49522,N_49733);
nor UO_2060 (O_2060,N_49609,N_49694);
and UO_2061 (O_2061,N_49635,N_49942);
xnor UO_2062 (O_2062,N_49697,N_49713);
nor UO_2063 (O_2063,N_49519,N_49651);
nor UO_2064 (O_2064,N_49613,N_49828);
xnor UO_2065 (O_2065,N_49891,N_49645);
nand UO_2066 (O_2066,N_49686,N_49843);
xnor UO_2067 (O_2067,N_49501,N_49581);
nor UO_2068 (O_2068,N_49824,N_49912);
xnor UO_2069 (O_2069,N_49929,N_49711);
and UO_2070 (O_2070,N_49790,N_49834);
nor UO_2071 (O_2071,N_49996,N_49623);
nand UO_2072 (O_2072,N_49807,N_49573);
nand UO_2073 (O_2073,N_49721,N_49653);
and UO_2074 (O_2074,N_49739,N_49884);
nor UO_2075 (O_2075,N_49844,N_49726);
and UO_2076 (O_2076,N_49818,N_49632);
xnor UO_2077 (O_2077,N_49888,N_49849);
nor UO_2078 (O_2078,N_49853,N_49645);
or UO_2079 (O_2079,N_49714,N_49536);
and UO_2080 (O_2080,N_49962,N_49510);
nor UO_2081 (O_2081,N_49988,N_49534);
nor UO_2082 (O_2082,N_49588,N_49789);
nor UO_2083 (O_2083,N_49606,N_49884);
xor UO_2084 (O_2084,N_49795,N_49810);
nand UO_2085 (O_2085,N_49737,N_49906);
and UO_2086 (O_2086,N_49531,N_49963);
nand UO_2087 (O_2087,N_49863,N_49781);
and UO_2088 (O_2088,N_49725,N_49768);
or UO_2089 (O_2089,N_49782,N_49555);
and UO_2090 (O_2090,N_49939,N_49637);
and UO_2091 (O_2091,N_49657,N_49805);
nand UO_2092 (O_2092,N_49574,N_49592);
nand UO_2093 (O_2093,N_49743,N_49800);
or UO_2094 (O_2094,N_49625,N_49745);
xor UO_2095 (O_2095,N_49629,N_49513);
nor UO_2096 (O_2096,N_49662,N_49947);
and UO_2097 (O_2097,N_49929,N_49895);
and UO_2098 (O_2098,N_49748,N_49710);
nand UO_2099 (O_2099,N_49521,N_49848);
xnor UO_2100 (O_2100,N_49891,N_49970);
or UO_2101 (O_2101,N_49841,N_49610);
or UO_2102 (O_2102,N_49713,N_49578);
xor UO_2103 (O_2103,N_49933,N_49777);
nand UO_2104 (O_2104,N_49915,N_49778);
nand UO_2105 (O_2105,N_49795,N_49701);
nand UO_2106 (O_2106,N_49999,N_49893);
nand UO_2107 (O_2107,N_49565,N_49843);
or UO_2108 (O_2108,N_49648,N_49633);
nand UO_2109 (O_2109,N_49793,N_49928);
nand UO_2110 (O_2110,N_49560,N_49702);
nand UO_2111 (O_2111,N_49508,N_49949);
nand UO_2112 (O_2112,N_49592,N_49898);
and UO_2113 (O_2113,N_49808,N_49604);
nor UO_2114 (O_2114,N_49580,N_49594);
nand UO_2115 (O_2115,N_49714,N_49542);
nand UO_2116 (O_2116,N_49872,N_49907);
xor UO_2117 (O_2117,N_49706,N_49566);
or UO_2118 (O_2118,N_49693,N_49673);
or UO_2119 (O_2119,N_49811,N_49805);
nor UO_2120 (O_2120,N_49973,N_49720);
nor UO_2121 (O_2121,N_49503,N_49840);
xor UO_2122 (O_2122,N_49524,N_49551);
or UO_2123 (O_2123,N_49958,N_49694);
xor UO_2124 (O_2124,N_49607,N_49553);
xor UO_2125 (O_2125,N_49644,N_49699);
nand UO_2126 (O_2126,N_49866,N_49767);
nor UO_2127 (O_2127,N_49808,N_49839);
nor UO_2128 (O_2128,N_49878,N_49723);
xnor UO_2129 (O_2129,N_49982,N_49702);
and UO_2130 (O_2130,N_49712,N_49983);
and UO_2131 (O_2131,N_49867,N_49507);
nand UO_2132 (O_2132,N_49856,N_49722);
and UO_2133 (O_2133,N_49745,N_49816);
nand UO_2134 (O_2134,N_49554,N_49582);
nand UO_2135 (O_2135,N_49801,N_49831);
nor UO_2136 (O_2136,N_49773,N_49620);
or UO_2137 (O_2137,N_49504,N_49736);
nand UO_2138 (O_2138,N_49757,N_49512);
nand UO_2139 (O_2139,N_49715,N_49547);
and UO_2140 (O_2140,N_49921,N_49989);
nand UO_2141 (O_2141,N_49998,N_49895);
nor UO_2142 (O_2142,N_49818,N_49686);
xor UO_2143 (O_2143,N_49827,N_49613);
nor UO_2144 (O_2144,N_49698,N_49563);
xnor UO_2145 (O_2145,N_49867,N_49984);
or UO_2146 (O_2146,N_49633,N_49954);
nor UO_2147 (O_2147,N_49810,N_49782);
nand UO_2148 (O_2148,N_49749,N_49614);
and UO_2149 (O_2149,N_49793,N_49511);
and UO_2150 (O_2150,N_49618,N_49637);
and UO_2151 (O_2151,N_49641,N_49924);
and UO_2152 (O_2152,N_49512,N_49600);
nor UO_2153 (O_2153,N_49682,N_49784);
nand UO_2154 (O_2154,N_49746,N_49945);
and UO_2155 (O_2155,N_49803,N_49866);
nand UO_2156 (O_2156,N_49959,N_49708);
or UO_2157 (O_2157,N_49577,N_49979);
nand UO_2158 (O_2158,N_49513,N_49960);
nor UO_2159 (O_2159,N_49539,N_49923);
xor UO_2160 (O_2160,N_49672,N_49533);
and UO_2161 (O_2161,N_49911,N_49545);
nand UO_2162 (O_2162,N_49822,N_49975);
nor UO_2163 (O_2163,N_49920,N_49992);
xor UO_2164 (O_2164,N_49981,N_49588);
and UO_2165 (O_2165,N_49594,N_49524);
and UO_2166 (O_2166,N_49562,N_49568);
xor UO_2167 (O_2167,N_49934,N_49734);
nor UO_2168 (O_2168,N_49941,N_49714);
nand UO_2169 (O_2169,N_49932,N_49637);
nor UO_2170 (O_2170,N_49794,N_49679);
xor UO_2171 (O_2171,N_49645,N_49646);
xor UO_2172 (O_2172,N_49766,N_49947);
xor UO_2173 (O_2173,N_49853,N_49878);
nand UO_2174 (O_2174,N_49827,N_49983);
nand UO_2175 (O_2175,N_49729,N_49509);
xnor UO_2176 (O_2176,N_49841,N_49580);
nand UO_2177 (O_2177,N_49583,N_49638);
xor UO_2178 (O_2178,N_49936,N_49690);
and UO_2179 (O_2179,N_49874,N_49822);
and UO_2180 (O_2180,N_49786,N_49630);
and UO_2181 (O_2181,N_49759,N_49742);
nand UO_2182 (O_2182,N_49582,N_49564);
nand UO_2183 (O_2183,N_49580,N_49916);
nand UO_2184 (O_2184,N_49614,N_49830);
xnor UO_2185 (O_2185,N_49792,N_49703);
nand UO_2186 (O_2186,N_49503,N_49591);
nand UO_2187 (O_2187,N_49589,N_49953);
xor UO_2188 (O_2188,N_49595,N_49678);
nor UO_2189 (O_2189,N_49680,N_49693);
nand UO_2190 (O_2190,N_49842,N_49768);
xor UO_2191 (O_2191,N_49941,N_49709);
and UO_2192 (O_2192,N_49840,N_49950);
and UO_2193 (O_2193,N_49667,N_49708);
and UO_2194 (O_2194,N_49758,N_49995);
and UO_2195 (O_2195,N_49712,N_49788);
nand UO_2196 (O_2196,N_49621,N_49681);
nand UO_2197 (O_2197,N_49762,N_49736);
nor UO_2198 (O_2198,N_49596,N_49543);
nor UO_2199 (O_2199,N_49556,N_49520);
and UO_2200 (O_2200,N_49861,N_49731);
nand UO_2201 (O_2201,N_49926,N_49839);
nand UO_2202 (O_2202,N_49570,N_49730);
nand UO_2203 (O_2203,N_49660,N_49693);
xnor UO_2204 (O_2204,N_49776,N_49714);
or UO_2205 (O_2205,N_49810,N_49809);
nand UO_2206 (O_2206,N_49801,N_49936);
and UO_2207 (O_2207,N_49978,N_49742);
and UO_2208 (O_2208,N_49506,N_49790);
xor UO_2209 (O_2209,N_49546,N_49755);
or UO_2210 (O_2210,N_49872,N_49646);
and UO_2211 (O_2211,N_49739,N_49899);
xnor UO_2212 (O_2212,N_49877,N_49563);
nor UO_2213 (O_2213,N_49543,N_49779);
nor UO_2214 (O_2214,N_49988,N_49761);
and UO_2215 (O_2215,N_49604,N_49547);
nand UO_2216 (O_2216,N_49634,N_49900);
xor UO_2217 (O_2217,N_49972,N_49736);
xnor UO_2218 (O_2218,N_49582,N_49793);
and UO_2219 (O_2219,N_49606,N_49737);
and UO_2220 (O_2220,N_49833,N_49575);
xnor UO_2221 (O_2221,N_49986,N_49722);
nor UO_2222 (O_2222,N_49573,N_49805);
nand UO_2223 (O_2223,N_49749,N_49729);
or UO_2224 (O_2224,N_49550,N_49577);
xor UO_2225 (O_2225,N_49918,N_49996);
and UO_2226 (O_2226,N_49664,N_49786);
and UO_2227 (O_2227,N_49592,N_49528);
nor UO_2228 (O_2228,N_49950,N_49506);
or UO_2229 (O_2229,N_49873,N_49742);
and UO_2230 (O_2230,N_49506,N_49741);
nand UO_2231 (O_2231,N_49808,N_49978);
or UO_2232 (O_2232,N_49939,N_49647);
nor UO_2233 (O_2233,N_49775,N_49983);
nor UO_2234 (O_2234,N_49943,N_49865);
and UO_2235 (O_2235,N_49974,N_49798);
nand UO_2236 (O_2236,N_49707,N_49543);
xor UO_2237 (O_2237,N_49787,N_49985);
nor UO_2238 (O_2238,N_49516,N_49820);
and UO_2239 (O_2239,N_49810,N_49956);
nand UO_2240 (O_2240,N_49948,N_49818);
and UO_2241 (O_2241,N_49732,N_49986);
nand UO_2242 (O_2242,N_49544,N_49692);
and UO_2243 (O_2243,N_49566,N_49682);
xor UO_2244 (O_2244,N_49932,N_49902);
and UO_2245 (O_2245,N_49911,N_49936);
and UO_2246 (O_2246,N_49904,N_49509);
nor UO_2247 (O_2247,N_49555,N_49785);
and UO_2248 (O_2248,N_49513,N_49926);
or UO_2249 (O_2249,N_49682,N_49888);
nand UO_2250 (O_2250,N_49768,N_49613);
nand UO_2251 (O_2251,N_49931,N_49708);
nor UO_2252 (O_2252,N_49844,N_49585);
nor UO_2253 (O_2253,N_49809,N_49914);
and UO_2254 (O_2254,N_49529,N_49710);
and UO_2255 (O_2255,N_49773,N_49654);
nor UO_2256 (O_2256,N_49832,N_49606);
or UO_2257 (O_2257,N_49616,N_49793);
nor UO_2258 (O_2258,N_49612,N_49720);
nand UO_2259 (O_2259,N_49616,N_49800);
nor UO_2260 (O_2260,N_49870,N_49735);
or UO_2261 (O_2261,N_49501,N_49532);
xnor UO_2262 (O_2262,N_49876,N_49961);
or UO_2263 (O_2263,N_49537,N_49786);
xnor UO_2264 (O_2264,N_49704,N_49679);
or UO_2265 (O_2265,N_49983,N_49723);
nand UO_2266 (O_2266,N_49633,N_49539);
or UO_2267 (O_2267,N_49955,N_49717);
xor UO_2268 (O_2268,N_49587,N_49876);
or UO_2269 (O_2269,N_49837,N_49610);
or UO_2270 (O_2270,N_49923,N_49568);
or UO_2271 (O_2271,N_49744,N_49654);
nand UO_2272 (O_2272,N_49805,N_49934);
nor UO_2273 (O_2273,N_49774,N_49994);
nor UO_2274 (O_2274,N_49616,N_49649);
xor UO_2275 (O_2275,N_49898,N_49848);
nand UO_2276 (O_2276,N_49511,N_49509);
xor UO_2277 (O_2277,N_49621,N_49968);
nor UO_2278 (O_2278,N_49941,N_49562);
and UO_2279 (O_2279,N_49928,N_49987);
xor UO_2280 (O_2280,N_49777,N_49996);
xor UO_2281 (O_2281,N_49676,N_49749);
nand UO_2282 (O_2282,N_49624,N_49865);
nor UO_2283 (O_2283,N_49730,N_49720);
xnor UO_2284 (O_2284,N_49835,N_49865);
and UO_2285 (O_2285,N_49777,N_49832);
nand UO_2286 (O_2286,N_49932,N_49908);
nor UO_2287 (O_2287,N_49974,N_49583);
and UO_2288 (O_2288,N_49732,N_49604);
xnor UO_2289 (O_2289,N_49795,N_49671);
nand UO_2290 (O_2290,N_49856,N_49517);
and UO_2291 (O_2291,N_49879,N_49851);
xnor UO_2292 (O_2292,N_49677,N_49652);
nand UO_2293 (O_2293,N_49743,N_49787);
or UO_2294 (O_2294,N_49787,N_49611);
and UO_2295 (O_2295,N_49835,N_49682);
nor UO_2296 (O_2296,N_49542,N_49640);
nor UO_2297 (O_2297,N_49569,N_49700);
nor UO_2298 (O_2298,N_49668,N_49947);
xor UO_2299 (O_2299,N_49633,N_49640);
nand UO_2300 (O_2300,N_49953,N_49577);
nand UO_2301 (O_2301,N_49562,N_49970);
xor UO_2302 (O_2302,N_49951,N_49730);
nor UO_2303 (O_2303,N_49594,N_49788);
nand UO_2304 (O_2304,N_49598,N_49728);
or UO_2305 (O_2305,N_49599,N_49968);
and UO_2306 (O_2306,N_49849,N_49859);
nor UO_2307 (O_2307,N_49625,N_49666);
nand UO_2308 (O_2308,N_49860,N_49509);
nor UO_2309 (O_2309,N_49864,N_49956);
nand UO_2310 (O_2310,N_49788,N_49657);
or UO_2311 (O_2311,N_49911,N_49882);
nor UO_2312 (O_2312,N_49746,N_49951);
nor UO_2313 (O_2313,N_49655,N_49661);
xnor UO_2314 (O_2314,N_49823,N_49746);
nand UO_2315 (O_2315,N_49519,N_49945);
or UO_2316 (O_2316,N_49703,N_49702);
nand UO_2317 (O_2317,N_49628,N_49860);
nor UO_2318 (O_2318,N_49677,N_49633);
and UO_2319 (O_2319,N_49516,N_49588);
xnor UO_2320 (O_2320,N_49572,N_49738);
xor UO_2321 (O_2321,N_49770,N_49823);
or UO_2322 (O_2322,N_49980,N_49732);
nand UO_2323 (O_2323,N_49607,N_49648);
nor UO_2324 (O_2324,N_49942,N_49708);
xor UO_2325 (O_2325,N_49908,N_49889);
nand UO_2326 (O_2326,N_49632,N_49835);
nand UO_2327 (O_2327,N_49552,N_49674);
or UO_2328 (O_2328,N_49933,N_49669);
and UO_2329 (O_2329,N_49723,N_49693);
xnor UO_2330 (O_2330,N_49586,N_49877);
nor UO_2331 (O_2331,N_49996,N_49654);
and UO_2332 (O_2332,N_49614,N_49971);
xor UO_2333 (O_2333,N_49691,N_49513);
nor UO_2334 (O_2334,N_49842,N_49891);
and UO_2335 (O_2335,N_49874,N_49825);
and UO_2336 (O_2336,N_49945,N_49809);
nor UO_2337 (O_2337,N_49761,N_49571);
nor UO_2338 (O_2338,N_49503,N_49816);
and UO_2339 (O_2339,N_49527,N_49830);
or UO_2340 (O_2340,N_49894,N_49952);
nand UO_2341 (O_2341,N_49599,N_49740);
nand UO_2342 (O_2342,N_49631,N_49727);
nor UO_2343 (O_2343,N_49723,N_49705);
xnor UO_2344 (O_2344,N_49892,N_49823);
nand UO_2345 (O_2345,N_49721,N_49943);
and UO_2346 (O_2346,N_49583,N_49764);
xnor UO_2347 (O_2347,N_49826,N_49748);
and UO_2348 (O_2348,N_49776,N_49578);
and UO_2349 (O_2349,N_49683,N_49622);
or UO_2350 (O_2350,N_49775,N_49835);
nand UO_2351 (O_2351,N_49923,N_49709);
xnor UO_2352 (O_2352,N_49829,N_49705);
nor UO_2353 (O_2353,N_49988,N_49898);
nor UO_2354 (O_2354,N_49509,N_49952);
and UO_2355 (O_2355,N_49508,N_49635);
and UO_2356 (O_2356,N_49801,N_49793);
xor UO_2357 (O_2357,N_49819,N_49525);
nor UO_2358 (O_2358,N_49672,N_49964);
and UO_2359 (O_2359,N_49977,N_49577);
and UO_2360 (O_2360,N_49576,N_49591);
xor UO_2361 (O_2361,N_49705,N_49918);
or UO_2362 (O_2362,N_49762,N_49862);
or UO_2363 (O_2363,N_49715,N_49944);
and UO_2364 (O_2364,N_49672,N_49740);
nand UO_2365 (O_2365,N_49695,N_49942);
or UO_2366 (O_2366,N_49612,N_49542);
or UO_2367 (O_2367,N_49847,N_49870);
and UO_2368 (O_2368,N_49802,N_49841);
nand UO_2369 (O_2369,N_49505,N_49645);
or UO_2370 (O_2370,N_49926,N_49857);
nand UO_2371 (O_2371,N_49506,N_49514);
xor UO_2372 (O_2372,N_49801,N_49728);
nor UO_2373 (O_2373,N_49993,N_49767);
and UO_2374 (O_2374,N_49983,N_49834);
nand UO_2375 (O_2375,N_49591,N_49811);
xor UO_2376 (O_2376,N_49519,N_49553);
nand UO_2377 (O_2377,N_49592,N_49740);
xnor UO_2378 (O_2378,N_49679,N_49681);
or UO_2379 (O_2379,N_49784,N_49967);
or UO_2380 (O_2380,N_49609,N_49672);
or UO_2381 (O_2381,N_49865,N_49922);
nor UO_2382 (O_2382,N_49526,N_49819);
xor UO_2383 (O_2383,N_49735,N_49888);
nor UO_2384 (O_2384,N_49785,N_49812);
and UO_2385 (O_2385,N_49605,N_49870);
nor UO_2386 (O_2386,N_49901,N_49830);
nor UO_2387 (O_2387,N_49795,N_49641);
or UO_2388 (O_2388,N_49650,N_49978);
or UO_2389 (O_2389,N_49968,N_49500);
or UO_2390 (O_2390,N_49551,N_49698);
and UO_2391 (O_2391,N_49914,N_49632);
or UO_2392 (O_2392,N_49558,N_49920);
nand UO_2393 (O_2393,N_49798,N_49666);
nand UO_2394 (O_2394,N_49534,N_49558);
or UO_2395 (O_2395,N_49936,N_49930);
or UO_2396 (O_2396,N_49577,N_49735);
xnor UO_2397 (O_2397,N_49755,N_49556);
and UO_2398 (O_2398,N_49767,N_49747);
xnor UO_2399 (O_2399,N_49773,N_49884);
xnor UO_2400 (O_2400,N_49781,N_49724);
nor UO_2401 (O_2401,N_49792,N_49737);
or UO_2402 (O_2402,N_49695,N_49948);
or UO_2403 (O_2403,N_49942,N_49583);
xnor UO_2404 (O_2404,N_49703,N_49909);
nor UO_2405 (O_2405,N_49779,N_49636);
xnor UO_2406 (O_2406,N_49527,N_49996);
nor UO_2407 (O_2407,N_49593,N_49846);
and UO_2408 (O_2408,N_49784,N_49656);
nor UO_2409 (O_2409,N_49918,N_49782);
nor UO_2410 (O_2410,N_49951,N_49656);
and UO_2411 (O_2411,N_49777,N_49679);
nand UO_2412 (O_2412,N_49907,N_49541);
or UO_2413 (O_2413,N_49533,N_49537);
and UO_2414 (O_2414,N_49903,N_49763);
nor UO_2415 (O_2415,N_49982,N_49710);
and UO_2416 (O_2416,N_49859,N_49825);
and UO_2417 (O_2417,N_49961,N_49567);
and UO_2418 (O_2418,N_49642,N_49521);
and UO_2419 (O_2419,N_49501,N_49972);
nand UO_2420 (O_2420,N_49645,N_49695);
xnor UO_2421 (O_2421,N_49811,N_49654);
or UO_2422 (O_2422,N_49797,N_49551);
and UO_2423 (O_2423,N_49696,N_49504);
and UO_2424 (O_2424,N_49645,N_49587);
or UO_2425 (O_2425,N_49715,N_49806);
or UO_2426 (O_2426,N_49958,N_49733);
nand UO_2427 (O_2427,N_49705,N_49500);
and UO_2428 (O_2428,N_49950,N_49639);
or UO_2429 (O_2429,N_49671,N_49754);
nand UO_2430 (O_2430,N_49606,N_49834);
nand UO_2431 (O_2431,N_49834,N_49881);
nor UO_2432 (O_2432,N_49787,N_49862);
nand UO_2433 (O_2433,N_49764,N_49818);
nor UO_2434 (O_2434,N_49839,N_49948);
nand UO_2435 (O_2435,N_49630,N_49911);
and UO_2436 (O_2436,N_49973,N_49532);
nand UO_2437 (O_2437,N_49984,N_49790);
xnor UO_2438 (O_2438,N_49615,N_49980);
xnor UO_2439 (O_2439,N_49687,N_49598);
nand UO_2440 (O_2440,N_49758,N_49998);
or UO_2441 (O_2441,N_49961,N_49895);
and UO_2442 (O_2442,N_49622,N_49842);
nor UO_2443 (O_2443,N_49895,N_49513);
xor UO_2444 (O_2444,N_49827,N_49806);
nand UO_2445 (O_2445,N_49678,N_49994);
or UO_2446 (O_2446,N_49743,N_49840);
and UO_2447 (O_2447,N_49687,N_49648);
or UO_2448 (O_2448,N_49817,N_49728);
xnor UO_2449 (O_2449,N_49512,N_49969);
and UO_2450 (O_2450,N_49887,N_49738);
xor UO_2451 (O_2451,N_49792,N_49780);
nand UO_2452 (O_2452,N_49573,N_49516);
xor UO_2453 (O_2453,N_49661,N_49571);
or UO_2454 (O_2454,N_49745,N_49630);
nor UO_2455 (O_2455,N_49506,N_49590);
or UO_2456 (O_2456,N_49812,N_49988);
xnor UO_2457 (O_2457,N_49852,N_49988);
and UO_2458 (O_2458,N_49869,N_49521);
nand UO_2459 (O_2459,N_49622,N_49790);
nor UO_2460 (O_2460,N_49541,N_49872);
and UO_2461 (O_2461,N_49717,N_49763);
or UO_2462 (O_2462,N_49519,N_49518);
or UO_2463 (O_2463,N_49633,N_49850);
and UO_2464 (O_2464,N_49970,N_49763);
xor UO_2465 (O_2465,N_49735,N_49872);
and UO_2466 (O_2466,N_49778,N_49777);
nor UO_2467 (O_2467,N_49834,N_49700);
nor UO_2468 (O_2468,N_49735,N_49646);
or UO_2469 (O_2469,N_49653,N_49642);
nand UO_2470 (O_2470,N_49941,N_49984);
nor UO_2471 (O_2471,N_49957,N_49916);
or UO_2472 (O_2472,N_49818,N_49580);
nand UO_2473 (O_2473,N_49636,N_49910);
nand UO_2474 (O_2474,N_49744,N_49786);
and UO_2475 (O_2475,N_49921,N_49889);
xor UO_2476 (O_2476,N_49723,N_49846);
xor UO_2477 (O_2477,N_49968,N_49639);
or UO_2478 (O_2478,N_49502,N_49925);
xor UO_2479 (O_2479,N_49775,N_49951);
nand UO_2480 (O_2480,N_49681,N_49941);
or UO_2481 (O_2481,N_49940,N_49575);
nor UO_2482 (O_2482,N_49879,N_49621);
nand UO_2483 (O_2483,N_49658,N_49660);
and UO_2484 (O_2484,N_49895,N_49826);
or UO_2485 (O_2485,N_49973,N_49601);
nand UO_2486 (O_2486,N_49844,N_49924);
or UO_2487 (O_2487,N_49716,N_49749);
xor UO_2488 (O_2488,N_49924,N_49685);
xor UO_2489 (O_2489,N_49728,N_49979);
nor UO_2490 (O_2490,N_49608,N_49883);
nor UO_2491 (O_2491,N_49782,N_49756);
xnor UO_2492 (O_2492,N_49806,N_49609);
nand UO_2493 (O_2493,N_49822,N_49846);
xor UO_2494 (O_2494,N_49732,N_49898);
xor UO_2495 (O_2495,N_49535,N_49510);
nand UO_2496 (O_2496,N_49530,N_49698);
xnor UO_2497 (O_2497,N_49835,N_49646);
nor UO_2498 (O_2498,N_49745,N_49758);
xor UO_2499 (O_2499,N_49931,N_49768);
or UO_2500 (O_2500,N_49756,N_49584);
or UO_2501 (O_2501,N_49510,N_49835);
or UO_2502 (O_2502,N_49835,N_49844);
and UO_2503 (O_2503,N_49700,N_49866);
xnor UO_2504 (O_2504,N_49938,N_49735);
or UO_2505 (O_2505,N_49518,N_49650);
nor UO_2506 (O_2506,N_49783,N_49904);
and UO_2507 (O_2507,N_49911,N_49799);
and UO_2508 (O_2508,N_49614,N_49727);
nor UO_2509 (O_2509,N_49564,N_49717);
xor UO_2510 (O_2510,N_49719,N_49551);
and UO_2511 (O_2511,N_49627,N_49615);
and UO_2512 (O_2512,N_49634,N_49764);
xnor UO_2513 (O_2513,N_49986,N_49977);
xor UO_2514 (O_2514,N_49508,N_49659);
or UO_2515 (O_2515,N_49527,N_49561);
nor UO_2516 (O_2516,N_49849,N_49712);
nor UO_2517 (O_2517,N_49738,N_49613);
nor UO_2518 (O_2518,N_49621,N_49700);
and UO_2519 (O_2519,N_49713,N_49874);
xnor UO_2520 (O_2520,N_49805,N_49640);
or UO_2521 (O_2521,N_49733,N_49939);
nand UO_2522 (O_2522,N_49535,N_49742);
xor UO_2523 (O_2523,N_49771,N_49893);
nand UO_2524 (O_2524,N_49895,N_49525);
nand UO_2525 (O_2525,N_49600,N_49855);
nor UO_2526 (O_2526,N_49772,N_49936);
xor UO_2527 (O_2527,N_49580,N_49965);
nand UO_2528 (O_2528,N_49868,N_49862);
or UO_2529 (O_2529,N_49641,N_49568);
and UO_2530 (O_2530,N_49881,N_49622);
nor UO_2531 (O_2531,N_49572,N_49855);
and UO_2532 (O_2532,N_49862,N_49932);
or UO_2533 (O_2533,N_49750,N_49689);
nor UO_2534 (O_2534,N_49593,N_49816);
nand UO_2535 (O_2535,N_49812,N_49875);
or UO_2536 (O_2536,N_49616,N_49861);
nor UO_2537 (O_2537,N_49602,N_49760);
nor UO_2538 (O_2538,N_49663,N_49637);
xor UO_2539 (O_2539,N_49685,N_49970);
nand UO_2540 (O_2540,N_49636,N_49583);
nand UO_2541 (O_2541,N_49610,N_49908);
nor UO_2542 (O_2542,N_49610,N_49592);
xnor UO_2543 (O_2543,N_49792,N_49674);
xnor UO_2544 (O_2544,N_49863,N_49716);
nand UO_2545 (O_2545,N_49670,N_49548);
nand UO_2546 (O_2546,N_49850,N_49911);
or UO_2547 (O_2547,N_49535,N_49621);
and UO_2548 (O_2548,N_49566,N_49556);
or UO_2549 (O_2549,N_49745,N_49619);
and UO_2550 (O_2550,N_49739,N_49799);
and UO_2551 (O_2551,N_49824,N_49651);
and UO_2552 (O_2552,N_49912,N_49588);
xor UO_2553 (O_2553,N_49564,N_49792);
nand UO_2554 (O_2554,N_49650,N_49574);
and UO_2555 (O_2555,N_49812,N_49810);
nand UO_2556 (O_2556,N_49824,N_49865);
nand UO_2557 (O_2557,N_49951,N_49829);
nor UO_2558 (O_2558,N_49749,N_49924);
nor UO_2559 (O_2559,N_49690,N_49845);
nor UO_2560 (O_2560,N_49603,N_49512);
and UO_2561 (O_2561,N_49897,N_49559);
and UO_2562 (O_2562,N_49890,N_49827);
xnor UO_2563 (O_2563,N_49889,N_49890);
or UO_2564 (O_2564,N_49603,N_49577);
nand UO_2565 (O_2565,N_49970,N_49624);
nand UO_2566 (O_2566,N_49759,N_49917);
xnor UO_2567 (O_2567,N_49940,N_49757);
nor UO_2568 (O_2568,N_49644,N_49777);
or UO_2569 (O_2569,N_49667,N_49546);
xnor UO_2570 (O_2570,N_49641,N_49831);
nand UO_2571 (O_2571,N_49565,N_49976);
xor UO_2572 (O_2572,N_49593,N_49700);
and UO_2573 (O_2573,N_49546,N_49729);
xor UO_2574 (O_2574,N_49604,N_49774);
nand UO_2575 (O_2575,N_49984,N_49506);
nand UO_2576 (O_2576,N_49806,N_49658);
nand UO_2577 (O_2577,N_49833,N_49561);
xnor UO_2578 (O_2578,N_49965,N_49540);
xnor UO_2579 (O_2579,N_49612,N_49733);
xnor UO_2580 (O_2580,N_49870,N_49679);
or UO_2581 (O_2581,N_49768,N_49525);
or UO_2582 (O_2582,N_49781,N_49599);
xnor UO_2583 (O_2583,N_49758,N_49684);
or UO_2584 (O_2584,N_49861,N_49515);
or UO_2585 (O_2585,N_49982,N_49547);
and UO_2586 (O_2586,N_49628,N_49822);
nor UO_2587 (O_2587,N_49958,N_49916);
and UO_2588 (O_2588,N_49796,N_49836);
nor UO_2589 (O_2589,N_49970,N_49583);
nand UO_2590 (O_2590,N_49511,N_49697);
xnor UO_2591 (O_2591,N_49608,N_49856);
or UO_2592 (O_2592,N_49988,N_49887);
xnor UO_2593 (O_2593,N_49587,N_49812);
nor UO_2594 (O_2594,N_49764,N_49561);
xnor UO_2595 (O_2595,N_49556,N_49954);
and UO_2596 (O_2596,N_49973,N_49627);
and UO_2597 (O_2597,N_49609,N_49916);
xor UO_2598 (O_2598,N_49905,N_49995);
or UO_2599 (O_2599,N_49574,N_49657);
or UO_2600 (O_2600,N_49947,N_49631);
nand UO_2601 (O_2601,N_49835,N_49608);
xnor UO_2602 (O_2602,N_49999,N_49843);
or UO_2603 (O_2603,N_49610,N_49687);
nand UO_2604 (O_2604,N_49819,N_49963);
and UO_2605 (O_2605,N_49819,N_49810);
xnor UO_2606 (O_2606,N_49744,N_49958);
xnor UO_2607 (O_2607,N_49715,N_49556);
nor UO_2608 (O_2608,N_49640,N_49840);
nand UO_2609 (O_2609,N_49980,N_49650);
or UO_2610 (O_2610,N_49665,N_49684);
or UO_2611 (O_2611,N_49657,N_49724);
or UO_2612 (O_2612,N_49866,N_49670);
nand UO_2613 (O_2613,N_49849,N_49664);
and UO_2614 (O_2614,N_49708,N_49800);
or UO_2615 (O_2615,N_49997,N_49526);
nand UO_2616 (O_2616,N_49982,N_49789);
nand UO_2617 (O_2617,N_49878,N_49815);
xor UO_2618 (O_2618,N_49808,N_49664);
xor UO_2619 (O_2619,N_49618,N_49841);
xnor UO_2620 (O_2620,N_49583,N_49713);
xor UO_2621 (O_2621,N_49900,N_49660);
or UO_2622 (O_2622,N_49764,N_49587);
or UO_2623 (O_2623,N_49576,N_49909);
nor UO_2624 (O_2624,N_49736,N_49924);
nand UO_2625 (O_2625,N_49736,N_49749);
xnor UO_2626 (O_2626,N_49578,N_49767);
and UO_2627 (O_2627,N_49876,N_49700);
and UO_2628 (O_2628,N_49554,N_49804);
or UO_2629 (O_2629,N_49900,N_49555);
nor UO_2630 (O_2630,N_49671,N_49957);
xor UO_2631 (O_2631,N_49555,N_49988);
xor UO_2632 (O_2632,N_49529,N_49674);
nand UO_2633 (O_2633,N_49871,N_49706);
nor UO_2634 (O_2634,N_49655,N_49676);
and UO_2635 (O_2635,N_49558,N_49687);
xor UO_2636 (O_2636,N_49897,N_49883);
nor UO_2637 (O_2637,N_49672,N_49725);
and UO_2638 (O_2638,N_49997,N_49963);
nand UO_2639 (O_2639,N_49922,N_49781);
and UO_2640 (O_2640,N_49761,N_49712);
nor UO_2641 (O_2641,N_49870,N_49741);
or UO_2642 (O_2642,N_49514,N_49927);
or UO_2643 (O_2643,N_49675,N_49807);
xor UO_2644 (O_2644,N_49864,N_49736);
and UO_2645 (O_2645,N_49797,N_49610);
xnor UO_2646 (O_2646,N_49693,N_49519);
or UO_2647 (O_2647,N_49659,N_49662);
xnor UO_2648 (O_2648,N_49944,N_49617);
nor UO_2649 (O_2649,N_49550,N_49753);
nor UO_2650 (O_2650,N_49776,N_49734);
and UO_2651 (O_2651,N_49553,N_49646);
or UO_2652 (O_2652,N_49852,N_49556);
nor UO_2653 (O_2653,N_49672,N_49977);
nor UO_2654 (O_2654,N_49519,N_49619);
nor UO_2655 (O_2655,N_49501,N_49695);
and UO_2656 (O_2656,N_49825,N_49923);
nor UO_2657 (O_2657,N_49737,N_49647);
and UO_2658 (O_2658,N_49606,N_49575);
xor UO_2659 (O_2659,N_49574,N_49756);
nor UO_2660 (O_2660,N_49613,N_49549);
and UO_2661 (O_2661,N_49824,N_49834);
nand UO_2662 (O_2662,N_49979,N_49913);
nor UO_2663 (O_2663,N_49620,N_49674);
nor UO_2664 (O_2664,N_49894,N_49513);
and UO_2665 (O_2665,N_49965,N_49522);
nor UO_2666 (O_2666,N_49949,N_49518);
and UO_2667 (O_2667,N_49896,N_49738);
nor UO_2668 (O_2668,N_49657,N_49686);
or UO_2669 (O_2669,N_49802,N_49961);
nor UO_2670 (O_2670,N_49740,N_49858);
and UO_2671 (O_2671,N_49920,N_49559);
nand UO_2672 (O_2672,N_49526,N_49548);
or UO_2673 (O_2673,N_49988,N_49806);
nand UO_2674 (O_2674,N_49817,N_49791);
and UO_2675 (O_2675,N_49525,N_49515);
or UO_2676 (O_2676,N_49755,N_49639);
nand UO_2677 (O_2677,N_49653,N_49766);
nor UO_2678 (O_2678,N_49866,N_49663);
xnor UO_2679 (O_2679,N_49823,N_49535);
xor UO_2680 (O_2680,N_49694,N_49906);
nand UO_2681 (O_2681,N_49641,N_49741);
nand UO_2682 (O_2682,N_49919,N_49711);
nor UO_2683 (O_2683,N_49878,N_49903);
xor UO_2684 (O_2684,N_49932,N_49979);
nor UO_2685 (O_2685,N_49842,N_49502);
nand UO_2686 (O_2686,N_49861,N_49990);
and UO_2687 (O_2687,N_49758,N_49704);
or UO_2688 (O_2688,N_49652,N_49565);
or UO_2689 (O_2689,N_49943,N_49900);
or UO_2690 (O_2690,N_49872,N_49621);
or UO_2691 (O_2691,N_49632,N_49986);
or UO_2692 (O_2692,N_49961,N_49542);
nor UO_2693 (O_2693,N_49766,N_49652);
or UO_2694 (O_2694,N_49529,N_49831);
and UO_2695 (O_2695,N_49922,N_49639);
or UO_2696 (O_2696,N_49878,N_49986);
or UO_2697 (O_2697,N_49541,N_49901);
xnor UO_2698 (O_2698,N_49817,N_49645);
nand UO_2699 (O_2699,N_49750,N_49505);
xnor UO_2700 (O_2700,N_49875,N_49644);
or UO_2701 (O_2701,N_49922,N_49890);
or UO_2702 (O_2702,N_49689,N_49988);
nor UO_2703 (O_2703,N_49818,N_49726);
xor UO_2704 (O_2704,N_49840,N_49554);
xor UO_2705 (O_2705,N_49642,N_49820);
nor UO_2706 (O_2706,N_49757,N_49907);
and UO_2707 (O_2707,N_49840,N_49910);
or UO_2708 (O_2708,N_49932,N_49745);
and UO_2709 (O_2709,N_49838,N_49846);
nand UO_2710 (O_2710,N_49576,N_49564);
and UO_2711 (O_2711,N_49515,N_49604);
nand UO_2712 (O_2712,N_49890,N_49558);
nor UO_2713 (O_2713,N_49599,N_49847);
nand UO_2714 (O_2714,N_49598,N_49940);
or UO_2715 (O_2715,N_49661,N_49844);
nor UO_2716 (O_2716,N_49868,N_49948);
nand UO_2717 (O_2717,N_49820,N_49987);
and UO_2718 (O_2718,N_49525,N_49704);
nand UO_2719 (O_2719,N_49601,N_49736);
or UO_2720 (O_2720,N_49725,N_49635);
xnor UO_2721 (O_2721,N_49582,N_49872);
xor UO_2722 (O_2722,N_49853,N_49786);
and UO_2723 (O_2723,N_49684,N_49949);
nor UO_2724 (O_2724,N_49836,N_49545);
nand UO_2725 (O_2725,N_49950,N_49583);
and UO_2726 (O_2726,N_49923,N_49706);
nor UO_2727 (O_2727,N_49931,N_49860);
or UO_2728 (O_2728,N_49925,N_49737);
nand UO_2729 (O_2729,N_49923,N_49723);
nor UO_2730 (O_2730,N_49895,N_49887);
and UO_2731 (O_2731,N_49628,N_49707);
nor UO_2732 (O_2732,N_49818,N_49896);
xor UO_2733 (O_2733,N_49947,N_49988);
and UO_2734 (O_2734,N_49897,N_49539);
or UO_2735 (O_2735,N_49511,N_49785);
and UO_2736 (O_2736,N_49526,N_49901);
nor UO_2737 (O_2737,N_49809,N_49739);
and UO_2738 (O_2738,N_49603,N_49802);
or UO_2739 (O_2739,N_49841,N_49903);
nor UO_2740 (O_2740,N_49757,N_49829);
nand UO_2741 (O_2741,N_49585,N_49734);
nand UO_2742 (O_2742,N_49540,N_49617);
nand UO_2743 (O_2743,N_49601,N_49855);
nor UO_2744 (O_2744,N_49824,N_49676);
xor UO_2745 (O_2745,N_49779,N_49885);
nand UO_2746 (O_2746,N_49911,N_49982);
xnor UO_2747 (O_2747,N_49629,N_49541);
and UO_2748 (O_2748,N_49756,N_49859);
xor UO_2749 (O_2749,N_49548,N_49691);
nand UO_2750 (O_2750,N_49670,N_49711);
or UO_2751 (O_2751,N_49961,N_49676);
nor UO_2752 (O_2752,N_49975,N_49730);
and UO_2753 (O_2753,N_49961,N_49902);
nor UO_2754 (O_2754,N_49568,N_49765);
or UO_2755 (O_2755,N_49855,N_49522);
or UO_2756 (O_2756,N_49884,N_49809);
xnor UO_2757 (O_2757,N_49903,N_49859);
nand UO_2758 (O_2758,N_49736,N_49681);
or UO_2759 (O_2759,N_49764,N_49907);
and UO_2760 (O_2760,N_49908,N_49801);
nor UO_2761 (O_2761,N_49715,N_49739);
and UO_2762 (O_2762,N_49755,N_49641);
nor UO_2763 (O_2763,N_49577,N_49551);
nor UO_2764 (O_2764,N_49615,N_49634);
nand UO_2765 (O_2765,N_49674,N_49839);
nor UO_2766 (O_2766,N_49594,N_49552);
xor UO_2767 (O_2767,N_49923,N_49745);
xor UO_2768 (O_2768,N_49858,N_49594);
nor UO_2769 (O_2769,N_49797,N_49767);
xor UO_2770 (O_2770,N_49793,N_49753);
nor UO_2771 (O_2771,N_49709,N_49702);
or UO_2772 (O_2772,N_49912,N_49614);
and UO_2773 (O_2773,N_49591,N_49917);
nor UO_2774 (O_2774,N_49971,N_49640);
nand UO_2775 (O_2775,N_49576,N_49799);
or UO_2776 (O_2776,N_49767,N_49908);
or UO_2777 (O_2777,N_49734,N_49559);
xnor UO_2778 (O_2778,N_49807,N_49906);
xnor UO_2779 (O_2779,N_49784,N_49624);
nor UO_2780 (O_2780,N_49868,N_49697);
xnor UO_2781 (O_2781,N_49650,N_49858);
nand UO_2782 (O_2782,N_49903,N_49625);
and UO_2783 (O_2783,N_49957,N_49895);
xnor UO_2784 (O_2784,N_49533,N_49598);
xor UO_2785 (O_2785,N_49730,N_49521);
nand UO_2786 (O_2786,N_49788,N_49894);
nand UO_2787 (O_2787,N_49816,N_49724);
xor UO_2788 (O_2788,N_49835,N_49610);
and UO_2789 (O_2789,N_49993,N_49929);
or UO_2790 (O_2790,N_49609,N_49569);
xor UO_2791 (O_2791,N_49953,N_49610);
nor UO_2792 (O_2792,N_49673,N_49988);
and UO_2793 (O_2793,N_49637,N_49925);
xor UO_2794 (O_2794,N_49713,N_49757);
or UO_2795 (O_2795,N_49803,N_49917);
and UO_2796 (O_2796,N_49891,N_49651);
xnor UO_2797 (O_2797,N_49895,N_49573);
or UO_2798 (O_2798,N_49953,N_49917);
or UO_2799 (O_2799,N_49925,N_49547);
xnor UO_2800 (O_2800,N_49631,N_49583);
and UO_2801 (O_2801,N_49810,N_49892);
nor UO_2802 (O_2802,N_49661,N_49500);
xor UO_2803 (O_2803,N_49641,N_49913);
nand UO_2804 (O_2804,N_49918,N_49530);
xnor UO_2805 (O_2805,N_49749,N_49759);
or UO_2806 (O_2806,N_49716,N_49755);
xnor UO_2807 (O_2807,N_49609,N_49805);
or UO_2808 (O_2808,N_49570,N_49885);
or UO_2809 (O_2809,N_49706,N_49683);
and UO_2810 (O_2810,N_49752,N_49850);
or UO_2811 (O_2811,N_49803,N_49678);
nor UO_2812 (O_2812,N_49672,N_49606);
nand UO_2813 (O_2813,N_49987,N_49500);
or UO_2814 (O_2814,N_49991,N_49747);
nand UO_2815 (O_2815,N_49581,N_49963);
or UO_2816 (O_2816,N_49889,N_49564);
nor UO_2817 (O_2817,N_49674,N_49569);
nor UO_2818 (O_2818,N_49952,N_49866);
nor UO_2819 (O_2819,N_49590,N_49703);
nor UO_2820 (O_2820,N_49689,N_49649);
nor UO_2821 (O_2821,N_49777,N_49545);
nor UO_2822 (O_2822,N_49926,N_49799);
nand UO_2823 (O_2823,N_49560,N_49988);
and UO_2824 (O_2824,N_49644,N_49856);
and UO_2825 (O_2825,N_49637,N_49983);
and UO_2826 (O_2826,N_49640,N_49810);
nand UO_2827 (O_2827,N_49771,N_49528);
xnor UO_2828 (O_2828,N_49866,N_49962);
nand UO_2829 (O_2829,N_49564,N_49964);
nor UO_2830 (O_2830,N_49956,N_49930);
or UO_2831 (O_2831,N_49909,N_49689);
and UO_2832 (O_2832,N_49725,N_49638);
nand UO_2833 (O_2833,N_49988,N_49886);
xnor UO_2834 (O_2834,N_49875,N_49630);
nor UO_2835 (O_2835,N_49905,N_49671);
nor UO_2836 (O_2836,N_49525,N_49566);
and UO_2837 (O_2837,N_49808,N_49556);
nand UO_2838 (O_2838,N_49902,N_49581);
and UO_2839 (O_2839,N_49609,N_49703);
nand UO_2840 (O_2840,N_49835,N_49506);
nand UO_2841 (O_2841,N_49852,N_49958);
nor UO_2842 (O_2842,N_49650,N_49626);
nand UO_2843 (O_2843,N_49680,N_49846);
and UO_2844 (O_2844,N_49679,N_49673);
nand UO_2845 (O_2845,N_49698,N_49614);
nand UO_2846 (O_2846,N_49719,N_49738);
and UO_2847 (O_2847,N_49788,N_49896);
nand UO_2848 (O_2848,N_49519,N_49681);
nor UO_2849 (O_2849,N_49843,N_49818);
and UO_2850 (O_2850,N_49896,N_49806);
xnor UO_2851 (O_2851,N_49801,N_49850);
xor UO_2852 (O_2852,N_49691,N_49871);
nor UO_2853 (O_2853,N_49983,N_49576);
or UO_2854 (O_2854,N_49998,N_49934);
or UO_2855 (O_2855,N_49622,N_49734);
xor UO_2856 (O_2856,N_49605,N_49674);
and UO_2857 (O_2857,N_49836,N_49589);
and UO_2858 (O_2858,N_49708,N_49692);
nor UO_2859 (O_2859,N_49549,N_49523);
and UO_2860 (O_2860,N_49748,N_49664);
nor UO_2861 (O_2861,N_49970,N_49859);
and UO_2862 (O_2862,N_49777,N_49634);
or UO_2863 (O_2863,N_49502,N_49915);
xor UO_2864 (O_2864,N_49503,N_49882);
nand UO_2865 (O_2865,N_49945,N_49756);
and UO_2866 (O_2866,N_49885,N_49971);
nor UO_2867 (O_2867,N_49678,N_49591);
and UO_2868 (O_2868,N_49551,N_49871);
or UO_2869 (O_2869,N_49964,N_49744);
or UO_2870 (O_2870,N_49671,N_49986);
xnor UO_2871 (O_2871,N_49852,N_49707);
xor UO_2872 (O_2872,N_49666,N_49622);
and UO_2873 (O_2873,N_49620,N_49745);
or UO_2874 (O_2874,N_49533,N_49647);
or UO_2875 (O_2875,N_49519,N_49928);
xnor UO_2876 (O_2876,N_49943,N_49941);
and UO_2877 (O_2877,N_49974,N_49985);
nor UO_2878 (O_2878,N_49586,N_49720);
and UO_2879 (O_2879,N_49635,N_49806);
nor UO_2880 (O_2880,N_49639,N_49887);
nand UO_2881 (O_2881,N_49812,N_49674);
xnor UO_2882 (O_2882,N_49912,N_49524);
nand UO_2883 (O_2883,N_49643,N_49787);
nor UO_2884 (O_2884,N_49834,N_49959);
and UO_2885 (O_2885,N_49923,N_49653);
xnor UO_2886 (O_2886,N_49714,N_49943);
xnor UO_2887 (O_2887,N_49940,N_49600);
or UO_2888 (O_2888,N_49793,N_49709);
nor UO_2889 (O_2889,N_49663,N_49538);
and UO_2890 (O_2890,N_49941,N_49602);
xor UO_2891 (O_2891,N_49510,N_49563);
xor UO_2892 (O_2892,N_49621,N_49625);
or UO_2893 (O_2893,N_49810,N_49751);
and UO_2894 (O_2894,N_49857,N_49648);
and UO_2895 (O_2895,N_49693,N_49533);
xor UO_2896 (O_2896,N_49825,N_49636);
xor UO_2897 (O_2897,N_49647,N_49665);
nand UO_2898 (O_2898,N_49733,N_49540);
nand UO_2899 (O_2899,N_49754,N_49913);
and UO_2900 (O_2900,N_49526,N_49900);
nor UO_2901 (O_2901,N_49514,N_49760);
nor UO_2902 (O_2902,N_49521,N_49653);
nand UO_2903 (O_2903,N_49932,N_49644);
nand UO_2904 (O_2904,N_49650,N_49544);
and UO_2905 (O_2905,N_49504,N_49784);
and UO_2906 (O_2906,N_49825,N_49676);
and UO_2907 (O_2907,N_49506,N_49721);
and UO_2908 (O_2908,N_49556,N_49679);
or UO_2909 (O_2909,N_49952,N_49678);
and UO_2910 (O_2910,N_49829,N_49749);
and UO_2911 (O_2911,N_49673,N_49750);
or UO_2912 (O_2912,N_49675,N_49669);
or UO_2913 (O_2913,N_49774,N_49907);
and UO_2914 (O_2914,N_49578,N_49601);
nor UO_2915 (O_2915,N_49836,N_49862);
and UO_2916 (O_2916,N_49681,N_49943);
or UO_2917 (O_2917,N_49988,N_49692);
or UO_2918 (O_2918,N_49955,N_49578);
and UO_2919 (O_2919,N_49838,N_49952);
or UO_2920 (O_2920,N_49674,N_49997);
xor UO_2921 (O_2921,N_49786,N_49751);
or UO_2922 (O_2922,N_49895,N_49538);
nand UO_2923 (O_2923,N_49668,N_49712);
nor UO_2924 (O_2924,N_49535,N_49639);
and UO_2925 (O_2925,N_49677,N_49922);
or UO_2926 (O_2926,N_49659,N_49938);
or UO_2927 (O_2927,N_49745,N_49710);
and UO_2928 (O_2928,N_49901,N_49667);
and UO_2929 (O_2929,N_49617,N_49535);
nor UO_2930 (O_2930,N_49826,N_49847);
xor UO_2931 (O_2931,N_49883,N_49671);
nor UO_2932 (O_2932,N_49859,N_49783);
or UO_2933 (O_2933,N_49915,N_49931);
or UO_2934 (O_2934,N_49923,N_49951);
nand UO_2935 (O_2935,N_49593,N_49528);
and UO_2936 (O_2936,N_49526,N_49544);
or UO_2937 (O_2937,N_49991,N_49556);
and UO_2938 (O_2938,N_49747,N_49878);
or UO_2939 (O_2939,N_49978,N_49786);
nor UO_2940 (O_2940,N_49921,N_49630);
nor UO_2941 (O_2941,N_49982,N_49810);
nand UO_2942 (O_2942,N_49555,N_49608);
xor UO_2943 (O_2943,N_49810,N_49581);
or UO_2944 (O_2944,N_49831,N_49740);
or UO_2945 (O_2945,N_49661,N_49921);
nand UO_2946 (O_2946,N_49909,N_49849);
or UO_2947 (O_2947,N_49743,N_49525);
xnor UO_2948 (O_2948,N_49582,N_49667);
xor UO_2949 (O_2949,N_49597,N_49778);
nand UO_2950 (O_2950,N_49644,N_49747);
nand UO_2951 (O_2951,N_49820,N_49631);
nor UO_2952 (O_2952,N_49921,N_49793);
nor UO_2953 (O_2953,N_49956,N_49659);
nand UO_2954 (O_2954,N_49884,N_49555);
xor UO_2955 (O_2955,N_49886,N_49579);
nor UO_2956 (O_2956,N_49906,N_49599);
or UO_2957 (O_2957,N_49680,N_49697);
and UO_2958 (O_2958,N_49779,N_49665);
nor UO_2959 (O_2959,N_49984,N_49640);
xnor UO_2960 (O_2960,N_49514,N_49607);
nand UO_2961 (O_2961,N_49897,N_49507);
nor UO_2962 (O_2962,N_49935,N_49936);
nand UO_2963 (O_2963,N_49501,N_49575);
or UO_2964 (O_2964,N_49929,N_49748);
xnor UO_2965 (O_2965,N_49565,N_49912);
nor UO_2966 (O_2966,N_49797,N_49848);
or UO_2967 (O_2967,N_49889,N_49955);
nand UO_2968 (O_2968,N_49764,N_49767);
or UO_2969 (O_2969,N_49894,N_49687);
and UO_2970 (O_2970,N_49669,N_49571);
or UO_2971 (O_2971,N_49866,N_49846);
xor UO_2972 (O_2972,N_49925,N_49974);
xnor UO_2973 (O_2973,N_49583,N_49946);
nor UO_2974 (O_2974,N_49599,N_49724);
nand UO_2975 (O_2975,N_49807,N_49674);
nor UO_2976 (O_2976,N_49560,N_49848);
or UO_2977 (O_2977,N_49616,N_49754);
xor UO_2978 (O_2978,N_49585,N_49984);
xor UO_2979 (O_2979,N_49844,N_49555);
and UO_2980 (O_2980,N_49824,N_49988);
and UO_2981 (O_2981,N_49662,N_49587);
and UO_2982 (O_2982,N_49540,N_49544);
xnor UO_2983 (O_2983,N_49770,N_49890);
xnor UO_2984 (O_2984,N_49718,N_49703);
and UO_2985 (O_2985,N_49890,N_49968);
nor UO_2986 (O_2986,N_49619,N_49998);
nand UO_2987 (O_2987,N_49709,N_49570);
nor UO_2988 (O_2988,N_49703,N_49519);
nand UO_2989 (O_2989,N_49894,N_49771);
or UO_2990 (O_2990,N_49605,N_49860);
and UO_2991 (O_2991,N_49615,N_49713);
xnor UO_2992 (O_2992,N_49830,N_49825);
or UO_2993 (O_2993,N_49970,N_49525);
nor UO_2994 (O_2994,N_49906,N_49777);
and UO_2995 (O_2995,N_49801,N_49737);
and UO_2996 (O_2996,N_49646,N_49873);
or UO_2997 (O_2997,N_49770,N_49660);
xor UO_2998 (O_2998,N_49556,N_49990);
or UO_2999 (O_2999,N_49934,N_49819);
nor UO_3000 (O_3000,N_49681,N_49741);
or UO_3001 (O_3001,N_49573,N_49560);
or UO_3002 (O_3002,N_49708,N_49568);
or UO_3003 (O_3003,N_49581,N_49515);
and UO_3004 (O_3004,N_49820,N_49666);
nor UO_3005 (O_3005,N_49890,N_49661);
or UO_3006 (O_3006,N_49507,N_49887);
nand UO_3007 (O_3007,N_49524,N_49970);
xnor UO_3008 (O_3008,N_49722,N_49807);
nand UO_3009 (O_3009,N_49665,N_49580);
or UO_3010 (O_3010,N_49506,N_49586);
nand UO_3011 (O_3011,N_49998,N_49799);
and UO_3012 (O_3012,N_49839,N_49927);
nand UO_3013 (O_3013,N_49579,N_49502);
nand UO_3014 (O_3014,N_49700,N_49631);
or UO_3015 (O_3015,N_49814,N_49717);
nor UO_3016 (O_3016,N_49899,N_49563);
nor UO_3017 (O_3017,N_49703,N_49559);
nor UO_3018 (O_3018,N_49645,N_49571);
or UO_3019 (O_3019,N_49569,N_49594);
or UO_3020 (O_3020,N_49716,N_49878);
and UO_3021 (O_3021,N_49609,N_49850);
nand UO_3022 (O_3022,N_49563,N_49806);
or UO_3023 (O_3023,N_49887,N_49956);
nand UO_3024 (O_3024,N_49873,N_49638);
and UO_3025 (O_3025,N_49808,N_49692);
nor UO_3026 (O_3026,N_49630,N_49621);
xor UO_3027 (O_3027,N_49629,N_49996);
or UO_3028 (O_3028,N_49555,N_49843);
nand UO_3029 (O_3029,N_49548,N_49518);
or UO_3030 (O_3030,N_49743,N_49747);
nor UO_3031 (O_3031,N_49627,N_49824);
xnor UO_3032 (O_3032,N_49748,N_49651);
and UO_3033 (O_3033,N_49893,N_49600);
nand UO_3034 (O_3034,N_49838,N_49766);
nor UO_3035 (O_3035,N_49678,N_49619);
and UO_3036 (O_3036,N_49926,N_49607);
or UO_3037 (O_3037,N_49770,N_49551);
or UO_3038 (O_3038,N_49816,N_49940);
nand UO_3039 (O_3039,N_49925,N_49866);
nor UO_3040 (O_3040,N_49596,N_49584);
xor UO_3041 (O_3041,N_49971,N_49759);
xor UO_3042 (O_3042,N_49984,N_49950);
nand UO_3043 (O_3043,N_49684,N_49588);
nand UO_3044 (O_3044,N_49900,N_49600);
xnor UO_3045 (O_3045,N_49767,N_49505);
xor UO_3046 (O_3046,N_49775,N_49986);
or UO_3047 (O_3047,N_49632,N_49611);
nand UO_3048 (O_3048,N_49648,N_49717);
xor UO_3049 (O_3049,N_49533,N_49847);
nor UO_3050 (O_3050,N_49879,N_49815);
and UO_3051 (O_3051,N_49883,N_49602);
nor UO_3052 (O_3052,N_49889,N_49707);
nor UO_3053 (O_3053,N_49587,N_49725);
or UO_3054 (O_3054,N_49936,N_49699);
or UO_3055 (O_3055,N_49719,N_49644);
xor UO_3056 (O_3056,N_49578,N_49519);
and UO_3057 (O_3057,N_49664,N_49502);
nor UO_3058 (O_3058,N_49601,N_49686);
nand UO_3059 (O_3059,N_49818,N_49776);
nand UO_3060 (O_3060,N_49542,N_49663);
and UO_3061 (O_3061,N_49957,N_49769);
or UO_3062 (O_3062,N_49565,N_49885);
or UO_3063 (O_3063,N_49592,N_49979);
nand UO_3064 (O_3064,N_49768,N_49557);
and UO_3065 (O_3065,N_49505,N_49584);
or UO_3066 (O_3066,N_49713,N_49747);
xnor UO_3067 (O_3067,N_49588,N_49671);
nand UO_3068 (O_3068,N_49770,N_49701);
nand UO_3069 (O_3069,N_49556,N_49588);
and UO_3070 (O_3070,N_49879,N_49830);
or UO_3071 (O_3071,N_49878,N_49977);
nand UO_3072 (O_3072,N_49621,N_49657);
and UO_3073 (O_3073,N_49929,N_49612);
nand UO_3074 (O_3074,N_49591,N_49737);
or UO_3075 (O_3075,N_49825,N_49503);
nand UO_3076 (O_3076,N_49786,N_49930);
xor UO_3077 (O_3077,N_49522,N_49653);
or UO_3078 (O_3078,N_49525,N_49567);
or UO_3079 (O_3079,N_49630,N_49986);
or UO_3080 (O_3080,N_49938,N_49645);
or UO_3081 (O_3081,N_49993,N_49636);
xor UO_3082 (O_3082,N_49908,N_49802);
nand UO_3083 (O_3083,N_49955,N_49755);
or UO_3084 (O_3084,N_49654,N_49503);
and UO_3085 (O_3085,N_49966,N_49844);
nor UO_3086 (O_3086,N_49907,N_49701);
and UO_3087 (O_3087,N_49983,N_49929);
or UO_3088 (O_3088,N_49955,N_49834);
nor UO_3089 (O_3089,N_49911,N_49716);
and UO_3090 (O_3090,N_49931,N_49734);
and UO_3091 (O_3091,N_49786,N_49506);
or UO_3092 (O_3092,N_49572,N_49969);
nand UO_3093 (O_3093,N_49760,N_49697);
nor UO_3094 (O_3094,N_49560,N_49703);
xor UO_3095 (O_3095,N_49666,N_49813);
nor UO_3096 (O_3096,N_49697,N_49960);
xor UO_3097 (O_3097,N_49839,N_49822);
nor UO_3098 (O_3098,N_49512,N_49807);
nor UO_3099 (O_3099,N_49681,N_49510);
or UO_3100 (O_3100,N_49832,N_49949);
nor UO_3101 (O_3101,N_49937,N_49955);
nand UO_3102 (O_3102,N_49534,N_49713);
or UO_3103 (O_3103,N_49903,N_49829);
and UO_3104 (O_3104,N_49710,N_49645);
nand UO_3105 (O_3105,N_49639,N_49719);
and UO_3106 (O_3106,N_49544,N_49808);
nor UO_3107 (O_3107,N_49625,N_49939);
nor UO_3108 (O_3108,N_49515,N_49628);
nor UO_3109 (O_3109,N_49864,N_49563);
or UO_3110 (O_3110,N_49774,N_49623);
xor UO_3111 (O_3111,N_49654,N_49764);
and UO_3112 (O_3112,N_49632,N_49970);
xnor UO_3113 (O_3113,N_49818,N_49528);
and UO_3114 (O_3114,N_49868,N_49671);
nor UO_3115 (O_3115,N_49755,N_49704);
and UO_3116 (O_3116,N_49952,N_49886);
xor UO_3117 (O_3117,N_49744,N_49724);
nand UO_3118 (O_3118,N_49536,N_49748);
nand UO_3119 (O_3119,N_49910,N_49656);
nor UO_3120 (O_3120,N_49927,N_49773);
nand UO_3121 (O_3121,N_49920,N_49993);
or UO_3122 (O_3122,N_49759,N_49979);
nand UO_3123 (O_3123,N_49808,N_49500);
or UO_3124 (O_3124,N_49997,N_49662);
nand UO_3125 (O_3125,N_49873,N_49609);
and UO_3126 (O_3126,N_49685,N_49670);
nand UO_3127 (O_3127,N_49586,N_49714);
or UO_3128 (O_3128,N_49539,N_49583);
nand UO_3129 (O_3129,N_49638,N_49635);
nand UO_3130 (O_3130,N_49748,N_49890);
nor UO_3131 (O_3131,N_49602,N_49571);
and UO_3132 (O_3132,N_49861,N_49804);
or UO_3133 (O_3133,N_49825,N_49651);
and UO_3134 (O_3134,N_49875,N_49825);
nor UO_3135 (O_3135,N_49880,N_49712);
xnor UO_3136 (O_3136,N_49589,N_49746);
nor UO_3137 (O_3137,N_49905,N_49910);
and UO_3138 (O_3138,N_49666,N_49806);
or UO_3139 (O_3139,N_49506,N_49745);
and UO_3140 (O_3140,N_49605,N_49978);
and UO_3141 (O_3141,N_49619,N_49739);
xor UO_3142 (O_3142,N_49725,N_49623);
and UO_3143 (O_3143,N_49568,N_49610);
xor UO_3144 (O_3144,N_49886,N_49677);
nor UO_3145 (O_3145,N_49986,N_49767);
nand UO_3146 (O_3146,N_49860,N_49723);
nand UO_3147 (O_3147,N_49846,N_49966);
nand UO_3148 (O_3148,N_49648,N_49632);
nor UO_3149 (O_3149,N_49988,N_49785);
or UO_3150 (O_3150,N_49737,N_49725);
nand UO_3151 (O_3151,N_49769,N_49873);
nor UO_3152 (O_3152,N_49859,N_49882);
nand UO_3153 (O_3153,N_49620,N_49573);
or UO_3154 (O_3154,N_49691,N_49660);
nand UO_3155 (O_3155,N_49524,N_49504);
xor UO_3156 (O_3156,N_49797,N_49894);
or UO_3157 (O_3157,N_49850,N_49998);
xor UO_3158 (O_3158,N_49858,N_49527);
nand UO_3159 (O_3159,N_49882,N_49998);
and UO_3160 (O_3160,N_49629,N_49569);
and UO_3161 (O_3161,N_49674,N_49713);
nand UO_3162 (O_3162,N_49737,N_49877);
or UO_3163 (O_3163,N_49690,N_49669);
and UO_3164 (O_3164,N_49581,N_49503);
or UO_3165 (O_3165,N_49548,N_49967);
or UO_3166 (O_3166,N_49518,N_49867);
or UO_3167 (O_3167,N_49775,N_49668);
or UO_3168 (O_3168,N_49659,N_49983);
or UO_3169 (O_3169,N_49709,N_49888);
and UO_3170 (O_3170,N_49804,N_49904);
or UO_3171 (O_3171,N_49884,N_49767);
or UO_3172 (O_3172,N_49895,N_49745);
or UO_3173 (O_3173,N_49703,N_49721);
or UO_3174 (O_3174,N_49576,N_49977);
nor UO_3175 (O_3175,N_49851,N_49907);
or UO_3176 (O_3176,N_49914,N_49969);
xnor UO_3177 (O_3177,N_49545,N_49680);
nand UO_3178 (O_3178,N_49619,N_49682);
or UO_3179 (O_3179,N_49826,N_49621);
and UO_3180 (O_3180,N_49624,N_49529);
and UO_3181 (O_3181,N_49855,N_49913);
xor UO_3182 (O_3182,N_49833,N_49686);
or UO_3183 (O_3183,N_49568,N_49925);
or UO_3184 (O_3184,N_49970,N_49846);
xnor UO_3185 (O_3185,N_49749,N_49675);
nand UO_3186 (O_3186,N_49796,N_49740);
xor UO_3187 (O_3187,N_49961,N_49777);
or UO_3188 (O_3188,N_49998,N_49553);
nor UO_3189 (O_3189,N_49693,N_49990);
nor UO_3190 (O_3190,N_49895,N_49860);
and UO_3191 (O_3191,N_49667,N_49820);
and UO_3192 (O_3192,N_49922,N_49845);
and UO_3193 (O_3193,N_49622,N_49878);
xor UO_3194 (O_3194,N_49563,N_49569);
or UO_3195 (O_3195,N_49692,N_49985);
nand UO_3196 (O_3196,N_49904,N_49860);
and UO_3197 (O_3197,N_49585,N_49542);
and UO_3198 (O_3198,N_49688,N_49789);
and UO_3199 (O_3199,N_49767,N_49804);
or UO_3200 (O_3200,N_49739,N_49574);
nor UO_3201 (O_3201,N_49987,N_49648);
and UO_3202 (O_3202,N_49543,N_49661);
or UO_3203 (O_3203,N_49840,N_49779);
or UO_3204 (O_3204,N_49531,N_49872);
and UO_3205 (O_3205,N_49854,N_49534);
nand UO_3206 (O_3206,N_49579,N_49626);
or UO_3207 (O_3207,N_49619,N_49637);
nand UO_3208 (O_3208,N_49518,N_49990);
nand UO_3209 (O_3209,N_49760,N_49879);
nor UO_3210 (O_3210,N_49940,N_49988);
and UO_3211 (O_3211,N_49513,N_49682);
nor UO_3212 (O_3212,N_49758,N_49748);
nand UO_3213 (O_3213,N_49544,N_49679);
xor UO_3214 (O_3214,N_49984,N_49850);
nor UO_3215 (O_3215,N_49838,N_49504);
xor UO_3216 (O_3216,N_49613,N_49843);
nor UO_3217 (O_3217,N_49670,N_49641);
or UO_3218 (O_3218,N_49906,N_49543);
nor UO_3219 (O_3219,N_49956,N_49613);
and UO_3220 (O_3220,N_49876,N_49955);
nand UO_3221 (O_3221,N_49949,N_49756);
and UO_3222 (O_3222,N_49717,N_49722);
and UO_3223 (O_3223,N_49952,N_49935);
or UO_3224 (O_3224,N_49599,N_49580);
xnor UO_3225 (O_3225,N_49900,N_49850);
xnor UO_3226 (O_3226,N_49565,N_49643);
and UO_3227 (O_3227,N_49533,N_49741);
or UO_3228 (O_3228,N_49909,N_49872);
nor UO_3229 (O_3229,N_49952,N_49588);
and UO_3230 (O_3230,N_49597,N_49988);
and UO_3231 (O_3231,N_49713,N_49904);
nand UO_3232 (O_3232,N_49869,N_49953);
nand UO_3233 (O_3233,N_49766,N_49502);
xor UO_3234 (O_3234,N_49809,N_49846);
or UO_3235 (O_3235,N_49648,N_49769);
xor UO_3236 (O_3236,N_49563,N_49711);
nand UO_3237 (O_3237,N_49893,N_49730);
and UO_3238 (O_3238,N_49655,N_49565);
nor UO_3239 (O_3239,N_49934,N_49989);
xnor UO_3240 (O_3240,N_49889,N_49970);
xor UO_3241 (O_3241,N_49874,N_49510);
nand UO_3242 (O_3242,N_49989,N_49732);
and UO_3243 (O_3243,N_49815,N_49668);
nor UO_3244 (O_3244,N_49706,N_49666);
nand UO_3245 (O_3245,N_49855,N_49669);
or UO_3246 (O_3246,N_49741,N_49736);
or UO_3247 (O_3247,N_49993,N_49696);
nand UO_3248 (O_3248,N_49946,N_49830);
nor UO_3249 (O_3249,N_49736,N_49991);
or UO_3250 (O_3250,N_49976,N_49610);
nand UO_3251 (O_3251,N_49785,N_49712);
xnor UO_3252 (O_3252,N_49536,N_49844);
nand UO_3253 (O_3253,N_49641,N_49935);
nand UO_3254 (O_3254,N_49996,N_49592);
and UO_3255 (O_3255,N_49505,N_49724);
xor UO_3256 (O_3256,N_49928,N_49603);
nor UO_3257 (O_3257,N_49767,N_49668);
xor UO_3258 (O_3258,N_49923,N_49645);
xor UO_3259 (O_3259,N_49526,N_49972);
or UO_3260 (O_3260,N_49799,N_49561);
nand UO_3261 (O_3261,N_49772,N_49662);
and UO_3262 (O_3262,N_49769,N_49927);
and UO_3263 (O_3263,N_49649,N_49808);
or UO_3264 (O_3264,N_49990,N_49745);
nand UO_3265 (O_3265,N_49602,N_49619);
nand UO_3266 (O_3266,N_49847,N_49883);
xnor UO_3267 (O_3267,N_49659,N_49895);
nor UO_3268 (O_3268,N_49710,N_49542);
or UO_3269 (O_3269,N_49557,N_49834);
xnor UO_3270 (O_3270,N_49897,N_49545);
nor UO_3271 (O_3271,N_49630,N_49878);
nand UO_3272 (O_3272,N_49992,N_49848);
nand UO_3273 (O_3273,N_49808,N_49602);
nor UO_3274 (O_3274,N_49611,N_49749);
nand UO_3275 (O_3275,N_49904,N_49835);
nor UO_3276 (O_3276,N_49778,N_49567);
and UO_3277 (O_3277,N_49634,N_49733);
xnor UO_3278 (O_3278,N_49583,N_49741);
and UO_3279 (O_3279,N_49522,N_49578);
xor UO_3280 (O_3280,N_49531,N_49537);
nand UO_3281 (O_3281,N_49583,N_49552);
and UO_3282 (O_3282,N_49980,N_49680);
nor UO_3283 (O_3283,N_49546,N_49699);
nand UO_3284 (O_3284,N_49557,N_49942);
nand UO_3285 (O_3285,N_49658,N_49679);
xor UO_3286 (O_3286,N_49844,N_49544);
nor UO_3287 (O_3287,N_49714,N_49593);
and UO_3288 (O_3288,N_49630,N_49723);
or UO_3289 (O_3289,N_49828,N_49902);
nand UO_3290 (O_3290,N_49876,N_49556);
and UO_3291 (O_3291,N_49999,N_49674);
nand UO_3292 (O_3292,N_49871,N_49566);
xor UO_3293 (O_3293,N_49908,N_49910);
nand UO_3294 (O_3294,N_49552,N_49830);
nor UO_3295 (O_3295,N_49868,N_49800);
xor UO_3296 (O_3296,N_49836,N_49617);
xnor UO_3297 (O_3297,N_49637,N_49843);
nor UO_3298 (O_3298,N_49898,N_49720);
and UO_3299 (O_3299,N_49684,N_49646);
or UO_3300 (O_3300,N_49628,N_49918);
xor UO_3301 (O_3301,N_49908,N_49542);
nand UO_3302 (O_3302,N_49903,N_49556);
xor UO_3303 (O_3303,N_49893,N_49777);
nor UO_3304 (O_3304,N_49760,N_49901);
xor UO_3305 (O_3305,N_49579,N_49569);
or UO_3306 (O_3306,N_49544,N_49785);
nand UO_3307 (O_3307,N_49821,N_49772);
xor UO_3308 (O_3308,N_49595,N_49839);
xnor UO_3309 (O_3309,N_49902,N_49735);
nor UO_3310 (O_3310,N_49974,N_49954);
or UO_3311 (O_3311,N_49817,N_49799);
nor UO_3312 (O_3312,N_49814,N_49673);
and UO_3313 (O_3313,N_49635,N_49634);
or UO_3314 (O_3314,N_49995,N_49682);
and UO_3315 (O_3315,N_49614,N_49760);
nand UO_3316 (O_3316,N_49811,N_49891);
xnor UO_3317 (O_3317,N_49761,N_49613);
xnor UO_3318 (O_3318,N_49584,N_49547);
and UO_3319 (O_3319,N_49616,N_49783);
xor UO_3320 (O_3320,N_49690,N_49753);
xnor UO_3321 (O_3321,N_49717,N_49732);
or UO_3322 (O_3322,N_49564,N_49852);
nor UO_3323 (O_3323,N_49520,N_49711);
nor UO_3324 (O_3324,N_49625,N_49520);
and UO_3325 (O_3325,N_49760,N_49847);
and UO_3326 (O_3326,N_49997,N_49568);
nor UO_3327 (O_3327,N_49929,N_49713);
xor UO_3328 (O_3328,N_49849,N_49716);
xor UO_3329 (O_3329,N_49777,N_49820);
nand UO_3330 (O_3330,N_49912,N_49849);
nor UO_3331 (O_3331,N_49878,N_49954);
nand UO_3332 (O_3332,N_49651,N_49859);
or UO_3333 (O_3333,N_49673,N_49815);
xnor UO_3334 (O_3334,N_49732,N_49516);
nor UO_3335 (O_3335,N_49507,N_49869);
or UO_3336 (O_3336,N_49691,N_49726);
or UO_3337 (O_3337,N_49784,N_49902);
and UO_3338 (O_3338,N_49648,N_49977);
nor UO_3339 (O_3339,N_49507,N_49936);
or UO_3340 (O_3340,N_49577,N_49606);
or UO_3341 (O_3341,N_49934,N_49824);
or UO_3342 (O_3342,N_49830,N_49849);
nand UO_3343 (O_3343,N_49824,N_49714);
nor UO_3344 (O_3344,N_49678,N_49531);
xnor UO_3345 (O_3345,N_49858,N_49794);
and UO_3346 (O_3346,N_49723,N_49643);
xnor UO_3347 (O_3347,N_49585,N_49742);
and UO_3348 (O_3348,N_49870,N_49767);
and UO_3349 (O_3349,N_49755,N_49781);
or UO_3350 (O_3350,N_49537,N_49881);
xnor UO_3351 (O_3351,N_49683,N_49648);
nand UO_3352 (O_3352,N_49646,N_49612);
xor UO_3353 (O_3353,N_49951,N_49986);
and UO_3354 (O_3354,N_49846,N_49644);
or UO_3355 (O_3355,N_49886,N_49702);
nand UO_3356 (O_3356,N_49699,N_49943);
xnor UO_3357 (O_3357,N_49576,N_49506);
xnor UO_3358 (O_3358,N_49584,N_49603);
nor UO_3359 (O_3359,N_49773,N_49995);
xnor UO_3360 (O_3360,N_49552,N_49739);
nand UO_3361 (O_3361,N_49664,N_49998);
or UO_3362 (O_3362,N_49556,N_49693);
or UO_3363 (O_3363,N_49657,N_49912);
or UO_3364 (O_3364,N_49745,N_49817);
and UO_3365 (O_3365,N_49736,N_49607);
nand UO_3366 (O_3366,N_49945,N_49525);
xnor UO_3367 (O_3367,N_49849,N_49856);
or UO_3368 (O_3368,N_49742,N_49631);
or UO_3369 (O_3369,N_49514,N_49649);
or UO_3370 (O_3370,N_49525,N_49985);
or UO_3371 (O_3371,N_49991,N_49685);
and UO_3372 (O_3372,N_49552,N_49538);
and UO_3373 (O_3373,N_49505,N_49893);
nor UO_3374 (O_3374,N_49896,N_49576);
xnor UO_3375 (O_3375,N_49872,N_49586);
nand UO_3376 (O_3376,N_49894,N_49569);
nand UO_3377 (O_3377,N_49677,N_49635);
xnor UO_3378 (O_3378,N_49948,N_49714);
or UO_3379 (O_3379,N_49963,N_49756);
nand UO_3380 (O_3380,N_49662,N_49677);
nand UO_3381 (O_3381,N_49677,N_49875);
xor UO_3382 (O_3382,N_49866,N_49976);
nand UO_3383 (O_3383,N_49669,N_49826);
nor UO_3384 (O_3384,N_49634,N_49993);
and UO_3385 (O_3385,N_49777,N_49506);
nand UO_3386 (O_3386,N_49740,N_49836);
nor UO_3387 (O_3387,N_49897,N_49826);
xor UO_3388 (O_3388,N_49771,N_49567);
or UO_3389 (O_3389,N_49946,N_49923);
or UO_3390 (O_3390,N_49766,N_49721);
and UO_3391 (O_3391,N_49503,N_49776);
or UO_3392 (O_3392,N_49567,N_49984);
and UO_3393 (O_3393,N_49842,N_49588);
and UO_3394 (O_3394,N_49973,N_49844);
and UO_3395 (O_3395,N_49785,N_49673);
xor UO_3396 (O_3396,N_49604,N_49861);
nor UO_3397 (O_3397,N_49763,N_49945);
nor UO_3398 (O_3398,N_49878,N_49797);
nand UO_3399 (O_3399,N_49603,N_49855);
xnor UO_3400 (O_3400,N_49607,N_49808);
nor UO_3401 (O_3401,N_49921,N_49857);
or UO_3402 (O_3402,N_49589,N_49608);
nor UO_3403 (O_3403,N_49585,N_49767);
and UO_3404 (O_3404,N_49529,N_49891);
nor UO_3405 (O_3405,N_49612,N_49556);
xnor UO_3406 (O_3406,N_49640,N_49969);
xor UO_3407 (O_3407,N_49998,N_49667);
nand UO_3408 (O_3408,N_49615,N_49725);
xor UO_3409 (O_3409,N_49520,N_49903);
xor UO_3410 (O_3410,N_49883,N_49659);
nor UO_3411 (O_3411,N_49500,N_49830);
and UO_3412 (O_3412,N_49978,N_49715);
nor UO_3413 (O_3413,N_49825,N_49749);
and UO_3414 (O_3414,N_49839,N_49835);
nor UO_3415 (O_3415,N_49674,N_49595);
nor UO_3416 (O_3416,N_49845,N_49623);
nor UO_3417 (O_3417,N_49626,N_49890);
xor UO_3418 (O_3418,N_49775,N_49619);
nor UO_3419 (O_3419,N_49753,N_49641);
nor UO_3420 (O_3420,N_49791,N_49777);
nand UO_3421 (O_3421,N_49843,N_49992);
and UO_3422 (O_3422,N_49762,N_49534);
and UO_3423 (O_3423,N_49578,N_49810);
and UO_3424 (O_3424,N_49740,N_49596);
nand UO_3425 (O_3425,N_49653,N_49574);
xor UO_3426 (O_3426,N_49843,N_49977);
xnor UO_3427 (O_3427,N_49862,N_49826);
and UO_3428 (O_3428,N_49629,N_49653);
xor UO_3429 (O_3429,N_49568,N_49683);
and UO_3430 (O_3430,N_49983,N_49590);
nand UO_3431 (O_3431,N_49714,N_49920);
or UO_3432 (O_3432,N_49628,N_49946);
and UO_3433 (O_3433,N_49886,N_49878);
or UO_3434 (O_3434,N_49501,N_49622);
nor UO_3435 (O_3435,N_49625,N_49746);
and UO_3436 (O_3436,N_49763,N_49943);
and UO_3437 (O_3437,N_49786,N_49806);
nor UO_3438 (O_3438,N_49729,N_49719);
xor UO_3439 (O_3439,N_49769,N_49976);
xnor UO_3440 (O_3440,N_49909,N_49659);
nand UO_3441 (O_3441,N_49823,N_49557);
nand UO_3442 (O_3442,N_49527,N_49950);
or UO_3443 (O_3443,N_49522,N_49958);
xnor UO_3444 (O_3444,N_49541,N_49893);
nand UO_3445 (O_3445,N_49779,N_49674);
nor UO_3446 (O_3446,N_49826,N_49591);
or UO_3447 (O_3447,N_49949,N_49794);
or UO_3448 (O_3448,N_49834,N_49810);
nand UO_3449 (O_3449,N_49665,N_49786);
nand UO_3450 (O_3450,N_49874,N_49513);
xnor UO_3451 (O_3451,N_49978,N_49520);
nand UO_3452 (O_3452,N_49502,N_49955);
nor UO_3453 (O_3453,N_49584,N_49665);
nand UO_3454 (O_3454,N_49582,N_49989);
and UO_3455 (O_3455,N_49835,N_49808);
or UO_3456 (O_3456,N_49612,N_49995);
or UO_3457 (O_3457,N_49966,N_49768);
nand UO_3458 (O_3458,N_49677,N_49910);
and UO_3459 (O_3459,N_49856,N_49994);
xor UO_3460 (O_3460,N_49691,N_49555);
or UO_3461 (O_3461,N_49625,N_49614);
or UO_3462 (O_3462,N_49585,N_49512);
or UO_3463 (O_3463,N_49881,N_49651);
or UO_3464 (O_3464,N_49995,N_49635);
nand UO_3465 (O_3465,N_49884,N_49859);
nand UO_3466 (O_3466,N_49677,N_49986);
nor UO_3467 (O_3467,N_49691,N_49803);
and UO_3468 (O_3468,N_49857,N_49799);
xor UO_3469 (O_3469,N_49696,N_49905);
xnor UO_3470 (O_3470,N_49942,N_49998);
nor UO_3471 (O_3471,N_49945,N_49745);
xnor UO_3472 (O_3472,N_49933,N_49751);
or UO_3473 (O_3473,N_49702,N_49780);
or UO_3474 (O_3474,N_49615,N_49631);
nor UO_3475 (O_3475,N_49872,N_49802);
nand UO_3476 (O_3476,N_49551,N_49560);
nor UO_3477 (O_3477,N_49870,N_49622);
nand UO_3478 (O_3478,N_49904,N_49572);
xor UO_3479 (O_3479,N_49883,N_49675);
nor UO_3480 (O_3480,N_49932,N_49640);
nand UO_3481 (O_3481,N_49548,N_49758);
nand UO_3482 (O_3482,N_49997,N_49525);
xor UO_3483 (O_3483,N_49560,N_49529);
or UO_3484 (O_3484,N_49600,N_49756);
nand UO_3485 (O_3485,N_49574,N_49799);
nor UO_3486 (O_3486,N_49729,N_49816);
xor UO_3487 (O_3487,N_49952,N_49951);
xor UO_3488 (O_3488,N_49759,N_49589);
xnor UO_3489 (O_3489,N_49849,N_49772);
nand UO_3490 (O_3490,N_49895,N_49726);
or UO_3491 (O_3491,N_49611,N_49563);
nor UO_3492 (O_3492,N_49778,N_49689);
xor UO_3493 (O_3493,N_49683,N_49541);
nand UO_3494 (O_3494,N_49596,N_49760);
xnor UO_3495 (O_3495,N_49513,N_49980);
nor UO_3496 (O_3496,N_49830,N_49934);
or UO_3497 (O_3497,N_49524,N_49592);
or UO_3498 (O_3498,N_49922,N_49812);
nand UO_3499 (O_3499,N_49738,N_49623);
xor UO_3500 (O_3500,N_49893,N_49503);
nor UO_3501 (O_3501,N_49534,N_49944);
or UO_3502 (O_3502,N_49537,N_49696);
xnor UO_3503 (O_3503,N_49727,N_49662);
or UO_3504 (O_3504,N_49635,N_49607);
or UO_3505 (O_3505,N_49844,N_49712);
nor UO_3506 (O_3506,N_49900,N_49774);
nand UO_3507 (O_3507,N_49755,N_49649);
or UO_3508 (O_3508,N_49751,N_49747);
or UO_3509 (O_3509,N_49673,N_49939);
xnor UO_3510 (O_3510,N_49852,N_49822);
and UO_3511 (O_3511,N_49733,N_49710);
and UO_3512 (O_3512,N_49533,N_49559);
nand UO_3513 (O_3513,N_49805,N_49514);
xor UO_3514 (O_3514,N_49690,N_49800);
or UO_3515 (O_3515,N_49549,N_49900);
and UO_3516 (O_3516,N_49821,N_49919);
and UO_3517 (O_3517,N_49928,N_49579);
nand UO_3518 (O_3518,N_49573,N_49948);
or UO_3519 (O_3519,N_49757,N_49562);
xnor UO_3520 (O_3520,N_49723,N_49844);
xnor UO_3521 (O_3521,N_49767,N_49867);
or UO_3522 (O_3522,N_49956,N_49534);
nor UO_3523 (O_3523,N_49649,N_49827);
nand UO_3524 (O_3524,N_49534,N_49828);
nor UO_3525 (O_3525,N_49819,N_49948);
nor UO_3526 (O_3526,N_49749,N_49950);
and UO_3527 (O_3527,N_49733,N_49653);
and UO_3528 (O_3528,N_49869,N_49780);
and UO_3529 (O_3529,N_49950,N_49582);
and UO_3530 (O_3530,N_49567,N_49715);
nand UO_3531 (O_3531,N_49975,N_49544);
nor UO_3532 (O_3532,N_49754,N_49542);
or UO_3533 (O_3533,N_49622,N_49709);
xor UO_3534 (O_3534,N_49837,N_49756);
and UO_3535 (O_3535,N_49911,N_49810);
or UO_3536 (O_3536,N_49896,N_49675);
xor UO_3537 (O_3537,N_49740,N_49588);
or UO_3538 (O_3538,N_49694,N_49942);
nand UO_3539 (O_3539,N_49631,N_49977);
nor UO_3540 (O_3540,N_49823,N_49944);
xnor UO_3541 (O_3541,N_49744,N_49676);
nand UO_3542 (O_3542,N_49872,N_49916);
xor UO_3543 (O_3543,N_49599,N_49856);
or UO_3544 (O_3544,N_49733,N_49848);
nor UO_3545 (O_3545,N_49889,N_49590);
xnor UO_3546 (O_3546,N_49642,N_49931);
or UO_3547 (O_3547,N_49971,N_49892);
and UO_3548 (O_3548,N_49615,N_49920);
and UO_3549 (O_3549,N_49561,N_49994);
nor UO_3550 (O_3550,N_49586,N_49608);
or UO_3551 (O_3551,N_49991,N_49585);
or UO_3552 (O_3552,N_49705,N_49726);
nand UO_3553 (O_3553,N_49741,N_49814);
or UO_3554 (O_3554,N_49547,N_49641);
nand UO_3555 (O_3555,N_49583,N_49646);
and UO_3556 (O_3556,N_49896,N_49746);
and UO_3557 (O_3557,N_49623,N_49735);
and UO_3558 (O_3558,N_49616,N_49583);
xnor UO_3559 (O_3559,N_49538,N_49965);
nor UO_3560 (O_3560,N_49637,N_49914);
or UO_3561 (O_3561,N_49718,N_49915);
or UO_3562 (O_3562,N_49868,N_49797);
nand UO_3563 (O_3563,N_49887,N_49898);
xor UO_3564 (O_3564,N_49976,N_49775);
nand UO_3565 (O_3565,N_49621,N_49669);
xnor UO_3566 (O_3566,N_49847,N_49723);
or UO_3567 (O_3567,N_49651,N_49909);
and UO_3568 (O_3568,N_49687,N_49988);
or UO_3569 (O_3569,N_49908,N_49561);
nor UO_3570 (O_3570,N_49520,N_49723);
and UO_3571 (O_3571,N_49990,N_49641);
nand UO_3572 (O_3572,N_49885,N_49947);
or UO_3573 (O_3573,N_49892,N_49630);
nor UO_3574 (O_3574,N_49532,N_49526);
and UO_3575 (O_3575,N_49871,N_49715);
and UO_3576 (O_3576,N_49542,N_49761);
xor UO_3577 (O_3577,N_49721,N_49529);
and UO_3578 (O_3578,N_49901,N_49832);
and UO_3579 (O_3579,N_49977,N_49530);
and UO_3580 (O_3580,N_49509,N_49950);
and UO_3581 (O_3581,N_49523,N_49684);
and UO_3582 (O_3582,N_49785,N_49553);
nand UO_3583 (O_3583,N_49993,N_49954);
nand UO_3584 (O_3584,N_49523,N_49991);
nand UO_3585 (O_3585,N_49947,N_49942);
and UO_3586 (O_3586,N_49743,N_49723);
nor UO_3587 (O_3587,N_49523,N_49982);
nand UO_3588 (O_3588,N_49684,N_49692);
nor UO_3589 (O_3589,N_49663,N_49760);
nand UO_3590 (O_3590,N_49817,N_49874);
or UO_3591 (O_3591,N_49747,N_49974);
nor UO_3592 (O_3592,N_49934,N_49736);
and UO_3593 (O_3593,N_49982,N_49723);
and UO_3594 (O_3594,N_49946,N_49562);
or UO_3595 (O_3595,N_49731,N_49987);
nand UO_3596 (O_3596,N_49722,N_49779);
nor UO_3597 (O_3597,N_49784,N_49766);
and UO_3598 (O_3598,N_49555,N_49930);
nand UO_3599 (O_3599,N_49885,N_49672);
nand UO_3600 (O_3600,N_49756,N_49784);
and UO_3601 (O_3601,N_49676,N_49567);
or UO_3602 (O_3602,N_49862,N_49850);
nand UO_3603 (O_3603,N_49743,N_49675);
or UO_3604 (O_3604,N_49854,N_49795);
nand UO_3605 (O_3605,N_49935,N_49917);
xnor UO_3606 (O_3606,N_49921,N_49844);
xnor UO_3607 (O_3607,N_49656,N_49935);
and UO_3608 (O_3608,N_49948,N_49709);
and UO_3609 (O_3609,N_49816,N_49735);
xor UO_3610 (O_3610,N_49596,N_49914);
nand UO_3611 (O_3611,N_49604,N_49714);
and UO_3612 (O_3612,N_49815,N_49655);
xor UO_3613 (O_3613,N_49649,N_49941);
or UO_3614 (O_3614,N_49885,N_49634);
xor UO_3615 (O_3615,N_49979,N_49610);
nand UO_3616 (O_3616,N_49762,N_49660);
xor UO_3617 (O_3617,N_49845,N_49512);
nor UO_3618 (O_3618,N_49947,N_49812);
nor UO_3619 (O_3619,N_49799,N_49551);
nand UO_3620 (O_3620,N_49661,N_49567);
or UO_3621 (O_3621,N_49756,N_49936);
or UO_3622 (O_3622,N_49669,N_49917);
and UO_3623 (O_3623,N_49567,N_49609);
xnor UO_3624 (O_3624,N_49671,N_49789);
or UO_3625 (O_3625,N_49874,N_49738);
nand UO_3626 (O_3626,N_49732,N_49931);
nand UO_3627 (O_3627,N_49844,N_49563);
xnor UO_3628 (O_3628,N_49867,N_49802);
or UO_3629 (O_3629,N_49960,N_49546);
nand UO_3630 (O_3630,N_49677,N_49715);
xnor UO_3631 (O_3631,N_49531,N_49923);
or UO_3632 (O_3632,N_49900,N_49798);
nand UO_3633 (O_3633,N_49852,N_49823);
and UO_3634 (O_3634,N_49997,N_49847);
or UO_3635 (O_3635,N_49614,N_49694);
nor UO_3636 (O_3636,N_49982,N_49729);
nor UO_3637 (O_3637,N_49952,N_49732);
nor UO_3638 (O_3638,N_49792,N_49983);
and UO_3639 (O_3639,N_49793,N_49639);
nor UO_3640 (O_3640,N_49992,N_49756);
or UO_3641 (O_3641,N_49834,N_49751);
nor UO_3642 (O_3642,N_49821,N_49845);
xnor UO_3643 (O_3643,N_49738,N_49568);
xnor UO_3644 (O_3644,N_49972,N_49568);
xor UO_3645 (O_3645,N_49748,N_49606);
nand UO_3646 (O_3646,N_49812,N_49566);
or UO_3647 (O_3647,N_49682,N_49501);
and UO_3648 (O_3648,N_49670,N_49583);
and UO_3649 (O_3649,N_49966,N_49605);
nor UO_3650 (O_3650,N_49686,N_49776);
nand UO_3651 (O_3651,N_49804,N_49703);
nor UO_3652 (O_3652,N_49583,N_49627);
and UO_3653 (O_3653,N_49513,N_49508);
or UO_3654 (O_3654,N_49967,N_49612);
and UO_3655 (O_3655,N_49752,N_49937);
and UO_3656 (O_3656,N_49921,N_49700);
nor UO_3657 (O_3657,N_49981,N_49936);
and UO_3658 (O_3658,N_49541,N_49775);
and UO_3659 (O_3659,N_49957,N_49828);
xor UO_3660 (O_3660,N_49682,N_49971);
or UO_3661 (O_3661,N_49849,N_49983);
or UO_3662 (O_3662,N_49701,N_49562);
xnor UO_3663 (O_3663,N_49502,N_49632);
nor UO_3664 (O_3664,N_49758,N_49842);
nor UO_3665 (O_3665,N_49781,N_49546);
xnor UO_3666 (O_3666,N_49746,N_49944);
xnor UO_3667 (O_3667,N_49512,N_49720);
xnor UO_3668 (O_3668,N_49514,N_49822);
or UO_3669 (O_3669,N_49550,N_49883);
and UO_3670 (O_3670,N_49697,N_49990);
and UO_3671 (O_3671,N_49712,N_49968);
nand UO_3672 (O_3672,N_49725,N_49851);
xnor UO_3673 (O_3673,N_49605,N_49619);
or UO_3674 (O_3674,N_49502,N_49880);
nand UO_3675 (O_3675,N_49959,N_49660);
xor UO_3676 (O_3676,N_49613,N_49573);
xor UO_3677 (O_3677,N_49525,N_49516);
or UO_3678 (O_3678,N_49885,N_49553);
and UO_3679 (O_3679,N_49577,N_49573);
or UO_3680 (O_3680,N_49813,N_49567);
nor UO_3681 (O_3681,N_49504,N_49709);
and UO_3682 (O_3682,N_49813,N_49891);
nor UO_3683 (O_3683,N_49795,N_49837);
nor UO_3684 (O_3684,N_49584,N_49739);
xor UO_3685 (O_3685,N_49969,N_49743);
and UO_3686 (O_3686,N_49551,N_49796);
xor UO_3687 (O_3687,N_49500,N_49592);
xor UO_3688 (O_3688,N_49729,N_49905);
or UO_3689 (O_3689,N_49814,N_49758);
nand UO_3690 (O_3690,N_49579,N_49698);
nand UO_3691 (O_3691,N_49538,N_49707);
and UO_3692 (O_3692,N_49739,N_49855);
nand UO_3693 (O_3693,N_49505,N_49764);
xor UO_3694 (O_3694,N_49580,N_49969);
nand UO_3695 (O_3695,N_49705,N_49797);
xor UO_3696 (O_3696,N_49747,N_49968);
and UO_3697 (O_3697,N_49902,N_49531);
nand UO_3698 (O_3698,N_49664,N_49964);
and UO_3699 (O_3699,N_49692,N_49698);
xnor UO_3700 (O_3700,N_49926,N_49528);
or UO_3701 (O_3701,N_49798,N_49525);
nand UO_3702 (O_3702,N_49875,N_49784);
xor UO_3703 (O_3703,N_49507,N_49670);
or UO_3704 (O_3704,N_49554,N_49656);
and UO_3705 (O_3705,N_49946,N_49513);
and UO_3706 (O_3706,N_49943,N_49617);
nor UO_3707 (O_3707,N_49765,N_49816);
nand UO_3708 (O_3708,N_49678,N_49504);
nor UO_3709 (O_3709,N_49534,N_49991);
xor UO_3710 (O_3710,N_49618,N_49659);
xnor UO_3711 (O_3711,N_49720,N_49874);
and UO_3712 (O_3712,N_49736,N_49647);
nor UO_3713 (O_3713,N_49666,N_49629);
or UO_3714 (O_3714,N_49733,N_49616);
and UO_3715 (O_3715,N_49845,N_49777);
nor UO_3716 (O_3716,N_49695,N_49658);
and UO_3717 (O_3717,N_49719,N_49950);
xnor UO_3718 (O_3718,N_49893,N_49501);
or UO_3719 (O_3719,N_49803,N_49867);
and UO_3720 (O_3720,N_49997,N_49987);
xor UO_3721 (O_3721,N_49986,N_49591);
and UO_3722 (O_3722,N_49954,N_49877);
xnor UO_3723 (O_3723,N_49983,N_49698);
or UO_3724 (O_3724,N_49695,N_49505);
nand UO_3725 (O_3725,N_49786,N_49548);
nand UO_3726 (O_3726,N_49871,N_49557);
or UO_3727 (O_3727,N_49691,N_49889);
and UO_3728 (O_3728,N_49701,N_49711);
and UO_3729 (O_3729,N_49685,N_49850);
nor UO_3730 (O_3730,N_49675,N_49603);
and UO_3731 (O_3731,N_49866,N_49604);
nand UO_3732 (O_3732,N_49609,N_49581);
nor UO_3733 (O_3733,N_49968,N_49614);
and UO_3734 (O_3734,N_49923,N_49642);
nor UO_3735 (O_3735,N_49917,N_49505);
or UO_3736 (O_3736,N_49978,N_49878);
nand UO_3737 (O_3737,N_49669,N_49604);
xor UO_3738 (O_3738,N_49738,N_49974);
nor UO_3739 (O_3739,N_49803,N_49984);
nand UO_3740 (O_3740,N_49627,N_49912);
or UO_3741 (O_3741,N_49695,N_49907);
nand UO_3742 (O_3742,N_49837,N_49508);
nor UO_3743 (O_3743,N_49663,N_49560);
and UO_3744 (O_3744,N_49848,N_49637);
xor UO_3745 (O_3745,N_49872,N_49928);
nand UO_3746 (O_3746,N_49510,N_49578);
and UO_3747 (O_3747,N_49971,N_49763);
or UO_3748 (O_3748,N_49911,N_49909);
nand UO_3749 (O_3749,N_49795,N_49545);
nand UO_3750 (O_3750,N_49673,N_49986);
and UO_3751 (O_3751,N_49898,N_49563);
and UO_3752 (O_3752,N_49771,N_49692);
xor UO_3753 (O_3753,N_49556,N_49851);
and UO_3754 (O_3754,N_49504,N_49522);
and UO_3755 (O_3755,N_49727,N_49630);
and UO_3756 (O_3756,N_49923,N_49779);
nor UO_3757 (O_3757,N_49642,N_49564);
nor UO_3758 (O_3758,N_49783,N_49545);
nand UO_3759 (O_3759,N_49926,N_49809);
or UO_3760 (O_3760,N_49647,N_49614);
or UO_3761 (O_3761,N_49943,N_49518);
and UO_3762 (O_3762,N_49518,N_49636);
nand UO_3763 (O_3763,N_49620,N_49770);
nor UO_3764 (O_3764,N_49753,N_49989);
nor UO_3765 (O_3765,N_49570,N_49753);
and UO_3766 (O_3766,N_49881,N_49500);
nor UO_3767 (O_3767,N_49926,N_49661);
or UO_3768 (O_3768,N_49535,N_49846);
nand UO_3769 (O_3769,N_49799,N_49515);
and UO_3770 (O_3770,N_49986,N_49694);
nor UO_3771 (O_3771,N_49765,N_49646);
xnor UO_3772 (O_3772,N_49942,N_49730);
nand UO_3773 (O_3773,N_49947,N_49959);
nand UO_3774 (O_3774,N_49788,N_49560);
xnor UO_3775 (O_3775,N_49867,N_49636);
nand UO_3776 (O_3776,N_49770,N_49927);
and UO_3777 (O_3777,N_49780,N_49665);
xor UO_3778 (O_3778,N_49559,N_49592);
xnor UO_3779 (O_3779,N_49740,N_49534);
or UO_3780 (O_3780,N_49768,N_49528);
and UO_3781 (O_3781,N_49851,N_49584);
nor UO_3782 (O_3782,N_49553,N_49621);
or UO_3783 (O_3783,N_49860,N_49922);
and UO_3784 (O_3784,N_49744,N_49825);
xor UO_3785 (O_3785,N_49775,N_49848);
nor UO_3786 (O_3786,N_49767,N_49584);
or UO_3787 (O_3787,N_49850,N_49773);
and UO_3788 (O_3788,N_49657,N_49731);
or UO_3789 (O_3789,N_49909,N_49807);
nand UO_3790 (O_3790,N_49789,N_49545);
or UO_3791 (O_3791,N_49920,N_49738);
nand UO_3792 (O_3792,N_49948,N_49673);
nand UO_3793 (O_3793,N_49752,N_49877);
xor UO_3794 (O_3794,N_49544,N_49877);
nand UO_3795 (O_3795,N_49816,N_49618);
and UO_3796 (O_3796,N_49781,N_49935);
xor UO_3797 (O_3797,N_49617,N_49518);
nand UO_3798 (O_3798,N_49782,N_49615);
xor UO_3799 (O_3799,N_49801,N_49812);
nor UO_3800 (O_3800,N_49918,N_49792);
nand UO_3801 (O_3801,N_49692,N_49786);
nor UO_3802 (O_3802,N_49642,N_49874);
or UO_3803 (O_3803,N_49707,N_49823);
nor UO_3804 (O_3804,N_49730,N_49905);
or UO_3805 (O_3805,N_49777,N_49668);
or UO_3806 (O_3806,N_49894,N_49618);
or UO_3807 (O_3807,N_49889,N_49678);
nor UO_3808 (O_3808,N_49571,N_49990);
nand UO_3809 (O_3809,N_49926,N_49739);
nor UO_3810 (O_3810,N_49963,N_49912);
xnor UO_3811 (O_3811,N_49514,N_49680);
and UO_3812 (O_3812,N_49741,N_49591);
and UO_3813 (O_3813,N_49760,N_49845);
nand UO_3814 (O_3814,N_49553,N_49970);
nor UO_3815 (O_3815,N_49587,N_49738);
nand UO_3816 (O_3816,N_49882,N_49630);
and UO_3817 (O_3817,N_49517,N_49973);
and UO_3818 (O_3818,N_49677,N_49795);
or UO_3819 (O_3819,N_49799,N_49983);
nand UO_3820 (O_3820,N_49944,N_49562);
and UO_3821 (O_3821,N_49533,N_49930);
and UO_3822 (O_3822,N_49803,N_49953);
and UO_3823 (O_3823,N_49992,N_49673);
and UO_3824 (O_3824,N_49727,N_49812);
nor UO_3825 (O_3825,N_49583,N_49633);
or UO_3826 (O_3826,N_49918,N_49720);
xor UO_3827 (O_3827,N_49739,N_49850);
and UO_3828 (O_3828,N_49841,N_49700);
or UO_3829 (O_3829,N_49902,N_49696);
nand UO_3830 (O_3830,N_49847,N_49954);
or UO_3831 (O_3831,N_49797,N_49970);
or UO_3832 (O_3832,N_49546,N_49573);
or UO_3833 (O_3833,N_49678,N_49712);
nor UO_3834 (O_3834,N_49960,N_49919);
and UO_3835 (O_3835,N_49585,N_49554);
nor UO_3836 (O_3836,N_49732,N_49707);
nor UO_3837 (O_3837,N_49525,N_49974);
nand UO_3838 (O_3838,N_49979,N_49843);
xnor UO_3839 (O_3839,N_49506,N_49742);
nor UO_3840 (O_3840,N_49650,N_49507);
nand UO_3841 (O_3841,N_49669,N_49679);
nor UO_3842 (O_3842,N_49691,N_49508);
nor UO_3843 (O_3843,N_49882,N_49576);
nand UO_3844 (O_3844,N_49750,N_49601);
and UO_3845 (O_3845,N_49708,N_49678);
and UO_3846 (O_3846,N_49925,N_49955);
and UO_3847 (O_3847,N_49995,N_49598);
or UO_3848 (O_3848,N_49816,N_49548);
and UO_3849 (O_3849,N_49506,N_49650);
and UO_3850 (O_3850,N_49793,N_49520);
xnor UO_3851 (O_3851,N_49522,N_49704);
nand UO_3852 (O_3852,N_49971,N_49672);
nand UO_3853 (O_3853,N_49952,N_49757);
or UO_3854 (O_3854,N_49796,N_49568);
nor UO_3855 (O_3855,N_49674,N_49543);
and UO_3856 (O_3856,N_49527,N_49603);
and UO_3857 (O_3857,N_49642,N_49750);
nand UO_3858 (O_3858,N_49806,N_49893);
nor UO_3859 (O_3859,N_49774,N_49723);
xnor UO_3860 (O_3860,N_49879,N_49596);
xor UO_3861 (O_3861,N_49506,N_49749);
nand UO_3862 (O_3862,N_49854,N_49711);
and UO_3863 (O_3863,N_49562,N_49500);
nor UO_3864 (O_3864,N_49718,N_49589);
or UO_3865 (O_3865,N_49663,N_49933);
nor UO_3866 (O_3866,N_49907,N_49666);
nand UO_3867 (O_3867,N_49944,N_49947);
and UO_3868 (O_3868,N_49848,N_49580);
and UO_3869 (O_3869,N_49779,N_49927);
nor UO_3870 (O_3870,N_49699,N_49534);
xor UO_3871 (O_3871,N_49954,N_49720);
xor UO_3872 (O_3872,N_49622,N_49745);
xnor UO_3873 (O_3873,N_49715,N_49669);
xor UO_3874 (O_3874,N_49740,N_49979);
and UO_3875 (O_3875,N_49526,N_49585);
and UO_3876 (O_3876,N_49501,N_49882);
or UO_3877 (O_3877,N_49748,N_49866);
xor UO_3878 (O_3878,N_49619,N_49902);
xnor UO_3879 (O_3879,N_49860,N_49793);
xor UO_3880 (O_3880,N_49869,N_49918);
xnor UO_3881 (O_3881,N_49689,N_49514);
xnor UO_3882 (O_3882,N_49996,N_49801);
nor UO_3883 (O_3883,N_49905,N_49594);
or UO_3884 (O_3884,N_49943,N_49596);
and UO_3885 (O_3885,N_49541,N_49891);
nand UO_3886 (O_3886,N_49770,N_49597);
xnor UO_3887 (O_3887,N_49684,N_49576);
or UO_3888 (O_3888,N_49518,N_49996);
xor UO_3889 (O_3889,N_49673,N_49741);
nand UO_3890 (O_3890,N_49889,N_49795);
nor UO_3891 (O_3891,N_49575,N_49815);
nor UO_3892 (O_3892,N_49961,N_49953);
xor UO_3893 (O_3893,N_49704,N_49545);
or UO_3894 (O_3894,N_49967,N_49707);
nor UO_3895 (O_3895,N_49628,N_49710);
and UO_3896 (O_3896,N_49830,N_49715);
nor UO_3897 (O_3897,N_49985,N_49732);
nor UO_3898 (O_3898,N_49818,N_49991);
nor UO_3899 (O_3899,N_49761,N_49635);
or UO_3900 (O_3900,N_49500,N_49643);
or UO_3901 (O_3901,N_49749,N_49681);
nand UO_3902 (O_3902,N_49699,N_49788);
nor UO_3903 (O_3903,N_49512,N_49764);
xnor UO_3904 (O_3904,N_49931,N_49508);
nand UO_3905 (O_3905,N_49967,N_49917);
xor UO_3906 (O_3906,N_49777,N_49731);
or UO_3907 (O_3907,N_49548,N_49678);
and UO_3908 (O_3908,N_49553,N_49609);
nand UO_3909 (O_3909,N_49782,N_49871);
and UO_3910 (O_3910,N_49593,N_49931);
xor UO_3911 (O_3911,N_49951,N_49617);
nor UO_3912 (O_3912,N_49941,N_49774);
and UO_3913 (O_3913,N_49932,N_49796);
or UO_3914 (O_3914,N_49822,N_49692);
nand UO_3915 (O_3915,N_49506,N_49852);
and UO_3916 (O_3916,N_49987,N_49691);
or UO_3917 (O_3917,N_49898,N_49955);
and UO_3918 (O_3918,N_49642,N_49607);
or UO_3919 (O_3919,N_49571,N_49979);
or UO_3920 (O_3920,N_49927,N_49751);
nor UO_3921 (O_3921,N_49557,N_49822);
nand UO_3922 (O_3922,N_49876,N_49706);
or UO_3923 (O_3923,N_49961,N_49772);
or UO_3924 (O_3924,N_49946,N_49656);
xnor UO_3925 (O_3925,N_49709,N_49805);
xnor UO_3926 (O_3926,N_49943,N_49627);
xor UO_3927 (O_3927,N_49570,N_49783);
xor UO_3928 (O_3928,N_49662,N_49852);
and UO_3929 (O_3929,N_49677,N_49932);
and UO_3930 (O_3930,N_49610,N_49614);
and UO_3931 (O_3931,N_49541,N_49643);
or UO_3932 (O_3932,N_49812,N_49945);
or UO_3933 (O_3933,N_49931,N_49771);
nor UO_3934 (O_3934,N_49825,N_49861);
and UO_3935 (O_3935,N_49996,N_49516);
nor UO_3936 (O_3936,N_49945,N_49609);
nand UO_3937 (O_3937,N_49791,N_49636);
or UO_3938 (O_3938,N_49933,N_49694);
and UO_3939 (O_3939,N_49857,N_49564);
xor UO_3940 (O_3940,N_49645,N_49799);
xor UO_3941 (O_3941,N_49803,N_49784);
or UO_3942 (O_3942,N_49507,N_49761);
nand UO_3943 (O_3943,N_49945,N_49838);
and UO_3944 (O_3944,N_49615,N_49993);
or UO_3945 (O_3945,N_49615,N_49864);
and UO_3946 (O_3946,N_49829,N_49723);
or UO_3947 (O_3947,N_49974,N_49863);
or UO_3948 (O_3948,N_49898,N_49960);
or UO_3949 (O_3949,N_49628,N_49795);
nand UO_3950 (O_3950,N_49953,N_49838);
or UO_3951 (O_3951,N_49537,N_49983);
nor UO_3952 (O_3952,N_49909,N_49779);
nor UO_3953 (O_3953,N_49558,N_49900);
nand UO_3954 (O_3954,N_49547,N_49884);
xor UO_3955 (O_3955,N_49788,N_49935);
nor UO_3956 (O_3956,N_49895,N_49862);
or UO_3957 (O_3957,N_49951,N_49991);
and UO_3958 (O_3958,N_49845,N_49766);
or UO_3959 (O_3959,N_49612,N_49885);
xor UO_3960 (O_3960,N_49818,N_49936);
nor UO_3961 (O_3961,N_49982,N_49962);
or UO_3962 (O_3962,N_49996,N_49740);
and UO_3963 (O_3963,N_49878,N_49676);
and UO_3964 (O_3964,N_49738,N_49942);
nor UO_3965 (O_3965,N_49935,N_49848);
xor UO_3966 (O_3966,N_49710,N_49752);
and UO_3967 (O_3967,N_49775,N_49713);
xor UO_3968 (O_3968,N_49770,N_49898);
or UO_3969 (O_3969,N_49752,N_49585);
nor UO_3970 (O_3970,N_49565,N_49568);
nand UO_3971 (O_3971,N_49919,N_49920);
and UO_3972 (O_3972,N_49766,N_49668);
xor UO_3973 (O_3973,N_49771,N_49726);
and UO_3974 (O_3974,N_49674,N_49936);
nand UO_3975 (O_3975,N_49860,N_49941);
xnor UO_3976 (O_3976,N_49872,N_49784);
or UO_3977 (O_3977,N_49904,N_49986);
nand UO_3978 (O_3978,N_49978,N_49575);
and UO_3979 (O_3979,N_49619,N_49828);
and UO_3980 (O_3980,N_49718,N_49878);
nand UO_3981 (O_3981,N_49718,N_49541);
and UO_3982 (O_3982,N_49578,N_49982);
nor UO_3983 (O_3983,N_49605,N_49924);
or UO_3984 (O_3984,N_49717,N_49926);
and UO_3985 (O_3985,N_49595,N_49715);
or UO_3986 (O_3986,N_49658,N_49591);
nor UO_3987 (O_3987,N_49522,N_49534);
nand UO_3988 (O_3988,N_49636,N_49878);
nor UO_3989 (O_3989,N_49701,N_49912);
xnor UO_3990 (O_3990,N_49687,N_49533);
nand UO_3991 (O_3991,N_49983,N_49882);
nor UO_3992 (O_3992,N_49872,N_49778);
or UO_3993 (O_3993,N_49593,N_49800);
nor UO_3994 (O_3994,N_49985,N_49584);
nor UO_3995 (O_3995,N_49574,N_49942);
nor UO_3996 (O_3996,N_49738,N_49928);
nand UO_3997 (O_3997,N_49516,N_49905);
nand UO_3998 (O_3998,N_49541,N_49851);
or UO_3999 (O_3999,N_49568,N_49586);
xnor UO_4000 (O_4000,N_49642,N_49672);
or UO_4001 (O_4001,N_49688,N_49862);
or UO_4002 (O_4002,N_49627,N_49512);
and UO_4003 (O_4003,N_49884,N_49881);
or UO_4004 (O_4004,N_49708,N_49763);
xor UO_4005 (O_4005,N_49602,N_49587);
nand UO_4006 (O_4006,N_49530,N_49616);
nor UO_4007 (O_4007,N_49884,N_49661);
or UO_4008 (O_4008,N_49541,N_49874);
nor UO_4009 (O_4009,N_49885,N_49911);
nor UO_4010 (O_4010,N_49766,N_49725);
nand UO_4011 (O_4011,N_49957,N_49934);
nor UO_4012 (O_4012,N_49878,N_49989);
nor UO_4013 (O_4013,N_49907,N_49611);
nand UO_4014 (O_4014,N_49705,N_49634);
nand UO_4015 (O_4015,N_49584,N_49866);
xor UO_4016 (O_4016,N_49533,N_49863);
nor UO_4017 (O_4017,N_49541,N_49665);
xnor UO_4018 (O_4018,N_49943,N_49521);
or UO_4019 (O_4019,N_49742,N_49794);
nor UO_4020 (O_4020,N_49600,N_49650);
nand UO_4021 (O_4021,N_49559,N_49567);
or UO_4022 (O_4022,N_49818,N_49619);
nand UO_4023 (O_4023,N_49935,N_49872);
nand UO_4024 (O_4024,N_49743,N_49539);
xnor UO_4025 (O_4025,N_49654,N_49947);
nor UO_4026 (O_4026,N_49852,N_49614);
nor UO_4027 (O_4027,N_49999,N_49544);
or UO_4028 (O_4028,N_49860,N_49672);
nand UO_4029 (O_4029,N_49928,N_49817);
nor UO_4030 (O_4030,N_49754,N_49585);
and UO_4031 (O_4031,N_49938,N_49684);
or UO_4032 (O_4032,N_49748,N_49936);
nor UO_4033 (O_4033,N_49729,N_49502);
xor UO_4034 (O_4034,N_49505,N_49996);
xor UO_4035 (O_4035,N_49963,N_49926);
nor UO_4036 (O_4036,N_49940,N_49724);
or UO_4037 (O_4037,N_49874,N_49943);
nor UO_4038 (O_4038,N_49768,N_49666);
nor UO_4039 (O_4039,N_49510,N_49968);
or UO_4040 (O_4040,N_49785,N_49842);
or UO_4041 (O_4041,N_49975,N_49540);
nand UO_4042 (O_4042,N_49567,N_49675);
or UO_4043 (O_4043,N_49665,N_49994);
xnor UO_4044 (O_4044,N_49896,N_49995);
nand UO_4045 (O_4045,N_49782,N_49910);
nand UO_4046 (O_4046,N_49548,N_49654);
and UO_4047 (O_4047,N_49565,N_49767);
nor UO_4048 (O_4048,N_49999,N_49926);
nor UO_4049 (O_4049,N_49958,N_49531);
nand UO_4050 (O_4050,N_49722,N_49743);
nor UO_4051 (O_4051,N_49507,N_49974);
xnor UO_4052 (O_4052,N_49845,N_49546);
xor UO_4053 (O_4053,N_49732,N_49568);
and UO_4054 (O_4054,N_49925,N_49510);
or UO_4055 (O_4055,N_49793,N_49724);
or UO_4056 (O_4056,N_49971,N_49930);
xor UO_4057 (O_4057,N_49608,N_49571);
nor UO_4058 (O_4058,N_49674,N_49939);
nor UO_4059 (O_4059,N_49713,N_49621);
xnor UO_4060 (O_4060,N_49830,N_49978);
or UO_4061 (O_4061,N_49518,N_49853);
and UO_4062 (O_4062,N_49855,N_49687);
or UO_4063 (O_4063,N_49748,N_49831);
xor UO_4064 (O_4064,N_49863,N_49528);
or UO_4065 (O_4065,N_49553,N_49778);
and UO_4066 (O_4066,N_49799,N_49978);
xor UO_4067 (O_4067,N_49543,N_49915);
nor UO_4068 (O_4068,N_49879,N_49536);
nand UO_4069 (O_4069,N_49841,N_49860);
nand UO_4070 (O_4070,N_49944,N_49514);
nor UO_4071 (O_4071,N_49518,N_49777);
nor UO_4072 (O_4072,N_49639,N_49629);
or UO_4073 (O_4073,N_49695,N_49571);
nor UO_4074 (O_4074,N_49569,N_49805);
and UO_4075 (O_4075,N_49564,N_49898);
nand UO_4076 (O_4076,N_49957,N_49749);
and UO_4077 (O_4077,N_49959,N_49963);
and UO_4078 (O_4078,N_49637,N_49793);
nor UO_4079 (O_4079,N_49975,N_49930);
or UO_4080 (O_4080,N_49756,N_49657);
xnor UO_4081 (O_4081,N_49796,N_49964);
and UO_4082 (O_4082,N_49894,N_49976);
nor UO_4083 (O_4083,N_49654,N_49722);
nor UO_4084 (O_4084,N_49692,N_49755);
nand UO_4085 (O_4085,N_49954,N_49941);
nor UO_4086 (O_4086,N_49753,N_49894);
xor UO_4087 (O_4087,N_49998,N_49575);
or UO_4088 (O_4088,N_49558,N_49541);
and UO_4089 (O_4089,N_49774,N_49698);
or UO_4090 (O_4090,N_49747,N_49504);
nor UO_4091 (O_4091,N_49962,N_49880);
nor UO_4092 (O_4092,N_49543,N_49721);
nor UO_4093 (O_4093,N_49969,N_49944);
nor UO_4094 (O_4094,N_49508,N_49641);
or UO_4095 (O_4095,N_49965,N_49543);
nand UO_4096 (O_4096,N_49748,N_49580);
nor UO_4097 (O_4097,N_49794,N_49700);
or UO_4098 (O_4098,N_49995,N_49906);
or UO_4099 (O_4099,N_49735,N_49773);
or UO_4100 (O_4100,N_49962,N_49870);
and UO_4101 (O_4101,N_49922,N_49681);
xor UO_4102 (O_4102,N_49624,N_49517);
and UO_4103 (O_4103,N_49945,N_49598);
or UO_4104 (O_4104,N_49899,N_49864);
and UO_4105 (O_4105,N_49711,N_49502);
nor UO_4106 (O_4106,N_49949,N_49936);
nor UO_4107 (O_4107,N_49740,N_49629);
nor UO_4108 (O_4108,N_49726,N_49980);
nand UO_4109 (O_4109,N_49796,N_49571);
nand UO_4110 (O_4110,N_49713,N_49828);
or UO_4111 (O_4111,N_49633,N_49939);
and UO_4112 (O_4112,N_49795,N_49527);
nand UO_4113 (O_4113,N_49830,N_49766);
and UO_4114 (O_4114,N_49598,N_49708);
and UO_4115 (O_4115,N_49518,N_49825);
nor UO_4116 (O_4116,N_49831,N_49544);
and UO_4117 (O_4117,N_49532,N_49789);
nor UO_4118 (O_4118,N_49581,N_49703);
or UO_4119 (O_4119,N_49822,N_49673);
xor UO_4120 (O_4120,N_49538,N_49586);
nand UO_4121 (O_4121,N_49739,N_49797);
nor UO_4122 (O_4122,N_49715,N_49921);
or UO_4123 (O_4123,N_49604,N_49929);
and UO_4124 (O_4124,N_49988,N_49626);
xor UO_4125 (O_4125,N_49833,N_49653);
and UO_4126 (O_4126,N_49617,N_49839);
or UO_4127 (O_4127,N_49654,N_49515);
xor UO_4128 (O_4128,N_49875,N_49659);
and UO_4129 (O_4129,N_49828,N_49768);
nor UO_4130 (O_4130,N_49926,N_49941);
and UO_4131 (O_4131,N_49770,N_49546);
nand UO_4132 (O_4132,N_49668,N_49812);
xor UO_4133 (O_4133,N_49767,N_49575);
nand UO_4134 (O_4134,N_49556,N_49924);
nor UO_4135 (O_4135,N_49593,N_49758);
xor UO_4136 (O_4136,N_49697,N_49593);
xnor UO_4137 (O_4137,N_49761,N_49855);
and UO_4138 (O_4138,N_49624,N_49767);
or UO_4139 (O_4139,N_49765,N_49709);
and UO_4140 (O_4140,N_49834,N_49535);
nor UO_4141 (O_4141,N_49624,N_49662);
or UO_4142 (O_4142,N_49847,N_49732);
nor UO_4143 (O_4143,N_49508,N_49713);
nand UO_4144 (O_4144,N_49955,N_49520);
or UO_4145 (O_4145,N_49945,N_49712);
or UO_4146 (O_4146,N_49854,N_49564);
nand UO_4147 (O_4147,N_49821,N_49955);
xnor UO_4148 (O_4148,N_49501,N_49814);
or UO_4149 (O_4149,N_49912,N_49569);
and UO_4150 (O_4150,N_49966,N_49977);
nor UO_4151 (O_4151,N_49946,N_49718);
xor UO_4152 (O_4152,N_49782,N_49732);
nor UO_4153 (O_4153,N_49941,N_49811);
and UO_4154 (O_4154,N_49563,N_49630);
xor UO_4155 (O_4155,N_49667,N_49686);
xnor UO_4156 (O_4156,N_49738,N_49831);
xnor UO_4157 (O_4157,N_49997,N_49611);
or UO_4158 (O_4158,N_49895,N_49934);
and UO_4159 (O_4159,N_49569,N_49850);
nand UO_4160 (O_4160,N_49994,N_49634);
xnor UO_4161 (O_4161,N_49597,N_49583);
nor UO_4162 (O_4162,N_49560,N_49905);
and UO_4163 (O_4163,N_49924,N_49841);
nor UO_4164 (O_4164,N_49524,N_49807);
and UO_4165 (O_4165,N_49934,N_49867);
or UO_4166 (O_4166,N_49758,N_49936);
nor UO_4167 (O_4167,N_49657,N_49921);
nor UO_4168 (O_4168,N_49786,N_49742);
and UO_4169 (O_4169,N_49726,N_49931);
nor UO_4170 (O_4170,N_49769,N_49787);
or UO_4171 (O_4171,N_49765,N_49503);
nor UO_4172 (O_4172,N_49863,N_49926);
nor UO_4173 (O_4173,N_49914,N_49981);
and UO_4174 (O_4174,N_49511,N_49786);
or UO_4175 (O_4175,N_49888,N_49570);
or UO_4176 (O_4176,N_49632,N_49805);
or UO_4177 (O_4177,N_49741,N_49820);
nor UO_4178 (O_4178,N_49831,N_49887);
nand UO_4179 (O_4179,N_49943,N_49541);
or UO_4180 (O_4180,N_49929,N_49979);
nand UO_4181 (O_4181,N_49921,N_49622);
nor UO_4182 (O_4182,N_49689,N_49639);
nor UO_4183 (O_4183,N_49756,N_49975);
xor UO_4184 (O_4184,N_49912,N_49709);
or UO_4185 (O_4185,N_49629,N_49931);
nor UO_4186 (O_4186,N_49943,N_49939);
nand UO_4187 (O_4187,N_49595,N_49957);
or UO_4188 (O_4188,N_49695,N_49778);
and UO_4189 (O_4189,N_49603,N_49967);
nand UO_4190 (O_4190,N_49539,N_49559);
and UO_4191 (O_4191,N_49751,N_49604);
and UO_4192 (O_4192,N_49830,N_49763);
xnor UO_4193 (O_4193,N_49827,N_49506);
and UO_4194 (O_4194,N_49693,N_49628);
or UO_4195 (O_4195,N_49947,N_49617);
nor UO_4196 (O_4196,N_49614,N_49917);
or UO_4197 (O_4197,N_49510,N_49919);
nand UO_4198 (O_4198,N_49945,N_49630);
nand UO_4199 (O_4199,N_49726,N_49807);
nand UO_4200 (O_4200,N_49636,N_49769);
xnor UO_4201 (O_4201,N_49621,N_49997);
nor UO_4202 (O_4202,N_49595,N_49741);
nand UO_4203 (O_4203,N_49900,N_49675);
xnor UO_4204 (O_4204,N_49616,N_49725);
nand UO_4205 (O_4205,N_49817,N_49743);
nor UO_4206 (O_4206,N_49676,N_49707);
nand UO_4207 (O_4207,N_49968,N_49858);
xnor UO_4208 (O_4208,N_49508,N_49797);
or UO_4209 (O_4209,N_49766,N_49723);
nor UO_4210 (O_4210,N_49508,N_49708);
or UO_4211 (O_4211,N_49870,N_49947);
nor UO_4212 (O_4212,N_49659,N_49845);
nor UO_4213 (O_4213,N_49699,N_49516);
and UO_4214 (O_4214,N_49945,N_49919);
and UO_4215 (O_4215,N_49881,N_49697);
and UO_4216 (O_4216,N_49661,N_49705);
and UO_4217 (O_4217,N_49846,N_49689);
nand UO_4218 (O_4218,N_49710,N_49864);
nor UO_4219 (O_4219,N_49793,N_49856);
or UO_4220 (O_4220,N_49772,N_49954);
nor UO_4221 (O_4221,N_49996,N_49823);
nor UO_4222 (O_4222,N_49526,N_49928);
xnor UO_4223 (O_4223,N_49588,N_49767);
and UO_4224 (O_4224,N_49694,N_49879);
or UO_4225 (O_4225,N_49781,N_49979);
nand UO_4226 (O_4226,N_49872,N_49825);
nand UO_4227 (O_4227,N_49825,N_49684);
nand UO_4228 (O_4228,N_49740,N_49924);
nand UO_4229 (O_4229,N_49780,N_49967);
nor UO_4230 (O_4230,N_49938,N_49617);
xnor UO_4231 (O_4231,N_49977,N_49744);
or UO_4232 (O_4232,N_49709,N_49580);
and UO_4233 (O_4233,N_49869,N_49973);
and UO_4234 (O_4234,N_49923,N_49978);
nand UO_4235 (O_4235,N_49586,N_49888);
xnor UO_4236 (O_4236,N_49919,N_49509);
and UO_4237 (O_4237,N_49698,N_49529);
xor UO_4238 (O_4238,N_49741,N_49902);
nor UO_4239 (O_4239,N_49573,N_49794);
nor UO_4240 (O_4240,N_49988,N_49784);
nor UO_4241 (O_4241,N_49557,N_49806);
xor UO_4242 (O_4242,N_49681,N_49952);
and UO_4243 (O_4243,N_49602,N_49864);
or UO_4244 (O_4244,N_49842,N_49529);
nand UO_4245 (O_4245,N_49919,N_49680);
xnor UO_4246 (O_4246,N_49884,N_49609);
nand UO_4247 (O_4247,N_49723,N_49929);
xnor UO_4248 (O_4248,N_49742,N_49717);
xor UO_4249 (O_4249,N_49535,N_49910);
nand UO_4250 (O_4250,N_49957,N_49949);
or UO_4251 (O_4251,N_49593,N_49598);
nand UO_4252 (O_4252,N_49734,N_49778);
nand UO_4253 (O_4253,N_49631,N_49546);
nand UO_4254 (O_4254,N_49888,N_49556);
nor UO_4255 (O_4255,N_49674,N_49989);
or UO_4256 (O_4256,N_49953,N_49738);
or UO_4257 (O_4257,N_49996,N_49598);
xor UO_4258 (O_4258,N_49760,N_49907);
or UO_4259 (O_4259,N_49872,N_49545);
or UO_4260 (O_4260,N_49613,N_49612);
or UO_4261 (O_4261,N_49973,N_49992);
xnor UO_4262 (O_4262,N_49959,N_49503);
and UO_4263 (O_4263,N_49979,N_49901);
or UO_4264 (O_4264,N_49647,N_49905);
nor UO_4265 (O_4265,N_49546,N_49637);
or UO_4266 (O_4266,N_49566,N_49912);
or UO_4267 (O_4267,N_49581,N_49641);
nand UO_4268 (O_4268,N_49579,N_49938);
and UO_4269 (O_4269,N_49770,N_49904);
nor UO_4270 (O_4270,N_49887,N_49978);
nor UO_4271 (O_4271,N_49838,N_49850);
nand UO_4272 (O_4272,N_49794,N_49544);
xor UO_4273 (O_4273,N_49676,N_49942);
or UO_4274 (O_4274,N_49923,N_49611);
and UO_4275 (O_4275,N_49977,N_49561);
nand UO_4276 (O_4276,N_49631,N_49697);
xnor UO_4277 (O_4277,N_49792,N_49547);
nand UO_4278 (O_4278,N_49942,N_49543);
or UO_4279 (O_4279,N_49535,N_49922);
and UO_4280 (O_4280,N_49697,N_49588);
or UO_4281 (O_4281,N_49777,N_49516);
or UO_4282 (O_4282,N_49503,N_49792);
nand UO_4283 (O_4283,N_49950,N_49559);
nand UO_4284 (O_4284,N_49692,N_49891);
or UO_4285 (O_4285,N_49524,N_49931);
nor UO_4286 (O_4286,N_49570,N_49504);
nor UO_4287 (O_4287,N_49539,N_49702);
or UO_4288 (O_4288,N_49620,N_49905);
xnor UO_4289 (O_4289,N_49643,N_49529);
and UO_4290 (O_4290,N_49959,N_49537);
nand UO_4291 (O_4291,N_49941,N_49731);
nand UO_4292 (O_4292,N_49790,N_49871);
nand UO_4293 (O_4293,N_49734,N_49732);
nand UO_4294 (O_4294,N_49861,N_49796);
nand UO_4295 (O_4295,N_49996,N_49537);
and UO_4296 (O_4296,N_49784,N_49849);
nor UO_4297 (O_4297,N_49792,N_49763);
and UO_4298 (O_4298,N_49758,N_49673);
and UO_4299 (O_4299,N_49660,N_49547);
nand UO_4300 (O_4300,N_49527,N_49597);
xnor UO_4301 (O_4301,N_49586,N_49851);
or UO_4302 (O_4302,N_49939,N_49617);
nand UO_4303 (O_4303,N_49631,N_49955);
or UO_4304 (O_4304,N_49570,N_49610);
and UO_4305 (O_4305,N_49527,N_49652);
or UO_4306 (O_4306,N_49951,N_49654);
and UO_4307 (O_4307,N_49567,N_49690);
nor UO_4308 (O_4308,N_49742,N_49650);
xnor UO_4309 (O_4309,N_49899,N_49539);
and UO_4310 (O_4310,N_49985,N_49949);
xnor UO_4311 (O_4311,N_49832,N_49827);
xnor UO_4312 (O_4312,N_49790,N_49910);
xor UO_4313 (O_4313,N_49664,N_49689);
or UO_4314 (O_4314,N_49941,N_49698);
or UO_4315 (O_4315,N_49845,N_49933);
nor UO_4316 (O_4316,N_49508,N_49895);
or UO_4317 (O_4317,N_49539,N_49755);
nor UO_4318 (O_4318,N_49919,N_49970);
nor UO_4319 (O_4319,N_49678,N_49815);
and UO_4320 (O_4320,N_49935,N_49900);
nand UO_4321 (O_4321,N_49943,N_49630);
xor UO_4322 (O_4322,N_49883,N_49830);
and UO_4323 (O_4323,N_49533,N_49833);
nor UO_4324 (O_4324,N_49867,N_49620);
nand UO_4325 (O_4325,N_49894,N_49738);
nand UO_4326 (O_4326,N_49777,N_49754);
and UO_4327 (O_4327,N_49829,N_49946);
nor UO_4328 (O_4328,N_49731,N_49619);
xnor UO_4329 (O_4329,N_49870,N_49939);
or UO_4330 (O_4330,N_49731,N_49669);
xor UO_4331 (O_4331,N_49626,N_49644);
or UO_4332 (O_4332,N_49685,N_49942);
or UO_4333 (O_4333,N_49712,N_49958);
nand UO_4334 (O_4334,N_49719,N_49779);
nor UO_4335 (O_4335,N_49554,N_49851);
xnor UO_4336 (O_4336,N_49683,N_49805);
or UO_4337 (O_4337,N_49949,N_49575);
xor UO_4338 (O_4338,N_49573,N_49713);
xor UO_4339 (O_4339,N_49932,N_49811);
nor UO_4340 (O_4340,N_49786,N_49702);
or UO_4341 (O_4341,N_49846,N_49973);
and UO_4342 (O_4342,N_49761,N_49830);
or UO_4343 (O_4343,N_49832,N_49809);
xor UO_4344 (O_4344,N_49898,N_49818);
or UO_4345 (O_4345,N_49565,N_49580);
xor UO_4346 (O_4346,N_49724,N_49881);
or UO_4347 (O_4347,N_49792,N_49764);
or UO_4348 (O_4348,N_49562,N_49756);
and UO_4349 (O_4349,N_49616,N_49986);
nor UO_4350 (O_4350,N_49575,N_49764);
nand UO_4351 (O_4351,N_49659,N_49606);
nor UO_4352 (O_4352,N_49811,N_49967);
xor UO_4353 (O_4353,N_49861,N_49961);
nand UO_4354 (O_4354,N_49914,N_49515);
or UO_4355 (O_4355,N_49967,N_49875);
nand UO_4356 (O_4356,N_49924,N_49715);
xor UO_4357 (O_4357,N_49712,N_49589);
nand UO_4358 (O_4358,N_49876,N_49520);
xor UO_4359 (O_4359,N_49812,N_49521);
nor UO_4360 (O_4360,N_49679,N_49636);
or UO_4361 (O_4361,N_49953,N_49641);
and UO_4362 (O_4362,N_49549,N_49862);
nor UO_4363 (O_4363,N_49510,N_49780);
nand UO_4364 (O_4364,N_49922,N_49866);
nor UO_4365 (O_4365,N_49669,N_49553);
xnor UO_4366 (O_4366,N_49765,N_49946);
nand UO_4367 (O_4367,N_49706,N_49570);
xor UO_4368 (O_4368,N_49798,N_49563);
nor UO_4369 (O_4369,N_49542,N_49844);
or UO_4370 (O_4370,N_49783,N_49920);
or UO_4371 (O_4371,N_49925,N_49561);
xor UO_4372 (O_4372,N_49683,N_49635);
and UO_4373 (O_4373,N_49746,N_49576);
nand UO_4374 (O_4374,N_49504,N_49741);
nand UO_4375 (O_4375,N_49643,N_49566);
xor UO_4376 (O_4376,N_49864,N_49586);
nor UO_4377 (O_4377,N_49660,N_49591);
xor UO_4378 (O_4378,N_49843,N_49515);
nand UO_4379 (O_4379,N_49714,N_49603);
nand UO_4380 (O_4380,N_49706,N_49763);
xor UO_4381 (O_4381,N_49762,N_49928);
and UO_4382 (O_4382,N_49740,N_49897);
or UO_4383 (O_4383,N_49826,N_49930);
and UO_4384 (O_4384,N_49780,N_49728);
xnor UO_4385 (O_4385,N_49823,N_49899);
nor UO_4386 (O_4386,N_49936,N_49952);
nor UO_4387 (O_4387,N_49978,N_49937);
nor UO_4388 (O_4388,N_49593,N_49835);
or UO_4389 (O_4389,N_49510,N_49833);
or UO_4390 (O_4390,N_49849,N_49657);
or UO_4391 (O_4391,N_49514,N_49857);
nand UO_4392 (O_4392,N_49986,N_49581);
or UO_4393 (O_4393,N_49970,N_49793);
and UO_4394 (O_4394,N_49813,N_49595);
or UO_4395 (O_4395,N_49832,N_49904);
xnor UO_4396 (O_4396,N_49822,N_49925);
and UO_4397 (O_4397,N_49902,N_49584);
xnor UO_4398 (O_4398,N_49951,N_49747);
nand UO_4399 (O_4399,N_49730,N_49886);
and UO_4400 (O_4400,N_49989,N_49936);
and UO_4401 (O_4401,N_49861,N_49652);
nor UO_4402 (O_4402,N_49702,N_49993);
xor UO_4403 (O_4403,N_49767,N_49948);
nand UO_4404 (O_4404,N_49735,N_49867);
nor UO_4405 (O_4405,N_49905,N_49794);
nand UO_4406 (O_4406,N_49579,N_49665);
or UO_4407 (O_4407,N_49501,N_49755);
or UO_4408 (O_4408,N_49764,N_49556);
xor UO_4409 (O_4409,N_49702,N_49976);
and UO_4410 (O_4410,N_49525,N_49746);
nor UO_4411 (O_4411,N_49577,N_49875);
or UO_4412 (O_4412,N_49831,N_49553);
xor UO_4413 (O_4413,N_49595,N_49830);
nand UO_4414 (O_4414,N_49722,N_49867);
nor UO_4415 (O_4415,N_49731,N_49609);
and UO_4416 (O_4416,N_49625,N_49755);
nor UO_4417 (O_4417,N_49654,N_49991);
and UO_4418 (O_4418,N_49882,N_49671);
xnor UO_4419 (O_4419,N_49503,N_49839);
nand UO_4420 (O_4420,N_49587,N_49677);
and UO_4421 (O_4421,N_49688,N_49889);
and UO_4422 (O_4422,N_49908,N_49755);
nor UO_4423 (O_4423,N_49836,N_49815);
and UO_4424 (O_4424,N_49620,N_49680);
and UO_4425 (O_4425,N_49671,N_49884);
xnor UO_4426 (O_4426,N_49959,N_49562);
or UO_4427 (O_4427,N_49985,N_49825);
nor UO_4428 (O_4428,N_49598,N_49758);
or UO_4429 (O_4429,N_49709,N_49673);
nand UO_4430 (O_4430,N_49870,N_49988);
or UO_4431 (O_4431,N_49819,N_49874);
nand UO_4432 (O_4432,N_49567,N_49743);
nand UO_4433 (O_4433,N_49930,N_49912);
nand UO_4434 (O_4434,N_49958,N_49832);
nand UO_4435 (O_4435,N_49716,N_49509);
nand UO_4436 (O_4436,N_49831,N_49878);
and UO_4437 (O_4437,N_49891,N_49501);
nor UO_4438 (O_4438,N_49826,N_49524);
xnor UO_4439 (O_4439,N_49617,N_49848);
and UO_4440 (O_4440,N_49827,N_49734);
nand UO_4441 (O_4441,N_49544,N_49848);
and UO_4442 (O_4442,N_49673,N_49788);
xnor UO_4443 (O_4443,N_49729,N_49701);
and UO_4444 (O_4444,N_49887,N_49974);
and UO_4445 (O_4445,N_49940,N_49992);
and UO_4446 (O_4446,N_49565,N_49506);
xor UO_4447 (O_4447,N_49651,N_49673);
nand UO_4448 (O_4448,N_49593,N_49755);
nand UO_4449 (O_4449,N_49765,N_49570);
and UO_4450 (O_4450,N_49778,N_49937);
nor UO_4451 (O_4451,N_49677,N_49936);
xnor UO_4452 (O_4452,N_49642,N_49856);
nor UO_4453 (O_4453,N_49866,N_49805);
nor UO_4454 (O_4454,N_49603,N_49841);
nand UO_4455 (O_4455,N_49821,N_49621);
xnor UO_4456 (O_4456,N_49523,N_49628);
nor UO_4457 (O_4457,N_49833,N_49742);
nand UO_4458 (O_4458,N_49506,N_49874);
nor UO_4459 (O_4459,N_49683,N_49727);
nand UO_4460 (O_4460,N_49552,N_49835);
or UO_4461 (O_4461,N_49888,N_49712);
nor UO_4462 (O_4462,N_49715,N_49817);
nand UO_4463 (O_4463,N_49503,N_49774);
nor UO_4464 (O_4464,N_49820,N_49601);
or UO_4465 (O_4465,N_49972,N_49876);
and UO_4466 (O_4466,N_49526,N_49926);
nor UO_4467 (O_4467,N_49570,N_49994);
nor UO_4468 (O_4468,N_49574,N_49734);
and UO_4469 (O_4469,N_49662,N_49683);
nand UO_4470 (O_4470,N_49585,N_49733);
nand UO_4471 (O_4471,N_49736,N_49559);
and UO_4472 (O_4472,N_49765,N_49976);
nand UO_4473 (O_4473,N_49577,N_49843);
and UO_4474 (O_4474,N_49836,N_49886);
nand UO_4475 (O_4475,N_49525,N_49583);
nor UO_4476 (O_4476,N_49735,N_49995);
nand UO_4477 (O_4477,N_49982,N_49979);
or UO_4478 (O_4478,N_49661,N_49566);
or UO_4479 (O_4479,N_49744,N_49523);
or UO_4480 (O_4480,N_49515,N_49524);
and UO_4481 (O_4481,N_49880,N_49848);
xnor UO_4482 (O_4482,N_49982,N_49932);
nand UO_4483 (O_4483,N_49775,N_49558);
and UO_4484 (O_4484,N_49959,N_49548);
nor UO_4485 (O_4485,N_49766,N_49563);
and UO_4486 (O_4486,N_49849,N_49824);
and UO_4487 (O_4487,N_49717,N_49987);
and UO_4488 (O_4488,N_49691,N_49955);
nor UO_4489 (O_4489,N_49797,N_49758);
nor UO_4490 (O_4490,N_49605,N_49780);
and UO_4491 (O_4491,N_49801,N_49955);
nand UO_4492 (O_4492,N_49994,N_49831);
or UO_4493 (O_4493,N_49839,N_49773);
nand UO_4494 (O_4494,N_49531,N_49851);
or UO_4495 (O_4495,N_49765,N_49712);
nand UO_4496 (O_4496,N_49998,N_49638);
xor UO_4497 (O_4497,N_49761,N_49512);
and UO_4498 (O_4498,N_49844,N_49981);
and UO_4499 (O_4499,N_49943,N_49650);
nand UO_4500 (O_4500,N_49977,N_49997);
nand UO_4501 (O_4501,N_49722,N_49929);
nor UO_4502 (O_4502,N_49599,N_49991);
or UO_4503 (O_4503,N_49507,N_49672);
and UO_4504 (O_4504,N_49980,N_49556);
or UO_4505 (O_4505,N_49677,N_49824);
or UO_4506 (O_4506,N_49755,N_49995);
nor UO_4507 (O_4507,N_49984,N_49992);
nand UO_4508 (O_4508,N_49698,N_49727);
xor UO_4509 (O_4509,N_49584,N_49612);
and UO_4510 (O_4510,N_49776,N_49742);
or UO_4511 (O_4511,N_49527,N_49879);
xor UO_4512 (O_4512,N_49755,N_49658);
and UO_4513 (O_4513,N_49844,N_49925);
nand UO_4514 (O_4514,N_49562,N_49705);
nor UO_4515 (O_4515,N_49558,N_49517);
and UO_4516 (O_4516,N_49755,N_49595);
and UO_4517 (O_4517,N_49957,N_49516);
xnor UO_4518 (O_4518,N_49569,N_49736);
nand UO_4519 (O_4519,N_49565,N_49696);
nor UO_4520 (O_4520,N_49906,N_49690);
nand UO_4521 (O_4521,N_49970,N_49729);
nor UO_4522 (O_4522,N_49903,N_49628);
or UO_4523 (O_4523,N_49603,N_49996);
or UO_4524 (O_4524,N_49575,N_49754);
xor UO_4525 (O_4525,N_49665,N_49927);
xor UO_4526 (O_4526,N_49927,N_49707);
and UO_4527 (O_4527,N_49561,N_49932);
nand UO_4528 (O_4528,N_49585,N_49879);
nor UO_4529 (O_4529,N_49744,N_49636);
nand UO_4530 (O_4530,N_49953,N_49899);
xnor UO_4531 (O_4531,N_49590,N_49604);
xnor UO_4532 (O_4532,N_49855,N_49518);
and UO_4533 (O_4533,N_49886,N_49849);
nor UO_4534 (O_4534,N_49642,N_49614);
or UO_4535 (O_4535,N_49819,N_49620);
xnor UO_4536 (O_4536,N_49583,N_49745);
nand UO_4537 (O_4537,N_49805,N_49945);
nor UO_4538 (O_4538,N_49807,N_49624);
nand UO_4539 (O_4539,N_49630,N_49644);
and UO_4540 (O_4540,N_49738,N_49994);
xor UO_4541 (O_4541,N_49944,N_49900);
or UO_4542 (O_4542,N_49575,N_49878);
and UO_4543 (O_4543,N_49846,N_49856);
xor UO_4544 (O_4544,N_49871,N_49825);
xor UO_4545 (O_4545,N_49532,N_49586);
xnor UO_4546 (O_4546,N_49837,N_49764);
and UO_4547 (O_4547,N_49756,N_49551);
and UO_4548 (O_4548,N_49714,N_49528);
and UO_4549 (O_4549,N_49746,N_49981);
or UO_4550 (O_4550,N_49927,N_49827);
and UO_4551 (O_4551,N_49851,N_49500);
nor UO_4552 (O_4552,N_49754,N_49567);
xnor UO_4553 (O_4553,N_49929,N_49933);
nand UO_4554 (O_4554,N_49582,N_49559);
nand UO_4555 (O_4555,N_49632,N_49619);
xor UO_4556 (O_4556,N_49881,N_49864);
and UO_4557 (O_4557,N_49883,N_49674);
nor UO_4558 (O_4558,N_49928,N_49541);
and UO_4559 (O_4559,N_49776,N_49531);
xor UO_4560 (O_4560,N_49850,N_49866);
nand UO_4561 (O_4561,N_49557,N_49660);
xnor UO_4562 (O_4562,N_49615,N_49751);
xor UO_4563 (O_4563,N_49589,N_49929);
or UO_4564 (O_4564,N_49671,N_49529);
and UO_4565 (O_4565,N_49851,N_49861);
and UO_4566 (O_4566,N_49932,N_49703);
xor UO_4567 (O_4567,N_49971,N_49807);
or UO_4568 (O_4568,N_49786,N_49864);
nand UO_4569 (O_4569,N_49758,N_49602);
nor UO_4570 (O_4570,N_49624,N_49648);
or UO_4571 (O_4571,N_49866,N_49702);
and UO_4572 (O_4572,N_49762,N_49873);
and UO_4573 (O_4573,N_49768,N_49530);
nand UO_4574 (O_4574,N_49802,N_49636);
nand UO_4575 (O_4575,N_49773,N_49574);
xnor UO_4576 (O_4576,N_49519,N_49921);
or UO_4577 (O_4577,N_49658,N_49535);
nand UO_4578 (O_4578,N_49707,N_49842);
or UO_4579 (O_4579,N_49723,N_49595);
xor UO_4580 (O_4580,N_49890,N_49510);
xor UO_4581 (O_4581,N_49558,N_49956);
nor UO_4582 (O_4582,N_49625,N_49759);
or UO_4583 (O_4583,N_49957,N_49985);
or UO_4584 (O_4584,N_49568,N_49842);
nand UO_4585 (O_4585,N_49621,N_49509);
or UO_4586 (O_4586,N_49501,N_49787);
nor UO_4587 (O_4587,N_49597,N_49685);
and UO_4588 (O_4588,N_49547,N_49944);
and UO_4589 (O_4589,N_49988,N_49536);
nand UO_4590 (O_4590,N_49862,N_49656);
xnor UO_4591 (O_4591,N_49679,N_49732);
and UO_4592 (O_4592,N_49719,N_49664);
nand UO_4593 (O_4593,N_49538,N_49876);
nand UO_4594 (O_4594,N_49916,N_49585);
or UO_4595 (O_4595,N_49595,N_49834);
and UO_4596 (O_4596,N_49958,N_49510);
nand UO_4597 (O_4597,N_49955,N_49844);
nand UO_4598 (O_4598,N_49841,N_49566);
and UO_4599 (O_4599,N_49982,N_49969);
nand UO_4600 (O_4600,N_49694,N_49680);
and UO_4601 (O_4601,N_49532,N_49665);
and UO_4602 (O_4602,N_49954,N_49818);
xor UO_4603 (O_4603,N_49816,N_49701);
nor UO_4604 (O_4604,N_49979,N_49654);
nor UO_4605 (O_4605,N_49962,N_49956);
xor UO_4606 (O_4606,N_49862,N_49715);
nor UO_4607 (O_4607,N_49695,N_49768);
nor UO_4608 (O_4608,N_49534,N_49948);
or UO_4609 (O_4609,N_49862,N_49922);
nand UO_4610 (O_4610,N_49876,N_49642);
nand UO_4611 (O_4611,N_49926,N_49879);
or UO_4612 (O_4612,N_49721,N_49585);
xnor UO_4613 (O_4613,N_49820,N_49550);
and UO_4614 (O_4614,N_49937,N_49516);
nor UO_4615 (O_4615,N_49951,N_49763);
and UO_4616 (O_4616,N_49870,N_49535);
and UO_4617 (O_4617,N_49550,N_49596);
and UO_4618 (O_4618,N_49680,N_49634);
or UO_4619 (O_4619,N_49922,N_49789);
or UO_4620 (O_4620,N_49876,N_49627);
nand UO_4621 (O_4621,N_49711,N_49641);
and UO_4622 (O_4622,N_49509,N_49570);
and UO_4623 (O_4623,N_49510,N_49883);
nor UO_4624 (O_4624,N_49611,N_49654);
or UO_4625 (O_4625,N_49517,N_49678);
or UO_4626 (O_4626,N_49959,N_49732);
nor UO_4627 (O_4627,N_49610,N_49960);
or UO_4628 (O_4628,N_49867,N_49834);
nor UO_4629 (O_4629,N_49745,N_49888);
xnor UO_4630 (O_4630,N_49715,N_49872);
xor UO_4631 (O_4631,N_49790,N_49686);
nand UO_4632 (O_4632,N_49837,N_49503);
nand UO_4633 (O_4633,N_49963,N_49720);
nor UO_4634 (O_4634,N_49798,N_49896);
xnor UO_4635 (O_4635,N_49924,N_49575);
or UO_4636 (O_4636,N_49873,N_49957);
nor UO_4637 (O_4637,N_49653,N_49575);
xnor UO_4638 (O_4638,N_49693,N_49635);
nor UO_4639 (O_4639,N_49697,N_49842);
nor UO_4640 (O_4640,N_49834,N_49861);
nor UO_4641 (O_4641,N_49790,N_49849);
xor UO_4642 (O_4642,N_49975,N_49878);
and UO_4643 (O_4643,N_49547,N_49879);
nand UO_4644 (O_4644,N_49652,N_49864);
xnor UO_4645 (O_4645,N_49971,N_49704);
and UO_4646 (O_4646,N_49837,N_49782);
xor UO_4647 (O_4647,N_49877,N_49579);
nor UO_4648 (O_4648,N_49976,N_49924);
and UO_4649 (O_4649,N_49538,N_49555);
nand UO_4650 (O_4650,N_49857,N_49551);
nor UO_4651 (O_4651,N_49836,N_49984);
and UO_4652 (O_4652,N_49906,N_49606);
nor UO_4653 (O_4653,N_49793,N_49610);
nand UO_4654 (O_4654,N_49522,N_49750);
or UO_4655 (O_4655,N_49680,N_49679);
nor UO_4656 (O_4656,N_49891,N_49540);
xnor UO_4657 (O_4657,N_49563,N_49663);
and UO_4658 (O_4658,N_49709,N_49986);
or UO_4659 (O_4659,N_49681,N_49678);
nand UO_4660 (O_4660,N_49931,N_49589);
nand UO_4661 (O_4661,N_49534,N_49672);
xnor UO_4662 (O_4662,N_49805,N_49740);
and UO_4663 (O_4663,N_49745,N_49787);
or UO_4664 (O_4664,N_49692,N_49875);
and UO_4665 (O_4665,N_49683,N_49506);
or UO_4666 (O_4666,N_49719,N_49755);
and UO_4667 (O_4667,N_49872,N_49896);
nand UO_4668 (O_4668,N_49911,N_49614);
nand UO_4669 (O_4669,N_49826,N_49689);
nand UO_4670 (O_4670,N_49927,N_49539);
xor UO_4671 (O_4671,N_49611,N_49769);
nand UO_4672 (O_4672,N_49568,N_49718);
xnor UO_4673 (O_4673,N_49782,N_49717);
and UO_4674 (O_4674,N_49972,N_49915);
xnor UO_4675 (O_4675,N_49858,N_49886);
xor UO_4676 (O_4676,N_49528,N_49507);
nand UO_4677 (O_4677,N_49940,N_49946);
nand UO_4678 (O_4678,N_49643,N_49851);
or UO_4679 (O_4679,N_49633,N_49678);
or UO_4680 (O_4680,N_49983,N_49867);
nor UO_4681 (O_4681,N_49740,N_49786);
or UO_4682 (O_4682,N_49679,N_49526);
nor UO_4683 (O_4683,N_49537,N_49793);
and UO_4684 (O_4684,N_49902,N_49778);
and UO_4685 (O_4685,N_49719,N_49815);
nand UO_4686 (O_4686,N_49971,N_49615);
or UO_4687 (O_4687,N_49502,N_49916);
nor UO_4688 (O_4688,N_49590,N_49992);
and UO_4689 (O_4689,N_49915,N_49683);
and UO_4690 (O_4690,N_49541,N_49940);
nand UO_4691 (O_4691,N_49667,N_49545);
or UO_4692 (O_4692,N_49768,N_49889);
or UO_4693 (O_4693,N_49998,N_49865);
and UO_4694 (O_4694,N_49949,N_49911);
nor UO_4695 (O_4695,N_49950,N_49977);
xor UO_4696 (O_4696,N_49507,N_49824);
nand UO_4697 (O_4697,N_49674,N_49908);
nor UO_4698 (O_4698,N_49960,N_49933);
and UO_4699 (O_4699,N_49966,N_49611);
xnor UO_4700 (O_4700,N_49760,N_49915);
nor UO_4701 (O_4701,N_49855,N_49681);
or UO_4702 (O_4702,N_49788,N_49724);
nor UO_4703 (O_4703,N_49552,N_49795);
nor UO_4704 (O_4704,N_49826,N_49519);
nand UO_4705 (O_4705,N_49556,N_49968);
nand UO_4706 (O_4706,N_49596,N_49573);
nor UO_4707 (O_4707,N_49650,N_49810);
or UO_4708 (O_4708,N_49850,N_49762);
or UO_4709 (O_4709,N_49540,N_49545);
nor UO_4710 (O_4710,N_49984,N_49669);
nor UO_4711 (O_4711,N_49554,N_49830);
or UO_4712 (O_4712,N_49849,N_49777);
xnor UO_4713 (O_4713,N_49839,N_49622);
or UO_4714 (O_4714,N_49805,N_49690);
xor UO_4715 (O_4715,N_49814,N_49976);
nor UO_4716 (O_4716,N_49774,N_49862);
nor UO_4717 (O_4717,N_49520,N_49505);
and UO_4718 (O_4718,N_49737,N_49582);
and UO_4719 (O_4719,N_49818,N_49723);
xnor UO_4720 (O_4720,N_49661,N_49750);
or UO_4721 (O_4721,N_49635,N_49741);
nand UO_4722 (O_4722,N_49836,N_49688);
and UO_4723 (O_4723,N_49722,N_49957);
xor UO_4724 (O_4724,N_49697,N_49949);
nor UO_4725 (O_4725,N_49574,N_49579);
nand UO_4726 (O_4726,N_49910,N_49978);
nand UO_4727 (O_4727,N_49876,N_49964);
or UO_4728 (O_4728,N_49946,N_49771);
xor UO_4729 (O_4729,N_49802,N_49610);
xnor UO_4730 (O_4730,N_49724,N_49697);
or UO_4731 (O_4731,N_49522,N_49949);
nor UO_4732 (O_4732,N_49744,N_49845);
nor UO_4733 (O_4733,N_49920,N_49640);
xor UO_4734 (O_4734,N_49681,N_49518);
nand UO_4735 (O_4735,N_49942,N_49555);
and UO_4736 (O_4736,N_49773,N_49701);
or UO_4737 (O_4737,N_49761,N_49871);
or UO_4738 (O_4738,N_49651,N_49643);
or UO_4739 (O_4739,N_49633,N_49908);
or UO_4740 (O_4740,N_49527,N_49598);
or UO_4741 (O_4741,N_49618,N_49940);
nor UO_4742 (O_4742,N_49500,N_49950);
xnor UO_4743 (O_4743,N_49566,N_49674);
nor UO_4744 (O_4744,N_49783,N_49789);
nand UO_4745 (O_4745,N_49861,N_49741);
or UO_4746 (O_4746,N_49529,N_49716);
or UO_4747 (O_4747,N_49684,N_49962);
xor UO_4748 (O_4748,N_49744,N_49782);
nor UO_4749 (O_4749,N_49723,N_49534);
or UO_4750 (O_4750,N_49868,N_49585);
and UO_4751 (O_4751,N_49731,N_49856);
or UO_4752 (O_4752,N_49784,N_49789);
xnor UO_4753 (O_4753,N_49753,N_49745);
nand UO_4754 (O_4754,N_49904,N_49731);
nor UO_4755 (O_4755,N_49949,N_49819);
xor UO_4756 (O_4756,N_49990,N_49620);
nor UO_4757 (O_4757,N_49503,N_49686);
nor UO_4758 (O_4758,N_49610,N_49579);
or UO_4759 (O_4759,N_49663,N_49921);
and UO_4760 (O_4760,N_49586,N_49647);
xnor UO_4761 (O_4761,N_49907,N_49751);
xnor UO_4762 (O_4762,N_49589,N_49672);
or UO_4763 (O_4763,N_49783,N_49557);
xor UO_4764 (O_4764,N_49644,N_49662);
or UO_4765 (O_4765,N_49628,N_49558);
xor UO_4766 (O_4766,N_49899,N_49553);
nor UO_4767 (O_4767,N_49566,N_49530);
nand UO_4768 (O_4768,N_49567,N_49663);
nor UO_4769 (O_4769,N_49869,N_49810);
and UO_4770 (O_4770,N_49919,N_49800);
nand UO_4771 (O_4771,N_49760,N_49656);
and UO_4772 (O_4772,N_49742,N_49827);
or UO_4773 (O_4773,N_49807,N_49742);
xnor UO_4774 (O_4774,N_49798,N_49516);
nor UO_4775 (O_4775,N_49502,N_49537);
nor UO_4776 (O_4776,N_49639,N_49540);
nor UO_4777 (O_4777,N_49514,N_49930);
nand UO_4778 (O_4778,N_49841,N_49559);
and UO_4779 (O_4779,N_49838,N_49677);
nor UO_4780 (O_4780,N_49547,N_49909);
and UO_4781 (O_4781,N_49897,N_49741);
and UO_4782 (O_4782,N_49845,N_49646);
nand UO_4783 (O_4783,N_49801,N_49887);
and UO_4784 (O_4784,N_49883,N_49644);
and UO_4785 (O_4785,N_49756,N_49513);
or UO_4786 (O_4786,N_49726,N_49646);
or UO_4787 (O_4787,N_49915,N_49884);
and UO_4788 (O_4788,N_49666,N_49941);
or UO_4789 (O_4789,N_49919,N_49576);
or UO_4790 (O_4790,N_49847,N_49641);
xor UO_4791 (O_4791,N_49511,N_49674);
nand UO_4792 (O_4792,N_49508,N_49875);
xnor UO_4793 (O_4793,N_49986,N_49979);
nand UO_4794 (O_4794,N_49858,N_49925);
or UO_4795 (O_4795,N_49927,N_49511);
nand UO_4796 (O_4796,N_49584,N_49681);
nand UO_4797 (O_4797,N_49712,N_49854);
nor UO_4798 (O_4798,N_49504,N_49647);
and UO_4799 (O_4799,N_49942,N_49696);
nor UO_4800 (O_4800,N_49708,N_49561);
nor UO_4801 (O_4801,N_49992,N_49548);
or UO_4802 (O_4802,N_49603,N_49537);
nand UO_4803 (O_4803,N_49811,N_49699);
nor UO_4804 (O_4804,N_49688,N_49906);
or UO_4805 (O_4805,N_49859,N_49747);
xnor UO_4806 (O_4806,N_49536,N_49781);
and UO_4807 (O_4807,N_49793,N_49557);
or UO_4808 (O_4808,N_49540,N_49669);
nor UO_4809 (O_4809,N_49584,N_49964);
or UO_4810 (O_4810,N_49992,N_49750);
nor UO_4811 (O_4811,N_49749,N_49870);
xnor UO_4812 (O_4812,N_49578,N_49630);
and UO_4813 (O_4813,N_49745,N_49848);
nand UO_4814 (O_4814,N_49634,N_49772);
or UO_4815 (O_4815,N_49500,N_49675);
or UO_4816 (O_4816,N_49763,N_49782);
nor UO_4817 (O_4817,N_49695,N_49921);
xnor UO_4818 (O_4818,N_49528,N_49740);
nor UO_4819 (O_4819,N_49644,N_49650);
nand UO_4820 (O_4820,N_49566,N_49574);
xnor UO_4821 (O_4821,N_49684,N_49504);
nand UO_4822 (O_4822,N_49509,N_49991);
or UO_4823 (O_4823,N_49536,N_49901);
nand UO_4824 (O_4824,N_49768,N_49856);
xor UO_4825 (O_4825,N_49599,N_49864);
or UO_4826 (O_4826,N_49583,N_49663);
xnor UO_4827 (O_4827,N_49989,N_49700);
xnor UO_4828 (O_4828,N_49599,N_49772);
nand UO_4829 (O_4829,N_49937,N_49664);
nand UO_4830 (O_4830,N_49807,N_49927);
or UO_4831 (O_4831,N_49634,N_49988);
xor UO_4832 (O_4832,N_49929,N_49559);
nand UO_4833 (O_4833,N_49717,N_49952);
xor UO_4834 (O_4834,N_49838,N_49762);
nand UO_4835 (O_4835,N_49727,N_49866);
nand UO_4836 (O_4836,N_49986,N_49513);
or UO_4837 (O_4837,N_49886,N_49587);
xnor UO_4838 (O_4838,N_49800,N_49665);
nand UO_4839 (O_4839,N_49773,N_49976);
and UO_4840 (O_4840,N_49754,N_49866);
nand UO_4841 (O_4841,N_49719,N_49831);
xnor UO_4842 (O_4842,N_49678,N_49793);
and UO_4843 (O_4843,N_49979,N_49671);
and UO_4844 (O_4844,N_49588,N_49899);
nor UO_4845 (O_4845,N_49712,N_49525);
and UO_4846 (O_4846,N_49970,N_49966);
xnor UO_4847 (O_4847,N_49989,N_49775);
and UO_4848 (O_4848,N_49539,N_49785);
nor UO_4849 (O_4849,N_49898,N_49535);
nor UO_4850 (O_4850,N_49777,N_49505);
nor UO_4851 (O_4851,N_49898,N_49587);
xor UO_4852 (O_4852,N_49579,N_49853);
nand UO_4853 (O_4853,N_49703,N_49873);
nor UO_4854 (O_4854,N_49972,N_49582);
nor UO_4855 (O_4855,N_49817,N_49677);
and UO_4856 (O_4856,N_49822,N_49884);
or UO_4857 (O_4857,N_49992,N_49586);
nand UO_4858 (O_4858,N_49647,N_49854);
nor UO_4859 (O_4859,N_49700,N_49595);
and UO_4860 (O_4860,N_49535,N_49681);
nor UO_4861 (O_4861,N_49820,N_49918);
and UO_4862 (O_4862,N_49550,N_49683);
nand UO_4863 (O_4863,N_49842,N_49686);
or UO_4864 (O_4864,N_49612,N_49972);
nor UO_4865 (O_4865,N_49984,N_49583);
and UO_4866 (O_4866,N_49813,N_49865);
nand UO_4867 (O_4867,N_49693,N_49906);
or UO_4868 (O_4868,N_49899,N_49660);
and UO_4869 (O_4869,N_49823,N_49659);
nand UO_4870 (O_4870,N_49669,N_49727);
or UO_4871 (O_4871,N_49526,N_49530);
xnor UO_4872 (O_4872,N_49814,N_49702);
and UO_4873 (O_4873,N_49529,N_49676);
xor UO_4874 (O_4874,N_49820,N_49676);
nor UO_4875 (O_4875,N_49965,N_49736);
xor UO_4876 (O_4876,N_49777,N_49749);
or UO_4877 (O_4877,N_49541,N_49835);
or UO_4878 (O_4878,N_49770,N_49645);
nor UO_4879 (O_4879,N_49718,N_49735);
and UO_4880 (O_4880,N_49927,N_49613);
nor UO_4881 (O_4881,N_49834,N_49890);
nor UO_4882 (O_4882,N_49913,N_49982);
or UO_4883 (O_4883,N_49829,N_49754);
or UO_4884 (O_4884,N_49984,N_49551);
nand UO_4885 (O_4885,N_49690,N_49907);
xor UO_4886 (O_4886,N_49527,N_49977);
and UO_4887 (O_4887,N_49750,N_49735);
nor UO_4888 (O_4888,N_49921,N_49748);
and UO_4889 (O_4889,N_49655,N_49994);
nand UO_4890 (O_4890,N_49965,N_49977);
xnor UO_4891 (O_4891,N_49802,N_49913);
nor UO_4892 (O_4892,N_49528,N_49793);
nand UO_4893 (O_4893,N_49958,N_49658);
or UO_4894 (O_4894,N_49590,N_49709);
nand UO_4895 (O_4895,N_49882,N_49634);
nand UO_4896 (O_4896,N_49788,N_49768);
xor UO_4897 (O_4897,N_49712,N_49562);
or UO_4898 (O_4898,N_49679,N_49957);
or UO_4899 (O_4899,N_49932,N_49847);
nor UO_4900 (O_4900,N_49728,N_49911);
nand UO_4901 (O_4901,N_49596,N_49700);
and UO_4902 (O_4902,N_49687,N_49591);
or UO_4903 (O_4903,N_49593,N_49607);
nor UO_4904 (O_4904,N_49572,N_49922);
nor UO_4905 (O_4905,N_49900,N_49970);
or UO_4906 (O_4906,N_49861,N_49797);
xor UO_4907 (O_4907,N_49629,N_49516);
and UO_4908 (O_4908,N_49514,N_49533);
nand UO_4909 (O_4909,N_49631,N_49596);
xor UO_4910 (O_4910,N_49602,N_49732);
xor UO_4911 (O_4911,N_49512,N_49903);
xnor UO_4912 (O_4912,N_49583,N_49514);
xnor UO_4913 (O_4913,N_49997,N_49584);
nand UO_4914 (O_4914,N_49788,N_49911);
or UO_4915 (O_4915,N_49947,N_49943);
and UO_4916 (O_4916,N_49967,N_49732);
or UO_4917 (O_4917,N_49615,N_49898);
and UO_4918 (O_4918,N_49753,N_49846);
nand UO_4919 (O_4919,N_49723,N_49735);
nand UO_4920 (O_4920,N_49647,N_49755);
and UO_4921 (O_4921,N_49819,N_49888);
nor UO_4922 (O_4922,N_49964,N_49641);
or UO_4923 (O_4923,N_49674,N_49759);
and UO_4924 (O_4924,N_49703,N_49647);
xor UO_4925 (O_4925,N_49928,N_49763);
nor UO_4926 (O_4926,N_49837,N_49904);
nor UO_4927 (O_4927,N_49502,N_49609);
or UO_4928 (O_4928,N_49533,N_49928);
nand UO_4929 (O_4929,N_49627,N_49729);
nor UO_4930 (O_4930,N_49814,N_49880);
or UO_4931 (O_4931,N_49942,N_49898);
nor UO_4932 (O_4932,N_49754,N_49930);
nor UO_4933 (O_4933,N_49920,N_49613);
nor UO_4934 (O_4934,N_49520,N_49671);
nor UO_4935 (O_4935,N_49836,N_49774);
xor UO_4936 (O_4936,N_49645,N_49983);
nand UO_4937 (O_4937,N_49952,N_49551);
and UO_4938 (O_4938,N_49665,N_49539);
nor UO_4939 (O_4939,N_49688,N_49696);
xor UO_4940 (O_4940,N_49654,N_49901);
xor UO_4941 (O_4941,N_49904,N_49947);
xnor UO_4942 (O_4942,N_49502,N_49645);
or UO_4943 (O_4943,N_49807,N_49520);
or UO_4944 (O_4944,N_49973,N_49819);
nand UO_4945 (O_4945,N_49614,N_49648);
or UO_4946 (O_4946,N_49930,N_49502);
nand UO_4947 (O_4947,N_49639,N_49726);
nand UO_4948 (O_4948,N_49864,N_49722);
or UO_4949 (O_4949,N_49551,N_49747);
and UO_4950 (O_4950,N_49854,N_49991);
nand UO_4951 (O_4951,N_49546,N_49869);
or UO_4952 (O_4952,N_49596,N_49942);
or UO_4953 (O_4953,N_49722,N_49567);
nand UO_4954 (O_4954,N_49917,N_49819);
nor UO_4955 (O_4955,N_49839,N_49829);
nor UO_4956 (O_4956,N_49785,N_49701);
and UO_4957 (O_4957,N_49662,N_49824);
nand UO_4958 (O_4958,N_49744,N_49743);
xnor UO_4959 (O_4959,N_49541,N_49506);
nor UO_4960 (O_4960,N_49646,N_49776);
or UO_4961 (O_4961,N_49606,N_49988);
and UO_4962 (O_4962,N_49945,N_49705);
xnor UO_4963 (O_4963,N_49524,N_49623);
or UO_4964 (O_4964,N_49522,N_49515);
xnor UO_4965 (O_4965,N_49605,N_49643);
nor UO_4966 (O_4966,N_49860,N_49826);
xnor UO_4967 (O_4967,N_49525,N_49710);
xnor UO_4968 (O_4968,N_49638,N_49574);
nand UO_4969 (O_4969,N_49913,N_49501);
and UO_4970 (O_4970,N_49988,N_49578);
xnor UO_4971 (O_4971,N_49716,N_49695);
nor UO_4972 (O_4972,N_49759,N_49827);
nand UO_4973 (O_4973,N_49938,N_49905);
xnor UO_4974 (O_4974,N_49961,N_49809);
nand UO_4975 (O_4975,N_49719,N_49703);
nor UO_4976 (O_4976,N_49768,N_49866);
and UO_4977 (O_4977,N_49913,N_49879);
nor UO_4978 (O_4978,N_49886,N_49866);
and UO_4979 (O_4979,N_49607,N_49579);
nor UO_4980 (O_4980,N_49750,N_49803);
or UO_4981 (O_4981,N_49649,N_49632);
and UO_4982 (O_4982,N_49787,N_49741);
nand UO_4983 (O_4983,N_49819,N_49589);
and UO_4984 (O_4984,N_49866,N_49823);
xor UO_4985 (O_4985,N_49770,N_49899);
and UO_4986 (O_4986,N_49551,N_49940);
nand UO_4987 (O_4987,N_49816,N_49915);
nand UO_4988 (O_4988,N_49797,N_49717);
and UO_4989 (O_4989,N_49936,N_49617);
nor UO_4990 (O_4990,N_49567,N_49843);
and UO_4991 (O_4991,N_49840,N_49789);
xor UO_4992 (O_4992,N_49626,N_49693);
nand UO_4993 (O_4993,N_49587,N_49824);
nor UO_4994 (O_4994,N_49628,N_49719);
xor UO_4995 (O_4995,N_49734,N_49523);
xnor UO_4996 (O_4996,N_49622,N_49674);
nand UO_4997 (O_4997,N_49716,N_49698);
nor UO_4998 (O_4998,N_49606,N_49677);
and UO_4999 (O_4999,N_49795,N_49757);
endmodule