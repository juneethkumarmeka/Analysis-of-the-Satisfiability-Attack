module basic_2500_25000_3000_4_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18841,N_18842,N_18843,N_18844,N_18845,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19098,N_19099,N_19100,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19189,N_19190,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19201,N_19202,N_19203,N_19204,N_19205,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19317,N_19318,N_19319,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19389,N_19390,N_19391,N_19392,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19634,N_19635,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19655,N_19656,N_19657,N_19658,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19760,N_19761,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20334,N_20335,N_20336,N_20337,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20527,N_20529,N_20530,N_20531,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20926,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21049,N_21050,N_21051,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21091,N_21092,N_21093,N_21094,N_21095,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21105,N_21106,N_21107,N_21108,N_21109,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21140,N_21141,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21217,N_21218,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21324,N_21325,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21802,N_21803,N_21804,N_21805,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22188,N_22189,N_22190,N_22191,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22230,N_22231,N_22232,N_22233,N_22234,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22277,N_22278,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22296,N_22297,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22505,N_22506,N_22507,N_22508,N_22509,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22548,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22565,N_22566,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22731,N_22732,N_22733,N_22734,N_22735,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22853,N_22854,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22899,N_22900,N_22901,N_22902,N_22903,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23001,N_23002,N_23003,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23284,N_23285,N_23286,N_23287,N_23288,N_23290,N_23291,N_23292,N_23293,N_23294,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23446,N_23447,N_23448,N_23450,N_23451,N_23452,N_23453,N_23454,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23463,N_23464,N_23465,N_23466,N_23467,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23522,N_23523,N_23524,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23548,N_23549,N_23550,N_23551,N_23552,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23575,N_23577,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24174,N_24175,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24184,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24411,N_24412,N_24414,N_24415,N_24416,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24931,N_24932,N_24934,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1216,In_2032);
or U1 (N_1,In_1465,In_1239);
nor U2 (N_2,In_2158,In_466);
and U3 (N_3,In_90,In_2391);
nand U4 (N_4,In_2442,In_2459);
and U5 (N_5,In_2084,In_694);
xnor U6 (N_6,In_1318,In_106);
and U7 (N_7,In_210,In_1417);
nand U8 (N_8,In_1549,In_1930);
xor U9 (N_9,In_2300,In_871);
nand U10 (N_10,In_2148,In_2468);
or U11 (N_11,In_224,In_617);
nor U12 (N_12,In_362,In_887);
and U13 (N_13,In_1160,In_1184);
nand U14 (N_14,In_260,In_101);
xor U15 (N_15,In_411,In_1776);
xnor U16 (N_16,In_2106,In_478);
nand U17 (N_17,In_1048,In_2423);
nand U18 (N_18,In_707,In_215);
nor U19 (N_19,In_288,In_229);
or U20 (N_20,In_304,In_451);
and U21 (N_21,In_636,In_666);
nor U22 (N_22,In_2050,In_510);
xnor U23 (N_23,In_345,In_1326);
nor U24 (N_24,In_113,In_1371);
nand U25 (N_25,In_1947,In_2455);
nand U26 (N_26,In_1992,In_1446);
nor U27 (N_27,In_2034,In_2002);
and U28 (N_28,In_2412,In_2046);
and U29 (N_29,In_401,In_1306);
and U30 (N_30,In_2233,In_2011);
nor U31 (N_31,In_1846,In_675);
or U32 (N_32,In_2260,In_2483);
nor U33 (N_33,In_2219,In_230);
nand U34 (N_34,In_1673,In_927);
xor U35 (N_35,In_1951,In_1849);
xnor U36 (N_36,In_1166,In_784);
nor U37 (N_37,In_1079,In_1000);
nand U38 (N_38,In_2301,In_1340);
nand U39 (N_39,In_1696,In_1090);
nand U40 (N_40,In_296,In_2013);
nor U41 (N_41,In_480,In_2196);
xnor U42 (N_42,In_269,In_1124);
nand U43 (N_43,In_1966,In_1368);
xnor U44 (N_44,In_1989,In_1256);
or U45 (N_45,In_290,In_2220);
nor U46 (N_46,In_2165,In_657);
nand U47 (N_47,In_1045,In_68);
and U48 (N_48,In_562,In_1134);
xnor U49 (N_49,In_356,In_1848);
xor U50 (N_50,In_1301,In_1407);
nor U51 (N_51,In_2316,In_531);
or U52 (N_52,In_1060,In_1578);
xnor U53 (N_53,In_844,In_365);
or U54 (N_54,In_1390,In_1743);
or U55 (N_55,In_2144,In_660);
xnor U56 (N_56,In_344,In_1603);
and U57 (N_57,In_2258,In_441);
xnor U58 (N_58,In_1171,In_1935);
nand U59 (N_59,In_1191,In_1772);
nor U60 (N_60,In_1194,In_997);
nand U61 (N_61,In_736,In_1339);
or U62 (N_62,In_1539,In_1029);
and U63 (N_63,In_541,In_1796);
nor U64 (N_64,In_1660,In_1);
and U65 (N_65,In_472,In_721);
and U66 (N_66,In_1058,In_2454);
and U67 (N_67,In_158,In_816);
nor U68 (N_68,In_543,In_157);
nor U69 (N_69,In_1033,In_397);
or U70 (N_70,In_1808,In_929);
xor U71 (N_71,In_2147,In_708);
and U72 (N_72,In_581,In_806);
nand U73 (N_73,In_900,In_61);
and U74 (N_74,In_991,In_430);
xor U75 (N_75,In_628,In_2397);
xnor U76 (N_76,In_670,In_257);
nand U77 (N_77,In_1290,In_2066);
nor U78 (N_78,In_563,In_847);
and U79 (N_79,In_1592,In_203);
nor U80 (N_80,In_897,In_2246);
or U81 (N_81,In_1584,In_240);
and U82 (N_82,In_1746,In_1019);
nor U83 (N_83,In_2346,In_1731);
xor U84 (N_84,In_2272,In_555);
and U85 (N_85,In_464,In_647);
and U86 (N_86,In_389,In_2323);
and U87 (N_87,In_2404,In_1934);
or U88 (N_88,In_457,In_1392);
nand U89 (N_89,In_593,In_1460);
nor U90 (N_90,In_2313,In_783);
nor U91 (N_91,In_1401,In_881);
nor U92 (N_92,In_741,In_195);
nand U93 (N_93,In_925,In_993);
or U94 (N_94,In_1593,In_1459);
nor U95 (N_95,In_201,In_2443);
nand U96 (N_96,In_650,In_1745);
and U97 (N_97,In_726,In_1346);
and U98 (N_98,In_1273,In_710);
or U99 (N_99,In_942,In_1978);
xor U100 (N_100,In_1081,In_974);
nor U101 (N_101,In_1697,In_2189);
nor U102 (N_102,In_1840,In_2488);
xor U103 (N_103,In_2164,In_2109);
nand U104 (N_104,In_2049,In_1604);
and U105 (N_105,In_970,In_69);
and U106 (N_106,In_1172,In_2067);
nand U107 (N_107,In_1856,In_1872);
nand U108 (N_108,In_1137,In_1320);
and U109 (N_109,In_1608,In_703);
and U110 (N_110,In_637,In_2324);
nor U111 (N_111,In_55,In_2010);
nand U112 (N_112,In_2469,In_2122);
nor U113 (N_113,In_2195,In_718);
nor U114 (N_114,In_1933,In_988);
xor U115 (N_115,In_1217,In_33);
nor U116 (N_116,In_360,In_771);
or U117 (N_117,In_74,In_1083);
and U118 (N_118,In_91,In_398);
and U119 (N_119,In_837,In_437);
nand U120 (N_120,In_870,In_1457);
xnor U121 (N_121,In_461,In_1244);
and U122 (N_122,In_1876,In_2386);
nor U123 (N_123,In_403,In_2473);
nor U124 (N_124,In_1990,In_1971);
or U125 (N_125,In_1068,In_1338);
xor U126 (N_126,In_273,In_2026);
nand U127 (N_127,In_0,In_627);
nand U128 (N_128,In_1558,In_279);
xnor U129 (N_129,In_420,In_616);
or U130 (N_130,In_1901,In_2353);
nand U131 (N_131,In_1694,In_323);
or U132 (N_132,In_455,In_1471);
or U133 (N_133,In_2270,In_264);
xnor U134 (N_134,In_1577,In_1730);
nand U135 (N_135,In_1158,In_213);
or U136 (N_136,In_1544,In_1499);
or U137 (N_137,In_2078,In_1268);
xnor U138 (N_138,In_1798,In_937);
nor U139 (N_139,In_1468,In_1777);
nand U140 (N_140,In_242,In_504);
and U141 (N_141,In_1429,In_2019);
xnor U142 (N_142,In_757,In_1823);
and U143 (N_143,In_313,In_1316);
and U144 (N_144,In_2486,In_1122);
nand U145 (N_145,In_978,In_1713);
nand U146 (N_146,In_2135,In_1051);
or U147 (N_147,In_262,In_1467);
and U148 (N_148,In_2410,In_1859);
or U149 (N_149,In_54,In_948);
nand U150 (N_150,In_891,In_1646);
and U151 (N_151,In_855,In_41);
nor U152 (N_152,In_1939,In_184);
nor U153 (N_153,In_1960,In_1587);
nand U154 (N_154,In_888,In_795);
or U155 (N_155,In_1212,In_1103);
and U156 (N_156,In_1485,In_1975);
nor U157 (N_157,In_1118,In_340);
xnor U158 (N_158,In_1864,In_286);
or U159 (N_159,In_1517,In_1758);
xor U160 (N_160,In_2250,In_2123);
xnor U161 (N_161,In_223,In_2274);
xor U162 (N_162,In_2361,In_1890);
and U163 (N_163,In_1594,In_1638);
nor U164 (N_164,In_959,In_1794);
and U165 (N_165,In_2341,In_1585);
nand U166 (N_166,In_2017,In_2303);
or U167 (N_167,In_532,In_120);
and U168 (N_168,In_2108,In_1159);
or U169 (N_169,In_1759,In_2467);
nand U170 (N_170,In_231,In_2177);
or U171 (N_171,In_1508,In_943);
or U172 (N_172,In_310,In_1204);
or U173 (N_173,In_1169,In_898);
nand U174 (N_174,In_695,In_1970);
xor U175 (N_175,In_2045,In_1658);
nand U176 (N_176,In_59,In_1748);
nand U177 (N_177,In_2161,In_1546);
xnor U178 (N_178,In_638,In_1432);
or U179 (N_179,In_646,In_2208);
nor U180 (N_180,In_475,In_921);
nor U181 (N_181,In_1997,In_2181);
and U182 (N_182,In_216,In_729);
nand U183 (N_183,In_1855,In_1061);
nor U184 (N_184,In_178,In_1783);
and U185 (N_185,In_957,In_2440);
xnor U186 (N_186,In_2001,In_1464);
and U187 (N_187,In_517,In_2381);
xor U188 (N_188,In_1961,In_727);
nand U189 (N_189,In_2298,In_515);
xor U190 (N_190,In_905,In_1909);
xor U191 (N_191,In_1055,In_2359);
and U192 (N_192,In_756,In_358);
nor U193 (N_193,In_526,In_348);
xnor U194 (N_194,In_573,In_1096);
nor U195 (N_195,In_984,In_94);
nor U196 (N_196,In_1703,In_2096);
xnor U197 (N_197,In_462,In_1580);
nand U198 (N_198,In_1599,In_1622);
nand U199 (N_199,In_2040,In_1001);
xor U200 (N_200,In_873,In_141);
and U201 (N_201,In_2,In_326);
nor U202 (N_202,In_508,In_1800);
and U203 (N_203,In_843,In_1867);
and U204 (N_204,In_1568,In_1722);
and U205 (N_205,In_1132,In_402);
nand U206 (N_206,In_2243,In_1949);
nor U207 (N_207,In_2043,In_2191);
nand U208 (N_208,In_1728,In_1811);
nand U209 (N_209,In_301,In_2024);
or U210 (N_210,In_2415,In_2432);
and U211 (N_211,In_2118,In_93);
or U212 (N_212,In_1538,In_1157);
nand U213 (N_213,In_1636,In_625);
nand U214 (N_214,In_261,In_1202);
nor U215 (N_215,In_1190,In_52);
xor U216 (N_216,In_388,In_412);
nor U217 (N_217,In_2490,In_1507);
and U218 (N_218,In_2439,In_357);
and U219 (N_219,In_2254,In_1140);
nand U220 (N_220,In_2349,In_1860);
nand U221 (N_221,In_1315,In_2041);
xor U222 (N_222,In_931,In_2428);
nand U223 (N_223,In_1297,In_172);
nor U224 (N_224,In_263,In_8);
nor U225 (N_225,In_1224,In_1742);
and U226 (N_226,In_546,In_1751);
and U227 (N_227,In_26,In_740);
and U228 (N_228,In_2087,In_1450);
nand U229 (N_229,In_271,In_2447);
nor U230 (N_230,In_2222,In_1600);
nor U231 (N_231,In_418,In_1550);
or U232 (N_232,In_603,In_2248);
or U233 (N_233,In_697,In_1152);
nor U234 (N_234,In_2103,In_2042);
xor U235 (N_235,In_2456,In_2344);
nand U236 (N_236,In_2425,In_1677);
or U237 (N_237,In_1312,In_1080);
xor U238 (N_238,In_64,In_1192);
and U239 (N_239,In_31,In_337);
nor U240 (N_240,In_1006,In_1929);
nand U241 (N_241,In_1705,In_1814);
and U242 (N_242,In_2097,In_176);
and U243 (N_243,In_209,In_511);
nor U244 (N_244,In_51,In_1619);
xnor U245 (N_245,In_2477,In_714);
nor U246 (N_246,In_1861,In_454);
and U247 (N_247,In_1489,In_1112);
nor U248 (N_248,In_706,In_665);
xor U249 (N_249,In_965,In_1040);
xnor U250 (N_250,In_1111,In_1084);
nand U251 (N_251,In_2230,In_228);
nand U252 (N_252,In_19,In_2056);
nand U253 (N_253,In_1591,In_249);
xnor U254 (N_254,In_2069,In_1945);
nand U255 (N_255,In_1440,In_2378);
xor U256 (N_256,In_1335,In_1691);
nor U257 (N_257,In_2168,In_440);
or U258 (N_258,In_2227,In_1780);
xnor U259 (N_259,In_309,In_2480);
nand U260 (N_260,In_2229,In_1551);
or U261 (N_261,In_234,In_731);
nor U262 (N_262,In_482,In_2400);
nand U263 (N_263,In_2036,In_2256);
and U264 (N_264,In_1667,In_1139);
or U265 (N_265,In_2235,In_768);
and U266 (N_266,In_2142,In_2116);
nand U267 (N_267,In_701,In_1908);
xnor U268 (N_268,In_1104,In_2487);
xor U269 (N_269,In_1784,In_1427);
xor U270 (N_270,In_2498,In_643);
nor U271 (N_271,In_1428,In_305);
nand U272 (N_272,In_624,In_587);
nor U273 (N_273,In_88,In_1125);
xnor U274 (N_274,In_2294,In_933);
nor U275 (N_275,In_85,In_27);
xnor U276 (N_276,In_2101,In_1706);
nand U277 (N_277,In_2427,In_2336);
and U278 (N_278,In_2188,In_471);
nor U279 (N_279,In_1889,In_2362);
and U280 (N_280,In_963,In_1113);
and U281 (N_281,In_1250,In_2285);
and U282 (N_282,In_2099,In_1816);
xnor U283 (N_283,In_489,In_932);
nand U284 (N_284,In_6,In_488);
or U285 (N_285,In_2242,In_1526);
nand U286 (N_286,In_376,In_1795);
and U287 (N_287,In_1133,In_1458);
or U288 (N_288,In_422,In_1376);
nor U289 (N_289,In_2281,In_1410);
and U290 (N_290,In_792,In_1209);
xor U291 (N_291,In_522,In_686);
and U292 (N_292,In_503,In_287);
or U293 (N_293,In_1053,In_552);
and U294 (N_294,In_1530,In_253);
and U295 (N_295,In_385,In_1529);
nor U296 (N_296,In_2197,In_1279);
xnor U297 (N_297,In_1294,In_2149);
and U298 (N_298,In_1560,In_429);
xor U299 (N_299,In_542,In_1813);
xnor U300 (N_300,In_513,In_1422);
xnor U301 (N_301,In_1399,In_312);
nor U302 (N_302,In_558,In_947);
xor U303 (N_303,In_1886,In_569);
nand U304 (N_304,In_191,In_1142);
nand U305 (N_305,In_519,In_571);
xnor U306 (N_306,In_1105,In_977);
xor U307 (N_307,In_1498,In_1976);
nand U308 (N_308,In_1547,In_1518);
nor U309 (N_309,In_2186,In_1559);
and U310 (N_310,In_16,In_319);
nand U311 (N_311,In_1519,In_208);
xnor U312 (N_312,In_2210,In_270);
or U313 (N_313,In_2139,In_1298);
nand U314 (N_314,In_1482,In_967);
and U315 (N_315,In_754,In_1779);
xor U316 (N_316,In_834,In_1411);
nor U317 (N_317,In_2051,In_1156);
nor U318 (N_318,In_1481,In_1452);
nor U319 (N_319,In_1097,In_656);
xnor U320 (N_320,In_2350,In_372);
nor U321 (N_321,In_1162,In_2499);
xor U322 (N_322,In_421,In_1302);
xor U323 (N_323,In_2299,In_621);
or U324 (N_324,In_996,In_415);
nand U325 (N_325,In_1072,In_893);
or U326 (N_326,In_1927,In_419);
nand U327 (N_327,In_1605,In_679);
xnor U328 (N_328,In_274,In_1623);
or U329 (N_329,In_1914,In_177);
or U330 (N_330,In_1803,In_527);
xor U331 (N_331,In_777,In_1222);
and U332 (N_332,In_1375,In_1625);
or U333 (N_333,In_605,In_610);
xnor U334 (N_334,In_1806,In_556);
xor U335 (N_335,In_2493,In_1098);
nand U336 (N_336,In_1299,In_880);
xnor U337 (N_337,In_119,In_2284);
or U338 (N_338,In_1838,In_493);
or U339 (N_339,In_2004,In_1437);
xor U340 (N_340,In_2022,In_1282);
nor U341 (N_341,In_1187,In_2224);
nand U342 (N_342,In_1420,In_769);
or U343 (N_343,In_2268,In_612);
nor U344 (N_344,In_1237,In_1366);
and U345 (N_345,In_1695,In_244);
or U346 (N_346,In_171,In_790);
xor U347 (N_347,In_112,In_1477);
or U348 (N_348,In_565,In_2044);
xor U349 (N_349,In_2436,In_2200);
nor U350 (N_350,In_1893,In_67);
and U351 (N_351,In_416,In_709);
and U352 (N_352,In_248,In_1369);
xnor U353 (N_353,In_1289,In_575);
xnor U354 (N_354,In_63,In_2420);
nand U355 (N_355,In_717,In_374);
nor U356 (N_356,In_1117,In_1403);
nor U357 (N_357,In_874,In_1750);
or U358 (N_358,In_1617,In_1851);
xor U359 (N_359,In_1324,In_153);
nor U360 (N_360,In_2183,In_1077);
and U361 (N_361,In_320,In_352);
nor U362 (N_362,In_704,In_1520);
nor U363 (N_363,In_425,In_131);
xnor U364 (N_364,In_1955,In_1881);
nand U365 (N_365,In_2283,In_225);
and U366 (N_366,In_2090,In_2431);
nor U367 (N_367,In_1425,In_1511);
or U368 (N_368,In_1664,In_2356);
or U369 (N_369,In_114,In_1092);
nand U370 (N_370,In_2430,In_144);
nor U371 (N_371,In_165,In_2365);
or U372 (N_372,In_767,In_1915);
nand U373 (N_373,In_456,In_826);
or U374 (N_374,In_2405,In_904);
or U375 (N_375,In_1356,In_139);
or U376 (N_376,In_2039,In_682);
xor U377 (N_377,In_1774,In_1321);
nor U378 (N_378,In_2184,In_2262);
nor U379 (N_379,In_600,In_276);
nor U380 (N_380,In_1136,In_431);
or U381 (N_381,In_1639,In_739);
and U382 (N_382,In_163,In_901);
xnor U383 (N_383,In_1649,In_200);
nand U384 (N_384,In_1678,In_1255);
nand U385 (N_385,In_1662,In_433);
nand U386 (N_386,In_1702,In_370);
nand U387 (N_387,In_291,In_659);
nor U388 (N_388,In_1030,In_86);
or U389 (N_389,In_2394,In_2472);
and U390 (N_390,In_1987,In_1887);
and U391 (N_391,In_2009,In_1671);
nand U392 (N_392,In_557,In_1141);
or U393 (N_393,In_1516,In_1114);
or U394 (N_394,In_50,In_1449);
xnor U395 (N_395,In_2126,In_1101);
or U396 (N_396,In_1296,In_835);
xor U397 (N_397,In_380,In_794);
and U398 (N_398,In_126,In_1314);
xnor U399 (N_399,In_878,In_378);
nand U400 (N_400,In_1189,In_1896);
nor U401 (N_401,In_1049,In_1488);
or U402 (N_402,In_1404,In_1229);
nand U403 (N_403,In_1210,In_413);
or U404 (N_404,In_486,In_1741);
nand U405 (N_405,In_2311,In_1441);
nand U406 (N_406,In_485,In_586);
or U407 (N_407,In_1534,In_2240);
nand U408 (N_408,In_2204,In_956);
and U409 (N_409,In_117,In_1337);
or U410 (N_410,In_324,In_805);
nand U411 (N_411,In_2411,In_379);
or U412 (N_412,In_692,In_1344);
nor U413 (N_413,In_2309,In_1762);
nand U414 (N_414,In_1888,In_1514);
and U415 (N_415,In_1963,In_550);
nand U416 (N_416,In_84,In_175);
nor U417 (N_417,In_382,In_1198);
and U418 (N_418,In_917,In_2155);
xor U419 (N_419,In_1261,In_2291);
or U420 (N_420,In_481,In_48);
xnor U421 (N_421,In_2271,In_1756);
xnor U422 (N_422,In_1657,In_47);
and U423 (N_423,In_672,In_2073);
nor U424 (N_424,In_1680,In_1904);
xor U425 (N_425,In_763,In_1793);
or U426 (N_426,In_589,In_236);
and U427 (N_427,In_65,In_1435);
xnor U428 (N_428,In_987,In_369);
nor U429 (N_429,In_470,In_1692);
xor U430 (N_430,In_658,In_151);
nand U431 (N_431,In_1388,In_2286);
or U432 (N_432,In_145,In_2471);
xnor U433 (N_433,In_1699,In_23);
nand U434 (N_434,In_1350,In_1193);
nor U435 (N_435,In_1616,In_393);
or U436 (N_436,In_1845,In_867);
xor U437 (N_437,In_934,In_1773);
nand U438 (N_438,In_1292,In_44);
nor U439 (N_439,In_469,In_1334);
xor U440 (N_440,In_1964,In_212);
nand U441 (N_441,In_1554,In_712);
and U442 (N_442,In_1698,In_992);
nor U443 (N_443,In_443,In_428);
and U444 (N_444,In_1004,In_1629);
xor U445 (N_445,In_1223,In_1866);
and U446 (N_446,In_2063,In_940);
nand U447 (N_447,In_747,In_160);
xor U448 (N_448,In_328,In_1329);
xnor U449 (N_449,In_1313,In_1494);
nor U450 (N_450,In_1822,In_1847);
and U451 (N_451,In_2020,In_452);
and U452 (N_452,In_2251,In_190);
nor U453 (N_453,In_908,In_2190);
or U454 (N_454,In_2216,In_9);
or U455 (N_455,In_725,In_281);
xnor U456 (N_456,In_1850,In_2061);
nand U457 (N_457,In_1057,In_1684);
nor U458 (N_458,In_671,In_1891);
or U459 (N_459,In_2185,In_2453);
and U460 (N_460,In_2363,In_2259);
xnor U461 (N_461,In_207,In_698);
xor U462 (N_462,In_2390,In_2322);
or U463 (N_463,In_235,In_2249);
nand U464 (N_464,In_1778,In_892);
xnor U465 (N_465,In_1601,In_1642);
and U466 (N_466,In_2055,In_1956);
xnor U467 (N_467,In_926,In_1597);
nor U468 (N_468,In_990,In_185);
and U469 (N_469,In_645,In_1512);
nor U470 (N_470,In_596,In_170);
nor U471 (N_471,In_1542,In_1821);
xor U472 (N_472,In_1870,In_1039);
nor U473 (N_473,In_100,In_108);
xnor U474 (N_474,In_1269,In_1123);
nor U475 (N_475,In_394,In_2290);
xor U476 (N_476,In_1386,In_341);
or U477 (N_477,In_1233,In_2115);
nand U478 (N_478,In_1739,In_1274);
and U479 (N_479,In_2052,In_1023);
nor U480 (N_480,In_179,In_968);
nor U481 (N_481,In_1595,In_28);
xor U482 (N_482,In_391,In_2282);
nor U483 (N_483,In_688,In_842);
or U484 (N_484,In_140,In_1506);
nor U485 (N_485,In_1374,In_267);
nor U486 (N_486,In_1853,In_807);
or U487 (N_487,In_720,In_1034);
nor U488 (N_488,In_1760,In_136);
or U489 (N_489,In_2337,In_1775);
or U490 (N_490,In_1270,In_919);
nor U491 (N_491,In_1353,In_49);
nand U492 (N_492,In_2244,In_1852);
nand U493 (N_493,In_1247,In_1025);
nor U494 (N_494,In_1785,In_2226);
xor U495 (N_495,In_355,In_1618);
nand U496 (N_496,In_155,In_400);
nor U497 (N_497,In_2209,In_1736);
or U498 (N_498,In_66,In_829);
nor U499 (N_499,In_1065,In_1612);
or U500 (N_500,In_183,In_800);
and U501 (N_501,In_2297,In_1243);
xor U502 (N_502,In_1383,In_1303);
nand U503 (N_503,In_1687,In_1094);
nor U504 (N_504,In_1483,In_1674);
and U505 (N_505,In_128,In_2277);
xor U506 (N_506,In_474,In_1128);
and U507 (N_507,In_654,In_773);
xor U508 (N_508,In_292,In_383);
nor U509 (N_509,In_949,In_1186);
and U510 (N_510,In_1535,In_473);
nand U511 (N_511,In_2476,In_349);
xor U512 (N_512,In_591,In_752);
xor U513 (N_513,In_2402,In_864);
nor U514 (N_514,In_1836,In_241);
or U515 (N_515,In_2319,In_2288);
and U516 (N_516,In_1028,In_860);
and U517 (N_517,In_2054,In_1154);
nand U518 (N_518,In_1682,In_134);
or U519 (N_519,In_499,In_869);
nand U520 (N_520,In_1490,In_1451);
or U521 (N_521,In_1724,In_1107);
and U522 (N_522,In_1562,In_2479);
nor U523 (N_523,In_1370,In_936);
and U524 (N_524,In_1714,In_748);
and U525 (N_525,In_1579,In_2238);
and U526 (N_526,In_1589,In_2077);
xor U527 (N_527,In_2315,In_733);
nor U528 (N_528,In_295,In_883);
nand U529 (N_529,In_590,In_245);
or U530 (N_530,In_239,In_1828);
xor U531 (N_531,In_734,In_1555);
nand U532 (N_532,In_607,In_137);
nand U533 (N_533,In_1287,In_1357);
xnor U534 (N_534,In_1236,In_702);
or U535 (N_535,In_1984,In_439);
nor U536 (N_536,In_1343,In_317);
or U537 (N_537,In_1632,In_1679);
and U538 (N_538,In_1280,In_1548);
nor U539 (N_539,In_2225,In_1442);
or U540 (N_540,In_162,In_945);
xnor U541 (N_541,In_1147,In_518);
xor U542 (N_542,In_639,In_760);
xnor U543 (N_543,In_368,In_570);
xnor U544 (N_544,In_220,In_1266);
nand U545 (N_545,In_180,In_716);
xor U546 (N_546,In_2308,In_588);
and U547 (N_547,In_669,In_1923);
nand U548 (N_548,In_250,In_1565);
xnor U549 (N_549,In_1278,In_2072);
nand U550 (N_550,In_1952,In_293);
nand U551 (N_551,In_498,In_83);
nor U552 (N_552,In_1844,In_2457);
nand U553 (N_553,In_1491,In_2446);
nand U554 (N_554,In_1946,In_1932);
xor U555 (N_555,In_1718,In_1382);
xor U556 (N_556,In_548,In_1126);
or U557 (N_557,In_1982,In_308);
xnor U558 (N_558,In_159,In_2333);
or U559 (N_559,In_361,In_14);
nand U560 (N_560,In_1026,In_2112);
nor U561 (N_561,In_2162,In_1824);
nor U562 (N_562,In_2173,In_387);
or U563 (N_563,In_567,In_447);
nor U564 (N_564,In_2213,In_685);
or U565 (N_565,In_226,In_404);
nor U566 (N_566,In_2198,In_1875);
nor U567 (N_567,In_2310,In_525);
nand U568 (N_568,In_1944,In_827);
or U569 (N_569,In_2201,In_912);
nor U570 (N_570,In_2214,In_505);
nor U571 (N_571,In_761,In_227);
and U572 (N_572,In_1252,In_1950);
xor U573 (N_573,In_477,In_2279);
or U574 (N_574,In_138,In_1119);
nand U575 (N_575,In_2491,In_2232);
and U576 (N_576,In_544,In_444);
nor U577 (N_577,In_1686,In_2413);
xor U578 (N_578,In_840,In_653);
nor U579 (N_579,In_632,In_1892);
nor U580 (N_580,In_1938,In_2289);
nor U581 (N_581,In_820,In_73);
nor U582 (N_582,In_1011,In_1021);
nor U583 (N_583,In_1688,In_831);
xor U584 (N_584,In_691,In_1240);
and U585 (N_585,In_651,In_1086);
xnor U586 (N_586,In_1564,In_1740);
nand U587 (N_587,In_449,In_78);
and U588 (N_588,In_1360,In_2489);
nor U589 (N_589,In_465,In_1461);
nand U590 (N_590,In_630,In_1017);
and U591 (N_591,In_450,In_2358);
nand U592 (N_592,In_1089,In_342);
nand U593 (N_593,In_1581,In_585);
or U594 (N_594,In_1054,In_318);
and U595 (N_595,In_540,In_1630);
and U596 (N_596,In_1153,In_580);
xnor U597 (N_597,In_2005,In_673);
nand U598 (N_598,In_1525,In_1470);
nor U599 (N_599,In_1827,In_1668);
nand U600 (N_600,In_1768,In_1996);
or U601 (N_601,In_502,In_467);
or U602 (N_602,In_2150,In_2202);
or U603 (N_603,In_1424,In_2292);
or U604 (N_604,In_982,In_2461);
or U605 (N_605,In_2088,In_969);
nand U606 (N_606,In_1799,In_1993);
nor U607 (N_607,In_964,In_1138);
xor U608 (N_608,In_875,In_879);
nand U609 (N_609,In_2015,In_386);
xor U610 (N_610,In_849,In_1835);
xnor U611 (N_611,In_1251,In_2451);
xnor U612 (N_612,In_1062,In_1880);
nor U613 (N_613,In_442,In_2380);
xor U614 (N_614,In_2160,In_1531);
xor U615 (N_615,In_899,In_1145);
and U616 (N_616,In_272,In_1218);
or U617 (N_617,In_1130,In_147);
nor U618 (N_618,In_1384,In_560);
or U619 (N_619,In_1036,In_2228);
nand U620 (N_620,In_2330,In_848);
or U621 (N_621,In_604,In_1643);
nand U622 (N_622,In_1358,In_1444);
or U623 (N_623,In_2433,In_283);
nand U624 (N_624,In_719,In_2369);
nand U625 (N_625,In_196,In_2143);
nand U626 (N_626,In_746,In_24);
or U627 (N_627,In_255,In_1150);
nor U628 (N_628,In_1868,In_1100);
and U629 (N_629,In_732,In_1309);
xor U630 (N_630,In_2421,In_2038);
or U631 (N_631,In_715,In_950);
nor U632 (N_632,In_1201,In_1910);
nand U633 (N_633,In_839,In_782);
and U634 (N_634,In_1834,In_193);
xor U635 (N_635,In_1115,In_284);
and U636 (N_636,In_152,In_2125);
xnor U637 (N_637,In_2388,In_1493);
nor U638 (N_638,In_1757,In_2070);
nor U639 (N_639,In_298,In_330);
nor U640 (N_640,In_1044,In_1998);
nand U641 (N_641,In_1022,In_2326);
nor U642 (N_642,In_1765,In_1317);
nor U643 (N_643,In_1865,In_2178);
or U644 (N_644,In_1448,In_2478);
nand U645 (N_645,In_1188,In_1095);
or U646 (N_646,In_278,In_857);
or U647 (N_647,In_613,In_664);
nor U648 (N_648,In_652,In_35);
or U649 (N_649,In_1487,In_1087);
nor U650 (N_650,In_2452,In_742);
nor U651 (N_651,In_58,In_2062);
xor U652 (N_652,In_1267,In_1075);
and U653 (N_653,In_597,In_118);
nor U654 (N_654,In_1174,In_772);
and U655 (N_655,In_608,In_2231);
xor U656 (N_656,In_1527,In_920);
or U657 (N_657,In_1211,In_1895);
nand U658 (N_658,In_2304,In_266);
xnor U659 (N_659,In_259,In_2152);
nor U660 (N_660,In_2367,In_221);
nor U661 (N_661,In_1277,In_533);
nand U662 (N_662,In_1328,In_1624);
nand U663 (N_663,In_955,In_765);
nor U664 (N_664,In_1786,In_232);
or U665 (N_665,In_1108,In_1903);
xnor U666 (N_666,In_10,In_886);
nand U667 (N_667,In_406,In_830);
and U668 (N_668,In_1258,In_2221);
nand U669 (N_669,In_1099,In_2494);
nand U670 (N_670,In_1931,In_668);
nand U671 (N_671,In_1726,In_1567);
xor U672 (N_672,In_2383,In_1727);
nand U673 (N_673,In_1501,In_923);
xnor U674 (N_674,In_809,In_1264);
and U675 (N_675,In_202,In_592);
or U676 (N_676,In_1110,In_735);
nand U677 (N_677,In_22,In_1734);
or U678 (N_678,In_833,In_2360);
nand U679 (N_679,In_944,In_396);
xor U680 (N_680,In_1645,In_1685);
xnor U681 (N_681,In_2095,In_110);
xor U682 (N_682,In_238,In_346);
and U683 (N_683,In_1412,In_2253);
nand U684 (N_684,In_80,In_311);
or U685 (N_685,In_2047,In_251);
nor U686 (N_686,In_1408,In_1478);
nor U687 (N_687,In_980,In_1377);
nand U688 (N_688,In_1819,In_572);
and U689 (N_689,In_1311,In_2348);
nor U690 (N_690,In_743,In_2470);
and U691 (N_691,In_2265,In_436);
or U692 (N_692,In_2137,In_2163);
nand U693 (N_693,In_2395,In_2385);
xnor U694 (N_694,In_1532,In_1288);
nor U695 (N_695,In_812,In_549);
nor U696 (N_696,In_2157,In_1681);
and U697 (N_697,In_2334,In_1701);
nor U698 (N_698,In_2403,In_1918);
or U699 (N_699,In_2317,In_166);
nand U700 (N_700,In_976,In_1504);
xor U701 (N_701,In_2124,In_174);
nand U702 (N_702,In_2239,In_2343);
nor U703 (N_703,In_169,In_2438);
and U704 (N_704,In_1920,In_1167);
xor U705 (N_705,In_856,In_1810);
and U706 (N_706,In_2366,In_1178);
nor U707 (N_707,In_787,In_2153);
nor U708 (N_708,In_811,In_2355);
nor U709 (N_709,In_1515,In_520);
xnor U710 (N_710,In_962,In_2376);
and U711 (N_711,In_1968,In_204);
nand U712 (N_712,In_635,In_1010);
xnor U713 (N_713,In_1071,In_1582);
or U714 (N_714,In_1333,In_1943);
and U715 (N_715,In_689,In_1615);
nand U716 (N_716,In_845,In_1131);
xnor U717 (N_717,In_2257,In_148);
and U718 (N_718,In_2092,In_2207);
nor U719 (N_719,In_1536,In_1413);
xnor U720 (N_720,In_353,In_2128);
or U721 (N_721,In_738,In_1431);
and U722 (N_722,In_410,In_1557);
xor U723 (N_723,In_808,In_1293);
nand U724 (N_724,In_1228,In_2305);
nor U725 (N_725,In_622,In_7);
and U726 (N_726,In_1473,In_1336);
and U727 (N_727,In_333,In_1199);
and U728 (N_728,In_861,In_680);
nand U729 (N_729,In_1839,In_2264);
or U730 (N_730,In_579,In_1257);
xnor U731 (N_731,In_1972,In_1754);
and U732 (N_732,In_1576,In_417);
and U733 (N_733,In_2495,In_1613);
nor U734 (N_734,In_2023,In_1752);
nor U735 (N_735,In_1472,In_1203);
nand U736 (N_736,In_2075,In_1253);
nand U737 (N_737,In_745,In_1717);
nor U738 (N_738,In_1263,In_2187);
nand U739 (N_739,In_1789,In_2098);
and U740 (N_740,In_619,In_1078);
and U741 (N_741,In_863,In_246);
nand U742 (N_742,In_676,In_534);
or U743 (N_743,In_314,In_2080);
and U744 (N_744,In_796,In_34);
nor U745 (N_745,In_435,In_1825);
or U746 (N_746,In_2466,In_1163);
xnor U747 (N_747,In_2351,In_1669);
nand U748 (N_748,In_2079,In_96);
xor U749 (N_749,In_690,In_2424);
and U750 (N_750,In_1502,In_1363);
nand U751 (N_751,In_1572,In_2145);
nand U752 (N_752,In_1723,In_1378);
nand U753 (N_753,In_817,In_1284);
nor U754 (N_754,In_611,In_1654);
or U755 (N_755,In_115,In_705);
nand U756 (N_756,In_564,In_1200);
nor U757 (N_757,In_946,In_1635);
nor U758 (N_758,In_1155,In_793);
nand U759 (N_759,In_1922,In_1419);
nand U760 (N_760,In_1858,In_2458);
xnor U761 (N_761,In_799,In_824);
xnor U762 (N_762,In_1919,In_427);
xnor U763 (N_763,In_615,In_2212);
and U764 (N_764,In_939,In_884);
and U765 (N_765,In_758,In_661);
nor U766 (N_766,In_359,In_1348);
or U767 (N_767,In_154,In_12);
nand U768 (N_768,In_375,In_2409);
or U769 (N_769,In_966,In_1991);
nand U770 (N_770,In_233,In_648);
nor U771 (N_771,In_2280,In_1355);
and U772 (N_772,In_2417,In_1484);
or U773 (N_773,In_1907,In_256);
and U774 (N_774,In_574,In_1185);
nand U775 (N_775,In_167,In_1648);
xnor U776 (N_776,In_2089,In_1711);
and U777 (N_777,In_1323,In_300);
or U778 (N_778,In_2342,In_1874);
xnor U779 (N_779,In_1259,In_2247);
and U780 (N_780,In_1545,In_1626);
or U781 (N_781,In_302,In_2236);
or U782 (N_782,In_866,In_20);
nor U783 (N_783,In_981,In_1102);
nand U784 (N_784,In_1330,In_1260);
nor U785 (N_785,In_1523,In_1653);
nor U786 (N_786,In_1737,In_192);
xnor U787 (N_787,In_168,In_1182);
nand U788 (N_788,In_294,In_82);
and U789 (N_789,In_1423,In_642);
and U790 (N_790,In_779,In_1009);
nand U791 (N_791,In_2406,In_1037);
and U792 (N_792,In_876,In_107);
or U793 (N_793,In_1633,In_985);
nor U794 (N_794,In_818,In_582);
nor U795 (N_795,In_759,In_1552);
nand U796 (N_796,In_434,In_1510);
or U797 (N_797,In_2102,In_2434);
and U798 (N_798,In_1073,In_2175);
xor U799 (N_799,In_1093,In_1345);
nor U800 (N_800,In_1008,In_1513);
nand U801 (N_801,In_751,In_914);
nor U802 (N_802,In_1663,In_2448);
or U803 (N_803,In_289,In_776);
nand U804 (N_804,In_1899,In_1898);
nand U805 (N_805,In_1307,In_2327);
nand U806 (N_806,In_2199,In_1070);
nor U807 (N_807,In_479,In_1941);
and U808 (N_808,In_1921,In_915);
nor U809 (N_809,In_1445,In_1012);
nor U810 (N_810,In_683,In_2081);
or U811 (N_811,In_896,In_2331);
xor U812 (N_812,In_961,In_1396);
nor U813 (N_813,In_2306,In_2445);
nor U814 (N_814,In_1032,In_2347);
nand U815 (N_815,In_2058,In_865);
or U816 (N_816,In_2114,In_1505);
and U817 (N_817,In_667,In_60);
nand U818 (N_818,In_2028,In_1177);
nand U819 (N_819,In_2307,In_1767);
nand U820 (N_820,In_1391,In_858);
or U821 (N_821,In_1606,In_535);
xnor U822 (N_822,In_841,In_509);
and U823 (N_823,In_744,In_414);
and U824 (N_824,In_1394,In_1180);
nand U825 (N_825,In_1016,In_1196);
xnor U826 (N_826,In_810,In_1042);
nor U827 (N_827,In_2482,In_2375);
nor U828 (N_828,In_1917,In_43);
nand U829 (N_829,In_252,In_1285);
xnor U830 (N_830,In_2107,In_1214);
nand U831 (N_831,In_633,In_2068);
xor U832 (N_832,In_753,In_89);
or U833 (N_833,In_335,In_392);
or U834 (N_834,In_21,In_687);
nor U835 (N_835,In_130,In_1925);
nand U836 (N_836,In_1319,In_2180);
nor U837 (N_837,In_275,In_909);
and U838 (N_838,In_1208,In_350);
xor U839 (N_839,In_1052,In_491);
nor U840 (N_840,In_2293,In_1817);
or U841 (N_841,In_2119,In_1729);
and U842 (N_842,In_960,In_1063);
nor U843 (N_843,In_2296,In_497);
or U844 (N_844,In_297,In_2007);
nor U845 (N_845,In_1528,In_98);
xnor U846 (N_846,In_1161,In_189);
nand U847 (N_847,In_1443,In_129);
and U848 (N_848,In_2329,In_1262);
nand U849 (N_849,In_1283,In_2223);
xnor U850 (N_850,In_907,In_426);
and U851 (N_851,In_998,In_2384);
and U852 (N_852,In_2352,In_1433);
or U853 (N_853,In_539,In_797);
nor U854 (N_854,In_2136,In_823);
xnor U855 (N_855,In_1059,In_868);
or U856 (N_856,In_602,In_2422);
nor U857 (N_857,In_836,In_329);
nand U858 (N_858,In_750,In_1305);
xnor U859 (N_859,In_1241,In_476);
and U860 (N_860,In_1271,In_156);
or U861 (N_861,In_1959,In_1553);
nand U862 (N_862,In_2245,In_468);
nand U863 (N_863,In_1983,In_1693);
nand U864 (N_864,In_1781,In_649);
or U865 (N_865,In_1771,In_1215);
or U866 (N_866,In_528,In_781);
nand U867 (N_867,In_2332,In_2387);
nand U868 (N_868,In_2138,In_1500);
or U869 (N_869,In_764,In_972);
and U870 (N_870,In_25,In_347);
nand U871 (N_871,In_1620,In_728);
or U872 (N_872,In_198,In_506);
and U873 (N_873,In_127,In_2321);
nor U874 (N_874,In_903,In_1275);
nand U875 (N_875,In_1596,In_1272);
nand U876 (N_876,In_1359,In_408);
or U877 (N_877,In_1637,In_711);
or U878 (N_878,In_1151,In_87);
xor U879 (N_879,In_846,In_1640);
nand U880 (N_880,In_889,In_1655);
or U881 (N_881,In_1715,In_1755);
nand U882 (N_882,In_490,In_852);
nor U883 (N_883,In_895,In_1325);
nand U884 (N_884,In_2094,In_2419);
nand U885 (N_885,In_1322,In_336);
nand U886 (N_886,In_537,In_321);
nor U887 (N_887,In_494,In_623);
or U888 (N_888,In_1936,In_1704);
and U889 (N_889,In_72,In_813);
nor U890 (N_890,In_181,In_995);
xnor U891 (N_891,In_1486,In_1885);
and U892 (N_892,In_1610,In_75);
nand U893 (N_893,In_1495,In_862);
nor U894 (N_894,In_30,In_1310);
or U895 (N_895,In_2171,In_1879);
xnor U896 (N_896,In_1496,In_36);
or U897 (N_897,In_1878,In_124);
or U898 (N_898,In_618,In_2474);
nand U899 (N_899,In_45,In_384);
xor U900 (N_900,In_815,In_2130);
and U901 (N_901,In_631,In_1650);
or U902 (N_902,In_1405,In_2371);
xor U903 (N_903,In_766,In_149);
xnor U904 (N_904,In_1670,In_551);
xor U905 (N_905,In_516,In_1843);
xnor U906 (N_906,In_2276,In_173);
xnor U907 (N_907,In_2008,In_1735);
nand U908 (N_908,In_1181,In_109);
nand U909 (N_909,In_1091,In_29);
nand U910 (N_910,In_2464,In_1802);
xnor U911 (N_911,In_1985,In_598);
or U912 (N_912,In_1207,In_2159);
or U913 (N_913,In_859,In_1364);
or U914 (N_914,In_1570,In_778);
xor U915 (N_915,In_1173,In_2263);
nand U916 (N_916,In_1659,In_1003);
xnor U917 (N_917,In_1197,In_1456);
or U918 (N_918,In_132,In_938);
xnor U919 (N_919,In_911,In_2059);
nand U920 (N_920,In_1469,In_1116);
nor U921 (N_921,In_958,In_325);
xnor U922 (N_922,In_432,In_243);
and U923 (N_923,In_367,In_2379);
and U924 (N_924,In_1466,In_803);
xnor U925 (N_925,In_838,In_77);
and U926 (N_926,In_1176,In_662);
or U927 (N_927,In_2082,In_595);
or U928 (N_928,In_678,In_629);
nor U929 (N_929,In_1397,In_979);
xor U930 (N_930,In_655,In_1144);
xnor U931 (N_931,In_1416,In_1331);
and U932 (N_932,In_2497,In_674);
nand U933 (N_933,In_2401,In_495);
nor U934 (N_934,In_882,In_1573);
xor U935 (N_935,In_2278,In_2328);
or U936 (N_936,In_1928,In_1609);
nand U937 (N_937,In_13,In_2093);
or U938 (N_938,In_755,In_463);
nand U939 (N_939,In_299,In_1833);
nand U940 (N_940,In_2340,In_135);
nor U941 (N_941,In_1897,In_2320);
or U942 (N_942,In_2100,In_2182);
or U943 (N_943,In_1175,In_1672);
nor U944 (N_944,In_1826,In_2429);
and U945 (N_945,In_910,In_737);
nor U946 (N_946,In_487,In_2441);
or U947 (N_947,In_2086,In_1805);
and U948 (N_948,In_57,In_1782);
nor U949 (N_949,In_116,In_872);
nand U950 (N_950,In_99,In_2127);
nand U951 (N_951,In_1958,In_722);
and U952 (N_952,In_105,In_1106);
nor U953 (N_953,In_15,In_164);
or U954 (N_954,In_1563,In_2025);
and U955 (N_955,In_1415,In_2302);
nand U956 (N_956,In_1013,In_1614);
and U957 (N_957,In_2374,In_303);
nand U958 (N_958,In_2484,In_1453);
xnor U959 (N_959,In_1168,In_723);
and U960 (N_960,In_1024,In_1937);
xnor U961 (N_961,In_2146,In_2372);
xor U962 (N_962,In_2006,In_1379);
nor U963 (N_963,In_1308,In_1708);
or U964 (N_964,In_2449,In_514);
and U965 (N_965,In_1969,In_954);
or U966 (N_966,In_194,In_70);
and U967 (N_967,In_1014,In_1911);
and U968 (N_968,In_1249,In_828);
nand U969 (N_969,In_853,In_423);
nor U970 (N_970,In_56,In_1744);
xor U971 (N_971,In_1611,In_1372);
nor U972 (N_972,In_1509,In_38);
xor U973 (N_973,In_1749,In_1787);
nor U974 (N_974,In_2399,In_2206);
nor U975 (N_975,In_523,In_1641);
nor U976 (N_976,In_315,In_1747);
nor U977 (N_977,In_2192,In_2172);
nor U978 (N_978,In_1143,In_1873);
nand U979 (N_979,In_1438,In_1954);
nor U980 (N_980,In_2496,In_1018);
nand U981 (N_981,In_1373,In_2141);
nand U982 (N_982,In_125,In_1815);
xnor U983 (N_983,In_1265,In_46);
and U984 (N_984,In_785,In_219);
xor U985 (N_985,In_18,In_713);
xnor U986 (N_986,In_81,In_1792);
or U987 (N_987,In_331,In_770);
or U988 (N_988,In_1769,In_2121);
nand U989 (N_989,In_798,In_529);
or U990 (N_990,In_1631,In_1148);
nor U991 (N_991,In_1069,In_2218);
or U992 (N_992,In_459,In_2120);
and U993 (N_993,In_916,In_2104);
or U994 (N_994,In_1015,In_161);
or U995 (N_995,In_1661,In_277);
and U996 (N_996,In_1720,In_663);
and U997 (N_997,In_1841,In_2357);
or U998 (N_998,In_1135,In_1863);
or U999 (N_999,In_832,In_2475);
or U1000 (N_1000,In_237,In_1195);
and U1001 (N_1001,In_890,In_2174);
nand U1002 (N_1002,In_2437,In_1221);
xor U1003 (N_1003,In_724,In_1906);
and U1004 (N_1004,In_1409,In_1689);
and U1005 (N_1005,In_521,In_2416);
or U1006 (N_1006,In_577,In_2105);
nor U1007 (N_1007,In_1725,In_409);
or U1008 (N_1008,In_1082,In_102);
xnor U1009 (N_1009,In_254,In_1883);
nor U1010 (N_1010,In_1533,In_1707);
xor U1011 (N_1011,In_559,In_1902);
nand U1012 (N_1012,In_2053,In_111);
or U1013 (N_1013,In_37,In_1436);
nor U1014 (N_1014,In_62,In_821);
xnor U1015 (N_1015,In_2450,In_547);
xnor U1016 (N_1016,In_407,In_334);
or U1017 (N_1017,In_1832,In_1146);
xor U1018 (N_1018,In_1414,In_2255);
or U1019 (N_1019,In_1385,In_1402);
and U1020 (N_1020,In_1046,In_1652);
nand U1021 (N_1021,In_483,In_2398);
and U1022 (N_1022,In_2133,In_1721);
or U1023 (N_1023,In_97,In_1393);
nor U1024 (N_1024,In_1020,In_1877);
nand U1025 (N_1025,In_1761,In_1804);
xor U1026 (N_1026,In_1035,In_2021);
nand U1027 (N_1027,In_1351,In_1300);
xnor U1028 (N_1028,In_576,In_1475);
nand U1029 (N_1029,In_1454,In_2408);
and U1030 (N_1030,In_1400,In_2074);
nor U1031 (N_1031,In_1733,In_1434);
nor U1032 (N_1032,In_1994,In_280);
nand U1033 (N_1033,In_40,In_2465);
or U1034 (N_1034,In_122,In_2382);
and U1035 (N_1035,In_1665,In_1571);
and U1036 (N_1036,In_1830,In_1809);
and U1037 (N_1037,In_1569,In_1913);
xnor U1038 (N_1038,In_2076,In_568);
nor U1039 (N_1039,In_1607,In_1387);
nor U1040 (N_1040,In_1254,In_2151);
nand U1041 (N_1041,In_819,In_2389);
nor U1042 (N_1042,In_2241,In_918);
or U1043 (N_1043,In_1219,In_749);
or U1044 (N_1044,In_2414,In_877);
or U1045 (N_1045,In_1074,In_609);
nand U1046 (N_1046,In_1521,In_1647);
and U1047 (N_1047,In_1766,In_1007);
nand U1048 (N_1048,In_1120,In_424);
nor U1049 (N_1049,In_1430,In_2339);
nand U1050 (N_1050,In_2027,In_1341);
nand U1051 (N_1051,In_1245,In_2057);
nor U1052 (N_1052,In_2435,In_2029);
or U1053 (N_1053,In_640,In_2134);
nand U1054 (N_1054,In_1980,In_1476);
and U1055 (N_1055,In_1246,In_2060);
nand U1056 (N_1056,In_983,In_1986);
nor U1057 (N_1057,In_2016,In_507);
nor U1058 (N_1058,In_786,In_1791);
nor U1059 (N_1059,In_405,In_1628);
and U1060 (N_1060,In_1926,In_218);
or U1061 (N_1061,In_2269,In_1842);
or U1062 (N_1062,In_2418,In_1474);
xnor U1063 (N_1063,In_1248,In_2237);
nand U1064 (N_1064,In_1862,In_1492);
nor U1065 (N_1065,In_814,In_338);
nor U1066 (N_1066,In_1002,In_2370);
xnor U1067 (N_1067,In_1406,In_802);
xnor U1068 (N_1068,In_584,In_95);
nand U1069 (N_1069,In_1447,In_2287);
or U1070 (N_1070,In_1165,In_307);
xor U1071 (N_1071,In_377,In_684);
xnor U1072 (N_1072,In_285,In_1940);
nor U1073 (N_1073,In_1988,In_1230);
nor U1074 (N_1074,In_1362,In_39);
nor U1075 (N_1075,In_17,In_1455);
or U1076 (N_1076,In_1066,In_199);
nor U1077 (N_1077,In_1543,In_2215);
and U1078 (N_1078,In_1462,In_339);
and U1079 (N_1079,In_1395,In_2318);
or U1080 (N_1080,In_924,In_1924);
nand U1081 (N_1081,In_1242,In_700);
nor U1082 (N_1082,In_804,In_935);
nand U1083 (N_1083,In_2312,In_2368);
xor U1084 (N_1084,In_1398,In_1977);
and U1085 (N_1085,In_1085,In_222);
and U1086 (N_1086,In_601,In_851);
nand U1087 (N_1087,In_973,In_2156);
and U1088 (N_1088,In_644,In_1900);
xnor U1089 (N_1089,In_123,In_32);
and U1090 (N_1090,In_1232,In_1675);
xor U1091 (N_1091,In_902,In_205);
or U1092 (N_1092,In_2003,In_696);
xnor U1093 (N_1093,In_1234,In_677);
nand U1094 (N_1094,In_1540,In_774);
nor U1095 (N_1095,In_1869,In_2035);
and U1096 (N_1096,In_1644,In_1634);
nand U1097 (N_1097,In_211,In_1295);
or U1098 (N_1098,In_2179,In_2000);
or U1099 (N_1099,In_1627,In_1164);
or U1100 (N_1100,In_1837,In_150);
nand U1101 (N_1101,In_1738,In_2314);
nand U1102 (N_1102,In_561,In_1764);
or U1103 (N_1103,In_1064,In_197);
xor U1104 (N_1104,In_1127,In_1238);
and U1105 (N_1105,In_1763,In_1541);
nand U1106 (N_1106,In_2266,In_2012);
nand U1107 (N_1107,In_2048,In_530);
nand U1108 (N_1108,In_448,In_1352);
nand U1109 (N_1109,In_2335,In_930);
xor U1110 (N_1110,In_1121,In_952);
and U1111 (N_1111,In_214,In_2110);
and U1112 (N_1112,In_2462,In_1574);
xor U1113 (N_1113,In_1905,In_1380);
or U1114 (N_1114,In_446,In_2485);
xnor U1115 (N_1115,In_1586,In_822);
nand U1116 (N_1116,In_363,In_641);
nand U1117 (N_1117,In_2167,In_500);
xor U1118 (N_1118,In_554,In_1894);
nor U1119 (N_1119,In_1566,In_371);
and U1120 (N_1120,In_2205,In_143);
or U1121 (N_1121,In_928,In_994);
xor U1122 (N_1122,In_1043,In_986);
nand U1123 (N_1123,In_2176,In_484);
and U1124 (N_1124,In_322,In_1332);
and U1125 (N_1125,In_351,In_306);
or U1126 (N_1126,In_453,In_941);
nor U1127 (N_1127,In_2031,In_366);
nand U1128 (N_1128,In_626,In_1965);
nand U1129 (N_1129,In_971,In_5);
and U1130 (N_1130,In_1231,In_217);
xor U1131 (N_1131,In_1732,In_1588);
or U1132 (N_1132,In_1524,In_730);
xor U1133 (N_1133,In_1957,In_2193);
and U1134 (N_1134,In_1149,In_2111);
nand U1135 (N_1135,In_1522,In_1281);
xnor U1136 (N_1136,In_2064,In_1354);
xor U1137 (N_1137,In_2091,In_2267);
nand U1138 (N_1138,In_951,In_1005);
nand U1139 (N_1139,In_922,In_2373);
nor U1140 (N_1140,In_1916,In_268);
nor U1141 (N_1141,In_2407,In_1227);
or U1142 (N_1142,In_524,In_1831);
and U1143 (N_1143,In_1183,In_1651);
and U1144 (N_1144,In_545,In_1857);
and U1145 (N_1145,In_1710,In_501);
xnor U1146 (N_1146,In_399,In_247);
nand U1147 (N_1147,In_354,In_1225);
and U1148 (N_1148,In_1047,In_1109);
xor U1149 (N_1149,In_1347,In_2338);
xnor U1150 (N_1150,In_1421,In_1912);
nor U1151 (N_1151,In_2325,In_1235);
nand U1152 (N_1152,In_2037,In_2170);
nor U1153 (N_1153,In_2083,In_913);
nand U1154 (N_1154,In_1656,In_606);
or U1155 (N_1155,In_2345,In_583);
nand U1156 (N_1156,In_850,In_1179);
xnor U1157 (N_1157,In_1981,In_1291);
nor U1158 (N_1158,In_762,In_142);
nand U1159 (N_1159,In_1953,In_1497);
nand U1160 (N_1160,In_1418,In_894);
and U1161 (N_1161,In_460,In_2261);
nor U1162 (N_1162,In_1676,In_1979);
nor U1163 (N_1163,In_2203,In_801);
nand U1164 (N_1164,In_2071,In_566);
nor U1165 (N_1165,In_1327,In_2463);
nor U1166 (N_1166,In_1076,In_2444);
or U1167 (N_1167,In_2033,In_1027);
xor U1168 (N_1168,In_2030,In_1342);
nor U1169 (N_1169,In_1361,In_1871);
or U1170 (N_1170,In_1801,In_2018);
or U1171 (N_1171,In_578,In_1479);
or U1172 (N_1172,In_1884,In_1556);
nor U1173 (N_1173,In_496,In_1973);
nand U1174 (N_1174,In_594,In_2481);
nand U1175 (N_1175,In_445,In_146);
and U1176 (N_1176,In_1503,In_2154);
nand U1177 (N_1177,In_1276,In_634);
nand U1178 (N_1178,In_788,In_2275);
nand U1179 (N_1179,In_2117,In_104);
xnor U1180 (N_1180,In_364,In_133);
or U1181 (N_1181,In_1205,In_854);
nor U1182 (N_1182,In_121,In_1948);
nor U1183 (N_1183,In_1967,In_1067);
nand U1184 (N_1184,In_1797,In_775);
and U1185 (N_1185,In_1820,In_1349);
and U1186 (N_1186,In_1367,In_1790);
xnor U1187 (N_1187,In_2460,In_1807);
nor U1188 (N_1188,In_2194,In_1788);
nor U1189 (N_1189,In_2364,In_1286);
xor U1190 (N_1190,In_1170,In_2234);
xor U1191 (N_1191,In_825,In_780);
or U1192 (N_1192,In_1829,In_2113);
nand U1193 (N_1193,In_614,In_2014);
nand U1194 (N_1194,In_2252,In_1590);
nand U1195 (N_1195,In_681,In_79);
and U1196 (N_1196,In_92,In_538);
and U1197 (N_1197,In_2085,In_1537);
or U1198 (N_1198,In_1962,In_390);
nand U1199 (N_1199,In_1709,In_1602);
or U1200 (N_1200,In_2354,In_103);
nand U1201 (N_1201,In_1683,In_1056);
nand U1202 (N_1202,In_693,In_1882);
nand U1203 (N_1203,In_699,In_1050);
nor U1204 (N_1204,In_1389,In_953);
or U1205 (N_1205,In_1753,In_789);
nand U1206 (N_1206,In_536,In_1999);
nand U1207 (N_1207,In_1561,In_458);
and U1208 (N_1208,In_2211,In_2131);
xor U1209 (N_1209,In_438,In_1038);
or U1210 (N_1210,In_2396,In_1598);
nor U1211 (N_1211,In_2065,In_2166);
xor U1212 (N_1212,In_258,In_2492);
xor U1213 (N_1213,In_332,In_343);
xor U1214 (N_1214,In_1365,In_2217);
and U1215 (N_1215,In_1719,In_316);
nand U1216 (N_1216,In_265,In_1575);
nand U1217 (N_1217,In_2132,In_188);
nor U1218 (N_1218,In_999,In_1463);
and U1219 (N_1219,In_11,In_1088);
nand U1220 (N_1220,In_2295,In_53);
nand U1221 (N_1221,In_1031,In_187);
nor U1222 (N_1222,In_620,In_989);
nor U1223 (N_1223,In_2393,In_553);
xnor U1224 (N_1224,In_1690,In_373);
and U1225 (N_1225,In_2140,In_1206);
nor U1226 (N_1226,In_206,In_1381);
nor U1227 (N_1227,In_71,In_1770);
nand U1228 (N_1228,In_512,In_381);
nor U1229 (N_1229,In_975,In_1812);
nor U1230 (N_1230,In_2426,In_1942);
xnor U1231 (N_1231,In_1712,In_186);
xor U1232 (N_1232,In_1666,In_1426);
nor U1233 (N_1233,In_2377,In_1700);
nand U1234 (N_1234,In_182,In_1226);
or U1235 (N_1235,In_1995,In_76);
nor U1236 (N_1236,In_2169,In_1716);
nand U1237 (N_1237,In_4,In_1220);
nand U1238 (N_1238,In_1304,In_791);
and U1239 (N_1239,In_395,In_1854);
nand U1240 (N_1240,In_599,In_2129);
nor U1241 (N_1241,In_1583,In_1213);
and U1242 (N_1242,In_1041,In_885);
and U1243 (N_1243,In_1480,In_327);
xnor U1244 (N_1244,In_1129,In_492);
and U1245 (N_1245,In_282,In_1818);
and U1246 (N_1246,In_3,In_1439);
xnor U1247 (N_1247,In_1621,In_2273);
xor U1248 (N_1248,In_906,In_2392);
nand U1249 (N_1249,In_42,In_1974);
and U1250 (N_1250,In_1207,In_1731);
or U1251 (N_1251,In_304,In_167);
nand U1252 (N_1252,In_2326,In_1694);
nor U1253 (N_1253,In_1843,In_1250);
xnor U1254 (N_1254,In_1040,In_980);
nor U1255 (N_1255,In_11,In_237);
xor U1256 (N_1256,In_1017,In_2324);
nor U1257 (N_1257,In_2214,In_914);
and U1258 (N_1258,In_2225,In_1704);
nor U1259 (N_1259,In_1478,In_1803);
nor U1260 (N_1260,In_1140,In_2433);
xnor U1261 (N_1261,In_1362,In_950);
and U1262 (N_1262,In_1487,In_25);
or U1263 (N_1263,In_993,In_1582);
nor U1264 (N_1264,In_716,In_116);
nand U1265 (N_1265,In_925,In_221);
nand U1266 (N_1266,In_2017,In_1751);
and U1267 (N_1267,In_1470,In_122);
nor U1268 (N_1268,In_1850,In_1670);
nor U1269 (N_1269,In_1710,In_2144);
and U1270 (N_1270,In_583,In_1880);
and U1271 (N_1271,In_256,In_414);
and U1272 (N_1272,In_350,In_2477);
xnor U1273 (N_1273,In_2298,In_1589);
xor U1274 (N_1274,In_57,In_1331);
nand U1275 (N_1275,In_1973,In_371);
and U1276 (N_1276,In_1102,In_12);
nand U1277 (N_1277,In_2304,In_2217);
nand U1278 (N_1278,In_229,In_1080);
xnor U1279 (N_1279,In_1030,In_1905);
nor U1280 (N_1280,In_1899,In_2100);
and U1281 (N_1281,In_2250,In_1885);
xnor U1282 (N_1282,In_1370,In_607);
nor U1283 (N_1283,In_1780,In_981);
or U1284 (N_1284,In_1104,In_616);
or U1285 (N_1285,In_617,In_290);
nand U1286 (N_1286,In_2348,In_1827);
xor U1287 (N_1287,In_723,In_749);
or U1288 (N_1288,In_838,In_369);
and U1289 (N_1289,In_555,In_2398);
xnor U1290 (N_1290,In_2499,In_508);
and U1291 (N_1291,In_2182,In_1236);
xnor U1292 (N_1292,In_855,In_1089);
nand U1293 (N_1293,In_1540,In_970);
or U1294 (N_1294,In_267,In_1164);
xnor U1295 (N_1295,In_2131,In_2462);
nor U1296 (N_1296,In_2385,In_1197);
xnor U1297 (N_1297,In_1734,In_1657);
and U1298 (N_1298,In_2413,In_1285);
nor U1299 (N_1299,In_89,In_1111);
and U1300 (N_1300,In_1843,In_1804);
or U1301 (N_1301,In_1852,In_587);
nor U1302 (N_1302,In_2322,In_1091);
xnor U1303 (N_1303,In_1192,In_2350);
nor U1304 (N_1304,In_201,In_1393);
nand U1305 (N_1305,In_542,In_523);
and U1306 (N_1306,In_662,In_143);
xnor U1307 (N_1307,In_136,In_1640);
and U1308 (N_1308,In_664,In_246);
and U1309 (N_1309,In_2188,In_2346);
and U1310 (N_1310,In_1199,In_68);
and U1311 (N_1311,In_765,In_2009);
xnor U1312 (N_1312,In_981,In_1448);
nor U1313 (N_1313,In_397,In_1926);
xor U1314 (N_1314,In_2313,In_2124);
nand U1315 (N_1315,In_1963,In_1418);
and U1316 (N_1316,In_542,In_1672);
xnor U1317 (N_1317,In_2180,In_821);
nor U1318 (N_1318,In_2253,In_2124);
or U1319 (N_1319,In_2395,In_68);
nor U1320 (N_1320,In_92,In_1654);
or U1321 (N_1321,In_278,In_1069);
xor U1322 (N_1322,In_1521,In_1892);
nand U1323 (N_1323,In_1983,In_2084);
xor U1324 (N_1324,In_1900,In_1684);
xnor U1325 (N_1325,In_304,In_694);
or U1326 (N_1326,In_590,In_2175);
xor U1327 (N_1327,In_172,In_503);
or U1328 (N_1328,In_374,In_1553);
xor U1329 (N_1329,In_2310,In_1691);
nor U1330 (N_1330,In_1011,In_130);
xor U1331 (N_1331,In_102,In_1532);
nand U1332 (N_1332,In_1663,In_2369);
nor U1333 (N_1333,In_1537,In_1808);
nor U1334 (N_1334,In_1320,In_2142);
or U1335 (N_1335,In_633,In_2052);
or U1336 (N_1336,In_308,In_352);
nand U1337 (N_1337,In_1700,In_1680);
and U1338 (N_1338,In_1287,In_800);
nor U1339 (N_1339,In_1002,In_169);
nor U1340 (N_1340,In_976,In_2425);
or U1341 (N_1341,In_2166,In_1438);
xor U1342 (N_1342,In_1457,In_1558);
xor U1343 (N_1343,In_31,In_1469);
xnor U1344 (N_1344,In_988,In_2358);
nand U1345 (N_1345,In_2156,In_1836);
xnor U1346 (N_1346,In_595,In_1552);
nor U1347 (N_1347,In_2116,In_967);
xnor U1348 (N_1348,In_647,In_621);
and U1349 (N_1349,In_2128,In_2286);
and U1350 (N_1350,In_261,In_476);
and U1351 (N_1351,In_1929,In_1662);
or U1352 (N_1352,In_2356,In_853);
and U1353 (N_1353,In_1737,In_1034);
xnor U1354 (N_1354,In_2100,In_1977);
xor U1355 (N_1355,In_2206,In_533);
or U1356 (N_1356,In_1692,In_2176);
and U1357 (N_1357,In_74,In_217);
or U1358 (N_1358,In_2100,In_995);
or U1359 (N_1359,In_2207,In_53);
nor U1360 (N_1360,In_1977,In_385);
nand U1361 (N_1361,In_2226,In_2209);
or U1362 (N_1362,In_1716,In_893);
or U1363 (N_1363,In_2272,In_445);
nand U1364 (N_1364,In_1202,In_1206);
xnor U1365 (N_1365,In_1919,In_1138);
or U1366 (N_1366,In_921,In_1864);
or U1367 (N_1367,In_26,In_1192);
or U1368 (N_1368,In_770,In_748);
or U1369 (N_1369,In_2194,In_854);
and U1370 (N_1370,In_481,In_608);
xor U1371 (N_1371,In_2382,In_493);
nor U1372 (N_1372,In_1594,In_782);
or U1373 (N_1373,In_1405,In_1176);
nand U1374 (N_1374,In_2298,In_1949);
or U1375 (N_1375,In_1586,In_2338);
xor U1376 (N_1376,In_1408,In_202);
or U1377 (N_1377,In_1376,In_2091);
nor U1378 (N_1378,In_2192,In_2111);
and U1379 (N_1379,In_1033,In_915);
nor U1380 (N_1380,In_329,In_2416);
xnor U1381 (N_1381,In_1976,In_446);
nor U1382 (N_1382,In_116,In_1767);
and U1383 (N_1383,In_678,In_165);
and U1384 (N_1384,In_2281,In_1468);
nand U1385 (N_1385,In_444,In_1722);
nand U1386 (N_1386,In_870,In_849);
xnor U1387 (N_1387,In_2036,In_850);
nand U1388 (N_1388,In_807,In_2476);
or U1389 (N_1389,In_541,In_1726);
nand U1390 (N_1390,In_1250,In_95);
nor U1391 (N_1391,In_717,In_749);
or U1392 (N_1392,In_2493,In_1925);
nand U1393 (N_1393,In_1162,In_2014);
xor U1394 (N_1394,In_608,In_943);
nand U1395 (N_1395,In_1824,In_2444);
and U1396 (N_1396,In_1501,In_1936);
or U1397 (N_1397,In_760,In_1379);
nor U1398 (N_1398,In_2164,In_983);
xnor U1399 (N_1399,In_208,In_2264);
and U1400 (N_1400,In_2223,In_2253);
xor U1401 (N_1401,In_2433,In_566);
nand U1402 (N_1402,In_412,In_2275);
xnor U1403 (N_1403,In_686,In_388);
or U1404 (N_1404,In_877,In_300);
xor U1405 (N_1405,In_2433,In_773);
nor U1406 (N_1406,In_287,In_2050);
nand U1407 (N_1407,In_758,In_2011);
and U1408 (N_1408,In_2043,In_2465);
or U1409 (N_1409,In_311,In_1815);
nand U1410 (N_1410,In_1036,In_1785);
or U1411 (N_1411,In_1629,In_405);
nor U1412 (N_1412,In_389,In_234);
xor U1413 (N_1413,In_570,In_680);
and U1414 (N_1414,In_1425,In_81);
and U1415 (N_1415,In_638,In_450);
or U1416 (N_1416,In_1128,In_127);
nand U1417 (N_1417,In_1584,In_1753);
xnor U1418 (N_1418,In_2138,In_1680);
xor U1419 (N_1419,In_1132,In_1728);
xor U1420 (N_1420,In_608,In_2440);
nor U1421 (N_1421,In_2423,In_799);
xnor U1422 (N_1422,In_57,In_2152);
nor U1423 (N_1423,In_1549,In_493);
or U1424 (N_1424,In_2357,In_6);
nand U1425 (N_1425,In_321,In_534);
nand U1426 (N_1426,In_2250,In_822);
and U1427 (N_1427,In_238,In_2432);
nand U1428 (N_1428,In_1902,In_1854);
and U1429 (N_1429,In_1356,In_1711);
and U1430 (N_1430,In_693,In_2370);
or U1431 (N_1431,In_2496,In_782);
or U1432 (N_1432,In_31,In_751);
and U1433 (N_1433,In_2477,In_911);
nor U1434 (N_1434,In_1370,In_1899);
nor U1435 (N_1435,In_1845,In_1420);
or U1436 (N_1436,In_441,In_826);
xor U1437 (N_1437,In_2164,In_2296);
nor U1438 (N_1438,In_896,In_539);
and U1439 (N_1439,In_1892,In_1530);
and U1440 (N_1440,In_147,In_533);
nor U1441 (N_1441,In_127,In_1785);
and U1442 (N_1442,In_1001,In_1013);
nand U1443 (N_1443,In_1251,In_1285);
nor U1444 (N_1444,In_1786,In_2152);
or U1445 (N_1445,In_631,In_2258);
nand U1446 (N_1446,In_1812,In_2183);
and U1447 (N_1447,In_24,In_691);
and U1448 (N_1448,In_898,In_404);
or U1449 (N_1449,In_600,In_1428);
and U1450 (N_1450,In_399,In_1257);
or U1451 (N_1451,In_775,In_1746);
nand U1452 (N_1452,In_1312,In_923);
nor U1453 (N_1453,In_1825,In_467);
or U1454 (N_1454,In_2367,In_926);
nand U1455 (N_1455,In_573,In_1201);
xor U1456 (N_1456,In_1690,In_125);
and U1457 (N_1457,In_1567,In_2048);
or U1458 (N_1458,In_1590,In_6);
or U1459 (N_1459,In_1731,In_611);
or U1460 (N_1460,In_1222,In_1355);
and U1461 (N_1461,In_1751,In_541);
and U1462 (N_1462,In_1712,In_1776);
xor U1463 (N_1463,In_1761,In_1507);
nand U1464 (N_1464,In_499,In_336);
nand U1465 (N_1465,In_1497,In_212);
nand U1466 (N_1466,In_150,In_562);
xnor U1467 (N_1467,In_2327,In_1739);
xnor U1468 (N_1468,In_2345,In_512);
xnor U1469 (N_1469,In_584,In_1569);
or U1470 (N_1470,In_2254,In_2495);
nand U1471 (N_1471,In_1361,In_905);
or U1472 (N_1472,In_1286,In_107);
nand U1473 (N_1473,In_1004,In_2349);
xnor U1474 (N_1474,In_919,In_225);
or U1475 (N_1475,In_1121,In_1428);
and U1476 (N_1476,In_1536,In_363);
nor U1477 (N_1477,In_2011,In_1214);
and U1478 (N_1478,In_1614,In_1342);
nor U1479 (N_1479,In_1726,In_1758);
or U1480 (N_1480,In_1889,In_1916);
nand U1481 (N_1481,In_1534,In_1841);
xnor U1482 (N_1482,In_1045,In_1953);
or U1483 (N_1483,In_393,In_2380);
or U1484 (N_1484,In_2488,In_972);
xor U1485 (N_1485,In_519,In_626);
nand U1486 (N_1486,In_1655,In_2046);
nand U1487 (N_1487,In_1361,In_439);
xor U1488 (N_1488,In_390,In_1114);
or U1489 (N_1489,In_2206,In_1332);
nor U1490 (N_1490,In_2264,In_417);
xnor U1491 (N_1491,In_2370,In_1164);
or U1492 (N_1492,In_44,In_299);
and U1493 (N_1493,In_2035,In_137);
nor U1494 (N_1494,In_1021,In_1471);
nand U1495 (N_1495,In_1590,In_1256);
and U1496 (N_1496,In_1337,In_1727);
and U1497 (N_1497,In_1927,In_1093);
and U1498 (N_1498,In_1426,In_2219);
nand U1499 (N_1499,In_1876,In_1971);
nor U1500 (N_1500,In_1049,In_172);
xor U1501 (N_1501,In_1078,In_271);
xor U1502 (N_1502,In_668,In_178);
nand U1503 (N_1503,In_2284,In_1778);
and U1504 (N_1504,In_1110,In_1373);
nand U1505 (N_1505,In_151,In_1106);
nand U1506 (N_1506,In_2412,In_2096);
nand U1507 (N_1507,In_984,In_1098);
xnor U1508 (N_1508,In_739,In_510);
and U1509 (N_1509,In_1016,In_245);
nor U1510 (N_1510,In_265,In_1919);
xor U1511 (N_1511,In_568,In_2466);
nor U1512 (N_1512,In_1456,In_1513);
and U1513 (N_1513,In_1007,In_1823);
or U1514 (N_1514,In_82,In_1689);
nand U1515 (N_1515,In_478,In_1655);
nand U1516 (N_1516,In_406,In_1094);
nor U1517 (N_1517,In_2483,In_773);
nand U1518 (N_1518,In_419,In_2155);
and U1519 (N_1519,In_1400,In_2245);
nand U1520 (N_1520,In_1451,In_795);
and U1521 (N_1521,In_1440,In_437);
or U1522 (N_1522,In_2129,In_1272);
or U1523 (N_1523,In_1414,In_1879);
and U1524 (N_1524,In_2340,In_356);
xnor U1525 (N_1525,In_842,In_572);
xnor U1526 (N_1526,In_2369,In_606);
or U1527 (N_1527,In_1432,In_1752);
and U1528 (N_1528,In_546,In_2153);
and U1529 (N_1529,In_2191,In_1187);
nor U1530 (N_1530,In_247,In_566);
nor U1531 (N_1531,In_1480,In_2262);
nor U1532 (N_1532,In_1126,In_2482);
nor U1533 (N_1533,In_317,In_1403);
and U1534 (N_1534,In_1093,In_290);
nand U1535 (N_1535,In_1176,In_2485);
nand U1536 (N_1536,In_2158,In_1417);
nor U1537 (N_1537,In_1527,In_407);
nor U1538 (N_1538,In_1999,In_2335);
nand U1539 (N_1539,In_1878,In_2196);
and U1540 (N_1540,In_2266,In_602);
nor U1541 (N_1541,In_496,In_2167);
nor U1542 (N_1542,In_1331,In_2076);
nor U1543 (N_1543,In_1768,In_244);
nand U1544 (N_1544,In_1421,In_323);
xor U1545 (N_1545,In_1114,In_926);
or U1546 (N_1546,In_460,In_1389);
xnor U1547 (N_1547,In_242,In_1926);
and U1548 (N_1548,In_1092,In_604);
or U1549 (N_1549,In_2005,In_1091);
nor U1550 (N_1550,In_1692,In_897);
or U1551 (N_1551,In_1531,In_2432);
xor U1552 (N_1552,In_2014,In_1534);
nor U1553 (N_1553,In_1541,In_1128);
xor U1554 (N_1554,In_2197,In_1191);
nor U1555 (N_1555,In_2230,In_271);
xor U1556 (N_1556,In_215,In_1532);
and U1557 (N_1557,In_2165,In_533);
and U1558 (N_1558,In_1172,In_2427);
and U1559 (N_1559,In_1224,In_1466);
xnor U1560 (N_1560,In_786,In_711);
or U1561 (N_1561,In_1653,In_2035);
xor U1562 (N_1562,In_1568,In_1070);
xnor U1563 (N_1563,In_1682,In_1703);
xor U1564 (N_1564,In_493,In_1418);
nor U1565 (N_1565,In_1871,In_819);
or U1566 (N_1566,In_2087,In_1018);
and U1567 (N_1567,In_954,In_2418);
and U1568 (N_1568,In_148,In_1477);
xor U1569 (N_1569,In_441,In_2108);
and U1570 (N_1570,In_665,In_917);
nor U1571 (N_1571,In_1961,In_2220);
nor U1572 (N_1572,In_451,In_2450);
and U1573 (N_1573,In_1967,In_1168);
xor U1574 (N_1574,In_1272,In_333);
nor U1575 (N_1575,In_1332,In_2347);
or U1576 (N_1576,In_1361,In_505);
or U1577 (N_1577,In_1593,In_341);
nand U1578 (N_1578,In_2370,In_1736);
nand U1579 (N_1579,In_2408,In_185);
nand U1580 (N_1580,In_1921,In_1372);
and U1581 (N_1581,In_749,In_1982);
nor U1582 (N_1582,In_2172,In_122);
and U1583 (N_1583,In_312,In_1594);
nor U1584 (N_1584,In_520,In_2248);
or U1585 (N_1585,In_238,In_78);
or U1586 (N_1586,In_1825,In_2176);
xor U1587 (N_1587,In_1589,In_2450);
or U1588 (N_1588,In_608,In_1011);
nand U1589 (N_1589,In_240,In_1206);
and U1590 (N_1590,In_1633,In_765);
nand U1591 (N_1591,In_2418,In_1352);
nor U1592 (N_1592,In_1201,In_1454);
nand U1593 (N_1593,In_657,In_836);
nor U1594 (N_1594,In_582,In_271);
nor U1595 (N_1595,In_2314,In_1263);
xnor U1596 (N_1596,In_2309,In_2019);
nor U1597 (N_1597,In_1356,In_1770);
nand U1598 (N_1598,In_538,In_474);
nor U1599 (N_1599,In_596,In_1920);
xnor U1600 (N_1600,In_1512,In_1292);
nand U1601 (N_1601,In_1925,In_1190);
and U1602 (N_1602,In_222,In_2361);
nand U1603 (N_1603,In_703,In_104);
and U1604 (N_1604,In_875,In_2063);
xor U1605 (N_1605,In_551,In_327);
nand U1606 (N_1606,In_2444,In_1813);
nor U1607 (N_1607,In_36,In_830);
or U1608 (N_1608,In_126,In_901);
and U1609 (N_1609,In_1434,In_777);
and U1610 (N_1610,In_1373,In_994);
or U1611 (N_1611,In_331,In_1837);
nor U1612 (N_1612,In_740,In_1594);
xor U1613 (N_1613,In_2257,In_94);
nand U1614 (N_1614,In_2445,In_662);
nand U1615 (N_1615,In_2049,In_1845);
and U1616 (N_1616,In_1769,In_171);
xor U1617 (N_1617,In_1755,In_2366);
and U1618 (N_1618,In_137,In_772);
or U1619 (N_1619,In_1555,In_273);
nand U1620 (N_1620,In_1653,In_44);
or U1621 (N_1621,In_1495,In_1164);
xnor U1622 (N_1622,In_261,In_1479);
xnor U1623 (N_1623,In_1317,In_617);
or U1624 (N_1624,In_2075,In_71);
or U1625 (N_1625,In_1003,In_268);
nand U1626 (N_1626,In_930,In_1835);
nor U1627 (N_1627,In_2236,In_798);
nand U1628 (N_1628,In_833,In_1309);
xor U1629 (N_1629,In_477,In_1414);
xnor U1630 (N_1630,In_921,In_1386);
nand U1631 (N_1631,In_2485,In_2406);
xnor U1632 (N_1632,In_1922,In_1390);
nor U1633 (N_1633,In_374,In_1255);
nand U1634 (N_1634,In_855,In_678);
or U1635 (N_1635,In_1520,In_672);
or U1636 (N_1636,In_889,In_160);
nand U1637 (N_1637,In_262,In_2030);
and U1638 (N_1638,In_458,In_1891);
nand U1639 (N_1639,In_1092,In_1744);
or U1640 (N_1640,In_436,In_480);
nand U1641 (N_1641,In_462,In_2137);
xnor U1642 (N_1642,In_1012,In_753);
or U1643 (N_1643,In_172,In_914);
and U1644 (N_1644,In_1881,In_2455);
xor U1645 (N_1645,In_2217,In_358);
and U1646 (N_1646,In_434,In_1827);
xor U1647 (N_1647,In_983,In_2363);
nand U1648 (N_1648,In_917,In_2300);
nor U1649 (N_1649,In_129,In_281);
or U1650 (N_1650,In_1104,In_1937);
nor U1651 (N_1651,In_2234,In_2163);
nand U1652 (N_1652,In_717,In_1230);
or U1653 (N_1653,In_1318,In_755);
nand U1654 (N_1654,In_1991,In_1921);
or U1655 (N_1655,In_1368,In_1569);
or U1656 (N_1656,In_1882,In_2246);
nor U1657 (N_1657,In_208,In_528);
and U1658 (N_1658,In_2057,In_2352);
and U1659 (N_1659,In_2408,In_1827);
nand U1660 (N_1660,In_2498,In_975);
or U1661 (N_1661,In_163,In_374);
or U1662 (N_1662,In_2207,In_1914);
and U1663 (N_1663,In_1351,In_2335);
and U1664 (N_1664,In_1700,In_234);
nand U1665 (N_1665,In_441,In_1878);
xnor U1666 (N_1666,In_1105,In_615);
xnor U1667 (N_1667,In_538,In_796);
and U1668 (N_1668,In_1914,In_1574);
or U1669 (N_1669,In_1121,In_1335);
xor U1670 (N_1670,In_2062,In_278);
nand U1671 (N_1671,In_1595,In_1844);
nand U1672 (N_1672,In_115,In_1138);
or U1673 (N_1673,In_1893,In_118);
or U1674 (N_1674,In_776,In_2293);
or U1675 (N_1675,In_2353,In_558);
and U1676 (N_1676,In_1201,In_519);
xor U1677 (N_1677,In_464,In_2258);
or U1678 (N_1678,In_2137,In_773);
and U1679 (N_1679,In_2075,In_216);
or U1680 (N_1680,In_1049,In_1267);
xnor U1681 (N_1681,In_1385,In_2042);
nand U1682 (N_1682,In_823,In_1828);
nor U1683 (N_1683,In_1128,In_23);
nand U1684 (N_1684,In_613,In_1126);
nand U1685 (N_1685,In_86,In_2199);
xor U1686 (N_1686,In_803,In_2201);
xnor U1687 (N_1687,In_414,In_1461);
and U1688 (N_1688,In_1823,In_2492);
nor U1689 (N_1689,In_690,In_763);
and U1690 (N_1690,In_1958,In_1740);
and U1691 (N_1691,In_2217,In_1719);
nand U1692 (N_1692,In_1202,In_1425);
xnor U1693 (N_1693,In_121,In_753);
nand U1694 (N_1694,In_416,In_1087);
xor U1695 (N_1695,In_1729,In_880);
nand U1696 (N_1696,In_905,In_665);
nor U1697 (N_1697,In_1785,In_730);
nand U1698 (N_1698,In_2467,In_777);
nand U1699 (N_1699,In_1376,In_1915);
nor U1700 (N_1700,In_2063,In_937);
nand U1701 (N_1701,In_711,In_1628);
or U1702 (N_1702,In_137,In_2148);
or U1703 (N_1703,In_693,In_653);
and U1704 (N_1704,In_778,In_919);
or U1705 (N_1705,In_1315,In_1398);
or U1706 (N_1706,In_1016,In_2129);
and U1707 (N_1707,In_190,In_108);
or U1708 (N_1708,In_2247,In_1470);
and U1709 (N_1709,In_1108,In_1648);
or U1710 (N_1710,In_1394,In_686);
or U1711 (N_1711,In_1648,In_706);
xor U1712 (N_1712,In_48,In_9);
and U1713 (N_1713,In_1848,In_1049);
xnor U1714 (N_1714,In_1733,In_1330);
xnor U1715 (N_1715,In_1011,In_706);
nor U1716 (N_1716,In_2499,In_842);
nor U1717 (N_1717,In_2110,In_459);
xor U1718 (N_1718,In_82,In_2183);
nand U1719 (N_1719,In_1062,In_2392);
nor U1720 (N_1720,In_1415,In_200);
xnor U1721 (N_1721,In_460,In_1596);
or U1722 (N_1722,In_1900,In_1586);
xnor U1723 (N_1723,In_1711,In_1435);
xnor U1724 (N_1724,In_842,In_2204);
nor U1725 (N_1725,In_2077,In_1682);
and U1726 (N_1726,In_1677,In_1749);
nor U1727 (N_1727,In_1917,In_873);
xor U1728 (N_1728,In_644,In_1445);
nand U1729 (N_1729,In_628,In_43);
nand U1730 (N_1730,In_2399,In_1511);
and U1731 (N_1731,In_1567,In_1944);
and U1732 (N_1732,In_1440,In_1978);
xnor U1733 (N_1733,In_2076,In_2312);
and U1734 (N_1734,In_762,In_2047);
xnor U1735 (N_1735,In_2164,In_1267);
xnor U1736 (N_1736,In_1202,In_2375);
or U1737 (N_1737,In_1585,In_1445);
or U1738 (N_1738,In_2422,In_1185);
nand U1739 (N_1739,In_1127,In_2303);
xor U1740 (N_1740,In_1818,In_1245);
nor U1741 (N_1741,In_984,In_2360);
nor U1742 (N_1742,In_29,In_2275);
nor U1743 (N_1743,In_900,In_2193);
nor U1744 (N_1744,In_2430,In_15);
xor U1745 (N_1745,In_1281,In_1618);
xor U1746 (N_1746,In_252,In_124);
and U1747 (N_1747,In_105,In_1816);
nor U1748 (N_1748,In_1985,In_654);
nor U1749 (N_1749,In_302,In_1468);
and U1750 (N_1750,In_930,In_1127);
nand U1751 (N_1751,In_727,In_602);
xor U1752 (N_1752,In_387,In_34);
or U1753 (N_1753,In_416,In_1526);
and U1754 (N_1754,In_2287,In_2360);
and U1755 (N_1755,In_2452,In_441);
nand U1756 (N_1756,In_2000,In_1589);
nand U1757 (N_1757,In_2208,In_170);
xor U1758 (N_1758,In_953,In_983);
nor U1759 (N_1759,In_1517,In_2321);
and U1760 (N_1760,In_63,In_2196);
nor U1761 (N_1761,In_1247,In_1800);
or U1762 (N_1762,In_2408,In_664);
nand U1763 (N_1763,In_2450,In_80);
nor U1764 (N_1764,In_2330,In_1460);
or U1765 (N_1765,In_742,In_2050);
nor U1766 (N_1766,In_1323,In_883);
and U1767 (N_1767,In_97,In_1638);
or U1768 (N_1768,In_2487,In_822);
and U1769 (N_1769,In_2343,In_1519);
nand U1770 (N_1770,In_1715,In_2415);
nor U1771 (N_1771,In_2475,In_259);
and U1772 (N_1772,In_268,In_1542);
or U1773 (N_1773,In_1848,In_796);
nand U1774 (N_1774,In_1671,In_1887);
nand U1775 (N_1775,In_128,In_2352);
and U1776 (N_1776,In_892,In_1127);
nor U1777 (N_1777,In_351,In_827);
nand U1778 (N_1778,In_738,In_1286);
or U1779 (N_1779,In_1569,In_2153);
or U1780 (N_1780,In_248,In_1039);
and U1781 (N_1781,In_2220,In_1221);
nand U1782 (N_1782,In_2164,In_511);
and U1783 (N_1783,In_2074,In_1712);
nor U1784 (N_1784,In_2288,In_853);
nor U1785 (N_1785,In_536,In_1743);
xor U1786 (N_1786,In_804,In_861);
and U1787 (N_1787,In_1729,In_543);
and U1788 (N_1788,In_30,In_1504);
or U1789 (N_1789,In_1192,In_589);
and U1790 (N_1790,In_289,In_1253);
nand U1791 (N_1791,In_859,In_294);
nor U1792 (N_1792,In_2258,In_1176);
nor U1793 (N_1793,In_2418,In_1037);
nand U1794 (N_1794,In_212,In_1763);
xnor U1795 (N_1795,In_1555,In_290);
or U1796 (N_1796,In_980,In_1602);
and U1797 (N_1797,In_2034,In_1601);
or U1798 (N_1798,In_1352,In_1040);
xor U1799 (N_1799,In_585,In_540);
nor U1800 (N_1800,In_235,In_1668);
nor U1801 (N_1801,In_2241,In_2278);
or U1802 (N_1802,In_2019,In_624);
xnor U1803 (N_1803,In_2234,In_1628);
xor U1804 (N_1804,In_1693,In_661);
and U1805 (N_1805,In_1369,In_736);
nor U1806 (N_1806,In_949,In_1794);
or U1807 (N_1807,In_512,In_1331);
xor U1808 (N_1808,In_1066,In_1172);
and U1809 (N_1809,In_929,In_1032);
and U1810 (N_1810,In_910,In_69);
nor U1811 (N_1811,In_231,In_291);
nor U1812 (N_1812,In_1895,In_1388);
and U1813 (N_1813,In_1378,In_1084);
and U1814 (N_1814,In_1909,In_923);
or U1815 (N_1815,In_335,In_981);
or U1816 (N_1816,In_2057,In_149);
nand U1817 (N_1817,In_1570,In_1643);
or U1818 (N_1818,In_815,In_2099);
and U1819 (N_1819,In_1275,In_684);
nand U1820 (N_1820,In_360,In_1391);
xor U1821 (N_1821,In_1791,In_1561);
or U1822 (N_1822,In_2367,In_825);
nor U1823 (N_1823,In_885,In_1474);
or U1824 (N_1824,In_270,In_1458);
xor U1825 (N_1825,In_656,In_2007);
xnor U1826 (N_1826,In_1638,In_643);
or U1827 (N_1827,In_31,In_2410);
nor U1828 (N_1828,In_2151,In_322);
or U1829 (N_1829,In_2252,In_1971);
nand U1830 (N_1830,In_1146,In_1311);
and U1831 (N_1831,In_1012,In_1743);
nor U1832 (N_1832,In_1310,In_181);
nor U1833 (N_1833,In_694,In_2289);
or U1834 (N_1834,In_189,In_1823);
or U1835 (N_1835,In_2361,In_2041);
xor U1836 (N_1836,In_1154,In_2071);
or U1837 (N_1837,In_1288,In_352);
or U1838 (N_1838,In_561,In_318);
xor U1839 (N_1839,In_1161,In_871);
nand U1840 (N_1840,In_887,In_1392);
nor U1841 (N_1841,In_1490,In_1661);
xor U1842 (N_1842,In_1010,In_37);
nand U1843 (N_1843,In_873,In_1798);
nand U1844 (N_1844,In_2079,In_1598);
xor U1845 (N_1845,In_320,In_1073);
or U1846 (N_1846,In_2125,In_608);
xnor U1847 (N_1847,In_999,In_829);
or U1848 (N_1848,In_830,In_1221);
xnor U1849 (N_1849,In_1687,In_1497);
or U1850 (N_1850,In_133,In_1466);
nor U1851 (N_1851,In_1763,In_1998);
nand U1852 (N_1852,In_1803,In_617);
and U1853 (N_1853,In_1493,In_72);
nor U1854 (N_1854,In_2170,In_349);
nor U1855 (N_1855,In_1853,In_669);
and U1856 (N_1856,In_201,In_1789);
and U1857 (N_1857,In_607,In_322);
or U1858 (N_1858,In_1666,In_2229);
or U1859 (N_1859,In_2329,In_1952);
or U1860 (N_1860,In_1674,In_1054);
and U1861 (N_1861,In_2298,In_223);
xor U1862 (N_1862,In_50,In_2200);
xnor U1863 (N_1863,In_1155,In_2434);
nand U1864 (N_1864,In_1180,In_1641);
nor U1865 (N_1865,In_513,In_2333);
or U1866 (N_1866,In_1312,In_2112);
and U1867 (N_1867,In_1732,In_2411);
xor U1868 (N_1868,In_1496,In_1333);
or U1869 (N_1869,In_344,In_1248);
and U1870 (N_1870,In_1277,In_1977);
and U1871 (N_1871,In_699,In_1072);
xnor U1872 (N_1872,In_2270,In_517);
or U1873 (N_1873,In_990,In_1383);
nor U1874 (N_1874,In_1388,In_1620);
nand U1875 (N_1875,In_1786,In_1801);
nand U1876 (N_1876,In_2402,In_86);
xor U1877 (N_1877,In_928,In_1806);
or U1878 (N_1878,In_1835,In_1008);
nor U1879 (N_1879,In_52,In_344);
or U1880 (N_1880,In_573,In_2135);
nor U1881 (N_1881,In_792,In_947);
xor U1882 (N_1882,In_2184,In_274);
and U1883 (N_1883,In_2089,In_1585);
or U1884 (N_1884,In_2372,In_312);
or U1885 (N_1885,In_2314,In_1848);
nor U1886 (N_1886,In_2395,In_960);
nand U1887 (N_1887,In_948,In_2492);
xnor U1888 (N_1888,In_2352,In_1801);
and U1889 (N_1889,In_1837,In_1954);
and U1890 (N_1890,In_3,In_525);
nor U1891 (N_1891,In_1981,In_1135);
or U1892 (N_1892,In_1629,In_25);
or U1893 (N_1893,In_1964,In_563);
and U1894 (N_1894,In_1148,In_1468);
nor U1895 (N_1895,In_1544,In_2398);
or U1896 (N_1896,In_1855,In_1558);
xor U1897 (N_1897,In_806,In_1588);
xor U1898 (N_1898,In_885,In_1529);
or U1899 (N_1899,In_230,In_684);
nor U1900 (N_1900,In_2355,In_2186);
xnor U1901 (N_1901,In_712,In_1055);
and U1902 (N_1902,In_330,In_303);
xnor U1903 (N_1903,In_795,In_528);
nand U1904 (N_1904,In_841,In_1278);
nand U1905 (N_1905,In_1818,In_1312);
or U1906 (N_1906,In_1417,In_1208);
and U1907 (N_1907,In_2196,In_782);
nand U1908 (N_1908,In_1907,In_1091);
nor U1909 (N_1909,In_1747,In_2346);
nand U1910 (N_1910,In_1713,In_662);
nor U1911 (N_1911,In_1993,In_1924);
or U1912 (N_1912,In_2258,In_995);
nor U1913 (N_1913,In_1178,In_1999);
nand U1914 (N_1914,In_950,In_948);
nand U1915 (N_1915,In_1562,In_975);
nor U1916 (N_1916,In_2314,In_398);
or U1917 (N_1917,In_2101,In_1106);
or U1918 (N_1918,In_1651,In_150);
nand U1919 (N_1919,In_413,In_1480);
or U1920 (N_1920,In_1952,In_596);
nand U1921 (N_1921,In_311,In_2034);
xnor U1922 (N_1922,In_1389,In_1502);
xor U1923 (N_1923,In_17,In_468);
nor U1924 (N_1924,In_2418,In_461);
xnor U1925 (N_1925,In_713,In_1489);
xnor U1926 (N_1926,In_805,In_83);
and U1927 (N_1927,In_73,In_2045);
or U1928 (N_1928,In_2268,In_1779);
nor U1929 (N_1929,In_876,In_1433);
and U1930 (N_1930,In_1035,In_1857);
nor U1931 (N_1931,In_2186,In_735);
nand U1932 (N_1932,In_1842,In_52);
xnor U1933 (N_1933,In_1056,In_1827);
and U1934 (N_1934,In_2097,In_415);
xnor U1935 (N_1935,In_391,In_715);
xnor U1936 (N_1936,In_695,In_1821);
xor U1937 (N_1937,In_403,In_2189);
nand U1938 (N_1938,In_321,In_269);
nand U1939 (N_1939,In_2028,In_294);
nor U1940 (N_1940,In_946,In_524);
or U1941 (N_1941,In_827,In_42);
nand U1942 (N_1942,In_1983,In_1320);
nand U1943 (N_1943,In_423,In_735);
nand U1944 (N_1944,In_257,In_1552);
xor U1945 (N_1945,In_699,In_1122);
xor U1946 (N_1946,In_2079,In_1638);
nor U1947 (N_1947,In_2452,In_403);
and U1948 (N_1948,In_86,In_2317);
and U1949 (N_1949,In_119,In_569);
nor U1950 (N_1950,In_2114,In_1988);
or U1951 (N_1951,In_1353,In_2435);
nand U1952 (N_1952,In_2356,In_2119);
or U1953 (N_1953,In_564,In_600);
xnor U1954 (N_1954,In_2051,In_108);
nand U1955 (N_1955,In_255,In_720);
nor U1956 (N_1956,In_1904,In_342);
nor U1957 (N_1957,In_1423,In_1850);
and U1958 (N_1958,In_1997,In_1803);
xor U1959 (N_1959,In_82,In_2215);
and U1960 (N_1960,In_2222,In_784);
or U1961 (N_1961,In_429,In_1401);
nor U1962 (N_1962,In_942,In_1832);
and U1963 (N_1963,In_2092,In_265);
xor U1964 (N_1964,In_608,In_832);
nor U1965 (N_1965,In_644,In_621);
and U1966 (N_1966,In_1977,In_463);
xor U1967 (N_1967,In_2019,In_2435);
or U1968 (N_1968,In_315,In_551);
xnor U1969 (N_1969,In_712,In_883);
and U1970 (N_1970,In_1210,In_804);
and U1971 (N_1971,In_1780,In_537);
and U1972 (N_1972,In_127,In_1540);
and U1973 (N_1973,In_2129,In_2223);
nor U1974 (N_1974,In_1056,In_1360);
nor U1975 (N_1975,In_1335,In_1312);
or U1976 (N_1976,In_1036,In_28);
or U1977 (N_1977,In_956,In_1246);
nand U1978 (N_1978,In_567,In_1212);
and U1979 (N_1979,In_964,In_2231);
nand U1980 (N_1980,In_2306,In_1496);
nand U1981 (N_1981,In_1406,In_1390);
xor U1982 (N_1982,In_489,In_2028);
nand U1983 (N_1983,In_1161,In_1623);
and U1984 (N_1984,In_127,In_1228);
nand U1985 (N_1985,In_813,In_710);
and U1986 (N_1986,In_2486,In_1685);
and U1987 (N_1987,In_526,In_941);
or U1988 (N_1988,In_1213,In_1436);
nor U1989 (N_1989,In_1705,In_213);
or U1990 (N_1990,In_787,In_1829);
nand U1991 (N_1991,In_195,In_1207);
nand U1992 (N_1992,In_1363,In_1963);
nand U1993 (N_1993,In_1559,In_422);
xor U1994 (N_1994,In_2388,In_2251);
nand U1995 (N_1995,In_279,In_634);
xnor U1996 (N_1996,In_1699,In_2066);
nor U1997 (N_1997,In_2257,In_1181);
nor U1998 (N_1998,In_1575,In_1643);
nand U1999 (N_1999,In_1863,In_168);
nand U2000 (N_2000,In_2392,In_1866);
or U2001 (N_2001,In_652,In_512);
xnor U2002 (N_2002,In_1299,In_422);
or U2003 (N_2003,In_1807,In_1399);
and U2004 (N_2004,In_2149,In_36);
nand U2005 (N_2005,In_472,In_2256);
xor U2006 (N_2006,In_445,In_1527);
or U2007 (N_2007,In_685,In_1443);
and U2008 (N_2008,In_1455,In_2102);
and U2009 (N_2009,In_2374,In_318);
nor U2010 (N_2010,In_939,In_1298);
nor U2011 (N_2011,In_422,In_1220);
and U2012 (N_2012,In_432,In_1409);
and U2013 (N_2013,In_1665,In_1425);
nor U2014 (N_2014,In_1091,In_2032);
nor U2015 (N_2015,In_1148,In_1902);
and U2016 (N_2016,In_342,In_830);
and U2017 (N_2017,In_1198,In_1669);
and U2018 (N_2018,In_1702,In_989);
nor U2019 (N_2019,In_1013,In_530);
or U2020 (N_2020,In_649,In_2338);
nor U2021 (N_2021,In_1720,In_1604);
nand U2022 (N_2022,In_1344,In_218);
nor U2023 (N_2023,In_2043,In_928);
nor U2024 (N_2024,In_1665,In_2078);
and U2025 (N_2025,In_1082,In_2129);
nand U2026 (N_2026,In_1371,In_439);
and U2027 (N_2027,In_798,In_366);
or U2028 (N_2028,In_2271,In_1369);
nand U2029 (N_2029,In_851,In_744);
and U2030 (N_2030,In_782,In_101);
or U2031 (N_2031,In_1282,In_583);
or U2032 (N_2032,In_1890,In_740);
nor U2033 (N_2033,In_121,In_156);
nand U2034 (N_2034,In_1493,In_1912);
nand U2035 (N_2035,In_2368,In_1253);
nor U2036 (N_2036,In_1334,In_987);
and U2037 (N_2037,In_501,In_480);
xor U2038 (N_2038,In_656,In_11);
or U2039 (N_2039,In_508,In_2031);
xnor U2040 (N_2040,In_1993,In_1995);
nor U2041 (N_2041,In_1422,In_2124);
or U2042 (N_2042,In_344,In_506);
nand U2043 (N_2043,In_471,In_1281);
nand U2044 (N_2044,In_372,In_1274);
nor U2045 (N_2045,In_306,In_2366);
nor U2046 (N_2046,In_2413,In_1542);
and U2047 (N_2047,In_142,In_1699);
and U2048 (N_2048,In_549,In_772);
nor U2049 (N_2049,In_1768,In_908);
or U2050 (N_2050,In_1072,In_414);
nand U2051 (N_2051,In_25,In_883);
or U2052 (N_2052,In_1382,In_2345);
nand U2053 (N_2053,In_258,In_2288);
nand U2054 (N_2054,In_1567,In_2340);
nand U2055 (N_2055,In_1697,In_249);
or U2056 (N_2056,In_421,In_1492);
and U2057 (N_2057,In_1763,In_2065);
and U2058 (N_2058,In_1609,In_1374);
xor U2059 (N_2059,In_1162,In_2104);
nor U2060 (N_2060,In_134,In_1168);
nand U2061 (N_2061,In_171,In_1042);
or U2062 (N_2062,In_893,In_1801);
nor U2063 (N_2063,In_2399,In_1134);
xnor U2064 (N_2064,In_789,In_1517);
or U2065 (N_2065,In_428,In_792);
and U2066 (N_2066,In_1217,In_1982);
nor U2067 (N_2067,In_643,In_1031);
nand U2068 (N_2068,In_1099,In_450);
nor U2069 (N_2069,In_994,In_1388);
and U2070 (N_2070,In_361,In_135);
xnor U2071 (N_2071,In_2085,In_2389);
nand U2072 (N_2072,In_900,In_1978);
and U2073 (N_2073,In_1837,In_1623);
or U2074 (N_2074,In_187,In_1995);
and U2075 (N_2075,In_669,In_1904);
and U2076 (N_2076,In_8,In_765);
and U2077 (N_2077,In_1198,In_1440);
xor U2078 (N_2078,In_1530,In_47);
nor U2079 (N_2079,In_1457,In_923);
or U2080 (N_2080,In_188,In_1782);
and U2081 (N_2081,In_1535,In_2134);
nor U2082 (N_2082,In_2102,In_2300);
or U2083 (N_2083,In_2282,In_503);
and U2084 (N_2084,In_494,In_1007);
xnor U2085 (N_2085,In_394,In_1022);
nor U2086 (N_2086,In_890,In_1832);
or U2087 (N_2087,In_610,In_2324);
or U2088 (N_2088,In_2499,In_1477);
nor U2089 (N_2089,In_1386,In_1243);
and U2090 (N_2090,In_2324,In_577);
nor U2091 (N_2091,In_833,In_629);
nor U2092 (N_2092,In_655,In_1145);
and U2093 (N_2093,In_1112,In_1212);
nand U2094 (N_2094,In_1847,In_2039);
or U2095 (N_2095,In_2317,In_2096);
nand U2096 (N_2096,In_1242,In_2368);
xnor U2097 (N_2097,In_942,In_1167);
and U2098 (N_2098,In_1554,In_1384);
xnor U2099 (N_2099,In_470,In_1121);
and U2100 (N_2100,In_1265,In_2033);
or U2101 (N_2101,In_1370,In_1031);
nor U2102 (N_2102,In_626,In_327);
nand U2103 (N_2103,In_483,In_624);
and U2104 (N_2104,In_2041,In_1277);
nor U2105 (N_2105,In_2051,In_1319);
xor U2106 (N_2106,In_2093,In_1099);
nand U2107 (N_2107,In_1035,In_820);
nand U2108 (N_2108,In_1490,In_510);
nand U2109 (N_2109,In_2213,In_123);
or U2110 (N_2110,In_1123,In_508);
xor U2111 (N_2111,In_595,In_1383);
xnor U2112 (N_2112,In_649,In_1298);
nor U2113 (N_2113,In_824,In_1092);
nand U2114 (N_2114,In_155,In_1023);
nand U2115 (N_2115,In_2378,In_269);
nor U2116 (N_2116,In_2025,In_2304);
and U2117 (N_2117,In_665,In_1034);
nor U2118 (N_2118,In_1232,In_826);
nor U2119 (N_2119,In_1726,In_2289);
nand U2120 (N_2120,In_1107,In_28);
xnor U2121 (N_2121,In_538,In_1116);
nand U2122 (N_2122,In_14,In_2180);
and U2123 (N_2123,In_163,In_1391);
or U2124 (N_2124,In_127,In_1627);
and U2125 (N_2125,In_581,In_1200);
nand U2126 (N_2126,In_21,In_1235);
xor U2127 (N_2127,In_63,In_908);
nand U2128 (N_2128,In_995,In_1872);
or U2129 (N_2129,In_1843,In_2077);
xor U2130 (N_2130,In_101,In_106);
nand U2131 (N_2131,In_982,In_2278);
nor U2132 (N_2132,In_642,In_2040);
and U2133 (N_2133,In_148,In_2232);
or U2134 (N_2134,In_2394,In_2251);
xnor U2135 (N_2135,In_711,In_1169);
nand U2136 (N_2136,In_1542,In_2352);
and U2137 (N_2137,In_647,In_1082);
or U2138 (N_2138,In_2301,In_863);
and U2139 (N_2139,In_305,In_2151);
or U2140 (N_2140,In_1460,In_2144);
nand U2141 (N_2141,In_1388,In_1035);
or U2142 (N_2142,In_2073,In_394);
xor U2143 (N_2143,In_131,In_19);
nand U2144 (N_2144,In_2037,In_1989);
and U2145 (N_2145,In_1460,In_680);
nor U2146 (N_2146,In_677,In_257);
xnor U2147 (N_2147,In_974,In_606);
xor U2148 (N_2148,In_1739,In_1938);
xor U2149 (N_2149,In_279,In_2213);
and U2150 (N_2150,In_465,In_2442);
xnor U2151 (N_2151,In_145,In_1159);
nor U2152 (N_2152,In_203,In_1420);
and U2153 (N_2153,In_1273,In_187);
nor U2154 (N_2154,In_214,In_1755);
nor U2155 (N_2155,In_1784,In_1857);
or U2156 (N_2156,In_1539,In_1648);
nor U2157 (N_2157,In_2409,In_1020);
and U2158 (N_2158,In_6,In_1228);
xnor U2159 (N_2159,In_2360,In_120);
or U2160 (N_2160,In_1270,In_638);
xor U2161 (N_2161,In_855,In_375);
nand U2162 (N_2162,In_1984,In_445);
xor U2163 (N_2163,In_1739,In_621);
xnor U2164 (N_2164,In_2389,In_1868);
or U2165 (N_2165,In_1237,In_643);
or U2166 (N_2166,In_2188,In_337);
and U2167 (N_2167,In_1619,In_1162);
xor U2168 (N_2168,In_432,In_1304);
nor U2169 (N_2169,In_2028,In_1259);
nor U2170 (N_2170,In_1185,In_882);
or U2171 (N_2171,In_1781,In_1557);
nor U2172 (N_2172,In_1611,In_1691);
or U2173 (N_2173,In_1328,In_1257);
and U2174 (N_2174,In_1878,In_1659);
and U2175 (N_2175,In_625,In_2439);
and U2176 (N_2176,In_2071,In_1669);
or U2177 (N_2177,In_2304,In_337);
nand U2178 (N_2178,In_95,In_2134);
and U2179 (N_2179,In_2227,In_92);
nand U2180 (N_2180,In_1238,In_474);
nand U2181 (N_2181,In_767,In_2211);
nand U2182 (N_2182,In_1999,In_1187);
or U2183 (N_2183,In_1944,In_968);
nor U2184 (N_2184,In_1286,In_1809);
or U2185 (N_2185,In_1616,In_2216);
nor U2186 (N_2186,In_1826,In_1693);
xnor U2187 (N_2187,In_165,In_1305);
or U2188 (N_2188,In_1970,In_1878);
and U2189 (N_2189,In_974,In_1752);
xnor U2190 (N_2190,In_1719,In_1936);
nand U2191 (N_2191,In_442,In_454);
nor U2192 (N_2192,In_1368,In_2001);
or U2193 (N_2193,In_1927,In_464);
or U2194 (N_2194,In_1204,In_2030);
or U2195 (N_2195,In_18,In_117);
nand U2196 (N_2196,In_599,In_1629);
nand U2197 (N_2197,In_1611,In_1938);
and U2198 (N_2198,In_1617,In_1523);
xnor U2199 (N_2199,In_1555,In_1194);
or U2200 (N_2200,In_1808,In_2459);
or U2201 (N_2201,In_6,In_1987);
or U2202 (N_2202,In_1516,In_546);
nand U2203 (N_2203,In_1719,In_1041);
xor U2204 (N_2204,In_818,In_2108);
or U2205 (N_2205,In_2099,In_817);
xor U2206 (N_2206,In_1917,In_490);
xnor U2207 (N_2207,In_890,In_1894);
xor U2208 (N_2208,In_1483,In_1966);
or U2209 (N_2209,In_2495,In_1604);
nor U2210 (N_2210,In_1237,In_262);
xor U2211 (N_2211,In_2023,In_1964);
nand U2212 (N_2212,In_467,In_1034);
and U2213 (N_2213,In_590,In_1930);
nor U2214 (N_2214,In_1426,In_1310);
nand U2215 (N_2215,In_1473,In_149);
xor U2216 (N_2216,In_1800,In_1036);
xor U2217 (N_2217,In_1084,In_618);
or U2218 (N_2218,In_123,In_2324);
nand U2219 (N_2219,In_1082,In_693);
and U2220 (N_2220,In_777,In_554);
or U2221 (N_2221,In_2408,In_806);
xor U2222 (N_2222,In_1296,In_250);
nand U2223 (N_2223,In_1679,In_86);
or U2224 (N_2224,In_943,In_2010);
xnor U2225 (N_2225,In_1182,In_262);
or U2226 (N_2226,In_989,In_588);
and U2227 (N_2227,In_1251,In_903);
or U2228 (N_2228,In_1706,In_2068);
or U2229 (N_2229,In_276,In_1453);
nand U2230 (N_2230,In_607,In_1836);
or U2231 (N_2231,In_2365,In_1215);
or U2232 (N_2232,In_984,In_1517);
and U2233 (N_2233,In_2397,In_1402);
nand U2234 (N_2234,In_2064,In_1972);
or U2235 (N_2235,In_510,In_1135);
or U2236 (N_2236,In_927,In_1098);
nor U2237 (N_2237,In_839,In_1892);
nand U2238 (N_2238,In_1541,In_898);
or U2239 (N_2239,In_1168,In_12);
xnor U2240 (N_2240,In_2040,In_1933);
or U2241 (N_2241,In_981,In_2274);
and U2242 (N_2242,In_534,In_1240);
nor U2243 (N_2243,In_1873,In_276);
xor U2244 (N_2244,In_98,In_588);
or U2245 (N_2245,In_532,In_955);
xor U2246 (N_2246,In_273,In_1827);
nor U2247 (N_2247,In_2145,In_71);
nand U2248 (N_2248,In_1655,In_708);
or U2249 (N_2249,In_2457,In_2011);
xnor U2250 (N_2250,In_2168,In_1960);
or U2251 (N_2251,In_1235,In_1326);
xor U2252 (N_2252,In_1796,In_2330);
xnor U2253 (N_2253,In_2221,In_232);
nand U2254 (N_2254,In_1154,In_467);
and U2255 (N_2255,In_703,In_2111);
nor U2256 (N_2256,In_682,In_1570);
xnor U2257 (N_2257,In_1649,In_2152);
nor U2258 (N_2258,In_2348,In_767);
nand U2259 (N_2259,In_2269,In_1755);
and U2260 (N_2260,In_468,In_1969);
xor U2261 (N_2261,In_1731,In_595);
nand U2262 (N_2262,In_46,In_1809);
and U2263 (N_2263,In_349,In_1508);
xor U2264 (N_2264,In_2108,In_1115);
or U2265 (N_2265,In_119,In_1853);
nor U2266 (N_2266,In_2319,In_1393);
and U2267 (N_2267,In_1873,In_1244);
and U2268 (N_2268,In_1815,In_669);
or U2269 (N_2269,In_731,In_404);
and U2270 (N_2270,In_1952,In_1073);
and U2271 (N_2271,In_1254,In_467);
xnor U2272 (N_2272,In_467,In_151);
or U2273 (N_2273,In_970,In_1780);
xor U2274 (N_2274,In_1632,In_773);
nor U2275 (N_2275,In_862,In_735);
and U2276 (N_2276,In_1483,In_118);
nand U2277 (N_2277,In_2193,In_1654);
nand U2278 (N_2278,In_750,In_292);
xnor U2279 (N_2279,In_1549,In_960);
xor U2280 (N_2280,In_1914,In_772);
and U2281 (N_2281,In_1950,In_2235);
nor U2282 (N_2282,In_2364,In_1658);
xnor U2283 (N_2283,In_2059,In_157);
nor U2284 (N_2284,In_498,In_2268);
or U2285 (N_2285,In_1348,In_1418);
xnor U2286 (N_2286,In_1013,In_819);
nand U2287 (N_2287,In_955,In_103);
nor U2288 (N_2288,In_261,In_589);
nor U2289 (N_2289,In_324,In_836);
nand U2290 (N_2290,In_1804,In_1127);
nand U2291 (N_2291,In_1725,In_638);
nand U2292 (N_2292,In_222,In_1803);
or U2293 (N_2293,In_1294,In_607);
and U2294 (N_2294,In_2451,In_2205);
nand U2295 (N_2295,In_682,In_35);
or U2296 (N_2296,In_603,In_764);
or U2297 (N_2297,In_1743,In_1187);
and U2298 (N_2298,In_2167,In_833);
nand U2299 (N_2299,In_1158,In_414);
or U2300 (N_2300,In_2344,In_1476);
or U2301 (N_2301,In_171,In_1747);
xnor U2302 (N_2302,In_134,In_1269);
and U2303 (N_2303,In_1176,In_2495);
xnor U2304 (N_2304,In_456,In_746);
or U2305 (N_2305,In_2102,In_794);
nor U2306 (N_2306,In_48,In_1952);
and U2307 (N_2307,In_915,In_1516);
nor U2308 (N_2308,In_671,In_1363);
xor U2309 (N_2309,In_1896,In_390);
and U2310 (N_2310,In_504,In_2090);
or U2311 (N_2311,In_1016,In_870);
nor U2312 (N_2312,In_845,In_1364);
nor U2313 (N_2313,In_1860,In_1639);
or U2314 (N_2314,In_1144,In_258);
or U2315 (N_2315,In_1377,In_806);
xnor U2316 (N_2316,In_1390,In_903);
and U2317 (N_2317,In_1256,In_160);
xor U2318 (N_2318,In_592,In_476);
nor U2319 (N_2319,In_2433,In_1116);
and U2320 (N_2320,In_1409,In_2300);
nand U2321 (N_2321,In_1749,In_1908);
and U2322 (N_2322,In_1695,In_624);
or U2323 (N_2323,In_1940,In_1505);
nand U2324 (N_2324,In_1381,In_1172);
and U2325 (N_2325,In_1731,In_1696);
nand U2326 (N_2326,In_133,In_938);
xor U2327 (N_2327,In_2227,In_1615);
xnor U2328 (N_2328,In_2460,In_1776);
nand U2329 (N_2329,In_531,In_701);
xor U2330 (N_2330,In_1472,In_799);
nand U2331 (N_2331,In_428,In_1393);
xor U2332 (N_2332,In_874,In_2443);
nand U2333 (N_2333,In_69,In_2411);
nand U2334 (N_2334,In_2317,In_1957);
nand U2335 (N_2335,In_218,In_848);
or U2336 (N_2336,In_2453,In_1083);
nor U2337 (N_2337,In_1562,In_840);
or U2338 (N_2338,In_2132,In_521);
nor U2339 (N_2339,In_1454,In_183);
or U2340 (N_2340,In_2488,In_1723);
xnor U2341 (N_2341,In_1246,In_1210);
and U2342 (N_2342,In_2158,In_676);
nand U2343 (N_2343,In_161,In_2015);
and U2344 (N_2344,In_822,In_521);
xor U2345 (N_2345,In_1947,In_1946);
and U2346 (N_2346,In_768,In_2467);
xor U2347 (N_2347,In_547,In_1305);
nand U2348 (N_2348,In_615,In_2344);
nor U2349 (N_2349,In_522,In_1572);
and U2350 (N_2350,In_224,In_1665);
and U2351 (N_2351,In_1496,In_143);
nand U2352 (N_2352,In_2438,In_1198);
nand U2353 (N_2353,In_1466,In_2065);
xnor U2354 (N_2354,In_1896,In_1188);
or U2355 (N_2355,In_1566,In_1397);
nor U2356 (N_2356,In_1815,In_1717);
nor U2357 (N_2357,In_2105,In_1431);
nor U2358 (N_2358,In_1535,In_2059);
nor U2359 (N_2359,In_976,In_2435);
nand U2360 (N_2360,In_1669,In_2427);
xor U2361 (N_2361,In_1158,In_1911);
nor U2362 (N_2362,In_630,In_209);
xnor U2363 (N_2363,In_739,In_1207);
or U2364 (N_2364,In_123,In_253);
or U2365 (N_2365,In_253,In_365);
and U2366 (N_2366,In_2275,In_2332);
and U2367 (N_2367,In_1646,In_893);
or U2368 (N_2368,In_951,In_339);
and U2369 (N_2369,In_779,In_2448);
nor U2370 (N_2370,In_10,In_346);
and U2371 (N_2371,In_1283,In_799);
nor U2372 (N_2372,In_2280,In_1006);
nand U2373 (N_2373,In_2397,In_560);
nor U2374 (N_2374,In_1749,In_2494);
and U2375 (N_2375,In_1562,In_851);
or U2376 (N_2376,In_329,In_1633);
xor U2377 (N_2377,In_1795,In_1100);
nand U2378 (N_2378,In_1379,In_1420);
xnor U2379 (N_2379,In_141,In_1347);
xnor U2380 (N_2380,In_790,In_2310);
xor U2381 (N_2381,In_427,In_1783);
and U2382 (N_2382,In_2329,In_1208);
and U2383 (N_2383,In_1950,In_152);
xnor U2384 (N_2384,In_2181,In_303);
or U2385 (N_2385,In_2089,In_1519);
xor U2386 (N_2386,In_2160,In_1935);
nand U2387 (N_2387,In_820,In_1086);
and U2388 (N_2388,In_774,In_1943);
or U2389 (N_2389,In_2464,In_112);
and U2390 (N_2390,In_1938,In_2106);
nor U2391 (N_2391,In_1658,In_1938);
nor U2392 (N_2392,In_1932,In_1188);
or U2393 (N_2393,In_912,In_2066);
nor U2394 (N_2394,In_2181,In_2456);
and U2395 (N_2395,In_450,In_477);
and U2396 (N_2396,In_2123,In_1500);
nand U2397 (N_2397,In_1919,In_1978);
and U2398 (N_2398,In_1190,In_1821);
and U2399 (N_2399,In_2276,In_1939);
or U2400 (N_2400,In_1751,In_1957);
xnor U2401 (N_2401,In_1977,In_361);
and U2402 (N_2402,In_355,In_555);
nand U2403 (N_2403,In_1437,In_1996);
nand U2404 (N_2404,In_1080,In_1202);
and U2405 (N_2405,In_1754,In_1988);
nor U2406 (N_2406,In_1767,In_1261);
nor U2407 (N_2407,In_2038,In_742);
nand U2408 (N_2408,In_2340,In_508);
xor U2409 (N_2409,In_208,In_81);
nor U2410 (N_2410,In_508,In_1164);
xor U2411 (N_2411,In_2495,In_1529);
xor U2412 (N_2412,In_780,In_1256);
xnor U2413 (N_2413,In_1123,In_615);
and U2414 (N_2414,In_1054,In_6);
xor U2415 (N_2415,In_2067,In_641);
and U2416 (N_2416,In_2059,In_1448);
nand U2417 (N_2417,In_361,In_1875);
and U2418 (N_2418,In_1770,In_884);
or U2419 (N_2419,In_615,In_761);
and U2420 (N_2420,In_903,In_1712);
xor U2421 (N_2421,In_427,In_271);
and U2422 (N_2422,In_1414,In_908);
nor U2423 (N_2423,In_549,In_1130);
nand U2424 (N_2424,In_490,In_1532);
and U2425 (N_2425,In_204,In_847);
or U2426 (N_2426,In_1331,In_756);
or U2427 (N_2427,In_1265,In_1377);
and U2428 (N_2428,In_2273,In_1334);
or U2429 (N_2429,In_1304,In_2301);
nor U2430 (N_2430,In_289,In_967);
nand U2431 (N_2431,In_1814,In_1467);
nor U2432 (N_2432,In_439,In_28);
xnor U2433 (N_2433,In_1107,In_1921);
nor U2434 (N_2434,In_1768,In_281);
nor U2435 (N_2435,In_1598,In_1297);
and U2436 (N_2436,In_2390,In_9);
xnor U2437 (N_2437,In_878,In_2128);
nand U2438 (N_2438,In_888,In_96);
nand U2439 (N_2439,In_2361,In_361);
xnor U2440 (N_2440,In_1021,In_1064);
and U2441 (N_2441,In_184,In_2439);
xnor U2442 (N_2442,In_1501,In_1506);
nand U2443 (N_2443,In_483,In_1212);
or U2444 (N_2444,In_6,In_667);
xnor U2445 (N_2445,In_609,In_1934);
nor U2446 (N_2446,In_1662,In_1157);
and U2447 (N_2447,In_2189,In_1524);
or U2448 (N_2448,In_1953,In_265);
and U2449 (N_2449,In_862,In_821);
or U2450 (N_2450,In_942,In_2234);
nor U2451 (N_2451,In_2162,In_129);
nand U2452 (N_2452,In_2472,In_1134);
nor U2453 (N_2453,In_898,In_1465);
nor U2454 (N_2454,In_2173,In_2401);
nor U2455 (N_2455,In_2402,In_223);
nor U2456 (N_2456,In_1045,In_111);
nor U2457 (N_2457,In_1961,In_1496);
or U2458 (N_2458,In_1397,In_491);
xor U2459 (N_2459,In_2095,In_612);
or U2460 (N_2460,In_1418,In_1806);
nor U2461 (N_2461,In_1669,In_591);
xnor U2462 (N_2462,In_1765,In_141);
or U2463 (N_2463,In_1642,In_1655);
nand U2464 (N_2464,In_2378,In_1890);
or U2465 (N_2465,In_115,In_1725);
or U2466 (N_2466,In_1090,In_149);
nor U2467 (N_2467,In_1213,In_2063);
nor U2468 (N_2468,In_983,In_2420);
nor U2469 (N_2469,In_395,In_1523);
nor U2470 (N_2470,In_340,In_2101);
or U2471 (N_2471,In_1872,In_1899);
nand U2472 (N_2472,In_1394,In_2447);
and U2473 (N_2473,In_333,In_340);
nor U2474 (N_2474,In_2208,In_1343);
nor U2475 (N_2475,In_76,In_1905);
and U2476 (N_2476,In_920,In_692);
and U2477 (N_2477,In_302,In_1734);
nand U2478 (N_2478,In_634,In_2178);
xor U2479 (N_2479,In_301,In_67);
xor U2480 (N_2480,In_701,In_351);
or U2481 (N_2481,In_2003,In_1213);
and U2482 (N_2482,In_2388,In_998);
nand U2483 (N_2483,In_2208,In_132);
and U2484 (N_2484,In_2296,In_2006);
and U2485 (N_2485,In_1454,In_2037);
xor U2486 (N_2486,In_147,In_1738);
xnor U2487 (N_2487,In_185,In_1516);
xor U2488 (N_2488,In_666,In_820);
or U2489 (N_2489,In_642,In_1448);
nand U2490 (N_2490,In_1435,In_803);
xnor U2491 (N_2491,In_2349,In_657);
xnor U2492 (N_2492,In_1817,In_1475);
nor U2493 (N_2493,In_1853,In_736);
xnor U2494 (N_2494,In_874,In_1188);
nor U2495 (N_2495,In_1335,In_1892);
nand U2496 (N_2496,In_1732,In_1234);
and U2497 (N_2497,In_70,In_1520);
xor U2498 (N_2498,In_2127,In_2405);
and U2499 (N_2499,In_788,In_1074);
or U2500 (N_2500,In_937,In_214);
or U2501 (N_2501,In_2375,In_902);
and U2502 (N_2502,In_1017,In_2269);
and U2503 (N_2503,In_648,In_1758);
nor U2504 (N_2504,In_1301,In_1092);
and U2505 (N_2505,In_1295,In_1921);
or U2506 (N_2506,In_197,In_658);
or U2507 (N_2507,In_893,In_1182);
and U2508 (N_2508,In_1794,In_178);
or U2509 (N_2509,In_2441,In_1337);
or U2510 (N_2510,In_227,In_1086);
xor U2511 (N_2511,In_2466,In_1002);
nand U2512 (N_2512,In_1738,In_571);
nor U2513 (N_2513,In_1819,In_685);
nand U2514 (N_2514,In_956,In_2210);
or U2515 (N_2515,In_1246,In_1527);
xnor U2516 (N_2516,In_1997,In_669);
xnor U2517 (N_2517,In_550,In_1828);
nand U2518 (N_2518,In_765,In_2404);
or U2519 (N_2519,In_1926,In_1857);
xor U2520 (N_2520,In_213,In_2456);
nand U2521 (N_2521,In_1327,In_904);
or U2522 (N_2522,In_1637,In_2101);
nor U2523 (N_2523,In_1888,In_1950);
nor U2524 (N_2524,In_308,In_419);
xnor U2525 (N_2525,In_1112,In_109);
or U2526 (N_2526,In_2423,In_2045);
or U2527 (N_2527,In_2285,In_238);
xor U2528 (N_2528,In_585,In_1752);
xor U2529 (N_2529,In_1163,In_2319);
xnor U2530 (N_2530,In_2245,In_1243);
nand U2531 (N_2531,In_1001,In_445);
nand U2532 (N_2532,In_617,In_954);
nand U2533 (N_2533,In_804,In_1332);
or U2534 (N_2534,In_1389,In_455);
or U2535 (N_2535,In_674,In_734);
nor U2536 (N_2536,In_2315,In_627);
or U2537 (N_2537,In_68,In_657);
xor U2538 (N_2538,In_1753,In_2169);
or U2539 (N_2539,In_158,In_1769);
nor U2540 (N_2540,In_2017,In_592);
xnor U2541 (N_2541,In_858,In_1713);
or U2542 (N_2542,In_1477,In_5);
nand U2543 (N_2543,In_2303,In_2407);
nor U2544 (N_2544,In_2267,In_2495);
and U2545 (N_2545,In_786,In_1257);
nor U2546 (N_2546,In_6,In_489);
or U2547 (N_2547,In_1462,In_1121);
or U2548 (N_2548,In_2451,In_678);
nor U2549 (N_2549,In_308,In_260);
nand U2550 (N_2550,In_388,In_2114);
or U2551 (N_2551,In_1848,In_1212);
nand U2552 (N_2552,In_2415,In_419);
and U2553 (N_2553,In_191,In_1319);
or U2554 (N_2554,In_1212,In_2002);
nand U2555 (N_2555,In_2142,In_766);
or U2556 (N_2556,In_2027,In_2131);
or U2557 (N_2557,In_2027,In_520);
nand U2558 (N_2558,In_1633,In_1595);
xnor U2559 (N_2559,In_1757,In_1987);
nand U2560 (N_2560,In_1809,In_1492);
and U2561 (N_2561,In_1482,In_1298);
nand U2562 (N_2562,In_1938,In_1252);
and U2563 (N_2563,In_1356,In_590);
or U2564 (N_2564,In_348,In_926);
xor U2565 (N_2565,In_230,In_1069);
and U2566 (N_2566,In_872,In_1572);
or U2567 (N_2567,In_1923,In_2032);
xor U2568 (N_2568,In_744,In_1195);
or U2569 (N_2569,In_1409,In_1385);
and U2570 (N_2570,In_1770,In_390);
or U2571 (N_2571,In_892,In_1707);
or U2572 (N_2572,In_1951,In_2024);
nor U2573 (N_2573,In_2491,In_1965);
xnor U2574 (N_2574,In_522,In_1394);
nand U2575 (N_2575,In_264,In_1757);
and U2576 (N_2576,In_537,In_285);
or U2577 (N_2577,In_913,In_1253);
and U2578 (N_2578,In_190,In_1397);
nor U2579 (N_2579,In_426,In_765);
nand U2580 (N_2580,In_2295,In_281);
nand U2581 (N_2581,In_1905,In_435);
nand U2582 (N_2582,In_1834,In_2037);
or U2583 (N_2583,In_2397,In_1443);
nor U2584 (N_2584,In_361,In_512);
or U2585 (N_2585,In_673,In_780);
and U2586 (N_2586,In_1088,In_2201);
nor U2587 (N_2587,In_571,In_1872);
nor U2588 (N_2588,In_1898,In_882);
or U2589 (N_2589,In_1836,In_2429);
nand U2590 (N_2590,In_2002,In_966);
nor U2591 (N_2591,In_2025,In_139);
or U2592 (N_2592,In_1284,In_1373);
nor U2593 (N_2593,In_1946,In_1228);
or U2594 (N_2594,In_1551,In_2406);
nor U2595 (N_2595,In_2072,In_486);
xor U2596 (N_2596,In_1527,In_641);
nand U2597 (N_2597,In_2354,In_2090);
xnor U2598 (N_2598,In_1989,In_918);
nor U2599 (N_2599,In_1588,In_798);
nand U2600 (N_2600,In_2144,In_1033);
xnor U2601 (N_2601,In_823,In_1252);
nor U2602 (N_2602,In_1657,In_1338);
nand U2603 (N_2603,In_1214,In_2297);
or U2604 (N_2604,In_1846,In_1615);
or U2605 (N_2605,In_1918,In_1737);
xnor U2606 (N_2606,In_2011,In_1236);
nand U2607 (N_2607,In_1493,In_715);
or U2608 (N_2608,In_1785,In_1615);
and U2609 (N_2609,In_2415,In_1351);
nand U2610 (N_2610,In_1693,In_2345);
or U2611 (N_2611,In_2122,In_1060);
or U2612 (N_2612,In_553,In_1189);
or U2613 (N_2613,In_2458,In_2331);
xnor U2614 (N_2614,In_1913,In_1000);
nand U2615 (N_2615,In_1137,In_970);
xor U2616 (N_2616,In_693,In_2463);
nand U2617 (N_2617,In_2,In_809);
nor U2618 (N_2618,In_1567,In_885);
and U2619 (N_2619,In_944,In_711);
and U2620 (N_2620,In_649,In_2243);
nand U2621 (N_2621,In_1057,In_751);
nand U2622 (N_2622,In_507,In_1052);
or U2623 (N_2623,In_915,In_1844);
and U2624 (N_2624,In_1814,In_1779);
or U2625 (N_2625,In_97,In_1898);
and U2626 (N_2626,In_2142,In_214);
nand U2627 (N_2627,In_966,In_2234);
or U2628 (N_2628,In_2054,In_982);
or U2629 (N_2629,In_793,In_395);
and U2630 (N_2630,In_578,In_305);
nor U2631 (N_2631,In_2100,In_729);
and U2632 (N_2632,In_795,In_2352);
and U2633 (N_2633,In_642,In_2054);
and U2634 (N_2634,In_1209,In_823);
nand U2635 (N_2635,In_1945,In_1677);
or U2636 (N_2636,In_1052,In_1086);
nand U2637 (N_2637,In_1961,In_825);
nand U2638 (N_2638,In_821,In_321);
nand U2639 (N_2639,In_2394,In_1177);
or U2640 (N_2640,In_1746,In_721);
and U2641 (N_2641,In_2171,In_1838);
xnor U2642 (N_2642,In_769,In_2254);
xnor U2643 (N_2643,In_590,In_350);
nand U2644 (N_2644,In_83,In_582);
and U2645 (N_2645,In_1134,In_2287);
or U2646 (N_2646,In_738,In_2403);
or U2647 (N_2647,In_935,In_1593);
nor U2648 (N_2648,In_2279,In_1370);
xor U2649 (N_2649,In_1382,In_934);
nor U2650 (N_2650,In_1484,In_2414);
nand U2651 (N_2651,In_1837,In_1436);
or U2652 (N_2652,In_350,In_361);
nor U2653 (N_2653,In_1069,In_752);
xor U2654 (N_2654,In_1304,In_1970);
nor U2655 (N_2655,In_1349,In_442);
xnor U2656 (N_2656,In_1097,In_722);
and U2657 (N_2657,In_1320,In_1673);
nor U2658 (N_2658,In_1457,In_2030);
nor U2659 (N_2659,In_1491,In_704);
nor U2660 (N_2660,In_979,In_207);
nand U2661 (N_2661,In_2078,In_557);
xor U2662 (N_2662,In_2312,In_35);
nor U2663 (N_2663,In_426,In_1922);
nand U2664 (N_2664,In_1760,In_1185);
xnor U2665 (N_2665,In_634,In_1805);
or U2666 (N_2666,In_1768,In_662);
xnor U2667 (N_2667,In_2466,In_218);
nor U2668 (N_2668,In_1360,In_1766);
and U2669 (N_2669,In_795,In_23);
and U2670 (N_2670,In_507,In_2403);
nand U2671 (N_2671,In_103,In_1389);
and U2672 (N_2672,In_759,In_569);
nor U2673 (N_2673,In_1731,In_2355);
xor U2674 (N_2674,In_1313,In_901);
nor U2675 (N_2675,In_863,In_1239);
nor U2676 (N_2676,In_114,In_1695);
xnor U2677 (N_2677,In_1010,In_2156);
nand U2678 (N_2678,In_905,In_2154);
nor U2679 (N_2679,In_686,In_1653);
or U2680 (N_2680,In_934,In_2480);
nor U2681 (N_2681,In_1752,In_996);
nor U2682 (N_2682,In_2043,In_2215);
nor U2683 (N_2683,In_168,In_559);
nor U2684 (N_2684,In_759,In_1497);
xnor U2685 (N_2685,In_2471,In_555);
nor U2686 (N_2686,In_2183,In_25);
xnor U2687 (N_2687,In_1655,In_1312);
xnor U2688 (N_2688,In_1176,In_1344);
xnor U2689 (N_2689,In_2411,In_2437);
nand U2690 (N_2690,In_552,In_1834);
nand U2691 (N_2691,In_84,In_1097);
nor U2692 (N_2692,In_991,In_740);
nand U2693 (N_2693,In_851,In_475);
or U2694 (N_2694,In_608,In_1361);
nor U2695 (N_2695,In_560,In_0);
xnor U2696 (N_2696,In_829,In_1612);
or U2697 (N_2697,In_1653,In_1486);
xor U2698 (N_2698,In_188,In_449);
or U2699 (N_2699,In_1439,In_2320);
or U2700 (N_2700,In_137,In_1490);
or U2701 (N_2701,In_971,In_1070);
xor U2702 (N_2702,In_1116,In_1322);
xnor U2703 (N_2703,In_1549,In_226);
or U2704 (N_2704,In_831,In_1533);
nor U2705 (N_2705,In_1737,In_394);
and U2706 (N_2706,In_969,In_282);
and U2707 (N_2707,In_1434,In_838);
nor U2708 (N_2708,In_1515,In_88);
nor U2709 (N_2709,In_559,In_1748);
or U2710 (N_2710,In_1198,In_1246);
or U2711 (N_2711,In_500,In_1304);
nand U2712 (N_2712,In_161,In_1598);
and U2713 (N_2713,In_1829,In_15);
nor U2714 (N_2714,In_2087,In_1575);
xnor U2715 (N_2715,In_2341,In_1469);
and U2716 (N_2716,In_1972,In_413);
and U2717 (N_2717,In_1375,In_1448);
xnor U2718 (N_2718,In_1477,In_2108);
nor U2719 (N_2719,In_738,In_1481);
xor U2720 (N_2720,In_674,In_1648);
xor U2721 (N_2721,In_860,In_2015);
or U2722 (N_2722,In_806,In_208);
and U2723 (N_2723,In_1758,In_923);
and U2724 (N_2724,In_1816,In_1360);
nor U2725 (N_2725,In_1536,In_1373);
nor U2726 (N_2726,In_2366,In_182);
nor U2727 (N_2727,In_195,In_1965);
xnor U2728 (N_2728,In_1622,In_1764);
nor U2729 (N_2729,In_106,In_1494);
or U2730 (N_2730,In_1872,In_677);
nor U2731 (N_2731,In_726,In_2470);
xor U2732 (N_2732,In_296,In_192);
xor U2733 (N_2733,In_2351,In_682);
nand U2734 (N_2734,In_1662,In_2341);
and U2735 (N_2735,In_570,In_499);
xor U2736 (N_2736,In_247,In_2097);
nand U2737 (N_2737,In_2279,In_1078);
xor U2738 (N_2738,In_772,In_1936);
xnor U2739 (N_2739,In_1179,In_753);
or U2740 (N_2740,In_2167,In_2358);
xnor U2741 (N_2741,In_970,In_510);
nand U2742 (N_2742,In_1600,In_1001);
nor U2743 (N_2743,In_2383,In_2268);
nor U2744 (N_2744,In_1811,In_2237);
nand U2745 (N_2745,In_2067,In_36);
nor U2746 (N_2746,In_2498,In_386);
or U2747 (N_2747,In_1251,In_422);
or U2748 (N_2748,In_2041,In_1098);
and U2749 (N_2749,In_2162,In_927);
nor U2750 (N_2750,In_1313,In_1683);
or U2751 (N_2751,In_2026,In_451);
and U2752 (N_2752,In_220,In_820);
xnor U2753 (N_2753,In_2012,In_14);
nand U2754 (N_2754,In_34,In_39);
or U2755 (N_2755,In_852,In_452);
or U2756 (N_2756,In_2209,In_1350);
nand U2757 (N_2757,In_222,In_1339);
nor U2758 (N_2758,In_846,In_307);
or U2759 (N_2759,In_70,In_484);
and U2760 (N_2760,In_79,In_827);
nand U2761 (N_2761,In_2355,In_1712);
nand U2762 (N_2762,In_492,In_931);
and U2763 (N_2763,In_2260,In_1869);
and U2764 (N_2764,In_2334,In_1361);
xor U2765 (N_2765,In_1329,In_530);
xor U2766 (N_2766,In_1951,In_2002);
xnor U2767 (N_2767,In_2002,In_843);
nand U2768 (N_2768,In_2497,In_170);
and U2769 (N_2769,In_2084,In_2047);
nor U2770 (N_2770,In_2124,In_1237);
nor U2771 (N_2771,In_726,In_1130);
and U2772 (N_2772,In_1204,In_471);
or U2773 (N_2773,In_2308,In_2395);
or U2774 (N_2774,In_2467,In_613);
and U2775 (N_2775,In_508,In_116);
nor U2776 (N_2776,In_147,In_232);
and U2777 (N_2777,In_2396,In_2175);
xor U2778 (N_2778,In_439,In_26);
xor U2779 (N_2779,In_779,In_509);
nand U2780 (N_2780,In_2355,In_951);
xnor U2781 (N_2781,In_427,In_1701);
nor U2782 (N_2782,In_2165,In_2392);
or U2783 (N_2783,In_1986,In_227);
nand U2784 (N_2784,In_882,In_1269);
and U2785 (N_2785,In_62,In_1286);
and U2786 (N_2786,In_511,In_2136);
and U2787 (N_2787,In_2203,In_1147);
nand U2788 (N_2788,In_1399,In_649);
or U2789 (N_2789,In_725,In_51);
xor U2790 (N_2790,In_1942,In_2162);
nand U2791 (N_2791,In_1070,In_997);
or U2792 (N_2792,In_1309,In_579);
or U2793 (N_2793,In_2038,In_1809);
nand U2794 (N_2794,In_493,In_771);
or U2795 (N_2795,In_103,In_1597);
xor U2796 (N_2796,In_1002,In_915);
nor U2797 (N_2797,In_808,In_757);
xor U2798 (N_2798,In_507,In_264);
nor U2799 (N_2799,In_302,In_152);
nand U2800 (N_2800,In_2257,In_325);
nor U2801 (N_2801,In_1837,In_1075);
or U2802 (N_2802,In_2200,In_667);
xnor U2803 (N_2803,In_630,In_1741);
nand U2804 (N_2804,In_277,In_1177);
and U2805 (N_2805,In_1974,In_1390);
nand U2806 (N_2806,In_1193,In_2306);
or U2807 (N_2807,In_1511,In_2430);
nand U2808 (N_2808,In_134,In_1286);
and U2809 (N_2809,In_779,In_94);
xnor U2810 (N_2810,In_2177,In_2250);
and U2811 (N_2811,In_850,In_2427);
and U2812 (N_2812,In_1002,In_1159);
or U2813 (N_2813,In_772,In_578);
or U2814 (N_2814,In_2177,In_1028);
xnor U2815 (N_2815,In_192,In_2085);
and U2816 (N_2816,In_2475,In_2301);
xor U2817 (N_2817,In_1400,In_847);
and U2818 (N_2818,In_667,In_2490);
or U2819 (N_2819,In_2316,In_2344);
or U2820 (N_2820,In_1668,In_637);
nand U2821 (N_2821,In_722,In_951);
xnor U2822 (N_2822,In_2176,In_1364);
xor U2823 (N_2823,In_220,In_2442);
nand U2824 (N_2824,In_2360,In_132);
or U2825 (N_2825,In_1726,In_597);
and U2826 (N_2826,In_1926,In_2175);
xor U2827 (N_2827,In_213,In_2122);
nand U2828 (N_2828,In_1896,In_2092);
and U2829 (N_2829,In_2044,In_2329);
nand U2830 (N_2830,In_1312,In_252);
or U2831 (N_2831,In_624,In_1905);
or U2832 (N_2832,In_904,In_1940);
nor U2833 (N_2833,In_2329,In_1235);
nor U2834 (N_2834,In_2202,In_956);
and U2835 (N_2835,In_368,In_2491);
nand U2836 (N_2836,In_2189,In_1086);
and U2837 (N_2837,In_527,In_2409);
and U2838 (N_2838,In_709,In_442);
nand U2839 (N_2839,In_1203,In_62);
xnor U2840 (N_2840,In_1914,In_2471);
nor U2841 (N_2841,In_1663,In_2133);
and U2842 (N_2842,In_1219,In_1522);
xor U2843 (N_2843,In_1087,In_714);
xnor U2844 (N_2844,In_2073,In_1466);
nor U2845 (N_2845,In_612,In_1947);
nand U2846 (N_2846,In_1015,In_809);
or U2847 (N_2847,In_2030,In_1754);
nor U2848 (N_2848,In_1640,In_1416);
and U2849 (N_2849,In_1197,In_1627);
or U2850 (N_2850,In_843,In_2247);
nor U2851 (N_2851,In_1678,In_2344);
or U2852 (N_2852,In_234,In_2312);
nand U2853 (N_2853,In_1816,In_366);
and U2854 (N_2854,In_2279,In_2057);
and U2855 (N_2855,In_1508,In_513);
and U2856 (N_2856,In_351,In_1973);
nand U2857 (N_2857,In_1589,In_2132);
and U2858 (N_2858,In_94,In_2320);
or U2859 (N_2859,In_1451,In_161);
or U2860 (N_2860,In_644,In_2055);
and U2861 (N_2861,In_1929,In_2267);
or U2862 (N_2862,In_595,In_1687);
nor U2863 (N_2863,In_913,In_1146);
nand U2864 (N_2864,In_944,In_1040);
and U2865 (N_2865,In_2490,In_2100);
xor U2866 (N_2866,In_2215,In_2412);
and U2867 (N_2867,In_2472,In_1760);
and U2868 (N_2868,In_2335,In_954);
and U2869 (N_2869,In_130,In_2177);
xnor U2870 (N_2870,In_1062,In_1313);
nand U2871 (N_2871,In_563,In_1941);
nor U2872 (N_2872,In_1316,In_605);
xor U2873 (N_2873,In_565,In_2413);
and U2874 (N_2874,In_1431,In_39);
or U2875 (N_2875,In_1108,In_2396);
xor U2876 (N_2876,In_1464,In_1078);
or U2877 (N_2877,In_1695,In_2359);
nor U2878 (N_2878,In_643,In_449);
xnor U2879 (N_2879,In_1588,In_48);
or U2880 (N_2880,In_2398,In_867);
or U2881 (N_2881,In_2353,In_1665);
xnor U2882 (N_2882,In_2024,In_1403);
xor U2883 (N_2883,In_299,In_1972);
nand U2884 (N_2884,In_148,In_1695);
xnor U2885 (N_2885,In_202,In_1793);
and U2886 (N_2886,In_2337,In_864);
and U2887 (N_2887,In_1632,In_189);
and U2888 (N_2888,In_1321,In_454);
xnor U2889 (N_2889,In_1943,In_1477);
nor U2890 (N_2890,In_371,In_74);
xnor U2891 (N_2891,In_2109,In_1473);
xor U2892 (N_2892,In_568,In_973);
nor U2893 (N_2893,In_878,In_741);
or U2894 (N_2894,In_2416,In_644);
and U2895 (N_2895,In_2462,In_2096);
nor U2896 (N_2896,In_1704,In_1184);
and U2897 (N_2897,In_1883,In_560);
and U2898 (N_2898,In_1138,In_831);
xor U2899 (N_2899,In_1886,In_2010);
or U2900 (N_2900,In_1444,In_277);
and U2901 (N_2901,In_1272,In_1924);
and U2902 (N_2902,In_2302,In_154);
or U2903 (N_2903,In_55,In_222);
nand U2904 (N_2904,In_2451,In_0);
or U2905 (N_2905,In_57,In_2326);
and U2906 (N_2906,In_1753,In_911);
nand U2907 (N_2907,In_1325,In_2474);
or U2908 (N_2908,In_1387,In_1939);
nor U2909 (N_2909,In_636,In_1340);
or U2910 (N_2910,In_315,In_2226);
nor U2911 (N_2911,In_844,In_429);
and U2912 (N_2912,In_1455,In_2273);
nor U2913 (N_2913,In_1653,In_699);
or U2914 (N_2914,In_1977,In_1537);
and U2915 (N_2915,In_6,In_1063);
or U2916 (N_2916,In_711,In_1643);
xnor U2917 (N_2917,In_1902,In_832);
nand U2918 (N_2918,In_168,In_1501);
nand U2919 (N_2919,In_1135,In_664);
nand U2920 (N_2920,In_1520,In_1788);
or U2921 (N_2921,In_1278,In_2000);
or U2922 (N_2922,In_2304,In_2189);
xor U2923 (N_2923,In_2026,In_1167);
or U2924 (N_2924,In_2463,In_2316);
xnor U2925 (N_2925,In_21,In_1232);
and U2926 (N_2926,In_2302,In_292);
nor U2927 (N_2927,In_325,In_1019);
or U2928 (N_2928,In_2100,In_2049);
xor U2929 (N_2929,In_980,In_1678);
xor U2930 (N_2930,In_568,In_1961);
xor U2931 (N_2931,In_176,In_950);
or U2932 (N_2932,In_1554,In_133);
nand U2933 (N_2933,In_2387,In_1998);
nor U2934 (N_2934,In_1825,In_2049);
or U2935 (N_2935,In_598,In_491);
and U2936 (N_2936,In_1303,In_1450);
or U2937 (N_2937,In_212,In_2108);
nor U2938 (N_2938,In_5,In_2339);
and U2939 (N_2939,In_859,In_1843);
nor U2940 (N_2940,In_1578,In_459);
nor U2941 (N_2941,In_258,In_1398);
or U2942 (N_2942,In_221,In_79);
nand U2943 (N_2943,In_774,In_1898);
and U2944 (N_2944,In_1428,In_1855);
and U2945 (N_2945,In_574,In_467);
or U2946 (N_2946,In_631,In_979);
or U2947 (N_2947,In_1824,In_1976);
and U2948 (N_2948,In_1226,In_49);
xor U2949 (N_2949,In_2416,In_968);
nand U2950 (N_2950,In_1002,In_25);
and U2951 (N_2951,In_2448,In_2099);
nand U2952 (N_2952,In_378,In_2100);
xor U2953 (N_2953,In_1959,In_750);
nor U2954 (N_2954,In_545,In_1379);
or U2955 (N_2955,In_1513,In_1284);
and U2956 (N_2956,In_135,In_1077);
and U2957 (N_2957,In_212,In_1854);
or U2958 (N_2958,In_1191,In_436);
and U2959 (N_2959,In_1144,In_1627);
or U2960 (N_2960,In_1729,In_1822);
and U2961 (N_2961,In_1735,In_1896);
nor U2962 (N_2962,In_816,In_2056);
nand U2963 (N_2963,In_933,In_1315);
xnor U2964 (N_2964,In_961,In_2211);
xnor U2965 (N_2965,In_2133,In_916);
and U2966 (N_2966,In_663,In_217);
nand U2967 (N_2967,In_2416,In_456);
or U2968 (N_2968,In_1938,In_1978);
and U2969 (N_2969,In_118,In_509);
nand U2970 (N_2970,In_2336,In_1494);
nor U2971 (N_2971,In_774,In_955);
or U2972 (N_2972,In_1973,In_668);
and U2973 (N_2973,In_1388,In_2212);
or U2974 (N_2974,In_346,In_211);
nor U2975 (N_2975,In_580,In_14);
or U2976 (N_2976,In_1105,In_716);
nand U2977 (N_2977,In_2383,In_635);
and U2978 (N_2978,In_2193,In_2035);
nor U2979 (N_2979,In_1375,In_736);
xnor U2980 (N_2980,In_1996,In_192);
and U2981 (N_2981,In_229,In_639);
nor U2982 (N_2982,In_394,In_308);
xnor U2983 (N_2983,In_2441,In_835);
or U2984 (N_2984,In_42,In_1730);
nor U2985 (N_2985,In_1759,In_1339);
and U2986 (N_2986,In_1822,In_957);
xor U2987 (N_2987,In_61,In_726);
nand U2988 (N_2988,In_1662,In_765);
or U2989 (N_2989,In_230,In_1615);
or U2990 (N_2990,In_2386,In_1265);
and U2991 (N_2991,In_647,In_162);
xnor U2992 (N_2992,In_434,In_430);
and U2993 (N_2993,In_267,In_1760);
nor U2994 (N_2994,In_1517,In_1055);
xor U2995 (N_2995,In_1098,In_1039);
xor U2996 (N_2996,In_1212,In_2293);
xor U2997 (N_2997,In_1665,In_410);
or U2998 (N_2998,In_814,In_2058);
or U2999 (N_2999,In_1626,In_2449);
nor U3000 (N_3000,In_1648,In_990);
nor U3001 (N_3001,In_1563,In_1497);
and U3002 (N_3002,In_273,In_84);
or U3003 (N_3003,In_19,In_660);
xor U3004 (N_3004,In_1126,In_569);
nand U3005 (N_3005,In_2041,In_268);
or U3006 (N_3006,In_2376,In_188);
or U3007 (N_3007,In_252,In_2341);
nand U3008 (N_3008,In_1220,In_1346);
nor U3009 (N_3009,In_863,In_1137);
nor U3010 (N_3010,In_472,In_1280);
nand U3011 (N_3011,In_729,In_2040);
nor U3012 (N_3012,In_811,In_1307);
and U3013 (N_3013,In_2071,In_2457);
and U3014 (N_3014,In_1323,In_2442);
nor U3015 (N_3015,In_165,In_747);
nand U3016 (N_3016,In_2431,In_228);
or U3017 (N_3017,In_1923,In_964);
and U3018 (N_3018,In_568,In_454);
nor U3019 (N_3019,In_1551,In_979);
xnor U3020 (N_3020,In_545,In_1933);
xnor U3021 (N_3021,In_1235,In_1569);
nand U3022 (N_3022,In_2291,In_1697);
xor U3023 (N_3023,In_249,In_1128);
and U3024 (N_3024,In_2302,In_534);
or U3025 (N_3025,In_2007,In_664);
nand U3026 (N_3026,In_2341,In_1712);
nand U3027 (N_3027,In_1365,In_1141);
or U3028 (N_3028,In_1381,In_884);
and U3029 (N_3029,In_1731,In_790);
nand U3030 (N_3030,In_1314,In_1784);
or U3031 (N_3031,In_333,In_1109);
xor U3032 (N_3032,In_2211,In_307);
and U3033 (N_3033,In_2467,In_6);
nand U3034 (N_3034,In_849,In_1991);
nand U3035 (N_3035,In_245,In_984);
or U3036 (N_3036,In_2157,In_176);
xnor U3037 (N_3037,In_1863,In_1439);
xnor U3038 (N_3038,In_1033,In_1246);
and U3039 (N_3039,In_744,In_791);
nor U3040 (N_3040,In_369,In_1414);
or U3041 (N_3041,In_725,In_233);
nor U3042 (N_3042,In_1566,In_1604);
nand U3043 (N_3043,In_222,In_2250);
xnor U3044 (N_3044,In_863,In_727);
and U3045 (N_3045,In_484,In_778);
nand U3046 (N_3046,In_337,In_2329);
nand U3047 (N_3047,In_440,In_2406);
or U3048 (N_3048,In_1553,In_1941);
nand U3049 (N_3049,In_68,In_1071);
nand U3050 (N_3050,In_1519,In_1687);
nor U3051 (N_3051,In_567,In_333);
nor U3052 (N_3052,In_1163,In_2310);
and U3053 (N_3053,In_675,In_1167);
or U3054 (N_3054,In_2162,In_1823);
nand U3055 (N_3055,In_2134,In_412);
and U3056 (N_3056,In_1935,In_1178);
and U3057 (N_3057,In_1099,In_1123);
xnor U3058 (N_3058,In_607,In_313);
nand U3059 (N_3059,In_328,In_1101);
nor U3060 (N_3060,In_503,In_473);
and U3061 (N_3061,In_2494,In_922);
nand U3062 (N_3062,In_1049,In_1343);
nand U3063 (N_3063,In_679,In_1056);
or U3064 (N_3064,In_186,In_2159);
nand U3065 (N_3065,In_1414,In_604);
or U3066 (N_3066,In_1898,In_1123);
and U3067 (N_3067,In_2003,In_1547);
nand U3068 (N_3068,In_975,In_530);
xor U3069 (N_3069,In_1920,In_1233);
xor U3070 (N_3070,In_1891,In_685);
xor U3071 (N_3071,In_1244,In_475);
or U3072 (N_3072,In_502,In_1232);
or U3073 (N_3073,In_1157,In_1547);
nand U3074 (N_3074,In_428,In_1258);
xor U3075 (N_3075,In_86,In_1946);
nand U3076 (N_3076,In_1403,In_429);
nor U3077 (N_3077,In_940,In_1667);
nor U3078 (N_3078,In_629,In_2266);
nand U3079 (N_3079,In_471,In_84);
and U3080 (N_3080,In_1552,In_1801);
and U3081 (N_3081,In_1562,In_1301);
xor U3082 (N_3082,In_2403,In_1326);
nor U3083 (N_3083,In_457,In_1669);
nor U3084 (N_3084,In_476,In_1897);
nand U3085 (N_3085,In_1731,In_1057);
nor U3086 (N_3086,In_1987,In_2169);
and U3087 (N_3087,In_360,In_138);
or U3088 (N_3088,In_825,In_824);
and U3089 (N_3089,In_1237,In_680);
nor U3090 (N_3090,In_1092,In_1812);
nand U3091 (N_3091,In_576,In_1518);
nor U3092 (N_3092,In_2053,In_98);
and U3093 (N_3093,In_425,In_982);
or U3094 (N_3094,In_2425,In_542);
nand U3095 (N_3095,In_1914,In_2279);
nand U3096 (N_3096,In_730,In_2312);
xnor U3097 (N_3097,In_370,In_2408);
nand U3098 (N_3098,In_2006,In_2324);
or U3099 (N_3099,In_2075,In_2174);
and U3100 (N_3100,In_2457,In_638);
and U3101 (N_3101,In_183,In_5);
and U3102 (N_3102,In_1887,In_1830);
nand U3103 (N_3103,In_979,In_1237);
nand U3104 (N_3104,In_761,In_2319);
nor U3105 (N_3105,In_529,In_1382);
nor U3106 (N_3106,In_1708,In_2397);
and U3107 (N_3107,In_317,In_1069);
xor U3108 (N_3108,In_235,In_1033);
or U3109 (N_3109,In_2282,In_284);
nor U3110 (N_3110,In_537,In_1083);
or U3111 (N_3111,In_882,In_1633);
or U3112 (N_3112,In_164,In_1560);
nor U3113 (N_3113,In_1104,In_2291);
nor U3114 (N_3114,In_2451,In_133);
or U3115 (N_3115,In_682,In_634);
and U3116 (N_3116,In_1251,In_190);
nand U3117 (N_3117,In_118,In_507);
xnor U3118 (N_3118,In_2036,In_829);
nand U3119 (N_3119,In_762,In_736);
xor U3120 (N_3120,In_2132,In_1083);
and U3121 (N_3121,In_946,In_1388);
and U3122 (N_3122,In_644,In_2251);
nor U3123 (N_3123,In_1775,In_2483);
nor U3124 (N_3124,In_1903,In_191);
xnor U3125 (N_3125,In_2125,In_1298);
nand U3126 (N_3126,In_1042,In_1926);
xnor U3127 (N_3127,In_2064,In_324);
nor U3128 (N_3128,In_1773,In_2483);
xnor U3129 (N_3129,In_2087,In_620);
and U3130 (N_3130,In_393,In_2496);
xnor U3131 (N_3131,In_1822,In_325);
or U3132 (N_3132,In_440,In_1220);
and U3133 (N_3133,In_1881,In_330);
nor U3134 (N_3134,In_11,In_1675);
xnor U3135 (N_3135,In_2097,In_1013);
and U3136 (N_3136,In_717,In_980);
nor U3137 (N_3137,In_242,In_1854);
nor U3138 (N_3138,In_2065,In_1241);
or U3139 (N_3139,In_1876,In_2156);
or U3140 (N_3140,In_2012,In_1052);
xnor U3141 (N_3141,In_2059,In_1696);
nor U3142 (N_3142,In_1600,In_1255);
xnor U3143 (N_3143,In_888,In_1290);
nand U3144 (N_3144,In_782,In_1010);
nand U3145 (N_3145,In_693,In_1819);
nor U3146 (N_3146,In_1214,In_2321);
nor U3147 (N_3147,In_2329,In_423);
and U3148 (N_3148,In_168,In_247);
nor U3149 (N_3149,In_24,In_387);
or U3150 (N_3150,In_272,In_2097);
or U3151 (N_3151,In_2248,In_1510);
and U3152 (N_3152,In_507,In_2295);
and U3153 (N_3153,In_226,In_517);
xnor U3154 (N_3154,In_381,In_1555);
and U3155 (N_3155,In_842,In_1082);
or U3156 (N_3156,In_120,In_2103);
nor U3157 (N_3157,In_1970,In_1959);
nor U3158 (N_3158,In_1952,In_457);
or U3159 (N_3159,In_2101,In_2291);
xnor U3160 (N_3160,In_2037,In_1116);
and U3161 (N_3161,In_1372,In_1860);
xnor U3162 (N_3162,In_462,In_2332);
nor U3163 (N_3163,In_1697,In_1187);
or U3164 (N_3164,In_265,In_2058);
and U3165 (N_3165,In_1237,In_2159);
or U3166 (N_3166,In_1776,In_2170);
and U3167 (N_3167,In_2007,In_592);
nand U3168 (N_3168,In_2042,In_465);
nor U3169 (N_3169,In_593,In_2134);
xor U3170 (N_3170,In_2266,In_1510);
nor U3171 (N_3171,In_305,In_2394);
nor U3172 (N_3172,In_218,In_2225);
or U3173 (N_3173,In_2308,In_457);
nor U3174 (N_3174,In_154,In_243);
nand U3175 (N_3175,In_2104,In_2310);
nand U3176 (N_3176,In_1573,In_1190);
and U3177 (N_3177,In_116,In_750);
and U3178 (N_3178,In_518,In_612);
xnor U3179 (N_3179,In_2203,In_19);
nor U3180 (N_3180,In_2313,In_259);
xnor U3181 (N_3181,In_2420,In_1054);
xnor U3182 (N_3182,In_928,In_1461);
nand U3183 (N_3183,In_2380,In_1448);
and U3184 (N_3184,In_1468,In_481);
nand U3185 (N_3185,In_1669,In_71);
xnor U3186 (N_3186,In_2245,In_1704);
xor U3187 (N_3187,In_1409,In_329);
nand U3188 (N_3188,In_2381,In_2221);
and U3189 (N_3189,In_1735,In_41);
xor U3190 (N_3190,In_1200,In_924);
or U3191 (N_3191,In_1568,In_846);
or U3192 (N_3192,In_630,In_1428);
and U3193 (N_3193,In_1397,In_2017);
and U3194 (N_3194,In_1175,In_1971);
nor U3195 (N_3195,In_1463,In_1386);
xnor U3196 (N_3196,In_1682,In_1259);
xnor U3197 (N_3197,In_1869,In_1258);
nand U3198 (N_3198,In_965,In_1009);
nand U3199 (N_3199,In_2387,In_263);
or U3200 (N_3200,In_1067,In_2291);
nor U3201 (N_3201,In_2490,In_1622);
xnor U3202 (N_3202,In_2455,In_1235);
nand U3203 (N_3203,In_1116,In_1982);
and U3204 (N_3204,In_449,In_1057);
xor U3205 (N_3205,In_2088,In_1195);
nor U3206 (N_3206,In_522,In_616);
and U3207 (N_3207,In_1882,In_1532);
or U3208 (N_3208,In_1550,In_1827);
xnor U3209 (N_3209,In_1088,In_1704);
xnor U3210 (N_3210,In_2327,In_1735);
xor U3211 (N_3211,In_1874,In_2164);
nor U3212 (N_3212,In_1208,In_1618);
nand U3213 (N_3213,In_1535,In_477);
xnor U3214 (N_3214,In_815,In_88);
xor U3215 (N_3215,In_1399,In_302);
or U3216 (N_3216,In_1885,In_1903);
nor U3217 (N_3217,In_372,In_953);
xnor U3218 (N_3218,In_755,In_1599);
xnor U3219 (N_3219,In_684,In_1970);
nor U3220 (N_3220,In_1520,In_495);
and U3221 (N_3221,In_1077,In_1937);
nor U3222 (N_3222,In_1192,In_132);
xnor U3223 (N_3223,In_736,In_1178);
or U3224 (N_3224,In_374,In_899);
and U3225 (N_3225,In_1004,In_1114);
xnor U3226 (N_3226,In_1956,In_2373);
and U3227 (N_3227,In_1309,In_1801);
or U3228 (N_3228,In_1252,In_107);
or U3229 (N_3229,In_1328,In_1063);
nor U3230 (N_3230,In_1206,In_215);
or U3231 (N_3231,In_1068,In_83);
and U3232 (N_3232,In_388,In_1018);
nand U3233 (N_3233,In_1330,In_692);
and U3234 (N_3234,In_2371,In_1643);
nand U3235 (N_3235,In_888,In_1888);
nand U3236 (N_3236,In_1135,In_2088);
xnor U3237 (N_3237,In_2087,In_1614);
nor U3238 (N_3238,In_1083,In_180);
and U3239 (N_3239,In_1660,In_1764);
or U3240 (N_3240,In_932,In_1542);
nand U3241 (N_3241,In_941,In_33);
and U3242 (N_3242,In_1933,In_1773);
nor U3243 (N_3243,In_736,In_1054);
xor U3244 (N_3244,In_1245,In_506);
and U3245 (N_3245,In_283,In_2136);
and U3246 (N_3246,In_2221,In_253);
nor U3247 (N_3247,In_596,In_760);
or U3248 (N_3248,In_322,In_1278);
nor U3249 (N_3249,In_1760,In_2437);
and U3250 (N_3250,In_1990,In_254);
and U3251 (N_3251,In_2018,In_1119);
and U3252 (N_3252,In_2438,In_910);
nor U3253 (N_3253,In_400,In_1930);
nand U3254 (N_3254,In_2464,In_494);
xnor U3255 (N_3255,In_2208,In_2023);
xnor U3256 (N_3256,In_2271,In_409);
or U3257 (N_3257,In_1914,In_1184);
or U3258 (N_3258,In_2074,In_98);
or U3259 (N_3259,In_2319,In_151);
xnor U3260 (N_3260,In_1942,In_1969);
or U3261 (N_3261,In_1907,In_987);
and U3262 (N_3262,In_2388,In_2038);
xnor U3263 (N_3263,In_824,In_1567);
nand U3264 (N_3264,In_2244,In_1673);
or U3265 (N_3265,In_2372,In_2400);
and U3266 (N_3266,In_2208,In_916);
nor U3267 (N_3267,In_1102,In_2117);
and U3268 (N_3268,In_935,In_2390);
xor U3269 (N_3269,In_1761,In_2305);
nand U3270 (N_3270,In_1163,In_191);
xor U3271 (N_3271,In_1903,In_223);
nor U3272 (N_3272,In_1267,In_2168);
nand U3273 (N_3273,In_2181,In_1900);
nand U3274 (N_3274,In_609,In_129);
and U3275 (N_3275,In_1827,In_373);
nor U3276 (N_3276,In_1117,In_1962);
or U3277 (N_3277,In_795,In_1471);
and U3278 (N_3278,In_983,In_567);
xnor U3279 (N_3279,In_1961,In_480);
and U3280 (N_3280,In_1688,In_1006);
nand U3281 (N_3281,In_770,In_1194);
or U3282 (N_3282,In_745,In_2302);
or U3283 (N_3283,In_1121,In_1475);
and U3284 (N_3284,In_447,In_2303);
and U3285 (N_3285,In_1676,In_1225);
nand U3286 (N_3286,In_1391,In_947);
nand U3287 (N_3287,In_2020,In_2127);
xor U3288 (N_3288,In_90,In_1805);
nor U3289 (N_3289,In_1282,In_114);
or U3290 (N_3290,In_189,In_2053);
nand U3291 (N_3291,In_2412,In_85);
nor U3292 (N_3292,In_1649,In_2351);
nor U3293 (N_3293,In_914,In_472);
or U3294 (N_3294,In_1405,In_454);
nand U3295 (N_3295,In_243,In_727);
and U3296 (N_3296,In_1779,In_1381);
xor U3297 (N_3297,In_172,In_1385);
nor U3298 (N_3298,In_902,In_1910);
nand U3299 (N_3299,In_1403,In_1808);
nand U3300 (N_3300,In_1205,In_392);
and U3301 (N_3301,In_1152,In_2177);
nor U3302 (N_3302,In_1340,In_2236);
xor U3303 (N_3303,In_2101,In_1756);
nor U3304 (N_3304,In_190,In_1168);
xor U3305 (N_3305,In_871,In_51);
nor U3306 (N_3306,In_1373,In_1939);
and U3307 (N_3307,In_2495,In_410);
and U3308 (N_3308,In_1589,In_1297);
or U3309 (N_3309,In_2258,In_183);
or U3310 (N_3310,In_526,In_504);
nor U3311 (N_3311,In_336,In_1133);
nor U3312 (N_3312,In_751,In_1556);
nand U3313 (N_3313,In_1428,In_2088);
and U3314 (N_3314,In_2104,In_598);
nand U3315 (N_3315,In_2219,In_411);
or U3316 (N_3316,In_1501,In_1504);
and U3317 (N_3317,In_434,In_1873);
and U3318 (N_3318,In_1616,In_991);
nand U3319 (N_3319,In_47,In_502);
nand U3320 (N_3320,In_1076,In_2293);
nand U3321 (N_3321,In_1971,In_2050);
and U3322 (N_3322,In_1424,In_2018);
or U3323 (N_3323,In_2343,In_1549);
and U3324 (N_3324,In_1536,In_826);
and U3325 (N_3325,In_582,In_1241);
nor U3326 (N_3326,In_1592,In_1534);
or U3327 (N_3327,In_2189,In_1537);
and U3328 (N_3328,In_1962,In_515);
nor U3329 (N_3329,In_1758,In_1544);
or U3330 (N_3330,In_1732,In_1218);
nand U3331 (N_3331,In_978,In_1098);
and U3332 (N_3332,In_2193,In_2107);
nor U3333 (N_3333,In_694,In_1792);
nor U3334 (N_3334,In_848,In_1858);
xor U3335 (N_3335,In_2094,In_2129);
or U3336 (N_3336,In_1448,In_1516);
or U3337 (N_3337,In_857,In_1748);
or U3338 (N_3338,In_179,In_1792);
or U3339 (N_3339,In_1893,In_2088);
xnor U3340 (N_3340,In_1493,In_1062);
xor U3341 (N_3341,In_2421,In_33);
xor U3342 (N_3342,In_1144,In_2379);
or U3343 (N_3343,In_866,In_963);
xnor U3344 (N_3344,In_1235,In_1213);
and U3345 (N_3345,In_730,In_2354);
nor U3346 (N_3346,In_1381,In_389);
xnor U3347 (N_3347,In_939,In_1224);
and U3348 (N_3348,In_766,In_2185);
or U3349 (N_3349,In_285,In_254);
nor U3350 (N_3350,In_971,In_440);
and U3351 (N_3351,In_812,In_57);
xnor U3352 (N_3352,In_169,In_718);
xor U3353 (N_3353,In_1547,In_1603);
xnor U3354 (N_3354,In_34,In_1192);
xor U3355 (N_3355,In_1082,In_849);
nor U3356 (N_3356,In_922,In_151);
nand U3357 (N_3357,In_2391,In_1984);
nor U3358 (N_3358,In_2014,In_697);
xor U3359 (N_3359,In_2374,In_2269);
nand U3360 (N_3360,In_1790,In_2331);
or U3361 (N_3361,In_1251,In_647);
nand U3362 (N_3362,In_2443,In_2108);
nand U3363 (N_3363,In_1743,In_1942);
xnor U3364 (N_3364,In_2434,In_1609);
xnor U3365 (N_3365,In_1163,In_1527);
xor U3366 (N_3366,In_882,In_2372);
xnor U3367 (N_3367,In_1592,In_773);
or U3368 (N_3368,In_485,In_632);
and U3369 (N_3369,In_604,In_1281);
and U3370 (N_3370,In_2138,In_1148);
nor U3371 (N_3371,In_1608,In_788);
nor U3372 (N_3372,In_1896,In_1256);
nor U3373 (N_3373,In_540,In_1970);
or U3374 (N_3374,In_948,In_1683);
nor U3375 (N_3375,In_2059,In_1792);
or U3376 (N_3376,In_589,In_925);
nand U3377 (N_3377,In_2300,In_103);
xor U3378 (N_3378,In_832,In_1429);
nand U3379 (N_3379,In_1613,In_238);
xnor U3380 (N_3380,In_1671,In_1788);
nor U3381 (N_3381,In_70,In_1072);
and U3382 (N_3382,In_1791,In_906);
xor U3383 (N_3383,In_440,In_1033);
or U3384 (N_3384,In_1785,In_1127);
nand U3385 (N_3385,In_72,In_1780);
nand U3386 (N_3386,In_1593,In_1257);
xnor U3387 (N_3387,In_2290,In_2328);
and U3388 (N_3388,In_81,In_100);
nor U3389 (N_3389,In_844,In_1189);
xor U3390 (N_3390,In_2249,In_2314);
or U3391 (N_3391,In_375,In_462);
nand U3392 (N_3392,In_406,In_855);
nor U3393 (N_3393,In_1821,In_1896);
xor U3394 (N_3394,In_26,In_260);
xnor U3395 (N_3395,In_1859,In_2245);
xnor U3396 (N_3396,In_1158,In_2064);
and U3397 (N_3397,In_1026,In_1192);
nand U3398 (N_3398,In_1266,In_1115);
nand U3399 (N_3399,In_687,In_2210);
or U3400 (N_3400,In_2365,In_213);
nor U3401 (N_3401,In_275,In_1737);
and U3402 (N_3402,In_1433,In_2005);
or U3403 (N_3403,In_2211,In_1381);
or U3404 (N_3404,In_2288,In_508);
xor U3405 (N_3405,In_689,In_1027);
nand U3406 (N_3406,In_1778,In_1604);
xnor U3407 (N_3407,In_1127,In_1714);
nor U3408 (N_3408,In_2413,In_1998);
xnor U3409 (N_3409,In_512,In_1922);
nor U3410 (N_3410,In_655,In_1743);
nand U3411 (N_3411,In_2321,In_1445);
or U3412 (N_3412,In_1227,In_2338);
xor U3413 (N_3413,In_1675,In_1133);
nand U3414 (N_3414,In_276,In_364);
nor U3415 (N_3415,In_636,In_2147);
nand U3416 (N_3416,In_692,In_874);
xor U3417 (N_3417,In_2246,In_462);
and U3418 (N_3418,In_1266,In_1705);
xor U3419 (N_3419,In_236,In_492);
xnor U3420 (N_3420,In_848,In_2064);
nand U3421 (N_3421,In_278,In_1958);
or U3422 (N_3422,In_2350,In_880);
nand U3423 (N_3423,In_576,In_803);
or U3424 (N_3424,In_343,In_1335);
xnor U3425 (N_3425,In_1328,In_2178);
and U3426 (N_3426,In_96,In_362);
and U3427 (N_3427,In_2394,In_1645);
and U3428 (N_3428,In_2393,In_484);
xor U3429 (N_3429,In_149,In_45);
xnor U3430 (N_3430,In_2225,In_2114);
nor U3431 (N_3431,In_109,In_1363);
nand U3432 (N_3432,In_1135,In_1087);
nand U3433 (N_3433,In_1736,In_1513);
nand U3434 (N_3434,In_1971,In_1767);
nor U3435 (N_3435,In_1055,In_282);
and U3436 (N_3436,In_2367,In_1072);
and U3437 (N_3437,In_1088,In_404);
and U3438 (N_3438,In_1076,In_21);
or U3439 (N_3439,In_1412,In_1775);
or U3440 (N_3440,In_236,In_1807);
and U3441 (N_3441,In_1878,In_556);
nor U3442 (N_3442,In_1572,In_1151);
xor U3443 (N_3443,In_2190,In_1306);
nor U3444 (N_3444,In_1295,In_319);
xor U3445 (N_3445,In_2349,In_676);
and U3446 (N_3446,In_1093,In_372);
nand U3447 (N_3447,In_852,In_2232);
xor U3448 (N_3448,In_1139,In_381);
nor U3449 (N_3449,In_1062,In_1632);
and U3450 (N_3450,In_948,In_2275);
xnor U3451 (N_3451,In_2168,In_1977);
or U3452 (N_3452,In_93,In_620);
and U3453 (N_3453,In_1635,In_362);
and U3454 (N_3454,In_1738,In_2317);
xnor U3455 (N_3455,In_1030,In_1428);
nor U3456 (N_3456,In_2327,In_15);
xor U3457 (N_3457,In_2393,In_1073);
and U3458 (N_3458,In_348,In_1124);
and U3459 (N_3459,In_2171,In_974);
or U3460 (N_3460,In_272,In_1399);
xor U3461 (N_3461,In_1296,In_323);
or U3462 (N_3462,In_534,In_188);
or U3463 (N_3463,In_926,In_1318);
nand U3464 (N_3464,In_2191,In_2208);
xnor U3465 (N_3465,In_1544,In_1472);
and U3466 (N_3466,In_1630,In_826);
and U3467 (N_3467,In_684,In_1723);
nand U3468 (N_3468,In_829,In_1780);
or U3469 (N_3469,In_2380,In_300);
nor U3470 (N_3470,In_1801,In_444);
xnor U3471 (N_3471,In_1662,In_2223);
nor U3472 (N_3472,In_730,In_700);
nor U3473 (N_3473,In_1223,In_123);
or U3474 (N_3474,In_1755,In_108);
and U3475 (N_3475,In_720,In_172);
nor U3476 (N_3476,In_2379,In_946);
nand U3477 (N_3477,In_419,In_1060);
xor U3478 (N_3478,In_1388,In_1181);
or U3479 (N_3479,In_2009,In_1565);
xor U3480 (N_3480,In_1802,In_1528);
nand U3481 (N_3481,In_1106,In_735);
xnor U3482 (N_3482,In_1022,In_144);
nand U3483 (N_3483,In_1761,In_2312);
and U3484 (N_3484,In_1019,In_293);
xnor U3485 (N_3485,In_34,In_641);
or U3486 (N_3486,In_1425,In_180);
nand U3487 (N_3487,In_1241,In_1376);
nand U3488 (N_3488,In_1150,In_756);
xnor U3489 (N_3489,In_172,In_841);
nand U3490 (N_3490,In_1849,In_661);
xnor U3491 (N_3491,In_1854,In_916);
or U3492 (N_3492,In_1116,In_437);
or U3493 (N_3493,In_659,In_1099);
and U3494 (N_3494,In_903,In_1824);
xor U3495 (N_3495,In_1805,In_2467);
xnor U3496 (N_3496,In_1949,In_2323);
nor U3497 (N_3497,In_2088,In_1665);
xor U3498 (N_3498,In_1096,In_285);
xor U3499 (N_3499,In_542,In_1499);
nand U3500 (N_3500,In_1158,In_2488);
or U3501 (N_3501,In_453,In_1286);
xor U3502 (N_3502,In_1650,In_1956);
nand U3503 (N_3503,In_1586,In_411);
nand U3504 (N_3504,In_2036,In_879);
or U3505 (N_3505,In_1609,In_1561);
nand U3506 (N_3506,In_676,In_1190);
nand U3507 (N_3507,In_746,In_1665);
and U3508 (N_3508,In_404,In_2205);
nor U3509 (N_3509,In_1314,In_2312);
nor U3510 (N_3510,In_53,In_1860);
and U3511 (N_3511,In_58,In_2173);
and U3512 (N_3512,In_1300,In_662);
and U3513 (N_3513,In_1721,In_2003);
nand U3514 (N_3514,In_1494,In_2495);
xor U3515 (N_3515,In_1025,In_1501);
nor U3516 (N_3516,In_638,In_808);
xnor U3517 (N_3517,In_611,In_1136);
and U3518 (N_3518,In_943,In_1250);
or U3519 (N_3519,In_1761,In_1341);
nand U3520 (N_3520,In_2212,In_549);
nand U3521 (N_3521,In_1756,In_541);
nor U3522 (N_3522,In_1130,In_1926);
or U3523 (N_3523,In_1542,In_1368);
nand U3524 (N_3524,In_807,In_503);
xnor U3525 (N_3525,In_528,In_2350);
and U3526 (N_3526,In_1730,In_1887);
or U3527 (N_3527,In_2037,In_646);
or U3528 (N_3528,In_408,In_338);
nand U3529 (N_3529,In_436,In_1939);
or U3530 (N_3530,In_1926,In_2283);
and U3531 (N_3531,In_380,In_1499);
nand U3532 (N_3532,In_2004,In_1532);
nor U3533 (N_3533,In_382,In_2167);
xnor U3534 (N_3534,In_1563,In_1394);
and U3535 (N_3535,In_1042,In_1054);
and U3536 (N_3536,In_2210,In_2065);
nor U3537 (N_3537,In_2243,In_393);
xnor U3538 (N_3538,In_723,In_2344);
xnor U3539 (N_3539,In_2052,In_12);
nand U3540 (N_3540,In_706,In_1691);
or U3541 (N_3541,In_255,In_1365);
or U3542 (N_3542,In_116,In_1689);
and U3543 (N_3543,In_1389,In_27);
xor U3544 (N_3544,In_1568,In_2322);
nand U3545 (N_3545,In_1467,In_2215);
and U3546 (N_3546,In_1047,In_833);
and U3547 (N_3547,In_995,In_1963);
xor U3548 (N_3548,In_567,In_1363);
xor U3549 (N_3549,In_257,In_1253);
xor U3550 (N_3550,In_58,In_1448);
or U3551 (N_3551,In_2185,In_53);
and U3552 (N_3552,In_126,In_575);
xnor U3553 (N_3553,In_906,In_374);
nand U3554 (N_3554,In_1006,In_1816);
xnor U3555 (N_3555,In_636,In_1160);
nand U3556 (N_3556,In_755,In_278);
and U3557 (N_3557,In_2221,In_475);
xor U3558 (N_3558,In_1674,In_963);
and U3559 (N_3559,In_2146,In_1775);
xor U3560 (N_3560,In_1234,In_618);
xnor U3561 (N_3561,In_2405,In_882);
xor U3562 (N_3562,In_2415,In_449);
nand U3563 (N_3563,In_987,In_5);
nor U3564 (N_3564,In_2179,In_1995);
or U3565 (N_3565,In_2436,In_673);
nor U3566 (N_3566,In_398,In_293);
nor U3567 (N_3567,In_827,In_1261);
nand U3568 (N_3568,In_1008,In_266);
and U3569 (N_3569,In_23,In_1682);
and U3570 (N_3570,In_372,In_1705);
nand U3571 (N_3571,In_812,In_582);
xor U3572 (N_3572,In_59,In_1146);
or U3573 (N_3573,In_1584,In_3);
or U3574 (N_3574,In_4,In_1388);
or U3575 (N_3575,In_1523,In_2351);
nor U3576 (N_3576,In_222,In_335);
and U3577 (N_3577,In_1755,In_770);
or U3578 (N_3578,In_2344,In_1908);
xor U3579 (N_3579,In_905,In_1695);
or U3580 (N_3580,In_859,In_781);
xnor U3581 (N_3581,In_1742,In_1127);
nor U3582 (N_3582,In_1984,In_2203);
or U3583 (N_3583,In_583,In_1513);
or U3584 (N_3584,In_403,In_995);
xor U3585 (N_3585,In_46,In_938);
nand U3586 (N_3586,In_1802,In_516);
nand U3587 (N_3587,In_330,In_851);
nand U3588 (N_3588,In_1498,In_622);
nand U3589 (N_3589,In_2365,In_1476);
xnor U3590 (N_3590,In_1186,In_865);
and U3591 (N_3591,In_1166,In_1009);
xnor U3592 (N_3592,In_1217,In_451);
and U3593 (N_3593,In_871,In_387);
or U3594 (N_3594,In_255,In_2266);
nor U3595 (N_3595,In_728,In_2098);
nor U3596 (N_3596,In_1969,In_614);
xor U3597 (N_3597,In_2243,In_939);
nor U3598 (N_3598,In_537,In_569);
nor U3599 (N_3599,In_1705,In_1341);
nor U3600 (N_3600,In_1288,In_1318);
xor U3601 (N_3601,In_2278,In_989);
nand U3602 (N_3602,In_843,In_316);
or U3603 (N_3603,In_2037,In_2461);
nor U3604 (N_3604,In_920,In_1297);
xnor U3605 (N_3605,In_2296,In_578);
or U3606 (N_3606,In_1661,In_2096);
and U3607 (N_3607,In_383,In_2359);
xor U3608 (N_3608,In_1137,In_1913);
or U3609 (N_3609,In_748,In_1124);
nand U3610 (N_3610,In_1635,In_471);
or U3611 (N_3611,In_492,In_1575);
nand U3612 (N_3612,In_2109,In_2451);
and U3613 (N_3613,In_1838,In_1290);
xnor U3614 (N_3614,In_1154,In_732);
xor U3615 (N_3615,In_379,In_170);
nand U3616 (N_3616,In_2370,In_1448);
nor U3617 (N_3617,In_2440,In_488);
xnor U3618 (N_3618,In_2178,In_1160);
nand U3619 (N_3619,In_1262,In_1610);
xor U3620 (N_3620,In_1024,In_1409);
or U3621 (N_3621,In_1985,In_963);
xnor U3622 (N_3622,In_864,In_765);
xnor U3623 (N_3623,In_927,In_1105);
or U3624 (N_3624,In_680,In_1523);
and U3625 (N_3625,In_1527,In_809);
nand U3626 (N_3626,In_126,In_362);
xnor U3627 (N_3627,In_1710,In_1150);
and U3628 (N_3628,In_144,In_2257);
xnor U3629 (N_3629,In_99,In_1265);
or U3630 (N_3630,In_2260,In_1303);
or U3631 (N_3631,In_2355,In_301);
nor U3632 (N_3632,In_97,In_1234);
nand U3633 (N_3633,In_1643,In_1161);
and U3634 (N_3634,In_907,In_164);
nand U3635 (N_3635,In_2329,In_1559);
nand U3636 (N_3636,In_1045,In_1051);
xor U3637 (N_3637,In_1959,In_597);
nor U3638 (N_3638,In_1204,In_1485);
or U3639 (N_3639,In_965,In_1565);
nor U3640 (N_3640,In_1535,In_2079);
nor U3641 (N_3641,In_1307,In_2057);
nor U3642 (N_3642,In_71,In_1972);
xnor U3643 (N_3643,In_1286,In_14);
nor U3644 (N_3644,In_1023,In_328);
nand U3645 (N_3645,In_1102,In_42);
nand U3646 (N_3646,In_1325,In_1914);
xnor U3647 (N_3647,In_2160,In_1801);
or U3648 (N_3648,In_1717,In_1945);
or U3649 (N_3649,In_556,In_445);
xor U3650 (N_3650,In_2305,In_2018);
or U3651 (N_3651,In_317,In_1878);
or U3652 (N_3652,In_70,In_1861);
nor U3653 (N_3653,In_1876,In_2129);
nor U3654 (N_3654,In_480,In_20);
or U3655 (N_3655,In_2414,In_635);
nand U3656 (N_3656,In_394,In_1800);
nand U3657 (N_3657,In_330,In_26);
and U3658 (N_3658,In_2060,In_715);
and U3659 (N_3659,In_981,In_954);
nor U3660 (N_3660,In_1460,In_35);
and U3661 (N_3661,In_2295,In_814);
nor U3662 (N_3662,In_437,In_434);
and U3663 (N_3663,In_678,In_1055);
xnor U3664 (N_3664,In_1993,In_2372);
xnor U3665 (N_3665,In_630,In_2350);
xnor U3666 (N_3666,In_451,In_1042);
and U3667 (N_3667,In_1297,In_543);
nand U3668 (N_3668,In_1407,In_135);
and U3669 (N_3669,In_1625,In_2328);
nor U3670 (N_3670,In_411,In_172);
or U3671 (N_3671,In_139,In_611);
nor U3672 (N_3672,In_1112,In_1420);
xor U3673 (N_3673,In_621,In_1120);
xor U3674 (N_3674,In_476,In_687);
nand U3675 (N_3675,In_742,In_1393);
and U3676 (N_3676,In_1950,In_1121);
nand U3677 (N_3677,In_922,In_1051);
and U3678 (N_3678,In_1970,In_897);
nand U3679 (N_3679,In_2181,In_1246);
xnor U3680 (N_3680,In_1345,In_1908);
nor U3681 (N_3681,In_1993,In_1298);
or U3682 (N_3682,In_615,In_1774);
or U3683 (N_3683,In_1383,In_2214);
or U3684 (N_3684,In_1472,In_629);
nand U3685 (N_3685,In_1539,In_1444);
and U3686 (N_3686,In_656,In_553);
or U3687 (N_3687,In_340,In_1339);
nand U3688 (N_3688,In_704,In_2200);
xnor U3689 (N_3689,In_1182,In_2112);
nand U3690 (N_3690,In_336,In_514);
and U3691 (N_3691,In_772,In_2379);
xnor U3692 (N_3692,In_1777,In_1896);
nand U3693 (N_3693,In_1130,In_639);
or U3694 (N_3694,In_730,In_1242);
nand U3695 (N_3695,In_1479,In_18);
nor U3696 (N_3696,In_1177,In_2189);
nor U3697 (N_3697,In_997,In_2469);
xnor U3698 (N_3698,In_1694,In_1168);
or U3699 (N_3699,In_2172,In_1002);
or U3700 (N_3700,In_1083,In_1903);
nand U3701 (N_3701,In_259,In_831);
nand U3702 (N_3702,In_109,In_2299);
xor U3703 (N_3703,In_1571,In_2257);
xnor U3704 (N_3704,In_711,In_1707);
and U3705 (N_3705,In_9,In_792);
nor U3706 (N_3706,In_2475,In_2008);
nand U3707 (N_3707,In_746,In_391);
xnor U3708 (N_3708,In_1063,In_656);
or U3709 (N_3709,In_2136,In_904);
xnor U3710 (N_3710,In_1752,In_1973);
and U3711 (N_3711,In_1732,In_1486);
xor U3712 (N_3712,In_1909,In_2089);
nand U3713 (N_3713,In_2063,In_88);
and U3714 (N_3714,In_200,In_399);
or U3715 (N_3715,In_469,In_742);
nor U3716 (N_3716,In_161,In_1170);
and U3717 (N_3717,In_997,In_2310);
xor U3718 (N_3718,In_974,In_1604);
xnor U3719 (N_3719,In_245,In_1251);
or U3720 (N_3720,In_513,In_2274);
and U3721 (N_3721,In_1778,In_2123);
or U3722 (N_3722,In_1171,In_671);
xor U3723 (N_3723,In_2322,In_771);
or U3724 (N_3724,In_136,In_1758);
and U3725 (N_3725,In_1949,In_204);
xor U3726 (N_3726,In_2028,In_224);
or U3727 (N_3727,In_964,In_1726);
nand U3728 (N_3728,In_414,In_1225);
or U3729 (N_3729,In_787,In_168);
xor U3730 (N_3730,In_22,In_710);
nand U3731 (N_3731,In_2441,In_1127);
or U3732 (N_3732,In_974,In_1426);
nor U3733 (N_3733,In_2396,In_2373);
nor U3734 (N_3734,In_2483,In_770);
or U3735 (N_3735,In_1851,In_1565);
nand U3736 (N_3736,In_2496,In_1789);
nand U3737 (N_3737,In_1389,In_2428);
or U3738 (N_3738,In_1454,In_584);
nand U3739 (N_3739,In_109,In_1848);
xnor U3740 (N_3740,In_1060,In_626);
nor U3741 (N_3741,In_674,In_1645);
nand U3742 (N_3742,In_142,In_2296);
xnor U3743 (N_3743,In_490,In_481);
xnor U3744 (N_3744,In_581,In_1008);
or U3745 (N_3745,In_774,In_849);
and U3746 (N_3746,In_1632,In_799);
nor U3747 (N_3747,In_1414,In_158);
xnor U3748 (N_3748,In_1893,In_1965);
or U3749 (N_3749,In_1750,In_1953);
xor U3750 (N_3750,In_33,In_1682);
nor U3751 (N_3751,In_768,In_1169);
nand U3752 (N_3752,In_2343,In_221);
and U3753 (N_3753,In_243,In_503);
and U3754 (N_3754,In_2345,In_56);
nor U3755 (N_3755,In_895,In_2216);
xnor U3756 (N_3756,In_1540,In_2403);
or U3757 (N_3757,In_2119,In_0);
xnor U3758 (N_3758,In_319,In_245);
and U3759 (N_3759,In_1426,In_1397);
xor U3760 (N_3760,In_2378,In_653);
and U3761 (N_3761,In_1155,In_724);
and U3762 (N_3762,In_826,In_1521);
or U3763 (N_3763,In_17,In_1804);
nor U3764 (N_3764,In_499,In_1559);
nand U3765 (N_3765,In_303,In_1871);
or U3766 (N_3766,In_1478,In_2184);
nor U3767 (N_3767,In_1173,In_1183);
xnor U3768 (N_3768,In_974,In_1213);
nand U3769 (N_3769,In_2453,In_1234);
xnor U3770 (N_3770,In_1486,In_2440);
or U3771 (N_3771,In_1873,In_208);
xor U3772 (N_3772,In_1999,In_1162);
nand U3773 (N_3773,In_589,In_1450);
or U3774 (N_3774,In_989,In_2338);
xor U3775 (N_3775,In_79,In_1395);
nand U3776 (N_3776,In_1509,In_1926);
nand U3777 (N_3777,In_1665,In_419);
nor U3778 (N_3778,In_2198,In_1064);
nor U3779 (N_3779,In_2459,In_869);
nand U3780 (N_3780,In_139,In_657);
nand U3781 (N_3781,In_187,In_1304);
nor U3782 (N_3782,In_1465,In_2247);
nor U3783 (N_3783,In_2306,In_1329);
xnor U3784 (N_3784,In_1845,In_2251);
and U3785 (N_3785,In_223,In_2014);
nand U3786 (N_3786,In_395,In_1925);
or U3787 (N_3787,In_1088,In_1800);
xor U3788 (N_3788,In_1660,In_1245);
nor U3789 (N_3789,In_68,In_2113);
nand U3790 (N_3790,In_229,In_697);
nor U3791 (N_3791,In_2102,In_336);
and U3792 (N_3792,In_2429,In_1075);
nor U3793 (N_3793,In_1332,In_625);
xnor U3794 (N_3794,In_1430,In_994);
nand U3795 (N_3795,In_2020,In_645);
and U3796 (N_3796,In_1433,In_1977);
nand U3797 (N_3797,In_1312,In_1814);
or U3798 (N_3798,In_373,In_217);
and U3799 (N_3799,In_281,In_638);
or U3800 (N_3800,In_876,In_2307);
nor U3801 (N_3801,In_751,In_1570);
xor U3802 (N_3802,In_165,In_577);
xnor U3803 (N_3803,In_1213,In_74);
xor U3804 (N_3804,In_2232,In_1857);
xor U3805 (N_3805,In_2091,In_952);
or U3806 (N_3806,In_2365,In_2011);
and U3807 (N_3807,In_1296,In_2357);
nor U3808 (N_3808,In_2347,In_62);
nor U3809 (N_3809,In_1143,In_267);
and U3810 (N_3810,In_1688,In_2058);
nor U3811 (N_3811,In_287,In_1348);
nor U3812 (N_3812,In_98,In_1902);
and U3813 (N_3813,In_611,In_322);
nand U3814 (N_3814,In_2230,In_2057);
and U3815 (N_3815,In_1876,In_1794);
xnor U3816 (N_3816,In_2415,In_1622);
nor U3817 (N_3817,In_467,In_2433);
xor U3818 (N_3818,In_325,In_1165);
and U3819 (N_3819,In_1369,In_2437);
nand U3820 (N_3820,In_255,In_963);
nor U3821 (N_3821,In_2469,In_2007);
nand U3822 (N_3822,In_1231,In_50);
and U3823 (N_3823,In_1965,In_559);
or U3824 (N_3824,In_1317,In_1634);
nor U3825 (N_3825,In_180,In_1089);
nor U3826 (N_3826,In_314,In_576);
xor U3827 (N_3827,In_350,In_5);
nand U3828 (N_3828,In_978,In_1076);
xor U3829 (N_3829,In_1175,In_846);
xor U3830 (N_3830,In_1878,In_367);
or U3831 (N_3831,In_912,In_505);
nor U3832 (N_3832,In_331,In_957);
nor U3833 (N_3833,In_2012,In_1675);
xor U3834 (N_3834,In_2376,In_1829);
or U3835 (N_3835,In_462,In_2466);
nor U3836 (N_3836,In_242,In_1565);
and U3837 (N_3837,In_1467,In_756);
or U3838 (N_3838,In_1653,In_1874);
xor U3839 (N_3839,In_1814,In_497);
nor U3840 (N_3840,In_2140,In_1755);
nor U3841 (N_3841,In_1320,In_389);
nand U3842 (N_3842,In_62,In_2418);
or U3843 (N_3843,In_767,In_466);
nand U3844 (N_3844,In_131,In_1245);
nand U3845 (N_3845,In_169,In_1246);
and U3846 (N_3846,In_2293,In_1287);
nand U3847 (N_3847,In_1027,In_748);
nand U3848 (N_3848,In_925,In_341);
or U3849 (N_3849,In_334,In_1632);
xnor U3850 (N_3850,In_2007,In_1385);
nor U3851 (N_3851,In_1960,In_751);
xnor U3852 (N_3852,In_862,In_295);
nand U3853 (N_3853,In_2272,In_1508);
and U3854 (N_3854,In_431,In_1892);
or U3855 (N_3855,In_729,In_1839);
nor U3856 (N_3856,In_870,In_553);
or U3857 (N_3857,In_360,In_2166);
xor U3858 (N_3858,In_570,In_697);
and U3859 (N_3859,In_1122,In_775);
nand U3860 (N_3860,In_1722,In_2384);
nand U3861 (N_3861,In_2306,In_1008);
xor U3862 (N_3862,In_934,In_1651);
nand U3863 (N_3863,In_1709,In_2286);
nand U3864 (N_3864,In_154,In_1041);
xnor U3865 (N_3865,In_777,In_1659);
nand U3866 (N_3866,In_350,In_1256);
nand U3867 (N_3867,In_251,In_2220);
xor U3868 (N_3868,In_2253,In_1617);
nor U3869 (N_3869,In_2050,In_2241);
nor U3870 (N_3870,In_439,In_2354);
or U3871 (N_3871,In_1420,In_801);
and U3872 (N_3872,In_1117,In_1621);
nand U3873 (N_3873,In_1200,In_257);
or U3874 (N_3874,In_1103,In_2201);
nand U3875 (N_3875,In_1808,In_174);
nor U3876 (N_3876,In_368,In_2482);
nand U3877 (N_3877,In_2072,In_145);
nand U3878 (N_3878,In_961,In_1525);
nor U3879 (N_3879,In_1578,In_1030);
or U3880 (N_3880,In_918,In_1158);
nand U3881 (N_3881,In_1661,In_2020);
or U3882 (N_3882,In_71,In_513);
xnor U3883 (N_3883,In_1838,In_728);
nor U3884 (N_3884,In_1775,In_220);
nor U3885 (N_3885,In_1148,In_572);
nand U3886 (N_3886,In_848,In_1339);
xor U3887 (N_3887,In_2414,In_256);
or U3888 (N_3888,In_1621,In_1541);
nand U3889 (N_3889,In_2401,In_86);
nor U3890 (N_3890,In_1923,In_1798);
nor U3891 (N_3891,In_987,In_2208);
nor U3892 (N_3892,In_46,In_617);
xor U3893 (N_3893,In_1680,In_2471);
xnor U3894 (N_3894,In_1891,In_1842);
or U3895 (N_3895,In_2065,In_865);
or U3896 (N_3896,In_2112,In_2190);
xnor U3897 (N_3897,In_1487,In_2222);
or U3898 (N_3898,In_646,In_2281);
nand U3899 (N_3899,In_1771,In_2439);
xor U3900 (N_3900,In_524,In_2083);
xor U3901 (N_3901,In_420,In_650);
nor U3902 (N_3902,In_884,In_1059);
or U3903 (N_3903,In_1995,In_2372);
nand U3904 (N_3904,In_1322,In_1926);
and U3905 (N_3905,In_1177,In_1830);
nor U3906 (N_3906,In_82,In_321);
nor U3907 (N_3907,In_1286,In_1477);
nor U3908 (N_3908,In_1796,In_1246);
xor U3909 (N_3909,In_652,In_2358);
xor U3910 (N_3910,In_1541,In_470);
nor U3911 (N_3911,In_222,In_1416);
and U3912 (N_3912,In_2335,In_1843);
and U3913 (N_3913,In_2243,In_900);
nor U3914 (N_3914,In_2085,In_2046);
xor U3915 (N_3915,In_10,In_2117);
nand U3916 (N_3916,In_2364,In_1793);
nand U3917 (N_3917,In_152,In_1208);
and U3918 (N_3918,In_40,In_405);
nand U3919 (N_3919,In_773,In_998);
nor U3920 (N_3920,In_234,In_1504);
nand U3921 (N_3921,In_1578,In_2043);
xnor U3922 (N_3922,In_1472,In_2254);
nand U3923 (N_3923,In_1023,In_823);
and U3924 (N_3924,In_1471,In_1676);
or U3925 (N_3925,In_2499,In_902);
or U3926 (N_3926,In_2057,In_174);
nor U3927 (N_3927,In_929,In_1494);
nand U3928 (N_3928,In_2184,In_1519);
xnor U3929 (N_3929,In_2087,In_2097);
nand U3930 (N_3930,In_895,In_239);
or U3931 (N_3931,In_390,In_1);
and U3932 (N_3932,In_2203,In_1126);
or U3933 (N_3933,In_1981,In_294);
xor U3934 (N_3934,In_535,In_863);
or U3935 (N_3935,In_1299,In_2470);
nand U3936 (N_3936,In_628,In_421);
xnor U3937 (N_3937,In_2220,In_2077);
nor U3938 (N_3938,In_1182,In_1787);
and U3939 (N_3939,In_1589,In_1571);
or U3940 (N_3940,In_243,In_1828);
nand U3941 (N_3941,In_1393,In_1281);
and U3942 (N_3942,In_2491,In_1657);
nand U3943 (N_3943,In_1868,In_19);
xnor U3944 (N_3944,In_87,In_1624);
nor U3945 (N_3945,In_2287,In_2147);
and U3946 (N_3946,In_2208,In_773);
or U3947 (N_3947,In_1568,In_752);
nor U3948 (N_3948,In_1347,In_1043);
nor U3949 (N_3949,In_1716,In_1270);
or U3950 (N_3950,In_401,In_774);
nand U3951 (N_3951,In_132,In_2225);
and U3952 (N_3952,In_2222,In_388);
or U3953 (N_3953,In_2064,In_89);
and U3954 (N_3954,In_2227,In_1100);
nor U3955 (N_3955,In_739,In_2124);
or U3956 (N_3956,In_1976,In_1328);
nand U3957 (N_3957,In_1106,In_2379);
nor U3958 (N_3958,In_1432,In_1210);
nor U3959 (N_3959,In_1364,In_1402);
and U3960 (N_3960,In_1311,In_543);
nand U3961 (N_3961,In_1601,In_1481);
xor U3962 (N_3962,In_928,In_2254);
xor U3963 (N_3963,In_1739,In_1138);
xor U3964 (N_3964,In_2072,In_1026);
and U3965 (N_3965,In_366,In_1076);
xor U3966 (N_3966,In_1096,In_1744);
and U3967 (N_3967,In_2403,In_809);
and U3968 (N_3968,In_1763,In_1397);
xor U3969 (N_3969,In_823,In_1227);
and U3970 (N_3970,In_1754,In_1492);
nor U3971 (N_3971,In_308,In_1592);
nor U3972 (N_3972,In_1639,In_1642);
nor U3973 (N_3973,In_312,In_972);
nor U3974 (N_3974,In_2147,In_488);
xnor U3975 (N_3975,In_1215,In_474);
and U3976 (N_3976,In_944,In_64);
xor U3977 (N_3977,In_749,In_2233);
nand U3978 (N_3978,In_281,In_1151);
and U3979 (N_3979,In_297,In_312);
or U3980 (N_3980,In_558,In_2227);
or U3981 (N_3981,In_2209,In_1687);
or U3982 (N_3982,In_1656,In_2018);
nand U3983 (N_3983,In_1287,In_283);
or U3984 (N_3984,In_541,In_2498);
and U3985 (N_3985,In_752,In_475);
and U3986 (N_3986,In_1606,In_1873);
xor U3987 (N_3987,In_1580,In_1315);
nand U3988 (N_3988,In_7,In_2189);
xnor U3989 (N_3989,In_1096,In_1416);
and U3990 (N_3990,In_9,In_1423);
xnor U3991 (N_3991,In_1300,In_1441);
nand U3992 (N_3992,In_2052,In_1036);
and U3993 (N_3993,In_2468,In_148);
nand U3994 (N_3994,In_1156,In_1115);
and U3995 (N_3995,In_857,In_246);
nand U3996 (N_3996,In_1461,In_436);
or U3997 (N_3997,In_1060,In_1382);
xnor U3998 (N_3998,In_1752,In_1293);
xor U3999 (N_3999,In_2010,In_2265);
nor U4000 (N_4000,In_1252,In_1089);
nand U4001 (N_4001,In_931,In_2113);
nor U4002 (N_4002,In_2487,In_856);
or U4003 (N_4003,In_1630,In_1296);
and U4004 (N_4004,In_846,In_64);
xor U4005 (N_4005,In_1250,In_929);
nor U4006 (N_4006,In_1108,In_2047);
nor U4007 (N_4007,In_2127,In_913);
and U4008 (N_4008,In_1169,In_1248);
or U4009 (N_4009,In_2176,In_2472);
nand U4010 (N_4010,In_1644,In_784);
nand U4011 (N_4011,In_479,In_495);
nor U4012 (N_4012,In_2197,In_110);
nand U4013 (N_4013,In_227,In_192);
or U4014 (N_4014,In_2190,In_984);
and U4015 (N_4015,In_2008,In_740);
xor U4016 (N_4016,In_450,In_1876);
nand U4017 (N_4017,In_2228,In_581);
xor U4018 (N_4018,In_843,In_180);
nor U4019 (N_4019,In_670,In_872);
xor U4020 (N_4020,In_102,In_2179);
nand U4021 (N_4021,In_1709,In_782);
xnor U4022 (N_4022,In_1174,In_1827);
nor U4023 (N_4023,In_2264,In_1821);
or U4024 (N_4024,In_1409,In_1298);
or U4025 (N_4025,In_1247,In_774);
nor U4026 (N_4026,In_1149,In_1683);
nand U4027 (N_4027,In_1413,In_2285);
xnor U4028 (N_4028,In_400,In_2012);
nand U4029 (N_4029,In_1063,In_1975);
and U4030 (N_4030,In_913,In_427);
xnor U4031 (N_4031,In_2079,In_1892);
or U4032 (N_4032,In_616,In_1334);
xnor U4033 (N_4033,In_1326,In_1007);
xor U4034 (N_4034,In_2299,In_925);
xnor U4035 (N_4035,In_301,In_314);
nand U4036 (N_4036,In_1543,In_662);
nor U4037 (N_4037,In_1657,In_974);
xor U4038 (N_4038,In_840,In_1158);
nor U4039 (N_4039,In_1992,In_1440);
nand U4040 (N_4040,In_300,In_788);
or U4041 (N_4041,In_1353,In_2056);
or U4042 (N_4042,In_1000,In_2003);
xor U4043 (N_4043,In_1961,In_1465);
and U4044 (N_4044,In_979,In_808);
nor U4045 (N_4045,In_445,In_1213);
nand U4046 (N_4046,In_1544,In_2092);
and U4047 (N_4047,In_144,In_684);
and U4048 (N_4048,In_245,In_2074);
or U4049 (N_4049,In_1203,In_2348);
nand U4050 (N_4050,In_2177,In_2456);
xor U4051 (N_4051,In_1746,In_2196);
or U4052 (N_4052,In_701,In_1167);
nor U4053 (N_4053,In_352,In_33);
and U4054 (N_4054,In_1625,In_2091);
nand U4055 (N_4055,In_2471,In_394);
or U4056 (N_4056,In_1603,In_305);
or U4057 (N_4057,In_1060,In_1936);
or U4058 (N_4058,In_2076,In_1115);
or U4059 (N_4059,In_595,In_1513);
nand U4060 (N_4060,In_727,In_1199);
nand U4061 (N_4061,In_898,In_1770);
and U4062 (N_4062,In_544,In_516);
or U4063 (N_4063,In_2080,In_1232);
and U4064 (N_4064,In_481,In_2486);
or U4065 (N_4065,In_541,In_2031);
and U4066 (N_4066,In_594,In_1152);
or U4067 (N_4067,In_2246,In_1447);
xor U4068 (N_4068,In_1038,In_1860);
xnor U4069 (N_4069,In_779,In_1605);
xnor U4070 (N_4070,In_2235,In_1430);
nand U4071 (N_4071,In_2267,In_1109);
xnor U4072 (N_4072,In_932,In_563);
nand U4073 (N_4073,In_2284,In_1633);
xnor U4074 (N_4074,In_1234,In_990);
nand U4075 (N_4075,In_1923,In_2230);
and U4076 (N_4076,In_1854,In_1909);
nor U4077 (N_4077,In_2089,In_1651);
nand U4078 (N_4078,In_2406,In_1404);
xnor U4079 (N_4079,In_1711,In_2074);
nand U4080 (N_4080,In_1618,In_770);
xnor U4081 (N_4081,In_1403,In_313);
nor U4082 (N_4082,In_2317,In_577);
nand U4083 (N_4083,In_1178,In_2240);
nand U4084 (N_4084,In_648,In_2194);
nand U4085 (N_4085,In_259,In_317);
or U4086 (N_4086,In_1987,In_1575);
xor U4087 (N_4087,In_1910,In_2195);
and U4088 (N_4088,In_1658,In_914);
and U4089 (N_4089,In_2077,In_626);
xnor U4090 (N_4090,In_947,In_1886);
nor U4091 (N_4091,In_1402,In_1064);
and U4092 (N_4092,In_985,In_552);
nor U4093 (N_4093,In_745,In_1425);
nor U4094 (N_4094,In_246,In_158);
xnor U4095 (N_4095,In_1933,In_600);
nor U4096 (N_4096,In_900,In_1281);
or U4097 (N_4097,In_285,In_2400);
nand U4098 (N_4098,In_1417,In_249);
nand U4099 (N_4099,In_45,In_103);
nor U4100 (N_4100,In_472,In_916);
nor U4101 (N_4101,In_2219,In_1916);
xnor U4102 (N_4102,In_1728,In_2128);
and U4103 (N_4103,In_1345,In_1334);
nand U4104 (N_4104,In_1304,In_2444);
nor U4105 (N_4105,In_2370,In_853);
nor U4106 (N_4106,In_469,In_1524);
xor U4107 (N_4107,In_975,In_1508);
or U4108 (N_4108,In_1022,In_1874);
or U4109 (N_4109,In_297,In_1090);
xor U4110 (N_4110,In_702,In_837);
nor U4111 (N_4111,In_30,In_1681);
or U4112 (N_4112,In_1742,In_1294);
or U4113 (N_4113,In_1491,In_839);
nor U4114 (N_4114,In_595,In_482);
nand U4115 (N_4115,In_399,In_577);
nand U4116 (N_4116,In_1305,In_1430);
and U4117 (N_4117,In_1263,In_1325);
xnor U4118 (N_4118,In_215,In_255);
or U4119 (N_4119,In_1187,In_434);
nand U4120 (N_4120,In_1323,In_1754);
xor U4121 (N_4121,In_1540,In_1775);
xor U4122 (N_4122,In_1415,In_462);
xnor U4123 (N_4123,In_891,In_2497);
nor U4124 (N_4124,In_1549,In_781);
or U4125 (N_4125,In_2457,In_1735);
or U4126 (N_4126,In_88,In_2479);
and U4127 (N_4127,In_2406,In_1312);
or U4128 (N_4128,In_1872,In_1110);
xnor U4129 (N_4129,In_2158,In_1019);
or U4130 (N_4130,In_196,In_1955);
nor U4131 (N_4131,In_2027,In_2367);
nor U4132 (N_4132,In_1617,In_2219);
and U4133 (N_4133,In_2037,In_1187);
and U4134 (N_4134,In_829,In_1597);
and U4135 (N_4135,In_348,In_1537);
nand U4136 (N_4136,In_698,In_1659);
or U4137 (N_4137,In_2103,In_1457);
xnor U4138 (N_4138,In_566,In_1139);
and U4139 (N_4139,In_727,In_31);
nor U4140 (N_4140,In_859,In_2071);
nand U4141 (N_4141,In_2348,In_815);
xor U4142 (N_4142,In_1562,In_2092);
or U4143 (N_4143,In_573,In_101);
nand U4144 (N_4144,In_2394,In_1493);
or U4145 (N_4145,In_982,In_961);
nor U4146 (N_4146,In_1270,In_1971);
and U4147 (N_4147,In_2149,In_1344);
or U4148 (N_4148,In_2444,In_47);
and U4149 (N_4149,In_851,In_2321);
nor U4150 (N_4150,In_981,In_2104);
nor U4151 (N_4151,In_1406,In_166);
and U4152 (N_4152,In_2091,In_1001);
xor U4153 (N_4153,In_1226,In_2055);
nand U4154 (N_4154,In_1732,In_1573);
and U4155 (N_4155,In_940,In_442);
xnor U4156 (N_4156,In_1775,In_1663);
nor U4157 (N_4157,In_2169,In_38);
nor U4158 (N_4158,In_1152,In_1434);
nor U4159 (N_4159,In_1728,In_191);
or U4160 (N_4160,In_1936,In_143);
xor U4161 (N_4161,In_1044,In_677);
or U4162 (N_4162,In_1711,In_813);
or U4163 (N_4163,In_2460,In_63);
nor U4164 (N_4164,In_929,In_1235);
and U4165 (N_4165,In_566,In_139);
and U4166 (N_4166,In_413,In_1275);
xor U4167 (N_4167,In_1196,In_684);
xnor U4168 (N_4168,In_2081,In_961);
xor U4169 (N_4169,In_2282,In_1585);
nor U4170 (N_4170,In_1623,In_1670);
nor U4171 (N_4171,In_1590,In_1462);
nor U4172 (N_4172,In_2215,In_1097);
or U4173 (N_4173,In_315,In_39);
nor U4174 (N_4174,In_1980,In_1552);
nor U4175 (N_4175,In_890,In_696);
nand U4176 (N_4176,In_1643,In_269);
or U4177 (N_4177,In_1275,In_1174);
xnor U4178 (N_4178,In_1131,In_1371);
xnor U4179 (N_4179,In_643,In_1184);
or U4180 (N_4180,In_1760,In_944);
nand U4181 (N_4181,In_525,In_1138);
xnor U4182 (N_4182,In_2169,In_1533);
or U4183 (N_4183,In_2198,In_704);
and U4184 (N_4184,In_1927,In_1364);
nand U4185 (N_4185,In_2347,In_903);
xor U4186 (N_4186,In_1966,In_706);
and U4187 (N_4187,In_2140,In_276);
nand U4188 (N_4188,In_79,In_1119);
nand U4189 (N_4189,In_1655,In_1995);
or U4190 (N_4190,In_114,In_639);
and U4191 (N_4191,In_986,In_2097);
xor U4192 (N_4192,In_1346,In_1292);
xor U4193 (N_4193,In_623,In_2425);
and U4194 (N_4194,In_1332,In_1300);
nor U4195 (N_4195,In_1087,In_1454);
xnor U4196 (N_4196,In_446,In_2187);
nand U4197 (N_4197,In_407,In_1590);
nor U4198 (N_4198,In_661,In_2187);
nand U4199 (N_4199,In_2258,In_1399);
xnor U4200 (N_4200,In_755,In_1641);
nor U4201 (N_4201,In_704,In_2403);
and U4202 (N_4202,In_244,In_1601);
or U4203 (N_4203,In_2405,In_1930);
and U4204 (N_4204,In_1321,In_541);
nand U4205 (N_4205,In_968,In_1058);
or U4206 (N_4206,In_1511,In_803);
or U4207 (N_4207,In_2151,In_1195);
or U4208 (N_4208,In_1136,In_1691);
nand U4209 (N_4209,In_334,In_874);
nand U4210 (N_4210,In_18,In_2096);
xor U4211 (N_4211,In_1114,In_937);
and U4212 (N_4212,In_2085,In_553);
or U4213 (N_4213,In_238,In_106);
nand U4214 (N_4214,In_858,In_1388);
xor U4215 (N_4215,In_1953,In_2430);
xor U4216 (N_4216,In_639,In_1648);
or U4217 (N_4217,In_1397,In_1493);
nor U4218 (N_4218,In_710,In_1807);
nand U4219 (N_4219,In_1350,In_1180);
and U4220 (N_4220,In_1375,In_1949);
nor U4221 (N_4221,In_1476,In_2248);
nand U4222 (N_4222,In_1151,In_2438);
nor U4223 (N_4223,In_344,In_702);
nor U4224 (N_4224,In_31,In_1944);
or U4225 (N_4225,In_1561,In_1974);
and U4226 (N_4226,In_613,In_2405);
nand U4227 (N_4227,In_1159,In_936);
xnor U4228 (N_4228,In_1370,In_1475);
nand U4229 (N_4229,In_1009,In_436);
nor U4230 (N_4230,In_160,In_2255);
or U4231 (N_4231,In_851,In_1348);
nor U4232 (N_4232,In_528,In_1757);
or U4233 (N_4233,In_1387,In_1308);
or U4234 (N_4234,In_1188,In_1901);
nand U4235 (N_4235,In_1392,In_1734);
xor U4236 (N_4236,In_530,In_288);
nor U4237 (N_4237,In_573,In_550);
nand U4238 (N_4238,In_2167,In_534);
and U4239 (N_4239,In_2454,In_323);
nor U4240 (N_4240,In_89,In_1992);
and U4241 (N_4241,In_1538,In_1121);
nand U4242 (N_4242,In_1764,In_2198);
and U4243 (N_4243,In_2311,In_1578);
nand U4244 (N_4244,In_1899,In_777);
or U4245 (N_4245,In_2199,In_1155);
nand U4246 (N_4246,In_1795,In_385);
xnor U4247 (N_4247,In_2304,In_1440);
nor U4248 (N_4248,In_1359,In_2296);
nor U4249 (N_4249,In_760,In_1054);
or U4250 (N_4250,In_402,In_89);
nand U4251 (N_4251,In_1615,In_1348);
nand U4252 (N_4252,In_2435,In_1165);
or U4253 (N_4253,In_519,In_2380);
and U4254 (N_4254,In_2391,In_2250);
and U4255 (N_4255,In_814,In_1090);
nand U4256 (N_4256,In_1402,In_1787);
xnor U4257 (N_4257,In_1948,In_212);
or U4258 (N_4258,In_2186,In_1596);
nand U4259 (N_4259,In_247,In_1998);
and U4260 (N_4260,In_1895,In_1698);
nor U4261 (N_4261,In_1647,In_1421);
nor U4262 (N_4262,In_1094,In_1751);
nor U4263 (N_4263,In_1436,In_1170);
nand U4264 (N_4264,In_2075,In_2179);
nand U4265 (N_4265,In_1620,In_495);
or U4266 (N_4266,In_1847,In_395);
nor U4267 (N_4267,In_2427,In_911);
nor U4268 (N_4268,In_722,In_1199);
xor U4269 (N_4269,In_1971,In_1522);
nor U4270 (N_4270,In_871,In_1744);
nor U4271 (N_4271,In_1726,In_1813);
and U4272 (N_4272,In_1929,In_1604);
xor U4273 (N_4273,In_1692,In_485);
nand U4274 (N_4274,In_1543,In_1915);
nand U4275 (N_4275,In_643,In_286);
nor U4276 (N_4276,In_131,In_2164);
xor U4277 (N_4277,In_1206,In_1096);
nor U4278 (N_4278,In_1524,In_1593);
nand U4279 (N_4279,In_1293,In_1769);
nor U4280 (N_4280,In_1516,In_2201);
or U4281 (N_4281,In_1886,In_2261);
nor U4282 (N_4282,In_2361,In_1892);
nor U4283 (N_4283,In_1520,In_572);
or U4284 (N_4284,In_1357,In_1751);
and U4285 (N_4285,In_487,In_494);
xor U4286 (N_4286,In_154,In_2120);
xor U4287 (N_4287,In_1744,In_359);
xor U4288 (N_4288,In_336,In_622);
nor U4289 (N_4289,In_1721,In_1442);
xnor U4290 (N_4290,In_1020,In_368);
or U4291 (N_4291,In_726,In_247);
or U4292 (N_4292,In_21,In_608);
or U4293 (N_4293,In_236,In_1638);
nor U4294 (N_4294,In_773,In_1653);
nor U4295 (N_4295,In_2248,In_216);
nor U4296 (N_4296,In_1518,In_376);
and U4297 (N_4297,In_1048,In_1289);
nor U4298 (N_4298,In_2247,In_1299);
nand U4299 (N_4299,In_272,In_1107);
nor U4300 (N_4300,In_608,In_2458);
nand U4301 (N_4301,In_2157,In_749);
nor U4302 (N_4302,In_170,In_2116);
nor U4303 (N_4303,In_2397,In_1257);
nand U4304 (N_4304,In_902,In_728);
and U4305 (N_4305,In_1718,In_1150);
xnor U4306 (N_4306,In_1986,In_853);
or U4307 (N_4307,In_912,In_565);
or U4308 (N_4308,In_2184,In_1970);
nor U4309 (N_4309,In_2174,In_731);
or U4310 (N_4310,In_344,In_648);
xnor U4311 (N_4311,In_662,In_1875);
nand U4312 (N_4312,In_1576,In_101);
and U4313 (N_4313,In_33,In_1764);
nor U4314 (N_4314,In_1790,In_382);
or U4315 (N_4315,In_701,In_2249);
nor U4316 (N_4316,In_359,In_1003);
nor U4317 (N_4317,In_916,In_1138);
and U4318 (N_4318,In_1183,In_2090);
xor U4319 (N_4319,In_1757,In_1073);
nor U4320 (N_4320,In_790,In_1554);
xnor U4321 (N_4321,In_1717,In_351);
nor U4322 (N_4322,In_348,In_69);
or U4323 (N_4323,In_438,In_1614);
and U4324 (N_4324,In_327,In_1816);
or U4325 (N_4325,In_2160,In_440);
nand U4326 (N_4326,In_1504,In_2227);
or U4327 (N_4327,In_1368,In_975);
nand U4328 (N_4328,In_1334,In_1290);
and U4329 (N_4329,In_370,In_1027);
and U4330 (N_4330,In_399,In_2494);
nor U4331 (N_4331,In_654,In_1360);
nor U4332 (N_4332,In_904,In_57);
nand U4333 (N_4333,In_267,In_2476);
nor U4334 (N_4334,In_1274,In_1671);
xor U4335 (N_4335,In_814,In_2233);
nor U4336 (N_4336,In_2177,In_1228);
or U4337 (N_4337,In_2127,In_323);
xor U4338 (N_4338,In_517,In_1671);
and U4339 (N_4339,In_2498,In_190);
and U4340 (N_4340,In_947,In_1633);
and U4341 (N_4341,In_1259,In_50);
nand U4342 (N_4342,In_2089,In_1382);
nand U4343 (N_4343,In_1599,In_1780);
nand U4344 (N_4344,In_1472,In_1608);
and U4345 (N_4345,In_995,In_1836);
or U4346 (N_4346,In_670,In_2432);
xnor U4347 (N_4347,In_1644,In_1476);
nor U4348 (N_4348,In_478,In_1850);
xnor U4349 (N_4349,In_196,In_1582);
nand U4350 (N_4350,In_1648,In_1445);
xnor U4351 (N_4351,In_1615,In_2107);
nor U4352 (N_4352,In_2315,In_488);
and U4353 (N_4353,In_1813,In_2477);
nor U4354 (N_4354,In_2029,In_2490);
or U4355 (N_4355,In_2486,In_1733);
nand U4356 (N_4356,In_514,In_2146);
nand U4357 (N_4357,In_1505,In_109);
or U4358 (N_4358,In_1193,In_152);
nand U4359 (N_4359,In_1699,In_1155);
xnor U4360 (N_4360,In_1273,In_2243);
nand U4361 (N_4361,In_457,In_201);
nor U4362 (N_4362,In_1554,In_733);
xnor U4363 (N_4363,In_1166,In_1792);
nor U4364 (N_4364,In_50,In_991);
xor U4365 (N_4365,In_883,In_1949);
nor U4366 (N_4366,In_1576,In_301);
xor U4367 (N_4367,In_1507,In_673);
xor U4368 (N_4368,In_2028,In_152);
nor U4369 (N_4369,In_1749,In_245);
nand U4370 (N_4370,In_1108,In_445);
nand U4371 (N_4371,In_766,In_1398);
or U4372 (N_4372,In_1275,In_680);
nor U4373 (N_4373,In_410,In_1196);
and U4374 (N_4374,In_494,In_2164);
xor U4375 (N_4375,In_319,In_2218);
xnor U4376 (N_4376,In_1281,In_470);
nand U4377 (N_4377,In_1328,In_63);
nand U4378 (N_4378,In_1450,In_1293);
or U4379 (N_4379,In_884,In_1558);
and U4380 (N_4380,In_2242,In_408);
and U4381 (N_4381,In_2106,In_602);
and U4382 (N_4382,In_1879,In_813);
xnor U4383 (N_4383,In_65,In_1209);
or U4384 (N_4384,In_1344,In_2483);
nor U4385 (N_4385,In_2040,In_546);
and U4386 (N_4386,In_1025,In_422);
nand U4387 (N_4387,In_1080,In_2098);
nand U4388 (N_4388,In_118,In_1476);
nand U4389 (N_4389,In_1387,In_566);
and U4390 (N_4390,In_2395,In_923);
and U4391 (N_4391,In_643,In_880);
nand U4392 (N_4392,In_928,In_1914);
nor U4393 (N_4393,In_842,In_1550);
or U4394 (N_4394,In_1934,In_1622);
xnor U4395 (N_4395,In_499,In_1863);
or U4396 (N_4396,In_1099,In_1524);
and U4397 (N_4397,In_1717,In_151);
nand U4398 (N_4398,In_2131,In_1594);
and U4399 (N_4399,In_374,In_566);
xor U4400 (N_4400,In_896,In_833);
and U4401 (N_4401,In_1228,In_1649);
and U4402 (N_4402,In_743,In_2170);
xnor U4403 (N_4403,In_2320,In_2258);
and U4404 (N_4404,In_631,In_2287);
xnor U4405 (N_4405,In_1120,In_2478);
xnor U4406 (N_4406,In_2451,In_806);
or U4407 (N_4407,In_1753,In_1523);
nand U4408 (N_4408,In_276,In_1368);
or U4409 (N_4409,In_1272,In_1610);
nor U4410 (N_4410,In_1005,In_2223);
or U4411 (N_4411,In_1418,In_19);
nand U4412 (N_4412,In_1844,In_2340);
nand U4413 (N_4413,In_923,In_671);
nand U4414 (N_4414,In_1542,In_1637);
and U4415 (N_4415,In_579,In_1322);
nand U4416 (N_4416,In_1895,In_2365);
nor U4417 (N_4417,In_546,In_2362);
nand U4418 (N_4418,In_745,In_1453);
and U4419 (N_4419,In_958,In_26);
nor U4420 (N_4420,In_535,In_1627);
and U4421 (N_4421,In_1497,In_2275);
nand U4422 (N_4422,In_988,In_304);
nand U4423 (N_4423,In_929,In_1108);
nor U4424 (N_4424,In_1884,In_322);
xnor U4425 (N_4425,In_1604,In_1008);
nand U4426 (N_4426,In_991,In_1368);
or U4427 (N_4427,In_1190,In_1673);
nor U4428 (N_4428,In_190,In_1451);
nor U4429 (N_4429,In_644,In_2121);
nor U4430 (N_4430,In_405,In_960);
nor U4431 (N_4431,In_1743,In_2237);
nor U4432 (N_4432,In_310,In_1833);
or U4433 (N_4433,In_754,In_722);
and U4434 (N_4434,In_1448,In_2179);
xnor U4435 (N_4435,In_356,In_1392);
and U4436 (N_4436,In_1385,In_1891);
xor U4437 (N_4437,In_2416,In_1532);
xor U4438 (N_4438,In_1610,In_498);
or U4439 (N_4439,In_325,In_1780);
nor U4440 (N_4440,In_357,In_1820);
or U4441 (N_4441,In_231,In_2125);
or U4442 (N_4442,In_1757,In_195);
nor U4443 (N_4443,In_338,In_2371);
nor U4444 (N_4444,In_1094,In_1407);
and U4445 (N_4445,In_2236,In_120);
nand U4446 (N_4446,In_1104,In_706);
xor U4447 (N_4447,In_727,In_1216);
nor U4448 (N_4448,In_1484,In_1078);
xnor U4449 (N_4449,In_1411,In_73);
nor U4450 (N_4450,In_61,In_1087);
or U4451 (N_4451,In_704,In_322);
xor U4452 (N_4452,In_1201,In_501);
or U4453 (N_4453,In_1627,In_2186);
nor U4454 (N_4454,In_1210,In_1490);
or U4455 (N_4455,In_1045,In_384);
or U4456 (N_4456,In_1521,In_1778);
nand U4457 (N_4457,In_2011,In_2035);
nor U4458 (N_4458,In_705,In_1586);
and U4459 (N_4459,In_1572,In_744);
or U4460 (N_4460,In_1255,In_2495);
xor U4461 (N_4461,In_2183,In_648);
xnor U4462 (N_4462,In_1492,In_668);
xor U4463 (N_4463,In_1910,In_2010);
or U4464 (N_4464,In_1020,In_1751);
and U4465 (N_4465,In_1370,In_1453);
nor U4466 (N_4466,In_686,In_593);
nand U4467 (N_4467,In_2462,In_984);
nor U4468 (N_4468,In_1754,In_358);
xnor U4469 (N_4469,In_1492,In_233);
xnor U4470 (N_4470,In_200,In_110);
nand U4471 (N_4471,In_1855,In_1181);
xnor U4472 (N_4472,In_1708,In_1554);
nor U4473 (N_4473,In_1609,In_1938);
nor U4474 (N_4474,In_824,In_2161);
nand U4475 (N_4475,In_192,In_1614);
xor U4476 (N_4476,In_480,In_1954);
or U4477 (N_4477,In_298,In_765);
and U4478 (N_4478,In_1257,In_2328);
or U4479 (N_4479,In_438,In_360);
and U4480 (N_4480,In_940,In_1804);
xor U4481 (N_4481,In_53,In_2073);
xor U4482 (N_4482,In_47,In_1319);
xnor U4483 (N_4483,In_32,In_1787);
nor U4484 (N_4484,In_2418,In_1727);
nand U4485 (N_4485,In_134,In_216);
or U4486 (N_4486,In_2054,In_82);
or U4487 (N_4487,In_1592,In_2034);
xnor U4488 (N_4488,In_2484,In_440);
nor U4489 (N_4489,In_2436,In_326);
and U4490 (N_4490,In_619,In_634);
or U4491 (N_4491,In_322,In_2334);
nor U4492 (N_4492,In_104,In_600);
xnor U4493 (N_4493,In_2082,In_205);
nor U4494 (N_4494,In_2278,In_1294);
and U4495 (N_4495,In_815,In_730);
nor U4496 (N_4496,In_2019,In_155);
xor U4497 (N_4497,In_318,In_1340);
and U4498 (N_4498,In_310,In_1368);
nand U4499 (N_4499,In_1856,In_2416);
nand U4500 (N_4500,In_166,In_1191);
nand U4501 (N_4501,In_2076,In_2342);
and U4502 (N_4502,In_603,In_369);
nand U4503 (N_4503,In_2311,In_1036);
and U4504 (N_4504,In_313,In_795);
or U4505 (N_4505,In_2253,In_1055);
or U4506 (N_4506,In_1267,In_1197);
nor U4507 (N_4507,In_1804,In_1227);
nand U4508 (N_4508,In_2384,In_404);
nand U4509 (N_4509,In_138,In_1024);
xnor U4510 (N_4510,In_780,In_467);
or U4511 (N_4511,In_1831,In_1645);
and U4512 (N_4512,In_929,In_1029);
xor U4513 (N_4513,In_1214,In_1752);
nand U4514 (N_4514,In_242,In_61);
and U4515 (N_4515,In_641,In_1407);
and U4516 (N_4516,In_1465,In_1391);
xor U4517 (N_4517,In_308,In_1205);
or U4518 (N_4518,In_427,In_1914);
and U4519 (N_4519,In_2014,In_622);
nor U4520 (N_4520,In_2054,In_1371);
nor U4521 (N_4521,In_422,In_252);
nand U4522 (N_4522,In_66,In_604);
nand U4523 (N_4523,In_850,In_202);
nor U4524 (N_4524,In_909,In_213);
xor U4525 (N_4525,In_464,In_2224);
or U4526 (N_4526,In_195,In_478);
and U4527 (N_4527,In_268,In_1495);
nand U4528 (N_4528,In_217,In_1822);
or U4529 (N_4529,In_2066,In_975);
or U4530 (N_4530,In_1175,In_132);
nor U4531 (N_4531,In_878,In_1443);
and U4532 (N_4532,In_1203,In_1884);
xor U4533 (N_4533,In_1742,In_1801);
and U4534 (N_4534,In_1601,In_1722);
nand U4535 (N_4535,In_234,In_1039);
nand U4536 (N_4536,In_2281,In_1134);
or U4537 (N_4537,In_2346,In_1776);
nor U4538 (N_4538,In_2185,In_570);
or U4539 (N_4539,In_451,In_1834);
nor U4540 (N_4540,In_552,In_1143);
and U4541 (N_4541,In_560,In_607);
or U4542 (N_4542,In_364,In_1909);
or U4543 (N_4543,In_151,In_2344);
and U4544 (N_4544,In_811,In_1188);
or U4545 (N_4545,In_2060,In_563);
or U4546 (N_4546,In_2413,In_1354);
xor U4547 (N_4547,In_1878,In_1530);
or U4548 (N_4548,In_776,In_586);
nor U4549 (N_4549,In_1311,In_2447);
nand U4550 (N_4550,In_447,In_468);
xor U4551 (N_4551,In_759,In_1945);
nor U4552 (N_4552,In_1076,In_2005);
or U4553 (N_4553,In_908,In_695);
nand U4554 (N_4554,In_556,In_1661);
xor U4555 (N_4555,In_2135,In_676);
and U4556 (N_4556,In_2467,In_2129);
or U4557 (N_4557,In_1204,In_1638);
xor U4558 (N_4558,In_1807,In_2456);
and U4559 (N_4559,In_717,In_7);
nor U4560 (N_4560,In_1503,In_1577);
nand U4561 (N_4561,In_108,In_235);
or U4562 (N_4562,In_1158,In_2217);
nor U4563 (N_4563,In_1633,In_1128);
and U4564 (N_4564,In_281,In_1729);
xor U4565 (N_4565,In_232,In_392);
or U4566 (N_4566,In_1877,In_957);
nor U4567 (N_4567,In_1623,In_1689);
and U4568 (N_4568,In_31,In_811);
and U4569 (N_4569,In_924,In_991);
or U4570 (N_4570,In_551,In_274);
or U4571 (N_4571,In_1942,In_902);
nand U4572 (N_4572,In_344,In_242);
nor U4573 (N_4573,In_1434,In_1393);
or U4574 (N_4574,In_2007,In_131);
or U4575 (N_4575,In_1985,In_2381);
nor U4576 (N_4576,In_259,In_1881);
and U4577 (N_4577,In_1018,In_602);
nand U4578 (N_4578,In_1655,In_2133);
nor U4579 (N_4579,In_2199,In_2283);
or U4580 (N_4580,In_1728,In_438);
nor U4581 (N_4581,In_1369,In_744);
and U4582 (N_4582,In_1425,In_1995);
and U4583 (N_4583,In_79,In_1088);
and U4584 (N_4584,In_979,In_1063);
xnor U4585 (N_4585,In_2295,In_1088);
or U4586 (N_4586,In_1734,In_1751);
xnor U4587 (N_4587,In_452,In_757);
and U4588 (N_4588,In_2371,In_1069);
nor U4589 (N_4589,In_2341,In_869);
nand U4590 (N_4590,In_1424,In_439);
xnor U4591 (N_4591,In_1967,In_2496);
nor U4592 (N_4592,In_1007,In_362);
or U4593 (N_4593,In_2335,In_2165);
nor U4594 (N_4594,In_1654,In_1783);
nor U4595 (N_4595,In_2476,In_1530);
xor U4596 (N_4596,In_369,In_379);
and U4597 (N_4597,In_27,In_488);
and U4598 (N_4598,In_148,In_1689);
xnor U4599 (N_4599,In_294,In_2458);
and U4600 (N_4600,In_2490,In_1490);
nor U4601 (N_4601,In_1381,In_1100);
and U4602 (N_4602,In_1604,In_2264);
nor U4603 (N_4603,In_1076,In_2318);
nor U4604 (N_4604,In_2157,In_1820);
and U4605 (N_4605,In_1784,In_1248);
nor U4606 (N_4606,In_214,In_474);
and U4607 (N_4607,In_285,In_745);
xnor U4608 (N_4608,In_64,In_616);
nand U4609 (N_4609,In_1973,In_1636);
and U4610 (N_4610,In_1397,In_494);
nor U4611 (N_4611,In_2430,In_639);
xnor U4612 (N_4612,In_797,In_1025);
xor U4613 (N_4613,In_632,In_2053);
nand U4614 (N_4614,In_625,In_235);
nor U4615 (N_4615,In_7,In_2134);
and U4616 (N_4616,In_1885,In_2304);
xor U4617 (N_4617,In_1797,In_2020);
nand U4618 (N_4618,In_174,In_210);
xnor U4619 (N_4619,In_2439,In_201);
nand U4620 (N_4620,In_1018,In_1579);
xnor U4621 (N_4621,In_315,In_446);
and U4622 (N_4622,In_1320,In_152);
xnor U4623 (N_4623,In_1267,In_2207);
or U4624 (N_4624,In_2380,In_576);
xor U4625 (N_4625,In_127,In_1582);
nor U4626 (N_4626,In_1608,In_252);
xor U4627 (N_4627,In_2316,In_2270);
or U4628 (N_4628,In_1232,In_974);
nand U4629 (N_4629,In_1431,In_1250);
nor U4630 (N_4630,In_1295,In_2412);
or U4631 (N_4631,In_1928,In_2408);
xnor U4632 (N_4632,In_231,In_816);
and U4633 (N_4633,In_2331,In_762);
nand U4634 (N_4634,In_29,In_1875);
nand U4635 (N_4635,In_1734,In_1995);
nand U4636 (N_4636,In_1706,In_222);
nor U4637 (N_4637,In_1433,In_1652);
and U4638 (N_4638,In_415,In_290);
xnor U4639 (N_4639,In_2192,In_639);
nand U4640 (N_4640,In_1134,In_771);
or U4641 (N_4641,In_809,In_698);
nand U4642 (N_4642,In_680,In_831);
and U4643 (N_4643,In_843,In_458);
xor U4644 (N_4644,In_2139,In_2158);
nor U4645 (N_4645,In_2201,In_1191);
xnor U4646 (N_4646,In_1350,In_1887);
nor U4647 (N_4647,In_2259,In_682);
and U4648 (N_4648,In_1749,In_2398);
or U4649 (N_4649,In_84,In_616);
nand U4650 (N_4650,In_1251,In_571);
or U4651 (N_4651,In_1536,In_257);
or U4652 (N_4652,In_1134,In_1548);
nand U4653 (N_4653,In_1590,In_1357);
nor U4654 (N_4654,In_403,In_2226);
or U4655 (N_4655,In_622,In_2145);
nor U4656 (N_4656,In_175,In_865);
or U4657 (N_4657,In_1540,In_1651);
and U4658 (N_4658,In_1149,In_445);
nand U4659 (N_4659,In_2461,In_2426);
and U4660 (N_4660,In_1341,In_284);
or U4661 (N_4661,In_724,In_247);
nor U4662 (N_4662,In_2406,In_406);
xor U4663 (N_4663,In_1992,In_1274);
xor U4664 (N_4664,In_1733,In_2020);
nand U4665 (N_4665,In_274,In_1795);
nor U4666 (N_4666,In_1387,In_1436);
nand U4667 (N_4667,In_1179,In_2119);
or U4668 (N_4668,In_572,In_2046);
or U4669 (N_4669,In_1760,In_2227);
nand U4670 (N_4670,In_1329,In_2329);
or U4671 (N_4671,In_982,In_2087);
nor U4672 (N_4672,In_1086,In_192);
or U4673 (N_4673,In_879,In_1526);
or U4674 (N_4674,In_475,In_750);
and U4675 (N_4675,In_320,In_1797);
xor U4676 (N_4676,In_603,In_2274);
and U4677 (N_4677,In_1195,In_2130);
nor U4678 (N_4678,In_1523,In_2182);
nor U4679 (N_4679,In_853,In_557);
or U4680 (N_4680,In_2178,In_330);
nand U4681 (N_4681,In_304,In_1345);
and U4682 (N_4682,In_1384,In_2310);
nor U4683 (N_4683,In_1850,In_2062);
xnor U4684 (N_4684,In_1728,In_2488);
and U4685 (N_4685,In_1057,In_1576);
and U4686 (N_4686,In_101,In_443);
nor U4687 (N_4687,In_1846,In_1164);
or U4688 (N_4688,In_785,In_316);
nor U4689 (N_4689,In_1949,In_653);
and U4690 (N_4690,In_1379,In_42);
or U4691 (N_4691,In_2451,In_1079);
xnor U4692 (N_4692,In_1378,In_1352);
and U4693 (N_4693,In_2421,In_2147);
nor U4694 (N_4694,In_1534,In_632);
or U4695 (N_4695,In_1262,In_2113);
nor U4696 (N_4696,In_928,In_826);
xor U4697 (N_4697,In_637,In_123);
or U4698 (N_4698,In_2131,In_2210);
nand U4699 (N_4699,In_756,In_515);
nor U4700 (N_4700,In_456,In_2409);
and U4701 (N_4701,In_2424,In_1284);
nand U4702 (N_4702,In_38,In_633);
and U4703 (N_4703,In_2017,In_1597);
nor U4704 (N_4704,In_18,In_84);
nand U4705 (N_4705,In_562,In_1007);
xnor U4706 (N_4706,In_954,In_1968);
or U4707 (N_4707,In_1861,In_2312);
xor U4708 (N_4708,In_1049,In_1990);
and U4709 (N_4709,In_306,In_1715);
nand U4710 (N_4710,In_2257,In_2186);
nor U4711 (N_4711,In_2395,In_1467);
or U4712 (N_4712,In_1982,In_442);
or U4713 (N_4713,In_1899,In_2261);
nand U4714 (N_4714,In_992,In_1776);
and U4715 (N_4715,In_1012,In_1086);
nor U4716 (N_4716,In_248,In_1619);
and U4717 (N_4717,In_2275,In_89);
xnor U4718 (N_4718,In_2269,In_1324);
nand U4719 (N_4719,In_2172,In_691);
and U4720 (N_4720,In_97,In_1933);
or U4721 (N_4721,In_1999,In_115);
nor U4722 (N_4722,In_2145,In_766);
nor U4723 (N_4723,In_1581,In_1035);
xnor U4724 (N_4724,In_829,In_2437);
or U4725 (N_4725,In_1150,In_2065);
or U4726 (N_4726,In_1441,In_1391);
or U4727 (N_4727,In_724,In_368);
xor U4728 (N_4728,In_683,In_836);
or U4729 (N_4729,In_1991,In_1840);
and U4730 (N_4730,In_357,In_235);
nand U4731 (N_4731,In_1110,In_1254);
and U4732 (N_4732,In_1515,In_882);
or U4733 (N_4733,In_1775,In_1502);
xnor U4734 (N_4734,In_1966,In_1181);
nor U4735 (N_4735,In_422,In_2235);
nand U4736 (N_4736,In_1351,In_634);
nand U4737 (N_4737,In_1815,In_1968);
or U4738 (N_4738,In_378,In_347);
xnor U4739 (N_4739,In_1629,In_1846);
nand U4740 (N_4740,In_1693,In_656);
nand U4741 (N_4741,In_299,In_2253);
or U4742 (N_4742,In_471,In_953);
xor U4743 (N_4743,In_496,In_386);
or U4744 (N_4744,In_1763,In_966);
and U4745 (N_4745,In_1431,In_14);
xnor U4746 (N_4746,In_1909,In_2411);
and U4747 (N_4747,In_2470,In_446);
or U4748 (N_4748,In_486,In_553);
or U4749 (N_4749,In_1562,In_213);
or U4750 (N_4750,In_241,In_901);
xor U4751 (N_4751,In_1637,In_597);
xnor U4752 (N_4752,In_1170,In_2018);
or U4753 (N_4753,In_948,In_1406);
nand U4754 (N_4754,In_2496,In_124);
or U4755 (N_4755,In_1294,In_530);
nor U4756 (N_4756,In_819,In_212);
and U4757 (N_4757,In_2485,In_642);
nand U4758 (N_4758,In_1077,In_996);
or U4759 (N_4759,In_1702,In_735);
xnor U4760 (N_4760,In_473,In_178);
or U4761 (N_4761,In_1863,In_167);
or U4762 (N_4762,In_681,In_2487);
or U4763 (N_4763,In_2411,In_933);
nand U4764 (N_4764,In_1869,In_992);
and U4765 (N_4765,In_481,In_434);
and U4766 (N_4766,In_2106,In_491);
nor U4767 (N_4767,In_1194,In_970);
xor U4768 (N_4768,In_1185,In_1415);
and U4769 (N_4769,In_334,In_442);
nor U4770 (N_4770,In_688,In_1898);
or U4771 (N_4771,In_94,In_740);
nor U4772 (N_4772,In_795,In_347);
xnor U4773 (N_4773,In_1534,In_731);
and U4774 (N_4774,In_1489,In_2496);
nor U4775 (N_4775,In_2087,In_2348);
and U4776 (N_4776,In_1338,In_2431);
nor U4777 (N_4777,In_1222,In_1629);
and U4778 (N_4778,In_2321,In_1129);
nand U4779 (N_4779,In_2009,In_1510);
nor U4780 (N_4780,In_1127,In_1757);
xnor U4781 (N_4781,In_1733,In_2229);
nand U4782 (N_4782,In_1963,In_1136);
or U4783 (N_4783,In_1274,In_349);
nor U4784 (N_4784,In_1737,In_197);
nand U4785 (N_4785,In_982,In_507);
xor U4786 (N_4786,In_151,In_2294);
nor U4787 (N_4787,In_751,In_2181);
xor U4788 (N_4788,In_1596,In_1762);
xor U4789 (N_4789,In_2395,In_652);
and U4790 (N_4790,In_2376,In_1045);
and U4791 (N_4791,In_758,In_612);
or U4792 (N_4792,In_1656,In_1818);
and U4793 (N_4793,In_128,In_214);
or U4794 (N_4794,In_1746,In_1662);
nor U4795 (N_4795,In_1033,In_2451);
nor U4796 (N_4796,In_1542,In_586);
nand U4797 (N_4797,In_322,In_202);
nand U4798 (N_4798,In_1710,In_794);
nand U4799 (N_4799,In_1273,In_267);
nor U4800 (N_4800,In_1209,In_1895);
nor U4801 (N_4801,In_1687,In_2427);
nor U4802 (N_4802,In_1992,In_1437);
and U4803 (N_4803,In_963,In_972);
xnor U4804 (N_4804,In_1623,In_2189);
nand U4805 (N_4805,In_2477,In_692);
xnor U4806 (N_4806,In_845,In_1589);
xnor U4807 (N_4807,In_525,In_609);
xnor U4808 (N_4808,In_1726,In_2491);
xnor U4809 (N_4809,In_1931,In_1785);
xor U4810 (N_4810,In_177,In_46);
and U4811 (N_4811,In_1039,In_2019);
xnor U4812 (N_4812,In_2084,In_1336);
nor U4813 (N_4813,In_1383,In_2253);
xor U4814 (N_4814,In_1476,In_1069);
xnor U4815 (N_4815,In_550,In_1201);
nor U4816 (N_4816,In_1045,In_91);
nor U4817 (N_4817,In_119,In_827);
or U4818 (N_4818,In_2287,In_443);
nand U4819 (N_4819,In_1810,In_182);
xnor U4820 (N_4820,In_444,In_1176);
nand U4821 (N_4821,In_982,In_855);
nand U4822 (N_4822,In_2198,In_901);
or U4823 (N_4823,In_1542,In_1415);
or U4824 (N_4824,In_1406,In_61);
nand U4825 (N_4825,In_1407,In_1322);
and U4826 (N_4826,In_1511,In_1769);
nor U4827 (N_4827,In_1564,In_908);
xnor U4828 (N_4828,In_1800,In_1297);
and U4829 (N_4829,In_1402,In_190);
nor U4830 (N_4830,In_1745,In_125);
or U4831 (N_4831,In_665,In_1654);
and U4832 (N_4832,In_1066,In_1067);
nand U4833 (N_4833,In_1314,In_38);
nor U4834 (N_4834,In_2311,In_2434);
xnor U4835 (N_4835,In_227,In_142);
xnor U4836 (N_4836,In_88,In_11);
xor U4837 (N_4837,In_1020,In_1656);
nand U4838 (N_4838,In_428,In_289);
or U4839 (N_4839,In_1925,In_1176);
nor U4840 (N_4840,In_1319,In_2042);
and U4841 (N_4841,In_2175,In_1965);
nand U4842 (N_4842,In_13,In_752);
nor U4843 (N_4843,In_133,In_1185);
nand U4844 (N_4844,In_1960,In_1013);
nor U4845 (N_4845,In_1399,In_1000);
and U4846 (N_4846,In_1358,In_1094);
nand U4847 (N_4847,In_1937,In_1262);
nand U4848 (N_4848,In_1026,In_342);
or U4849 (N_4849,In_1429,In_1978);
nand U4850 (N_4850,In_2278,In_306);
nand U4851 (N_4851,In_2101,In_687);
nor U4852 (N_4852,In_1637,In_712);
nor U4853 (N_4853,In_1410,In_691);
or U4854 (N_4854,In_619,In_2116);
nor U4855 (N_4855,In_509,In_308);
nor U4856 (N_4856,In_992,In_493);
nand U4857 (N_4857,In_1864,In_1234);
or U4858 (N_4858,In_649,In_1427);
xnor U4859 (N_4859,In_1613,In_2296);
and U4860 (N_4860,In_850,In_1439);
nor U4861 (N_4861,In_740,In_1672);
nor U4862 (N_4862,In_233,In_792);
nor U4863 (N_4863,In_1518,In_554);
nand U4864 (N_4864,In_1416,In_2441);
xor U4865 (N_4865,In_2290,In_775);
and U4866 (N_4866,In_2112,In_981);
or U4867 (N_4867,In_2077,In_1098);
nand U4868 (N_4868,In_2195,In_1246);
nor U4869 (N_4869,In_185,In_1771);
nand U4870 (N_4870,In_1780,In_10);
and U4871 (N_4871,In_782,In_1511);
xor U4872 (N_4872,In_1020,In_1766);
and U4873 (N_4873,In_865,In_869);
and U4874 (N_4874,In_1865,In_2146);
or U4875 (N_4875,In_1297,In_641);
nand U4876 (N_4876,In_709,In_2071);
and U4877 (N_4877,In_318,In_2109);
or U4878 (N_4878,In_2104,In_1714);
or U4879 (N_4879,In_862,In_891);
xnor U4880 (N_4880,In_867,In_312);
or U4881 (N_4881,In_657,In_983);
xnor U4882 (N_4882,In_539,In_876);
or U4883 (N_4883,In_1927,In_2387);
nor U4884 (N_4884,In_2366,In_1049);
and U4885 (N_4885,In_1307,In_1242);
nand U4886 (N_4886,In_1268,In_234);
nand U4887 (N_4887,In_2119,In_2169);
or U4888 (N_4888,In_58,In_775);
or U4889 (N_4889,In_2345,In_1700);
nor U4890 (N_4890,In_1202,In_2334);
nand U4891 (N_4891,In_2163,In_296);
nand U4892 (N_4892,In_2385,In_1122);
or U4893 (N_4893,In_2499,In_955);
and U4894 (N_4894,In_2309,In_1803);
or U4895 (N_4895,In_1442,In_1332);
or U4896 (N_4896,In_965,In_2006);
and U4897 (N_4897,In_599,In_906);
nor U4898 (N_4898,In_1957,In_1256);
nor U4899 (N_4899,In_322,In_1472);
or U4900 (N_4900,In_1337,In_1202);
and U4901 (N_4901,In_912,In_713);
nand U4902 (N_4902,In_800,In_1170);
nor U4903 (N_4903,In_2268,In_1552);
and U4904 (N_4904,In_93,In_2343);
or U4905 (N_4905,In_2465,In_1186);
or U4906 (N_4906,In_1851,In_2363);
nand U4907 (N_4907,In_567,In_2032);
or U4908 (N_4908,In_1766,In_2436);
and U4909 (N_4909,In_2295,In_1935);
nor U4910 (N_4910,In_636,In_55);
or U4911 (N_4911,In_1911,In_2033);
xnor U4912 (N_4912,In_2373,In_1563);
or U4913 (N_4913,In_619,In_2493);
nand U4914 (N_4914,In_2405,In_2407);
xor U4915 (N_4915,In_2242,In_533);
or U4916 (N_4916,In_2438,In_1233);
nor U4917 (N_4917,In_1416,In_1678);
xor U4918 (N_4918,In_341,In_1569);
nor U4919 (N_4919,In_461,In_1945);
and U4920 (N_4920,In_894,In_580);
nand U4921 (N_4921,In_182,In_667);
or U4922 (N_4922,In_2480,In_2204);
and U4923 (N_4923,In_1720,In_2441);
and U4924 (N_4924,In_614,In_1927);
nand U4925 (N_4925,In_1049,In_2466);
nor U4926 (N_4926,In_1742,In_984);
and U4927 (N_4927,In_1837,In_1660);
and U4928 (N_4928,In_1200,In_1131);
or U4929 (N_4929,In_1662,In_62);
nand U4930 (N_4930,In_485,In_321);
or U4931 (N_4931,In_2393,In_2281);
or U4932 (N_4932,In_2068,In_1842);
nand U4933 (N_4933,In_123,In_657);
nand U4934 (N_4934,In_400,In_1257);
xor U4935 (N_4935,In_1206,In_1249);
and U4936 (N_4936,In_1419,In_2466);
or U4937 (N_4937,In_1752,In_1755);
xor U4938 (N_4938,In_1937,In_1815);
nand U4939 (N_4939,In_987,In_847);
nor U4940 (N_4940,In_1745,In_636);
or U4941 (N_4941,In_1321,In_1586);
and U4942 (N_4942,In_1804,In_886);
xor U4943 (N_4943,In_680,In_1894);
and U4944 (N_4944,In_273,In_2474);
nor U4945 (N_4945,In_1724,In_1113);
and U4946 (N_4946,In_1537,In_1217);
or U4947 (N_4947,In_760,In_2414);
xnor U4948 (N_4948,In_592,In_1772);
nor U4949 (N_4949,In_316,In_840);
nor U4950 (N_4950,In_1267,In_69);
or U4951 (N_4951,In_2137,In_1951);
nand U4952 (N_4952,In_1958,In_1733);
or U4953 (N_4953,In_2291,In_1842);
nor U4954 (N_4954,In_2393,In_1683);
xnor U4955 (N_4955,In_375,In_123);
nor U4956 (N_4956,In_1786,In_444);
nor U4957 (N_4957,In_949,In_2065);
nand U4958 (N_4958,In_2013,In_558);
or U4959 (N_4959,In_275,In_2483);
nand U4960 (N_4960,In_131,In_830);
nor U4961 (N_4961,In_1620,In_705);
or U4962 (N_4962,In_2385,In_2339);
or U4963 (N_4963,In_2158,In_2203);
and U4964 (N_4964,In_126,In_2119);
xnor U4965 (N_4965,In_1531,In_971);
nor U4966 (N_4966,In_1568,In_1229);
nand U4967 (N_4967,In_358,In_619);
nand U4968 (N_4968,In_648,In_170);
or U4969 (N_4969,In_1714,In_1982);
xor U4970 (N_4970,In_870,In_2444);
or U4971 (N_4971,In_289,In_1631);
nand U4972 (N_4972,In_2268,In_2035);
and U4973 (N_4973,In_374,In_1453);
or U4974 (N_4974,In_1197,In_1653);
or U4975 (N_4975,In_219,In_177);
nor U4976 (N_4976,In_2120,In_816);
nand U4977 (N_4977,In_351,In_1944);
nor U4978 (N_4978,In_1390,In_624);
or U4979 (N_4979,In_1453,In_61);
xnor U4980 (N_4980,In_1633,In_711);
or U4981 (N_4981,In_1670,In_7);
nand U4982 (N_4982,In_156,In_1135);
nor U4983 (N_4983,In_587,In_2048);
xor U4984 (N_4984,In_1559,In_1668);
nand U4985 (N_4985,In_2093,In_367);
or U4986 (N_4986,In_1850,In_1945);
nor U4987 (N_4987,In_1979,In_1919);
or U4988 (N_4988,In_2111,In_1212);
nor U4989 (N_4989,In_603,In_712);
nor U4990 (N_4990,In_142,In_2266);
nor U4991 (N_4991,In_2099,In_1061);
nand U4992 (N_4992,In_1980,In_1913);
or U4993 (N_4993,In_479,In_2022);
nand U4994 (N_4994,In_1990,In_2230);
nand U4995 (N_4995,In_339,In_2149);
or U4996 (N_4996,In_236,In_963);
and U4997 (N_4997,In_552,In_2252);
and U4998 (N_4998,In_315,In_103);
xnor U4999 (N_4999,In_2452,In_1695);
nor U5000 (N_5000,In_1958,In_2410);
xnor U5001 (N_5001,In_1939,In_2439);
and U5002 (N_5002,In_1191,In_2143);
nor U5003 (N_5003,In_2174,In_1086);
and U5004 (N_5004,In_1263,In_1367);
xor U5005 (N_5005,In_291,In_1942);
nor U5006 (N_5006,In_796,In_1554);
nand U5007 (N_5007,In_295,In_697);
xor U5008 (N_5008,In_1998,In_505);
and U5009 (N_5009,In_2121,In_1983);
xor U5010 (N_5010,In_727,In_1229);
nand U5011 (N_5011,In_1010,In_12);
or U5012 (N_5012,In_647,In_574);
nand U5013 (N_5013,In_1060,In_995);
nor U5014 (N_5014,In_1206,In_1510);
nor U5015 (N_5015,In_2249,In_426);
nor U5016 (N_5016,In_1955,In_969);
nor U5017 (N_5017,In_410,In_1448);
xor U5018 (N_5018,In_1353,In_1271);
nand U5019 (N_5019,In_2159,In_1603);
and U5020 (N_5020,In_388,In_2083);
and U5021 (N_5021,In_2075,In_15);
nand U5022 (N_5022,In_1470,In_644);
or U5023 (N_5023,In_982,In_2320);
or U5024 (N_5024,In_773,In_77);
nor U5025 (N_5025,In_2097,In_292);
nand U5026 (N_5026,In_536,In_1067);
and U5027 (N_5027,In_118,In_1417);
xor U5028 (N_5028,In_394,In_1600);
nand U5029 (N_5029,In_1948,In_2153);
and U5030 (N_5030,In_221,In_1162);
and U5031 (N_5031,In_122,In_1626);
xor U5032 (N_5032,In_88,In_1524);
nor U5033 (N_5033,In_2162,In_2115);
nor U5034 (N_5034,In_1486,In_391);
and U5035 (N_5035,In_1601,In_1603);
and U5036 (N_5036,In_551,In_2387);
and U5037 (N_5037,In_1050,In_2258);
xor U5038 (N_5038,In_606,In_2172);
or U5039 (N_5039,In_542,In_497);
or U5040 (N_5040,In_479,In_1936);
xor U5041 (N_5041,In_578,In_1093);
nand U5042 (N_5042,In_880,In_1396);
and U5043 (N_5043,In_848,In_615);
nor U5044 (N_5044,In_1038,In_996);
xor U5045 (N_5045,In_1774,In_62);
nand U5046 (N_5046,In_1058,In_1688);
xor U5047 (N_5047,In_675,In_1676);
or U5048 (N_5048,In_1298,In_886);
nand U5049 (N_5049,In_2165,In_259);
nor U5050 (N_5050,In_952,In_401);
and U5051 (N_5051,In_2,In_2443);
and U5052 (N_5052,In_1171,In_1213);
nand U5053 (N_5053,In_1912,In_2218);
nand U5054 (N_5054,In_407,In_351);
nor U5055 (N_5055,In_121,In_1037);
nor U5056 (N_5056,In_705,In_1660);
nand U5057 (N_5057,In_1833,In_1911);
nor U5058 (N_5058,In_918,In_1094);
xnor U5059 (N_5059,In_1035,In_1209);
xnor U5060 (N_5060,In_133,In_2299);
or U5061 (N_5061,In_1709,In_839);
and U5062 (N_5062,In_105,In_2179);
xor U5063 (N_5063,In_1685,In_1803);
or U5064 (N_5064,In_1231,In_307);
nand U5065 (N_5065,In_216,In_1195);
nand U5066 (N_5066,In_1537,In_1580);
xor U5067 (N_5067,In_1234,In_2457);
nor U5068 (N_5068,In_1908,In_1611);
and U5069 (N_5069,In_2306,In_127);
or U5070 (N_5070,In_2200,In_737);
and U5071 (N_5071,In_1611,In_610);
and U5072 (N_5072,In_147,In_1548);
nand U5073 (N_5073,In_2289,In_1583);
nor U5074 (N_5074,In_1245,In_2446);
nor U5075 (N_5075,In_457,In_2327);
or U5076 (N_5076,In_1000,In_2307);
or U5077 (N_5077,In_1616,In_739);
nand U5078 (N_5078,In_1732,In_32);
nand U5079 (N_5079,In_488,In_491);
nor U5080 (N_5080,In_796,In_512);
xnor U5081 (N_5081,In_484,In_122);
nor U5082 (N_5082,In_982,In_1382);
xor U5083 (N_5083,In_1913,In_1805);
nand U5084 (N_5084,In_2399,In_2047);
or U5085 (N_5085,In_2059,In_2354);
nand U5086 (N_5086,In_1845,In_2194);
and U5087 (N_5087,In_820,In_1576);
nand U5088 (N_5088,In_367,In_1546);
and U5089 (N_5089,In_907,In_375);
xor U5090 (N_5090,In_2337,In_1580);
nand U5091 (N_5091,In_580,In_816);
or U5092 (N_5092,In_1978,In_542);
or U5093 (N_5093,In_555,In_697);
nand U5094 (N_5094,In_1732,In_1853);
nor U5095 (N_5095,In_1887,In_860);
and U5096 (N_5096,In_2134,In_2421);
xor U5097 (N_5097,In_1892,In_2486);
nor U5098 (N_5098,In_2158,In_257);
nand U5099 (N_5099,In_229,In_848);
or U5100 (N_5100,In_1448,In_1967);
xor U5101 (N_5101,In_742,In_1415);
nand U5102 (N_5102,In_516,In_1406);
or U5103 (N_5103,In_880,In_252);
nor U5104 (N_5104,In_1482,In_2079);
nor U5105 (N_5105,In_2461,In_1195);
xnor U5106 (N_5106,In_577,In_1678);
and U5107 (N_5107,In_2312,In_893);
xnor U5108 (N_5108,In_1870,In_933);
or U5109 (N_5109,In_2015,In_1483);
nor U5110 (N_5110,In_374,In_263);
nor U5111 (N_5111,In_161,In_145);
nor U5112 (N_5112,In_1303,In_2437);
nand U5113 (N_5113,In_1264,In_1344);
or U5114 (N_5114,In_2113,In_137);
nor U5115 (N_5115,In_1102,In_1992);
xor U5116 (N_5116,In_1479,In_1200);
xor U5117 (N_5117,In_401,In_2165);
xor U5118 (N_5118,In_52,In_1407);
or U5119 (N_5119,In_501,In_185);
nor U5120 (N_5120,In_1864,In_900);
or U5121 (N_5121,In_1419,In_983);
xor U5122 (N_5122,In_1406,In_1141);
and U5123 (N_5123,In_1383,In_28);
or U5124 (N_5124,In_55,In_1230);
nor U5125 (N_5125,In_1590,In_1724);
xor U5126 (N_5126,In_1804,In_162);
xnor U5127 (N_5127,In_605,In_1055);
nand U5128 (N_5128,In_1909,In_626);
nor U5129 (N_5129,In_957,In_2274);
or U5130 (N_5130,In_13,In_11);
nand U5131 (N_5131,In_1646,In_1227);
or U5132 (N_5132,In_490,In_1707);
nor U5133 (N_5133,In_326,In_65);
xor U5134 (N_5134,In_2005,In_2057);
or U5135 (N_5135,In_1208,In_702);
and U5136 (N_5136,In_692,In_825);
and U5137 (N_5137,In_2464,In_2142);
and U5138 (N_5138,In_1229,In_757);
and U5139 (N_5139,In_2013,In_723);
nand U5140 (N_5140,In_1052,In_139);
xnor U5141 (N_5141,In_1078,In_1327);
xnor U5142 (N_5142,In_2129,In_1483);
and U5143 (N_5143,In_2128,In_555);
nand U5144 (N_5144,In_2063,In_1685);
and U5145 (N_5145,In_1766,In_1045);
xnor U5146 (N_5146,In_449,In_105);
nand U5147 (N_5147,In_1492,In_487);
xor U5148 (N_5148,In_176,In_1526);
or U5149 (N_5149,In_929,In_1563);
or U5150 (N_5150,In_1637,In_1974);
xor U5151 (N_5151,In_2129,In_1839);
nor U5152 (N_5152,In_1372,In_1947);
nand U5153 (N_5153,In_1851,In_106);
nand U5154 (N_5154,In_1172,In_1466);
or U5155 (N_5155,In_1239,In_1175);
nor U5156 (N_5156,In_2433,In_1147);
nand U5157 (N_5157,In_2498,In_1336);
or U5158 (N_5158,In_599,In_1510);
nor U5159 (N_5159,In_1610,In_740);
nor U5160 (N_5160,In_1063,In_726);
nor U5161 (N_5161,In_224,In_381);
xor U5162 (N_5162,In_1478,In_1889);
xor U5163 (N_5163,In_748,In_638);
xnor U5164 (N_5164,In_717,In_2293);
nand U5165 (N_5165,In_1763,In_1279);
nor U5166 (N_5166,In_1781,In_1438);
xnor U5167 (N_5167,In_556,In_2179);
nor U5168 (N_5168,In_1384,In_182);
and U5169 (N_5169,In_1442,In_805);
or U5170 (N_5170,In_984,In_1515);
and U5171 (N_5171,In_2277,In_279);
xor U5172 (N_5172,In_2077,In_326);
xor U5173 (N_5173,In_1986,In_968);
and U5174 (N_5174,In_535,In_1411);
xor U5175 (N_5175,In_1349,In_2010);
nand U5176 (N_5176,In_957,In_1955);
nor U5177 (N_5177,In_514,In_1658);
nand U5178 (N_5178,In_198,In_2425);
or U5179 (N_5179,In_639,In_1509);
or U5180 (N_5180,In_34,In_820);
or U5181 (N_5181,In_1283,In_497);
and U5182 (N_5182,In_1561,In_2337);
nor U5183 (N_5183,In_191,In_1402);
nand U5184 (N_5184,In_1178,In_1710);
and U5185 (N_5185,In_2350,In_1511);
nand U5186 (N_5186,In_414,In_1784);
and U5187 (N_5187,In_2346,In_540);
or U5188 (N_5188,In_247,In_883);
nor U5189 (N_5189,In_631,In_1545);
and U5190 (N_5190,In_2145,In_1721);
nand U5191 (N_5191,In_2473,In_1781);
nor U5192 (N_5192,In_1415,In_905);
and U5193 (N_5193,In_1996,In_1051);
or U5194 (N_5194,In_1278,In_1608);
or U5195 (N_5195,In_2114,In_1506);
or U5196 (N_5196,In_790,In_1581);
or U5197 (N_5197,In_2082,In_2067);
nand U5198 (N_5198,In_862,In_1050);
or U5199 (N_5199,In_1452,In_2367);
nor U5200 (N_5200,In_739,In_20);
nand U5201 (N_5201,In_1767,In_839);
or U5202 (N_5202,In_383,In_408);
or U5203 (N_5203,In_2223,In_628);
and U5204 (N_5204,In_528,In_1560);
nand U5205 (N_5205,In_1480,In_849);
nor U5206 (N_5206,In_1085,In_431);
nor U5207 (N_5207,In_1656,In_568);
nor U5208 (N_5208,In_130,In_507);
xor U5209 (N_5209,In_2302,In_429);
xnor U5210 (N_5210,In_1304,In_2008);
xnor U5211 (N_5211,In_1658,In_628);
and U5212 (N_5212,In_2285,In_2275);
nor U5213 (N_5213,In_2330,In_1105);
or U5214 (N_5214,In_2310,In_1704);
nor U5215 (N_5215,In_492,In_1309);
nor U5216 (N_5216,In_50,In_1949);
or U5217 (N_5217,In_286,In_1821);
nand U5218 (N_5218,In_329,In_2126);
nor U5219 (N_5219,In_2339,In_168);
and U5220 (N_5220,In_1751,In_2056);
nand U5221 (N_5221,In_1573,In_1544);
nor U5222 (N_5222,In_183,In_1999);
xnor U5223 (N_5223,In_814,In_2289);
xor U5224 (N_5224,In_1819,In_281);
nor U5225 (N_5225,In_18,In_1671);
nor U5226 (N_5226,In_919,In_2166);
nand U5227 (N_5227,In_79,In_408);
or U5228 (N_5228,In_608,In_244);
and U5229 (N_5229,In_1679,In_1793);
xor U5230 (N_5230,In_1445,In_1572);
xor U5231 (N_5231,In_1351,In_1289);
xnor U5232 (N_5232,In_886,In_390);
nand U5233 (N_5233,In_1242,In_540);
or U5234 (N_5234,In_775,In_638);
nand U5235 (N_5235,In_1726,In_337);
xor U5236 (N_5236,In_2024,In_1976);
nand U5237 (N_5237,In_508,In_756);
and U5238 (N_5238,In_594,In_1600);
nor U5239 (N_5239,In_1558,In_2471);
and U5240 (N_5240,In_210,In_513);
nand U5241 (N_5241,In_1442,In_546);
xnor U5242 (N_5242,In_1270,In_661);
xor U5243 (N_5243,In_1449,In_769);
nand U5244 (N_5244,In_500,In_1259);
and U5245 (N_5245,In_194,In_346);
nand U5246 (N_5246,In_2472,In_1554);
nor U5247 (N_5247,In_216,In_1242);
and U5248 (N_5248,In_2018,In_1981);
nor U5249 (N_5249,In_2358,In_1949);
nor U5250 (N_5250,In_404,In_1145);
or U5251 (N_5251,In_1988,In_1163);
xor U5252 (N_5252,In_1166,In_1893);
xnor U5253 (N_5253,In_426,In_1735);
nor U5254 (N_5254,In_2428,In_1039);
nor U5255 (N_5255,In_1318,In_409);
nor U5256 (N_5256,In_558,In_1088);
nor U5257 (N_5257,In_1204,In_1572);
nand U5258 (N_5258,In_917,In_2334);
or U5259 (N_5259,In_897,In_527);
or U5260 (N_5260,In_1765,In_1197);
nor U5261 (N_5261,In_1727,In_2012);
or U5262 (N_5262,In_113,In_1032);
and U5263 (N_5263,In_349,In_1062);
or U5264 (N_5264,In_1508,In_1826);
nand U5265 (N_5265,In_2141,In_1344);
nand U5266 (N_5266,In_1731,In_1320);
xor U5267 (N_5267,In_195,In_1733);
and U5268 (N_5268,In_616,In_154);
nor U5269 (N_5269,In_1588,In_845);
or U5270 (N_5270,In_1466,In_978);
nand U5271 (N_5271,In_2411,In_1204);
nand U5272 (N_5272,In_127,In_1446);
nor U5273 (N_5273,In_555,In_1579);
nand U5274 (N_5274,In_480,In_1350);
and U5275 (N_5275,In_1938,In_1473);
nand U5276 (N_5276,In_1935,In_141);
nand U5277 (N_5277,In_1539,In_1728);
and U5278 (N_5278,In_1406,In_2445);
or U5279 (N_5279,In_1036,In_998);
or U5280 (N_5280,In_218,In_653);
nor U5281 (N_5281,In_1360,In_2395);
and U5282 (N_5282,In_2028,In_25);
or U5283 (N_5283,In_2499,In_2213);
xor U5284 (N_5284,In_2146,In_269);
nor U5285 (N_5285,In_1826,In_1750);
and U5286 (N_5286,In_637,In_163);
or U5287 (N_5287,In_12,In_2320);
nor U5288 (N_5288,In_2186,In_246);
nand U5289 (N_5289,In_544,In_330);
nor U5290 (N_5290,In_116,In_1144);
or U5291 (N_5291,In_998,In_2100);
or U5292 (N_5292,In_2470,In_1541);
nor U5293 (N_5293,In_2033,In_563);
and U5294 (N_5294,In_1346,In_1253);
xnor U5295 (N_5295,In_1234,In_414);
nor U5296 (N_5296,In_2339,In_1117);
nand U5297 (N_5297,In_1553,In_1307);
and U5298 (N_5298,In_2305,In_1006);
or U5299 (N_5299,In_1321,In_156);
or U5300 (N_5300,In_2059,In_1282);
or U5301 (N_5301,In_2249,In_1080);
nand U5302 (N_5302,In_2047,In_922);
and U5303 (N_5303,In_1677,In_1797);
nand U5304 (N_5304,In_1882,In_1958);
xnor U5305 (N_5305,In_2092,In_770);
or U5306 (N_5306,In_290,In_1377);
xnor U5307 (N_5307,In_872,In_1379);
nor U5308 (N_5308,In_1623,In_1204);
and U5309 (N_5309,In_2176,In_1832);
and U5310 (N_5310,In_717,In_647);
or U5311 (N_5311,In_1055,In_1638);
nor U5312 (N_5312,In_1303,In_1018);
or U5313 (N_5313,In_1728,In_1996);
nor U5314 (N_5314,In_118,In_670);
xor U5315 (N_5315,In_2064,In_1191);
or U5316 (N_5316,In_1878,In_1621);
nand U5317 (N_5317,In_800,In_201);
xor U5318 (N_5318,In_2208,In_662);
nor U5319 (N_5319,In_1610,In_1794);
and U5320 (N_5320,In_2425,In_2481);
or U5321 (N_5321,In_2438,In_1920);
and U5322 (N_5322,In_2366,In_1947);
nor U5323 (N_5323,In_1267,In_78);
or U5324 (N_5324,In_1976,In_2315);
nor U5325 (N_5325,In_1307,In_1481);
xnor U5326 (N_5326,In_942,In_2041);
nor U5327 (N_5327,In_2328,In_1005);
nand U5328 (N_5328,In_2367,In_1974);
nor U5329 (N_5329,In_1313,In_117);
nor U5330 (N_5330,In_1189,In_1443);
xor U5331 (N_5331,In_2219,In_1824);
nor U5332 (N_5332,In_191,In_2479);
nand U5333 (N_5333,In_1004,In_1979);
nand U5334 (N_5334,In_1006,In_2079);
xnor U5335 (N_5335,In_713,In_2229);
or U5336 (N_5336,In_1965,In_645);
xor U5337 (N_5337,In_2342,In_1224);
and U5338 (N_5338,In_640,In_1126);
xnor U5339 (N_5339,In_924,In_2038);
xor U5340 (N_5340,In_690,In_422);
and U5341 (N_5341,In_387,In_2372);
nand U5342 (N_5342,In_515,In_203);
or U5343 (N_5343,In_290,In_463);
xnor U5344 (N_5344,In_1341,In_2321);
nand U5345 (N_5345,In_1835,In_2250);
xor U5346 (N_5346,In_979,In_2254);
xor U5347 (N_5347,In_507,In_1886);
or U5348 (N_5348,In_2489,In_1924);
and U5349 (N_5349,In_558,In_1044);
or U5350 (N_5350,In_2453,In_964);
nand U5351 (N_5351,In_433,In_682);
nand U5352 (N_5352,In_1958,In_885);
and U5353 (N_5353,In_332,In_2402);
nor U5354 (N_5354,In_268,In_2004);
nand U5355 (N_5355,In_1382,In_1999);
nand U5356 (N_5356,In_682,In_1338);
or U5357 (N_5357,In_2036,In_1857);
nor U5358 (N_5358,In_812,In_862);
or U5359 (N_5359,In_795,In_2338);
nand U5360 (N_5360,In_305,In_975);
nand U5361 (N_5361,In_458,In_936);
and U5362 (N_5362,In_497,In_1989);
nor U5363 (N_5363,In_2390,In_2293);
nand U5364 (N_5364,In_392,In_195);
nand U5365 (N_5365,In_1332,In_1202);
nand U5366 (N_5366,In_1398,In_1665);
xor U5367 (N_5367,In_1068,In_26);
nand U5368 (N_5368,In_1514,In_392);
and U5369 (N_5369,In_1900,In_330);
or U5370 (N_5370,In_1992,In_715);
or U5371 (N_5371,In_1722,In_1488);
nor U5372 (N_5372,In_861,In_823);
nor U5373 (N_5373,In_1023,In_2041);
or U5374 (N_5374,In_2115,In_1860);
nand U5375 (N_5375,In_2449,In_2436);
and U5376 (N_5376,In_2067,In_665);
nand U5377 (N_5377,In_2198,In_1194);
nand U5378 (N_5378,In_931,In_1627);
nor U5379 (N_5379,In_871,In_1350);
xnor U5380 (N_5380,In_237,In_370);
nor U5381 (N_5381,In_1252,In_2068);
nor U5382 (N_5382,In_1664,In_2051);
and U5383 (N_5383,In_2401,In_766);
and U5384 (N_5384,In_1667,In_40);
or U5385 (N_5385,In_1545,In_1469);
or U5386 (N_5386,In_69,In_1355);
and U5387 (N_5387,In_839,In_2007);
or U5388 (N_5388,In_2433,In_1988);
or U5389 (N_5389,In_2254,In_43);
xnor U5390 (N_5390,In_228,In_786);
nand U5391 (N_5391,In_556,In_272);
or U5392 (N_5392,In_2026,In_2114);
xnor U5393 (N_5393,In_2391,In_828);
xnor U5394 (N_5394,In_514,In_323);
nand U5395 (N_5395,In_1725,In_635);
and U5396 (N_5396,In_1068,In_910);
nor U5397 (N_5397,In_1716,In_1115);
xnor U5398 (N_5398,In_597,In_1971);
or U5399 (N_5399,In_507,In_1210);
or U5400 (N_5400,In_928,In_2368);
and U5401 (N_5401,In_960,In_530);
xor U5402 (N_5402,In_1412,In_55);
nor U5403 (N_5403,In_1139,In_1339);
nor U5404 (N_5404,In_402,In_2148);
or U5405 (N_5405,In_1126,In_1557);
nor U5406 (N_5406,In_362,In_1803);
and U5407 (N_5407,In_932,In_1634);
nor U5408 (N_5408,In_2403,In_705);
nand U5409 (N_5409,In_2436,In_940);
and U5410 (N_5410,In_876,In_945);
nand U5411 (N_5411,In_2351,In_997);
nor U5412 (N_5412,In_1647,In_1916);
or U5413 (N_5413,In_755,In_131);
nor U5414 (N_5414,In_1316,In_928);
nand U5415 (N_5415,In_97,In_1470);
or U5416 (N_5416,In_2249,In_1000);
xnor U5417 (N_5417,In_2493,In_395);
xor U5418 (N_5418,In_577,In_2080);
nor U5419 (N_5419,In_441,In_1496);
and U5420 (N_5420,In_1652,In_366);
nand U5421 (N_5421,In_698,In_64);
nor U5422 (N_5422,In_2026,In_474);
xor U5423 (N_5423,In_401,In_994);
nand U5424 (N_5424,In_1131,In_852);
xnor U5425 (N_5425,In_933,In_428);
xor U5426 (N_5426,In_1357,In_865);
and U5427 (N_5427,In_2446,In_801);
nor U5428 (N_5428,In_597,In_1385);
nor U5429 (N_5429,In_232,In_61);
xor U5430 (N_5430,In_1213,In_706);
nand U5431 (N_5431,In_310,In_2271);
xor U5432 (N_5432,In_511,In_711);
nor U5433 (N_5433,In_621,In_2362);
or U5434 (N_5434,In_266,In_1593);
nand U5435 (N_5435,In_2013,In_1107);
xnor U5436 (N_5436,In_1739,In_2482);
xor U5437 (N_5437,In_909,In_1904);
and U5438 (N_5438,In_1364,In_111);
or U5439 (N_5439,In_598,In_2217);
nor U5440 (N_5440,In_2395,In_749);
nand U5441 (N_5441,In_810,In_149);
and U5442 (N_5442,In_1283,In_1320);
xnor U5443 (N_5443,In_327,In_1742);
nand U5444 (N_5444,In_1317,In_1287);
nor U5445 (N_5445,In_183,In_354);
nand U5446 (N_5446,In_2490,In_1028);
xor U5447 (N_5447,In_669,In_1050);
nand U5448 (N_5448,In_744,In_2104);
nand U5449 (N_5449,In_2306,In_2310);
and U5450 (N_5450,In_320,In_1006);
xnor U5451 (N_5451,In_1062,In_1498);
xnor U5452 (N_5452,In_1818,In_253);
xnor U5453 (N_5453,In_946,In_1146);
and U5454 (N_5454,In_1785,In_449);
nor U5455 (N_5455,In_836,In_2285);
nor U5456 (N_5456,In_1633,In_18);
nor U5457 (N_5457,In_936,In_2196);
nor U5458 (N_5458,In_1493,In_33);
xor U5459 (N_5459,In_504,In_1575);
or U5460 (N_5460,In_1956,In_2068);
and U5461 (N_5461,In_436,In_1411);
and U5462 (N_5462,In_1255,In_1930);
or U5463 (N_5463,In_2476,In_658);
nor U5464 (N_5464,In_563,In_2249);
and U5465 (N_5465,In_667,In_1849);
or U5466 (N_5466,In_545,In_1151);
and U5467 (N_5467,In_990,In_423);
xnor U5468 (N_5468,In_884,In_2094);
xor U5469 (N_5469,In_1652,In_2141);
nor U5470 (N_5470,In_1011,In_734);
or U5471 (N_5471,In_175,In_735);
and U5472 (N_5472,In_76,In_1284);
xnor U5473 (N_5473,In_1063,In_1914);
xnor U5474 (N_5474,In_120,In_1111);
nor U5475 (N_5475,In_446,In_1869);
nor U5476 (N_5476,In_2303,In_459);
nor U5477 (N_5477,In_2200,In_581);
nand U5478 (N_5478,In_495,In_2090);
and U5479 (N_5479,In_2257,In_567);
nor U5480 (N_5480,In_520,In_1886);
nand U5481 (N_5481,In_2171,In_613);
or U5482 (N_5482,In_627,In_2460);
and U5483 (N_5483,In_2312,In_885);
or U5484 (N_5484,In_1796,In_1652);
xnor U5485 (N_5485,In_2235,In_2217);
and U5486 (N_5486,In_1875,In_950);
xnor U5487 (N_5487,In_2193,In_636);
nor U5488 (N_5488,In_2178,In_996);
nand U5489 (N_5489,In_385,In_1548);
and U5490 (N_5490,In_1197,In_92);
or U5491 (N_5491,In_2336,In_1709);
or U5492 (N_5492,In_1090,In_319);
nand U5493 (N_5493,In_1868,In_85);
xnor U5494 (N_5494,In_1294,In_2375);
xnor U5495 (N_5495,In_655,In_96);
or U5496 (N_5496,In_20,In_1063);
nand U5497 (N_5497,In_534,In_140);
xor U5498 (N_5498,In_1663,In_1829);
nand U5499 (N_5499,In_1614,In_2106);
and U5500 (N_5500,In_1699,In_912);
xor U5501 (N_5501,In_230,In_2409);
or U5502 (N_5502,In_854,In_692);
nand U5503 (N_5503,In_274,In_375);
or U5504 (N_5504,In_1242,In_139);
nand U5505 (N_5505,In_2121,In_856);
nor U5506 (N_5506,In_169,In_914);
and U5507 (N_5507,In_2063,In_2269);
or U5508 (N_5508,In_906,In_182);
or U5509 (N_5509,In_1148,In_2495);
xnor U5510 (N_5510,In_2071,In_21);
or U5511 (N_5511,In_1846,In_910);
nand U5512 (N_5512,In_152,In_773);
nand U5513 (N_5513,In_422,In_2209);
or U5514 (N_5514,In_1641,In_2111);
or U5515 (N_5515,In_1834,In_386);
nand U5516 (N_5516,In_1058,In_2194);
xnor U5517 (N_5517,In_2220,In_2324);
nor U5518 (N_5518,In_105,In_2070);
nor U5519 (N_5519,In_1834,In_60);
nor U5520 (N_5520,In_807,In_2149);
nand U5521 (N_5521,In_605,In_885);
nand U5522 (N_5522,In_1310,In_1499);
and U5523 (N_5523,In_2245,In_1313);
or U5524 (N_5524,In_1466,In_804);
or U5525 (N_5525,In_1678,In_593);
nor U5526 (N_5526,In_831,In_219);
nand U5527 (N_5527,In_1632,In_2367);
and U5528 (N_5528,In_2151,In_291);
or U5529 (N_5529,In_1263,In_1644);
xor U5530 (N_5530,In_664,In_1913);
or U5531 (N_5531,In_1770,In_2297);
or U5532 (N_5532,In_2133,In_66);
and U5533 (N_5533,In_1593,In_2263);
nand U5534 (N_5534,In_1518,In_337);
nand U5535 (N_5535,In_1715,In_1389);
xor U5536 (N_5536,In_761,In_426);
or U5537 (N_5537,In_1647,In_1756);
or U5538 (N_5538,In_837,In_1741);
nor U5539 (N_5539,In_1059,In_2002);
or U5540 (N_5540,In_914,In_56);
nor U5541 (N_5541,In_1989,In_1063);
or U5542 (N_5542,In_1425,In_1318);
xor U5543 (N_5543,In_1114,In_2091);
xnor U5544 (N_5544,In_1308,In_38);
xnor U5545 (N_5545,In_2046,In_948);
nand U5546 (N_5546,In_1413,In_2047);
nor U5547 (N_5547,In_1060,In_403);
xor U5548 (N_5548,In_1421,In_2435);
and U5549 (N_5549,In_391,In_740);
or U5550 (N_5550,In_438,In_2307);
nor U5551 (N_5551,In_8,In_786);
nor U5552 (N_5552,In_1668,In_1446);
and U5553 (N_5553,In_945,In_2175);
and U5554 (N_5554,In_939,In_1880);
and U5555 (N_5555,In_423,In_173);
or U5556 (N_5556,In_2262,In_2332);
nor U5557 (N_5557,In_1897,In_1104);
xnor U5558 (N_5558,In_529,In_245);
nor U5559 (N_5559,In_2443,In_1575);
nand U5560 (N_5560,In_2470,In_1570);
nor U5561 (N_5561,In_1168,In_712);
nor U5562 (N_5562,In_863,In_842);
xnor U5563 (N_5563,In_2400,In_2352);
xor U5564 (N_5564,In_1785,In_718);
nor U5565 (N_5565,In_696,In_1562);
and U5566 (N_5566,In_2111,In_255);
xor U5567 (N_5567,In_2126,In_2089);
or U5568 (N_5568,In_415,In_1386);
or U5569 (N_5569,In_1215,In_2302);
nor U5570 (N_5570,In_1958,In_213);
nand U5571 (N_5571,In_2021,In_362);
or U5572 (N_5572,In_161,In_2180);
nand U5573 (N_5573,In_2228,In_327);
nor U5574 (N_5574,In_1045,In_725);
or U5575 (N_5575,In_1518,In_251);
xor U5576 (N_5576,In_301,In_225);
or U5577 (N_5577,In_692,In_189);
xor U5578 (N_5578,In_1622,In_1658);
or U5579 (N_5579,In_54,In_1576);
and U5580 (N_5580,In_2097,In_1164);
or U5581 (N_5581,In_1601,In_1094);
nor U5582 (N_5582,In_1989,In_1446);
nand U5583 (N_5583,In_1179,In_60);
nor U5584 (N_5584,In_1704,In_2147);
nand U5585 (N_5585,In_1336,In_2355);
nand U5586 (N_5586,In_1910,In_53);
nor U5587 (N_5587,In_1977,In_1002);
xor U5588 (N_5588,In_473,In_1877);
nand U5589 (N_5589,In_1973,In_1391);
nand U5590 (N_5590,In_74,In_864);
xnor U5591 (N_5591,In_2301,In_958);
nor U5592 (N_5592,In_2418,In_65);
nand U5593 (N_5593,In_1659,In_185);
xor U5594 (N_5594,In_437,In_1670);
and U5595 (N_5595,In_1783,In_1434);
nand U5596 (N_5596,In_1006,In_15);
and U5597 (N_5597,In_1602,In_857);
nand U5598 (N_5598,In_1501,In_123);
nor U5599 (N_5599,In_1181,In_2017);
xnor U5600 (N_5600,In_42,In_2381);
nand U5601 (N_5601,In_1474,In_1760);
nand U5602 (N_5602,In_2190,In_875);
nor U5603 (N_5603,In_2045,In_2067);
and U5604 (N_5604,In_206,In_106);
xnor U5605 (N_5605,In_1784,In_1066);
nor U5606 (N_5606,In_878,In_864);
nor U5607 (N_5607,In_878,In_1747);
xnor U5608 (N_5608,In_1266,In_1004);
nor U5609 (N_5609,In_511,In_333);
xnor U5610 (N_5610,In_358,In_1500);
and U5611 (N_5611,In_2193,In_2121);
or U5612 (N_5612,In_935,In_2271);
xnor U5613 (N_5613,In_2167,In_736);
xnor U5614 (N_5614,In_1417,In_756);
xnor U5615 (N_5615,In_1304,In_753);
xnor U5616 (N_5616,In_1807,In_918);
or U5617 (N_5617,In_188,In_798);
nor U5618 (N_5618,In_2363,In_1165);
or U5619 (N_5619,In_2200,In_2256);
or U5620 (N_5620,In_1783,In_1925);
or U5621 (N_5621,In_1998,In_172);
and U5622 (N_5622,In_813,In_2304);
nand U5623 (N_5623,In_2251,In_588);
xnor U5624 (N_5624,In_1488,In_249);
nand U5625 (N_5625,In_813,In_2309);
nor U5626 (N_5626,In_1521,In_1421);
or U5627 (N_5627,In_172,In_2196);
xor U5628 (N_5628,In_2365,In_2319);
or U5629 (N_5629,In_1245,In_687);
nand U5630 (N_5630,In_658,In_1384);
and U5631 (N_5631,In_1766,In_1717);
nand U5632 (N_5632,In_2081,In_2132);
and U5633 (N_5633,In_244,In_463);
nor U5634 (N_5634,In_1273,In_1708);
and U5635 (N_5635,In_939,In_271);
or U5636 (N_5636,In_996,In_375);
and U5637 (N_5637,In_30,In_1176);
or U5638 (N_5638,In_2197,In_469);
or U5639 (N_5639,In_2439,In_1271);
xnor U5640 (N_5640,In_634,In_1130);
nand U5641 (N_5641,In_530,In_1850);
nor U5642 (N_5642,In_1783,In_1779);
or U5643 (N_5643,In_1739,In_1423);
nand U5644 (N_5644,In_248,In_1185);
and U5645 (N_5645,In_1087,In_164);
xor U5646 (N_5646,In_2018,In_1423);
and U5647 (N_5647,In_1455,In_68);
nor U5648 (N_5648,In_852,In_658);
xnor U5649 (N_5649,In_61,In_70);
or U5650 (N_5650,In_1127,In_1661);
or U5651 (N_5651,In_2070,In_993);
nor U5652 (N_5652,In_709,In_1760);
nor U5653 (N_5653,In_111,In_1803);
xnor U5654 (N_5654,In_307,In_1425);
and U5655 (N_5655,In_2395,In_1321);
or U5656 (N_5656,In_1476,In_2332);
nor U5657 (N_5657,In_2102,In_162);
or U5658 (N_5658,In_1508,In_296);
nor U5659 (N_5659,In_111,In_990);
nor U5660 (N_5660,In_559,In_841);
and U5661 (N_5661,In_2357,In_672);
xnor U5662 (N_5662,In_2129,In_423);
and U5663 (N_5663,In_1427,In_613);
nor U5664 (N_5664,In_2474,In_2124);
or U5665 (N_5665,In_602,In_1170);
or U5666 (N_5666,In_1277,In_860);
or U5667 (N_5667,In_1323,In_1784);
nor U5668 (N_5668,In_977,In_44);
nor U5669 (N_5669,In_2183,In_685);
nand U5670 (N_5670,In_2150,In_2350);
or U5671 (N_5671,In_1347,In_359);
nand U5672 (N_5672,In_770,In_1284);
or U5673 (N_5673,In_1191,In_1166);
xor U5674 (N_5674,In_598,In_171);
nand U5675 (N_5675,In_2420,In_940);
and U5676 (N_5676,In_2422,In_920);
nor U5677 (N_5677,In_193,In_2031);
nand U5678 (N_5678,In_181,In_1564);
and U5679 (N_5679,In_1130,In_1227);
xor U5680 (N_5680,In_537,In_1598);
and U5681 (N_5681,In_2245,In_2002);
or U5682 (N_5682,In_1102,In_477);
or U5683 (N_5683,In_1773,In_1550);
xnor U5684 (N_5684,In_835,In_639);
xor U5685 (N_5685,In_163,In_2191);
and U5686 (N_5686,In_1106,In_1173);
nand U5687 (N_5687,In_620,In_1337);
and U5688 (N_5688,In_139,In_2168);
nand U5689 (N_5689,In_2349,In_878);
nor U5690 (N_5690,In_107,In_339);
and U5691 (N_5691,In_169,In_1336);
xor U5692 (N_5692,In_916,In_1453);
and U5693 (N_5693,In_2365,In_823);
or U5694 (N_5694,In_327,In_1219);
nand U5695 (N_5695,In_929,In_557);
or U5696 (N_5696,In_704,In_1112);
nand U5697 (N_5697,In_1155,In_106);
nor U5698 (N_5698,In_1610,In_2052);
nor U5699 (N_5699,In_1294,In_2484);
nor U5700 (N_5700,In_2133,In_1737);
or U5701 (N_5701,In_963,In_2021);
xnor U5702 (N_5702,In_179,In_1544);
or U5703 (N_5703,In_23,In_1886);
xor U5704 (N_5704,In_441,In_2075);
or U5705 (N_5705,In_2302,In_2156);
nand U5706 (N_5706,In_1023,In_622);
and U5707 (N_5707,In_782,In_1733);
or U5708 (N_5708,In_758,In_1298);
nor U5709 (N_5709,In_732,In_938);
or U5710 (N_5710,In_650,In_1545);
or U5711 (N_5711,In_1761,In_340);
and U5712 (N_5712,In_864,In_299);
nand U5713 (N_5713,In_42,In_38);
or U5714 (N_5714,In_2308,In_2120);
and U5715 (N_5715,In_2489,In_1542);
nand U5716 (N_5716,In_2246,In_814);
nor U5717 (N_5717,In_146,In_950);
or U5718 (N_5718,In_1943,In_238);
nor U5719 (N_5719,In_1070,In_974);
or U5720 (N_5720,In_1243,In_371);
nor U5721 (N_5721,In_1462,In_220);
nand U5722 (N_5722,In_1675,In_2181);
nand U5723 (N_5723,In_2282,In_2225);
and U5724 (N_5724,In_317,In_440);
nor U5725 (N_5725,In_466,In_366);
and U5726 (N_5726,In_844,In_1386);
and U5727 (N_5727,In_1040,In_1653);
or U5728 (N_5728,In_1091,In_782);
or U5729 (N_5729,In_5,In_2300);
nand U5730 (N_5730,In_494,In_2091);
nor U5731 (N_5731,In_1651,In_1826);
nor U5732 (N_5732,In_983,In_1627);
or U5733 (N_5733,In_1604,In_1659);
nand U5734 (N_5734,In_1762,In_263);
or U5735 (N_5735,In_470,In_349);
nor U5736 (N_5736,In_1670,In_1146);
xor U5737 (N_5737,In_1552,In_363);
and U5738 (N_5738,In_723,In_128);
xor U5739 (N_5739,In_924,In_698);
nor U5740 (N_5740,In_2306,In_1181);
nor U5741 (N_5741,In_572,In_1722);
or U5742 (N_5742,In_763,In_1154);
and U5743 (N_5743,In_569,In_512);
nor U5744 (N_5744,In_2393,In_489);
or U5745 (N_5745,In_1271,In_1045);
nor U5746 (N_5746,In_2172,In_1844);
and U5747 (N_5747,In_667,In_1709);
xor U5748 (N_5748,In_1370,In_638);
and U5749 (N_5749,In_326,In_1028);
and U5750 (N_5750,In_1607,In_660);
xor U5751 (N_5751,In_921,In_1525);
nand U5752 (N_5752,In_1721,In_648);
nand U5753 (N_5753,In_1701,In_1456);
xor U5754 (N_5754,In_176,In_1125);
or U5755 (N_5755,In_759,In_398);
nand U5756 (N_5756,In_92,In_1841);
and U5757 (N_5757,In_1831,In_781);
and U5758 (N_5758,In_2267,In_1980);
and U5759 (N_5759,In_1925,In_1533);
xor U5760 (N_5760,In_919,In_1433);
and U5761 (N_5761,In_1252,In_1768);
xnor U5762 (N_5762,In_455,In_710);
and U5763 (N_5763,In_2186,In_1527);
nor U5764 (N_5764,In_99,In_602);
nand U5765 (N_5765,In_1706,In_1587);
nand U5766 (N_5766,In_735,In_1989);
nand U5767 (N_5767,In_992,In_450);
nor U5768 (N_5768,In_2239,In_2469);
xnor U5769 (N_5769,In_227,In_1473);
nor U5770 (N_5770,In_2436,In_693);
nand U5771 (N_5771,In_1941,In_1737);
and U5772 (N_5772,In_1794,In_2476);
nand U5773 (N_5773,In_1824,In_1725);
nor U5774 (N_5774,In_1873,In_2210);
and U5775 (N_5775,In_298,In_593);
or U5776 (N_5776,In_2005,In_2388);
or U5777 (N_5777,In_110,In_798);
nand U5778 (N_5778,In_161,In_627);
nor U5779 (N_5779,In_2024,In_2357);
xor U5780 (N_5780,In_1955,In_1626);
nor U5781 (N_5781,In_1630,In_228);
xnor U5782 (N_5782,In_2328,In_1343);
xnor U5783 (N_5783,In_1391,In_1118);
and U5784 (N_5784,In_1405,In_2452);
xnor U5785 (N_5785,In_1847,In_756);
or U5786 (N_5786,In_535,In_99);
nand U5787 (N_5787,In_83,In_1890);
or U5788 (N_5788,In_981,In_2245);
or U5789 (N_5789,In_398,In_2338);
or U5790 (N_5790,In_1432,In_1588);
nor U5791 (N_5791,In_1401,In_2091);
and U5792 (N_5792,In_2304,In_2156);
xor U5793 (N_5793,In_1987,In_405);
nor U5794 (N_5794,In_2171,In_647);
nor U5795 (N_5795,In_1407,In_655);
and U5796 (N_5796,In_498,In_1648);
nand U5797 (N_5797,In_476,In_78);
and U5798 (N_5798,In_1914,In_414);
or U5799 (N_5799,In_973,In_2270);
nor U5800 (N_5800,In_2182,In_932);
and U5801 (N_5801,In_1917,In_1145);
nand U5802 (N_5802,In_915,In_2488);
or U5803 (N_5803,In_1837,In_763);
nand U5804 (N_5804,In_1652,In_2195);
and U5805 (N_5805,In_641,In_1863);
and U5806 (N_5806,In_2235,In_6);
xor U5807 (N_5807,In_126,In_1551);
xnor U5808 (N_5808,In_1261,In_2380);
nand U5809 (N_5809,In_109,In_183);
nor U5810 (N_5810,In_374,In_1663);
nand U5811 (N_5811,In_1521,In_1747);
xnor U5812 (N_5812,In_1023,In_1263);
nor U5813 (N_5813,In_978,In_1619);
and U5814 (N_5814,In_655,In_1273);
nor U5815 (N_5815,In_1035,In_1189);
xnor U5816 (N_5816,In_1312,In_818);
and U5817 (N_5817,In_2400,In_243);
nor U5818 (N_5818,In_1232,In_1600);
nand U5819 (N_5819,In_1572,In_1040);
and U5820 (N_5820,In_1580,In_1415);
and U5821 (N_5821,In_393,In_638);
xor U5822 (N_5822,In_1503,In_235);
and U5823 (N_5823,In_2438,In_1703);
and U5824 (N_5824,In_626,In_417);
nor U5825 (N_5825,In_1858,In_1393);
xor U5826 (N_5826,In_1699,In_575);
nor U5827 (N_5827,In_1859,In_228);
and U5828 (N_5828,In_1505,In_2145);
or U5829 (N_5829,In_1482,In_929);
xor U5830 (N_5830,In_380,In_2128);
or U5831 (N_5831,In_645,In_267);
and U5832 (N_5832,In_2284,In_1628);
xnor U5833 (N_5833,In_17,In_952);
and U5834 (N_5834,In_631,In_2283);
xnor U5835 (N_5835,In_1991,In_1380);
and U5836 (N_5836,In_1937,In_645);
nand U5837 (N_5837,In_1043,In_1647);
nand U5838 (N_5838,In_2023,In_470);
nor U5839 (N_5839,In_449,In_2156);
xor U5840 (N_5840,In_949,In_578);
nor U5841 (N_5841,In_2090,In_782);
nor U5842 (N_5842,In_763,In_911);
and U5843 (N_5843,In_2366,In_89);
and U5844 (N_5844,In_965,In_647);
nor U5845 (N_5845,In_1453,In_1281);
xor U5846 (N_5846,In_2453,In_228);
nand U5847 (N_5847,In_170,In_1358);
nor U5848 (N_5848,In_498,In_1368);
xor U5849 (N_5849,In_800,In_595);
nand U5850 (N_5850,In_2196,In_669);
xor U5851 (N_5851,In_265,In_951);
nand U5852 (N_5852,In_1246,In_2008);
nand U5853 (N_5853,In_117,In_511);
xor U5854 (N_5854,In_246,In_23);
nor U5855 (N_5855,In_1817,In_1778);
or U5856 (N_5856,In_1998,In_1058);
and U5857 (N_5857,In_2258,In_2408);
nor U5858 (N_5858,In_1635,In_682);
or U5859 (N_5859,In_983,In_1017);
nand U5860 (N_5860,In_1393,In_2192);
nand U5861 (N_5861,In_192,In_1473);
xnor U5862 (N_5862,In_1749,In_880);
nor U5863 (N_5863,In_344,In_166);
nor U5864 (N_5864,In_405,In_1765);
nor U5865 (N_5865,In_1159,In_1235);
nand U5866 (N_5866,In_995,In_388);
nand U5867 (N_5867,In_1527,In_698);
xor U5868 (N_5868,In_912,In_800);
nor U5869 (N_5869,In_1883,In_1599);
nand U5870 (N_5870,In_1344,In_1061);
nand U5871 (N_5871,In_1169,In_827);
nand U5872 (N_5872,In_1478,In_906);
or U5873 (N_5873,In_2361,In_2060);
or U5874 (N_5874,In_1478,In_1604);
and U5875 (N_5875,In_120,In_2485);
xor U5876 (N_5876,In_2367,In_2390);
or U5877 (N_5877,In_2390,In_1283);
or U5878 (N_5878,In_1940,In_489);
and U5879 (N_5879,In_1053,In_1244);
nand U5880 (N_5880,In_1233,In_2047);
xnor U5881 (N_5881,In_738,In_2047);
nor U5882 (N_5882,In_1651,In_2264);
nand U5883 (N_5883,In_2258,In_271);
xnor U5884 (N_5884,In_1233,In_636);
xor U5885 (N_5885,In_2029,In_1955);
nand U5886 (N_5886,In_1705,In_2104);
xor U5887 (N_5887,In_1181,In_569);
or U5888 (N_5888,In_675,In_546);
nor U5889 (N_5889,In_1822,In_62);
xor U5890 (N_5890,In_198,In_0);
or U5891 (N_5891,In_2481,In_1840);
nand U5892 (N_5892,In_1431,In_1207);
nor U5893 (N_5893,In_2050,In_1883);
nor U5894 (N_5894,In_931,In_100);
and U5895 (N_5895,In_1094,In_1116);
nand U5896 (N_5896,In_282,In_455);
nand U5897 (N_5897,In_2420,In_2478);
xor U5898 (N_5898,In_595,In_1507);
xnor U5899 (N_5899,In_1285,In_472);
nand U5900 (N_5900,In_1076,In_1381);
nor U5901 (N_5901,In_1366,In_1358);
nor U5902 (N_5902,In_883,In_2287);
nand U5903 (N_5903,In_1337,In_411);
and U5904 (N_5904,In_1887,In_1939);
nand U5905 (N_5905,In_17,In_1445);
and U5906 (N_5906,In_442,In_2078);
nand U5907 (N_5907,In_1652,In_558);
or U5908 (N_5908,In_1735,In_893);
nor U5909 (N_5909,In_938,In_960);
nor U5910 (N_5910,In_2108,In_1972);
and U5911 (N_5911,In_2304,In_2477);
nand U5912 (N_5912,In_2074,In_1408);
and U5913 (N_5913,In_904,In_285);
nor U5914 (N_5914,In_895,In_2481);
or U5915 (N_5915,In_239,In_1785);
nor U5916 (N_5916,In_1167,In_818);
xor U5917 (N_5917,In_1320,In_809);
nor U5918 (N_5918,In_33,In_956);
nor U5919 (N_5919,In_2378,In_2184);
nor U5920 (N_5920,In_1570,In_1098);
nor U5921 (N_5921,In_266,In_1670);
nand U5922 (N_5922,In_91,In_1766);
xnor U5923 (N_5923,In_1622,In_76);
nand U5924 (N_5924,In_446,In_2291);
xnor U5925 (N_5925,In_1104,In_629);
and U5926 (N_5926,In_1993,In_1442);
or U5927 (N_5927,In_772,In_530);
or U5928 (N_5928,In_941,In_285);
nand U5929 (N_5929,In_1979,In_971);
and U5930 (N_5930,In_1872,In_1590);
xnor U5931 (N_5931,In_1894,In_902);
xor U5932 (N_5932,In_164,In_1798);
or U5933 (N_5933,In_1414,In_2435);
nor U5934 (N_5934,In_867,In_774);
and U5935 (N_5935,In_2339,In_1402);
nor U5936 (N_5936,In_480,In_1696);
xnor U5937 (N_5937,In_1321,In_1987);
xor U5938 (N_5938,In_1521,In_656);
or U5939 (N_5939,In_2292,In_1423);
and U5940 (N_5940,In_1810,In_1395);
and U5941 (N_5941,In_1798,In_1519);
xor U5942 (N_5942,In_851,In_623);
xnor U5943 (N_5943,In_372,In_435);
or U5944 (N_5944,In_265,In_1620);
or U5945 (N_5945,In_1076,In_427);
nand U5946 (N_5946,In_2080,In_1412);
and U5947 (N_5947,In_977,In_185);
nor U5948 (N_5948,In_2415,In_1144);
nand U5949 (N_5949,In_1867,In_687);
and U5950 (N_5950,In_2063,In_907);
and U5951 (N_5951,In_2423,In_2132);
and U5952 (N_5952,In_53,In_2178);
nand U5953 (N_5953,In_1928,In_334);
xor U5954 (N_5954,In_1719,In_861);
or U5955 (N_5955,In_727,In_1873);
xnor U5956 (N_5956,In_2048,In_1538);
xor U5957 (N_5957,In_2158,In_1370);
nor U5958 (N_5958,In_189,In_1423);
nor U5959 (N_5959,In_2155,In_587);
or U5960 (N_5960,In_782,In_2151);
nor U5961 (N_5961,In_2118,In_2414);
or U5962 (N_5962,In_164,In_1398);
or U5963 (N_5963,In_1601,In_751);
nor U5964 (N_5964,In_1406,In_464);
and U5965 (N_5965,In_1084,In_206);
and U5966 (N_5966,In_822,In_2383);
xnor U5967 (N_5967,In_852,In_1406);
nand U5968 (N_5968,In_1485,In_2301);
xnor U5969 (N_5969,In_1692,In_705);
or U5970 (N_5970,In_1588,In_477);
or U5971 (N_5971,In_435,In_295);
nand U5972 (N_5972,In_1538,In_238);
xor U5973 (N_5973,In_1520,In_1722);
nor U5974 (N_5974,In_2313,In_1059);
xor U5975 (N_5975,In_945,In_1795);
and U5976 (N_5976,In_473,In_807);
and U5977 (N_5977,In_810,In_1539);
and U5978 (N_5978,In_892,In_876);
xor U5979 (N_5979,In_897,In_3);
nand U5980 (N_5980,In_1656,In_159);
and U5981 (N_5981,In_2044,In_812);
nand U5982 (N_5982,In_13,In_1103);
and U5983 (N_5983,In_1141,In_1673);
nor U5984 (N_5984,In_1817,In_131);
nand U5985 (N_5985,In_2290,In_1296);
or U5986 (N_5986,In_1225,In_2473);
or U5987 (N_5987,In_1623,In_882);
nand U5988 (N_5988,In_1469,In_2209);
nor U5989 (N_5989,In_808,In_1471);
xor U5990 (N_5990,In_152,In_1258);
nor U5991 (N_5991,In_1319,In_1591);
nor U5992 (N_5992,In_2433,In_97);
and U5993 (N_5993,In_1077,In_2475);
xnor U5994 (N_5994,In_1986,In_511);
nand U5995 (N_5995,In_2384,In_1745);
or U5996 (N_5996,In_873,In_111);
xor U5997 (N_5997,In_2032,In_388);
nor U5998 (N_5998,In_2284,In_861);
xnor U5999 (N_5999,In_928,In_1260);
nand U6000 (N_6000,In_2348,In_1577);
and U6001 (N_6001,In_1227,In_1400);
nand U6002 (N_6002,In_1790,In_1106);
nand U6003 (N_6003,In_1819,In_1111);
nor U6004 (N_6004,In_290,In_1772);
and U6005 (N_6005,In_2038,In_1019);
and U6006 (N_6006,In_284,In_2415);
nand U6007 (N_6007,In_836,In_2431);
and U6008 (N_6008,In_590,In_422);
xor U6009 (N_6009,In_1645,In_507);
xor U6010 (N_6010,In_268,In_1941);
xor U6011 (N_6011,In_1252,In_1864);
nor U6012 (N_6012,In_905,In_2260);
nand U6013 (N_6013,In_840,In_1911);
or U6014 (N_6014,In_178,In_1892);
and U6015 (N_6015,In_1345,In_699);
nor U6016 (N_6016,In_2078,In_1881);
or U6017 (N_6017,In_580,In_1138);
and U6018 (N_6018,In_720,In_1041);
nand U6019 (N_6019,In_683,In_218);
xor U6020 (N_6020,In_1474,In_612);
xor U6021 (N_6021,In_2005,In_1927);
xnor U6022 (N_6022,In_1058,In_1233);
or U6023 (N_6023,In_399,In_2378);
and U6024 (N_6024,In_1759,In_1591);
nor U6025 (N_6025,In_599,In_947);
xnor U6026 (N_6026,In_1470,In_762);
and U6027 (N_6027,In_1943,In_502);
and U6028 (N_6028,In_2174,In_361);
and U6029 (N_6029,In_448,In_357);
and U6030 (N_6030,In_2317,In_1572);
or U6031 (N_6031,In_348,In_2141);
nor U6032 (N_6032,In_1790,In_213);
and U6033 (N_6033,In_1926,In_899);
nor U6034 (N_6034,In_2154,In_799);
xor U6035 (N_6035,In_2215,In_272);
nand U6036 (N_6036,In_573,In_402);
nor U6037 (N_6037,In_1050,In_2014);
xor U6038 (N_6038,In_1163,In_475);
nor U6039 (N_6039,In_201,In_862);
nor U6040 (N_6040,In_1707,In_2190);
nand U6041 (N_6041,In_1484,In_2355);
or U6042 (N_6042,In_361,In_225);
and U6043 (N_6043,In_2123,In_256);
nand U6044 (N_6044,In_1982,In_1636);
nand U6045 (N_6045,In_1843,In_11);
nand U6046 (N_6046,In_2344,In_2251);
and U6047 (N_6047,In_1234,In_2202);
nor U6048 (N_6048,In_2156,In_2436);
nand U6049 (N_6049,In_614,In_705);
nor U6050 (N_6050,In_521,In_2330);
nand U6051 (N_6051,In_1062,In_1450);
nand U6052 (N_6052,In_414,In_1687);
or U6053 (N_6053,In_285,In_991);
nand U6054 (N_6054,In_321,In_521);
xor U6055 (N_6055,In_183,In_1321);
xnor U6056 (N_6056,In_667,In_592);
xnor U6057 (N_6057,In_297,In_2107);
nor U6058 (N_6058,In_40,In_2392);
nand U6059 (N_6059,In_2416,In_1991);
nand U6060 (N_6060,In_693,In_1770);
and U6061 (N_6061,In_1147,In_1121);
and U6062 (N_6062,In_832,In_2204);
nand U6063 (N_6063,In_283,In_1658);
xor U6064 (N_6064,In_119,In_2035);
xor U6065 (N_6065,In_1750,In_314);
nand U6066 (N_6066,In_804,In_1376);
and U6067 (N_6067,In_1269,In_725);
xnor U6068 (N_6068,In_1504,In_738);
and U6069 (N_6069,In_1942,In_681);
xor U6070 (N_6070,In_1101,In_577);
xnor U6071 (N_6071,In_1892,In_2277);
nand U6072 (N_6072,In_973,In_403);
nor U6073 (N_6073,In_2282,In_2062);
and U6074 (N_6074,In_1034,In_1942);
xor U6075 (N_6075,In_1671,In_1131);
nand U6076 (N_6076,In_200,In_115);
nor U6077 (N_6077,In_18,In_1576);
xnor U6078 (N_6078,In_443,In_336);
xor U6079 (N_6079,In_1376,In_1723);
xnor U6080 (N_6080,In_1261,In_1970);
or U6081 (N_6081,In_1410,In_61);
nor U6082 (N_6082,In_1411,In_1448);
or U6083 (N_6083,In_2445,In_1077);
nor U6084 (N_6084,In_231,In_1519);
nand U6085 (N_6085,In_2198,In_555);
xor U6086 (N_6086,In_2305,In_1503);
and U6087 (N_6087,In_2241,In_42);
xor U6088 (N_6088,In_1819,In_2218);
nor U6089 (N_6089,In_2395,In_2170);
nor U6090 (N_6090,In_416,In_176);
nand U6091 (N_6091,In_810,In_792);
nand U6092 (N_6092,In_1324,In_531);
nand U6093 (N_6093,In_1783,In_328);
nand U6094 (N_6094,In_995,In_2267);
nor U6095 (N_6095,In_158,In_1798);
xor U6096 (N_6096,In_136,In_878);
xnor U6097 (N_6097,In_1660,In_1214);
nand U6098 (N_6098,In_857,In_1819);
nand U6099 (N_6099,In_1322,In_950);
and U6100 (N_6100,In_0,In_2195);
nor U6101 (N_6101,In_1977,In_364);
or U6102 (N_6102,In_1899,In_2151);
and U6103 (N_6103,In_739,In_1236);
nand U6104 (N_6104,In_1582,In_885);
nor U6105 (N_6105,In_1792,In_169);
and U6106 (N_6106,In_782,In_310);
nand U6107 (N_6107,In_1811,In_113);
and U6108 (N_6108,In_2183,In_304);
and U6109 (N_6109,In_1848,In_1872);
or U6110 (N_6110,In_1282,In_399);
or U6111 (N_6111,In_1518,In_120);
xnor U6112 (N_6112,In_161,In_1578);
nand U6113 (N_6113,In_2263,In_181);
and U6114 (N_6114,In_657,In_2143);
and U6115 (N_6115,In_469,In_2377);
xnor U6116 (N_6116,In_1767,In_1596);
nand U6117 (N_6117,In_1105,In_2046);
and U6118 (N_6118,In_678,In_1605);
or U6119 (N_6119,In_793,In_588);
or U6120 (N_6120,In_745,In_1635);
and U6121 (N_6121,In_1501,In_453);
nand U6122 (N_6122,In_1998,In_1331);
nand U6123 (N_6123,In_1431,In_2487);
nand U6124 (N_6124,In_1694,In_1615);
xnor U6125 (N_6125,In_2107,In_1029);
or U6126 (N_6126,In_1794,In_511);
nand U6127 (N_6127,In_1822,In_128);
or U6128 (N_6128,In_2155,In_1091);
nor U6129 (N_6129,In_777,In_964);
xnor U6130 (N_6130,In_1688,In_190);
nand U6131 (N_6131,In_884,In_578);
and U6132 (N_6132,In_2169,In_850);
and U6133 (N_6133,In_100,In_305);
or U6134 (N_6134,In_2095,In_2327);
nand U6135 (N_6135,In_1953,In_802);
nor U6136 (N_6136,In_1990,In_888);
and U6137 (N_6137,In_79,In_1262);
nand U6138 (N_6138,In_1639,In_1809);
nor U6139 (N_6139,In_979,In_827);
or U6140 (N_6140,In_2390,In_1439);
xnor U6141 (N_6141,In_1293,In_1126);
nor U6142 (N_6142,In_1313,In_540);
and U6143 (N_6143,In_673,In_2296);
nand U6144 (N_6144,In_2326,In_293);
nor U6145 (N_6145,In_472,In_948);
nor U6146 (N_6146,In_2195,In_194);
or U6147 (N_6147,In_143,In_1861);
nand U6148 (N_6148,In_1219,In_1297);
nor U6149 (N_6149,In_1309,In_2462);
or U6150 (N_6150,In_649,In_887);
and U6151 (N_6151,In_958,In_307);
nor U6152 (N_6152,In_2192,In_1850);
nor U6153 (N_6153,In_668,In_931);
xor U6154 (N_6154,In_339,In_1285);
nand U6155 (N_6155,In_2014,In_2375);
xor U6156 (N_6156,In_1822,In_1001);
nand U6157 (N_6157,In_508,In_1394);
or U6158 (N_6158,In_2267,In_2452);
xor U6159 (N_6159,In_1261,In_1513);
nand U6160 (N_6160,In_1515,In_784);
xnor U6161 (N_6161,In_2038,In_291);
nor U6162 (N_6162,In_902,In_1015);
and U6163 (N_6163,In_1152,In_511);
nand U6164 (N_6164,In_2133,In_1733);
nand U6165 (N_6165,In_1816,In_5);
nand U6166 (N_6166,In_2270,In_1027);
nor U6167 (N_6167,In_2093,In_1489);
nand U6168 (N_6168,In_2265,In_1878);
xor U6169 (N_6169,In_2326,In_2098);
xnor U6170 (N_6170,In_1111,In_2370);
nor U6171 (N_6171,In_1647,In_728);
nor U6172 (N_6172,In_1452,In_1356);
and U6173 (N_6173,In_2433,In_2447);
nor U6174 (N_6174,In_724,In_1382);
nor U6175 (N_6175,In_2045,In_179);
or U6176 (N_6176,In_2105,In_799);
nand U6177 (N_6177,In_1907,In_877);
xnor U6178 (N_6178,In_1027,In_186);
nand U6179 (N_6179,In_734,In_913);
or U6180 (N_6180,In_2072,In_363);
xnor U6181 (N_6181,In_262,In_1953);
nor U6182 (N_6182,In_715,In_931);
or U6183 (N_6183,In_1206,In_577);
xnor U6184 (N_6184,In_1739,In_2120);
xnor U6185 (N_6185,In_677,In_27);
or U6186 (N_6186,In_1611,In_1747);
nor U6187 (N_6187,In_1022,In_1105);
or U6188 (N_6188,In_2214,In_234);
nor U6189 (N_6189,In_2230,In_2422);
nor U6190 (N_6190,In_2121,In_112);
or U6191 (N_6191,In_1735,In_2492);
xnor U6192 (N_6192,In_1424,In_1935);
or U6193 (N_6193,In_333,In_1051);
nor U6194 (N_6194,In_367,In_2422);
and U6195 (N_6195,In_141,In_310);
nand U6196 (N_6196,In_1057,In_235);
xor U6197 (N_6197,In_213,In_1441);
nand U6198 (N_6198,In_1437,In_1630);
or U6199 (N_6199,In_994,In_1345);
nor U6200 (N_6200,In_2196,In_2368);
or U6201 (N_6201,In_1715,In_1792);
xor U6202 (N_6202,In_154,In_1696);
nand U6203 (N_6203,In_2370,In_78);
and U6204 (N_6204,In_1247,In_1717);
nor U6205 (N_6205,In_2434,In_2451);
nand U6206 (N_6206,In_1588,In_934);
nor U6207 (N_6207,In_30,In_1834);
nor U6208 (N_6208,In_1898,In_416);
nor U6209 (N_6209,In_1472,In_554);
nand U6210 (N_6210,In_948,In_1717);
nand U6211 (N_6211,In_2152,In_652);
nor U6212 (N_6212,In_1227,In_2206);
nand U6213 (N_6213,In_2464,In_1987);
xor U6214 (N_6214,In_1465,In_810);
nor U6215 (N_6215,In_1669,In_1685);
xor U6216 (N_6216,In_2058,In_2473);
and U6217 (N_6217,In_788,In_157);
nor U6218 (N_6218,In_1050,In_989);
xnor U6219 (N_6219,In_190,In_576);
nand U6220 (N_6220,In_114,In_291);
nor U6221 (N_6221,In_1733,In_2472);
or U6222 (N_6222,In_2236,In_196);
nor U6223 (N_6223,In_1790,In_1472);
or U6224 (N_6224,In_64,In_2119);
nand U6225 (N_6225,In_1636,In_1543);
nand U6226 (N_6226,In_796,In_1059);
nor U6227 (N_6227,In_648,In_144);
or U6228 (N_6228,In_309,In_2399);
and U6229 (N_6229,In_944,In_839);
xnor U6230 (N_6230,In_73,In_1351);
nand U6231 (N_6231,In_1558,In_1016);
nor U6232 (N_6232,In_2377,In_1345);
or U6233 (N_6233,In_1298,In_1150);
and U6234 (N_6234,In_2370,In_365);
nor U6235 (N_6235,In_1911,In_138);
and U6236 (N_6236,In_1620,In_931);
xor U6237 (N_6237,In_1484,In_756);
nand U6238 (N_6238,In_544,In_655);
or U6239 (N_6239,In_245,In_1214);
or U6240 (N_6240,In_1722,In_274);
xnor U6241 (N_6241,In_2235,In_1518);
and U6242 (N_6242,In_1656,In_533);
and U6243 (N_6243,In_2230,In_1343);
or U6244 (N_6244,In_252,In_1165);
or U6245 (N_6245,In_34,In_1961);
or U6246 (N_6246,In_1762,In_1918);
nand U6247 (N_6247,In_373,In_2092);
xor U6248 (N_6248,In_2085,In_267);
and U6249 (N_6249,In_2158,In_103);
nand U6250 (N_6250,N_5195,N_4861);
and U6251 (N_6251,N_3436,N_5465);
or U6252 (N_6252,N_136,N_2413);
xor U6253 (N_6253,N_3109,N_5709);
xnor U6254 (N_6254,N_44,N_3459);
nor U6255 (N_6255,N_1290,N_2773);
xor U6256 (N_6256,N_5668,N_3418);
and U6257 (N_6257,N_2749,N_3449);
and U6258 (N_6258,N_1331,N_1791);
and U6259 (N_6259,N_5513,N_5415);
nor U6260 (N_6260,N_3899,N_5702);
nand U6261 (N_6261,N_4267,N_5205);
nand U6262 (N_6262,N_276,N_797);
or U6263 (N_6263,N_3304,N_5834);
nand U6264 (N_6264,N_3918,N_807);
or U6265 (N_6265,N_357,N_1536);
xor U6266 (N_6266,N_3367,N_5231);
or U6267 (N_6267,N_370,N_3249);
xor U6268 (N_6268,N_4795,N_4057);
nand U6269 (N_6269,N_509,N_4231);
or U6270 (N_6270,N_606,N_5487);
nor U6271 (N_6271,N_4473,N_2448);
nor U6272 (N_6272,N_2213,N_1169);
nor U6273 (N_6273,N_6169,N_5295);
xnor U6274 (N_6274,N_5457,N_5896);
and U6275 (N_6275,N_474,N_5237);
xor U6276 (N_6276,N_2732,N_5555);
nor U6277 (N_6277,N_1888,N_5478);
nand U6278 (N_6278,N_2912,N_4818);
nor U6279 (N_6279,N_3706,N_5197);
nor U6280 (N_6280,N_892,N_2753);
xor U6281 (N_6281,N_3906,N_5249);
nor U6282 (N_6282,N_5637,N_5119);
xor U6283 (N_6283,N_2716,N_91);
nand U6284 (N_6284,N_5945,N_1292);
nor U6285 (N_6285,N_5845,N_225);
and U6286 (N_6286,N_2065,N_1371);
or U6287 (N_6287,N_2000,N_5813);
xnor U6288 (N_6288,N_3802,N_6086);
nor U6289 (N_6289,N_1058,N_3402);
or U6290 (N_6290,N_6225,N_5838);
xor U6291 (N_6291,N_5646,N_5752);
nand U6292 (N_6292,N_5152,N_3161);
and U6293 (N_6293,N_2860,N_1684);
or U6294 (N_6294,N_882,N_3447);
and U6295 (N_6295,N_3273,N_4242);
nor U6296 (N_6296,N_5610,N_475);
and U6297 (N_6297,N_3631,N_4723);
or U6298 (N_6298,N_1668,N_5037);
or U6299 (N_6299,N_4645,N_2987);
xor U6300 (N_6300,N_518,N_3919);
nor U6301 (N_6301,N_3505,N_4004);
or U6302 (N_6302,N_3704,N_2003);
and U6303 (N_6303,N_1573,N_404);
nand U6304 (N_6304,N_1367,N_3708);
xnor U6305 (N_6305,N_3026,N_2824);
nor U6306 (N_6306,N_6245,N_1679);
nor U6307 (N_6307,N_5638,N_1080);
and U6308 (N_6308,N_2052,N_2900);
nor U6309 (N_6309,N_4143,N_247);
nor U6310 (N_6310,N_344,N_46);
and U6311 (N_6311,N_1769,N_3935);
and U6312 (N_6312,N_431,N_2996);
xor U6313 (N_6313,N_5819,N_1146);
or U6314 (N_6314,N_4197,N_4009);
xnor U6315 (N_6315,N_5942,N_1175);
and U6316 (N_6316,N_2477,N_2901);
nand U6317 (N_6317,N_5674,N_5737);
nor U6318 (N_6318,N_2330,N_4283);
or U6319 (N_6319,N_4737,N_3471);
and U6320 (N_6320,N_1232,N_760);
and U6321 (N_6321,N_97,N_4256);
nand U6322 (N_6322,N_3050,N_5281);
or U6323 (N_6323,N_164,N_1115);
or U6324 (N_6324,N_2663,N_3084);
xor U6325 (N_6325,N_723,N_2490);
and U6326 (N_6326,N_1079,N_4435);
and U6327 (N_6327,N_3769,N_3636);
nor U6328 (N_6328,N_1036,N_3430);
nand U6329 (N_6329,N_6107,N_3393);
nand U6330 (N_6330,N_3669,N_3309);
or U6331 (N_6331,N_5875,N_1754);
or U6332 (N_6332,N_2576,N_3588);
nand U6333 (N_6333,N_957,N_1337);
and U6334 (N_6334,N_2817,N_5228);
nor U6335 (N_6335,N_5366,N_3477);
or U6336 (N_6336,N_4603,N_4718);
xnor U6337 (N_6337,N_3850,N_5512);
nor U6338 (N_6338,N_1980,N_5770);
xnor U6339 (N_6339,N_3241,N_3403);
xnor U6340 (N_6340,N_3743,N_2256);
and U6341 (N_6341,N_1520,N_4495);
or U6342 (N_6342,N_1207,N_196);
nand U6343 (N_6343,N_3360,N_1582);
or U6344 (N_6344,N_2364,N_2592);
nand U6345 (N_6345,N_1843,N_6128);
nor U6346 (N_6346,N_5252,N_59);
and U6347 (N_6347,N_5578,N_11);
or U6348 (N_6348,N_2652,N_3328);
nand U6349 (N_6349,N_4301,N_1496);
xor U6350 (N_6350,N_3446,N_5891);
nand U6351 (N_6351,N_3791,N_325);
nor U6352 (N_6352,N_338,N_4949);
and U6353 (N_6353,N_2971,N_1841);
xnor U6354 (N_6354,N_1360,N_3325);
nand U6355 (N_6355,N_2724,N_2394);
and U6356 (N_6356,N_2367,N_489);
and U6357 (N_6357,N_1690,N_3845);
xor U6358 (N_6358,N_4416,N_3853);
xnor U6359 (N_6359,N_2227,N_724);
or U6360 (N_6360,N_342,N_2104);
nand U6361 (N_6361,N_6077,N_5695);
nor U6362 (N_6362,N_4280,N_5910);
or U6363 (N_6363,N_4679,N_5396);
and U6364 (N_6364,N_1701,N_3330);
and U6365 (N_6365,N_4801,N_5572);
nand U6366 (N_6366,N_5144,N_5977);
nor U6367 (N_6367,N_5703,N_457);
and U6368 (N_6368,N_741,N_6237);
nand U6369 (N_6369,N_2243,N_1749);
nand U6370 (N_6370,N_5211,N_429);
and U6371 (N_6371,N_3587,N_937);
nor U6372 (N_6372,N_1858,N_452);
nor U6373 (N_6373,N_4391,N_2435);
or U6374 (N_6374,N_5530,N_4664);
xnor U6375 (N_6375,N_5081,N_3336);
xnor U6376 (N_6376,N_689,N_4299);
xnor U6377 (N_6377,N_2211,N_5567);
or U6378 (N_6378,N_2492,N_662);
nand U6379 (N_6379,N_2896,N_5755);
nor U6380 (N_6380,N_966,N_4052);
or U6381 (N_6381,N_3198,N_4255);
xor U6382 (N_6382,N_5257,N_2048);
or U6383 (N_6383,N_4483,N_2591);
nand U6384 (N_6384,N_4397,N_2271);
nor U6385 (N_6385,N_3346,N_324);
and U6386 (N_6386,N_1104,N_2923);
and U6387 (N_6387,N_2069,N_3680);
nand U6388 (N_6388,N_954,N_1482);
or U6389 (N_6389,N_2905,N_3282);
xnor U6390 (N_6390,N_3856,N_5063);
nand U6391 (N_6391,N_3373,N_540);
nand U6392 (N_6392,N_2739,N_1896);
xnor U6393 (N_6393,N_4121,N_5794);
nor U6394 (N_6394,N_648,N_1258);
or U6395 (N_6395,N_3132,N_5908);
nor U6396 (N_6396,N_2059,N_5730);
and U6397 (N_6397,N_5289,N_5587);
and U6398 (N_6398,N_5851,N_5583);
nand U6399 (N_6399,N_4225,N_4479);
or U6400 (N_6400,N_6018,N_4431);
or U6401 (N_6401,N_1665,N_2347);
xnor U6402 (N_6402,N_5275,N_2745);
nor U6403 (N_6403,N_1043,N_6109);
and U6404 (N_6404,N_2254,N_4434);
nand U6405 (N_6405,N_165,N_542);
or U6406 (N_6406,N_2633,N_2056);
xnor U6407 (N_6407,N_2341,N_3469);
xnor U6408 (N_6408,N_2604,N_5715);
and U6409 (N_6409,N_2160,N_5874);
or U6410 (N_6410,N_3970,N_2185);
nor U6411 (N_6411,N_5436,N_515);
and U6412 (N_6412,N_4497,N_6006);
nand U6413 (N_6413,N_4675,N_3349);
and U6414 (N_6414,N_997,N_1645);
xor U6415 (N_6415,N_3484,N_4565);
or U6416 (N_6416,N_5057,N_1765);
xor U6417 (N_6417,N_6087,N_4567);
and U6418 (N_6418,N_1188,N_2297);
nor U6419 (N_6419,N_2176,N_4165);
and U6420 (N_6420,N_1265,N_1413);
nor U6421 (N_6421,N_6137,N_4928);
nor U6422 (N_6422,N_1866,N_361);
and U6423 (N_6423,N_5322,N_1762);
or U6424 (N_6424,N_2555,N_2007);
nand U6425 (N_6425,N_1148,N_5611);
nor U6426 (N_6426,N_6209,N_2875);
and U6427 (N_6427,N_5290,N_6075);
or U6428 (N_6428,N_1880,N_498);
nor U6429 (N_6429,N_2720,N_5336);
nor U6430 (N_6430,N_1103,N_888);
xnor U6431 (N_6431,N_5016,N_2661);
or U6432 (N_6432,N_2990,N_871);
nand U6433 (N_6433,N_855,N_1353);
and U6434 (N_6434,N_3285,N_788);
nor U6435 (N_6435,N_2070,N_5230);
and U6436 (N_6436,N_3147,N_637);
nor U6437 (N_6437,N_4788,N_1268);
nand U6438 (N_6438,N_2726,N_2289);
or U6439 (N_6439,N_4780,N_2643);
and U6440 (N_6440,N_500,N_5262);
and U6441 (N_6441,N_3535,N_624);
and U6442 (N_6442,N_2674,N_3585);
nor U6443 (N_6443,N_820,N_5189);
nor U6444 (N_6444,N_4760,N_1630);
or U6445 (N_6445,N_2866,N_446);
xor U6446 (N_6446,N_2650,N_4187);
or U6447 (N_6447,N_2463,N_677);
nand U6448 (N_6448,N_4507,N_4900);
nand U6449 (N_6449,N_4335,N_3733);
nor U6450 (N_6450,N_5599,N_4164);
and U6451 (N_6451,N_215,N_1391);
nor U6452 (N_6452,N_2879,N_3259);
nor U6453 (N_6453,N_4348,N_2340);
or U6454 (N_6454,N_5486,N_1488);
nand U6455 (N_6455,N_2457,N_3583);
nor U6456 (N_6456,N_4471,N_780);
xor U6457 (N_6457,N_2630,N_5991);
nor U6458 (N_6458,N_2665,N_5129);
nor U6459 (N_6459,N_3960,N_1910);
nor U6460 (N_6460,N_4712,N_5849);
and U6461 (N_6461,N_5269,N_4040);
xnor U6462 (N_6462,N_4827,N_4219);
and U6463 (N_6463,N_3852,N_4881);
nand U6464 (N_6464,N_811,N_5995);
nand U6465 (N_6465,N_894,N_5753);
xor U6466 (N_6466,N_228,N_2727);
and U6467 (N_6467,N_4292,N_237);
xor U6468 (N_6468,N_1972,N_1348);
xor U6469 (N_6469,N_1672,N_4761);
nor U6470 (N_6470,N_5601,N_1859);
nand U6471 (N_6471,N_561,N_2151);
xor U6472 (N_6472,N_3376,N_3838);
nor U6473 (N_6473,N_1689,N_2001);
nor U6474 (N_6474,N_3539,N_3977);
and U6475 (N_6475,N_3700,N_3732);
xnor U6476 (N_6476,N_978,N_3542);
or U6477 (N_6477,N_5238,N_1914);
xor U6478 (N_6478,N_698,N_5623);
nor U6479 (N_6479,N_4960,N_4743);
nand U6480 (N_6480,N_2257,N_2025);
or U6481 (N_6481,N_2608,N_4033);
or U6482 (N_6482,N_735,N_577);
nand U6483 (N_6483,N_5681,N_848);
xor U6484 (N_6484,N_5088,N_280);
and U6485 (N_6485,N_1817,N_413);
xnor U6486 (N_6486,N_987,N_5020);
xor U6487 (N_6487,N_2606,N_4919);
or U6488 (N_6488,N_4996,N_6021);
xor U6489 (N_6489,N_3964,N_1244);
or U6490 (N_6490,N_3288,N_3875);
or U6491 (N_6491,N_2778,N_2155);
or U6492 (N_6492,N_2770,N_3450);
nor U6493 (N_6493,N_1707,N_5390);
xor U6494 (N_6494,N_5319,N_4215);
and U6495 (N_6495,N_6080,N_4465);
xnor U6496 (N_6496,N_288,N_3605);
nor U6497 (N_6497,N_1428,N_200);
xor U6498 (N_6498,N_4226,N_589);
nand U6499 (N_6499,N_3379,N_2237);
nand U6500 (N_6500,N_1465,N_1463);
and U6501 (N_6501,N_2887,N_4105);
nand U6502 (N_6502,N_5589,N_4285);
and U6503 (N_6503,N_1849,N_1119);
or U6504 (N_6504,N_646,N_1751);
xor U6505 (N_6505,N_3002,N_1472);
or U6506 (N_6506,N_113,N_5045);
and U6507 (N_6507,N_299,N_2623);
nor U6508 (N_6508,N_982,N_4037);
or U6509 (N_6509,N_4769,N_2156);
or U6510 (N_6510,N_2404,N_4045);
nor U6511 (N_6511,N_1341,N_1906);
nand U6512 (N_6512,N_5018,N_1592);
nand U6513 (N_6513,N_2090,N_5179);
and U6514 (N_6514,N_3258,N_5856);
or U6515 (N_6515,N_319,N_4287);
or U6516 (N_6516,N_833,N_5952);
xor U6517 (N_6517,N_5376,N_4854);
or U6518 (N_6518,N_6144,N_1270);
nor U6519 (N_6519,N_536,N_3174);
xnor U6520 (N_6520,N_5377,N_1004);
nand U6521 (N_6521,N_4825,N_66);
or U6522 (N_6522,N_263,N_4363);
and U6523 (N_6523,N_2332,N_3406);
nand U6524 (N_6524,N_1539,N_347);
and U6525 (N_6525,N_303,N_4205);
and U6526 (N_6526,N_5516,N_3164);
nor U6527 (N_6527,N_4281,N_5294);
and U6528 (N_6528,N_1793,N_3885);
xor U6529 (N_6529,N_5007,N_3668);
and U6530 (N_6530,N_2962,N_4012);
nor U6531 (N_6531,N_3740,N_5245);
nor U6532 (N_6532,N_1189,N_3413);
or U6533 (N_6533,N_2468,N_3490);
nand U6534 (N_6534,N_5647,N_6180);
nand U6535 (N_6535,N_390,N_5676);
nor U6536 (N_6536,N_559,N_3486);
nor U6537 (N_6537,N_3959,N_4936);
or U6538 (N_6538,N_3480,N_5268);
and U6539 (N_6539,N_3180,N_2951);
nor U6540 (N_6540,N_4302,N_1087);
xnor U6541 (N_6541,N_4583,N_2159);
nand U6542 (N_6542,N_3257,N_316);
nor U6543 (N_6543,N_499,N_6055);
nor U6544 (N_6544,N_4811,N_2798);
xnor U6545 (N_6545,N_2101,N_6168);
xor U6546 (N_6546,N_1173,N_3881);
and U6547 (N_6547,N_1796,N_5375);
nor U6548 (N_6548,N_5073,N_2312);
nand U6549 (N_6549,N_5680,N_3685);
or U6550 (N_6550,N_5187,N_2983);
or U6551 (N_6551,N_4261,N_298);
and U6552 (N_6552,N_3054,N_2396);
nor U6553 (N_6553,N_4439,N_3621);
nor U6554 (N_6554,N_5405,N_5127);
or U6555 (N_6555,N_2789,N_331);
xor U6556 (N_6556,N_2936,N_2966);
and U6557 (N_6557,N_5943,N_1008);
or U6558 (N_6558,N_534,N_2558);
or U6559 (N_6559,N_3256,N_3411);
xnor U6560 (N_6560,N_1015,N_990);
xnor U6561 (N_6561,N_1800,N_5345);
nor U6562 (N_6562,N_3274,N_4901);
nor U6563 (N_6563,N_3628,N_5938);
and U6564 (N_6564,N_3606,N_1435);
or U6565 (N_6565,N_3291,N_3519);
or U6566 (N_6566,N_1343,N_3133);
nor U6567 (N_6567,N_4976,N_3389);
or U6568 (N_6568,N_5065,N_5070);
xor U6569 (N_6569,N_1143,N_893);
xor U6570 (N_6570,N_2042,N_1801);
xor U6571 (N_6571,N_4332,N_4819);
xnor U6572 (N_6572,N_3812,N_4359);
xnor U6573 (N_6573,N_6040,N_4724);
nand U6574 (N_6574,N_1228,N_2715);
and U6575 (N_6575,N_5220,N_5644);
or U6576 (N_6576,N_2189,N_4719);
xnor U6577 (N_6577,N_1351,N_67);
or U6578 (N_6578,N_3872,N_3032);
nand U6579 (N_6579,N_682,N_2384);
or U6580 (N_6580,N_753,N_4550);
or U6581 (N_6581,N_2190,N_5864);
xor U6582 (N_6582,N_2970,N_2475);
xor U6583 (N_6583,N_2497,N_985);
nand U6584 (N_6584,N_6085,N_4371);
nand U6585 (N_6585,N_2370,N_4166);
or U6586 (N_6586,N_488,N_1437);
nor U6587 (N_6587,N_934,N_4566);
nor U6588 (N_6588,N_5782,N_1006);
nand U6589 (N_6589,N_4328,N_4875);
and U6590 (N_6590,N_6113,N_4845);
nand U6591 (N_6591,N_759,N_607);
nor U6592 (N_6592,N_1187,N_3135);
nor U6593 (N_6593,N_366,N_1154);
or U6594 (N_6594,N_4584,N_76);
nor U6595 (N_6595,N_1168,N_227);
nand U6596 (N_6596,N_3208,N_3412);
xnor U6597 (N_6597,N_4392,N_5075);
and U6598 (N_6598,N_3949,N_40);
or U6599 (N_6599,N_3182,N_4171);
nand U6600 (N_6600,N_3238,N_2333);
and U6601 (N_6601,N_5287,N_2410);
or U6602 (N_6602,N_6223,N_557);
nor U6603 (N_6603,N_1240,N_2294);
or U6604 (N_6604,N_4677,N_3059);
nor U6605 (N_6605,N_2486,N_4094);
nand U6606 (N_6606,N_6131,N_808);
and U6607 (N_6607,N_5357,N_5098);
nand U6608 (N_6608,N_266,N_3110);
and U6609 (N_6609,N_4145,N_1490);
and U6610 (N_6610,N_4943,N_1020);
or U6611 (N_6611,N_1518,N_244);
nor U6612 (N_6612,N_4103,N_5824);
and U6613 (N_6613,N_3644,N_3571);
nand U6614 (N_6614,N_4864,N_2038);
nor U6615 (N_6615,N_1656,N_1741);
or U6616 (N_6616,N_2952,N_3496);
nand U6617 (N_6617,N_3515,N_504);
xor U6618 (N_6618,N_803,N_2219);
or U6619 (N_6619,N_1022,N_6112);
and U6620 (N_6620,N_5207,N_3522);
or U6621 (N_6621,N_5886,N_4568);
or U6622 (N_6622,N_4717,N_4699);
and U6623 (N_6623,N_573,N_1863);
xor U6624 (N_6624,N_672,N_6190);
and U6625 (N_6625,N_953,N_638);
or U6626 (N_6626,N_2822,N_3319);
and U6627 (N_6627,N_6039,N_455);
and U6628 (N_6628,N_4611,N_4730);
or U6629 (N_6629,N_5103,N_4373);
and U6630 (N_6630,N_2488,N_752);
xnor U6631 (N_6631,N_1547,N_4025);
xor U6632 (N_6632,N_2051,N_3814);
nor U6633 (N_6633,N_1394,N_626);
xnor U6634 (N_6634,N_5725,N_2316);
and U6635 (N_6635,N_962,N_5441);
nor U6636 (N_6636,N_442,N_179);
and U6637 (N_6637,N_6060,N_936);
nand U6638 (N_6638,N_3239,N_2019);
xor U6639 (N_6639,N_1132,N_5193);
or U6640 (N_6640,N_4781,N_3504);
nand U6641 (N_6641,N_3653,N_368);
xor U6642 (N_6642,N_553,N_558);
or U6643 (N_6643,N_6095,N_4569);
nor U6644 (N_6644,N_3658,N_2679);
nand U6645 (N_6645,N_5557,N_4074);
nand U6646 (N_6646,N_268,N_4366);
xnor U6647 (N_6647,N_1566,N_4108);
nor U6648 (N_6648,N_251,N_2262);
nand U6649 (N_6649,N_1452,N_991);
and U6650 (N_6650,N_1067,N_467);
and U6651 (N_6651,N_3765,N_4379);
xor U6652 (N_6652,N_458,N_2164);
and U6653 (N_6653,N_1504,N_3524);
nand U6654 (N_6654,N_4742,N_4920);
and U6655 (N_6655,N_1342,N_722);
or U6656 (N_6656,N_1159,N_2361);
xor U6657 (N_6657,N_2016,N_1678);
nand U6658 (N_6658,N_4310,N_2234);
and U6659 (N_6659,N_2355,N_1653);
xnor U6660 (N_6660,N_3162,N_3011);
xnor U6661 (N_6661,N_4690,N_3362);
nand U6662 (N_6662,N_868,N_2682);
nand U6663 (N_6663,N_1949,N_3705);
and U6664 (N_6664,N_3893,N_221);
or U6665 (N_6665,N_2422,N_3896);
nor U6666 (N_6666,N_6152,N_1813);
and U6667 (N_6667,N_2761,N_528);
xor U6668 (N_6668,N_897,N_809);
nand U6669 (N_6669,N_5959,N_5130);
and U6670 (N_6670,N_1836,N_2685);
xnor U6671 (N_6671,N_4003,N_5165);
nand U6672 (N_6672,N_1542,N_1449);
xnor U6673 (N_6673,N_1944,N_4015);
nand U6674 (N_6674,N_2676,N_5421);
or U6675 (N_6675,N_2554,N_3038);
and U6676 (N_6676,N_5139,N_618);
and U6677 (N_6677,N_754,N_3777);
nand U6678 (N_6678,N_1983,N_5641);
xor U6679 (N_6679,N_3399,N_1591);
xor U6680 (N_6680,N_4214,N_4071);
nor U6681 (N_6681,N_3029,N_4834);
nand U6682 (N_6682,N_804,N_2018);
or U6683 (N_6683,N_1283,N_2245);
and U6684 (N_6684,N_5663,N_1108);
or U6685 (N_6685,N_2429,N_590);
or U6686 (N_6686,N_4779,N_3499);
or U6687 (N_6687,N_5461,N_785);
nor U6688 (N_6688,N_4563,N_562);
and U6689 (N_6689,N_1646,N_1038);
nor U6690 (N_6690,N_3094,N_3865);
or U6691 (N_6691,N_1911,N_5206);
and U6692 (N_6692,N_4752,N_6238);
or U6693 (N_6693,N_906,N_2821);
nor U6694 (N_6694,N_400,N_4602);
and U6695 (N_6695,N_1512,N_965);
or U6696 (N_6696,N_4721,N_5499);
or U6697 (N_6697,N_4929,N_2915);
nor U6698 (N_6698,N_1195,N_4078);
nand U6699 (N_6699,N_478,N_4184);
and U6700 (N_6700,N_4453,N_245);
or U6701 (N_6701,N_2705,N_5600);
nor U6702 (N_6702,N_454,N_6027);
and U6703 (N_6703,N_3410,N_4026);
nor U6704 (N_6704,N_4802,N_3437);
and U6705 (N_6705,N_424,N_5126);
xnor U6706 (N_6706,N_58,N_1210);
nand U6707 (N_6707,N_4194,N_1985);
or U6708 (N_6708,N_3693,N_1965);
nand U6709 (N_6709,N_5263,N_5151);
and U6710 (N_6710,N_2636,N_2765);
and U6711 (N_6711,N_3989,N_2550);
nand U6712 (N_6712,N_2169,N_4237);
or U6713 (N_6713,N_5535,N_2310);
and U6714 (N_6714,N_1190,N_3574);
and U6715 (N_6715,N_925,N_4462);
or U6716 (N_6716,N_173,N_710);
or U6717 (N_6717,N_199,N_2265);
nand U6718 (N_6718,N_2858,N_781);
nand U6719 (N_6719,N_2178,N_2470);
nand U6720 (N_6720,N_3092,N_5540);
nand U6721 (N_6721,N_5112,N_6160);
nor U6722 (N_6722,N_486,N_2984);
or U6723 (N_6723,N_5613,N_5010);
nor U6724 (N_6724,N_3409,N_6138);
nor U6725 (N_6725,N_3622,N_3564);
nor U6726 (N_6726,N_1315,N_4652);
nand U6727 (N_6727,N_2081,N_1651);
and U6728 (N_6728,N_667,N_2327);
and U6729 (N_6729,N_2907,N_5705);
nand U6730 (N_6730,N_2419,N_4433);
or U6731 (N_6731,N_2939,N_5720);
xnor U6732 (N_6732,N_4520,N_2482);
and U6733 (N_6733,N_3698,N_5391);
or U6734 (N_6734,N_3965,N_2105);
xnor U6735 (N_6735,N_4701,N_4182);
nand U6736 (N_6736,N_693,N_72);
or U6737 (N_6737,N_4981,N_1018);
and U6738 (N_6738,N_5538,N_2450);
and U6739 (N_6739,N_1112,N_4461);
and U6740 (N_6740,N_4179,N_2578);
xor U6741 (N_6741,N_845,N_2233);
and U6742 (N_6742,N_233,N_80);
or U6743 (N_6743,N_4297,N_1101);
nand U6744 (N_6744,N_4036,N_4740);
xor U6745 (N_6745,N_3516,N_4440);
or U6746 (N_6746,N_703,N_5763);
or U6747 (N_6747,N_5315,N_9);
or U6748 (N_6748,N_502,N_160);
and U6749 (N_6749,N_2718,N_4658);
nor U6750 (N_6750,N_1047,N_2218);
xnor U6751 (N_6751,N_4749,N_3108);
xnor U6752 (N_6752,N_744,N_2165);
xor U6753 (N_6753,N_4432,N_4774);
nand U6754 (N_6754,N_1634,N_5547);
nand U6755 (N_6755,N_1323,N_6167);
and U6756 (N_6756,N_2496,N_2639);
xnor U6757 (N_6757,N_5409,N_5698);
xor U6758 (N_6758,N_3159,N_3711);
xnor U6759 (N_6759,N_4269,N_1788);
nor U6760 (N_6760,N_2957,N_202);
and U6761 (N_6761,N_4449,N_1588);
nand U6762 (N_6762,N_2417,N_3003);
nor U6763 (N_6763,N_2182,N_2153);
xor U6764 (N_6764,N_908,N_2342);
nand U6765 (N_6765,N_278,N_3312);
nor U6766 (N_6766,N_612,N_1460);
and U6767 (N_6767,N_4755,N_4122);
nor U6768 (N_6768,N_3737,N_3276);
nor U6769 (N_6769,N_4174,N_4931);
or U6770 (N_6770,N_5041,N_3136);
xor U6771 (N_6771,N_4748,N_5356);
xnor U6772 (N_6772,N_1155,N_102);
or U6773 (N_6773,N_5687,N_3457);
and U6774 (N_6774,N_6036,N_3581);
xor U6775 (N_6775,N_2110,N_1297);
nand U6776 (N_6776,N_261,N_3314);
nor U6777 (N_6777,N_4238,N_4357);
and U6778 (N_6778,N_5802,N_4523);
nor U6779 (N_6779,N_5327,N_823);
xor U6780 (N_6780,N_547,N_3167);
xnor U6781 (N_6781,N_691,N_5645);
or U6782 (N_6782,N_5004,N_5579);
and U6783 (N_6783,N_1727,N_1537);
and U6784 (N_6784,N_2942,N_2637);
nand U6785 (N_6785,N_6207,N_2434);
nand U6786 (N_6786,N_1110,N_5899);
and U6787 (N_6787,N_1277,N_3886);
nand U6788 (N_6788,N_3530,N_4538);
xor U6789 (N_6789,N_4980,N_1638);
and U6790 (N_6790,N_3520,N_1164);
nor U6791 (N_6791,N_50,N_5086);
or U6792 (N_6792,N_1321,N_4381);
nor U6793 (N_6793,N_4131,N_2712);
nor U6794 (N_6794,N_4700,N_3316);
nor U6795 (N_6795,N_595,N_3646);
xor U6796 (N_6796,N_5531,N_212);
or U6797 (N_6797,N_1485,N_3400);
or U6798 (N_6798,N_5798,N_5491);
and U6799 (N_6799,N_5799,N_5905);
nand U6800 (N_6800,N_2658,N_787);
nand U6801 (N_6801,N_792,N_4532);
nor U6802 (N_6802,N_1469,N_4072);
or U6803 (N_6803,N_5458,N_1898);
nor U6804 (N_6804,N_3560,N_2882);
or U6805 (N_6805,N_1248,N_620);
xor U6806 (N_6806,N_5083,N_226);
nor U6807 (N_6807,N_4727,N_2744);
xnor U6808 (N_6808,N_3981,N_1682);
and U6809 (N_6809,N_422,N_4758);
nand U6810 (N_6810,N_5648,N_354);
or U6811 (N_6811,N_5015,N_4333);
nand U6812 (N_6812,N_1712,N_1920);
and U6813 (N_6813,N_4263,N_2740);
nor U6814 (N_6814,N_5387,N_3586);
xnor U6815 (N_6815,N_5332,N_4407);
or U6816 (N_6816,N_1586,N_5113);
or U6817 (N_6817,N_4419,N_3684);
xnor U6818 (N_6818,N_1430,N_6162);
or U6819 (N_6819,N_2388,N_5740);
xor U6820 (N_6820,N_3892,N_3112);
nand U6821 (N_6821,N_6046,N_3442);
or U6822 (N_6822,N_1293,N_926);
or U6823 (N_6823,N_4726,N_5964);
xnor U6824 (N_6824,N_5378,N_108);
xor U6825 (N_6825,N_214,N_1538);
and U6826 (N_6826,N_4653,N_3828);
and U6827 (N_6827,N_4189,N_4766);
nor U6828 (N_6828,N_1919,N_5198);
and U6829 (N_6829,N_2673,N_2741);
and U6830 (N_6830,N_3408,N_1025);
xor U6831 (N_6831,N_5622,N_4672);
and U6832 (N_6832,N_2023,N_2024);
or U6833 (N_6833,N_5359,N_5397);
nor U6834 (N_6834,N_5467,N_706);
xor U6835 (N_6835,N_4210,N_2572);
nand U6836 (N_6836,N_4589,N_891);
or U6837 (N_6837,N_3934,N_5506);
xnor U6838 (N_6838,N_3597,N_2632);
nand U6839 (N_6839,N_6206,N_6189);
and U6840 (N_6840,N_4659,N_5392);
xor U6841 (N_6841,N_5825,N_3141);
or U6842 (N_6842,N_1199,N_2738);
xor U6843 (N_6843,N_6059,N_5217);
or U6844 (N_6844,N_2614,N_2746);
xor U6845 (N_6845,N_5679,N_1064);
or U6846 (N_6846,N_4358,N_1434);
and U6847 (N_6847,N_2174,N_1137);
nand U6848 (N_6848,N_2964,N_5906);
xor U6849 (N_6849,N_3,N_4632);
nand U6850 (N_6850,N_3537,N_117);
xor U6851 (N_6851,N_3844,N_5003);
or U6852 (N_6852,N_5312,N_5367);
xor U6853 (N_6853,N_3811,N_1959);
nand U6854 (N_6854,N_3331,N_1737);
nand U6855 (N_6855,N_4591,N_5526);
or U6856 (N_6856,N_1288,N_1743);
nand U6857 (N_6857,N_4202,N_3230);
or U6858 (N_6858,N_4494,N_5051);
and U6859 (N_6859,N_1694,N_1017);
xnor U6860 (N_6860,N_523,N_1026);
nand U6861 (N_6861,N_5903,N_2390);
xor U6862 (N_6862,N_3523,N_3582);
nand U6863 (N_6863,N_4153,N_5347);
or U6864 (N_6864,N_4409,N_1226);
xor U6865 (N_6865,N_3649,N_2747);
nand U6866 (N_6866,N_2945,N_1696);
nand U6867 (N_6867,N_1074,N_757);
or U6868 (N_6868,N_5946,N_3183);
xnor U6869 (N_6869,N_4062,N_4579);
and U6870 (N_6870,N_1541,N_3272);
xnor U6871 (N_6871,N_5892,N_2114);
or U6872 (N_6872,N_3296,N_2456);
nor U6873 (N_6873,N_5767,N_4091);
and U6874 (N_6874,N_983,N_406);
and U6875 (N_6875,N_1388,N_3633);
or U6876 (N_6876,N_4270,N_2756);
xor U6877 (N_6877,N_5597,N_4676);
nor U6878 (N_6878,N_625,N_6165);
or U6879 (N_6879,N_3203,N_1354);
or U6880 (N_6880,N_1814,N_4065);
and U6881 (N_6881,N_4955,N_5097);
and U6882 (N_6882,N_4654,N_2510);
xor U6883 (N_6883,N_3361,N_5880);
and U6884 (N_6884,N_2138,N_5829);
or U6885 (N_6885,N_841,N_569);
and U6886 (N_6886,N_5940,N_2842);
xor U6887 (N_6887,N_5895,N_4200);
and U6888 (N_6888,N_1346,N_6171);
xnor U6889 (N_6889,N_5299,N_3154);
nor U6890 (N_6890,N_1185,N_2696);
or U6891 (N_6891,N_3172,N_1365);
nand U6892 (N_6892,N_913,N_3359);
or U6893 (N_6893,N_2060,N_2683);
and U6894 (N_6894,N_5867,N_4954);
and U6895 (N_6895,N_6247,N_2357);
xnor U6896 (N_6896,N_3613,N_1414);
and U6897 (N_6897,N_1279,N_3641);
nand U6898 (N_6898,N_621,N_3584);
nor U6899 (N_6899,N_1997,N_2757);
xnor U6900 (N_6900,N_3380,N_3315);
nand U6901 (N_6901,N_635,N_4794);
nor U6902 (N_6902,N_3173,N_5434);
or U6903 (N_6903,N_5412,N_5954);
nand U6904 (N_6904,N_2574,N_3169);
nand U6905 (N_6905,N_4463,N_5244);
and U6906 (N_6906,N_448,N_623);
nor U6907 (N_6907,N_863,N_4141);
or U6908 (N_6908,N_4486,N_5210);
nand U6909 (N_6909,N_1100,N_3255);
nor U6910 (N_6910,N_2045,N_1357);
or U6911 (N_6911,N_2517,N_6248);
or U6912 (N_6912,N_5806,N_5712);
and U6913 (N_6913,N_1613,N_4878);
xor U6914 (N_6914,N_3235,N_4290);
xnor U6915 (N_6915,N_3659,N_532);
or U6916 (N_6916,N_2803,N_1984);
nand U6917 (N_6917,N_4046,N_5326);
and U6918 (N_6918,N_2932,N_4629);
and U6919 (N_6919,N_1954,N_1402);
and U6920 (N_6920,N_2445,N_1931);
nand U6921 (N_6921,N_654,N_2489);
or U6922 (N_6922,N_5935,N_5044);
xor U6923 (N_6923,N_3106,N_3047);
and U6924 (N_6924,N_2992,N_1075);
nor U6925 (N_6925,N_5427,N_5748);
xor U6926 (N_6926,N_712,N_2818);
or U6927 (N_6927,N_2401,N_6020);
xnor U6928 (N_6928,N_2826,N_1016);
nand U6929 (N_6929,N_4161,N_3035);
xnor U6930 (N_6930,N_3416,N_4889);
xor U6931 (N_6931,N_3297,N_5076);
nor U6932 (N_6932,N_3064,N_3248);
xnor U6933 (N_6933,N_416,N_3688);
and U6934 (N_6934,N_377,N_5335);
and U6935 (N_6935,N_5371,N_2666);
and U6936 (N_6936,N_1392,N_1680);
or U6937 (N_6937,N_914,N_203);
nor U6938 (N_6938,N_996,N_4711);
xnor U6939 (N_6939,N_4627,N_2505);
nand U6940 (N_6940,N_1239,N_551);
xnor U6941 (N_6941,N_2197,N_4396);
or U6942 (N_6942,N_3647,N_2345);
nand U6943 (N_6943,N_875,N_4925);
nand U6944 (N_6944,N_2794,N_2043);
and U6945 (N_6945,N_4908,N_1318);
and U6946 (N_6946,N_951,N_5493);
nand U6947 (N_6947,N_3417,N_6084);
xor U6948 (N_6948,N_5194,N_2702);
xor U6949 (N_6949,N_4320,N_4100);
nor U6950 (N_6950,N_4912,N_1744);
nand U6951 (N_6951,N_75,N_501);
xor U6952 (N_6952,N_2118,N_191);
xor U6953 (N_6953,N_1407,N_5537);
or U6954 (N_6954,N_5562,N_6010);
and U6955 (N_6955,N_3513,N_217);
nand U6956 (N_6956,N_28,N_1879);
xnor U6957 (N_6957,N_1269,N_5285);
nor U6958 (N_6958,N_282,N_3694);
xnor U6959 (N_6959,N_5352,N_2473);
xnor U6960 (N_6960,N_4932,N_1060);
xor U6961 (N_6961,N_6210,N_2758);
and U6962 (N_6962,N_4420,N_47);
and U6963 (N_6963,N_1675,N_3240);
nor U6964 (N_6964,N_2725,N_5809);
and U6965 (N_6965,N_633,N_1420);
nor U6966 (N_6966,N_4886,N_4369);
and U6967 (N_6967,N_1118,N_4312);
xnor U6968 (N_6968,N_3137,N_1894);
and U6969 (N_6969,N_3292,N_2180);
nand U6970 (N_6970,N_3797,N_5455);
xor U6971 (N_6971,N_4666,N_3264);
or U6972 (N_6972,N_4725,N_5576);
xnor U6973 (N_6973,N_4883,N_1167);
or U6974 (N_6974,N_4832,N_5999);
nor U6975 (N_6975,N_5523,N_1885);
or U6976 (N_6976,N_3170,N_5149);
or U6977 (N_6977,N_5068,N_2548);
or U6978 (N_6978,N_1505,N_5214);
or U6979 (N_6979,N_4185,N_1010);
and U6980 (N_6980,N_879,N_4830);
or U6981 (N_6981,N_4180,N_5544);
nor U6982 (N_6982,N_4293,N_4810);
nand U6983 (N_6983,N_4775,N_5963);
or U6984 (N_6984,N_5990,N_4414);
nor U6985 (N_6985,N_5212,N_3057);
or U6986 (N_6986,N_1728,N_4298);
nand U6987 (N_6987,N_786,N_3916);
and U6988 (N_6988,N_5640,N_5408);
nand U6989 (N_6989,N_601,N_1963);
or U6990 (N_6990,N_5620,N_1850);
or U6991 (N_6991,N_1372,N_2167);
or U6992 (N_6992,N_928,N_4317);
and U6993 (N_6993,N_1907,N_4646);
and U6994 (N_6994,N_3962,N_3690);
or U6995 (N_6995,N_393,N_4600);
xor U6996 (N_6996,N_5559,N_18);
nor U6997 (N_6997,N_1317,N_1238);
xor U6998 (N_6998,N_3563,N_4456);
or U6999 (N_6999,N_529,N_1909);
or U7000 (N_7000,N_3905,N_60);
nand U7001 (N_7001,N_371,N_1877);
and U7002 (N_7002,N_873,N_3358);
nor U7003 (N_7003,N_1853,N_1549);
nand U7004 (N_7004,N_5163,N_2545);
or U7005 (N_7005,N_5060,N_2328);
xnor U7006 (N_7006,N_3150,N_4147);
nand U7007 (N_7007,N_3595,N_3983);
nand U7008 (N_7008,N_4064,N_6233);
nor U7009 (N_7009,N_1489,N_5700);
xor U7010 (N_7010,N_5815,N_3067);
nor U7011 (N_7011,N_5012,N_2759);
and U7012 (N_7012,N_5868,N_2807);
nor U7013 (N_7013,N_3901,N_3924);
xnor U7014 (N_7014,N_5568,N_5604);
nand U7015 (N_7015,N_4436,N_5417);
and U7016 (N_7016,N_3419,N_977);
nor U7017 (N_7017,N_4809,N_3554);
xor U7018 (N_7018,N_1719,N_3576);
xnor U7019 (N_7019,N_2276,N_3018);
nand U7020 (N_7020,N_1641,N_4389);
or U7021 (N_7021,N_1385,N_1097);
and U7022 (N_7022,N_4814,N_1453);
nor U7023 (N_7023,N_334,N_2050);
or U7024 (N_7024,N_1056,N_4111);
and U7025 (N_7025,N_2930,N_5121);
or U7026 (N_7026,N_3381,N_1379);
nor U7027 (N_7027,N_2293,N_3929);
xnor U7028 (N_7028,N_3324,N_3500);
nor U7029 (N_7029,N_4501,N_1338);
nand U7030 (N_7030,N_3263,N_6019);
or U7031 (N_7031,N_974,N_5574);
nor U7032 (N_7032,N_6008,N_1923);
and U7033 (N_7033,N_1454,N_3821);
nand U7034 (N_7034,N_2238,N_4887);
xor U7035 (N_7035,N_84,N_4860);
and U7036 (N_7036,N_3903,N_3253);
xnor U7037 (N_7037,N_4316,N_2953);
xnor U7038 (N_7038,N_3096,N_4828);
xor U7039 (N_7039,N_3833,N_3761);
and U7040 (N_7040,N_5525,N_1802);
and U7041 (N_7041,N_2981,N_3770);
xor U7042 (N_7042,N_1364,N_945);
and U7043 (N_7043,N_1948,N_127);
or U7044 (N_7044,N_3472,N_4119);
nor U7045 (N_7045,N_4253,N_4597);
nor U7046 (N_7046,N_784,N_1726);
nor U7047 (N_7047,N_899,N_3113);
nor U7048 (N_7048,N_3143,N_3327);
nand U7049 (N_7049,N_5173,N_3579);
and U7050 (N_7050,N_2799,N_2671);
xnor U7051 (N_7051,N_6133,N_77);
xnor U7052 (N_7052,N_3069,N_5514);
nor U7053 (N_7053,N_4093,N_2844);
nor U7054 (N_7054,N_1039,N_1135);
or U7055 (N_7055,N_858,N_1932);
nor U7056 (N_7056,N_153,N_5912);
xnor U7057 (N_7057,N_3283,N_4913);
or U7058 (N_7058,N_5504,N_4481);
xor U7059 (N_7059,N_2598,N_4384);
and U7060 (N_7060,N_4786,N_4594);
xnor U7061 (N_7061,N_2041,N_3424);
nor U7062 (N_7062,N_4559,N_3701);
nand U7063 (N_7063,N_205,N_805);
nand U7064 (N_7064,N_4013,N_4362);
or U7065 (N_7065,N_1815,N_2177);
or U7066 (N_7066,N_2678,N_1217);
or U7067 (N_7067,N_5692,N_3549);
nand U7068 (N_7068,N_2378,N_645);
and U7069 (N_7069,N_3873,N_2564);
or U7070 (N_7070,N_6153,N_4642);
nand U7071 (N_7071,N_4762,N_849);
nor U7072 (N_7072,N_519,N_4115);
nand U7073 (N_7073,N_4916,N_6111);
nor U7074 (N_7074,N_89,N_1052);
nor U7075 (N_7075,N_4872,N_1349);
and U7076 (N_7076,N_653,N_2567);
and U7077 (N_7077,N_3603,N_1116);
and U7078 (N_7078,N_2212,N_3654);
nor U7079 (N_7079,N_4354,N_2699);
nor U7080 (N_7080,N_5154,N_3829);
and U7081 (N_7081,N_328,N_2129);
xnor U7082 (N_7082,N_1298,N_3895);
nand U7083 (N_7083,N_6073,N_1519);
and U7084 (N_7084,N_385,N_3799);
xnor U7085 (N_7085,N_3443,N_1900);
and U7086 (N_7086,N_2693,N_3712);
or U7087 (N_7087,N_4476,N_3171);
nand U7088 (N_7088,N_2386,N_1623);
nand U7089 (N_7089,N_5080,N_3275);
or U7090 (N_7090,N_5612,N_2166);
nand U7091 (N_7091,N_238,N_1713);
or U7092 (N_7092,N_2222,N_2793);
and U7093 (N_7093,N_3270,N_2249);
nand U7094 (N_7094,N_4813,N_359);
and U7095 (N_7095,N_1499,N_602);
or U7096 (N_7096,N_889,N_505);
xor U7097 (N_7097,N_4641,N_1229);
xnor U7098 (N_7098,N_265,N_2498);
or U7099 (N_7099,N_1053,N_1427);
nand U7100 (N_7100,N_3807,N_2398);
or U7101 (N_7101,N_4423,N_1221);
and U7102 (N_7102,N_5719,N_719);
or U7103 (N_7103,N_993,N_4241);
or U7104 (N_7104,N_5479,N_2892);
nand U7105 (N_7105,N_388,N_1356);
xnor U7106 (N_7106,N_1249,N_5071);
nand U7107 (N_7107,N_2978,N_927);
or U7108 (N_7108,N_919,N_1943);
and U7109 (N_7109,N_3805,N_1380);
nor U7110 (N_7110,N_4343,N_4211);
nor U7111 (N_7111,N_295,N_1868);
or U7112 (N_7112,N_6092,N_3810);
xnor U7113 (N_7113,N_438,N_5743);
and U7114 (N_7114,N_4276,N_1576);
nand U7115 (N_7115,N_3078,N_1412);
nand U7116 (N_7116,N_5582,N_1241);
and U7117 (N_7117,N_2767,N_1165);
nor U7118 (N_7118,N_1181,N_1237);
xor U7119 (N_7119,N_2838,N_5756);
xnor U7120 (N_7120,N_615,N_2995);
or U7121 (N_7121,N_3280,N_5793);
xnor U7122 (N_7122,N_5333,N_3958);
and U7123 (N_7123,N_1470,N_3445);
and U7124 (N_7124,N_5072,N_3952);
xor U7125 (N_7125,N_5509,N_1410);
xnor U7126 (N_7126,N_4388,N_4738);
xor U7127 (N_7127,N_5474,N_2688);
nand U7128 (N_7128,N_4217,N_4443);
nand U7129 (N_7129,N_1131,N_4154);
nand U7130 (N_7130,N_2175,N_3105);
nand U7131 (N_7131,N_112,N_3825);
nor U7132 (N_7132,N_5662,N_2827);
nor U7133 (N_7133,N_4468,N_167);
nor U7134 (N_7134,N_1399,N_1747);
or U7135 (N_7135,N_1927,N_609);
xor U7136 (N_7136,N_3061,N_2815);
nand U7137 (N_7137,N_145,N_600);
nor U7138 (N_7138,N_1973,N_7);
and U7139 (N_7139,N_6240,N_6230);
and U7140 (N_7140,N_3005,N_4992);
and U7141 (N_7141,N_2600,N_2339);
nand U7142 (N_7142,N_4323,N_2231);
xnor U7143 (N_7143,N_5814,N_195);
xor U7144 (N_7144,N_1446,N_1462);
or U7145 (N_7145,N_2351,N_326);
nor U7146 (N_7146,N_5803,N_1621);
nor U7147 (N_7147,N_5303,N_943);
or U7148 (N_7148,N_5410,N_2569);
xnor U7149 (N_7149,N_5025,N_2267);
and U7150 (N_7150,N_564,N_3339);
nor U7151 (N_7151,N_1034,N_4206);
xnor U7152 (N_7152,N_6200,N_5900);
and U7153 (N_7153,N_3908,N_307);
nor U7154 (N_7154,N_5017,N_3772);
xor U7155 (N_7155,N_3087,N_3365);
and U7156 (N_7156,N_687,N_5032);
xor U7157 (N_7157,N_4286,N_4616);
and U7158 (N_7158,N_636,N_2976);
or U7159 (N_7159,N_2956,N_4059);
xor U7160 (N_7160,N_3223,N_1214);
nor U7161 (N_7161,N_3277,N_408);
xor U7162 (N_7162,N_538,N_3933);
or U7163 (N_7163,N_2768,N_6234);
and U7164 (N_7164,N_4516,N_4998);
or U7165 (N_7165,N_3391,N_4596);
and U7166 (N_7166,N_5881,N_5751);
nand U7167 (N_7167,N_1552,N_5757);
or U7168 (N_7168,N_1996,N_5816);
or U7169 (N_7169,N_1692,N_5496);
and U7170 (N_7170,N_920,N_5440);
nand U7171 (N_7171,N_1609,N_3823);
or U7172 (N_7172,N_4896,N_2399);
nand U7173 (N_7173,N_1637,N_5971);
or U7174 (N_7174,N_1153,N_3998);
or U7175 (N_7175,N_2791,N_2020);
nor U7176 (N_7176,N_5690,N_2621);
nor U7177 (N_7177,N_4689,N_2172);
xnor U7178 (N_7178,N_4356,N_2183);
and U7179 (N_7179,N_5833,N_2993);
xor U7180 (N_7180,N_4984,N_657);
nor U7181 (N_7181,N_2709,N_3991);
and U7182 (N_7182,N_64,N_4638);
nand U7183 (N_7183,N_3142,N_4714);
or U7184 (N_7184,N_3986,N_5628);
or U7185 (N_7185,N_4622,N_4570);
nor U7186 (N_7186,N_1502,N_3427);
nor U7187 (N_7187,N_4370,N_4682);
nor U7188 (N_7188,N_121,N_2743);
nand U7189 (N_7189,N_208,N_2440);
nand U7190 (N_7190,N_3681,N_778);
xnor U7191 (N_7191,N_4800,N_2337);
xor U7192 (N_7192,N_6194,N_6186);
nor U7193 (N_7193,N_1585,N_5177);
nor U7194 (N_7194,N_860,N_5984);
or U7195 (N_7195,N_6132,N_5841);
nand U7196 (N_7196,N_5921,N_2026);
xnor U7197 (N_7197,N_4163,N_133);
xor U7198 (N_7198,N_1174,N_989);
nand U7199 (N_7199,N_599,N_1059);
or U7200 (N_7200,N_679,N_3052);
xor U7201 (N_7201,N_2525,N_3779);
nor U7202 (N_7202,N_4049,N_3664);
xnor U7203 (N_7203,N_427,N_6239);
nor U7204 (N_7204,N_1917,N_1231);
or U7205 (N_7205,N_5236,N_3936);
and U7206 (N_7206,N_2524,N_4706);
and U7207 (N_7207,N_6001,N_2928);
nand U7208 (N_7208,N_5769,N_4741);
or U7209 (N_7209,N_3577,N_3997);
or U7210 (N_7210,N_4986,N_3076);
nor U7211 (N_7211,N_5054,N_1424);
nor U7212 (N_7212,N_5314,N_4368);
nor U7213 (N_7213,N_1055,N_2480);
nor U7214 (N_7214,N_1783,N_2346);
nor U7215 (N_7215,N_1976,N_3033);
or U7216 (N_7216,N_109,N_5666);
or U7217 (N_7217,N_5775,N_2418);
nor U7218 (N_7218,N_5524,N_747);
nand U7219 (N_7219,N_2369,N_175);
nor U7220 (N_7220,N_2128,N_1893);
or U7221 (N_7221,N_3548,N_3601);
and U7222 (N_7222,N_2692,N_1358);
nor U7223 (N_7223,N_1565,N_1742);
xnor U7224 (N_7224,N_1771,N_1686);
xor U7225 (N_7225,N_5339,N_1251);
nand U7226 (N_7226,N_4138,N_1378);
and U7227 (N_7227,N_1770,N_2668);
and U7228 (N_7228,N_110,N_2522);
or U7229 (N_7229,N_2622,N_4948);
nor U7230 (N_7230,N_775,N_3609);
nor U7231 (N_7231,N_3165,N_1501);
and U7232 (N_7232,N_2058,N_1534);
nor U7233 (N_7233,N_4192,N_2811);
nand U7234 (N_7234,N_1905,N_5800);
xor U7235 (N_7235,N_994,N_3689);
and U7236 (N_7236,N_697,N_5592);
and U7237 (N_7237,N_4577,N_5573);
nand U7238 (N_7238,N_3909,N_3666);
and U7239 (N_7239,N_4848,N_2202);
xor U7240 (N_7240,N_1642,N_3479);
nand U7241 (N_7241,N_5384,N_3074);
and U7242 (N_7242,N_5492,N_1001);
or U7243 (N_7243,N_3322,N_4958);
and U7244 (N_7244,N_5758,N_3979);
or U7245 (N_7245,N_4704,N_5286);
nor U7246 (N_7246,N_4782,N_1659);
xor U7247 (N_7247,N_1447,N_4457);
xnor U7248 (N_7248,N_1797,N_5528);
nor U7249 (N_7249,N_4678,N_887);
nand U7250 (N_7250,N_2210,N_5014);
xnor U7251 (N_7251,N_1497,N_3190);
and U7252 (N_7252,N_1425,N_3278);
nand U7253 (N_7253,N_6249,N_5955);
and U7254 (N_7254,N_2729,N_4867);
nand U7255 (N_7255,N_4096,N_5053);
xor U7256 (N_7256,N_4451,N_5160);
nor U7257 (N_7257,N_5801,N_737);
or U7258 (N_7258,N_2008,N_6216);
nor U7259 (N_7259,N_473,N_494);
and U7260 (N_7260,N_6053,N_2610);
xnor U7261 (N_7261,N_5697,N_3476);
or U7262 (N_7262,N_647,N_676);
nand U7263 (N_7263,N_2960,N_6246);
xor U7264 (N_7264,N_5200,N_104);
xnor U7265 (N_7265,N_2975,N_769);
nor U7266 (N_7266,N_132,N_918);
and U7267 (N_7267,N_5655,N_1445);
xnor U7268 (N_7268,N_6197,N_3247);
nand U7269 (N_7269,N_5428,N_1835);
nand U7270 (N_7270,N_3394,N_267);
nor U7271 (N_7271,N_2344,N_580);
nand U7272 (N_7272,N_2948,N_3900);
or U7273 (N_7273,N_5580,N_6062);
or U7274 (N_7274,N_5701,N_1309);
nand U7275 (N_7275,N_1822,N_3160);
nand U7276 (N_7276,N_352,N_1551);
nor U7277 (N_7277,N_5473,N_2471);
nand U7278 (N_7278,N_6235,N_3485);
nand U7279 (N_7279,N_5532,N_900);
or U7280 (N_7280,N_1577,N_3789);
or U7281 (N_7281,N_5796,N_5364);
nor U7282 (N_7282,N_4888,N_1172);
and U7283 (N_7283,N_896,N_5865);
nor U7284 (N_7284,N_2836,N_1250);
and U7285 (N_7285,N_4649,N_468);
and U7286 (N_7286,N_3225,N_2288);
nor U7287 (N_7287,N_1076,N_3451);
or U7288 (N_7288,N_4554,N_4467);
xor U7289 (N_7289,N_4252,N_3553);
or U7290 (N_7290,N_6214,N_818);
and U7291 (N_7291,N_4626,N_1395);
xnor U7292 (N_7292,N_2601,N_4874);
nor U7293 (N_7293,N_5049,N_2501);
or U7294 (N_7294,N_5256,N_1142);
nand U7295 (N_7295,N_1295,N_2072);
and U7296 (N_7296,N_180,N_2358);
nand U7297 (N_7297,N_3822,N_2982);
and U7298 (N_7298,N_2568,N_904);
and U7299 (N_7299,N_5430,N_1386);
xnor U7300 (N_7300,N_684,N_4835);
or U7301 (N_7301,N_4191,N_341);
and U7302 (N_7302,N_5399,N_4337);
nor U7303 (N_7303,N_6121,N_3874);
nor U7304 (N_7304,N_3337,N_1966);
nand U7305 (N_7305,N_4833,N_5422);
nand U7306 (N_7306,N_6066,N_738);
xor U7307 (N_7307,N_4515,N_1508);
or U7308 (N_7308,N_2259,N_5840);
and U7309 (N_7309,N_5342,N_4983);
xnor U7310 (N_7310,N_2359,N_1308);
nand U7311 (N_7311,N_43,N_294);
or U7312 (N_7312,N_4858,N_2061);
and U7313 (N_7313,N_4879,N_5626);
or U7314 (N_7314,N_700,N_5873);
nand U7315 (N_7315,N_2898,N_2837);
and U7316 (N_7316,N_4869,N_527);
or U7317 (N_7317,N_372,N_3529);
or U7318 (N_7318,N_5120,N_1282);
xnor U7319 (N_7319,N_3650,N_2651);
nor U7320 (N_7320,N_1090,N_4530);
nor U7321 (N_7321,N_1507,N_5291);
and U7322 (N_7322,N_641,N_5111);
and U7323 (N_7323,N_2521,N_979);
nor U7324 (N_7324,N_2904,N_3234);
and U7325 (N_7325,N_1882,N_3425);
nor U7326 (N_7326,N_3048,N_3065);
or U7327 (N_7327,N_2520,N_4926);
nand U7328 (N_7328,N_924,N_2494);
or U7329 (N_7329,N_2331,N_4921);
xnor U7330 (N_7330,N_1784,N_632);
or U7331 (N_7331,N_4904,N_3244);
or U7332 (N_7332,N_5148,N_4360);
nand U7333 (N_7333,N_608,N_4993);
or U7334 (N_7334,N_3607,N_1096);
xor U7335 (N_7335,N_5508,N_1533);
or U7336 (N_7336,N_5221,N_4985);
and U7337 (N_7337,N_4995,N_3773);
nor U7338 (N_7338,N_63,N_6057);
and U7339 (N_7339,N_5386,N_4662);
and U7340 (N_7340,N_3215,N_5176);
and U7341 (N_7341,N_2881,N_5092);
nor U7342 (N_7342,N_4181,N_6149);
nor U7343 (N_7343,N_1205,N_2449);
nor U7344 (N_7344,N_576,N_281);
and U7345 (N_7345,N_1939,N_1319);
or U7346 (N_7346,N_4266,N_1264);
xnor U7347 (N_7347,N_4613,N_720);
or U7348 (N_7348,N_4125,N_1555);
or U7349 (N_7349,N_1820,N_4445);
or U7350 (N_7350,N_5052,N_4365);
and U7351 (N_7351,N_1384,N_2295);
and U7352 (N_7352,N_1345,N_6005);
nor U7353 (N_7353,N_736,N_800);
and U7354 (N_7354,N_3384,N_6094);
xnor U7355 (N_7355,N_1544,N_946);
nand U7356 (N_7356,N_3332,N_322);
or U7357 (N_7357,N_4315,N_1774);
and U7358 (N_7358,N_3941,N_2057);
nor U7359 (N_7359,N_2989,N_4385);
and U7360 (N_7360,N_4464,N_980);
and U7361 (N_7361,N_776,N_2777);
and U7362 (N_7362,N_3843,N_4376);
xnor U7363 (N_7363,N_6007,N_4051);
nor U7364 (N_7364,N_3869,N_4446);
nor U7365 (N_7365,N_4850,N_1629);
nand U7366 (N_7366,N_2299,N_3206);
nor U7367 (N_7367,N_4086,N_1677);
or U7368 (N_7368,N_1990,N_3098);
nor U7369 (N_7369,N_119,N_854);
or U7370 (N_7370,N_3677,N_103);
nor U7371 (N_7371,N_4254,N_5330);
nand U7372 (N_7372,N_4159,N_3194);
xor U7373 (N_7373,N_3610,N_2619);
nor U7374 (N_7374,N_4491,N_2861);
xnor U7375 (N_7375,N_4444,N_1865);
and U7376 (N_7376,N_853,N_435);
or U7377 (N_7377,N_124,N_1511);
and U7378 (N_7378,N_323,N_1851);
or U7379 (N_7379,N_4917,N_4553);
or U7380 (N_7380,N_1366,N_95);
nor U7381 (N_7381,N_3082,N_5893);
xor U7382 (N_7382,N_4807,N_4475);
or U7383 (N_7383,N_3036,N_2430);
or U7384 (N_7384,N_4868,N_3102);
nand U7385 (N_7385,N_3269,N_2810);
nor U7386 (N_7386,N_1554,N_5146);
nor U7387 (N_7387,N_3009,N_4288);
xor U7388 (N_7388,N_3062,N_5229);
nand U7389 (N_7389,N_5066,N_4144);
xnor U7390 (N_7390,N_1652,N_895);
xnor U7391 (N_7391,N_3488,N_4245);
and U7392 (N_7392,N_552,N_2063);
and U7393 (N_7393,N_3993,N_2979);
nand U7394 (N_7394,N_3458,N_5821);
or U7395 (N_7395,N_2535,N_767);
nand U7396 (N_7396,N_2142,N_4408);
or U7397 (N_7397,N_1062,N_4282);
or U7398 (N_7398,N_4527,N_5624);
nor U7399 (N_7399,N_1699,N_4599);
nor U7400 (N_7400,N_5331,N_4710);
nand U7401 (N_7401,N_1091,N_740);
or U7402 (N_7402,N_2782,N_4812);
nor U7403 (N_7403,N_2988,N_1922);
nand U7404 (N_7404,N_409,N_5745);
xor U7405 (N_7405,N_1752,N_3184);
or U7406 (N_7406,N_2268,N_4895);
nor U7407 (N_7407,N_5546,N_5180);
nor U7408 (N_7408,N_5321,N_5554);
nand U7409 (N_7409,N_2163,N_5246);
nor U7410 (N_7410,N_4247,N_6228);
and U7411 (N_7411,N_2469,N_1421);
nor U7412 (N_7412,N_289,N_2073);
nor U7413 (N_7413,N_6089,N_5914);
and U7414 (N_7414,N_192,N_1969);
nand U7415 (N_7415,N_6048,N_2068);
nor U7416 (N_7416,N_2891,N_3083);
or U7417 (N_7417,N_2870,N_147);
or U7418 (N_7418,N_5453,N_3857);
or U7419 (N_7419,N_5099,N_1583);
nand U7420 (N_7420,N_1806,N_1332);
and U7421 (N_7421,N_5569,N_5298);
and U7422 (N_7422,N_4042,N_1440);
nand U7423 (N_7423,N_714,N_5739);
nor U7424 (N_7424,N_5002,N_2570);
and U7425 (N_7425,N_5485,N_4221);
nor U7426 (N_7426,N_4961,N_1160);
or U7427 (N_7427,N_1693,N_630);
nor U7428 (N_7428,N_5928,N_476);
or U7429 (N_7429,N_4127,N_2857);
nor U7430 (N_7430,N_1683,N_4628);
xnor U7431 (N_7431,N_2149,N_3343);
nor U7432 (N_7432,N_3943,N_1045);
xnor U7433 (N_7433,N_5095,N_3846);
xnor U7434 (N_7434,N_1991,N_3766);
nor U7435 (N_7435,N_5742,N_5247);
and U7436 (N_7436,N_4089,N_1604);
nand U7437 (N_7437,N_670,N_5191);
or U7438 (N_7438,N_249,N_1522);
and U7439 (N_7439,N_1595,N_5178);
nand U7440 (N_7440,N_3672,N_1149);
nand U7441 (N_7441,N_3086,N_586);
nand U7442 (N_7442,N_19,N_5264);
xnor U7443 (N_7443,N_2537,N_2319);
xnor U7444 (N_7444,N_4692,N_2616);
or U7445 (N_7445,N_3912,N_3073);
nand U7446 (N_7446,N_2563,N_2684);
nor U7447 (N_7447,N_3994,N_1999);
nor U7448 (N_7448,N_4558,N_6241);
and U7449 (N_7449,N_2620,N_262);
and U7450 (N_7450,N_1614,N_1140);
or U7451 (N_7451,N_4142,N_4784);
nor U7452 (N_7452,N_1952,N_4448);
nand U7453 (N_7453,N_1464,N_4756);
nor U7454 (N_7454,N_2380,N_3898);
or U7455 (N_7455,N_5871,N_4305);
nand U7456 (N_7456,N_5278,N_3969);
nand U7457 (N_7457,N_3861,N_627);
nor U7458 (N_7458,N_5358,N_2596);
xor U7459 (N_7459,N_4101,N_2270);
nand U7460 (N_7460,N_4853,N_5381);
and U7461 (N_7461,N_2033,N_4032);
or U7462 (N_7462,N_6213,N_1029);
xor U7463 (N_7463,N_5866,N_4671);
or U7464 (N_7464,N_1776,N_2933);
and U7465 (N_7465,N_4106,N_5433);
or U7466 (N_7466,N_5031,N_956);
xor U7467 (N_7467,N_434,N_1657);
and U7468 (N_7468,N_4823,N_2377);
xor U7469 (N_7469,N_115,N_358);
or U7470 (N_7470,N_2922,N_5653);
nand U7471 (N_7471,N_57,N_5021);
or U7472 (N_7472,N_4633,N_128);
and U7473 (N_7473,N_2329,N_4557);
or U7474 (N_7474,N_4284,N_3008);
xnor U7475 (N_7475,N_1736,N_32);
nand U7476 (N_7476,N_3975,N_1475);
nor U7477 (N_7477,N_2292,N_5028);
nor U7478 (N_7478,N_3569,N_5608);
xor U7479 (N_7479,N_1120,N_4020);
nand U7480 (N_7480,N_5619,N_2804);
or U7481 (N_7481,N_3913,N_157);
nor U7482 (N_7482,N_1122,N_2593);
nand U7483 (N_7483,N_6201,N_4364);
xnor U7484 (N_7484,N_2354,N_2352);
xnor U7485 (N_7485,N_2760,N_4137);
or U7486 (N_7486,N_4971,N_4933);
nand U7487 (N_7487,N_4412,N_2751);
xor U7488 (N_7488,N_3511,N_3387);
nand U7489 (N_7489,N_1704,N_2066);
nor U7490 (N_7490,N_2366,N_733);
xor U7491 (N_7491,N_5418,N_5169);
or U7492 (N_7492,N_2491,N_5729);
xor U7493 (N_7493,N_3946,N_1397);
nor U7494 (N_7494,N_3927,N_4797);
or U7495 (N_7495,N_3207,N_3079);
or U7496 (N_7496,N_3557,N_395);
xor U7497 (N_7497,N_4585,N_6208);
nor U7498 (N_7498,N_1459,N_4209);
or U7499 (N_7499,N_1738,N_1785);
and U7500 (N_7500,N_4489,N_2835);
xnor U7501 (N_7501,N_220,N_1109);
and U7502 (N_7502,N_1746,N_998);
or U7503 (N_7503,N_5301,N_6220);
and U7504 (N_7504,N_1368,N_750);
nand U7505 (N_7505,N_3510,N_190);
nor U7506 (N_7506,N_5362,N_2689);
xnor U7507 (N_7507,N_1916,N_910);
and U7508 (N_7508,N_5534,N_4129);
or U7509 (N_7509,N_4190,N_6173);
or U7510 (N_7510,N_4213,N_661);
or U7511 (N_7511,N_6159,N_4271);
or U7512 (N_7512,N_2314,N_5374);
xor U7513 (N_7513,N_3075,N_696);
nand U7514 (N_7514,N_2283,N_3103);
nor U7515 (N_7515,N_1724,N_678);
nor U7516 (N_7516,N_5484,N_3662);
or U7517 (N_7517,N_3368,N_1758);
or U7518 (N_7518,N_3817,N_1107);
xor U7519 (N_7519,N_2124,N_4499);
nand U7520 (N_7520,N_1698,N_5760);
nor U7521 (N_7521,N_2203,N_4273);
and U7522 (N_7522,N_3870,N_283);
nor U7523 (N_7523,N_3572,N_12);
nand U7524 (N_7524,N_4946,N_5683);
nor U7525 (N_7525,N_1271,N_1183);
or U7526 (N_7526,N_3858,N_511);
and U7527 (N_7527,N_4959,N_2755);
or U7528 (N_7528,N_2136,N_1967);
nand U7529 (N_7529,N_1325,N_3156);
nand U7530 (N_7530,N_1327,N_3468);
and U7531 (N_7531,N_5685,N_3625);
nand U7532 (N_7532,N_3623,N_1389);
and U7533 (N_7533,N_2941,N_236);
nand U7534 (N_7534,N_239,N_2774);
xor U7535 (N_7535,N_2748,N_1951);
nand U7536 (N_7536,N_2053,N_1186);
nor U7537 (N_7537,N_6122,N_329);
and U7538 (N_7538,N_391,N_2780);
nand U7539 (N_7539,N_1562,N_5337);
and U7540 (N_7540,N_1262,N_2371);
nor U7541 (N_7541,N_1287,N_5961);
nand U7542 (N_7542,N_4855,N_216);
and U7543 (N_7543,N_828,N_2044);
nor U7544 (N_7544,N_1902,N_3474);
or U7545 (N_7545,N_4452,N_2205);
nor U7546 (N_7546,N_3864,N_0);
or U7547 (N_7547,N_444,N_5009);
or U7548 (N_7548,N_2431,N_2506);
nand U7549 (N_7549,N_1942,N_2258);
nor U7550 (N_7550,N_2423,N_4927);
nor U7551 (N_7551,N_2762,N_1429);
and U7552 (N_7552,N_2495,N_3847);
xnor U7553 (N_7553,N_3453,N_24);
or U7554 (N_7554,N_484,N_82);
and U7555 (N_7555,N_727,N_5402);
and U7556 (N_7556,N_6100,N_4640);
xnor U7557 (N_7557,N_2544,N_1021);
nand U7558 (N_7558,N_2036,N_4382);
xor U7559 (N_7559,N_1935,N_3715);
or U7560 (N_7560,N_1245,N_2634);
or U7561 (N_7561,N_2402,N_5026);
nand U7562 (N_7562,N_5087,N_5706);
or U7563 (N_7563,N_3095,N_81);
xor U7564 (N_7564,N_335,N_2707);
nand U7565 (N_7565,N_6217,N_4513);
nand U7566 (N_7566,N_2571,N_2139);
nor U7567 (N_7567,N_3140,N_5419);
or U7568 (N_7568,N_2560,N_3626);
nand U7569 (N_7569,N_1032,N_4387);
nand U7570 (N_7570,N_1432,N_2853);
nor U7571 (N_7571,N_3444,N_2706);
and U7572 (N_7572,N_5202,N_5788);
and U7573 (N_7573,N_1703,N_907);
nand U7574 (N_7574,N_3842,N_898);
and U7575 (N_7575,N_1509,N_1831);
nand U7576 (N_7576,N_151,N_6093);
or U7577 (N_7577,N_2426,N_4314);
and U7578 (N_7578,N_376,N_5471);
or U7579 (N_7579,N_1223,N_2750);
nor U7580 (N_7580,N_4024,N_4634);
xnor U7581 (N_7581,N_3784,N_568);
or U7582 (N_7582,N_4744,N_680);
nand U7583 (N_7583,N_1124,N_3126);
or U7584 (N_7584,N_1669,N_2890);
nand U7585 (N_7585,N_5772,N_1768);
and U7586 (N_7586,N_2144,N_5388);
nand U7587 (N_7587,N_480,N_3985);
and U7588 (N_7588,N_5167,N_3902);
and U7589 (N_7589,N_4910,N_2071);
nor U7590 (N_7590,N_3724,N_4773);
nand U7591 (N_7591,N_1590,N_6229);
nand U7592 (N_7592,N_2062,N_1500);
nor U7593 (N_7593,N_2323,N_2420);
nor U7594 (N_7594,N_4005,N_5505);
nor U7595 (N_7595,N_5398,N_1580);
nand U7596 (N_7596,N_1730,N_401);
nor U7597 (N_7597,N_2395,N_2035);
xor U7598 (N_7598,N_3482,N_94);
nor U7599 (N_7599,N_1498,N_5654);
and U7600 (N_7600,N_317,N_5721);
nor U7601 (N_7601,N_51,N_5598);
or U7602 (N_7602,N_3809,N_2626);
and U7603 (N_7603,N_649,N_822);
nor U7604 (N_7604,N_2446,N_2921);
nor U7605 (N_7605,N_604,N_3199);
xor U7606 (N_7606,N_1396,N_5348);
nor U7607 (N_7607,N_1382,N_449);
xor U7608 (N_7608,N_286,N_5078);
or U7609 (N_7609,N_4016,N_4702);
and U7610 (N_7610,N_3390,N_6176);
and U7611 (N_7611,N_466,N_1028);
nor U7612 (N_7612,N_3883,N_2080);
and U7613 (N_7613,N_3146,N_2868);
xnor U7614 (N_7614,N_99,N_170);
nand U7615 (N_7615,N_4429,N_5464);
nor U7616 (N_7616,N_3723,N_25);
and U7617 (N_7617,N_4019,N_421);
xnor U7618 (N_7618,N_1599,N_4605);
xnor U7619 (N_7619,N_705,N_5233);
and U7620 (N_7620,N_1596,N_4081);
and U7621 (N_7621,N_1810,N_5561);
xor U7622 (N_7622,N_2004,N_186);
or U7623 (N_7623,N_1375,N_138);
nand U7624 (N_7624,N_2320,N_277);
nor U7625 (N_7625,N_5147,N_5671);
xnor U7626 (N_7626,N_4778,N_3518);
or U7627 (N_7627,N_4176,N_1759);
nor U7628 (N_7628,N_3992,N_4624);
xor U7629 (N_7629,N_4967,N_2628);
and U7630 (N_7630,N_5951,N_1941);
nand U7631 (N_7631,N_4934,N_970);
or U7632 (N_7632,N_2145,N_3655);
nor U7633 (N_7633,N_2049,N_1322);
nor U7634 (N_7634,N_5185,N_2968);
and U7635 (N_7635,N_2552,N_2698);
or U7636 (N_7636,N_4156,N_3220);
xnor U7637 (N_7637,N_885,N_2248);
nor U7638 (N_7638,N_3675,N_5609);
and U7639 (N_7639,N_1213,N_614);
xnor U7640 (N_7640,N_1691,N_3987);
nor U7641 (N_7641,N_5416,N_3707);
xnor U7642 (N_7642,N_2954,N_1622);
nor U7643 (N_7643,N_4514,N_6203);
and U7644 (N_7644,N_5156,N_796);
or U7645 (N_7645,N_3097,N_2040);
or U7646 (N_7646,N_5266,N_5411);
xnor U7647 (N_7647,N_4862,N_2091);
and U7648 (N_7648,N_3025,N_5642);
or U7649 (N_7649,N_690,N_2353);
nor U7650 (N_7650,N_2230,N_2224);
nand U7651 (N_7651,N_5857,N_2078);
xor U7652 (N_7652,N_2792,N_1995);
nand U7653 (N_7653,N_1303,N_308);
or U7654 (N_7654,N_2195,N_3686);
and U7655 (N_7655,N_5584,N_3487);
and U7656 (N_7656,N_2287,N_4262);
and U7657 (N_7657,N_96,N_5981);
and U7658 (N_7658,N_3955,N_6012);
xor U7659 (N_7659,N_6064,N_2083);
or U7660 (N_7660,N_4747,N_3060);
or U7661 (N_7661,N_6063,N_931);
xnor U7662 (N_7662,N_1875,N_2897);
nand U7663 (N_7663,N_297,N_3730);
and U7664 (N_7664,N_158,N_4080);
nor U7665 (N_7665,N_3742,N_1946);
nor U7666 (N_7666,N_2531,N_3914);
xnor U7667 (N_7667,N_3531,N_414);
nor U7668 (N_7668,N_3219,N_1417);
xnor U7669 (N_7669,N_3910,N_3880);
and U7670 (N_7670,N_1418,N_5543);
xor U7671 (N_7671,N_1714,N_309);
nor U7672 (N_7672,N_2529,N_1953);
nor U7673 (N_7673,N_658,N_2781);
and U7674 (N_7674,N_219,N_2910);
or U7675 (N_7675,N_4683,N_5196);
xor U7676 (N_7676,N_3267,N_1992);
xnor U7677 (N_7677,N_5284,N_3840);
nor U7678 (N_7678,N_436,N_4450);
or U7679 (N_7679,N_3590,N_6033);
or U7680 (N_7680,N_4265,N_810);
or U7681 (N_7681,N_4586,N_4085);
and U7682 (N_7682,N_783,N_643);
nor U7683 (N_7683,N_1611,N_224);
nand U7684 (N_7684,N_5260,N_33);
or U7685 (N_7685,N_2588,N_6145);
and U7686 (N_7686,N_4560,N_1921);
nand U7687 (N_7687,N_3455,N_886);
and U7688 (N_7688,N_1177,N_4574);
nand U7689 (N_7689,N_1070,N_4608);
or U7690 (N_7690,N_1869,N_4803);
or U7691 (N_7691,N_510,N_1779);
or U7692 (N_7692,N_2638,N_4837);
and U7693 (N_7693,N_5517,N_1215);
and U7694 (N_7694,N_6215,N_2926);
or U7695 (N_7695,N_403,N_5575);
nand U7696 (N_7696,N_1387,N_5001);
nand U7697 (N_7697,N_4167,N_3824);
nor U7698 (N_7698,N_465,N_41);
or U7699 (N_7699,N_1895,N_1065);
and U7700 (N_7700,N_363,N_2415);
nor U7701 (N_7701,N_4697,N_5907);
and U7702 (N_7702,N_3441,N_5279);
and U7703 (N_7703,N_1128,N_545);
nand U7704 (N_7704,N_5122,N_5658);
nand U7705 (N_7705,N_5975,N_5027);
and U7706 (N_7706,N_4006,N_34);
and U7707 (N_7707,N_273,N_5401);
or U7708 (N_7708,N_5522,N_4776);
xor U7709 (N_7709,N_2126,N_1790);
xor U7710 (N_7710,N_3197,N_197);
xor U7711 (N_7711,N_2389,N_1852);
nand U7712 (N_7712,N_4669,N_4487);
xnor U7713 (N_7713,N_240,N_2184);
and U7714 (N_7714,N_4309,N_4720);
nand U7715 (N_7715,N_6188,N_6191);
and U7716 (N_7716,N_5636,N_4386);
nor U7717 (N_7717,N_5616,N_4684);
xor U7718 (N_7718,N_206,N_5872);
xor U7719 (N_7719,N_2959,N_2565);
nor U7720 (N_7720,N_2438,N_517);
xnor U7721 (N_7721,N_2878,N_5570);
or U7722 (N_7722,N_3040,N_3090);
nor U7723 (N_7723,N_1581,N_1484);
nor U7724 (N_7724,N_1587,N_1753);
xnor U7725 (N_7725,N_5778,N_4410);
xor U7726 (N_7726,N_2752,N_944);
xnor U7727 (N_7727,N_3894,N_4975);
nor U7728 (N_7728,N_4492,N_3728);
xnor U7729 (N_7729,N_1139,N_1157);
xor U7730 (N_7730,N_493,N_5960);
or U7731 (N_7731,N_3214,N_6016);
xnor U7732 (N_7732,N_4405,N_3044);
xnor U7733 (N_7733,N_1780,N_4050);
or U7734 (N_7734,N_4694,N_5901);
xor U7735 (N_7735,N_2523,N_2917);
nor U7736 (N_7736,N_2103,N_4651);
nand U7737 (N_7737,N_2478,N_1809);
and U7738 (N_7738,N_867,N_613);
or U7739 (N_7739,N_4764,N_5283);
xor U7740 (N_7740,N_5107,N_824);
and U7741 (N_7741,N_4757,N_850);
nand U7742 (N_7742,N_2736,N_2577);
and U7743 (N_7743,N_1133,N_4668);
nand U7744 (N_7744,N_6067,N_4915);
and U7745 (N_7745,N_3750,N_1804);
xor U7746 (N_7746,N_1957,N_4334);
nand U7747 (N_7747,N_3301,N_4400);
nand U7748 (N_7748,N_4170,N_725);
xor U7749 (N_7749,N_1632,N_1557);
nand U7750 (N_7750,N_6017,N_2047);
nor U7751 (N_7751,N_1594,N_4029);
nand U7752 (N_7752,N_3687,N_2584);
or U7753 (N_7753,N_3317,N_588);
xnor U7754 (N_7754,N_4656,N_1302);
xor U7755 (N_7755,N_4007,N_3148);
or U7756 (N_7756,N_3186,N_5305);
nor U7757 (N_7757,N_2,N_2192);
or U7758 (N_7758,N_2929,N_2217);
and U7759 (N_7759,N_373,N_13);
nand U7760 (N_7760,N_5372,N_1546);
xnor U7761 (N_7761,N_4799,N_4114);
and U7762 (N_7762,N_5889,N_6172);
or U7763 (N_7763,N_579,N_6041);
or U7764 (N_7764,N_100,N_572);
nor U7765 (N_7765,N_172,N_2225);
and U7766 (N_7766,N_2046,N_1401);
or U7767 (N_7767,N_471,N_4607);
xor U7768 (N_7768,N_2242,N_5091);
xor U7769 (N_7769,N_1209,N_5993);
nand U7770 (N_7770,N_5125,N_4892);
nand U7771 (N_7771,N_3691,N_1901);
or U7772 (N_7772,N_1313,N_2504);
and U7773 (N_7773,N_2994,N_451);
nand U7774 (N_7774,N_1639,N_836);
nand U7775 (N_7775,N_3540,N_4128);
or U7776 (N_7776,N_5334,N_668);
or U7777 (N_7777,N_5786,N_5716);
xnor U7778 (N_7778,N_4544,N_4957);
xnor U7779 (N_7779,N_1733,N_5771);
xor U7780 (N_7780,N_611,N_2304);
nor U7781 (N_7781,N_3932,N_4564);
nand U7782 (N_7782,N_4863,N_5313);
nand U7783 (N_7783,N_4404,N_1745);
nand U7784 (N_7784,N_1125,N_5019);
nor U7785 (N_7785,N_2556,N_3024);
and U7786 (N_7786,N_1825,N_550);
or U7787 (N_7787,N_2251,N_1553);
nand U7788 (N_7788,N_1687,N_4061);
nor U7789 (N_7789,N_5675,N_1208);
nand U7790 (N_7790,N_3676,N_6124);
nor U7791 (N_7791,N_1740,N_2376);
or U7792 (N_7792,N_3101,N_3594);
nand U7793 (N_7793,N_1842,N_964);
or U7794 (N_7794,N_3308,N_1655);
or U7795 (N_7795,N_2961,N_2627);
nand U7796 (N_7796,N_2649,N_2963);
and U7797 (N_7797,N_1314,N_1068);
and U7798 (N_7798,N_5153,N_1617);
xor U7799 (N_7799,N_2786,N_3999);
xnor U7800 (N_7800,N_5560,N_1763);
and U7801 (N_7801,N_350,N_6163);
nor U7802 (N_7802,N_3421,N_4537);
nand U7803 (N_7803,N_3395,N_4587);
or U7804 (N_7804,N_3787,N_2308);
and U7805 (N_7805,N_5168,N_4614);
nand U7806 (N_7806,N_1078,N_3503);
xnor U7807 (N_7807,N_2232,N_3562);
xor U7808 (N_7808,N_671,N_3697);
and U7809 (N_7809,N_5318,N_3678);
nor U7810 (N_7810,N_1050,N_3386);
nand U7811 (N_7811,N_1166,N_5656);
xor U7812 (N_7812,N_5925,N_2335);
nand U7813 (N_7813,N_3104,N_5451);
and U7814 (N_7814,N_4406,N_5048);
or U7815 (N_7815,N_4485,N_4196);
nor U7816 (N_7816,N_4028,N_6170);
and U7817 (N_7817,N_869,N_5780);
and U7818 (N_7818,N_2764,N_1574);
or U7819 (N_7819,N_1767,N_337);
nor U7820 (N_7820,N_1938,N_3435);
and U7821 (N_7821,N_2108,N_30);
or U7822 (N_7822,N_5150,N_1811);
nor U7823 (N_7823,N_1982,N_3228);
nor U7824 (N_7824,N_1855,N_567);
or U7825 (N_7825,N_5627,N_3800);
xor U7826 (N_7826,N_3637,N_1981);
xnor U7827 (N_7827,N_4295,N_3130);
nor U7828 (N_7828,N_5324,N_2883);
nor U7829 (N_7829,N_1088,N_3938);
nand U7830 (N_7830,N_6028,N_1051);
nor U7831 (N_7831,N_2409,N_5243);
xnor U7832 (N_7832,N_2547,N_2874);
xnor U7833 (N_7833,N_675,N_6135);
or U7834 (N_7834,N_742,N_6108);
nand U7835 (N_7835,N_905,N_2499);
and U7836 (N_7836,N_4149,N_4229);
or U7837 (N_7837,N_3058,N_3213);
xnor U7838 (N_7838,N_6081,N_5311);
nor U7839 (N_7839,N_1786,N_3721);
nor U7840 (N_7840,N_578,N_3867);
xnor U7841 (N_7841,N_995,N_4318);
nor U7842 (N_7842,N_5917,N_746);
xor U7843 (N_7843,N_3080,N_2093);
xor U7844 (N_7844,N_3034,N_2130);
nand U7845 (N_7845,N_1136,N_5972);
and U7846 (N_7846,N_35,N_2113);
and U7847 (N_7847,N_1198,N_4578);
nand U7848 (N_7848,N_1532,N_5242);
and U7849 (N_7849,N_4162,N_1129);
nor U7850 (N_7850,N_5511,N_2220);
or U7851 (N_7851,N_3122,N_5498);
nand U7852 (N_7852,N_4383,N_4398);
nor U7853 (N_7853,N_5747,N_2460);
nor U7854 (N_7854,N_3851,N_4728);
nand U7855 (N_7855,N_2307,N_3671);
or U7856 (N_7856,N_6024,N_4021);
or U7857 (N_7857,N_516,N_5463);
and U7858 (N_7858,N_4573,N_4571);
nand U7859 (N_7859,N_246,N_4551);
and U7860 (N_7860,N_2255,N_2931);
or U7861 (N_7861,N_846,N_10);
and U7862 (N_7862,N_3221,N_4018);
nand U7863 (N_7863,N_5738,N_2559);
and U7864 (N_7864,N_407,N_5711);
nor U7865 (N_7865,N_5213,N_1426);
xnor U7866 (N_7866,N_4731,N_1236);
nand U7867 (N_7867,N_5459,N_1002);
xnor U7868 (N_7868,N_3961,N_1887);
and U7869 (N_7869,N_4321,N_2611);
and U7870 (N_7870,N_2106,N_5669);
nor U7871 (N_7871,N_5551,N_1092);
xor U7872 (N_7872,N_3342,N_5890);
xnor U7873 (N_7873,N_795,N_958);
nor U7874 (N_7874,N_5953,N_332);
or U7875 (N_7875,N_3778,N_3727);
nand U7876 (N_7876,N_651,N_874);
nand U7877 (N_7877,N_6097,N_1127);
nand U7878 (N_7878,N_2141,N_5199);
nand U7879 (N_7879,N_5835,N_5957);
nor U7880 (N_7880,N_2481,N_5435);
or U7881 (N_7881,N_1644,N_5621);
nand U7882 (N_7882,N_2551,N_5686);
and U7883 (N_7883,N_2640,N_142);
nand U7884 (N_7884,N_2974,N_154);
nand U7885 (N_7885,N_3201,N_5446);
nand U7886 (N_7886,N_4944,N_1816);
nor U7887 (N_7887,N_4531,N_1799);
nor U7888 (N_7888,N_3744,N_4319);
nand U7889 (N_7889,N_503,N_1235);
nor U7890 (N_7890,N_4962,N_3222);
or U7891 (N_7891,N_748,N_3775);
nand U7892 (N_7892,N_2820,N_2109);
xor U7893 (N_7893,N_3370,N_1370);
xnor U7894 (N_7894,N_5726,N_4643);
nor U7895 (N_7895,N_2092,N_2416);
and U7896 (N_7896,N_541,N_665);
nor U7897 (N_7897,N_6035,N_5766);
xor U7898 (N_7898,N_2595,N_5370);
xor U7899 (N_7899,N_1839,N_3944);
nand U7900 (N_7900,N_5395,N_5714);
nand U7901 (N_7901,N_3396,N_622);
and U7902 (N_7902,N_4228,N_5909);
nor U7903 (N_7903,N_3340,N_3246);
or U7904 (N_7904,N_1441,N_5614);
and U7905 (N_7905,N_2235,N_2313);
or U7906 (N_7906,N_318,N_2382);
or U7907 (N_7907,N_6219,N_477);
xnor U7908 (N_7908,N_543,N_5219);
nor U7909 (N_7909,N_546,N_1558);
nor U7910 (N_7910,N_2543,N_5437);
xnor U7911 (N_7911,N_460,N_1376);
nand U7912 (N_7912,N_4534,N_3460);
and U7913 (N_7913,N_5992,N_2877);
and U7914 (N_7914,N_3333,N_3152);
or U7915 (N_7915,N_201,N_1760);
or U7916 (N_7916,N_5379,N_507);
nor U7917 (N_7917,N_5781,N_1857);
nor U7918 (N_7918,N_4893,N_3123);
nand U7919 (N_7919,N_3318,N_248);
nor U7920 (N_7920,N_2451,N_2424);
nor U7921 (N_7921,N_2132,N_5650);
and U7922 (N_7922,N_4857,N_3599);
and U7923 (N_7923,N_5442,N_5591);
or U7924 (N_7924,N_592,N_2561);
nand U7925 (N_7925,N_2250,N_3731);
nor U7926 (N_7926,N_1674,N_4311);
nor U7927 (N_7927,N_932,N_3878);
xnor U7928 (N_7928,N_3820,N_3501);
nand U7929 (N_7929,N_5307,N_1390);
nand U7930 (N_7930,N_4636,N_2779);
or U7931 (N_7931,N_2958,N_1789);
xnor U7932 (N_7932,N_16,N_5633);
and U7933 (N_7933,N_5828,N_5542);
xnor U7934 (N_7934,N_556,N_5947);
xor U7935 (N_7935,N_4048,N_688);
xor U7936 (N_7936,N_5141,N_4935);
nor U7937 (N_7937,N_799,N_5717);
nand U7938 (N_7938,N_6013,N_1138);
nor U7939 (N_7939,N_4790,N_4325);
and U7940 (N_7940,N_1256,N_522);
xnor U7941 (N_7941,N_1433,N_5043);
xor U7942 (N_7942,N_4841,N_5354);
or U7943 (N_7943,N_598,N_6096);
and U7944 (N_7944,N_4997,N_4460);
xor U7945 (N_7945,N_5882,N_3072);
xor U7946 (N_7946,N_5529,N_5792);
nand U7947 (N_7947,N_250,N_581);
and U7948 (N_7948,N_2318,N_2360);
or U7949 (N_7949,N_425,N_3534);
or U7950 (N_7950,N_2214,N_842);
nand U7951 (N_7951,N_5888,N_432);
or U7952 (N_7952,N_3904,N_1977);
nand U7953 (N_7953,N_4598,N_5360);
and U7954 (N_7954,N_1571,N_4657);
or U7955 (N_7955,N_1273,N_1956);
or U7956 (N_7956,N_5651,N_2787);
nand U7957 (N_7957,N_6175,N_23);
nor U7958 (N_7958,N_1506,N_3338);
and U7959 (N_7959,N_5424,N_2462);
xor U7960 (N_7960,N_2938,N_2797);
nor U7961 (N_7961,N_3502,N_695);
nand U7962 (N_7962,N_2852,N_4808);
nand U7963 (N_7963,N_4236,N_4793);
or U7964 (N_7964,N_6222,N_1301);
nand U7965 (N_7965,N_4488,N_1654);
nor U7966 (N_7966,N_3699,N_1383);
and U7967 (N_7967,N_5837,N_5201);
or U7968 (N_7968,N_1627,N_2414);
and U7969 (N_7969,N_5808,N_4593);
nand U7970 (N_7970,N_3928,N_2728);
xor U7971 (N_7971,N_3982,N_530);
xor U7972 (N_7972,N_2775,N_2133);
nor U7973 (N_7973,N_1688,N_4240);
nor U7974 (N_7974,N_2135,N_5967);
xnor U7975 (N_7975,N_2834,N_3988);
and U7976 (N_7976,N_5853,N_2228);
or U7977 (N_7977,N_533,N_2590);
nand U7978 (N_7978,N_4556,N_305);
and U7979 (N_7979,N_984,N_1054);
nand U7980 (N_7980,N_571,N_6202);
xnor U7981 (N_7981,N_1095,N_4084);
nand U7982 (N_7982,N_4157,N_5096);
xor U7983 (N_7983,N_4308,N_972);
xnor U7984 (N_7984,N_4504,N_3056);
and U7985 (N_7985,N_5732,N_2700);
or U7986 (N_7986,N_2015,N_4736);
nor U7987 (N_7987,N_1847,N_150);
or U7988 (N_7988,N_2518,N_4417);
or U7989 (N_7989,N_3536,N_1643);
and U7990 (N_7990,N_1913,N_634);
nand U7991 (N_7991,N_1281,N_5832);
xnor U7992 (N_7992,N_284,N_492);
nor U7993 (N_7993,N_743,N_2150);
xnor U7994 (N_7994,N_5368,N_2472);
or U7995 (N_7995,N_728,N_603);
nor U7996 (N_7996,N_3615,N_2512);
nand U7997 (N_7997,N_5563,N_3661);
xnor U7998 (N_7998,N_4000,N_1350);
xor U7999 (N_7999,N_1310,N_4765);
and U8000 (N_8000,N_4474,N_6105);
xnor U8001 (N_8001,N_4871,N_5652);
and U8002 (N_8002,N_5030,N_2527);
or U8003 (N_8003,N_2146,N_2605);
nand U8004 (N_8004,N_566,N_3051);
and U8005 (N_8005,N_1918,N_5074);
nor U8006 (N_8006,N_2464,N_4345);
nor U8007 (N_8007,N_3245,N_5128);
xor U8008 (N_8008,N_3860,N_1787);
nor U8009 (N_8009,N_773,N_2125);
and U8010 (N_8010,N_2631,N_3815);
and U8011 (N_8011,N_6051,N_5672);
and U8012 (N_8012,N_1821,N_5659);
nand U8013 (N_8013,N_1216,N_6083);
and U8014 (N_8014,N_2443,N_437);
or U8015 (N_8015,N_520,N_327);
xor U8016 (N_8016,N_2147,N_5443);
nand U8017 (N_8017,N_631,N_92);
nand U8018 (N_8018,N_1333,N_3600);
xor U8019 (N_8019,N_2087,N_4506);
or U8020 (N_8020,N_39,N_2290);
nor U8021 (N_8021,N_1480,N_1373);
and U8022 (N_8022,N_3016,N_2763);
xnor U8023 (N_8023,N_3046,N_2557);
nor U8024 (N_8024,N_1915,N_1369);
and U8025 (N_8025,N_5462,N_2284);
nor U8026 (N_8026,N_15,N_6052);
nor U8027 (N_8027,N_2452,N_312);
nand U8028 (N_8028,N_1755,N_2116);
xnor U8029 (N_8029,N_1819,N_2021);
nand U8030 (N_8030,N_1048,N_5325);
or U8031 (N_8031,N_146,N_3837);
and U8032 (N_8032,N_495,N_2532);
or U8033 (N_8033,N_1326,N_5665);
nand U8034 (N_8034,N_2266,N_5404);
nand U8035 (N_8035,N_5519,N_3144);
xor U8036 (N_8036,N_2115,N_2940);
nor U8037 (N_8037,N_1040,N_1450);
and U8038 (N_8038,N_560,N_293);
xor U8039 (N_8039,N_3295,N_2485);
nand U8040 (N_8040,N_3652,N_986);
xnor U8041 (N_8041,N_4734,N_5439);
and U8042 (N_8042,N_5140,N_4177);
xnor U8043 (N_8043,N_5722,N_1516);
nand U8044 (N_8044,N_2439,N_204);
and U8045 (N_8045,N_5536,N_213);
nand U8046 (N_8046,N_1848,N_5861);
or U8047 (N_8047,N_5296,N_4188);
nor U8048 (N_8048,N_2795,N_554);
xnor U8049 (N_8049,N_2583,N_4095);
xnor U8050 (N_8050,N_2349,N_763);
or U8051 (N_8051,N_3491,N_1257);
nand U8052 (N_8052,N_4092,N_6043);
nand U8053 (N_8053,N_3725,N_1647);
nor U8054 (N_8054,N_4097,N_6185);
nand U8055 (N_8055,N_491,N_4768);
and U8056 (N_8056,N_3043,N_4272);
and U8057 (N_8057,N_5162,N_5034);
and U8058 (N_8058,N_3351,N_4856);
and U8059 (N_8059,N_2102,N_1242);
and U8060 (N_8060,N_453,N_3155);
nor U8061 (N_8061,N_2695,N_765);
or U8062 (N_8062,N_5172,N_1994);
and U8063 (N_8063,N_3205,N_2530);
nand U8064 (N_8064,N_5084,N_139);
nor U8065 (N_8065,N_2437,N_4623);
nor U8066 (N_8066,N_38,N_1766);
xor U8067 (N_8067,N_3260,N_832);
xor U8068 (N_8068,N_5615,N_333);
nand U8069 (N_8069,N_5109,N_5691);
nor U8070 (N_8070,N_3667,N_4098);
nor U8071 (N_8071,N_5723,N_4415);
and U8072 (N_8072,N_3012,N_1098);
or U8073 (N_8073,N_5515,N_5248);
and U8074 (N_8074,N_3714,N_5497);
nor U8075 (N_8075,N_79,N_56);
nor U8076 (N_8076,N_5927,N_3031);
nand U8077 (N_8077,N_1014,N_2869);
nor U8078 (N_8078,N_1778,N_3719);
and U8079 (N_8079,N_5426,N_3473);
nor U8080 (N_8080,N_5764,N_4039);
or U8081 (N_8081,N_1881,N_2168);
xor U8082 (N_8082,N_5490,N_1266);
nor U8083 (N_8083,N_315,N_1600);
nand U8084 (N_8084,N_2493,N_3149);
nand U8085 (N_8085,N_1970,N_1530);
nand U8086 (N_8086,N_508,N_6140);
xnor U8087 (N_8087,N_2635,N_3429);
or U8088 (N_8088,N_1296,N_3077);
xor U8089 (N_8089,N_2880,N_5552);
and U8090 (N_8090,N_3279,N_1681);
nand U8091 (N_8091,N_2010,N_1676);
or U8092 (N_8092,N_6029,N_3042);
or U8093 (N_8093,N_4767,N_14);
and U8094 (N_8094,N_692,N_4644);
xor U8095 (N_8095,N_2274,N_5727);
nor U8096 (N_8096,N_5270,N_241);
or U8097 (N_8097,N_6227,N_5797);
and U8098 (N_8098,N_3158,N_4966);
xor U8099 (N_8099,N_4425,N_2343);
xor U8100 (N_8100,N_5707,N_1700);
nand U8101 (N_8101,N_6243,N_125);
xnor U8102 (N_8102,N_1891,N_1524);
nor U8103 (N_8103,N_617,N_5101);
and U8104 (N_8104,N_3405,N_4851);
and U8105 (N_8105,N_2839,N_865);
nor U8106 (N_8106,N_4034,N_2686);
nand U8107 (N_8107,N_2454,N_4621);
xor U8108 (N_8108,N_5956,N_2226);
or U8109 (N_8109,N_4839,N_2906);
or U8110 (N_8110,N_1066,N_2127);
xor U8111 (N_8111,N_1063,N_2849);
or U8112 (N_8112,N_861,N_3673);
nor U8113 (N_8113,N_52,N_4401);
nand U8114 (N_8114,N_2539,N_6023);
nand U8115 (N_8115,N_5297,N_1114);
and U8116 (N_8116,N_1862,N_1603);
xor U8117 (N_8117,N_4978,N_5115);
xor U8118 (N_8118,N_1987,N_5023);
nand U8119 (N_8119,N_1377,N_4549);
nand U8120 (N_8120,N_1415,N_3407);
or U8121 (N_8121,N_3093,N_1722);
or U8122 (N_8122,N_2646,N_3120);
nand U8123 (N_8123,N_5067,N_4008);
nor U8124 (N_8124,N_3138,N_628);
and U8125 (N_8125,N_3611,N_5902);
nand U8126 (N_8126,N_734,N_4703);
nand U8127 (N_8127,N_2411,N_1495);
xor U8128 (N_8128,N_3341,N_5594);
or U8129 (N_8129,N_2805,N_4898);
nor U8130 (N_8130,N_6151,N_4964);
or U8131 (N_8131,N_4099,N_5877);
nand U8132 (N_8132,N_3995,N_3722);
and U8133 (N_8133,N_1517,N_3236);
or U8134 (N_8134,N_4274,N_274);
nor U8135 (N_8135,N_999,N_2730);
nand U8136 (N_8136,N_3589,N_2162);
nor U8137 (N_8137,N_3926,N_1204);
and U8138 (N_8138,N_2476,N_2814);
and U8139 (N_8139,N_1312,N_5431);
xnor U8140 (N_8140,N_3353,N_2356);
xnor U8141 (N_8141,N_3726,N_770);
and U8142 (N_8142,N_5805,N_5338);
nor U8143 (N_8143,N_3528,N_2625);
nand U8144 (N_8144,N_351,N_5272);
or U8145 (N_8145,N_1974,N_3578);
xnor U8146 (N_8146,N_3226,N_5302);
and U8147 (N_8147,N_5503,N_3931);
nand U8148 (N_8148,N_1263,N_3382);
xor U8149 (N_8149,N_2754,N_2272);
or U8150 (N_8150,N_5843,N_3717);
nor U8151 (N_8151,N_5137,N_4053);
and U8152 (N_8152,N_2077,N_2055);
or U8153 (N_8153,N_4552,N_6117);
and U8154 (N_8154,N_2196,N_2965);
or U8155 (N_8155,N_4866,N_3153);
xor U8156 (N_8156,N_4509,N_1720);
or U8157 (N_8157,N_5157,N_3300);
nand U8158 (N_8158,N_1734,N_5688);
xnor U8159 (N_8159,N_2579,N_3426);
nor U8160 (N_8160,N_3157,N_4070);
nand U8161 (N_8161,N_5110,N_774);
nor U8162 (N_8162,N_2187,N_768);
nor U8163 (N_8163,N_5948,N_5885);
xnor U8164 (N_8164,N_5085,N_4937);
xor U8165 (N_8165,N_866,N_1864);
and U8166 (N_8166,N_6082,N_794);
nand U8167 (N_8167,N_2206,N_5131);
or U8168 (N_8168,N_3311,N_4178);
nor U8169 (N_8169,N_674,N_3559);
and U8170 (N_8170,N_5452,N_1924);
or U8171 (N_8171,N_6146,N_2708);
nand U8172 (N_8172,N_3834,N_386);
xnor U8173 (N_8173,N_2846,N_6126);
xnor U8174 (N_8174,N_4989,N_4836);
xor U8175 (N_8175,N_3286,N_3930);
xor U8176 (N_8176,N_1403,N_279);
nand U8177 (N_8177,N_3306,N_4001);
nor U8178 (N_8178,N_3088,N_2300);
or U8179 (N_8179,N_3517,N_851);
and U8180 (N_8180,N_4035,N_4517);
xnor U8181 (N_8181,N_3352,N_1709);
xnor U8182 (N_8182,N_3378,N_4350);
nor U8183 (N_8183,N_835,N_5222);
nand U8184 (N_8184,N_88,N_883);
nor U8185 (N_8185,N_6102,N_379);
and U8186 (N_8186,N_5858,N_3996);
or U8187 (N_8187,N_5933,N_6002);
and U8188 (N_8188,N_806,N_1328);
nand U8189 (N_8189,N_1458,N_1664);
xor U8190 (N_8190,N_3521,N_320);
and U8191 (N_8191,N_2677,N_3854);
nor U8192 (N_8192,N_4524,N_4539);
and U8193 (N_8193,N_445,N_2393);
or U8194 (N_8194,N_3738,N_4505);
and U8195 (N_8195,N_5226,N_3604);
or U8196 (N_8196,N_1649,N_3464);
nand U8197 (N_8197,N_4663,N_3939);
or U8198 (N_8198,N_2082,N_3374);
or U8199 (N_8199,N_4038,N_2662);
and U8200 (N_8200,N_4707,N_3388);
xnor U8201 (N_8201,N_4521,N_2350);
nor U8202 (N_8202,N_3957,N_4951);
nor U8203 (N_8203,N_1339,N_1926);
xnor U8204 (N_8204,N_1398,N_433);
nor U8205 (N_8205,N_5632,N_655);
nand U8206 (N_8206,N_5000,N_4079);
xor U8207 (N_8207,N_2199,N_948);
xnor U8208 (N_8208,N_864,N_4352);
nor U8209 (N_8209,N_5182,N_5831);
nor U8210 (N_8210,N_1723,N_5341);
xor U8211 (N_8211,N_3467,N_3179);
xor U8212 (N_8212,N_1280,N_5564);
or U8213 (N_8213,N_3591,N_3489);
and U8214 (N_8214,N_2546,N_2581);
and U8215 (N_8215,N_3397,N_3210);
nor U8216 (N_8216,N_2484,N_5596);
nor U8217 (N_8217,N_3250,N_969);
xor U8218 (N_8218,N_4988,N_4498);
xor U8219 (N_8219,N_5970,N_5472);
nand U8220 (N_8220,N_479,N_923);
and U8221 (N_8221,N_2899,N_793);
xor U8222 (N_8222,N_2985,N_819);
xor U8223 (N_8223,N_2911,N_1567);
and U8224 (N_8224,N_3021,N_1359);
or U8225 (N_8225,N_3448,N_5618);
nand U8226 (N_8226,N_666,N_450);
xnor U8227 (N_8227,N_275,N_3716);
nand U8228 (N_8228,N_310,N_188);
nand U8229 (N_8229,N_5241,N_1291);
nor U8230 (N_8230,N_3216,N_1937);
or U8231 (N_8231,N_862,N_2014);
or U8232 (N_8232,N_5011,N_6221);
nor U8233 (N_8233,N_1988,N_791);
xor U8234 (N_8234,N_6091,N_5470);
nor U8235 (N_8235,N_5548,N_5056);
and U8236 (N_8236,N_2269,N_5852);
nand U8237 (N_8237,N_1260,N_4234);
xor U8238 (N_8238,N_3211,N_3166);
and U8239 (N_8239,N_1525,N_3951);
or U8240 (N_8240,N_4548,N_4172);
nor U8241 (N_8241,N_1933,N_4610);
nor U8242 (N_8242,N_5860,N_2277);
xnor U8243 (N_8243,N_5350,N_4110);
nand U8244 (N_8244,N_2816,N_4673);
or U8245 (N_8245,N_2253,N_525);
nor U8246 (N_8246,N_2363,N_3729);
nor U8247 (N_8247,N_3192,N_2500);
nand U8248 (N_8248,N_3115,N_105);
nand U8249 (N_8249,N_2796,N_1072);
and U8250 (N_8250,N_412,N_660);
or U8251 (N_8251,N_1993,N_4512);
and U8252 (N_8252,N_4942,N_4843);
nand U8253 (N_8253,N_5744,N_1347);
nand U8254 (N_8254,N_1667,N_53);
and U8255 (N_8255,N_5879,N_2819);
and U8256 (N_8256,N_3648,N_2885);
nor U8257 (N_8257,N_223,N_1807);
xor U8258 (N_8258,N_4493,N_5750);
and U8259 (N_8259,N_3004,N_5818);
or U8260 (N_8260,N_2856,N_1467);
xor U8261 (N_8261,N_3670,N_3803);
xor U8262 (N_8262,N_1540,N_3432);
nor U8263 (N_8263,N_4846,N_1971);
or U8264 (N_8264,N_4132,N_1870);
nor U8265 (N_8265,N_3568,N_1404);
nor U8266 (N_8266,N_1438,N_3546);
xnor U8267 (N_8267,N_582,N_3922);
nand U8268 (N_8268,N_1940,N_5694);
or U8269 (N_8269,N_3907,N_2972);
xor U8270 (N_8270,N_2721,N_87);
nand U8271 (N_8271,N_816,N_857);
nand U8272 (N_8272,N_1461,N_5777);
nand U8273 (N_8273,N_1840,N_4227);
or U8274 (N_8274,N_3383,N_831);
xor U8275 (N_8275,N_4907,N_441);
nor U8276 (N_8276,N_5209,N_5132);
or U8277 (N_8277,N_1289,N_4502);
nor U8278 (N_8278,N_1113,N_3570);
nor U8279 (N_8279,N_2812,N_4313);
or U8280 (N_8280,N_877,N_2408);
nand U8281 (N_8281,N_1253,N_114);
and U8282 (N_8282,N_3299,N_2458);
nor U8283 (N_8283,N_1708,N_340);
nor U8284 (N_8284,N_2400,N_6065);
or U8285 (N_8285,N_1077,N_4511);
and U8286 (N_8286,N_4482,N_6072);
xor U8287 (N_8287,N_6205,N_5657);
or U8288 (N_8288,N_5588,N_6079);
and U8289 (N_8289,N_2717,N_5998);
and U8290 (N_8290,N_162,N_5776);
or U8291 (N_8291,N_856,N_5304);
nand U8292 (N_8292,N_6195,N_2005);
xnor U8293 (N_8293,N_1635,N_4472);
and U8294 (N_8294,N_5949,N_5218);
or U8295 (N_8295,N_2275,N_2241);
xor U8296 (N_8296,N_755,N_2502);
or U8297 (N_8297,N_111,N_2997);
xor U8298 (N_8298,N_209,N_5863);
and U8299 (N_8299,N_4186,N_4340);
and U8300 (N_8300,N_1011,N_5203);
or U8301 (N_8301,N_513,N_6110);
nor U8302 (N_8302,N_2067,N_1147);
and U8303 (N_8303,N_290,N_3545);
or U8304 (N_8304,N_1082,N_5038);
xor U8305 (N_8305,N_1084,N_4258);
or U8306 (N_8306,N_1442,N_715);
nand U8307 (N_8307,N_1812,N_3252);
nor U8308 (N_8308,N_1234,N_4763);
nand U8309 (N_8309,N_1663,N_4947);
and U8310 (N_8310,N_5261,N_193);
or U8311 (N_8311,N_717,N_713);
or U8312 (N_8312,N_872,N_3798);
nand U8313 (N_8313,N_526,N_2654);
and U8314 (N_8314,N_396,N_2325);
nand U8315 (N_8315,N_2017,N_4750);
and U8316 (N_8316,N_3974,N_3639);
and U8317 (N_8317,N_4430,N_2246);
nor U8318 (N_8318,N_4199,N_5363);
or U8319 (N_8319,N_6101,N_1598);
nor U8320 (N_8320,N_839,N_4555);
xor U8321 (N_8321,N_1330,N_4735);
and U8322 (N_8322,N_4746,N_1833);
xnor U8323 (N_8323,N_2514,N_5678);
xor U8324 (N_8324,N_5976,N_2373);
nand U8325 (N_8325,N_840,N_211);
xnor U8326 (N_8326,N_5077,N_3616);
xnor U8327 (N_8327,N_3757,N_2301);
and U8328 (N_8328,N_483,N_2582);
or U8329 (N_8329,N_285,N_2012);
and U8330 (N_8330,N_762,N_3781);
or U8331 (N_8331,N_5134,N_1526);
xor U8332 (N_8332,N_881,N_439);
or U8333 (N_8333,N_4787,N_1828);
nor U8334 (N_8334,N_3526,N_3683);
and U8335 (N_8335,N_4840,N_699);
and U8336 (N_8336,N_2916,N_169);
or U8337 (N_8337,N_3839,N_3627);
xnor U8338 (N_8338,N_1255,N_3774);
nand U8339 (N_8339,N_5445,N_843);
or U8340 (N_8340,N_155,N_3091);
nor U8341 (N_8341,N_1468,N_5380);
xor U8342 (N_8342,N_3187,N_1201);
and U8343 (N_8343,N_1219,N_2862);
xor U8344 (N_8344,N_2884,N_4695);
or U8345 (N_8345,N_126,N_6014);
nand U8346 (N_8346,N_4974,N_1845);
nand U8347 (N_8347,N_1527,N_3302);
and U8348 (N_8348,N_2519,N_3710);
xnor U8349 (N_8349,N_6068,N_356);
nand U8350 (N_8350,N_5924,N_5215);
nand U8351 (N_8351,N_4168,N_4022);
and U8352 (N_8352,N_4083,N_4972);
or U8353 (N_8353,N_6090,N_5962);
xor U8354 (N_8354,N_3334,N_4688);
nand U8355 (N_8355,N_1456,N_5649);
or U8356 (N_8356,N_6000,N_178);
xnor U8357 (N_8357,N_4023,N_4250);
nand U8358 (N_8358,N_2379,N_4438);
or U8359 (N_8359,N_584,N_2737);
or U8360 (N_8360,N_83,N_348);
and U8361 (N_8361,N_3401,N_1503);
nand U8362 (N_8362,N_3762,N_2859);
nor U8363 (N_8363,N_5181,N_2487);
and U8364 (N_8364,N_1285,N_6032);
nor U8365 (N_8365,N_1756,N_1626);
xor U8366 (N_8366,N_2918,N_5500);
and U8367 (N_8367,N_5749,N_4729);
nor U8368 (N_8368,N_4503,N_1960);
and U8369 (N_8369,N_5022,N_5783);
and U8370 (N_8370,N_539,N_1272);
nand U8371 (N_8371,N_4422,N_6147);
xnor U8372 (N_8372,N_5930,N_5240);
nor U8373 (N_8373,N_31,N_821);
xnor U8374 (N_8374,N_5064,N_739);
nand U8375 (N_8375,N_6193,N_70);
xnor U8376 (N_8376,N_642,N_1007);
nand U8377 (N_8377,N_367,N_5789);
and U8378 (N_8378,N_3313,N_3287);
and U8379 (N_8379,N_5539,N_4390);
nand U8380 (N_8380,N_5308,N_5114);
nor U8381 (N_8381,N_5631,N_5254);
nand U8382 (N_8382,N_2657,N_1739);
nor U8383 (N_8383,N_756,N_1860);
and U8384 (N_8384,N_4466,N_5731);
xnor U8385 (N_8385,N_5667,N_2920);
and U8386 (N_8386,N_5293,N_5929);
or U8387 (N_8387,N_4815,N_5188);
or U8388 (N_8388,N_3266,N_702);
or U8389 (N_8389,N_5407,N_210);
nand U8390 (N_8390,N_397,N_681);
and U8391 (N_8391,N_2120,N_610);
nand U8392 (N_8392,N_1794,N_5482);
xor U8393 (N_8393,N_2009,N_5480);
nor U8394 (N_8394,N_4148,N_2099);
or U8395 (N_8395,N_1405,N_1111);
nor U8396 (N_8396,N_1083,N_1584);
xnor U8397 (N_8397,N_1619,N_73);
and U8398 (N_8398,N_4353,N_605);
nor U8399 (N_8399,N_5773,N_1024);
and U8400 (N_8400,N_6231,N_1089);
nand U8401 (N_8401,N_2840,N_4442);
nand U8402 (N_8402,N_4124,N_4235);
or U8403 (N_8403,N_5931,N_2580);
and U8404 (N_8404,N_1493,N_3293);
nor U8405 (N_8405,N_2209,N_4459);
or U8406 (N_8406,N_3651,N_2629);
and U8407 (N_8407,N_2193,N_387);
and U8408 (N_8408,N_3506,N_3290);
and U8409 (N_8409,N_4372,N_5040);
nor U8410 (N_8410,N_4130,N_4601);
or U8411 (N_8411,N_5276,N_1979);
and U8412 (N_8412,N_4268,N_1406);
and U8413 (N_8413,N_4246,N_707);
nand U8414 (N_8414,N_1832,N_4838);
and U8415 (N_8415,N_6061,N_1775);
and U8416 (N_8416,N_1798,N_1856);
nand U8417 (N_8417,N_5846,N_4339);
xnor U8418 (N_8418,N_497,N_2924);
or U8419 (N_8419,N_5980,N_5035);
nor U8420 (N_8420,N_4047,N_313);
and U8421 (N_8421,N_1711,N_6164);
or U8422 (N_8422,N_456,N_4158);
or U8423 (N_8423,N_6104,N_4798);
nor U8424 (N_8424,N_5394,N_3129);
nor U8425 (N_8425,N_3117,N_8);
and U8426 (N_8426,N_4344,N_1899);
and U8427 (N_8427,N_5664,N_4010);
nor U8428 (N_8428,N_1393,N_3440);
nor U8429 (N_8429,N_369,N_652);
and U8430 (N_8430,N_5100,N_3305);
nand U8431 (N_8431,N_4413,N_1658);
nand U8432 (N_8432,N_4120,N_3756);
nor U8433 (N_8433,N_4540,N_5820);
and U8434 (N_8434,N_3456,N_3118);
nor U8435 (N_8435,N_2562,N_521);
xnor U8436 (N_8436,N_1883,N_2823);
and U8437 (N_8437,N_2944,N_2889);
xor U8438 (N_8438,N_2208,N_5549);
nor U8439 (N_8439,N_3000,N_5566);
xor U8440 (N_8440,N_472,N_2239);
xor U8441 (N_8441,N_3786,N_1620);
nand U8442 (N_8442,N_3879,N_4043);
nor U8443 (N_8443,N_134,N_3718);
xor U8444 (N_8444,N_3168,N_1545);
nor U8445 (N_8445,N_3660,N_4650);
and U8446 (N_8446,N_1009,N_1448);
xor U8447 (N_8447,N_3945,N_1019);
nand U8448 (N_8448,N_4275,N_4198);
nor U8449 (N_8449,N_1890,N_5192);
nor U8450 (N_8450,N_2201,N_6218);
or U8451 (N_8451,N_2865,N_4322);
xor U8452 (N_8452,N_852,N_2200);
nor U8453 (N_8453,N_1732,N_4732);
and U8454 (N_8454,N_3014,N_4118);
or U8455 (N_8455,N_1033,N_3243);
nor U8456 (N_8456,N_4294,N_4620);
and U8457 (N_8457,N_826,N_5639);
xor U8458 (N_8458,N_3323,N_5423);
xnor U8459 (N_8459,N_5124,N_5429);
xnor U8460 (N_8460,N_3632,N_2603);
nor U8461 (N_8461,N_6078,N_4535);
xnor U8462 (N_8462,N_3794,N_2054);
nand U8463 (N_8463,N_4195,N_1483);
and U8464 (N_8464,N_2609,N_5502);
nor U8465 (N_8465,N_1962,N_5913);
or U8466 (N_8466,N_3593,N_1267);
nor U8467 (N_8467,N_2772,N_4249);
nand U8468 (N_8468,N_2864,N_4546);
or U8469 (N_8469,N_6184,N_6178);
nor U8470 (N_8470,N_1361,N_6141);
nand U8471 (N_8471,N_2851,N_2742);
or U8472 (N_8472,N_5765,N_1161);
nor U8473 (N_8473,N_2710,N_3868);
nand U8474 (N_8474,N_4447,N_384);
nand U8475 (N_8475,N_2032,N_5413);
nor U8476 (N_8476,N_5774,N_5790);
nor U8477 (N_8477,N_3836,N_222);
and U8478 (N_8478,N_4789,N_4685);
xnor U8479 (N_8479,N_1023,N_802);
and U8480 (N_8480,N_4606,N_1486);
and U8481 (N_8481,N_1662,N_5239);
nand U8482 (N_8482,N_2776,N_4011);
xnor U8483 (N_8483,N_2615,N_2157);
or U8484 (N_8484,N_3547,N_1150);
and U8485 (N_8485,N_5710,N_4002);
xnor U8486 (N_8486,N_5349,N_2131);
or U8487 (N_8487,N_3917,N_4956);
nand U8488 (N_8488,N_1945,N_968);
xor U8489 (N_8489,N_4945,N_260);
and U8490 (N_8490,N_4224,N_1564);
and U8491 (N_8491,N_1162,N_2735);
or U8492 (N_8492,N_3189,N_4882);
xnor U8493 (N_8493,N_5965,N_940);
and U8494 (N_8494,N_640,N_917);
xor U8495 (N_8495,N_5432,N_229);
nor U8496 (N_8496,N_2925,N_1145);
nand U8497 (N_8497,N_3178,N_5724);
or U8498 (N_8498,N_4374,N_2186);
nor U8499 (N_8499,N_5400,N_1121);
and U8500 (N_8500,N_535,N_6204);
xnor U8501 (N_8501,N_685,N_1731);
nand U8502 (N_8502,N_1102,N_381);
nand U8503 (N_8503,N_5340,N_2374);
xor U8504 (N_8504,N_253,N_1284);
nand U8505 (N_8505,N_29,N_4891);
or U8506 (N_8506,N_1163,N_5008);
and U8507 (N_8507,N_4378,N_3366);
or U8508 (N_8508,N_5171,N_2589);
and U8509 (N_8509,N_2766,N_3013);
and U8510 (N_8510,N_4902,N_2507);
or U8511 (N_8511,N_664,N_5208);
nor U8512 (N_8512,N_5791,N_2986);
nand U8513 (N_8513,N_876,N_1305);
and U8514 (N_8514,N_3202,N_5055);
nor U8515 (N_8515,N_3369,N_5046);
xnor U8516 (N_8516,N_27,N_1344);
xnor U8517 (N_8517,N_942,N_428);
xor U8518 (N_8518,N_242,N_1196);
nand U8519 (N_8519,N_3041,N_5585);
nand U8520 (N_8520,N_5754,N_4991);
and U8521 (N_8521,N_447,N_6154);
and U8522 (N_8522,N_5733,N_2428);
and U8523 (N_8523,N_2194,N_4529);
nor U8524 (N_8524,N_5259,N_3830);
nor U8525 (N_8525,N_935,N_5602);
nand U8526 (N_8526,N_1671,N_798);
or U8527 (N_8527,N_360,N_1761);
or U8528 (N_8528,N_772,N_1830);
and U8529 (N_8529,N_271,N_4580);
nand U8530 (N_8530,N_4056,N_2474);
and U8531 (N_8531,N_3229,N_461);
nor U8532 (N_8532,N_2540,N_4588);
and U8533 (N_8533,N_4938,N_1925);
and U8534 (N_8534,N_2934,N_5382);
nor U8535 (N_8535,N_4792,N_5661);
xor U8536 (N_8536,N_143,N_364);
nor U8537 (N_8537,N_1012,N_4977);
and U8538 (N_8538,N_1151,N_2687);
nand U8539 (N_8539,N_2575,N_1123);
xor U8540 (N_8540,N_2888,N_1306);
nor U8541 (N_8541,N_1194,N_3131);
xor U8542 (N_8542,N_5059,N_2526);
nor U8543 (N_8543,N_3303,N_1352);
and U8544 (N_8544,N_4899,N_5607);
nor U8545 (N_8545,N_1099,N_3551);
nor U8546 (N_8546,N_3614,N_4655);
and U8547 (N_8547,N_1930,N_4914);
or U8548 (N_8548,N_6115,N_3224);
nand U8549 (N_8549,N_3037,N_5224);
xnor U8550 (N_8550,N_5812,N_1593);
and U8551 (N_8551,N_941,N_122);
xnor U8552 (N_8552,N_3127,N_5155);
xnor U8553 (N_8553,N_3344,N_5741);
nand U8554 (N_8554,N_5469,N_1252);
nand U8555 (N_8555,N_5693,N_22);
nor U8556 (N_8556,N_5827,N_2441);
or U8557 (N_8557,N_2784,N_1781);
xor U8558 (N_8558,N_2850,N_423);
xor U8559 (N_8559,N_3813,N_6226);
xnor U8560 (N_8560,N_4326,N_3463);
or U8561 (N_8561,N_1808,N_4426);
or U8562 (N_8562,N_2845,N_5787);
xor U8563 (N_8563,N_6244,N_4924);
and U8564 (N_8564,N_3763,N_1897);
or U8565 (N_8565,N_3404,N_2306);
nor U8566 (N_8566,N_3695,N_2503);
and U8567 (N_8567,N_4592,N_3017);
and U8568 (N_8568,N_1606,N_4279);
xnor U8569 (N_8569,N_4152,N_1494);
nand U8570 (N_8570,N_4183,N_4770);
or U8571 (N_8571,N_2733,N_5420);
nor U8572 (N_8572,N_4686,N_264);
and U8573 (N_8573,N_2154,N_4829);
nor U8574 (N_8574,N_3967,N_3298);
nand U8575 (N_8575,N_3749,N_6199);
xnor U8576 (N_8576,N_3023,N_2788);
nand U8577 (N_8577,N_1543,N_902);
nor U8578 (N_8578,N_3776,N_411);
nor U8579 (N_8579,N_2037,N_3841);
or U8580 (N_8580,N_3454,N_947);
nand U8581 (N_8581,N_721,N_3643);
nor U8582 (N_8582,N_36,N_5855);
xor U8583 (N_8583,N_1117,N_5184);
and U8584 (N_8584,N_6034,N_2895);
and U8585 (N_8585,N_78,N_5235);
nand U8586 (N_8586,N_3634,N_3431);
nor U8587 (N_8587,N_2403,N_1837);
nor U8588 (N_8588,N_2973,N_3755);
nor U8589 (N_8589,N_3556,N_6150);
xor U8590 (N_8590,N_2913,N_3620);
and U8591 (N_8591,N_5518,N_4604);
nor U8592 (N_8592,N_2511,N_2022);
and U8593 (N_8593,N_718,N_410);
nor U8594 (N_8594,N_3826,N_69);
or U8595 (N_8595,N_6004,N_3541);
nor U8596 (N_8596,N_1171,N_301);
and U8597 (N_8597,N_2121,N_2236);
or U8598 (N_8598,N_4342,N_2950);
and U8599 (N_8599,N_321,N_2368);
xnor U8600 (N_8600,N_230,N_4393);
nor U8601 (N_8601,N_4648,N_4069);
xor U8602 (N_8602,N_3855,N_3265);
and U8603 (N_8603,N_174,N_939);
nor U8604 (N_8604,N_1436,N_1531);
xnor U8605 (N_8605,N_4884,N_2534);
and U8606 (N_8606,N_3555,N_2011);
nand U8607 (N_8607,N_4329,N_4201);
and U8608 (N_8608,N_4905,N_5444);
nand U8609 (N_8609,N_4112,N_5460);
and U8610 (N_8610,N_4733,N_5024);
and U8611 (N_8611,N_4068,N_3420);
nor U8612 (N_8612,N_4239,N_5385);
nand U8613 (N_8613,N_4847,N_745);
nor U8614 (N_8614,N_4522,N_4116);
and U8615 (N_8615,N_3377,N_5488);
nor U8616 (N_8616,N_4525,N_1575);
and U8617 (N_8617,N_4923,N_5383);
xnor U8618 (N_8618,N_269,N_5232);
nor U8619 (N_8619,N_1521,N_814);
xnor U8620 (N_8620,N_2644,N_1335);
or U8621 (N_8621,N_3831,N_4804);
nand U8622 (N_8622,N_419,N_4609);
nand U8623 (N_8623,N_5310,N_1695);
nor U8624 (N_8624,N_2459,N_6120);
xor U8625 (N_8625,N_2669,N_1334);
xor U8626 (N_8626,N_3188,N_1955);
xnor U8627 (N_8627,N_1299,N_801);
nand U8628 (N_8628,N_232,N_1782);
and U8629 (N_8629,N_2783,N_1307);
xor U8630 (N_8630,N_2095,N_4346);
and U8631 (N_8631,N_2278,N_4590);
or U8632 (N_8632,N_4458,N_4660);
nor U8633 (N_8633,N_2536,N_380);
nor U8634 (N_8634,N_4939,N_4306);
or U8635 (N_8635,N_4865,N_596);
nor U8636 (N_8636,N_402,N_1206);
or U8637 (N_8637,N_1487,N_981);
nor U8638 (N_8638,N_4519,N_304);
nor U8639 (N_8639,N_5944,N_4542);
nor U8640 (N_8640,N_1706,N_3785);
nor U8641 (N_8641,N_3196,N_131);
nor U8642 (N_8642,N_5033,N_243);
xnor U8643 (N_8643,N_5118,N_3392);
or U8644 (N_8644,N_3320,N_3818);
and U8645 (N_8645,N_3355,N_417);
nor U8646 (N_8646,N_1873,N_4088);
or U8647 (N_8647,N_3481,N_3580);
xnor U8648 (N_8648,N_5306,N_3478);
and U8649 (N_8649,N_915,N_6103);
nor U8650 (N_8650,N_3630,N_3849);
nor U8651 (N_8651,N_2655,N_1838);
or U8652 (N_8652,N_4361,N_2260);
or U8653 (N_8653,N_1479,N_4791);
nand U8654 (N_8654,N_2221,N_375);
xor U8655 (N_8655,N_2397,N_3703);
xnor U8656 (N_8656,N_5785,N_4151);
nand U8657 (N_8657,N_5922,N_5456);
and U8658 (N_8658,N_4031,N_4897);
nand U8659 (N_8659,N_1773,N_4691);
or U8660 (N_8660,N_5950,N_2802);
xor U8661 (N_8661,N_394,N_4705);
nor U8662 (N_8662,N_4484,N_3793);
and U8663 (N_8663,N_4500,N_859);
xnor U8664 (N_8664,N_3596,N_1548);
nor U8665 (N_8665,N_314,N_4877);
and U8666 (N_8666,N_1294,N_838);
and U8667 (N_8667,N_5898,N_3801);
or U8668 (N_8668,N_911,N_3289);
xnor U8669 (N_8669,N_1640,N_6106);
nand U8670 (N_8670,N_4536,N_6114);
nor U8671 (N_8671,N_2980,N_3819);
nor U8672 (N_8672,N_26,N_2075);
and U8673 (N_8673,N_4123,N_2096);
and U8674 (N_8674,N_1607,N_3028);
nand U8675 (N_8675,N_2181,N_933);
and U8676 (N_8676,N_1491,N_4639);
xor U8677 (N_8677,N_2914,N_420);
xor U8678 (N_8678,N_1340,N_4117);
or U8679 (N_8679,N_4826,N_5477);
and U8680 (N_8680,N_4753,N_6224);
xnor U8681 (N_8681,N_123,N_878);
and U8682 (N_8682,N_2244,N_4082);
or U8683 (N_8683,N_766,N_4541);
xnor U8684 (N_8684,N_3495,N_2074);
nor U8685 (N_8685,N_1601,N_4693);
xnor U8686 (N_8686,N_3897,N_644);
nor U8687 (N_8687,N_761,N_2453);
nor U8688 (N_8688,N_5039,N_3887);
nand U8689 (N_8689,N_2566,N_3780);
and U8690 (N_8690,N_2612,N_4930);
nand U8691 (N_8691,N_4367,N_1514);
nor U8692 (N_8692,N_1535,N_4545);
xor U8693 (N_8693,N_107,N_2143);
or U8694 (N_8694,N_884,N_2479);
nor U8695 (N_8695,N_4785,N_4510);
or U8696 (N_8696,N_3176,N_5916);
or U8697 (N_8697,N_3310,N_1685);
xor U8698 (N_8698,N_711,N_3423);
and U8699 (N_8699,N_144,N_74);
xor U8700 (N_8700,N_5734,N_2385);
or U8701 (N_8701,N_2832,N_3492);
or U8702 (N_8702,N_3827,N_1515);
or U8703 (N_8703,N_1721,N_5069);
nor U8704 (N_8704,N_2122,N_6069);
nand U8705 (N_8705,N_3001,N_5768);
or U8706 (N_8706,N_4349,N_4680);
and U8707 (N_8707,N_255,N_3514);
or U8708 (N_8708,N_5545,N_3204);
and U8709 (N_8709,N_5489,N_2508);
and U8710 (N_8710,N_2670,N_3507);
and U8711 (N_8711,N_2444,N_3657);
xor U8712 (N_8712,N_3227,N_2365);
or U8713 (N_8713,N_4054,N_3783);
xor U8714 (N_8714,N_6074,N_2967);
nor U8715 (N_8715,N_3665,N_4338);
or U8716 (N_8716,N_1729,N_2894);
or U8717 (N_8717,N_3470,N_890);
nand U8718 (N_8718,N_5277,N_3937);
and U8719 (N_8719,N_4681,N_1027);
nor U8720 (N_8720,N_963,N_5848);
nand U8721 (N_8721,N_3494,N_3543);
nor U8722 (N_8722,N_4341,N_2806);
nand U8723 (N_8723,N_4260,N_3006);
and U8724 (N_8724,N_1170,N_3525);
nand U8725 (N_8725,N_3475,N_2107);
nor U8726 (N_8726,N_967,N_4133);
nor U8727 (N_8727,N_2086,N_4528);
or U8728 (N_8728,N_4722,N_5979);
or U8729 (N_8729,N_1042,N_291);
and U8730 (N_8730,N_619,N_3335);
nor U8731 (N_8731,N_2903,N_570);
nor U8732 (N_8732,N_5292,N_4950);
and U8733 (N_8733,N_4073,N_3561);
or U8734 (N_8734,N_844,N_3640);
nor U8735 (N_8735,N_3915,N_549);
nor U8736 (N_8736,N_101,N_3433);
or U8737 (N_8737,N_4230,N_5373);
or U8738 (N_8738,N_1476,N_130);
or U8739 (N_8739,N_921,N_1628);
nand U8740 (N_8740,N_2467,N_4940);
xnor U8741 (N_8741,N_272,N_2148);
or U8742 (N_8742,N_4661,N_5346);
xor U8743 (N_8743,N_5989,N_3414);
or U8744 (N_8744,N_2100,N_120);
and U8745 (N_8745,N_1069,N_415);
nor U8746 (N_8746,N_1416,N_6196);
nand U8747 (N_8747,N_2263,N_1492);
or U8748 (N_8748,N_2392,N_3980);
or U8749 (N_8749,N_3947,N_3978);
xnor U8750 (N_8750,N_3796,N_4490);
nor U8751 (N_8751,N_5253,N_481);
xnor U8752 (N_8752,N_4885,N_181);
and U8753 (N_8753,N_1363,N_6049);
or U8754 (N_8754,N_3053,N_2902);
nand U8755 (N_8755,N_5586,N_929);
nor U8756 (N_8756,N_270,N_2771);
and U8757 (N_8757,N_3713,N_5556);
nor U8758 (N_8758,N_4739,N_1570);
and U8759 (N_8759,N_311,N_5635);
nor U8760 (N_8760,N_5344,N_6009);
nand U8761 (N_8761,N_152,N_2587);
and U8762 (N_8762,N_5316,N_1457);
or U8763 (N_8763,N_2111,N_3107);
nor U8764 (N_8764,N_959,N_3099);
or U8765 (N_8765,N_4987,N_2387);
or U8766 (N_8766,N_3242,N_4160);
nand U8767 (N_8767,N_961,N_3261);
or U8768 (N_8768,N_5175,N_3019);
or U8769 (N_8769,N_2123,N_5142);
nor U8770 (N_8770,N_5982,N_3984);
nand U8771 (N_8771,N_1423,N_2642);
or U8772 (N_8772,N_5258,N_85);
or U8773 (N_8773,N_3816,N_45);
or U8774 (N_8774,N_5227,N_1227);
nand U8775 (N_8775,N_392,N_5850);
and U8776 (N_8776,N_1947,N_4547);
and U8777 (N_8777,N_5481,N_2714);
nand U8778 (N_8778,N_3217,N_4146);
nor U8779 (N_8779,N_3573,N_1422);
nor U8780 (N_8780,N_3972,N_4155);
nand U8781 (N_8781,N_1073,N_4);
xor U8782 (N_8782,N_3948,N_1823);
or U8783 (N_8783,N_5795,N_1569);
nand U8784 (N_8784,N_5839,N_2919);
or U8785 (N_8785,N_2597,N_4259);
nand U8786 (N_8786,N_5595,N_4330);
nor U8787 (N_8787,N_5138,N_218);
nor U8788 (N_8788,N_6038,N_4754);
nor U8789 (N_8789,N_1316,N_3452);
nand U8790 (N_8790,N_1035,N_256);
nor U8791 (N_8791,N_2830,N_21);
nor U8792 (N_8792,N_5978,N_3602);
and U8793 (N_8793,N_1777,N_4844);
nor U8794 (N_8794,N_2407,N_6056);
or U8795 (N_8795,N_5565,N_5475);
or U8796 (N_8796,N_1031,N_4427);
and U8797 (N_8797,N_2028,N_469);
nand U8798 (N_8798,N_3751,N_3100);
and U8799 (N_8799,N_2641,N_812);
nor U8800 (N_8800,N_2946,N_2298);
and U8801 (N_8801,N_1748,N_2286);
nand U8802 (N_8802,N_135,N_656);
nor U8803 (N_8803,N_4455,N_5317);
or U8804 (N_8804,N_106,N_2285);
nand U8805 (N_8805,N_4667,N_2613);
nor U8806 (N_8806,N_731,N_440);
nor U8807 (N_8807,N_575,N_2483);
and U8808 (N_8808,N_1182,N_6030);
nand U8809 (N_8809,N_4918,N_2955);
or U8810 (N_8810,N_5108,N_5143);
nor U8811 (N_8811,N_3790,N_3385);
nor U8812 (N_8812,N_5136,N_5987);
nand U8813 (N_8813,N_1904,N_4618);
or U8814 (N_8814,N_4300,N_166);
nand U8815 (N_8815,N_3268,N_4625);
nor U8816 (N_8816,N_2515,N_2412);
nand U8817 (N_8817,N_148,N_5920);
nand U8818 (N_8818,N_183,N_3422);
and U8819 (N_8819,N_5581,N_5932);
nor U8820 (N_8820,N_3345,N_1320);
nand U8821 (N_8821,N_4575,N_3089);
xnor U8822 (N_8822,N_459,N_5830);
nor U8823 (N_8823,N_1805,N_3795);
nand U8824 (N_8824,N_4561,N_960);
xnor U8825 (N_8825,N_3375,N_2809);
and U8826 (N_8826,N_6026,N_3085);
or U8827 (N_8827,N_2873,N_2324);
nor U8828 (N_8828,N_2991,N_779);
nand U8829 (N_8829,N_2704,N_4670);
nand U8830 (N_8830,N_3195,N_336);
and U8831 (N_8831,N_5660,N_1975);
or U8832 (N_8832,N_6118,N_1005);
nand U8833 (N_8833,N_4395,N_3806);
nor U8834 (N_8834,N_1431,N_2433);
or U8835 (N_8835,N_231,N_1455);
nand U8836 (N_8836,N_1044,N_6071);
and U8837 (N_8837,N_650,N_5106);
xnor U8838 (N_8838,N_815,N_2653);
nand U8839 (N_8839,N_5826,N_591);
or U8840 (N_8840,N_1156,N_6236);
and U8841 (N_8841,N_4990,N_4581);
or U8842 (N_8842,N_355,N_3835);
and U8843 (N_8843,N_1037,N_4852);
xnor U8844 (N_8844,N_2034,N_2076);
and U8845 (N_8845,N_531,N_5996);
and U8846 (N_8846,N_708,N_3231);
and U8847 (N_8847,N_187,N_5425);
nand U8848 (N_8848,N_5448,N_3055);
and U8849 (N_8849,N_1612,N_3281);
nand U8850 (N_8850,N_2645,N_1000);
and U8851 (N_8851,N_2533,N_3598);
and U8852 (N_8852,N_5862,N_6025);
xor U8853 (N_8853,N_1618,N_5603);
nor U8854 (N_8854,N_5454,N_1300);
and U8855 (N_8855,N_4055,N_1602);
and U8856 (N_8856,N_5093,N_1854);
xor U8857 (N_8857,N_6011,N_5577);
and U8858 (N_8858,N_156,N_2311);
or U8859 (N_8859,N_4063,N_5936);
and U8860 (N_8860,N_4208,N_726);
or U8861 (N_8861,N_847,N_4582);
and U8862 (N_8862,N_4496,N_4336);
xor U8863 (N_8863,N_3200,N_5670);
nor U8864 (N_8864,N_4698,N_1529);
or U8865 (N_8865,N_3357,N_4411);
nand U8866 (N_8866,N_5403,N_5822);
nor U8867 (N_8867,N_2302,N_3461);
xnor U8868 (N_8868,N_2322,N_5450);
and U8869 (N_8869,N_790,N_4304);
and U8870 (N_8870,N_2617,N_2466);
nand U8871 (N_8871,N_909,N_4772);
or U8872 (N_8872,N_3923,N_971);
nand U8873 (N_8873,N_2391,N_5696);
nor U8874 (N_8874,N_487,N_4665);
nor U8875 (N_8875,N_2027,N_4612);
xnor U8876 (N_8876,N_4216,N_3920);
xor U8877 (N_8877,N_1964,N_3973);
nor U8878 (N_8878,N_1929,N_383);
and U8879 (N_8879,N_398,N_2722);
nor U8880 (N_8880,N_5495,N_234);
xnor U8881 (N_8881,N_3356,N_5050);
and U8882 (N_8882,N_922,N_2088);
xnor U8883 (N_8883,N_3364,N_5836);
nor U8884 (N_8884,N_4619,N_4203);
nor U8885 (N_8885,N_5699,N_583);
nand U8886 (N_8886,N_1878,N_5309);
or U8887 (N_8887,N_6155,N_1844);
and U8888 (N_8888,N_2863,N_1871);
nand U8889 (N_8889,N_2188,N_1246);
or U8890 (N_8890,N_1624,N_2847);
and U8891 (N_8891,N_3294,N_1176);
nand U8892 (N_8892,N_3538,N_48);
and U8893 (N_8893,N_777,N_405);
nor U8894 (N_8894,N_1477,N_4331);
nor U8895 (N_8895,N_6047,N_4771);
nand U8896 (N_8896,N_4870,N_4421);
or U8897 (N_8897,N_6003,N_5784);
or U8898 (N_8898,N_2247,N_5870);
and U8899 (N_8899,N_5761,N_716);
nand U8900 (N_8900,N_5823,N_1311);
xnor U8901 (N_8901,N_4441,N_1324);
nand U8902 (N_8902,N_2790,N_1792);
xor U8903 (N_8903,N_1989,N_683);
or U8904 (N_8904,N_2273,N_6042);
nand U8905 (N_8905,N_5058,N_2829);
xnor U8906 (N_8906,N_4477,N_2171);
nor U8907 (N_8907,N_4999,N_1608);
xor U8908 (N_8908,N_5684,N_3663);
xnor U8909 (N_8909,N_1928,N_949);
nand U8910 (N_8910,N_1443,N_5510);
and U8911 (N_8911,N_5520,N_1144);
xor U8912 (N_8912,N_3193,N_1212);
and U8913 (N_8913,N_1478,N_4140);
or U8914 (N_8914,N_1572,N_1408);
nand U8915 (N_8915,N_5973,N_5643);
nor U8916 (N_8916,N_3329,N_382);
or U8917 (N_8917,N_2161,N_2198);
or U8918 (N_8918,N_1834,N_830);
nor U8919 (N_8919,N_3771,N_694);
nand U8920 (N_8920,N_62,N_5449);
or U8921 (N_8921,N_5267,N_4526);
or U8922 (N_8922,N_4572,N_1876);
xor U8923 (N_8923,N_4973,N_2719);
nor U8924 (N_8924,N_149,N_1061);
nand U8925 (N_8925,N_5550,N_2013);
or U8926 (N_8926,N_496,N_4175);
and U8927 (N_8927,N_5988,N_116);
xnor U8928 (N_8928,N_2691,N_2697);
xor U8929 (N_8929,N_1998,N_343);
xnor U8930 (N_8930,N_817,N_3575);
nand U8931 (N_8931,N_5,N_5682);
nor U8932 (N_8932,N_3788,N_3466);
nor U8933 (N_8933,N_1886,N_171);
and U8934 (N_8934,N_1718,N_730);
nand U8935 (N_8935,N_3233,N_6156);
and U8936 (N_8936,N_5677,N_2509);
and U8937 (N_8937,N_5029,N_2872);
xnor U8938 (N_8938,N_2282,N_1106);
nor U8939 (N_8939,N_1861,N_4777);
or U8940 (N_8940,N_3848,N_2425);
and U8941 (N_8941,N_4562,N_3398);
nand U8942 (N_8942,N_5274,N_2876);
nand U8943 (N_8943,N_3039,N_3151);
nor U8944 (N_8944,N_3371,N_3020);
xnor U8945 (N_8945,N_6119,N_3963);
nor U8946 (N_8946,N_5593,N_663);
xor U8947 (N_8947,N_4264,N_3741);
xnor U8948 (N_8948,N_3921,N_3617);
and U8949 (N_8949,N_4637,N_2002);
or U8950 (N_8950,N_3218,N_1409);
or U8951 (N_8951,N_3871,N_6211);
xnor U8952 (N_8952,N_6187,N_659);
nor U8953 (N_8953,N_2006,N_4355);
or U8954 (N_8954,N_5170,N_4058);
xor U8955 (N_8955,N_2223,N_2421);
nand U8956 (N_8956,N_2317,N_378);
nor U8957 (N_8957,N_1224,N_1568);
or U8958 (N_8958,N_177,N_5854);
and U8959 (N_8959,N_4375,N_5941);
xor U8960 (N_8960,N_2432,N_3508);
nor U8961 (N_8961,N_2315,N_4347);
xnor U8962 (N_8962,N_4222,N_3782);
or U8963 (N_8963,N_4713,N_3558);
and U8964 (N_8964,N_1093,N_4880);
nor U8965 (N_8965,N_5606,N_1846);
or U8966 (N_8966,N_4994,N_1278);
or U8967 (N_8967,N_4454,N_2321);
nand U8968 (N_8968,N_5250,N_5842);
nor U8969 (N_8969,N_6139,N_1158);
nand U8970 (N_8970,N_194,N_5869);
nor U8971 (N_8971,N_3181,N_6127);
nand U8972 (N_8972,N_159,N_3145);
or U8973 (N_8973,N_5937,N_3832);
or U8974 (N_8974,N_4173,N_1950);
nor U8975 (N_8975,N_2937,N_5605);
and U8976 (N_8976,N_2039,N_5630);
nand U8977 (N_8977,N_302,N_55);
or U8978 (N_8978,N_3745,N_2969);
xor U8979 (N_8979,N_3752,N_4674);
or U8980 (N_8980,N_880,N_6058);
or U8981 (N_8981,N_4478,N_140);
xnor U8982 (N_8982,N_825,N_1908);
and U8983 (N_8983,N_4251,N_1867);
or U8984 (N_8984,N_2690,N_4377);
nand U8985 (N_8985,N_2436,N_4982);
and U8986 (N_8986,N_5447,N_2660);
nand U8987 (N_8987,N_1750,N_2461);
or U8988 (N_8988,N_4615,N_1152);
and U8989 (N_8989,N_3889,N_3010);
nand U8990 (N_8990,N_5974,N_1230);
and U8991 (N_8991,N_5047,N_2908);
xnor U8992 (N_8992,N_976,N_3859);
and U8993 (N_8993,N_1597,N_4820);
and U8994 (N_8994,N_2375,N_3720);
nand U8995 (N_8995,N_6174,N_4480);
and U8996 (N_8996,N_5817,N_1134);
and U8997 (N_8997,N_3185,N_3284);
or U8998 (N_8998,N_3696,N_5082);
or U8999 (N_8999,N_1550,N_2935);
xnor U9000 (N_9000,N_3942,N_3465);
and U9001 (N_9001,N_2085,N_5629);
nand U9002 (N_9002,N_3177,N_5282);
xor U9003 (N_9003,N_3254,N_4876);
or U9004 (N_9004,N_5923,N_4635);
or U9005 (N_9005,N_1374,N_3877);
nand U9006 (N_9006,N_3747,N_5393);
and U9007 (N_9007,N_3768,N_1829);
nor U9008 (N_9008,N_555,N_1705);
and U9009 (N_9009,N_4469,N_6050);
xor U9010 (N_9010,N_4220,N_1013);
and U9011 (N_9011,N_3212,N_2140);
nor U9012 (N_9012,N_1049,N_789);
xor U9013 (N_9013,N_5728,N_5166);
nor U9014 (N_9014,N_1884,N_5859);
xor U9015 (N_9015,N_5617,N_1764);
nor U9016 (N_9016,N_2999,N_3682);
nor U9017 (N_9017,N_362,N_1473);
nand U9018 (N_9018,N_2538,N_3347);
nand U9019 (N_9019,N_5533,N_4953);
and U9020 (N_9020,N_4576,N_3565);
or U9021 (N_9021,N_2769,N_4307);
and U9022 (N_9022,N_1735,N_1041);
nor U9023 (N_9023,N_2703,N_4821);
and U9024 (N_9024,N_463,N_1648);
or U9025 (N_9025,N_2848,N_4647);
nand U9026 (N_9026,N_834,N_3354);
xnor U9027 (N_9027,N_6031,N_3950);
and U9028 (N_9028,N_4243,N_2406);
nand U9029 (N_9029,N_1202,N_1184);
and U9030 (N_9030,N_5251,N_2031);
xnor U9031 (N_9031,N_3679,N_2098);
nand U9032 (N_9032,N_5625,N_5365);
and U9033 (N_9033,N_6198,N_6242);
xnor U9034 (N_9034,N_2675,N_5541);
and U9035 (N_9035,N_639,N_3971);
xor U9036 (N_9036,N_2800,N_137);
xor U9037 (N_9037,N_3307,N_2179);
and U9038 (N_9038,N_1336,N_98);
nand U9039 (N_9039,N_5174,N_1579);
and U9040 (N_9040,N_5704,N_992);
xnor U9041 (N_9041,N_3735,N_2029);
or U9042 (N_9042,N_2831,N_2427);
xnor U9043 (N_9043,N_1513,N_3022);
and U9044 (N_9044,N_1329,N_2204);
and U9045 (N_9045,N_3759,N_6037);
nor U9046 (N_9046,N_5918,N_93);
or U9047 (N_9047,N_2280,N_2252);
or U9048 (N_9048,N_5736,N_1978);
and U9049 (N_9049,N_4631,N_4859);
and U9050 (N_9050,N_5468,N_207);
nand U9051 (N_9051,N_161,N_2336);
xor U9052 (N_9052,N_1824,N_1474);
xor U9053 (N_9053,N_2998,N_5746);
xor U9054 (N_9054,N_3552,N_5969);
or U9055 (N_9055,N_300,N_4041);
nand U9056 (N_9056,N_1451,N_6130);
nand U9057 (N_9057,N_1203,N_4109);
and U9058 (N_9058,N_1986,N_4193);
and U9059 (N_9059,N_1636,N_2170);
nand U9060 (N_9060,N_1605,N_782);
nor U9061 (N_9061,N_4135,N_4709);
nor U9062 (N_9062,N_1481,N_2542);
xnor U9063 (N_9063,N_4257,N_1772);
nor U9064 (N_9064,N_1827,N_903);
xor U9065 (N_9065,N_349,N_2854);
xnor U9066 (N_9066,N_732,N_2291);
or U9067 (N_9067,N_254,N_5062);
or U9068 (N_9068,N_2841,N_176);
and U9069 (N_9069,N_6181,N_2338);
nor U9070 (N_9070,N_2516,N_3114);
nand U9071 (N_9071,N_2731,N_2664);
xor U9072 (N_9072,N_771,N_6116);
nand U9073 (N_9073,N_3070,N_2097);
xnor U9074 (N_9074,N_3175,N_870);
nor U9075 (N_9075,N_2624,N_3739);
nor U9076 (N_9076,N_4424,N_2372);
nor U9077 (N_9077,N_6045,N_1934);
nor U9078 (N_9078,N_4796,N_5223);
xnor U9079 (N_9079,N_1411,N_1697);
or U9080 (N_9080,N_1559,N_4232);
nor U9081 (N_9081,N_3509,N_1523);
nor U9082 (N_9082,N_5005,N_2549);
xnor U9083 (N_9083,N_5271,N_673);
xnor U9084 (N_9084,N_901,N_389);
nor U9085 (N_9085,N_5414,N_2334);
xor U9086 (N_9086,N_5190,N_5090);
nor U9087 (N_9087,N_6148,N_353);
or U9088 (N_9088,N_5527,N_2465);
and U9089 (N_9089,N_1660,N_1057);
nor U9090 (N_9090,N_5507,N_5689);
nor U9091 (N_9091,N_4278,N_3124);
nand U9092 (N_9092,N_259,N_252);
nand U9093 (N_9093,N_470,N_5939);
nor U9094 (N_9094,N_1046,N_3350);
xnor U9095 (N_9095,N_764,N_4965);
xnor U9096 (N_9096,N_5811,N_345);
or U9097 (N_9097,N_5897,N_813);
nand U9098 (N_9098,N_5876,N_4533);
nand U9099 (N_9099,N_5553,N_5807);
and U9100 (N_9100,N_3748,N_3764);
or U9101 (N_9101,N_1725,N_2594);
nor U9102 (N_9102,N_5353,N_1892);
nand U9103 (N_9103,N_54,N_5708);
and U9104 (N_9104,N_1670,N_5501);
and U9105 (N_9105,N_3483,N_1126);
nor U9106 (N_9106,N_2326,N_90);
nor U9107 (N_9107,N_5105,N_1439);
nand U9108 (N_9108,N_4212,N_1818);
xor U9109 (N_9109,N_287,N_2867);
and U9110 (N_9110,N_4745,N_2089);
or U9111 (N_9111,N_3692,N_6098);
xnor U9112 (N_9112,N_1259,N_2264);
nand U9113 (N_9113,N_5288,N_4139);
nor U9114 (N_9114,N_2813,N_4941);
xnor U9115 (N_9115,N_306,N_6182);
nand U9116 (N_9116,N_544,N_4806);
xor U9117 (N_9117,N_4922,N_1631);
or U9118 (N_9118,N_3635,N_1936);
xnor U9119 (N_9119,N_2158,N_2513);
nor U9120 (N_9120,N_4303,N_4759);
or U9121 (N_9121,N_4204,N_829);
nor U9122 (N_9122,N_3063,N_1141);
nor U9123 (N_9123,N_5164,N_4617);
xor U9124 (N_9124,N_418,N_2215);
nand U9125 (N_9125,N_1650,N_1274);
xor U9126 (N_9126,N_4418,N_4291);
and U9127 (N_9127,N_524,N_1563);
or U9128 (N_9128,N_3612,N_3462);
or U9129 (N_9129,N_49,N_3882);
xnor U9130 (N_9130,N_629,N_5915);
xnor U9131 (N_9131,N_1702,N_4277);
nand U9132 (N_9132,N_1094,N_5036);
nand U9133 (N_9133,N_4906,N_2681);
nor U9134 (N_9134,N_1444,N_3326);
nand U9135 (N_9135,N_4077,N_426);
nand U9136 (N_9136,N_2585,N_5061);
and U9137 (N_9137,N_3866,N_482);
xnor U9138 (N_9138,N_4060,N_4044);
and U9139 (N_9139,N_3139,N_5911);
xor U9140 (N_9140,N_4968,N_574);
xor U9141 (N_9141,N_4817,N_5343);
xor U9142 (N_9142,N_5225,N_129);
and U9143 (N_9143,N_4630,N_5983);
xnor U9144 (N_9144,N_3890,N_837);
and U9145 (N_9145,N_5123,N_1715);
nand U9146 (N_9146,N_4470,N_5323);
nor U9147 (N_9147,N_6212,N_5161);
xor U9148 (N_9148,N_3163,N_3134);
xnor U9149 (N_9149,N_3645,N_5265);
xor U9150 (N_9150,N_1286,N_5847);
nor U9151 (N_9151,N_3071,N_701);
or U9152 (N_9152,N_2672,N_3116);
or U9153 (N_9153,N_1466,N_5089);
or U9154 (N_9154,N_1958,N_2134);
nand U9155 (N_9155,N_5904,N_4687);
and U9156 (N_9156,N_5966,N_118);
or U9157 (N_9157,N_3527,N_3940);
nor U9158 (N_9158,N_4067,N_3758);
and U9159 (N_9159,N_2383,N_4380);
xnor U9160 (N_9160,N_4402,N_3049);
or U9161 (N_9161,N_952,N_4248);
or U9162 (N_9162,N_2694,N_4244);
xor U9163 (N_9163,N_2296,N_4428);
nor U9164 (N_9164,N_1222,N_1275);
nor U9165 (N_9165,N_5406,N_5466);
and U9166 (N_9166,N_5673,N_3045);
and U9167 (N_9167,N_3862,N_2808);
nand U9168 (N_9168,N_4134,N_3066);
nor U9169 (N_9169,N_2119,N_1192);
nand U9170 (N_9170,N_2833,N_6076);
xnor U9171 (N_9171,N_4849,N_1968);
and U9172 (N_9172,N_5494,N_2947);
nor U9173 (N_9173,N_4963,N_5934);
nand U9174 (N_9174,N_616,N_6157);
or U9175 (N_9175,N_3638,N_5361);
nor U9176 (N_9176,N_3953,N_827);
and U9177 (N_9177,N_4113,N_3753);
or U9178 (N_9178,N_4399,N_1304);
nor U9179 (N_9179,N_3512,N_189);
nand U9180 (N_9180,N_2825,N_1589);
and U9181 (N_9181,N_346,N_257);
and U9182 (N_9182,N_597,N_3438);
xnor U9183 (N_9183,N_2216,N_4107);
nand U9184 (N_9184,N_1757,N_704);
nor U9185 (N_9185,N_330,N_3925);
nor U9186 (N_9186,N_2117,N_4169);
xnor U9187 (N_9187,N_5204,N_296);
or U9188 (N_9188,N_3497,N_3533);
or U9189 (N_9189,N_1086,N_537);
nor U9190 (N_9190,N_443,N_6070);
xor U9191 (N_9191,N_5369,N_3372);
xnor U9192 (N_9192,N_916,N_1528);
and U9193 (N_9193,N_1610,N_4014);
xor U9194 (N_9194,N_5986,N_3709);
xnor U9195 (N_9195,N_5558,N_1625);
xnor U9196 (N_9196,N_3911,N_938);
xor U9197 (N_9197,N_430,N_2528);
nor U9198 (N_9198,N_2362,N_1673);
or U9199 (N_9199,N_2927,N_4289);
xnor U9200 (N_9200,N_5804,N_3439);
and U9201 (N_9201,N_3251,N_2030);
or U9202 (N_9202,N_1666,N_3767);
xor U9203 (N_9203,N_2647,N_4126);
and U9204 (N_9204,N_5329,N_6143);
and U9205 (N_9205,N_4150,N_2173);
nor U9206 (N_9206,N_3030,N_68);
and U9207 (N_9207,N_2405,N_2064);
nor U9208 (N_9208,N_6015,N_4842);
or U9209 (N_9209,N_4403,N_709);
nand U9210 (N_9210,N_2553,N_184);
or U9211 (N_9211,N_1510,N_2828);
xor U9212 (N_9212,N_5759,N_2680);
xnor U9213 (N_9213,N_5483,N_4890);
and U9214 (N_9214,N_1616,N_6142);
xor U9215 (N_9215,N_548,N_365);
xor U9216 (N_9216,N_2723,N_2618);
nor U9217 (N_9217,N_6192,N_2541);
nor U9218 (N_9218,N_1912,N_399);
nand U9219 (N_9219,N_6125,N_1874);
or U9220 (N_9220,N_3015,N_3262);
xor U9221 (N_9221,N_2713,N_3702);
or U9222 (N_9222,N_163,N_3608);
xor U9223 (N_9223,N_4903,N_4351);
nand U9224 (N_9224,N_1826,N_3804);
or U9225 (N_9225,N_4970,N_6136);
nor U9226 (N_9226,N_4708,N_2348);
xnor U9227 (N_9227,N_3956,N_2447);
nand U9228 (N_9228,N_5634,N_6099);
or U9229 (N_9229,N_1276,N_462);
and U9230 (N_9230,N_5884,N_17);
and U9231 (N_9231,N_5994,N_141);
and U9232 (N_9232,N_3111,N_3321);
nor U9233 (N_9233,N_6129,N_3348);
nand U9234 (N_9234,N_2573,N_5590);
xor U9235 (N_9235,N_5351,N_1254);
xnor U9236 (N_9236,N_485,N_3619);
nor U9237 (N_9237,N_1193,N_2659);
and U9238 (N_9238,N_3121,N_5320);
and U9239 (N_9239,N_3888,N_4816);
xor U9240 (N_9240,N_4394,N_6088);
nand U9241 (N_9241,N_2801,N_4911);
nor U9242 (N_9242,N_1261,N_2261);
xor U9243 (N_9243,N_1085,N_2305);
nor U9244 (N_9244,N_4233,N_4952);
xor U9245 (N_9245,N_686,N_6232);
nand U9246 (N_9246,N_6166,N_3415);
nor U9247 (N_9247,N_4696,N_2303);
nand U9248 (N_9248,N_2648,N_2229);
and U9249 (N_9249,N_3232,N_1179);
nor U9250 (N_9250,N_2943,N_2084);
nand U9251 (N_9251,N_3544,N_2079);
nand U9252 (N_9252,N_464,N_4136);
nor U9253 (N_9253,N_5389,N_593);
nor U9254 (N_9254,N_20,N_2152);
xor U9255 (N_9255,N_1889,N_3968);
nand U9256 (N_9256,N_4751,N_4831);
or U9257 (N_9257,N_2871,N_3498);
nor U9258 (N_9258,N_5079,N_5883);
nand U9259 (N_9259,N_5158,N_1710);
nor U9260 (N_9260,N_3808,N_1633);
nand U9261 (N_9261,N_4104,N_6022);
nand U9262 (N_9262,N_1560,N_3792);
or U9263 (N_9263,N_4324,N_168);
nor U9264 (N_9264,N_5762,N_5713);
nor U9265 (N_9265,N_3746,N_5985);
nor U9266 (N_9266,N_4090,N_1225);
and U9267 (N_9267,N_1105,N_4030);
nor U9268 (N_9268,N_1400,N_3876);
and U9269 (N_9269,N_1355,N_1903);
xor U9270 (N_9270,N_1615,N_1795);
nand U9271 (N_9271,N_4075,N_5159);
xor U9272 (N_9272,N_4207,N_758);
and U9273 (N_9273,N_1247,N_1362);
nor U9274 (N_9274,N_1419,N_1003);
and U9275 (N_9275,N_5718,N_4437);
and U9276 (N_9276,N_3884,N_5779);
or U9277 (N_9277,N_5117,N_198);
and U9278 (N_9278,N_1178,N_514);
nor U9279 (N_9279,N_749,N_3760);
nand U9280 (N_9280,N_3125,N_988);
or U9281 (N_9281,N_3891,N_3428);
or U9282 (N_9282,N_5133,N_1471);
nand U9283 (N_9283,N_4327,N_1381);
or U9284 (N_9284,N_4066,N_6123);
and U9285 (N_9285,N_1661,N_2893);
or U9286 (N_9286,N_6,N_2381);
nand U9287 (N_9287,N_729,N_3642);
xnor U9288 (N_9288,N_5094,N_5968);
xnor U9289 (N_9289,N_512,N_751);
nand U9290 (N_9290,N_5186,N_2442);
nand U9291 (N_9291,N_2586,N_5810);
or U9292 (N_9292,N_3532,N_3237);
xor U9293 (N_9293,N_182,N_6158);
or U9294 (N_9294,N_4076,N_2949);
nor U9295 (N_9295,N_3592,N_235);
or U9296 (N_9296,N_1180,N_2281);
or U9297 (N_9297,N_5234,N_3119);
xor U9298 (N_9298,N_4873,N_973);
or U9299 (N_9299,N_506,N_6177);
or U9300 (N_9300,N_669,N_4716);
nand U9301 (N_9301,N_3674,N_5216);
and U9302 (N_9302,N_2785,N_2909);
nor U9303 (N_9303,N_5878,N_6161);
nor U9304 (N_9304,N_4969,N_1081);
or U9305 (N_9305,N_5997,N_37);
xor U9306 (N_9306,N_5183,N_1130);
xor U9307 (N_9307,N_339,N_1233);
or U9308 (N_9308,N_65,N_490);
xor U9309 (N_9309,N_2701,N_2602);
nor U9310 (N_9310,N_2667,N_3976);
xnor U9311 (N_9311,N_5894,N_3966);
nor U9312 (N_9312,N_6134,N_5571);
nand U9313 (N_9313,N_975,N_5255);
or U9314 (N_9314,N_3656,N_5919);
xor U9315 (N_9315,N_6183,N_3363);
or U9316 (N_9316,N_3128,N_2207);
or U9317 (N_9317,N_1243,N_1717);
or U9318 (N_9318,N_3209,N_258);
nand U9319 (N_9319,N_3629,N_86);
or U9320 (N_9320,N_1803,N_2734);
and U9321 (N_9321,N_587,N_5328);
or U9322 (N_9322,N_1211,N_3068);
xnor U9323 (N_9323,N_4909,N_5476);
and U9324 (N_9324,N_4296,N_2599);
nand U9325 (N_9325,N_930,N_3734);
and U9326 (N_9326,N_3493,N_1071);
xor U9327 (N_9327,N_3624,N_6044);
or U9328 (N_9328,N_1561,N_1030);
or U9329 (N_9329,N_1218,N_594);
and U9330 (N_9330,N_565,N_2455);
and U9331 (N_9331,N_5280,N_1716);
nor U9332 (N_9332,N_3566,N_3990);
or U9333 (N_9333,N_1220,N_4027);
or U9334 (N_9334,N_5735,N_2607);
nand U9335 (N_9335,N_912,N_71);
or U9336 (N_9336,N_2309,N_5104);
nor U9337 (N_9337,N_2137,N_2112);
nor U9338 (N_9338,N_2977,N_4518);
nand U9339 (N_9339,N_5135,N_5355);
xor U9340 (N_9340,N_6179,N_1872);
or U9341 (N_9341,N_4715,N_4822);
nor U9342 (N_9342,N_1578,N_4805);
nand U9343 (N_9343,N_5521,N_3618);
or U9344 (N_9344,N_5844,N_1);
nand U9345 (N_9345,N_3271,N_2240);
nor U9346 (N_9346,N_374,N_3567);
xnor U9347 (N_9347,N_5116,N_585);
and U9348 (N_9348,N_955,N_3863);
and U9349 (N_9349,N_2279,N_3434);
nor U9350 (N_9350,N_563,N_5145);
nor U9351 (N_9351,N_61,N_4017);
xor U9352 (N_9352,N_5102,N_4824);
xor U9353 (N_9353,N_5013,N_4894);
nor U9354 (N_9354,N_5958,N_4508);
nand U9355 (N_9355,N_2094,N_2656);
and U9356 (N_9356,N_3550,N_2843);
nor U9357 (N_9357,N_5006,N_4218);
xnor U9358 (N_9358,N_2711,N_1200);
or U9359 (N_9359,N_4595,N_5438);
and U9360 (N_9360,N_4223,N_42);
or U9361 (N_9361,N_2886,N_4979);
nand U9362 (N_9362,N_3007,N_2191);
xnor U9363 (N_9363,N_2855,N_6054);
nand U9364 (N_9364,N_4543,N_4087);
nor U9365 (N_9365,N_3081,N_3736);
xnor U9366 (N_9366,N_3954,N_3754);
nand U9367 (N_9367,N_1556,N_5887);
and U9368 (N_9368,N_292,N_5042);
nor U9369 (N_9369,N_4783,N_185);
nand U9370 (N_9370,N_3191,N_3027);
xor U9371 (N_9371,N_5273,N_1961);
or U9372 (N_9372,N_5300,N_1191);
and U9373 (N_9373,N_1197,N_950);
and U9374 (N_9374,N_4102,N_5926);
or U9375 (N_9375,N_343,N_3872);
nor U9376 (N_9376,N_1386,N_2405);
or U9377 (N_9377,N_1939,N_5200);
xor U9378 (N_9378,N_4377,N_5749);
xor U9379 (N_9379,N_280,N_3417);
and U9380 (N_9380,N_4631,N_3189);
and U9381 (N_9381,N_4460,N_765);
or U9382 (N_9382,N_1452,N_5694);
xor U9383 (N_9383,N_2029,N_2598);
and U9384 (N_9384,N_1934,N_1572);
or U9385 (N_9385,N_52,N_5747);
nor U9386 (N_9386,N_4109,N_2018);
nor U9387 (N_9387,N_2475,N_4147);
nor U9388 (N_9388,N_5180,N_3954);
and U9389 (N_9389,N_1361,N_2138);
nor U9390 (N_9390,N_3389,N_3154);
nor U9391 (N_9391,N_891,N_5246);
nor U9392 (N_9392,N_5656,N_3066);
and U9393 (N_9393,N_2074,N_5002);
nor U9394 (N_9394,N_3073,N_5582);
or U9395 (N_9395,N_507,N_5836);
nor U9396 (N_9396,N_4686,N_2944);
or U9397 (N_9397,N_5278,N_5376);
nor U9398 (N_9398,N_1918,N_50);
nand U9399 (N_9399,N_5554,N_2223);
xnor U9400 (N_9400,N_44,N_2819);
or U9401 (N_9401,N_805,N_5039);
or U9402 (N_9402,N_5197,N_4840);
and U9403 (N_9403,N_3017,N_4945);
nand U9404 (N_9404,N_260,N_4552);
or U9405 (N_9405,N_1966,N_5639);
nor U9406 (N_9406,N_3146,N_1221);
and U9407 (N_9407,N_2061,N_813);
xnor U9408 (N_9408,N_5363,N_3846);
nor U9409 (N_9409,N_2095,N_4335);
nand U9410 (N_9410,N_81,N_5560);
nor U9411 (N_9411,N_5984,N_5427);
or U9412 (N_9412,N_4178,N_3413);
and U9413 (N_9413,N_2823,N_2115);
nand U9414 (N_9414,N_3710,N_1769);
nor U9415 (N_9415,N_5360,N_258);
or U9416 (N_9416,N_5056,N_3607);
or U9417 (N_9417,N_4840,N_3141);
or U9418 (N_9418,N_2356,N_621);
or U9419 (N_9419,N_1900,N_597);
nand U9420 (N_9420,N_5802,N_5033);
nor U9421 (N_9421,N_1016,N_5107);
nand U9422 (N_9422,N_2412,N_2756);
nand U9423 (N_9423,N_2380,N_2741);
nor U9424 (N_9424,N_1481,N_4636);
nor U9425 (N_9425,N_1612,N_2453);
and U9426 (N_9426,N_3391,N_3694);
xor U9427 (N_9427,N_4454,N_216);
nand U9428 (N_9428,N_3663,N_4004);
or U9429 (N_9429,N_1604,N_669);
and U9430 (N_9430,N_3789,N_5645);
nor U9431 (N_9431,N_5938,N_5130);
nand U9432 (N_9432,N_1695,N_4228);
nand U9433 (N_9433,N_126,N_3716);
nor U9434 (N_9434,N_1341,N_3328);
nor U9435 (N_9435,N_2235,N_3432);
or U9436 (N_9436,N_348,N_3624);
nor U9437 (N_9437,N_1109,N_2991);
xnor U9438 (N_9438,N_2214,N_4494);
nor U9439 (N_9439,N_4172,N_113);
nand U9440 (N_9440,N_4856,N_5657);
xor U9441 (N_9441,N_4321,N_1862);
nand U9442 (N_9442,N_1266,N_641);
xnor U9443 (N_9443,N_3949,N_4261);
nand U9444 (N_9444,N_2470,N_2744);
nor U9445 (N_9445,N_512,N_2684);
nor U9446 (N_9446,N_3746,N_3128);
nor U9447 (N_9447,N_3161,N_144);
nor U9448 (N_9448,N_4025,N_5852);
nand U9449 (N_9449,N_2172,N_4564);
or U9450 (N_9450,N_229,N_1670);
nor U9451 (N_9451,N_1425,N_5872);
xnor U9452 (N_9452,N_2174,N_4496);
nand U9453 (N_9453,N_5358,N_5112);
and U9454 (N_9454,N_2348,N_6153);
xnor U9455 (N_9455,N_116,N_4617);
xnor U9456 (N_9456,N_4686,N_303);
xor U9457 (N_9457,N_3240,N_5363);
nand U9458 (N_9458,N_3202,N_3119);
xnor U9459 (N_9459,N_85,N_2888);
nand U9460 (N_9460,N_5168,N_213);
or U9461 (N_9461,N_1964,N_2350);
or U9462 (N_9462,N_4273,N_2852);
nand U9463 (N_9463,N_5395,N_3399);
or U9464 (N_9464,N_2447,N_3552);
and U9465 (N_9465,N_2897,N_1499);
or U9466 (N_9466,N_3038,N_616);
nand U9467 (N_9467,N_5448,N_3925);
nor U9468 (N_9468,N_6128,N_1692);
xor U9469 (N_9469,N_3630,N_5313);
or U9470 (N_9470,N_3429,N_2946);
nor U9471 (N_9471,N_3105,N_4862);
and U9472 (N_9472,N_2561,N_282);
nor U9473 (N_9473,N_1918,N_5827);
or U9474 (N_9474,N_2404,N_317);
or U9475 (N_9475,N_2977,N_1012);
nand U9476 (N_9476,N_1682,N_5595);
nand U9477 (N_9477,N_3852,N_3440);
nand U9478 (N_9478,N_5345,N_5920);
or U9479 (N_9479,N_4128,N_1704);
and U9480 (N_9480,N_3019,N_803);
xnor U9481 (N_9481,N_1981,N_1038);
nor U9482 (N_9482,N_5514,N_1846);
xor U9483 (N_9483,N_4075,N_5963);
and U9484 (N_9484,N_1601,N_5028);
nand U9485 (N_9485,N_4569,N_2669);
or U9486 (N_9486,N_5351,N_1998);
nand U9487 (N_9487,N_895,N_3112);
or U9488 (N_9488,N_4935,N_3993);
xor U9489 (N_9489,N_3574,N_202);
xor U9490 (N_9490,N_1079,N_3846);
xnor U9491 (N_9491,N_915,N_5693);
nand U9492 (N_9492,N_3449,N_4325);
or U9493 (N_9493,N_2097,N_550);
xnor U9494 (N_9494,N_5400,N_2530);
or U9495 (N_9495,N_5754,N_1373);
and U9496 (N_9496,N_586,N_657);
and U9497 (N_9497,N_1107,N_1051);
xnor U9498 (N_9498,N_2663,N_4048);
nand U9499 (N_9499,N_2695,N_4689);
xnor U9500 (N_9500,N_4437,N_5575);
or U9501 (N_9501,N_4122,N_5035);
and U9502 (N_9502,N_5578,N_3569);
or U9503 (N_9503,N_2742,N_4197);
nand U9504 (N_9504,N_5927,N_5591);
and U9505 (N_9505,N_4628,N_4800);
and U9506 (N_9506,N_2547,N_3285);
nand U9507 (N_9507,N_52,N_2631);
nor U9508 (N_9508,N_3574,N_2985);
and U9509 (N_9509,N_1110,N_3651);
and U9510 (N_9510,N_1413,N_1173);
nor U9511 (N_9511,N_1778,N_895);
or U9512 (N_9512,N_5623,N_5194);
nand U9513 (N_9513,N_4644,N_3420);
nand U9514 (N_9514,N_1091,N_4174);
nor U9515 (N_9515,N_3670,N_1435);
or U9516 (N_9516,N_5098,N_5262);
nand U9517 (N_9517,N_710,N_5113);
and U9518 (N_9518,N_3302,N_194);
nand U9519 (N_9519,N_1735,N_3951);
or U9520 (N_9520,N_1709,N_1473);
or U9521 (N_9521,N_3124,N_4081);
and U9522 (N_9522,N_5185,N_490);
or U9523 (N_9523,N_189,N_4754);
nor U9524 (N_9524,N_1809,N_5000);
nand U9525 (N_9525,N_1955,N_1841);
xnor U9526 (N_9526,N_727,N_3271);
nor U9527 (N_9527,N_1311,N_74);
or U9528 (N_9528,N_5325,N_5827);
and U9529 (N_9529,N_4664,N_3870);
or U9530 (N_9530,N_2220,N_93);
or U9531 (N_9531,N_1845,N_6005);
nor U9532 (N_9532,N_3064,N_3884);
or U9533 (N_9533,N_4291,N_3744);
xnor U9534 (N_9534,N_5552,N_2840);
xor U9535 (N_9535,N_3359,N_2319);
xnor U9536 (N_9536,N_3559,N_3046);
nand U9537 (N_9537,N_479,N_4968);
nor U9538 (N_9538,N_4287,N_4787);
xnor U9539 (N_9539,N_3907,N_3703);
and U9540 (N_9540,N_4985,N_3369);
or U9541 (N_9541,N_2876,N_5706);
nor U9542 (N_9542,N_2999,N_4420);
nor U9543 (N_9543,N_2676,N_6211);
xor U9544 (N_9544,N_251,N_2284);
or U9545 (N_9545,N_5895,N_1162);
nor U9546 (N_9546,N_4198,N_1056);
nor U9547 (N_9547,N_4596,N_4552);
nand U9548 (N_9548,N_4060,N_4225);
nor U9549 (N_9549,N_3173,N_317);
and U9550 (N_9550,N_3844,N_6168);
or U9551 (N_9551,N_2765,N_4707);
or U9552 (N_9552,N_4932,N_5066);
nand U9553 (N_9553,N_534,N_4534);
nand U9554 (N_9554,N_635,N_4228);
and U9555 (N_9555,N_1764,N_361);
or U9556 (N_9556,N_2631,N_4300);
or U9557 (N_9557,N_1466,N_1075);
nor U9558 (N_9558,N_2809,N_6038);
nor U9559 (N_9559,N_4818,N_2896);
or U9560 (N_9560,N_4684,N_4589);
and U9561 (N_9561,N_4176,N_2710);
and U9562 (N_9562,N_4118,N_1820);
nand U9563 (N_9563,N_1195,N_2162);
or U9564 (N_9564,N_4350,N_3952);
xnor U9565 (N_9565,N_1061,N_3596);
nor U9566 (N_9566,N_806,N_5376);
or U9567 (N_9567,N_2468,N_553);
or U9568 (N_9568,N_959,N_1803);
nand U9569 (N_9569,N_3196,N_239);
nor U9570 (N_9570,N_3140,N_4128);
xnor U9571 (N_9571,N_3261,N_1291);
nor U9572 (N_9572,N_384,N_2521);
nand U9573 (N_9573,N_2583,N_507);
or U9574 (N_9574,N_1565,N_3026);
and U9575 (N_9575,N_4478,N_4158);
and U9576 (N_9576,N_1108,N_3740);
nand U9577 (N_9577,N_2408,N_6051);
or U9578 (N_9578,N_3208,N_1685);
nor U9579 (N_9579,N_2186,N_463);
nand U9580 (N_9580,N_4631,N_2908);
nand U9581 (N_9581,N_3928,N_5459);
or U9582 (N_9582,N_5684,N_3742);
or U9583 (N_9583,N_5757,N_4779);
xor U9584 (N_9584,N_3476,N_3893);
nand U9585 (N_9585,N_3589,N_2201);
nand U9586 (N_9586,N_2875,N_4081);
nand U9587 (N_9587,N_3888,N_2004);
or U9588 (N_9588,N_5387,N_5295);
xnor U9589 (N_9589,N_3813,N_2800);
xnor U9590 (N_9590,N_4642,N_2438);
xor U9591 (N_9591,N_5349,N_808);
xor U9592 (N_9592,N_3038,N_161);
nor U9593 (N_9593,N_2106,N_2373);
xnor U9594 (N_9594,N_2958,N_2615);
and U9595 (N_9595,N_4288,N_1451);
or U9596 (N_9596,N_2014,N_4309);
nand U9597 (N_9597,N_2800,N_1387);
and U9598 (N_9598,N_1421,N_3673);
xor U9599 (N_9599,N_4938,N_3489);
nand U9600 (N_9600,N_60,N_1073);
or U9601 (N_9601,N_3393,N_2973);
nor U9602 (N_9602,N_4111,N_123);
nand U9603 (N_9603,N_39,N_2023);
nand U9604 (N_9604,N_1156,N_1712);
nand U9605 (N_9605,N_5439,N_80);
and U9606 (N_9606,N_3252,N_1268);
xnor U9607 (N_9607,N_4038,N_5009);
and U9608 (N_9608,N_1792,N_1244);
nand U9609 (N_9609,N_4338,N_262);
and U9610 (N_9610,N_6140,N_5283);
nand U9611 (N_9611,N_3026,N_3476);
nand U9612 (N_9612,N_2167,N_2647);
nor U9613 (N_9613,N_551,N_3302);
or U9614 (N_9614,N_5838,N_4390);
xor U9615 (N_9615,N_3046,N_1955);
and U9616 (N_9616,N_1348,N_6020);
nand U9617 (N_9617,N_942,N_5529);
and U9618 (N_9618,N_4555,N_2984);
nor U9619 (N_9619,N_679,N_6235);
xnor U9620 (N_9620,N_4346,N_5289);
nor U9621 (N_9621,N_6027,N_1507);
and U9622 (N_9622,N_5575,N_591);
nand U9623 (N_9623,N_4835,N_840);
nor U9624 (N_9624,N_96,N_5105);
or U9625 (N_9625,N_1373,N_829);
nor U9626 (N_9626,N_710,N_5821);
nor U9627 (N_9627,N_1518,N_613);
or U9628 (N_9628,N_4439,N_3604);
or U9629 (N_9629,N_714,N_3042);
and U9630 (N_9630,N_1891,N_3934);
nor U9631 (N_9631,N_3246,N_4873);
nor U9632 (N_9632,N_4310,N_1930);
or U9633 (N_9633,N_664,N_4210);
nand U9634 (N_9634,N_3944,N_5466);
xor U9635 (N_9635,N_5202,N_3522);
xnor U9636 (N_9636,N_886,N_760);
and U9637 (N_9637,N_5881,N_1610);
and U9638 (N_9638,N_2032,N_5476);
xor U9639 (N_9639,N_4585,N_6160);
xnor U9640 (N_9640,N_4191,N_1877);
nor U9641 (N_9641,N_4575,N_2393);
and U9642 (N_9642,N_5850,N_1594);
nand U9643 (N_9643,N_3660,N_3170);
and U9644 (N_9644,N_4947,N_3218);
nor U9645 (N_9645,N_3837,N_561);
nor U9646 (N_9646,N_3046,N_1638);
xor U9647 (N_9647,N_5612,N_3049);
nor U9648 (N_9648,N_982,N_4804);
and U9649 (N_9649,N_1869,N_5328);
xor U9650 (N_9650,N_5028,N_1090);
nand U9651 (N_9651,N_3030,N_1410);
and U9652 (N_9652,N_306,N_5381);
nand U9653 (N_9653,N_5371,N_5062);
and U9654 (N_9654,N_3092,N_2615);
and U9655 (N_9655,N_4773,N_115);
nor U9656 (N_9656,N_665,N_5129);
and U9657 (N_9657,N_5984,N_5484);
nor U9658 (N_9658,N_6197,N_5985);
nor U9659 (N_9659,N_2035,N_2527);
nor U9660 (N_9660,N_1457,N_5255);
or U9661 (N_9661,N_3939,N_2846);
xor U9662 (N_9662,N_2963,N_2548);
nand U9663 (N_9663,N_5881,N_682);
nor U9664 (N_9664,N_2224,N_254);
or U9665 (N_9665,N_1333,N_5790);
xor U9666 (N_9666,N_3792,N_3686);
nand U9667 (N_9667,N_4447,N_4224);
or U9668 (N_9668,N_1113,N_2099);
xnor U9669 (N_9669,N_5694,N_4595);
nand U9670 (N_9670,N_6247,N_3602);
xnor U9671 (N_9671,N_2302,N_4313);
and U9672 (N_9672,N_834,N_5914);
xor U9673 (N_9673,N_4167,N_6065);
nand U9674 (N_9674,N_5594,N_5574);
nor U9675 (N_9675,N_6213,N_1299);
nand U9676 (N_9676,N_783,N_1286);
xnor U9677 (N_9677,N_4224,N_785);
or U9678 (N_9678,N_782,N_2083);
nor U9679 (N_9679,N_6198,N_972);
and U9680 (N_9680,N_5132,N_3564);
nand U9681 (N_9681,N_2385,N_5779);
nand U9682 (N_9682,N_5590,N_1690);
nand U9683 (N_9683,N_407,N_4139);
nand U9684 (N_9684,N_3916,N_3512);
xor U9685 (N_9685,N_5513,N_4072);
and U9686 (N_9686,N_3143,N_415);
or U9687 (N_9687,N_2743,N_2556);
nor U9688 (N_9688,N_3397,N_5859);
xor U9689 (N_9689,N_3168,N_24);
xor U9690 (N_9690,N_2548,N_2478);
nor U9691 (N_9691,N_1255,N_1892);
nand U9692 (N_9692,N_1454,N_4556);
or U9693 (N_9693,N_3422,N_1290);
or U9694 (N_9694,N_1910,N_5253);
nand U9695 (N_9695,N_3991,N_3001);
nor U9696 (N_9696,N_2843,N_2916);
xor U9697 (N_9697,N_1268,N_3435);
and U9698 (N_9698,N_4409,N_6146);
and U9699 (N_9699,N_3383,N_1658);
or U9700 (N_9700,N_3427,N_4068);
nor U9701 (N_9701,N_1474,N_1856);
xnor U9702 (N_9702,N_1194,N_2262);
xnor U9703 (N_9703,N_2567,N_2251);
nor U9704 (N_9704,N_1551,N_5806);
nand U9705 (N_9705,N_3774,N_585);
nor U9706 (N_9706,N_4380,N_984);
or U9707 (N_9707,N_5625,N_5460);
nand U9708 (N_9708,N_2890,N_4876);
and U9709 (N_9709,N_1397,N_1099);
and U9710 (N_9710,N_2467,N_984);
and U9711 (N_9711,N_873,N_1171);
and U9712 (N_9712,N_3584,N_2636);
or U9713 (N_9713,N_435,N_1256);
nand U9714 (N_9714,N_5564,N_461);
nand U9715 (N_9715,N_810,N_2789);
or U9716 (N_9716,N_2550,N_5347);
or U9717 (N_9717,N_4230,N_4280);
xor U9718 (N_9718,N_5728,N_1991);
nor U9719 (N_9719,N_2107,N_5814);
or U9720 (N_9720,N_1498,N_4232);
nor U9721 (N_9721,N_6244,N_3119);
and U9722 (N_9722,N_3005,N_537);
nand U9723 (N_9723,N_5926,N_2228);
nor U9724 (N_9724,N_3117,N_5453);
nand U9725 (N_9725,N_3246,N_4492);
nand U9726 (N_9726,N_1120,N_4242);
or U9727 (N_9727,N_1584,N_1979);
nand U9728 (N_9728,N_4926,N_3599);
or U9729 (N_9729,N_4378,N_4783);
nor U9730 (N_9730,N_6235,N_346);
nand U9731 (N_9731,N_3605,N_5777);
and U9732 (N_9732,N_73,N_712);
nor U9733 (N_9733,N_5870,N_1223);
xnor U9734 (N_9734,N_5877,N_4683);
nor U9735 (N_9735,N_5440,N_3012);
nor U9736 (N_9736,N_2058,N_1209);
nand U9737 (N_9737,N_3384,N_975);
or U9738 (N_9738,N_1310,N_6000);
nor U9739 (N_9739,N_3003,N_2703);
nor U9740 (N_9740,N_4076,N_4069);
nor U9741 (N_9741,N_1941,N_6020);
nor U9742 (N_9742,N_1526,N_3223);
nor U9743 (N_9743,N_248,N_4277);
xnor U9744 (N_9744,N_1955,N_5181);
and U9745 (N_9745,N_5311,N_2285);
nor U9746 (N_9746,N_221,N_5312);
and U9747 (N_9747,N_4930,N_2166);
nand U9748 (N_9748,N_4811,N_4057);
xnor U9749 (N_9749,N_1101,N_3780);
or U9750 (N_9750,N_3432,N_5541);
or U9751 (N_9751,N_2932,N_307);
nor U9752 (N_9752,N_5636,N_5220);
or U9753 (N_9753,N_6087,N_3531);
and U9754 (N_9754,N_199,N_3906);
xor U9755 (N_9755,N_1855,N_532);
or U9756 (N_9756,N_737,N_4079);
nand U9757 (N_9757,N_1641,N_1166);
and U9758 (N_9758,N_4001,N_4155);
nor U9759 (N_9759,N_4343,N_2833);
xor U9760 (N_9760,N_5018,N_2549);
nor U9761 (N_9761,N_3223,N_5713);
nand U9762 (N_9762,N_2484,N_345);
and U9763 (N_9763,N_3561,N_1562);
nor U9764 (N_9764,N_5591,N_2218);
nor U9765 (N_9765,N_195,N_3681);
and U9766 (N_9766,N_2915,N_499);
nand U9767 (N_9767,N_4645,N_5064);
or U9768 (N_9768,N_117,N_5890);
and U9769 (N_9769,N_3888,N_3893);
xor U9770 (N_9770,N_2003,N_5209);
or U9771 (N_9771,N_5964,N_597);
nor U9772 (N_9772,N_1003,N_348);
or U9773 (N_9773,N_4669,N_1204);
or U9774 (N_9774,N_3083,N_5792);
or U9775 (N_9775,N_4147,N_5703);
nand U9776 (N_9776,N_1651,N_2346);
or U9777 (N_9777,N_770,N_1358);
or U9778 (N_9778,N_5514,N_4416);
nor U9779 (N_9779,N_1486,N_5722);
nand U9780 (N_9780,N_1003,N_2500);
and U9781 (N_9781,N_1005,N_2866);
xor U9782 (N_9782,N_4979,N_5501);
xnor U9783 (N_9783,N_6224,N_4649);
xor U9784 (N_9784,N_469,N_5133);
and U9785 (N_9785,N_2500,N_218);
nor U9786 (N_9786,N_1545,N_4036);
nor U9787 (N_9787,N_5777,N_3810);
and U9788 (N_9788,N_2633,N_1396);
nor U9789 (N_9789,N_3191,N_4427);
nor U9790 (N_9790,N_3157,N_2768);
nor U9791 (N_9791,N_959,N_3507);
or U9792 (N_9792,N_5370,N_2514);
or U9793 (N_9793,N_3380,N_2423);
and U9794 (N_9794,N_1677,N_3131);
nand U9795 (N_9795,N_2516,N_532);
and U9796 (N_9796,N_2276,N_6010);
nand U9797 (N_9797,N_2654,N_5278);
or U9798 (N_9798,N_2536,N_1097);
xor U9799 (N_9799,N_1151,N_3632);
nor U9800 (N_9800,N_3242,N_1358);
or U9801 (N_9801,N_3368,N_2965);
or U9802 (N_9802,N_725,N_5502);
xnor U9803 (N_9803,N_5556,N_4109);
and U9804 (N_9804,N_5873,N_2941);
or U9805 (N_9805,N_6167,N_2854);
nor U9806 (N_9806,N_3022,N_2143);
and U9807 (N_9807,N_1282,N_1745);
nor U9808 (N_9808,N_1146,N_2931);
nor U9809 (N_9809,N_1583,N_3531);
xnor U9810 (N_9810,N_5462,N_805);
and U9811 (N_9811,N_3084,N_5651);
xor U9812 (N_9812,N_5281,N_5901);
nor U9813 (N_9813,N_4536,N_3611);
or U9814 (N_9814,N_5319,N_338);
and U9815 (N_9815,N_4225,N_2020);
and U9816 (N_9816,N_4838,N_2372);
nor U9817 (N_9817,N_3150,N_1143);
or U9818 (N_9818,N_2515,N_406);
nor U9819 (N_9819,N_3937,N_3610);
nor U9820 (N_9820,N_2043,N_2234);
nor U9821 (N_9821,N_4502,N_1892);
nor U9822 (N_9822,N_2900,N_471);
and U9823 (N_9823,N_5760,N_4541);
nor U9824 (N_9824,N_4037,N_1241);
nor U9825 (N_9825,N_5255,N_1054);
xnor U9826 (N_9826,N_4886,N_253);
or U9827 (N_9827,N_4519,N_2583);
or U9828 (N_9828,N_6030,N_5731);
xor U9829 (N_9829,N_3473,N_3913);
xor U9830 (N_9830,N_3415,N_38);
nand U9831 (N_9831,N_3584,N_644);
xnor U9832 (N_9832,N_1070,N_3343);
or U9833 (N_9833,N_5813,N_3252);
xnor U9834 (N_9834,N_518,N_118);
xnor U9835 (N_9835,N_2870,N_3340);
nand U9836 (N_9836,N_3529,N_913);
nor U9837 (N_9837,N_2238,N_5778);
xor U9838 (N_9838,N_4620,N_4595);
or U9839 (N_9839,N_3599,N_3960);
and U9840 (N_9840,N_2610,N_1521);
nand U9841 (N_9841,N_3858,N_883);
xor U9842 (N_9842,N_841,N_948);
xnor U9843 (N_9843,N_5030,N_3241);
xor U9844 (N_9844,N_4082,N_2160);
or U9845 (N_9845,N_2252,N_3354);
nand U9846 (N_9846,N_5792,N_5453);
and U9847 (N_9847,N_4105,N_3928);
xnor U9848 (N_9848,N_945,N_3174);
xnor U9849 (N_9849,N_1336,N_4976);
or U9850 (N_9850,N_1446,N_2817);
or U9851 (N_9851,N_5995,N_5923);
nor U9852 (N_9852,N_403,N_3699);
nand U9853 (N_9853,N_2172,N_5073);
and U9854 (N_9854,N_3117,N_4216);
nor U9855 (N_9855,N_2783,N_1644);
nand U9856 (N_9856,N_3060,N_5964);
xnor U9857 (N_9857,N_4889,N_6188);
nand U9858 (N_9858,N_5997,N_3934);
nor U9859 (N_9859,N_2285,N_4682);
xnor U9860 (N_9860,N_2939,N_4683);
xor U9861 (N_9861,N_1387,N_3984);
or U9862 (N_9862,N_59,N_3728);
nor U9863 (N_9863,N_2146,N_3794);
nand U9864 (N_9864,N_3504,N_373);
nand U9865 (N_9865,N_2464,N_1266);
nand U9866 (N_9866,N_1361,N_2872);
nand U9867 (N_9867,N_4699,N_353);
nor U9868 (N_9868,N_3733,N_6024);
or U9869 (N_9869,N_3747,N_208);
and U9870 (N_9870,N_2009,N_3981);
and U9871 (N_9871,N_4432,N_6210);
nand U9872 (N_9872,N_5326,N_3738);
nor U9873 (N_9873,N_3083,N_4398);
nand U9874 (N_9874,N_5204,N_4848);
or U9875 (N_9875,N_902,N_4169);
nand U9876 (N_9876,N_5937,N_5704);
xor U9877 (N_9877,N_2478,N_4018);
nor U9878 (N_9878,N_2031,N_4916);
xor U9879 (N_9879,N_2845,N_2886);
and U9880 (N_9880,N_4695,N_4033);
nand U9881 (N_9881,N_4852,N_3445);
nor U9882 (N_9882,N_893,N_2391);
xnor U9883 (N_9883,N_6002,N_3611);
nand U9884 (N_9884,N_2929,N_3371);
xor U9885 (N_9885,N_4960,N_3980);
nor U9886 (N_9886,N_5564,N_1875);
and U9887 (N_9887,N_4624,N_4589);
or U9888 (N_9888,N_2095,N_1233);
nor U9889 (N_9889,N_2834,N_4728);
or U9890 (N_9890,N_1032,N_671);
nor U9891 (N_9891,N_1406,N_603);
xnor U9892 (N_9892,N_2000,N_4056);
xnor U9893 (N_9893,N_859,N_5457);
nand U9894 (N_9894,N_3045,N_4655);
or U9895 (N_9895,N_4788,N_3186);
or U9896 (N_9896,N_6177,N_771);
xnor U9897 (N_9897,N_5465,N_6000);
nor U9898 (N_9898,N_6082,N_5933);
nor U9899 (N_9899,N_5264,N_5998);
or U9900 (N_9900,N_4151,N_5916);
xnor U9901 (N_9901,N_5215,N_214);
nand U9902 (N_9902,N_5250,N_2431);
xor U9903 (N_9903,N_781,N_4290);
and U9904 (N_9904,N_1812,N_4963);
xor U9905 (N_9905,N_5100,N_216);
or U9906 (N_9906,N_3017,N_4876);
and U9907 (N_9907,N_5575,N_97);
or U9908 (N_9908,N_2219,N_5539);
or U9909 (N_9909,N_5422,N_2323);
nand U9910 (N_9910,N_6208,N_4555);
and U9911 (N_9911,N_3516,N_6151);
or U9912 (N_9912,N_3456,N_4295);
or U9913 (N_9913,N_1280,N_1997);
nand U9914 (N_9914,N_544,N_4204);
or U9915 (N_9915,N_1043,N_5995);
nand U9916 (N_9916,N_1411,N_311);
or U9917 (N_9917,N_1517,N_3191);
nor U9918 (N_9918,N_2228,N_4867);
xor U9919 (N_9919,N_2445,N_1075);
xor U9920 (N_9920,N_5470,N_2314);
or U9921 (N_9921,N_892,N_3741);
nand U9922 (N_9922,N_206,N_3516);
or U9923 (N_9923,N_1891,N_2230);
nand U9924 (N_9924,N_5519,N_4400);
xnor U9925 (N_9925,N_1419,N_1647);
nor U9926 (N_9926,N_1497,N_2800);
and U9927 (N_9927,N_3066,N_3870);
xor U9928 (N_9928,N_1877,N_1459);
nor U9929 (N_9929,N_2683,N_511);
or U9930 (N_9930,N_6210,N_2439);
nand U9931 (N_9931,N_4433,N_2081);
nor U9932 (N_9932,N_1267,N_5486);
or U9933 (N_9933,N_1783,N_2030);
nor U9934 (N_9934,N_1656,N_1554);
nand U9935 (N_9935,N_2214,N_1267);
and U9936 (N_9936,N_1303,N_3303);
and U9937 (N_9937,N_2724,N_2131);
or U9938 (N_9938,N_5444,N_3526);
xor U9939 (N_9939,N_5495,N_383);
or U9940 (N_9940,N_300,N_3390);
nor U9941 (N_9941,N_1523,N_1481);
nand U9942 (N_9942,N_2337,N_1640);
xnor U9943 (N_9943,N_5729,N_4598);
or U9944 (N_9944,N_1789,N_3726);
nand U9945 (N_9945,N_2272,N_5857);
nand U9946 (N_9946,N_2944,N_4107);
or U9947 (N_9947,N_1023,N_1723);
nor U9948 (N_9948,N_3219,N_3943);
and U9949 (N_9949,N_1285,N_1258);
nor U9950 (N_9950,N_2037,N_1150);
nor U9951 (N_9951,N_2233,N_219);
nor U9952 (N_9952,N_3768,N_4049);
xnor U9953 (N_9953,N_2336,N_1675);
and U9954 (N_9954,N_4590,N_3264);
xor U9955 (N_9955,N_2234,N_3373);
nor U9956 (N_9956,N_4121,N_616);
nor U9957 (N_9957,N_5288,N_3647);
nor U9958 (N_9958,N_3716,N_1651);
xnor U9959 (N_9959,N_1965,N_1583);
nor U9960 (N_9960,N_4444,N_1825);
nor U9961 (N_9961,N_3906,N_4800);
nand U9962 (N_9962,N_4720,N_4861);
nand U9963 (N_9963,N_717,N_1924);
xnor U9964 (N_9964,N_1953,N_4257);
nand U9965 (N_9965,N_6106,N_4060);
and U9966 (N_9966,N_4626,N_5778);
or U9967 (N_9967,N_5921,N_2202);
nor U9968 (N_9968,N_4106,N_4935);
or U9969 (N_9969,N_5440,N_4996);
nand U9970 (N_9970,N_1056,N_3158);
and U9971 (N_9971,N_3603,N_260);
xnor U9972 (N_9972,N_2557,N_399);
xnor U9973 (N_9973,N_932,N_5625);
and U9974 (N_9974,N_3169,N_4929);
nor U9975 (N_9975,N_35,N_1428);
xor U9976 (N_9976,N_857,N_4139);
nand U9977 (N_9977,N_947,N_4883);
nor U9978 (N_9978,N_5547,N_749);
nor U9979 (N_9979,N_1097,N_2167);
nand U9980 (N_9980,N_5234,N_5274);
or U9981 (N_9981,N_1071,N_3373);
or U9982 (N_9982,N_3537,N_6201);
xor U9983 (N_9983,N_3741,N_1767);
nand U9984 (N_9984,N_337,N_4018);
or U9985 (N_9985,N_1266,N_2829);
xor U9986 (N_9986,N_2650,N_1500);
nand U9987 (N_9987,N_5466,N_1994);
nand U9988 (N_9988,N_5312,N_2687);
nor U9989 (N_9989,N_4609,N_1440);
and U9990 (N_9990,N_1668,N_4394);
nand U9991 (N_9991,N_2647,N_3043);
xor U9992 (N_9992,N_575,N_5473);
nand U9993 (N_9993,N_5024,N_5279);
xnor U9994 (N_9994,N_3726,N_1959);
xnor U9995 (N_9995,N_642,N_3346);
and U9996 (N_9996,N_2443,N_2955);
nand U9997 (N_9997,N_182,N_721);
nor U9998 (N_9998,N_4689,N_784);
or U9999 (N_9999,N_1899,N_3138);
xor U10000 (N_10000,N_2186,N_5106);
nor U10001 (N_10001,N_2860,N_5121);
nor U10002 (N_10002,N_5642,N_5294);
and U10003 (N_10003,N_5281,N_4013);
nor U10004 (N_10004,N_959,N_239);
nand U10005 (N_10005,N_6071,N_989);
nand U10006 (N_10006,N_1036,N_6063);
xnor U10007 (N_10007,N_2845,N_895);
nor U10008 (N_10008,N_4366,N_4944);
nand U10009 (N_10009,N_5443,N_858);
or U10010 (N_10010,N_3387,N_322);
nor U10011 (N_10011,N_2066,N_1287);
nand U10012 (N_10012,N_1022,N_3615);
or U10013 (N_10013,N_4769,N_1679);
or U10014 (N_10014,N_1150,N_5068);
or U10015 (N_10015,N_5602,N_796);
or U10016 (N_10016,N_1672,N_524);
and U10017 (N_10017,N_806,N_188);
nand U10018 (N_10018,N_6036,N_1252);
nand U10019 (N_10019,N_4886,N_3639);
and U10020 (N_10020,N_814,N_2398);
xor U10021 (N_10021,N_2632,N_55);
xor U10022 (N_10022,N_6050,N_4111);
and U10023 (N_10023,N_165,N_702);
or U10024 (N_10024,N_4811,N_1927);
and U10025 (N_10025,N_416,N_2430);
or U10026 (N_10026,N_2141,N_4979);
nor U10027 (N_10027,N_3676,N_3188);
nand U10028 (N_10028,N_3543,N_5439);
nand U10029 (N_10029,N_3756,N_294);
and U10030 (N_10030,N_3139,N_370);
nand U10031 (N_10031,N_3247,N_4891);
xnor U10032 (N_10032,N_3551,N_5168);
nor U10033 (N_10033,N_450,N_3562);
xor U10034 (N_10034,N_2449,N_5095);
and U10035 (N_10035,N_2573,N_5283);
nor U10036 (N_10036,N_4828,N_6099);
xnor U10037 (N_10037,N_2942,N_5071);
or U10038 (N_10038,N_4965,N_90);
nand U10039 (N_10039,N_6192,N_1771);
nand U10040 (N_10040,N_4397,N_3495);
and U10041 (N_10041,N_1367,N_5982);
xor U10042 (N_10042,N_1715,N_4847);
or U10043 (N_10043,N_849,N_56);
nor U10044 (N_10044,N_5849,N_6243);
nor U10045 (N_10045,N_2839,N_530);
nor U10046 (N_10046,N_4963,N_4750);
xor U10047 (N_10047,N_134,N_4475);
nor U10048 (N_10048,N_1752,N_2786);
or U10049 (N_10049,N_1332,N_1078);
and U10050 (N_10050,N_4758,N_5686);
xnor U10051 (N_10051,N_6137,N_4624);
nand U10052 (N_10052,N_3389,N_2742);
nor U10053 (N_10053,N_3058,N_5644);
nand U10054 (N_10054,N_5546,N_6107);
xor U10055 (N_10055,N_2186,N_3112);
and U10056 (N_10056,N_2713,N_2336);
nor U10057 (N_10057,N_4219,N_2972);
nor U10058 (N_10058,N_4663,N_3184);
or U10059 (N_10059,N_3727,N_304);
nand U10060 (N_10060,N_1505,N_1922);
or U10061 (N_10061,N_5547,N_4279);
xor U10062 (N_10062,N_3418,N_647);
xor U10063 (N_10063,N_1309,N_2998);
xnor U10064 (N_10064,N_1194,N_5448);
nor U10065 (N_10065,N_1457,N_3487);
xnor U10066 (N_10066,N_6051,N_5830);
or U10067 (N_10067,N_3285,N_4378);
or U10068 (N_10068,N_5969,N_5801);
and U10069 (N_10069,N_4853,N_2629);
nand U10070 (N_10070,N_3916,N_109);
nor U10071 (N_10071,N_6125,N_3265);
nor U10072 (N_10072,N_4362,N_4053);
and U10073 (N_10073,N_2609,N_2350);
nand U10074 (N_10074,N_2238,N_5062);
nor U10075 (N_10075,N_4970,N_2620);
or U10076 (N_10076,N_4730,N_3507);
and U10077 (N_10077,N_2965,N_3062);
xnor U10078 (N_10078,N_1489,N_2843);
or U10079 (N_10079,N_2295,N_2840);
xor U10080 (N_10080,N_2902,N_2054);
or U10081 (N_10081,N_1503,N_6016);
xor U10082 (N_10082,N_5513,N_4705);
and U10083 (N_10083,N_408,N_4422);
nor U10084 (N_10084,N_4445,N_2862);
nor U10085 (N_10085,N_946,N_1792);
nor U10086 (N_10086,N_2386,N_2532);
xnor U10087 (N_10087,N_5402,N_1075);
xnor U10088 (N_10088,N_3583,N_5114);
nor U10089 (N_10089,N_5515,N_6155);
nor U10090 (N_10090,N_673,N_3887);
xnor U10091 (N_10091,N_1615,N_1906);
xnor U10092 (N_10092,N_2898,N_3668);
and U10093 (N_10093,N_4104,N_1670);
nor U10094 (N_10094,N_3457,N_5594);
and U10095 (N_10095,N_5956,N_4988);
or U10096 (N_10096,N_1205,N_1520);
nor U10097 (N_10097,N_5190,N_3857);
nand U10098 (N_10098,N_3314,N_4132);
or U10099 (N_10099,N_1948,N_946);
nand U10100 (N_10100,N_3655,N_2572);
xor U10101 (N_10101,N_249,N_4677);
nand U10102 (N_10102,N_5586,N_1235);
nand U10103 (N_10103,N_4495,N_5647);
or U10104 (N_10104,N_5059,N_1636);
nand U10105 (N_10105,N_6010,N_3259);
nor U10106 (N_10106,N_2861,N_1762);
xor U10107 (N_10107,N_5077,N_6128);
nor U10108 (N_10108,N_6232,N_6098);
nor U10109 (N_10109,N_3238,N_686);
xor U10110 (N_10110,N_12,N_2900);
xnor U10111 (N_10111,N_2973,N_2915);
xor U10112 (N_10112,N_3308,N_4187);
or U10113 (N_10113,N_5470,N_741);
xor U10114 (N_10114,N_5901,N_2480);
and U10115 (N_10115,N_1280,N_3835);
nor U10116 (N_10116,N_4945,N_232);
or U10117 (N_10117,N_6125,N_2449);
and U10118 (N_10118,N_603,N_5631);
xor U10119 (N_10119,N_2162,N_4920);
or U10120 (N_10120,N_314,N_455);
nand U10121 (N_10121,N_1183,N_1458);
or U10122 (N_10122,N_83,N_3268);
nand U10123 (N_10123,N_2274,N_2975);
and U10124 (N_10124,N_764,N_2946);
xor U10125 (N_10125,N_160,N_5226);
and U10126 (N_10126,N_4153,N_2953);
or U10127 (N_10127,N_5616,N_2752);
or U10128 (N_10128,N_2283,N_3730);
nand U10129 (N_10129,N_1132,N_2885);
or U10130 (N_10130,N_3441,N_2061);
nor U10131 (N_10131,N_3710,N_3886);
nand U10132 (N_10132,N_1886,N_2509);
or U10133 (N_10133,N_1011,N_2738);
or U10134 (N_10134,N_2845,N_3412);
xor U10135 (N_10135,N_1933,N_3232);
xor U10136 (N_10136,N_3226,N_3695);
nand U10137 (N_10137,N_227,N_5839);
nand U10138 (N_10138,N_5536,N_1876);
and U10139 (N_10139,N_3370,N_2383);
nor U10140 (N_10140,N_671,N_266);
or U10141 (N_10141,N_216,N_5933);
or U10142 (N_10142,N_1453,N_5340);
or U10143 (N_10143,N_2026,N_1959);
xnor U10144 (N_10144,N_5935,N_663);
xnor U10145 (N_10145,N_3522,N_1289);
xor U10146 (N_10146,N_1726,N_3973);
and U10147 (N_10147,N_5046,N_3440);
or U10148 (N_10148,N_4419,N_5971);
or U10149 (N_10149,N_3553,N_1480);
nor U10150 (N_10150,N_3461,N_4959);
xor U10151 (N_10151,N_4796,N_2949);
nand U10152 (N_10152,N_4814,N_1360);
xor U10153 (N_10153,N_1753,N_4880);
and U10154 (N_10154,N_6123,N_87);
and U10155 (N_10155,N_301,N_5708);
nand U10156 (N_10156,N_3803,N_4841);
or U10157 (N_10157,N_236,N_4766);
xor U10158 (N_10158,N_876,N_4426);
nor U10159 (N_10159,N_461,N_3822);
nor U10160 (N_10160,N_1434,N_3746);
nand U10161 (N_10161,N_1326,N_1327);
nand U10162 (N_10162,N_1674,N_6124);
nor U10163 (N_10163,N_2493,N_4459);
and U10164 (N_10164,N_3729,N_5436);
nand U10165 (N_10165,N_1080,N_3904);
nand U10166 (N_10166,N_5872,N_291);
or U10167 (N_10167,N_3725,N_1544);
xor U10168 (N_10168,N_1579,N_3349);
xor U10169 (N_10169,N_1735,N_4818);
nor U10170 (N_10170,N_5248,N_3312);
or U10171 (N_10171,N_4955,N_3438);
nand U10172 (N_10172,N_348,N_3303);
xnor U10173 (N_10173,N_881,N_741);
nor U10174 (N_10174,N_4516,N_4529);
nand U10175 (N_10175,N_4661,N_318);
nand U10176 (N_10176,N_5189,N_5141);
nand U10177 (N_10177,N_6137,N_133);
and U10178 (N_10178,N_6197,N_5088);
xnor U10179 (N_10179,N_6246,N_1707);
or U10180 (N_10180,N_1001,N_2308);
and U10181 (N_10181,N_2551,N_3832);
or U10182 (N_10182,N_2039,N_4299);
xor U10183 (N_10183,N_4726,N_4759);
or U10184 (N_10184,N_856,N_758);
and U10185 (N_10185,N_3133,N_1480);
xor U10186 (N_10186,N_5252,N_1504);
xnor U10187 (N_10187,N_527,N_1734);
and U10188 (N_10188,N_5683,N_1855);
nand U10189 (N_10189,N_296,N_4577);
nand U10190 (N_10190,N_3633,N_1250);
nor U10191 (N_10191,N_574,N_60);
nand U10192 (N_10192,N_513,N_3033);
or U10193 (N_10193,N_6140,N_287);
xor U10194 (N_10194,N_5411,N_3036);
nor U10195 (N_10195,N_4379,N_4164);
nand U10196 (N_10196,N_2701,N_3929);
nor U10197 (N_10197,N_623,N_3662);
nor U10198 (N_10198,N_4340,N_4042);
xor U10199 (N_10199,N_4075,N_4004);
or U10200 (N_10200,N_2899,N_4001);
or U10201 (N_10201,N_472,N_402);
nand U10202 (N_10202,N_1553,N_3231);
nand U10203 (N_10203,N_3442,N_1999);
and U10204 (N_10204,N_3830,N_1856);
or U10205 (N_10205,N_1927,N_4052);
and U10206 (N_10206,N_5093,N_6000);
and U10207 (N_10207,N_2568,N_3867);
or U10208 (N_10208,N_2223,N_3080);
nand U10209 (N_10209,N_2289,N_3828);
and U10210 (N_10210,N_4742,N_3803);
or U10211 (N_10211,N_3734,N_5126);
and U10212 (N_10212,N_2220,N_6046);
xnor U10213 (N_10213,N_4499,N_5553);
nand U10214 (N_10214,N_288,N_5492);
or U10215 (N_10215,N_4504,N_5722);
xor U10216 (N_10216,N_5378,N_1440);
or U10217 (N_10217,N_760,N_5052);
xnor U10218 (N_10218,N_3459,N_3529);
xor U10219 (N_10219,N_1824,N_1301);
or U10220 (N_10220,N_4370,N_6078);
and U10221 (N_10221,N_5671,N_4071);
nand U10222 (N_10222,N_1369,N_128);
and U10223 (N_10223,N_2313,N_87);
xnor U10224 (N_10224,N_2746,N_1924);
nor U10225 (N_10225,N_2521,N_396);
nor U10226 (N_10226,N_55,N_2372);
xnor U10227 (N_10227,N_1971,N_5585);
or U10228 (N_10228,N_4878,N_3436);
nand U10229 (N_10229,N_5219,N_2148);
nor U10230 (N_10230,N_5387,N_3214);
xor U10231 (N_10231,N_1221,N_4090);
and U10232 (N_10232,N_1470,N_4307);
xor U10233 (N_10233,N_3187,N_2434);
or U10234 (N_10234,N_1636,N_4402);
nand U10235 (N_10235,N_2861,N_3387);
nand U10236 (N_10236,N_2290,N_2712);
xor U10237 (N_10237,N_4553,N_3620);
and U10238 (N_10238,N_4573,N_6222);
nor U10239 (N_10239,N_87,N_4775);
or U10240 (N_10240,N_1665,N_4184);
and U10241 (N_10241,N_4273,N_3906);
and U10242 (N_10242,N_1388,N_1155);
or U10243 (N_10243,N_645,N_6144);
and U10244 (N_10244,N_5303,N_1634);
nor U10245 (N_10245,N_5980,N_1096);
nor U10246 (N_10246,N_244,N_4069);
nor U10247 (N_10247,N_5850,N_2371);
xnor U10248 (N_10248,N_4173,N_3038);
or U10249 (N_10249,N_4084,N_3523);
or U10250 (N_10250,N_1199,N_1634);
or U10251 (N_10251,N_910,N_3353);
or U10252 (N_10252,N_4939,N_3118);
nand U10253 (N_10253,N_2960,N_4920);
nor U10254 (N_10254,N_6045,N_3501);
or U10255 (N_10255,N_4763,N_2371);
xor U10256 (N_10256,N_5455,N_5290);
or U10257 (N_10257,N_5876,N_2330);
xor U10258 (N_10258,N_285,N_1696);
nor U10259 (N_10259,N_626,N_4732);
or U10260 (N_10260,N_2268,N_4394);
nand U10261 (N_10261,N_483,N_5334);
and U10262 (N_10262,N_4284,N_1);
nor U10263 (N_10263,N_3784,N_1192);
nor U10264 (N_10264,N_571,N_1930);
and U10265 (N_10265,N_126,N_2592);
and U10266 (N_10266,N_211,N_3691);
nand U10267 (N_10267,N_5438,N_2843);
xnor U10268 (N_10268,N_2210,N_5084);
and U10269 (N_10269,N_3469,N_5447);
nand U10270 (N_10270,N_5194,N_3276);
nand U10271 (N_10271,N_114,N_4369);
xor U10272 (N_10272,N_1686,N_1764);
nand U10273 (N_10273,N_2023,N_2006);
nor U10274 (N_10274,N_3834,N_3591);
and U10275 (N_10275,N_1932,N_3173);
xnor U10276 (N_10276,N_2123,N_5623);
nand U10277 (N_10277,N_4652,N_459);
nand U10278 (N_10278,N_4774,N_3331);
nor U10279 (N_10279,N_1515,N_5114);
or U10280 (N_10280,N_2599,N_2744);
nand U10281 (N_10281,N_1086,N_5186);
xor U10282 (N_10282,N_1351,N_601);
or U10283 (N_10283,N_498,N_1846);
or U10284 (N_10284,N_5267,N_5750);
or U10285 (N_10285,N_1468,N_1034);
and U10286 (N_10286,N_5696,N_6073);
nor U10287 (N_10287,N_5879,N_5096);
xor U10288 (N_10288,N_514,N_4113);
and U10289 (N_10289,N_4568,N_5627);
nor U10290 (N_10290,N_4839,N_5691);
xor U10291 (N_10291,N_4557,N_162);
nor U10292 (N_10292,N_4591,N_5607);
or U10293 (N_10293,N_4543,N_5110);
nor U10294 (N_10294,N_2697,N_2916);
or U10295 (N_10295,N_3036,N_5379);
and U10296 (N_10296,N_4638,N_547);
nor U10297 (N_10297,N_1671,N_5479);
and U10298 (N_10298,N_3122,N_6199);
nand U10299 (N_10299,N_3378,N_5354);
xor U10300 (N_10300,N_1251,N_2842);
and U10301 (N_10301,N_5166,N_54);
nand U10302 (N_10302,N_2048,N_722);
or U10303 (N_10303,N_1571,N_4870);
nand U10304 (N_10304,N_3607,N_2299);
and U10305 (N_10305,N_4959,N_667);
xnor U10306 (N_10306,N_1764,N_4485);
xnor U10307 (N_10307,N_5916,N_1436);
and U10308 (N_10308,N_4407,N_4004);
nand U10309 (N_10309,N_5778,N_5045);
xor U10310 (N_10310,N_4131,N_2253);
or U10311 (N_10311,N_3118,N_4422);
nand U10312 (N_10312,N_5359,N_3842);
and U10313 (N_10313,N_3814,N_3715);
nor U10314 (N_10314,N_2917,N_2984);
nand U10315 (N_10315,N_3850,N_5634);
xor U10316 (N_10316,N_4314,N_4513);
or U10317 (N_10317,N_5002,N_3555);
or U10318 (N_10318,N_2269,N_1292);
nor U10319 (N_10319,N_1262,N_4966);
and U10320 (N_10320,N_3260,N_3884);
xor U10321 (N_10321,N_1260,N_4186);
or U10322 (N_10322,N_3082,N_272);
and U10323 (N_10323,N_2954,N_5389);
xnor U10324 (N_10324,N_351,N_2912);
nor U10325 (N_10325,N_6214,N_1010);
xor U10326 (N_10326,N_1545,N_94);
and U10327 (N_10327,N_3432,N_5142);
nor U10328 (N_10328,N_2917,N_4921);
nand U10329 (N_10329,N_2855,N_5622);
or U10330 (N_10330,N_5085,N_2131);
xor U10331 (N_10331,N_3173,N_4698);
or U10332 (N_10332,N_1543,N_972);
xnor U10333 (N_10333,N_602,N_4771);
and U10334 (N_10334,N_1829,N_6041);
nand U10335 (N_10335,N_1736,N_1915);
nor U10336 (N_10336,N_692,N_3882);
nand U10337 (N_10337,N_2540,N_3818);
nand U10338 (N_10338,N_5006,N_1334);
nor U10339 (N_10339,N_3195,N_2479);
xor U10340 (N_10340,N_3524,N_3432);
nand U10341 (N_10341,N_2714,N_3271);
xnor U10342 (N_10342,N_1736,N_1562);
or U10343 (N_10343,N_2293,N_5981);
nand U10344 (N_10344,N_2039,N_904);
nor U10345 (N_10345,N_4541,N_417);
or U10346 (N_10346,N_3069,N_1866);
nand U10347 (N_10347,N_1174,N_3585);
nand U10348 (N_10348,N_978,N_556);
nor U10349 (N_10349,N_3618,N_424);
and U10350 (N_10350,N_2165,N_5473);
xor U10351 (N_10351,N_4816,N_1890);
nand U10352 (N_10352,N_3577,N_1990);
nand U10353 (N_10353,N_6246,N_1634);
nor U10354 (N_10354,N_4953,N_5849);
nor U10355 (N_10355,N_587,N_306);
xor U10356 (N_10356,N_157,N_4506);
or U10357 (N_10357,N_5581,N_1033);
xor U10358 (N_10358,N_3406,N_5075);
and U10359 (N_10359,N_4665,N_3757);
xnor U10360 (N_10360,N_92,N_433);
nand U10361 (N_10361,N_5206,N_3091);
xnor U10362 (N_10362,N_1468,N_3470);
and U10363 (N_10363,N_3715,N_5865);
and U10364 (N_10364,N_1681,N_2696);
and U10365 (N_10365,N_3483,N_2904);
and U10366 (N_10366,N_5460,N_3239);
xnor U10367 (N_10367,N_446,N_3875);
and U10368 (N_10368,N_5541,N_3532);
xnor U10369 (N_10369,N_304,N_5421);
xnor U10370 (N_10370,N_3190,N_1977);
nor U10371 (N_10371,N_4980,N_1514);
nor U10372 (N_10372,N_4899,N_6040);
or U10373 (N_10373,N_4422,N_6014);
nor U10374 (N_10374,N_5021,N_3627);
and U10375 (N_10375,N_4605,N_4602);
or U10376 (N_10376,N_4481,N_4724);
xor U10377 (N_10377,N_5317,N_4536);
nor U10378 (N_10378,N_380,N_1942);
or U10379 (N_10379,N_3752,N_2918);
or U10380 (N_10380,N_5406,N_501);
nand U10381 (N_10381,N_619,N_3872);
nor U10382 (N_10382,N_4748,N_5238);
xor U10383 (N_10383,N_20,N_5183);
and U10384 (N_10384,N_584,N_634);
nor U10385 (N_10385,N_1993,N_3569);
xnor U10386 (N_10386,N_1804,N_5090);
nor U10387 (N_10387,N_3272,N_4408);
xnor U10388 (N_10388,N_1234,N_4967);
nor U10389 (N_10389,N_2262,N_163);
xor U10390 (N_10390,N_5739,N_834);
or U10391 (N_10391,N_5913,N_5817);
nor U10392 (N_10392,N_937,N_2781);
and U10393 (N_10393,N_753,N_2754);
and U10394 (N_10394,N_2657,N_3539);
xnor U10395 (N_10395,N_1688,N_654);
nand U10396 (N_10396,N_1221,N_3046);
and U10397 (N_10397,N_3610,N_1180);
nand U10398 (N_10398,N_105,N_3867);
or U10399 (N_10399,N_5512,N_5794);
nand U10400 (N_10400,N_5504,N_1330);
or U10401 (N_10401,N_953,N_168);
and U10402 (N_10402,N_4374,N_814);
nor U10403 (N_10403,N_3266,N_3156);
xor U10404 (N_10404,N_4402,N_5449);
nand U10405 (N_10405,N_5582,N_4465);
xnor U10406 (N_10406,N_3472,N_3799);
xor U10407 (N_10407,N_1089,N_3201);
nand U10408 (N_10408,N_2447,N_3713);
nor U10409 (N_10409,N_335,N_1924);
or U10410 (N_10410,N_3166,N_1049);
or U10411 (N_10411,N_4105,N_1741);
or U10412 (N_10412,N_3844,N_2868);
nor U10413 (N_10413,N_247,N_4429);
nand U10414 (N_10414,N_1307,N_3362);
nor U10415 (N_10415,N_1003,N_1775);
nand U10416 (N_10416,N_340,N_5721);
and U10417 (N_10417,N_5201,N_2665);
or U10418 (N_10418,N_3506,N_5707);
and U10419 (N_10419,N_3230,N_2608);
nor U10420 (N_10420,N_4307,N_6169);
xnor U10421 (N_10421,N_135,N_3823);
nand U10422 (N_10422,N_4851,N_3727);
nand U10423 (N_10423,N_5933,N_4265);
and U10424 (N_10424,N_285,N_4470);
xnor U10425 (N_10425,N_1227,N_2124);
xnor U10426 (N_10426,N_1399,N_2695);
nor U10427 (N_10427,N_4593,N_5340);
or U10428 (N_10428,N_1557,N_3846);
nand U10429 (N_10429,N_5263,N_5344);
and U10430 (N_10430,N_4606,N_5285);
nand U10431 (N_10431,N_3383,N_2775);
nand U10432 (N_10432,N_1692,N_4877);
nor U10433 (N_10433,N_4321,N_4859);
nand U10434 (N_10434,N_2811,N_2777);
xor U10435 (N_10435,N_427,N_155);
nor U10436 (N_10436,N_4194,N_4154);
xnor U10437 (N_10437,N_1770,N_5236);
xor U10438 (N_10438,N_238,N_332);
nand U10439 (N_10439,N_2374,N_374);
or U10440 (N_10440,N_1039,N_5586);
xnor U10441 (N_10441,N_4729,N_453);
and U10442 (N_10442,N_6130,N_939);
and U10443 (N_10443,N_2260,N_3520);
xnor U10444 (N_10444,N_4785,N_2433);
nor U10445 (N_10445,N_4155,N_5974);
or U10446 (N_10446,N_766,N_1350);
nand U10447 (N_10447,N_5314,N_936);
nor U10448 (N_10448,N_5408,N_2765);
xor U10449 (N_10449,N_3206,N_3738);
nand U10450 (N_10450,N_4759,N_2484);
or U10451 (N_10451,N_2124,N_6);
or U10452 (N_10452,N_3441,N_3379);
nor U10453 (N_10453,N_1507,N_536);
xor U10454 (N_10454,N_2399,N_2851);
or U10455 (N_10455,N_5941,N_4037);
and U10456 (N_10456,N_2198,N_3643);
and U10457 (N_10457,N_1119,N_2499);
and U10458 (N_10458,N_1151,N_4412);
nand U10459 (N_10459,N_1114,N_5150);
and U10460 (N_10460,N_4885,N_184);
nand U10461 (N_10461,N_539,N_3527);
nand U10462 (N_10462,N_1396,N_4226);
or U10463 (N_10463,N_336,N_1252);
nand U10464 (N_10464,N_5630,N_221);
nand U10465 (N_10465,N_3182,N_523);
nand U10466 (N_10466,N_4026,N_6072);
or U10467 (N_10467,N_2950,N_4569);
and U10468 (N_10468,N_3868,N_3460);
nor U10469 (N_10469,N_1884,N_3961);
and U10470 (N_10470,N_582,N_4775);
nand U10471 (N_10471,N_1361,N_4022);
nor U10472 (N_10472,N_969,N_5823);
xnor U10473 (N_10473,N_3331,N_2580);
nor U10474 (N_10474,N_3539,N_2173);
xnor U10475 (N_10475,N_5400,N_3813);
and U10476 (N_10476,N_512,N_3986);
and U10477 (N_10477,N_3011,N_1117);
or U10478 (N_10478,N_4774,N_2526);
and U10479 (N_10479,N_5345,N_172);
nand U10480 (N_10480,N_435,N_2418);
and U10481 (N_10481,N_2952,N_490);
nand U10482 (N_10482,N_3672,N_3423);
xnor U10483 (N_10483,N_4845,N_5785);
or U10484 (N_10484,N_3200,N_4006);
xor U10485 (N_10485,N_2104,N_6231);
and U10486 (N_10486,N_5848,N_2243);
or U10487 (N_10487,N_5747,N_5671);
or U10488 (N_10488,N_3227,N_4303);
and U10489 (N_10489,N_4632,N_5298);
nand U10490 (N_10490,N_2243,N_1277);
nand U10491 (N_10491,N_6171,N_3133);
nor U10492 (N_10492,N_2342,N_826);
nor U10493 (N_10493,N_2402,N_3734);
and U10494 (N_10494,N_2879,N_5696);
or U10495 (N_10495,N_5810,N_2982);
nand U10496 (N_10496,N_1448,N_3954);
nand U10497 (N_10497,N_6065,N_3268);
nor U10498 (N_10498,N_4729,N_5330);
xnor U10499 (N_10499,N_1725,N_240);
nand U10500 (N_10500,N_4827,N_2914);
nor U10501 (N_10501,N_5406,N_4872);
nor U10502 (N_10502,N_3382,N_4324);
and U10503 (N_10503,N_1706,N_5021);
or U10504 (N_10504,N_1797,N_2156);
nor U10505 (N_10505,N_2349,N_1543);
xor U10506 (N_10506,N_3911,N_1988);
and U10507 (N_10507,N_574,N_176);
nand U10508 (N_10508,N_1236,N_1140);
nand U10509 (N_10509,N_4980,N_2607);
nor U10510 (N_10510,N_5860,N_3003);
or U10511 (N_10511,N_3144,N_4966);
nor U10512 (N_10512,N_2199,N_5879);
and U10513 (N_10513,N_949,N_1836);
or U10514 (N_10514,N_1757,N_3447);
nand U10515 (N_10515,N_981,N_719);
nor U10516 (N_10516,N_2367,N_1569);
and U10517 (N_10517,N_1613,N_4423);
nand U10518 (N_10518,N_5405,N_4950);
nand U10519 (N_10519,N_2520,N_3112);
and U10520 (N_10520,N_1330,N_2692);
xnor U10521 (N_10521,N_4848,N_3865);
xor U10522 (N_10522,N_3439,N_2502);
nor U10523 (N_10523,N_2690,N_4926);
nor U10524 (N_10524,N_3944,N_1479);
and U10525 (N_10525,N_4746,N_1841);
nand U10526 (N_10526,N_33,N_5013);
nor U10527 (N_10527,N_458,N_2982);
nand U10528 (N_10528,N_188,N_2832);
or U10529 (N_10529,N_1700,N_1144);
nand U10530 (N_10530,N_2318,N_1598);
xnor U10531 (N_10531,N_5890,N_2004);
or U10532 (N_10532,N_1118,N_283);
or U10533 (N_10533,N_3625,N_346);
nor U10534 (N_10534,N_3710,N_1840);
xnor U10535 (N_10535,N_4939,N_265);
and U10536 (N_10536,N_3092,N_2120);
or U10537 (N_10537,N_210,N_1691);
or U10538 (N_10538,N_5142,N_5379);
xnor U10539 (N_10539,N_3648,N_4171);
xnor U10540 (N_10540,N_5229,N_623);
nor U10541 (N_10541,N_2983,N_5328);
xnor U10542 (N_10542,N_54,N_4722);
and U10543 (N_10543,N_4407,N_3795);
nand U10544 (N_10544,N_155,N_25);
nor U10545 (N_10545,N_2574,N_5707);
and U10546 (N_10546,N_4109,N_5066);
xor U10547 (N_10547,N_3293,N_6006);
nor U10548 (N_10548,N_5328,N_4204);
and U10549 (N_10549,N_5149,N_6008);
and U10550 (N_10550,N_5137,N_469);
xor U10551 (N_10551,N_2300,N_2868);
and U10552 (N_10552,N_4418,N_2329);
and U10553 (N_10553,N_3183,N_2313);
and U10554 (N_10554,N_5921,N_2123);
or U10555 (N_10555,N_3439,N_4029);
and U10556 (N_10556,N_2367,N_4397);
xnor U10557 (N_10557,N_2513,N_1513);
nand U10558 (N_10558,N_2558,N_1831);
nand U10559 (N_10559,N_4143,N_3156);
nor U10560 (N_10560,N_5013,N_5700);
and U10561 (N_10561,N_1922,N_758);
or U10562 (N_10562,N_2938,N_5846);
and U10563 (N_10563,N_5003,N_235);
and U10564 (N_10564,N_1101,N_3985);
and U10565 (N_10565,N_5370,N_5092);
xnor U10566 (N_10566,N_2378,N_297);
xor U10567 (N_10567,N_2754,N_2893);
nand U10568 (N_10568,N_437,N_1478);
nand U10569 (N_10569,N_5499,N_2903);
nor U10570 (N_10570,N_1398,N_4792);
xnor U10571 (N_10571,N_2205,N_819);
nor U10572 (N_10572,N_1980,N_1545);
nor U10573 (N_10573,N_622,N_1762);
or U10574 (N_10574,N_3185,N_388);
and U10575 (N_10575,N_4230,N_366);
xnor U10576 (N_10576,N_2945,N_2861);
xnor U10577 (N_10577,N_57,N_3039);
and U10578 (N_10578,N_3108,N_2501);
xor U10579 (N_10579,N_3208,N_5560);
xnor U10580 (N_10580,N_704,N_1875);
nor U10581 (N_10581,N_2839,N_4680);
or U10582 (N_10582,N_2593,N_3006);
nand U10583 (N_10583,N_2279,N_5220);
or U10584 (N_10584,N_610,N_5446);
nand U10585 (N_10585,N_3741,N_3812);
nor U10586 (N_10586,N_2001,N_4051);
and U10587 (N_10587,N_2353,N_23);
xor U10588 (N_10588,N_3266,N_5889);
nor U10589 (N_10589,N_1875,N_97);
or U10590 (N_10590,N_507,N_2545);
or U10591 (N_10591,N_5966,N_5842);
nor U10592 (N_10592,N_3183,N_4488);
and U10593 (N_10593,N_2160,N_1188);
nand U10594 (N_10594,N_6036,N_1470);
or U10595 (N_10595,N_1357,N_1709);
and U10596 (N_10596,N_4705,N_2632);
nor U10597 (N_10597,N_278,N_1178);
nand U10598 (N_10598,N_1712,N_1242);
xnor U10599 (N_10599,N_2737,N_3852);
nand U10600 (N_10600,N_2993,N_1522);
nand U10601 (N_10601,N_5563,N_1447);
and U10602 (N_10602,N_5416,N_3423);
nand U10603 (N_10603,N_4695,N_5624);
nor U10604 (N_10604,N_5433,N_5521);
nor U10605 (N_10605,N_3978,N_1846);
nand U10606 (N_10606,N_2359,N_4669);
and U10607 (N_10607,N_2789,N_5499);
or U10608 (N_10608,N_4231,N_4377);
xor U10609 (N_10609,N_5896,N_5515);
or U10610 (N_10610,N_5246,N_2881);
and U10611 (N_10611,N_5824,N_5339);
nand U10612 (N_10612,N_4322,N_4532);
and U10613 (N_10613,N_5062,N_4145);
and U10614 (N_10614,N_5312,N_4313);
or U10615 (N_10615,N_5264,N_1440);
nor U10616 (N_10616,N_3053,N_4624);
or U10617 (N_10617,N_2636,N_6114);
or U10618 (N_10618,N_3691,N_5677);
or U10619 (N_10619,N_3464,N_2186);
and U10620 (N_10620,N_319,N_2836);
xor U10621 (N_10621,N_3295,N_4765);
nor U10622 (N_10622,N_880,N_4466);
xor U10623 (N_10623,N_3925,N_3502);
or U10624 (N_10624,N_2108,N_2309);
and U10625 (N_10625,N_4385,N_1583);
xor U10626 (N_10626,N_5574,N_3090);
or U10627 (N_10627,N_5184,N_3666);
xor U10628 (N_10628,N_4076,N_2830);
and U10629 (N_10629,N_2163,N_2907);
xnor U10630 (N_10630,N_5671,N_1303);
and U10631 (N_10631,N_5896,N_2383);
or U10632 (N_10632,N_5501,N_1108);
nand U10633 (N_10633,N_2162,N_432);
nor U10634 (N_10634,N_3782,N_1158);
nand U10635 (N_10635,N_1709,N_3081);
nand U10636 (N_10636,N_5089,N_4993);
or U10637 (N_10637,N_4026,N_4482);
nor U10638 (N_10638,N_3451,N_4958);
and U10639 (N_10639,N_1924,N_4820);
and U10640 (N_10640,N_5185,N_1092);
nor U10641 (N_10641,N_4238,N_1741);
and U10642 (N_10642,N_1621,N_4770);
xnor U10643 (N_10643,N_4982,N_5848);
or U10644 (N_10644,N_445,N_58);
or U10645 (N_10645,N_617,N_1540);
nor U10646 (N_10646,N_503,N_1632);
nor U10647 (N_10647,N_279,N_985);
xnor U10648 (N_10648,N_5908,N_2180);
xnor U10649 (N_10649,N_1061,N_4012);
nor U10650 (N_10650,N_5524,N_1436);
and U10651 (N_10651,N_5538,N_237);
and U10652 (N_10652,N_867,N_5438);
or U10653 (N_10653,N_3767,N_6027);
nor U10654 (N_10654,N_5328,N_4289);
nand U10655 (N_10655,N_5926,N_2882);
or U10656 (N_10656,N_3545,N_6220);
nor U10657 (N_10657,N_3454,N_668);
xnor U10658 (N_10658,N_5612,N_5658);
xor U10659 (N_10659,N_2231,N_4177);
and U10660 (N_10660,N_3736,N_667);
nor U10661 (N_10661,N_3026,N_2111);
and U10662 (N_10662,N_3823,N_5442);
or U10663 (N_10663,N_497,N_458);
nand U10664 (N_10664,N_20,N_1950);
xor U10665 (N_10665,N_5595,N_3185);
or U10666 (N_10666,N_4256,N_2306);
nor U10667 (N_10667,N_5811,N_311);
nor U10668 (N_10668,N_1753,N_3379);
xnor U10669 (N_10669,N_2843,N_3643);
xnor U10670 (N_10670,N_2132,N_4122);
and U10671 (N_10671,N_1307,N_4614);
nand U10672 (N_10672,N_2198,N_2194);
nor U10673 (N_10673,N_1406,N_1576);
or U10674 (N_10674,N_1294,N_5492);
and U10675 (N_10675,N_1720,N_1581);
or U10676 (N_10676,N_2942,N_3246);
xor U10677 (N_10677,N_2580,N_5783);
xor U10678 (N_10678,N_5372,N_4859);
nor U10679 (N_10679,N_4072,N_495);
nand U10680 (N_10680,N_3723,N_3408);
nand U10681 (N_10681,N_3405,N_2981);
or U10682 (N_10682,N_4388,N_5511);
and U10683 (N_10683,N_1732,N_5181);
nor U10684 (N_10684,N_6091,N_1289);
or U10685 (N_10685,N_1778,N_1624);
and U10686 (N_10686,N_2019,N_2261);
xor U10687 (N_10687,N_399,N_192);
and U10688 (N_10688,N_4488,N_256);
or U10689 (N_10689,N_4523,N_5762);
and U10690 (N_10690,N_3412,N_3257);
nor U10691 (N_10691,N_2660,N_3934);
and U10692 (N_10692,N_924,N_3953);
and U10693 (N_10693,N_5534,N_4047);
and U10694 (N_10694,N_2220,N_3190);
xnor U10695 (N_10695,N_673,N_4782);
nand U10696 (N_10696,N_305,N_4812);
nor U10697 (N_10697,N_1789,N_1768);
and U10698 (N_10698,N_5081,N_5588);
nand U10699 (N_10699,N_397,N_5678);
xor U10700 (N_10700,N_4201,N_2899);
xnor U10701 (N_10701,N_2209,N_4508);
nand U10702 (N_10702,N_4324,N_146);
nor U10703 (N_10703,N_393,N_5053);
and U10704 (N_10704,N_2479,N_4983);
xor U10705 (N_10705,N_1525,N_3157);
nor U10706 (N_10706,N_6044,N_4327);
nand U10707 (N_10707,N_4971,N_2289);
nor U10708 (N_10708,N_2186,N_526);
xor U10709 (N_10709,N_3369,N_951);
xor U10710 (N_10710,N_5763,N_6002);
nand U10711 (N_10711,N_877,N_6152);
nand U10712 (N_10712,N_1074,N_1834);
nor U10713 (N_10713,N_3280,N_1680);
nor U10714 (N_10714,N_1032,N_5637);
xor U10715 (N_10715,N_3941,N_1184);
nand U10716 (N_10716,N_1193,N_974);
or U10717 (N_10717,N_2466,N_3370);
xnor U10718 (N_10718,N_4527,N_3516);
and U10719 (N_10719,N_4488,N_3042);
and U10720 (N_10720,N_1031,N_126);
or U10721 (N_10721,N_1556,N_5167);
xnor U10722 (N_10722,N_4733,N_4076);
nand U10723 (N_10723,N_1946,N_4868);
nand U10724 (N_10724,N_1741,N_3964);
xor U10725 (N_10725,N_1608,N_5994);
xor U10726 (N_10726,N_6083,N_60);
or U10727 (N_10727,N_2016,N_5436);
and U10728 (N_10728,N_2699,N_1947);
and U10729 (N_10729,N_4656,N_1085);
or U10730 (N_10730,N_401,N_2451);
and U10731 (N_10731,N_3139,N_5046);
xor U10732 (N_10732,N_1160,N_5740);
or U10733 (N_10733,N_5644,N_4043);
and U10734 (N_10734,N_518,N_5518);
or U10735 (N_10735,N_5790,N_3013);
nor U10736 (N_10736,N_3509,N_3310);
nor U10737 (N_10737,N_4419,N_1809);
nand U10738 (N_10738,N_2844,N_768);
or U10739 (N_10739,N_2567,N_3109);
and U10740 (N_10740,N_3401,N_5826);
and U10741 (N_10741,N_425,N_2408);
and U10742 (N_10742,N_5866,N_5515);
nand U10743 (N_10743,N_1033,N_3809);
xor U10744 (N_10744,N_4119,N_1611);
nor U10745 (N_10745,N_4200,N_5034);
and U10746 (N_10746,N_1506,N_3439);
xnor U10747 (N_10747,N_1014,N_953);
xnor U10748 (N_10748,N_2717,N_1488);
or U10749 (N_10749,N_4182,N_966);
nand U10750 (N_10750,N_500,N_1159);
and U10751 (N_10751,N_811,N_3003);
and U10752 (N_10752,N_555,N_5431);
or U10753 (N_10753,N_2147,N_3207);
and U10754 (N_10754,N_4380,N_593);
nand U10755 (N_10755,N_4528,N_174);
and U10756 (N_10756,N_4793,N_109);
and U10757 (N_10757,N_4179,N_1838);
or U10758 (N_10758,N_3539,N_1899);
or U10759 (N_10759,N_5178,N_3569);
nor U10760 (N_10760,N_143,N_94);
and U10761 (N_10761,N_6143,N_1206);
xnor U10762 (N_10762,N_5370,N_3204);
nand U10763 (N_10763,N_869,N_1378);
or U10764 (N_10764,N_3734,N_2112);
xnor U10765 (N_10765,N_5370,N_5673);
xnor U10766 (N_10766,N_881,N_4013);
nor U10767 (N_10767,N_2384,N_5548);
nand U10768 (N_10768,N_2273,N_5036);
or U10769 (N_10769,N_1821,N_636);
and U10770 (N_10770,N_728,N_155);
nand U10771 (N_10771,N_4526,N_2196);
nand U10772 (N_10772,N_3904,N_2702);
or U10773 (N_10773,N_5170,N_4949);
xor U10774 (N_10774,N_5679,N_2911);
nor U10775 (N_10775,N_2962,N_3438);
and U10776 (N_10776,N_3888,N_4632);
and U10777 (N_10777,N_5262,N_1590);
or U10778 (N_10778,N_2546,N_3895);
nor U10779 (N_10779,N_809,N_1790);
nor U10780 (N_10780,N_2541,N_6125);
or U10781 (N_10781,N_1114,N_6129);
or U10782 (N_10782,N_4190,N_4873);
or U10783 (N_10783,N_706,N_5234);
xnor U10784 (N_10784,N_2134,N_2112);
nand U10785 (N_10785,N_864,N_2510);
nor U10786 (N_10786,N_5813,N_4901);
nor U10787 (N_10787,N_3237,N_6121);
and U10788 (N_10788,N_3740,N_565);
nor U10789 (N_10789,N_2698,N_2441);
or U10790 (N_10790,N_5490,N_1170);
and U10791 (N_10791,N_4107,N_2028);
and U10792 (N_10792,N_2070,N_149);
xnor U10793 (N_10793,N_1577,N_3772);
xnor U10794 (N_10794,N_2530,N_5367);
xor U10795 (N_10795,N_3273,N_3442);
and U10796 (N_10796,N_268,N_5267);
nand U10797 (N_10797,N_6072,N_4737);
or U10798 (N_10798,N_5092,N_185);
xnor U10799 (N_10799,N_5087,N_5775);
xnor U10800 (N_10800,N_3843,N_5000);
or U10801 (N_10801,N_2783,N_296);
nand U10802 (N_10802,N_1660,N_2950);
nand U10803 (N_10803,N_4196,N_979);
nor U10804 (N_10804,N_1233,N_5436);
nand U10805 (N_10805,N_631,N_949);
or U10806 (N_10806,N_4902,N_1438);
nor U10807 (N_10807,N_3642,N_5796);
and U10808 (N_10808,N_2195,N_4329);
nor U10809 (N_10809,N_2632,N_5057);
nand U10810 (N_10810,N_5632,N_4378);
or U10811 (N_10811,N_1901,N_70);
xor U10812 (N_10812,N_6171,N_2678);
xor U10813 (N_10813,N_5521,N_4727);
nor U10814 (N_10814,N_5177,N_3866);
nor U10815 (N_10815,N_1517,N_5352);
nor U10816 (N_10816,N_6039,N_3236);
and U10817 (N_10817,N_5151,N_3908);
and U10818 (N_10818,N_1647,N_1227);
or U10819 (N_10819,N_109,N_3835);
and U10820 (N_10820,N_141,N_5006);
xor U10821 (N_10821,N_2248,N_3247);
and U10822 (N_10822,N_4558,N_6120);
and U10823 (N_10823,N_1877,N_2605);
and U10824 (N_10824,N_678,N_668);
xnor U10825 (N_10825,N_2813,N_2788);
and U10826 (N_10826,N_1871,N_5201);
nor U10827 (N_10827,N_3851,N_248);
nor U10828 (N_10828,N_3057,N_2073);
and U10829 (N_10829,N_690,N_1446);
xor U10830 (N_10830,N_1043,N_5898);
or U10831 (N_10831,N_2042,N_3400);
nand U10832 (N_10832,N_5287,N_1107);
and U10833 (N_10833,N_323,N_439);
or U10834 (N_10834,N_4866,N_1342);
nand U10835 (N_10835,N_4921,N_4441);
or U10836 (N_10836,N_4686,N_2027);
nor U10837 (N_10837,N_643,N_1363);
nor U10838 (N_10838,N_5745,N_5436);
nand U10839 (N_10839,N_2279,N_4805);
or U10840 (N_10840,N_5720,N_5351);
and U10841 (N_10841,N_1640,N_2844);
nand U10842 (N_10842,N_3622,N_2256);
xnor U10843 (N_10843,N_3758,N_762);
and U10844 (N_10844,N_316,N_163);
nand U10845 (N_10845,N_452,N_2737);
nor U10846 (N_10846,N_1253,N_2375);
nand U10847 (N_10847,N_1691,N_4700);
nand U10848 (N_10848,N_4558,N_2632);
xnor U10849 (N_10849,N_240,N_5930);
and U10850 (N_10850,N_4384,N_4806);
nor U10851 (N_10851,N_244,N_2782);
nor U10852 (N_10852,N_3899,N_5409);
and U10853 (N_10853,N_6003,N_1196);
nor U10854 (N_10854,N_2086,N_308);
xor U10855 (N_10855,N_175,N_2581);
and U10856 (N_10856,N_4949,N_4409);
nand U10857 (N_10857,N_101,N_717);
and U10858 (N_10858,N_4972,N_56);
nor U10859 (N_10859,N_4196,N_562);
and U10860 (N_10860,N_5506,N_1447);
nor U10861 (N_10861,N_1289,N_2779);
or U10862 (N_10862,N_1687,N_1879);
and U10863 (N_10863,N_913,N_4525);
nand U10864 (N_10864,N_1725,N_1520);
or U10865 (N_10865,N_2234,N_5597);
nor U10866 (N_10866,N_3414,N_302);
xnor U10867 (N_10867,N_3940,N_1831);
nor U10868 (N_10868,N_2905,N_6175);
or U10869 (N_10869,N_3984,N_3740);
nor U10870 (N_10870,N_3330,N_3506);
or U10871 (N_10871,N_562,N_4535);
or U10872 (N_10872,N_4262,N_1186);
xor U10873 (N_10873,N_6076,N_1460);
or U10874 (N_10874,N_1402,N_4094);
xnor U10875 (N_10875,N_5318,N_5710);
and U10876 (N_10876,N_1354,N_526);
nand U10877 (N_10877,N_5291,N_963);
xnor U10878 (N_10878,N_1301,N_1338);
xnor U10879 (N_10879,N_1095,N_4917);
xor U10880 (N_10880,N_2384,N_1579);
and U10881 (N_10881,N_272,N_324);
or U10882 (N_10882,N_4187,N_3516);
or U10883 (N_10883,N_5174,N_1999);
or U10884 (N_10884,N_4753,N_1907);
xnor U10885 (N_10885,N_2453,N_3312);
or U10886 (N_10886,N_3811,N_4975);
nand U10887 (N_10887,N_389,N_6106);
nor U10888 (N_10888,N_6068,N_4300);
or U10889 (N_10889,N_223,N_2072);
or U10890 (N_10890,N_6012,N_4949);
or U10891 (N_10891,N_4486,N_808);
nand U10892 (N_10892,N_2383,N_2737);
xnor U10893 (N_10893,N_2080,N_2163);
xnor U10894 (N_10894,N_747,N_3512);
nand U10895 (N_10895,N_3346,N_3924);
nor U10896 (N_10896,N_2448,N_3949);
nand U10897 (N_10897,N_2061,N_1004);
or U10898 (N_10898,N_4055,N_5904);
nor U10899 (N_10899,N_2377,N_5672);
or U10900 (N_10900,N_2682,N_2579);
and U10901 (N_10901,N_2195,N_2525);
nor U10902 (N_10902,N_3276,N_3592);
nand U10903 (N_10903,N_5499,N_1275);
xnor U10904 (N_10904,N_2773,N_3455);
xnor U10905 (N_10905,N_5145,N_98);
xor U10906 (N_10906,N_149,N_1384);
nand U10907 (N_10907,N_5340,N_1321);
nor U10908 (N_10908,N_4993,N_901);
nand U10909 (N_10909,N_2397,N_3699);
nor U10910 (N_10910,N_6045,N_1672);
nor U10911 (N_10911,N_6068,N_1043);
nand U10912 (N_10912,N_368,N_2433);
or U10913 (N_10913,N_4259,N_5153);
nor U10914 (N_10914,N_865,N_2426);
xor U10915 (N_10915,N_375,N_4653);
xnor U10916 (N_10916,N_3812,N_2780);
or U10917 (N_10917,N_2913,N_4875);
nor U10918 (N_10918,N_935,N_4892);
xnor U10919 (N_10919,N_2773,N_5970);
and U10920 (N_10920,N_5336,N_4395);
nand U10921 (N_10921,N_13,N_1860);
and U10922 (N_10922,N_3277,N_1244);
and U10923 (N_10923,N_242,N_4211);
xnor U10924 (N_10924,N_6184,N_5814);
nor U10925 (N_10925,N_639,N_4360);
nand U10926 (N_10926,N_244,N_3732);
and U10927 (N_10927,N_4460,N_1949);
and U10928 (N_10928,N_2932,N_2128);
nand U10929 (N_10929,N_6198,N_5985);
xnor U10930 (N_10930,N_1566,N_5382);
nor U10931 (N_10931,N_3283,N_4572);
nor U10932 (N_10932,N_4264,N_3797);
nor U10933 (N_10933,N_113,N_2812);
nor U10934 (N_10934,N_3779,N_5420);
and U10935 (N_10935,N_6172,N_3390);
xor U10936 (N_10936,N_614,N_1055);
xor U10937 (N_10937,N_2026,N_5628);
xnor U10938 (N_10938,N_717,N_1554);
xor U10939 (N_10939,N_4526,N_4960);
xnor U10940 (N_10940,N_4593,N_1169);
xnor U10941 (N_10941,N_10,N_5107);
nor U10942 (N_10942,N_4316,N_2784);
and U10943 (N_10943,N_2209,N_4950);
nor U10944 (N_10944,N_3044,N_4994);
xor U10945 (N_10945,N_3274,N_1139);
nor U10946 (N_10946,N_2696,N_1096);
nand U10947 (N_10947,N_4005,N_628);
xor U10948 (N_10948,N_1243,N_5162);
or U10949 (N_10949,N_1964,N_2644);
xnor U10950 (N_10950,N_172,N_1365);
or U10951 (N_10951,N_5759,N_4331);
and U10952 (N_10952,N_2921,N_5327);
nand U10953 (N_10953,N_3624,N_6209);
and U10954 (N_10954,N_884,N_2907);
and U10955 (N_10955,N_3321,N_3685);
nor U10956 (N_10956,N_4542,N_4653);
and U10957 (N_10957,N_2361,N_1375);
and U10958 (N_10958,N_4867,N_1270);
nand U10959 (N_10959,N_5376,N_3435);
xor U10960 (N_10960,N_3681,N_5538);
nand U10961 (N_10961,N_2634,N_1705);
nand U10962 (N_10962,N_796,N_5408);
xor U10963 (N_10963,N_304,N_6078);
xnor U10964 (N_10964,N_256,N_1207);
nor U10965 (N_10965,N_3675,N_3111);
nand U10966 (N_10966,N_5432,N_1462);
nor U10967 (N_10967,N_393,N_1849);
nor U10968 (N_10968,N_5173,N_1272);
and U10969 (N_10969,N_2572,N_1047);
nand U10970 (N_10970,N_97,N_6108);
nor U10971 (N_10971,N_2789,N_2954);
or U10972 (N_10972,N_2110,N_4090);
or U10973 (N_10973,N_1290,N_5812);
nor U10974 (N_10974,N_1792,N_3409);
nor U10975 (N_10975,N_5635,N_2571);
nor U10976 (N_10976,N_6230,N_299);
xnor U10977 (N_10977,N_1937,N_5487);
or U10978 (N_10978,N_3055,N_1999);
nor U10979 (N_10979,N_1537,N_5065);
and U10980 (N_10980,N_1277,N_4080);
xnor U10981 (N_10981,N_5316,N_2991);
and U10982 (N_10982,N_5602,N_4610);
xnor U10983 (N_10983,N_4030,N_2680);
or U10984 (N_10984,N_5283,N_5679);
and U10985 (N_10985,N_1501,N_2468);
or U10986 (N_10986,N_2611,N_5568);
or U10987 (N_10987,N_381,N_1186);
and U10988 (N_10988,N_6085,N_1619);
or U10989 (N_10989,N_4300,N_5054);
nor U10990 (N_10990,N_1538,N_1977);
or U10991 (N_10991,N_3517,N_4582);
nor U10992 (N_10992,N_1634,N_5161);
or U10993 (N_10993,N_3214,N_4759);
and U10994 (N_10994,N_4749,N_3634);
xor U10995 (N_10995,N_3161,N_4106);
or U10996 (N_10996,N_3718,N_3846);
nor U10997 (N_10997,N_3862,N_925);
xor U10998 (N_10998,N_457,N_4370);
and U10999 (N_10999,N_5517,N_1280);
nand U11000 (N_11000,N_3953,N_4423);
and U11001 (N_11001,N_5944,N_3513);
xnor U11002 (N_11002,N_6109,N_5068);
xor U11003 (N_11003,N_1766,N_1934);
xnor U11004 (N_11004,N_1289,N_4277);
xnor U11005 (N_11005,N_5263,N_5863);
and U11006 (N_11006,N_5011,N_3321);
and U11007 (N_11007,N_5292,N_3496);
nor U11008 (N_11008,N_986,N_4235);
nand U11009 (N_11009,N_214,N_2721);
nand U11010 (N_11010,N_4575,N_3500);
nand U11011 (N_11011,N_4874,N_5204);
xnor U11012 (N_11012,N_5872,N_4559);
or U11013 (N_11013,N_5096,N_5368);
nand U11014 (N_11014,N_783,N_3008);
nand U11015 (N_11015,N_2403,N_5142);
and U11016 (N_11016,N_2063,N_2758);
or U11017 (N_11017,N_298,N_1322);
or U11018 (N_11018,N_4269,N_1115);
and U11019 (N_11019,N_71,N_3742);
and U11020 (N_11020,N_2175,N_2679);
and U11021 (N_11021,N_266,N_1153);
xor U11022 (N_11022,N_982,N_1642);
nand U11023 (N_11023,N_4995,N_433);
nand U11024 (N_11024,N_48,N_1887);
xnor U11025 (N_11025,N_809,N_32);
nand U11026 (N_11026,N_4875,N_2671);
xor U11027 (N_11027,N_3999,N_4731);
nor U11028 (N_11028,N_5024,N_2135);
and U11029 (N_11029,N_910,N_2039);
nand U11030 (N_11030,N_2915,N_2593);
nor U11031 (N_11031,N_4930,N_1268);
or U11032 (N_11032,N_227,N_3675);
nand U11033 (N_11033,N_4058,N_4014);
nor U11034 (N_11034,N_5647,N_3359);
and U11035 (N_11035,N_2020,N_5376);
xor U11036 (N_11036,N_1261,N_6216);
and U11037 (N_11037,N_5224,N_887);
or U11038 (N_11038,N_5599,N_699);
and U11039 (N_11039,N_5286,N_1569);
xnor U11040 (N_11040,N_5592,N_4626);
and U11041 (N_11041,N_20,N_4161);
nand U11042 (N_11042,N_152,N_1096);
or U11043 (N_11043,N_2279,N_3123);
and U11044 (N_11044,N_3575,N_4531);
nand U11045 (N_11045,N_4226,N_914);
or U11046 (N_11046,N_3509,N_5683);
xnor U11047 (N_11047,N_1760,N_401);
or U11048 (N_11048,N_6143,N_2308);
and U11049 (N_11049,N_4296,N_3940);
or U11050 (N_11050,N_5000,N_3061);
nand U11051 (N_11051,N_2434,N_5971);
xnor U11052 (N_11052,N_3747,N_1838);
or U11053 (N_11053,N_1198,N_352);
xnor U11054 (N_11054,N_2342,N_3764);
xor U11055 (N_11055,N_5451,N_4738);
xor U11056 (N_11056,N_1733,N_1232);
or U11057 (N_11057,N_1014,N_3842);
nand U11058 (N_11058,N_4964,N_5999);
nor U11059 (N_11059,N_2199,N_272);
nor U11060 (N_11060,N_2048,N_14);
nand U11061 (N_11061,N_4989,N_2816);
nor U11062 (N_11062,N_5646,N_1684);
nand U11063 (N_11063,N_3409,N_2544);
and U11064 (N_11064,N_2793,N_3849);
nand U11065 (N_11065,N_588,N_5053);
xnor U11066 (N_11066,N_5984,N_5736);
nor U11067 (N_11067,N_5767,N_5999);
xor U11068 (N_11068,N_2476,N_4691);
xor U11069 (N_11069,N_681,N_5248);
xor U11070 (N_11070,N_1350,N_202);
nand U11071 (N_11071,N_5001,N_1831);
or U11072 (N_11072,N_5790,N_5144);
nand U11073 (N_11073,N_4108,N_497);
nor U11074 (N_11074,N_5956,N_1463);
nand U11075 (N_11075,N_1820,N_1139);
nand U11076 (N_11076,N_5841,N_4671);
or U11077 (N_11077,N_1330,N_2158);
nor U11078 (N_11078,N_5822,N_2831);
nor U11079 (N_11079,N_3843,N_2314);
xnor U11080 (N_11080,N_656,N_1579);
and U11081 (N_11081,N_4347,N_2869);
nand U11082 (N_11082,N_2909,N_5581);
or U11083 (N_11083,N_1925,N_3149);
or U11084 (N_11084,N_6201,N_1701);
xnor U11085 (N_11085,N_3133,N_3478);
and U11086 (N_11086,N_309,N_481);
nand U11087 (N_11087,N_3102,N_1385);
nand U11088 (N_11088,N_3605,N_1480);
nor U11089 (N_11089,N_2021,N_1831);
nor U11090 (N_11090,N_472,N_3676);
nand U11091 (N_11091,N_4377,N_2205);
xor U11092 (N_11092,N_395,N_4605);
or U11093 (N_11093,N_3348,N_3562);
nand U11094 (N_11094,N_1169,N_2142);
xor U11095 (N_11095,N_3119,N_1022);
nand U11096 (N_11096,N_2146,N_3441);
or U11097 (N_11097,N_204,N_1359);
and U11098 (N_11098,N_6240,N_4460);
or U11099 (N_11099,N_3986,N_5472);
nand U11100 (N_11100,N_459,N_1254);
or U11101 (N_11101,N_340,N_1058);
nor U11102 (N_11102,N_984,N_2982);
nand U11103 (N_11103,N_290,N_1154);
and U11104 (N_11104,N_1247,N_3857);
or U11105 (N_11105,N_3057,N_5131);
or U11106 (N_11106,N_5019,N_5893);
or U11107 (N_11107,N_5925,N_2536);
nor U11108 (N_11108,N_4937,N_1318);
or U11109 (N_11109,N_2857,N_2134);
or U11110 (N_11110,N_1266,N_6167);
or U11111 (N_11111,N_3461,N_4645);
nand U11112 (N_11112,N_879,N_2643);
and U11113 (N_11113,N_4646,N_5156);
xnor U11114 (N_11114,N_5973,N_2241);
nor U11115 (N_11115,N_2814,N_5383);
xnor U11116 (N_11116,N_1058,N_3427);
nand U11117 (N_11117,N_415,N_3785);
and U11118 (N_11118,N_5993,N_3122);
nor U11119 (N_11119,N_729,N_3800);
or U11120 (N_11120,N_1021,N_3759);
nand U11121 (N_11121,N_1028,N_3565);
xor U11122 (N_11122,N_6204,N_837);
nand U11123 (N_11123,N_4453,N_1137);
nand U11124 (N_11124,N_3127,N_302);
or U11125 (N_11125,N_2549,N_3992);
xor U11126 (N_11126,N_4516,N_6028);
nor U11127 (N_11127,N_944,N_6218);
and U11128 (N_11128,N_4410,N_4213);
xnor U11129 (N_11129,N_3122,N_4429);
xnor U11130 (N_11130,N_270,N_3982);
nor U11131 (N_11131,N_1322,N_891);
nor U11132 (N_11132,N_3291,N_1454);
nand U11133 (N_11133,N_170,N_662);
or U11134 (N_11134,N_286,N_5559);
or U11135 (N_11135,N_6189,N_1896);
nand U11136 (N_11136,N_3715,N_4336);
xnor U11137 (N_11137,N_30,N_5857);
and U11138 (N_11138,N_5775,N_5859);
xor U11139 (N_11139,N_2071,N_3211);
nand U11140 (N_11140,N_4950,N_1778);
or U11141 (N_11141,N_2432,N_3638);
or U11142 (N_11142,N_4736,N_2801);
nor U11143 (N_11143,N_2251,N_5287);
nand U11144 (N_11144,N_2259,N_1962);
xor U11145 (N_11145,N_3694,N_4239);
nor U11146 (N_11146,N_2707,N_3521);
nand U11147 (N_11147,N_3188,N_4785);
nand U11148 (N_11148,N_3565,N_543);
nand U11149 (N_11149,N_5783,N_905);
xor U11150 (N_11150,N_6055,N_1831);
xor U11151 (N_11151,N_2164,N_2523);
nor U11152 (N_11152,N_6123,N_5740);
nand U11153 (N_11153,N_5301,N_744);
xor U11154 (N_11154,N_649,N_3821);
xor U11155 (N_11155,N_1473,N_3154);
xor U11156 (N_11156,N_2376,N_1927);
nand U11157 (N_11157,N_6161,N_1218);
and U11158 (N_11158,N_1936,N_1688);
and U11159 (N_11159,N_1792,N_4492);
xnor U11160 (N_11160,N_3036,N_2061);
and U11161 (N_11161,N_4225,N_4208);
and U11162 (N_11162,N_905,N_3961);
and U11163 (N_11163,N_3031,N_1969);
or U11164 (N_11164,N_1250,N_6025);
and U11165 (N_11165,N_3725,N_3026);
and U11166 (N_11166,N_984,N_4893);
and U11167 (N_11167,N_2154,N_2102);
xnor U11168 (N_11168,N_3927,N_4200);
nand U11169 (N_11169,N_423,N_2393);
or U11170 (N_11170,N_39,N_565);
nor U11171 (N_11171,N_3497,N_4236);
nor U11172 (N_11172,N_3507,N_5350);
or U11173 (N_11173,N_2405,N_5176);
and U11174 (N_11174,N_1994,N_717);
nand U11175 (N_11175,N_2196,N_2190);
nor U11176 (N_11176,N_2459,N_1438);
xnor U11177 (N_11177,N_5374,N_3823);
or U11178 (N_11178,N_3752,N_296);
nand U11179 (N_11179,N_3433,N_3404);
and U11180 (N_11180,N_5332,N_2437);
nand U11181 (N_11181,N_5329,N_3234);
xor U11182 (N_11182,N_5532,N_4478);
and U11183 (N_11183,N_3005,N_4220);
nand U11184 (N_11184,N_1827,N_4682);
or U11185 (N_11185,N_2690,N_5642);
xor U11186 (N_11186,N_5288,N_3065);
xor U11187 (N_11187,N_1668,N_1233);
nor U11188 (N_11188,N_276,N_2516);
and U11189 (N_11189,N_2032,N_697);
xnor U11190 (N_11190,N_4963,N_1070);
or U11191 (N_11191,N_5962,N_1286);
or U11192 (N_11192,N_2179,N_2424);
nor U11193 (N_11193,N_2895,N_1012);
nand U11194 (N_11194,N_995,N_2708);
or U11195 (N_11195,N_3980,N_427);
nor U11196 (N_11196,N_4947,N_3263);
nor U11197 (N_11197,N_3365,N_5101);
nor U11198 (N_11198,N_994,N_3806);
nand U11199 (N_11199,N_5831,N_3774);
or U11200 (N_11200,N_476,N_2811);
nor U11201 (N_11201,N_3694,N_5205);
and U11202 (N_11202,N_2382,N_4027);
nand U11203 (N_11203,N_319,N_3017);
nor U11204 (N_11204,N_1173,N_5023);
xnor U11205 (N_11205,N_3291,N_2272);
or U11206 (N_11206,N_5047,N_3120);
or U11207 (N_11207,N_4562,N_3169);
nand U11208 (N_11208,N_4810,N_1560);
and U11209 (N_11209,N_5120,N_2891);
nand U11210 (N_11210,N_407,N_3348);
xor U11211 (N_11211,N_4385,N_1642);
or U11212 (N_11212,N_3522,N_3761);
nor U11213 (N_11213,N_4630,N_2991);
nor U11214 (N_11214,N_3121,N_481);
and U11215 (N_11215,N_3523,N_1589);
and U11216 (N_11216,N_5480,N_1702);
and U11217 (N_11217,N_4886,N_1882);
and U11218 (N_11218,N_2107,N_5047);
and U11219 (N_11219,N_4305,N_3971);
and U11220 (N_11220,N_1398,N_3099);
nand U11221 (N_11221,N_4521,N_1796);
or U11222 (N_11222,N_3417,N_1535);
or U11223 (N_11223,N_1498,N_1489);
nand U11224 (N_11224,N_1357,N_5484);
and U11225 (N_11225,N_62,N_5183);
and U11226 (N_11226,N_141,N_3094);
xor U11227 (N_11227,N_1273,N_274);
and U11228 (N_11228,N_5814,N_4947);
xor U11229 (N_11229,N_2640,N_515);
nand U11230 (N_11230,N_1588,N_6044);
nand U11231 (N_11231,N_4054,N_4926);
and U11232 (N_11232,N_1962,N_2606);
xnor U11233 (N_11233,N_2110,N_4997);
nand U11234 (N_11234,N_1311,N_4586);
nor U11235 (N_11235,N_5995,N_5512);
nand U11236 (N_11236,N_5449,N_6181);
nand U11237 (N_11237,N_2904,N_3306);
xnor U11238 (N_11238,N_2489,N_3412);
and U11239 (N_11239,N_6224,N_1993);
or U11240 (N_11240,N_4497,N_4241);
and U11241 (N_11241,N_2430,N_925);
xnor U11242 (N_11242,N_2793,N_3230);
and U11243 (N_11243,N_4030,N_2858);
nand U11244 (N_11244,N_2454,N_2411);
nand U11245 (N_11245,N_4282,N_2974);
or U11246 (N_11246,N_5785,N_4867);
xnor U11247 (N_11247,N_5686,N_2968);
nor U11248 (N_11248,N_1881,N_4322);
nor U11249 (N_11249,N_5816,N_2986);
nand U11250 (N_11250,N_2949,N_3037);
nor U11251 (N_11251,N_230,N_5374);
nand U11252 (N_11252,N_5747,N_6051);
xnor U11253 (N_11253,N_2547,N_5275);
xnor U11254 (N_11254,N_2652,N_6123);
and U11255 (N_11255,N_3287,N_5907);
and U11256 (N_11256,N_5763,N_2515);
or U11257 (N_11257,N_5453,N_3035);
nor U11258 (N_11258,N_186,N_637);
nand U11259 (N_11259,N_3855,N_180);
xnor U11260 (N_11260,N_3172,N_5442);
nand U11261 (N_11261,N_6077,N_4643);
xnor U11262 (N_11262,N_475,N_2342);
or U11263 (N_11263,N_504,N_4878);
xnor U11264 (N_11264,N_39,N_5867);
and U11265 (N_11265,N_5024,N_4696);
xor U11266 (N_11266,N_677,N_668);
and U11267 (N_11267,N_615,N_1469);
or U11268 (N_11268,N_900,N_1197);
or U11269 (N_11269,N_4607,N_3909);
nor U11270 (N_11270,N_2050,N_3451);
nand U11271 (N_11271,N_101,N_324);
nand U11272 (N_11272,N_3830,N_2537);
nand U11273 (N_11273,N_650,N_4667);
nand U11274 (N_11274,N_21,N_4289);
xnor U11275 (N_11275,N_5703,N_4907);
or U11276 (N_11276,N_4723,N_1124);
and U11277 (N_11277,N_479,N_2368);
nand U11278 (N_11278,N_5754,N_5394);
xor U11279 (N_11279,N_907,N_20);
nor U11280 (N_11280,N_5390,N_1894);
and U11281 (N_11281,N_3467,N_3089);
nand U11282 (N_11282,N_3140,N_3269);
and U11283 (N_11283,N_3361,N_631);
xor U11284 (N_11284,N_3105,N_5558);
or U11285 (N_11285,N_2226,N_6048);
and U11286 (N_11286,N_1344,N_1007);
nand U11287 (N_11287,N_3366,N_4537);
nand U11288 (N_11288,N_5692,N_2395);
and U11289 (N_11289,N_5940,N_2762);
and U11290 (N_11290,N_738,N_846);
and U11291 (N_11291,N_1164,N_1724);
and U11292 (N_11292,N_5279,N_5445);
nor U11293 (N_11293,N_3832,N_2524);
xor U11294 (N_11294,N_4046,N_5146);
xor U11295 (N_11295,N_3235,N_2621);
nand U11296 (N_11296,N_1396,N_1926);
xnor U11297 (N_11297,N_4897,N_1759);
and U11298 (N_11298,N_427,N_5812);
or U11299 (N_11299,N_1306,N_1360);
nand U11300 (N_11300,N_6082,N_6039);
nand U11301 (N_11301,N_5388,N_1690);
or U11302 (N_11302,N_5330,N_5201);
or U11303 (N_11303,N_790,N_87);
nand U11304 (N_11304,N_2317,N_742);
nand U11305 (N_11305,N_3661,N_1068);
xor U11306 (N_11306,N_762,N_3381);
nor U11307 (N_11307,N_4704,N_733);
nor U11308 (N_11308,N_2244,N_3338);
nand U11309 (N_11309,N_441,N_5589);
nand U11310 (N_11310,N_262,N_2370);
nand U11311 (N_11311,N_1812,N_3610);
xnor U11312 (N_11312,N_3371,N_2404);
xor U11313 (N_11313,N_5007,N_4342);
or U11314 (N_11314,N_2506,N_3594);
or U11315 (N_11315,N_6008,N_6218);
and U11316 (N_11316,N_5782,N_3399);
xor U11317 (N_11317,N_5260,N_4289);
and U11318 (N_11318,N_4171,N_5694);
or U11319 (N_11319,N_2231,N_1833);
or U11320 (N_11320,N_704,N_158);
nor U11321 (N_11321,N_848,N_3772);
nand U11322 (N_11322,N_4248,N_6069);
nand U11323 (N_11323,N_5701,N_5421);
or U11324 (N_11324,N_492,N_795);
xnor U11325 (N_11325,N_1224,N_499);
nand U11326 (N_11326,N_4845,N_4095);
nor U11327 (N_11327,N_1159,N_700);
or U11328 (N_11328,N_6025,N_1680);
or U11329 (N_11329,N_1083,N_4927);
and U11330 (N_11330,N_2106,N_5067);
and U11331 (N_11331,N_1035,N_6154);
or U11332 (N_11332,N_4654,N_5980);
or U11333 (N_11333,N_1338,N_138);
and U11334 (N_11334,N_5379,N_944);
nand U11335 (N_11335,N_970,N_1808);
and U11336 (N_11336,N_902,N_2867);
and U11337 (N_11337,N_5842,N_1160);
xnor U11338 (N_11338,N_2322,N_1885);
and U11339 (N_11339,N_5989,N_4303);
nand U11340 (N_11340,N_4370,N_1919);
nor U11341 (N_11341,N_627,N_6022);
nand U11342 (N_11342,N_337,N_4486);
xor U11343 (N_11343,N_1519,N_4144);
nand U11344 (N_11344,N_2232,N_1695);
or U11345 (N_11345,N_580,N_1333);
nor U11346 (N_11346,N_3963,N_2392);
nor U11347 (N_11347,N_297,N_1435);
and U11348 (N_11348,N_5801,N_45);
xnor U11349 (N_11349,N_3058,N_3745);
nand U11350 (N_11350,N_2620,N_1075);
nor U11351 (N_11351,N_5802,N_3505);
nand U11352 (N_11352,N_599,N_1540);
or U11353 (N_11353,N_2591,N_3047);
or U11354 (N_11354,N_4338,N_3836);
and U11355 (N_11355,N_912,N_565);
xor U11356 (N_11356,N_6163,N_5225);
and U11357 (N_11357,N_2795,N_3519);
nor U11358 (N_11358,N_4551,N_4775);
nor U11359 (N_11359,N_6006,N_2281);
nand U11360 (N_11360,N_956,N_2614);
and U11361 (N_11361,N_1438,N_1907);
xor U11362 (N_11362,N_387,N_2924);
xnor U11363 (N_11363,N_786,N_5528);
and U11364 (N_11364,N_4923,N_5822);
or U11365 (N_11365,N_5771,N_1535);
nand U11366 (N_11366,N_1714,N_787);
and U11367 (N_11367,N_5908,N_2928);
xnor U11368 (N_11368,N_6247,N_1669);
xnor U11369 (N_11369,N_1050,N_2609);
and U11370 (N_11370,N_4082,N_5993);
nor U11371 (N_11371,N_4173,N_4947);
nor U11372 (N_11372,N_259,N_1323);
nor U11373 (N_11373,N_6083,N_4424);
nor U11374 (N_11374,N_3283,N_533);
and U11375 (N_11375,N_2367,N_2278);
xor U11376 (N_11376,N_3593,N_2756);
or U11377 (N_11377,N_4567,N_1888);
and U11378 (N_11378,N_277,N_1094);
nand U11379 (N_11379,N_2539,N_1135);
and U11380 (N_11380,N_2505,N_3976);
xor U11381 (N_11381,N_405,N_1750);
xnor U11382 (N_11382,N_5990,N_2186);
and U11383 (N_11383,N_1878,N_842);
or U11384 (N_11384,N_4967,N_5162);
nor U11385 (N_11385,N_5417,N_2343);
nand U11386 (N_11386,N_4987,N_115);
or U11387 (N_11387,N_480,N_4114);
or U11388 (N_11388,N_3191,N_849);
nor U11389 (N_11389,N_129,N_5827);
nand U11390 (N_11390,N_2715,N_3941);
and U11391 (N_11391,N_5610,N_1376);
nor U11392 (N_11392,N_4182,N_1559);
nor U11393 (N_11393,N_4176,N_4082);
nand U11394 (N_11394,N_1477,N_920);
or U11395 (N_11395,N_6207,N_2888);
and U11396 (N_11396,N_2400,N_5489);
and U11397 (N_11397,N_1787,N_2310);
and U11398 (N_11398,N_5038,N_5072);
xnor U11399 (N_11399,N_5801,N_1922);
nand U11400 (N_11400,N_2623,N_2711);
or U11401 (N_11401,N_2909,N_992);
and U11402 (N_11402,N_6102,N_2862);
and U11403 (N_11403,N_234,N_4989);
and U11404 (N_11404,N_2176,N_4004);
nand U11405 (N_11405,N_50,N_3975);
nor U11406 (N_11406,N_4716,N_5029);
nor U11407 (N_11407,N_5804,N_225);
or U11408 (N_11408,N_4204,N_2052);
nor U11409 (N_11409,N_1465,N_4344);
xor U11410 (N_11410,N_19,N_4427);
and U11411 (N_11411,N_3599,N_1639);
nor U11412 (N_11412,N_4248,N_5041);
nand U11413 (N_11413,N_3611,N_5526);
or U11414 (N_11414,N_689,N_4300);
xnor U11415 (N_11415,N_286,N_5726);
and U11416 (N_11416,N_1562,N_224);
nor U11417 (N_11417,N_5529,N_5630);
and U11418 (N_11418,N_322,N_3404);
xnor U11419 (N_11419,N_3329,N_5913);
nand U11420 (N_11420,N_3932,N_1719);
or U11421 (N_11421,N_4654,N_184);
xnor U11422 (N_11422,N_1395,N_1926);
xor U11423 (N_11423,N_3589,N_4328);
nor U11424 (N_11424,N_1597,N_5571);
nor U11425 (N_11425,N_1231,N_3455);
and U11426 (N_11426,N_3266,N_668);
and U11427 (N_11427,N_3953,N_4907);
or U11428 (N_11428,N_4411,N_4496);
or U11429 (N_11429,N_2903,N_1955);
nand U11430 (N_11430,N_151,N_5083);
or U11431 (N_11431,N_5415,N_5531);
or U11432 (N_11432,N_3247,N_2869);
nand U11433 (N_11433,N_5367,N_1434);
nor U11434 (N_11434,N_147,N_3713);
or U11435 (N_11435,N_4809,N_5029);
nand U11436 (N_11436,N_2940,N_5227);
and U11437 (N_11437,N_1573,N_2901);
nor U11438 (N_11438,N_5688,N_3820);
or U11439 (N_11439,N_815,N_2937);
nor U11440 (N_11440,N_3130,N_2049);
xnor U11441 (N_11441,N_68,N_3728);
nor U11442 (N_11442,N_646,N_1536);
xnor U11443 (N_11443,N_5442,N_5256);
nor U11444 (N_11444,N_1194,N_4317);
and U11445 (N_11445,N_958,N_2477);
xor U11446 (N_11446,N_1860,N_1639);
nor U11447 (N_11447,N_5370,N_4570);
xnor U11448 (N_11448,N_1711,N_1218);
or U11449 (N_11449,N_1748,N_2215);
xor U11450 (N_11450,N_5865,N_4763);
nor U11451 (N_11451,N_2595,N_2570);
nand U11452 (N_11452,N_1709,N_252);
xnor U11453 (N_11453,N_517,N_4914);
xnor U11454 (N_11454,N_2566,N_288);
nand U11455 (N_11455,N_2941,N_5109);
and U11456 (N_11456,N_2558,N_3778);
xnor U11457 (N_11457,N_1540,N_5016);
nand U11458 (N_11458,N_2120,N_3508);
or U11459 (N_11459,N_720,N_3279);
or U11460 (N_11460,N_4606,N_3824);
nand U11461 (N_11461,N_1635,N_3678);
xnor U11462 (N_11462,N_3394,N_3313);
xor U11463 (N_11463,N_3628,N_5010);
nand U11464 (N_11464,N_1553,N_2151);
nor U11465 (N_11465,N_4562,N_886);
and U11466 (N_11466,N_5467,N_358);
nor U11467 (N_11467,N_5253,N_2759);
and U11468 (N_11468,N_2514,N_4367);
nor U11469 (N_11469,N_2655,N_5142);
and U11470 (N_11470,N_2627,N_1565);
and U11471 (N_11471,N_3204,N_4053);
or U11472 (N_11472,N_5039,N_5024);
nor U11473 (N_11473,N_5798,N_4408);
xnor U11474 (N_11474,N_354,N_4809);
nand U11475 (N_11475,N_4023,N_223);
xnor U11476 (N_11476,N_5120,N_5279);
nor U11477 (N_11477,N_3340,N_5121);
xor U11478 (N_11478,N_6212,N_3686);
or U11479 (N_11479,N_5654,N_4780);
nand U11480 (N_11480,N_5601,N_2771);
nor U11481 (N_11481,N_777,N_1065);
or U11482 (N_11482,N_259,N_3757);
and U11483 (N_11483,N_3591,N_5144);
or U11484 (N_11484,N_5629,N_2144);
and U11485 (N_11485,N_5110,N_1563);
or U11486 (N_11486,N_4608,N_4848);
nor U11487 (N_11487,N_644,N_2712);
nand U11488 (N_11488,N_1894,N_1043);
nand U11489 (N_11489,N_4555,N_4437);
or U11490 (N_11490,N_2244,N_3774);
nand U11491 (N_11491,N_326,N_1584);
nand U11492 (N_11492,N_708,N_976);
xnor U11493 (N_11493,N_3064,N_5754);
or U11494 (N_11494,N_6202,N_2521);
xnor U11495 (N_11495,N_3063,N_5408);
or U11496 (N_11496,N_5421,N_4881);
nor U11497 (N_11497,N_1875,N_6018);
and U11498 (N_11498,N_1234,N_2244);
or U11499 (N_11499,N_1791,N_650);
nand U11500 (N_11500,N_2557,N_1814);
xnor U11501 (N_11501,N_3854,N_5141);
or U11502 (N_11502,N_1804,N_2177);
nand U11503 (N_11503,N_3107,N_5161);
xnor U11504 (N_11504,N_328,N_4862);
and U11505 (N_11505,N_1467,N_1120);
or U11506 (N_11506,N_1651,N_3440);
nor U11507 (N_11507,N_1985,N_3646);
nand U11508 (N_11508,N_5928,N_723);
or U11509 (N_11509,N_5578,N_1062);
or U11510 (N_11510,N_2203,N_3882);
nand U11511 (N_11511,N_578,N_4065);
or U11512 (N_11512,N_594,N_189);
nand U11513 (N_11513,N_2101,N_1988);
nor U11514 (N_11514,N_1188,N_2987);
and U11515 (N_11515,N_3278,N_5998);
and U11516 (N_11516,N_4688,N_5407);
or U11517 (N_11517,N_305,N_4414);
xnor U11518 (N_11518,N_653,N_4045);
or U11519 (N_11519,N_1278,N_63);
or U11520 (N_11520,N_2128,N_1219);
nor U11521 (N_11521,N_969,N_2217);
or U11522 (N_11522,N_1836,N_720);
and U11523 (N_11523,N_407,N_4304);
and U11524 (N_11524,N_1956,N_3068);
nor U11525 (N_11525,N_414,N_2238);
nor U11526 (N_11526,N_534,N_558);
nor U11527 (N_11527,N_1931,N_1011);
nor U11528 (N_11528,N_4447,N_5693);
nor U11529 (N_11529,N_2111,N_356);
or U11530 (N_11530,N_3208,N_5146);
nor U11531 (N_11531,N_2704,N_5087);
xor U11532 (N_11532,N_2152,N_3914);
nor U11533 (N_11533,N_930,N_2590);
or U11534 (N_11534,N_45,N_5259);
or U11535 (N_11535,N_2065,N_4269);
and U11536 (N_11536,N_4084,N_2807);
or U11537 (N_11537,N_228,N_216);
nor U11538 (N_11538,N_2353,N_5385);
xnor U11539 (N_11539,N_4479,N_5477);
or U11540 (N_11540,N_3464,N_3537);
xor U11541 (N_11541,N_871,N_5110);
xor U11542 (N_11542,N_2506,N_2612);
nand U11543 (N_11543,N_444,N_5670);
or U11544 (N_11544,N_4222,N_634);
nor U11545 (N_11545,N_4288,N_3894);
nor U11546 (N_11546,N_4960,N_5352);
nand U11547 (N_11547,N_761,N_5441);
and U11548 (N_11548,N_2731,N_1038);
or U11549 (N_11549,N_5753,N_1022);
and U11550 (N_11550,N_338,N_1563);
nor U11551 (N_11551,N_480,N_3412);
and U11552 (N_11552,N_6158,N_358);
nand U11553 (N_11553,N_2871,N_6034);
xor U11554 (N_11554,N_4850,N_5010);
and U11555 (N_11555,N_2228,N_3797);
nor U11556 (N_11556,N_3189,N_639);
nand U11557 (N_11557,N_647,N_3953);
or U11558 (N_11558,N_893,N_1477);
and U11559 (N_11559,N_4547,N_2935);
nand U11560 (N_11560,N_3790,N_3908);
xnor U11561 (N_11561,N_826,N_2771);
nor U11562 (N_11562,N_3954,N_4375);
or U11563 (N_11563,N_6157,N_582);
or U11564 (N_11564,N_3532,N_3371);
nand U11565 (N_11565,N_1977,N_6114);
nor U11566 (N_11566,N_3330,N_2099);
and U11567 (N_11567,N_508,N_920);
nor U11568 (N_11568,N_4778,N_3992);
and U11569 (N_11569,N_3043,N_4390);
or U11570 (N_11570,N_3543,N_2814);
xnor U11571 (N_11571,N_4834,N_5838);
nor U11572 (N_11572,N_3079,N_1005);
xor U11573 (N_11573,N_2128,N_5716);
xnor U11574 (N_11574,N_930,N_4279);
and U11575 (N_11575,N_2511,N_382);
or U11576 (N_11576,N_996,N_5827);
or U11577 (N_11577,N_3358,N_5173);
xor U11578 (N_11578,N_290,N_5469);
nand U11579 (N_11579,N_2871,N_3630);
and U11580 (N_11580,N_3897,N_214);
nor U11581 (N_11581,N_4826,N_1302);
or U11582 (N_11582,N_4804,N_5141);
nand U11583 (N_11583,N_5552,N_365);
nor U11584 (N_11584,N_5199,N_598);
nor U11585 (N_11585,N_3591,N_508);
nor U11586 (N_11586,N_3405,N_4664);
and U11587 (N_11587,N_2459,N_2849);
or U11588 (N_11588,N_3622,N_1203);
xor U11589 (N_11589,N_612,N_4939);
nand U11590 (N_11590,N_1541,N_1744);
nor U11591 (N_11591,N_4256,N_2309);
or U11592 (N_11592,N_4449,N_807);
and U11593 (N_11593,N_2640,N_4615);
nand U11594 (N_11594,N_1933,N_1921);
xnor U11595 (N_11595,N_4181,N_1103);
xor U11596 (N_11596,N_565,N_3483);
nand U11597 (N_11597,N_1960,N_1605);
nor U11598 (N_11598,N_1301,N_5498);
xor U11599 (N_11599,N_4805,N_1558);
or U11600 (N_11600,N_3940,N_4119);
and U11601 (N_11601,N_3724,N_2730);
or U11602 (N_11602,N_4617,N_4420);
xnor U11603 (N_11603,N_237,N_1855);
nand U11604 (N_11604,N_4192,N_3468);
nand U11605 (N_11605,N_5674,N_5384);
xnor U11606 (N_11606,N_2307,N_1786);
nor U11607 (N_11607,N_5030,N_4222);
and U11608 (N_11608,N_2146,N_1230);
xnor U11609 (N_11609,N_5266,N_4052);
or U11610 (N_11610,N_512,N_1898);
and U11611 (N_11611,N_2845,N_4366);
nand U11612 (N_11612,N_2112,N_2167);
or U11613 (N_11613,N_287,N_1152);
xnor U11614 (N_11614,N_2411,N_2146);
nand U11615 (N_11615,N_763,N_5356);
nand U11616 (N_11616,N_2989,N_4402);
or U11617 (N_11617,N_124,N_5567);
nand U11618 (N_11618,N_5115,N_2227);
nor U11619 (N_11619,N_4639,N_2150);
or U11620 (N_11620,N_4594,N_4326);
and U11621 (N_11621,N_5739,N_5708);
nand U11622 (N_11622,N_1752,N_6193);
nand U11623 (N_11623,N_103,N_4532);
nor U11624 (N_11624,N_726,N_581);
nand U11625 (N_11625,N_3748,N_2528);
nor U11626 (N_11626,N_5813,N_3120);
and U11627 (N_11627,N_3816,N_5368);
and U11628 (N_11628,N_2131,N_4253);
nor U11629 (N_11629,N_4265,N_5842);
nor U11630 (N_11630,N_441,N_2308);
nor U11631 (N_11631,N_872,N_1620);
xor U11632 (N_11632,N_1101,N_1561);
xnor U11633 (N_11633,N_4436,N_4145);
and U11634 (N_11634,N_4650,N_3247);
nand U11635 (N_11635,N_2645,N_1638);
and U11636 (N_11636,N_2358,N_5628);
and U11637 (N_11637,N_916,N_3718);
nor U11638 (N_11638,N_92,N_1503);
and U11639 (N_11639,N_2030,N_4102);
nor U11640 (N_11640,N_3290,N_1634);
and U11641 (N_11641,N_364,N_4646);
nor U11642 (N_11642,N_1528,N_4686);
xnor U11643 (N_11643,N_3993,N_5860);
nor U11644 (N_11644,N_1725,N_2863);
nand U11645 (N_11645,N_199,N_2982);
nor U11646 (N_11646,N_2813,N_5854);
nor U11647 (N_11647,N_2351,N_7);
or U11648 (N_11648,N_1579,N_5920);
xnor U11649 (N_11649,N_939,N_5103);
and U11650 (N_11650,N_5431,N_376);
nor U11651 (N_11651,N_4082,N_4642);
nand U11652 (N_11652,N_332,N_5489);
nor U11653 (N_11653,N_5336,N_2798);
nor U11654 (N_11654,N_3769,N_1005);
or U11655 (N_11655,N_879,N_3177);
and U11656 (N_11656,N_3864,N_6101);
xor U11657 (N_11657,N_1652,N_632);
or U11658 (N_11658,N_4878,N_78);
nand U11659 (N_11659,N_3883,N_2608);
or U11660 (N_11660,N_1471,N_3953);
nor U11661 (N_11661,N_4804,N_3505);
xor U11662 (N_11662,N_4328,N_5794);
xnor U11663 (N_11663,N_5387,N_4646);
xor U11664 (N_11664,N_1553,N_655);
xnor U11665 (N_11665,N_4287,N_4190);
nand U11666 (N_11666,N_5317,N_1832);
and U11667 (N_11667,N_516,N_3421);
nor U11668 (N_11668,N_1199,N_3480);
xnor U11669 (N_11669,N_3233,N_3736);
nand U11670 (N_11670,N_1778,N_6130);
nor U11671 (N_11671,N_4836,N_2475);
nand U11672 (N_11672,N_3373,N_5695);
or U11673 (N_11673,N_637,N_1287);
xnor U11674 (N_11674,N_2934,N_3847);
nand U11675 (N_11675,N_4627,N_2922);
or U11676 (N_11676,N_268,N_5048);
nor U11677 (N_11677,N_4622,N_680);
nand U11678 (N_11678,N_4626,N_2956);
and U11679 (N_11679,N_2159,N_916);
xor U11680 (N_11680,N_5866,N_1507);
xor U11681 (N_11681,N_1618,N_4598);
or U11682 (N_11682,N_3142,N_5178);
nor U11683 (N_11683,N_4723,N_2273);
xor U11684 (N_11684,N_5280,N_2827);
and U11685 (N_11685,N_5988,N_2047);
nand U11686 (N_11686,N_2466,N_5030);
xor U11687 (N_11687,N_1541,N_5968);
nand U11688 (N_11688,N_2941,N_2354);
nand U11689 (N_11689,N_6095,N_5815);
or U11690 (N_11690,N_2050,N_4691);
or U11691 (N_11691,N_4464,N_3734);
nor U11692 (N_11692,N_3730,N_4051);
and U11693 (N_11693,N_3904,N_2653);
or U11694 (N_11694,N_3710,N_1723);
xnor U11695 (N_11695,N_2101,N_2580);
xnor U11696 (N_11696,N_5245,N_371);
and U11697 (N_11697,N_3492,N_4839);
and U11698 (N_11698,N_136,N_1776);
xor U11699 (N_11699,N_485,N_4238);
and U11700 (N_11700,N_3192,N_4323);
and U11701 (N_11701,N_2426,N_4216);
or U11702 (N_11702,N_2576,N_542);
or U11703 (N_11703,N_321,N_5518);
xnor U11704 (N_11704,N_5268,N_3741);
xor U11705 (N_11705,N_6210,N_1482);
and U11706 (N_11706,N_4303,N_6042);
nor U11707 (N_11707,N_597,N_5680);
or U11708 (N_11708,N_5374,N_4511);
and U11709 (N_11709,N_5554,N_3893);
and U11710 (N_11710,N_4136,N_4060);
xnor U11711 (N_11711,N_2842,N_1803);
nor U11712 (N_11712,N_1882,N_4810);
nor U11713 (N_11713,N_2382,N_323);
nand U11714 (N_11714,N_1474,N_3148);
or U11715 (N_11715,N_4838,N_2254);
and U11716 (N_11716,N_2571,N_5067);
or U11717 (N_11717,N_1330,N_686);
nor U11718 (N_11718,N_6167,N_3687);
nor U11719 (N_11719,N_5869,N_3716);
or U11720 (N_11720,N_3959,N_5237);
or U11721 (N_11721,N_4148,N_3552);
or U11722 (N_11722,N_663,N_5565);
or U11723 (N_11723,N_4445,N_4997);
nor U11724 (N_11724,N_1137,N_62);
xor U11725 (N_11725,N_3401,N_181);
and U11726 (N_11726,N_555,N_5501);
or U11727 (N_11727,N_3972,N_4192);
or U11728 (N_11728,N_1800,N_1569);
xor U11729 (N_11729,N_3938,N_1725);
and U11730 (N_11730,N_4723,N_1883);
and U11731 (N_11731,N_823,N_5492);
nand U11732 (N_11732,N_129,N_597);
nor U11733 (N_11733,N_4364,N_1802);
nor U11734 (N_11734,N_142,N_4343);
and U11735 (N_11735,N_4773,N_3368);
xor U11736 (N_11736,N_2915,N_4128);
nand U11737 (N_11737,N_3652,N_3451);
nor U11738 (N_11738,N_2432,N_5010);
and U11739 (N_11739,N_2346,N_844);
xnor U11740 (N_11740,N_5196,N_4095);
xnor U11741 (N_11741,N_1263,N_839);
nor U11742 (N_11742,N_4355,N_5729);
or U11743 (N_11743,N_4265,N_2749);
and U11744 (N_11744,N_2168,N_2117);
nor U11745 (N_11745,N_5634,N_663);
or U11746 (N_11746,N_4447,N_3773);
xor U11747 (N_11747,N_1443,N_2255);
or U11748 (N_11748,N_4930,N_138);
xor U11749 (N_11749,N_1253,N_5468);
nand U11750 (N_11750,N_5666,N_3480);
nand U11751 (N_11751,N_2848,N_2094);
or U11752 (N_11752,N_5031,N_1972);
and U11753 (N_11753,N_5526,N_6160);
nor U11754 (N_11754,N_1772,N_2808);
xnor U11755 (N_11755,N_1414,N_1428);
nand U11756 (N_11756,N_6189,N_4512);
and U11757 (N_11757,N_1222,N_3616);
xor U11758 (N_11758,N_3715,N_2788);
xnor U11759 (N_11759,N_2133,N_765);
xnor U11760 (N_11760,N_2155,N_1667);
or U11761 (N_11761,N_4068,N_3044);
xnor U11762 (N_11762,N_1788,N_1636);
or U11763 (N_11763,N_5792,N_1921);
nor U11764 (N_11764,N_1646,N_2228);
nand U11765 (N_11765,N_4963,N_4025);
or U11766 (N_11766,N_4673,N_4273);
xor U11767 (N_11767,N_3999,N_931);
and U11768 (N_11768,N_5200,N_1428);
and U11769 (N_11769,N_2106,N_2108);
nand U11770 (N_11770,N_2168,N_3579);
and U11771 (N_11771,N_5633,N_2306);
and U11772 (N_11772,N_5526,N_1140);
and U11773 (N_11773,N_1549,N_1693);
nor U11774 (N_11774,N_2314,N_1479);
nor U11775 (N_11775,N_3759,N_1072);
nand U11776 (N_11776,N_1866,N_2845);
and U11777 (N_11777,N_2528,N_769);
or U11778 (N_11778,N_5961,N_5736);
and U11779 (N_11779,N_3444,N_2217);
nand U11780 (N_11780,N_4381,N_33);
xnor U11781 (N_11781,N_1696,N_662);
nand U11782 (N_11782,N_2605,N_5063);
nor U11783 (N_11783,N_2866,N_4837);
xnor U11784 (N_11784,N_2426,N_1126);
and U11785 (N_11785,N_5178,N_5413);
or U11786 (N_11786,N_4317,N_5420);
or U11787 (N_11787,N_3951,N_43);
xnor U11788 (N_11788,N_412,N_5070);
nand U11789 (N_11789,N_604,N_5705);
nand U11790 (N_11790,N_2561,N_6159);
and U11791 (N_11791,N_3102,N_507);
xnor U11792 (N_11792,N_5959,N_889);
xnor U11793 (N_11793,N_5680,N_1131);
nor U11794 (N_11794,N_4561,N_4266);
xor U11795 (N_11795,N_3901,N_4410);
xnor U11796 (N_11796,N_4727,N_3210);
nor U11797 (N_11797,N_3275,N_2980);
xor U11798 (N_11798,N_3625,N_98);
and U11799 (N_11799,N_6156,N_2778);
and U11800 (N_11800,N_3014,N_4804);
and U11801 (N_11801,N_6190,N_1458);
nand U11802 (N_11802,N_2945,N_205);
and U11803 (N_11803,N_4162,N_1484);
or U11804 (N_11804,N_1650,N_4099);
nor U11805 (N_11805,N_4841,N_5875);
and U11806 (N_11806,N_894,N_1136);
or U11807 (N_11807,N_2197,N_1377);
or U11808 (N_11808,N_5356,N_2343);
and U11809 (N_11809,N_1571,N_2571);
and U11810 (N_11810,N_80,N_5119);
or U11811 (N_11811,N_4624,N_3359);
nor U11812 (N_11812,N_727,N_5152);
nand U11813 (N_11813,N_3,N_3743);
nor U11814 (N_11814,N_1180,N_3456);
xnor U11815 (N_11815,N_2238,N_2183);
nor U11816 (N_11816,N_996,N_5884);
and U11817 (N_11817,N_5602,N_1098);
nand U11818 (N_11818,N_3885,N_1536);
and U11819 (N_11819,N_2824,N_798);
xnor U11820 (N_11820,N_1956,N_41);
xor U11821 (N_11821,N_1434,N_4863);
nor U11822 (N_11822,N_1223,N_1657);
nor U11823 (N_11823,N_2224,N_4639);
nand U11824 (N_11824,N_4019,N_47);
xnor U11825 (N_11825,N_196,N_5695);
nand U11826 (N_11826,N_1228,N_5572);
or U11827 (N_11827,N_1251,N_3236);
nand U11828 (N_11828,N_5122,N_1918);
nor U11829 (N_11829,N_2618,N_1512);
xnor U11830 (N_11830,N_4615,N_2891);
or U11831 (N_11831,N_4564,N_313);
and U11832 (N_11832,N_1776,N_750);
nand U11833 (N_11833,N_2648,N_2656);
nor U11834 (N_11834,N_5389,N_3513);
nand U11835 (N_11835,N_4071,N_3422);
xnor U11836 (N_11836,N_2696,N_223);
and U11837 (N_11837,N_900,N_5752);
nand U11838 (N_11838,N_833,N_5939);
and U11839 (N_11839,N_254,N_1104);
or U11840 (N_11840,N_2684,N_1289);
and U11841 (N_11841,N_5351,N_3168);
xnor U11842 (N_11842,N_4447,N_6061);
or U11843 (N_11843,N_3395,N_2561);
nor U11844 (N_11844,N_4724,N_771);
or U11845 (N_11845,N_3308,N_4053);
and U11846 (N_11846,N_2829,N_2669);
nand U11847 (N_11847,N_2580,N_5001);
xor U11848 (N_11848,N_3157,N_959);
xor U11849 (N_11849,N_2734,N_4790);
nor U11850 (N_11850,N_4318,N_2721);
or U11851 (N_11851,N_1840,N_2382);
and U11852 (N_11852,N_3785,N_3460);
nand U11853 (N_11853,N_4743,N_2949);
xor U11854 (N_11854,N_5336,N_3061);
nand U11855 (N_11855,N_3101,N_744);
nor U11856 (N_11856,N_4300,N_4045);
or U11857 (N_11857,N_5713,N_2879);
or U11858 (N_11858,N_420,N_3532);
xnor U11859 (N_11859,N_3507,N_969);
nor U11860 (N_11860,N_168,N_5470);
xnor U11861 (N_11861,N_4871,N_2426);
or U11862 (N_11862,N_5052,N_648);
and U11863 (N_11863,N_301,N_5986);
nand U11864 (N_11864,N_2737,N_3095);
or U11865 (N_11865,N_5429,N_2956);
nand U11866 (N_11866,N_2328,N_4408);
and U11867 (N_11867,N_1434,N_2950);
and U11868 (N_11868,N_4754,N_5552);
nand U11869 (N_11869,N_3300,N_4110);
xor U11870 (N_11870,N_5436,N_6234);
nand U11871 (N_11871,N_2151,N_4026);
and U11872 (N_11872,N_3489,N_5272);
xnor U11873 (N_11873,N_87,N_1734);
nand U11874 (N_11874,N_445,N_1205);
nand U11875 (N_11875,N_1722,N_3753);
nand U11876 (N_11876,N_2678,N_5507);
and U11877 (N_11877,N_6174,N_484);
and U11878 (N_11878,N_2619,N_3439);
or U11879 (N_11879,N_2826,N_4396);
nor U11880 (N_11880,N_2838,N_3834);
nand U11881 (N_11881,N_271,N_3198);
and U11882 (N_11882,N_734,N_4783);
xor U11883 (N_11883,N_48,N_3677);
and U11884 (N_11884,N_1698,N_2127);
nor U11885 (N_11885,N_1123,N_1645);
nor U11886 (N_11886,N_6180,N_1136);
xor U11887 (N_11887,N_3658,N_5300);
and U11888 (N_11888,N_5710,N_2417);
or U11889 (N_11889,N_2480,N_4797);
nand U11890 (N_11890,N_320,N_2891);
or U11891 (N_11891,N_3576,N_2097);
nor U11892 (N_11892,N_2923,N_2733);
and U11893 (N_11893,N_1114,N_5587);
nor U11894 (N_11894,N_1852,N_5431);
or U11895 (N_11895,N_3298,N_1703);
xor U11896 (N_11896,N_5552,N_1707);
xnor U11897 (N_11897,N_1184,N_4373);
nand U11898 (N_11898,N_5063,N_5908);
nor U11899 (N_11899,N_6177,N_4966);
xor U11900 (N_11900,N_1575,N_4472);
or U11901 (N_11901,N_4764,N_1090);
or U11902 (N_11902,N_3765,N_4373);
or U11903 (N_11903,N_2499,N_2859);
nand U11904 (N_11904,N_4847,N_4264);
xor U11905 (N_11905,N_6235,N_3584);
xnor U11906 (N_11906,N_3793,N_1458);
xnor U11907 (N_11907,N_587,N_2687);
and U11908 (N_11908,N_3308,N_3526);
and U11909 (N_11909,N_947,N_3800);
xnor U11910 (N_11910,N_3846,N_6173);
xnor U11911 (N_11911,N_1292,N_5373);
or U11912 (N_11912,N_4578,N_2201);
nand U11913 (N_11913,N_5707,N_490);
or U11914 (N_11914,N_5015,N_5751);
or U11915 (N_11915,N_4746,N_4192);
nor U11916 (N_11916,N_5160,N_448);
nor U11917 (N_11917,N_706,N_5314);
nor U11918 (N_11918,N_4601,N_817);
nor U11919 (N_11919,N_4981,N_3847);
and U11920 (N_11920,N_3870,N_5276);
and U11921 (N_11921,N_6154,N_1914);
xor U11922 (N_11922,N_1131,N_1503);
or U11923 (N_11923,N_5762,N_2100);
nor U11924 (N_11924,N_1509,N_51);
nor U11925 (N_11925,N_5537,N_3192);
or U11926 (N_11926,N_544,N_3644);
xor U11927 (N_11927,N_4659,N_2491);
or U11928 (N_11928,N_5458,N_915);
or U11929 (N_11929,N_4486,N_5047);
nand U11930 (N_11930,N_5384,N_2896);
or U11931 (N_11931,N_3834,N_2796);
or U11932 (N_11932,N_3375,N_3150);
nand U11933 (N_11933,N_5852,N_4530);
nand U11934 (N_11934,N_3743,N_6210);
or U11935 (N_11935,N_770,N_327);
or U11936 (N_11936,N_1039,N_5332);
nand U11937 (N_11937,N_3337,N_3515);
xnor U11938 (N_11938,N_3185,N_4085);
xor U11939 (N_11939,N_5900,N_2954);
nor U11940 (N_11940,N_64,N_1232);
nor U11941 (N_11941,N_6069,N_4282);
and U11942 (N_11942,N_3546,N_2721);
xor U11943 (N_11943,N_3791,N_4204);
and U11944 (N_11944,N_2725,N_3945);
nand U11945 (N_11945,N_3947,N_943);
or U11946 (N_11946,N_4260,N_1250);
or U11947 (N_11947,N_5626,N_318);
nand U11948 (N_11948,N_5213,N_3741);
or U11949 (N_11949,N_99,N_1098);
and U11950 (N_11950,N_5745,N_1325);
and U11951 (N_11951,N_1029,N_648);
and U11952 (N_11952,N_1358,N_5566);
nor U11953 (N_11953,N_5624,N_4908);
and U11954 (N_11954,N_3571,N_3898);
and U11955 (N_11955,N_5575,N_3817);
nand U11956 (N_11956,N_562,N_1546);
nand U11957 (N_11957,N_2275,N_5550);
nand U11958 (N_11958,N_1994,N_2388);
xor U11959 (N_11959,N_2600,N_1171);
and U11960 (N_11960,N_5667,N_855);
and U11961 (N_11961,N_4579,N_4294);
and U11962 (N_11962,N_316,N_5141);
nor U11963 (N_11963,N_2575,N_2633);
nand U11964 (N_11964,N_4460,N_6101);
or U11965 (N_11965,N_4318,N_3382);
nor U11966 (N_11966,N_6132,N_190);
nor U11967 (N_11967,N_6046,N_3383);
or U11968 (N_11968,N_4286,N_1087);
xor U11969 (N_11969,N_605,N_3245);
xor U11970 (N_11970,N_2673,N_5583);
nor U11971 (N_11971,N_4802,N_1473);
and U11972 (N_11972,N_4179,N_690);
and U11973 (N_11973,N_4330,N_1592);
and U11974 (N_11974,N_5035,N_1999);
or U11975 (N_11975,N_2997,N_5667);
nand U11976 (N_11976,N_555,N_4135);
xnor U11977 (N_11977,N_1533,N_3785);
nor U11978 (N_11978,N_5492,N_4332);
nand U11979 (N_11979,N_5912,N_6193);
nand U11980 (N_11980,N_2564,N_3940);
or U11981 (N_11981,N_2838,N_1590);
xnor U11982 (N_11982,N_1764,N_2421);
nand U11983 (N_11983,N_1401,N_3057);
xor U11984 (N_11984,N_3184,N_2518);
nor U11985 (N_11985,N_5220,N_3971);
nor U11986 (N_11986,N_703,N_1654);
nor U11987 (N_11987,N_4851,N_5485);
nor U11988 (N_11988,N_1564,N_5648);
xnor U11989 (N_11989,N_1313,N_1798);
xor U11990 (N_11990,N_1497,N_2570);
and U11991 (N_11991,N_3081,N_834);
nor U11992 (N_11992,N_1910,N_6161);
xnor U11993 (N_11993,N_316,N_1679);
or U11994 (N_11994,N_5106,N_143);
nand U11995 (N_11995,N_4118,N_1836);
and U11996 (N_11996,N_6101,N_544);
or U11997 (N_11997,N_332,N_3801);
and U11998 (N_11998,N_5362,N_5863);
and U11999 (N_11999,N_1863,N_274);
and U12000 (N_12000,N_1820,N_5942);
xnor U12001 (N_12001,N_3526,N_2043);
xor U12002 (N_12002,N_3899,N_5742);
or U12003 (N_12003,N_5622,N_4729);
xnor U12004 (N_12004,N_288,N_4863);
and U12005 (N_12005,N_106,N_5630);
or U12006 (N_12006,N_4841,N_3590);
nand U12007 (N_12007,N_5976,N_1038);
and U12008 (N_12008,N_4764,N_3255);
or U12009 (N_12009,N_1165,N_268);
nand U12010 (N_12010,N_1125,N_3238);
nand U12011 (N_12011,N_3867,N_3112);
and U12012 (N_12012,N_1345,N_244);
nand U12013 (N_12013,N_2387,N_2570);
and U12014 (N_12014,N_4414,N_3184);
and U12015 (N_12015,N_4086,N_1672);
or U12016 (N_12016,N_4062,N_4086);
or U12017 (N_12017,N_235,N_1075);
nand U12018 (N_12018,N_6,N_3930);
or U12019 (N_12019,N_1301,N_869);
or U12020 (N_12020,N_1256,N_3408);
and U12021 (N_12021,N_1270,N_3597);
and U12022 (N_12022,N_2052,N_5069);
nor U12023 (N_12023,N_1416,N_150);
and U12024 (N_12024,N_4041,N_2060);
nand U12025 (N_12025,N_2415,N_3765);
xor U12026 (N_12026,N_2848,N_4391);
nand U12027 (N_12027,N_4299,N_1524);
xnor U12028 (N_12028,N_5792,N_1068);
xnor U12029 (N_12029,N_1170,N_3140);
nand U12030 (N_12030,N_4999,N_2408);
nor U12031 (N_12031,N_4492,N_2595);
nor U12032 (N_12032,N_2710,N_2270);
or U12033 (N_12033,N_2839,N_5683);
or U12034 (N_12034,N_3712,N_2502);
nor U12035 (N_12035,N_5992,N_890);
xnor U12036 (N_12036,N_3480,N_1348);
xor U12037 (N_12037,N_5517,N_168);
nor U12038 (N_12038,N_2029,N_2160);
and U12039 (N_12039,N_5780,N_1924);
nor U12040 (N_12040,N_4913,N_4929);
xor U12041 (N_12041,N_5043,N_3177);
xor U12042 (N_12042,N_464,N_3730);
or U12043 (N_12043,N_710,N_3147);
nand U12044 (N_12044,N_1039,N_5337);
nand U12045 (N_12045,N_615,N_3607);
nand U12046 (N_12046,N_1531,N_2918);
nor U12047 (N_12047,N_3117,N_2628);
and U12048 (N_12048,N_5719,N_5428);
nand U12049 (N_12049,N_1159,N_1753);
xor U12050 (N_12050,N_3286,N_3228);
nor U12051 (N_12051,N_2247,N_2526);
xnor U12052 (N_12052,N_5487,N_3144);
and U12053 (N_12053,N_2626,N_1063);
xor U12054 (N_12054,N_1002,N_2055);
or U12055 (N_12055,N_1566,N_4788);
nor U12056 (N_12056,N_1940,N_4154);
nand U12057 (N_12057,N_5004,N_3453);
xnor U12058 (N_12058,N_2319,N_3217);
nand U12059 (N_12059,N_800,N_5214);
or U12060 (N_12060,N_1643,N_2660);
nand U12061 (N_12061,N_3736,N_63);
or U12062 (N_12062,N_3023,N_2630);
and U12063 (N_12063,N_5442,N_4392);
nor U12064 (N_12064,N_1276,N_2851);
nand U12065 (N_12065,N_2827,N_4373);
and U12066 (N_12066,N_5964,N_1712);
nor U12067 (N_12067,N_397,N_3956);
or U12068 (N_12068,N_606,N_4809);
or U12069 (N_12069,N_4871,N_4822);
and U12070 (N_12070,N_1295,N_5231);
nor U12071 (N_12071,N_1997,N_3560);
nor U12072 (N_12072,N_1398,N_4073);
xnor U12073 (N_12073,N_4102,N_757);
nor U12074 (N_12074,N_1769,N_5605);
nand U12075 (N_12075,N_3524,N_5114);
nor U12076 (N_12076,N_4809,N_2334);
or U12077 (N_12077,N_4606,N_1875);
nor U12078 (N_12078,N_2130,N_1416);
nor U12079 (N_12079,N_3939,N_2125);
or U12080 (N_12080,N_814,N_5237);
xor U12081 (N_12081,N_3035,N_5579);
xnor U12082 (N_12082,N_927,N_6094);
nand U12083 (N_12083,N_1282,N_1497);
nand U12084 (N_12084,N_834,N_5732);
or U12085 (N_12085,N_3444,N_2789);
nor U12086 (N_12086,N_2110,N_1004);
and U12087 (N_12087,N_1140,N_2917);
nand U12088 (N_12088,N_739,N_5496);
and U12089 (N_12089,N_3340,N_5858);
xor U12090 (N_12090,N_4472,N_4595);
and U12091 (N_12091,N_4446,N_301);
nor U12092 (N_12092,N_2575,N_3595);
or U12093 (N_12093,N_1991,N_3205);
xnor U12094 (N_12094,N_2347,N_1577);
or U12095 (N_12095,N_5213,N_4779);
and U12096 (N_12096,N_628,N_5477);
nor U12097 (N_12097,N_3468,N_2003);
nand U12098 (N_12098,N_391,N_3657);
or U12099 (N_12099,N_5723,N_1244);
or U12100 (N_12100,N_738,N_245);
nand U12101 (N_12101,N_1765,N_912);
nand U12102 (N_12102,N_5102,N_6137);
xnor U12103 (N_12103,N_29,N_427);
or U12104 (N_12104,N_4861,N_4002);
xor U12105 (N_12105,N_5983,N_973);
nand U12106 (N_12106,N_1501,N_5018);
nor U12107 (N_12107,N_1102,N_3355);
xor U12108 (N_12108,N_831,N_5440);
xnor U12109 (N_12109,N_112,N_1457);
xor U12110 (N_12110,N_6103,N_3851);
nor U12111 (N_12111,N_1135,N_2014);
or U12112 (N_12112,N_5691,N_919);
nor U12113 (N_12113,N_2835,N_5218);
xnor U12114 (N_12114,N_16,N_22);
xnor U12115 (N_12115,N_781,N_4928);
and U12116 (N_12116,N_1023,N_3263);
xnor U12117 (N_12117,N_3971,N_5327);
or U12118 (N_12118,N_1002,N_2895);
xor U12119 (N_12119,N_4750,N_3743);
xnor U12120 (N_12120,N_956,N_352);
or U12121 (N_12121,N_2598,N_679);
xor U12122 (N_12122,N_6217,N_1625);
or U12123 (N_12123,N_5265,N_4253);
xor U12124 (N_12124,N_5874,N_4560);
xnor U12125 (N_12125,N_4142,N_2556);
nand U12126 (N_12126,N_5706,N_6197);
or U12127 (N_12127,N_5454,N_3447);
xor U12128 (N_12128,N_3339,N_4332);
and U12129 (N_12129,N_5468,N_4995);
or U12130 (N_12130,N_493,N_7);
nand U12131 (N_12131,N_3382,N_5134);
xnor U12132 (N_12132,N_2954,N_182);
xor U12133 (N_12133,N_3389,N_4693);
and U12134 (N_12134,N_4611,N_1687);
or U12135 (N_12135,N_4671,N_2378);
or U12136 (N_12136,N_1710,N_3855);
xor U12137 (N_12137,N_4135,N_3566);
nand U12138 (N_12138,N_2301,N_2686);
xnor U12139 (N_12139,N_5352,N_1514);
and U12140 (N_12140,N_1376,N_4370);
or U12141 (N_12141,N_4088,N_795);
and U12142 (N_12142,N_5633,N_2449);
xnor U12143 (N_12143,N_944,N_376);
xnor U12144 (N_12144,N_5693,N_1064);
nand U12145 (N_12145,N_3450,N_6112);
or U12146 (N_12146,N_4988,N_5378);
and U12147 (N_12147,N_2299,N_1949);
xnor U12148 (N_12148,N_2867,N_3577);
or U12149 (N_12149,N_4531,N_1791);
and U12150 (N_12150,N_5270,N_4347);
xor U12151 (N_12151,N_2723,N_4590);
nor U12152 (N_12152,N_3611,N_955);
nor U12153 (N_12153,N_501,N_2788);
nor U12154 (N_12154,N_3059,N_4477);
xnor U12155 (N_12155,N_3569,N_1937);
and U12156 (N_12156,N_5759,N_1473);
nor U12157 (N_12157,N_4360,N_2988);
xor U12158 (N_12158,N_4089,N_4339);
nand U12159 (N_12159,N_1415,N_276);
and U12160 (N_12160,N_4238,N_1623);
and U12161 (N_12161,N_4535,N_2353);
nor U12162 (N_12162,N_3104,N_5048);
xnor U12163 (N_12163,N_4625,N_2643);
nand U12164 (N_12164,N_5132,N_4811);
or U12165 (N_12165,N_4388,N_2134);
and U12166 (N_12166,N_4078,N_3630);
and U12167 (N_12167,N_2880,N_5722);
xor U12168 (N_12168,N_3787,N_6026);
nor U12169 (N_12169,N_1570,N_2430);
nor U12170 (N_12170,N_3799,N_1113);
nand U12171 (N_12171,N_4679,N_5922);
xor U12172 (N_12172,N_5892,N_3580);
xnor U12173 (N_12173,N_1504,N_1559);
or U12174 (N_12174,N_10,N_5774);
or U12175 (N_12175,N_2105,N_2316);
or U12176 (N_12176,N_5874,N_749);
or U12177 (N_12177,N_3836,N_2411);
or U12178 (N_12178,N_1592,N_3555);
and U12179 (N_12179,N_2928,N_2842);
xor U12180 (N_12180,N_1298,N_1240);
xnor U12181 (N_12181,N_2108,N_5803);
nor U12182 (N_12182,N_4085,N_1414);
or U12183 (N_12183,N_324,N_1917);
or U12184 (N_12184,N_743,N_3603);
xnor U12185 (N_12185,N_1041,N_3225);
nor U12186 (N_12186,N_2224,N_1705);
or U12187 (N_12187,N_5378,N_1564);
nand U12188 (N_12188,N_4709,N_4771);
nand U12189 (N_12189,N_6092,N_2962);
nor U12190 (N_12190,N_5921,N_1636);
nand U12191 (N_12191,N_4233,N_1159);
nand U12192 (N_12192,N_2874,N_6113);
or U12193 (N_12193,N_6210,N_669);
or U12194 (N_12194,N_2835,N_2393);
and U12195 (N_12195,N_1750,N_2332);
nor U12196 (N_12196,N_664,N_5614);
nor U12197 (N_12197,N_4290,N_3071);
xor U12198 (N_12198,N_5430,N_1393);
or U12199 (N_12199,N_3430,N_1816);
or U12200 (N_12200,N_5114,N_1253);
or U12201 (N_12201,N_3357,N_2019);
nor U12202 (N_12202,N_554,N_457);
nor U12203 (N_12203,N_2812,N_1890);
nand U12204 (N_12204,N_5304,N_3979);
xnor U12205 (N_12205,N_5629,N_6204);
and U12206 (N_12206,N_5164,N_5338);
xnor U12207 (N_12207,N_5930,N_5416);
or U12208 (N_12208,N_4184,N_4883);
or U12209 (N_12209,N_361,N_220);
nand U12210 (N_12210,N_4612,N_1808);
nand U12211 (N_12211,N_5947,N_2598);
nand U12212 (N_12212,N_1204,N_2047);
nor U12213 (N_12213,N_1109,N_583);
nand U12214 (N_12214,N_1793,N_911);
or U12215 (N_12215,N_2532,N_428);
or U12216 (N_12216,N_2565,N_1620);
nand U12217 (N_12217,N_2337,N_4389);
xnor U12218 (N_12218,N_4093,N_2659);
nand U12219 (N_12219,N_4884,N_2389);
and U12220 (N_12220,N_2190,N_3367);
and U12221 (N_12221,N_4186,N_4815);
or U12222 (N_12222,N_2910,N_4490);
and U12223 (N_12223,N_1252,N_4641);
or U12224 (N_12224,N_3264,N_2023);
and U12225 (N_12225,N_3205,N_1);
and U12226 (N_12226,N_986,N_1705);
xor U12227 (N_12227,N_3834,N_3213);
nand U12228 (N_12228,N_5427,N_2282);
and U12229 (N_12229,N_4644,N_1943);
xnor U12230 (N_12230,N_2277,N_1303);
nand U12231 (N_12231,N_2749,N_5933);
or U12232 (N_12232,N_1235,N_3202);
nand U12233 (N_12233,N_5488,N_864);
or U12234 (N_12234,N_5254,N_63);
nand U12235 (N_12235,N_1516,N_2743);
xor U12236 (N_12236,N_3658,N_4219);
nand U12237 (N_12237,N_591,N_3168);
nor U12238 (N_12238,N_695,N_4604);
or U12239 (N_12239,N_2428,N_153);
nor U12240 (N_12240,N_511,N_1826);
or U12241 (N_12241,N_1849,N_4879);
nor U12242 (N_12242,N_6078,N_1791);
and U12243 (N_12243,N_3920,N_435);
and U12244 (N_12244,N_4995,N_2059);
xnor U12245 (N_12245,N_1317,N_399);
nor U12246 (N_12246,N_1552,N_1228);
or U12247 (N_12247,N_4684,N_2452);
nand U12248 (N_12248,N_3986,N_4340);
nand U12249 (N_12249,N_577,N_2373);
nor U12250 (N_12250,N_5570,N_1006);
xor U12251 (N_12251,N_5926,N_1341);
nand U12252 (N_12252,N_5837,N_5027);
nor U12253 (N_12253,N_4426,N_3387);
xor U12254 (N_12254,N_2158,N_4429);
nor U12255 (N_12255,N_3039,N_78);
and U12256 (N_12256,N_5404,N_674);
nor U12257 (N_12257,N_4970,N_5973);
and U12258 (N_12258,N_4886,N_2195);
nand U12259 (N_12259,N_3363,N_2598);
nand U12260 (N_12260,N_6247,N_4042);
xor U12261 (N_12261,N_1724,N_4957);
and U12262 (N_12262,N_1036,N_1835);
xor U12263 (N_12263,N_1812,N_4599);
xnor U12264 (N_12264,N_460,N_6139);
nor U12265 (N_12265,N_5599,N_5393);
or U12266 (N_12266,N_4335,N_302);
nor U12267 (N_12267,N_6017,N_5766);
nand U12268 (N_12268,N_1689,N_4826);
nor U12269 (N_12269,N_4042,N_1723);
xor U12270 (N_12270,N_3018,N_1343);
nand U12271 (N_12271,N_2337,N_318);
and U12272 (N_12272,N_4040,N_3779);
nor U12273 (N_12273,N_1284,N_5520);
xnor U12274 (N_12274,N_5839,N_658);
or U12275 (N_12275,N_3489,N_1914);
or U12276 (N_12276,N_3838,N_3997);
nand U12277 (N_12277,N_3775,N_3953);
xor U12278 (N_12278,N_5329,N_1972);
nand U12279 (N_12279,N_4748,N_2381);
nor U12280 (N_12280,N_5906,N_1964);
xor U12281 (N_12281,N_2907,N_1293);
nand U12282 (N_12282,N_4253,N_3988);
nand U12283 (N_12283,N_1190,N_2192);
nor U12284 (N_12284,N_1073,N_1146);
and U12285 (N_12285,N_130,N_526);
or U12286 (N_12286,N_5703,N_3833);
nor U12287 (N_12287,N_525,N_5595);
and U12288 (N_12288,N_5142,N_1114);
xor U12289 (N_12289,N_334,N_4725);
xnor U12290 (N_12290,N_4492,N_3281);
and U12291 (N_12291,N_5075,N_1158);
xor U12292 (N_12292,N_1737,N_138);
nand U12293 (N_12293,N_4816,N_5776);
xor U12294 (N_12294,N_5993,N_6088);
xor U12295 (N_12295,N_3939,N_291);
or U12296 (N_12296,N_167,N_1613);
or U12297 (N_12297,N_1562,N_3576);
nand U12298 (N_12298,N_3593,N_3300);
xnor U12299 (N_12299,N_5862,N_3023);
nand U12300 (N_12300,N_1491,N_1140);
nand U12301 (N_12301,N_1532,N_634);
nor U12302 (N_12302,N_3364,N_1992);
xor U12303 (N_12303,N_3870,N_2187);
nand U12304 (N_12304,N_4285,N_1185);
nor U12305 (N_12305,N_2782,N_17);
and U12306 (N_12306,N_5537,N_546);
and U12307 (N_12307,N_3816,N_4996);
nand U12308 (N_12308,N_5606,N_2537);
nor U12309 (N_12309,N_3333,N_2696);
nand U12310 (N_12310,N_2955,N_782);
nor U12311 (N_12311,N_2789,N_1757);
and U12312 (N_12312,N_5513,N_2889);
nor U12313 (N_12313,N_1446,N_2759);
nor U12314 (N_12314,N_1175,N_1830);
or U12315 (N_12315,N_776,N_4769);
xnor U12316 (N_12316,N_3363,N_6060);
xor U12317 (N_12317,N_1466,N_973);
or U12318 (N_12318,N_5145,N_3435);
or U12319 (N_12319,N_1827,N_2414);
xnor U12320 (N_12320,N_3938,N_857);
xor U12321 (N_12321,N_154,N_886);
xnor U12322 (N_12322,N_4295,N_1773);
xor U12323 (N_12323,N_1254,N_4187);
or U12324 (N_12324,N_2076,N_4078);
nor U12325 (N_12325,N_4821,N_4053);
nand U12326 (N_12326,N_4386,N_5657);
nor U12327 (N_12327,N_1066,N_3061);
xnor U12328 (N_12328,N_6075,N_2363);
and U12329 (N_12329,N_2010,N_940);
nor U12330 (N_12330,N_5568,N_1372);
or U12331 (N_12331,N_2228,N_4611);
xor U12332 (N_12332,N_4279,N_1065);
and U12333 (N_12333,N_1431,N_5972);
nand U12334 (N_12334,N_6045,N_4914);
xnor U12335 (N_12335,N_2563,N_3820);
nand U12336 (N_12336,N_4040,N_2303);
and U12337 (N_12337,N_3181,N_1946);
or U12338 (N_12338,N_6002,N_4842);
nand U12339 (N_12339,N_4669,N_5064);
or U12340 (N_12340,N_746,N_370);
xor U12341 (N_12341,N_2115,N_932);
or U12342 (N_12342,N_3895,N_2467);
nor U12343 (N_12343,N_1662,N_3598);
or U12344 (N_12344,N_5888,N_5045);
nand U12345 (N_12345,N_1856,N_3313);
nand U12346 (N_12346,N_229,N_3360);
or U12347 (N_12347,N_1758,N_1410);
and U12348 (N_12348,N_5052,N_6020);
xnor U12349 (N_12349,N_3924,N_1607);
and U12350 (N_12350,N_5859,N_5494);
or U12351 (N_12351,N_925,N_5725);
and U12352 (N_12352,N_5520,N_678);
or U12353 (N_12353,N_4414,N_4809);
or U12354 (N_12354,N_5431,N_2362);
nand U12355 (N_12355,N_4642,N_2237);
xor U12356 (N_12356,N_5112,N_1819);
nand U12357 (N_12357,N_1668,N_6005);
or U12358 (N_12358,N_919,N_4770);
nor U12359 (N_12359,N_4177,N_1745);
xnor U12360 (N_12360,N_5503,N_969);
or U12361 (N_12361,N_5644,N_3632);
xor U12362 (N_12362,N_5994,N_4632);
xnor U12363 (N_12363,N_1467,N_4348);
or U12364 (N_12364,N_5646,N_1829);
nand U12365 (N_12365,N_4213,N_4037);
nor U12366 (N_12366,N_3576,N_952);
or U12367 (N_12367,N_1548,N_4563);
nand U12368 (N_12368,N_5078,N_1476);
and U12369 (N_12369,N_5405,N_2729);
or U12370 (N_12370,N_2086,N_4433);
or U12371 (N_12371,N_5410,N_626);
nand U12372 (N_12372,N_1123,N_17);
and U12373 (N_12373,N_4933,N_307);
nor U12374 (N_12374,N_5856,N_4335);
nand U12375 (N_12375,N_547,N_4453);
nand U12376 (N_12376,N_397,N_2192);
xnor U12377 (N_12377,N_436,N_2684);
nand U12378 (N_12378,N_2970,N_2538);
nand U12379 (N_12379,N_4191,N_689);
or U12380 (N_12380,N_5380,N_4191);
and U12381 (N_12381,N_3607,N_791);
nand U12382 (N_12382,N_3926,N_3323);
nand U12383 (N_12383,N_3848,N_470);
xnor U12384 (N_12384,N_4218,N_5928);
or U12385 (N_12385,N_1719,N_706);
nor U12386 (N_12386,N_2541,N_1185);
nor U12387 (N_12387,N_4820,N_5626);
xor U12388 (N_12388,N_2150,N_225);
nor U12389 (N_12389,N_4607,N_2651);
xnor U12390 (N_12390,N_4702,N_2839);
nor U12391 (N_12391,N_5865,N_5206);
nor U12392 (N_12392,N_26,N_3003);
or U12393 (N_12393,N_5811,N_1568);
nor U12394 (N_12394,N_5143,N_3571);
or U12395 (N_12395,N_3614,N_5847);
xnor U12396 (N_12396,N_1346,N_4070);
and U12397 (N_12397,N_333,N_2596);
xnor U12398 (N_12398,N_5298,N_1949);
xnor U12399 (N_12399,N_5739,N_5491);
nand U12400 (N_12400,N_2017,N_467);
and U12401 (N_12401,N_2053,N_696);
nand U12402 (N_12402,N_4195,N_89);
nand U12403 (N_12403,N_4212,N_3125);
nor U12404 (N_12404,N_2738,N_1505);
or U12405 (N_12405,N_3764,N_4218);
nand U12406 (N_12406,N_3105,N_5023);
or U12407 (N_12407,N_6157,N_878);
or U12408 (N_12408,N_6145,N_1683);
xor U12409 (N_12409,N_484,N_1320);
nor U12410 (N_12410,N_6180,N_5429);
nand U12411 (N_12411,N_1169,N_2993);
nand U12412 (N_12412,N_6076,N_1349);
or U12413 (N_12413,N_2504,N_5767);
and U12414 (N_12414,N_3458,N_1120);
and U12415 (N_12415,N_441,N_5665);
or U12416 (N_12416,N_3094,N_4004);
and U12417 (N_12417,N_2449,N_1340);
nor U12418 (N_12418,N_4212,N_4044);
or U12419 (N_12419,N_1721,N_774);
and U12420 (N_12420,N_1521,N_1431);
nand U12421 (N_12421,N_9,N_1577);
or U12422 (N_12422,N_1469,N_1285);
or U12423 (N_12423,N_2257,N_419);
or U12424 (N_12424,N_44,N_2263);
and U12425 (N_12425,N_656,N_6247);
nor U12426 (N_12426,N_5448,N_3191);
xnor U12427 (N_12427,N_3041,N_4824);
and U12428 (N_12428,N_2642,N_1984);
and U12429 (N_12429,N_496,N_4930);
or U12430 (N_12430,N_5547,N_2239);
or U12431 (N_12431,N_3935,N_4956);
xor U12432 (N_12432,N_5915,N_6092);
nor U12433 (N_12433,N_362,N_3994);
nand U12434 (N_12434,N_894,N_4866);
and U12435 (N_12435,N_136,N_2952);
and U12436 (N_12436,N_1575,N_382);
nand U12437 (N_12437,N_1482,N_3962);
and U12438 (N_12438,N_2698,N_2237);
nand U12439 (N_12439,N_2678,N_1020);
xnor U12440 (N_12440,N_501,N_4231);
xnor U12441 (N_12441,N_1441,N_3701);
or U12442 (N_12442,N_4276,N_3551);
and U12443 (N_12443,N_4062,N_6091);
nand U12444 (N_12444,N_2430,N_1032);
and U12445 (N_12445,N_271,N_328);
or U12446 (N_12446,N_3600,N_4943);
nand U12447 (N_12447,N_1444,N_4056);
xor U12448 (N_12448,N_3070,N_1940);
nand U12449 (N_12449,N_1073,N_4099);
nor U12450 (N_12450,N_3040,N_5047);
and U12451 (N_12451,N_1932,N_3608);
xor U12452 (N_12452,N_3186,N_1522);
xor U12453 (N_12453,N_4971,N_4833);
and U12454 (N_12454,N_1300,N_2849);
xnor U12455 (N_12455,N_2617,N_4513);
nand U12456 (N_12456,N_5003,N_4965);
or U12457 (N_12457,N_6004,N_724);
nand U12458 (N_12458,N_1838,N_3122);
or U12459 (N_12459,N_5614,N_5311);
nor U12460 (N_12460,N_372,N_6045);
or U12461 (N_12461,N_5056,N_1597);
and U12462 (N_12462,N_5151,N_1102);
and U12463 (N_12463,N_3999,N_2966);
or U12464 (N_12464,N_713,N_2260);
nand U12465 (N_12465,N_5487,N_4387);
xnor U12466 (N_12466,N_5610,N_1149);
nor U12467 (N_12467,N_4886,N_592);
nand U12468 (N_12468,N_80,N_4564);
nand U12469 (N_12469,N_5331,N_5193);
and U12470 (N_12470,N_5634,N_3486);
or U12471 (N_12471,N_2095,N_3178);
or U12472 (N_12472,N_646,N_3921);
xor U12473 (N_12473,N_3118,N_4963);
nand U12474 (N_12474,N_5332,N_831);
xor U12475 (N_12475,N_5184,N_2128);
xnor U12476 (N_12476,N_5416,N_5150);
xnor U12477 (N_12477,N_3445,N_5593);
xor U12478 (N_12478,N_3527,N_5938);
and U12479 (N_12479,N_6175,N_3122);
nor U12480 (N_12480,N_3415,N_3126);
xnor U12481 (N_12481,N_5767,N_3081);
xor U12482 (N_12482,N_3852,N_4737);
nand U12483 (N_12483,N_5586,N_3856);
xor U12484 (N_12484,N_5864,N_2384);
xor U12485 (N_12485,N_1415,N_827);
and U12486 (N_12486,N_4469,N_334);
or U12487 (N_12487,N_4918,N_1926);
nand U12488 (N_12488,N_4670,N_3489);
xor U12489 (N_12489,N_1222,N_10);
nor U12490 (N_12490,N_929,N_71);
nand U12491 (N_12491,N_1501,N_4054);
nor U12492 (N_12492,N_5694,N_2690);
nand U12493 (N_12493,N_1482,N_559);
nor U12494 (N_12494,N_5518,N_2663);
and U12495 (N_12495,N_876,N_2997);
nand U12496 (N_12496,N_5693,N_6142);
and U12497 (N_12497,N_2799,N_6119);
nor U12498 (N_12498,N_4884,N_2013);
or U12499 (N_12499,N_658,N_4988);
xnor U12500 (N_12500,N_10510,N_6695);
xnor U12501 (N_12501,N_9052,N_6626);
or U12502 (N_12502,N_10004,N_9939);
xnor U12503 (N_12503,N_7923,N_8384);
nor U12504 (N_12504,N_12149,N_11983);
nand U12505 (N_12505,N_7408,N_7730);
and U12506 (N_12506,N_11605,N_12495);
nor U12507 (N_12507,N_8900,N_8662);
or U12508 (N_12508,N_8204,N_6919);
or U12509 (N_12509,N_8884,N_9018);
or U12510 (N_12510,N_10549,N_7057);
nand U12511 (N_12511,N_6740,N_11132);
nand U12512 (N_12512,N_7982,N_8284);
and U12513 (N_12513,N_6388,N_9949);
nand U12514 (N_12514,N_7744,N_9361);
and U12515 (N_12515,N_11315,N_9155);
or U12516 (N_12516,N_8944,N_8534);
or U12517 (N_12517,N_12062,N_8345);
and U12518 (N_12518,N_12081,N_10643);
and U12519 (N_12519,N_10214,N_7221);
xor U12520 (N_12520,N_7513,N_9754);
and U12521 (N_12521,N_9844,N_7196);
and U12522 (N_12522,N_11706,N_7604);
or U12523 (N_12523,N_6384,N_9071);
and U12524 (N_12524,N_6535,N_8748);
nor U12525 (N_12525,N_8160,N_6266);
nor U12526 (N_12526,N_6389,N_8268);
or U12527 (N_12527,N_6811,N_11876);
nor U12528 (N_12528,N_10270,N_6513);
xor U12529 (N_12529,N_11211,N_12443);
and U12530 (N_12530,N_7470,N_12209);
nor U12531 (N_12531,N_10915,N_9792);
xnor U12532 (N_12532,N_10357,N_7825);
and U12533 (N_12533,N_10425,N_9930);
xor U12534 (N_12534,N_6428,N_8706);
nor U12535 (N_12535,N_10031,N_11367);
or U12536 (N_12536,N_11375,N_11860);
xnor U12537 (N_12537,N_11448,N_6478);
nand U12538 (N_12538,N_8048,N_8556);
or U12539 (N_12539,N_12009,N_8723);
and U12540 (N_12540,N_7211,N_10500);
nand U12541 (N_12541,N_11297,N_9408);
or U12542 (N_12542,N_8100,N_10252);
nor U12543 (N_12543,N_12195,N_9055);
and U12544 (N_12544,N_12322,N_11589);
nor U12545 (N_12545,N_7950,N_9958);
nor U12546 (N_12546,N_11334,N_12039);
nand U12547 (N_12547,N_11823,N_8796);
xor U12548 (N_12548,N_7208,N_6824);
or U12549 (N_12549,N_6550,N_8734);
or U12550 (N_12550,N_7350,N_9468);
xnor U12551 (N_12551,N_9800,N_11759);
nand U12552 (N_12552,N_11900,N_10275);
nor U12553 (N_12553,N_6840,N_6312);
nand U12554 (N_12554,N_12437,N_6296);
xnor U12555 (N_12555,N_11598,N_11463);
xnor U12556 (N_12556,N_8569,N_11433);
nor U12557 (N_12557,N_7724,N_11370);
nand U12558 (N_12558,N_11677,N_10021);
xor U12559 (N_12559,N_6771,N_10746);
nand U12560 (N_12560,N_10015,N_6650);
nand U12561 (N_12561,N_11692,N_7125);
or U12562 (N_12562,N_10736,N_11953);
nor U12563 (N_12563,N_8770,N_7410);
nand U12564 (N_12564,N_10088,N_9385);
and U12565 (N_12565,N_11870,N_12091);
and U12566 (N_12566,N_7426,N_10895);
xor U12567 (N_12567,N_8372,N_10162);
or U12568 (N_12568,N_10817,N_10314);
nor U12569 (N_12569,N_8450,N_7404);
and U12570 (N_12570,N_8609,N_12256);
or U12571 (N_12571,N_8524,N_9223);
nor U12572 (N_12572,N_6619,N_7231);
nand U12573 (N_12573,N_11176,N_11063);
nor U12574 (N_12574,N_11635,N_12139);
nor U12575 (N_12575,N_9216,N_10366);
and U12576 (N_12576,N_8459,N_11928);
or U12577 (N_12577,N_9301,N_11806);
and U12578 (N_12578,N_9138,N_8039);
and U12579 (N_12579,N_11630,N_8879);
xor U12580 (N_12580,N_11530,N_9245);
xor U12581 (N_12581,N_10731,N_7786);
or U12582 (N_12582,N_11972,N_10960);
or U12583 (N_12583,N_10637,N_7465);
nor U12584 (N_12584,N_11970,N_10049);
and U12585 (N_12585,N_10507,N_7083);
or U12586 (N_12586,N_11144,N_12033);
xnor U12587 (N_12587,N_7941,N_10452);
nor U12588 (N_12588,N_9684,N_9236);
and U12589 (N_12589,N_9940,N_6863);
xor U12590 (N_12590,N_11331,N_11414);
nand U12591 (N_12591,N_10904,N_9523);
and U12592 (N_12592,N_10139,N_10145);
or U12593 (N_12593,N_8830,N_7387);
xor U12594 (N_12594,N_8259,N_10970);
nor U12595 (N_12595,N_10212,N_9397);
or U12596 (N_12596,N_8820,N_7713);
nor U12597 (N_12597,N_7314,N_6806);
and U12598 (N_12598,N_8171,N_8907);
and U12599 (N_12599,N_11381,N_11724);
or U12600 (N_12600,N_12023,N_10665);
nor U12601 (N_12601,N_6892,N_11417);
nand U12602 (N_12602,N_11950,N_8727);
and U12603 (N_12603,N_6782,N_8547);
nand U12604 (N_12604,N_11425,N_6589);
nor U12605 (N_12605,N_8050,N_7640);
and U12606 (N_12606,N_8823,N_6802);
nand U12607 (N_12607,N_7137,N_11701);
xor U12608 (N_12608,N_6670,N_12113);
or U12609 (N_12609,N_6257,N_8894);
nand U12610 (N_12610,N_11384,N_7702);
or U12611 (N_12611,N_6313,N_6653);
nand U12612 (N_12612,N_10773,N_7178);
and U12613 (N_12613,N_10435,N_12153);
or U12614 (N_12614,N_10753,N_9588);
and U12615 (N_12615,N_10278,N_11411);
or U12616 (N_12616,N_11632,N_9547);
xor U12617 (N_12617,N_10563,N_9276);
nand U12618 (N_12618,N_8242,N_6505);
nand U12619 (N_12619,N_12066,N_6768);
or U12620 (N_12620,N_8883,N_12211);
xor U12621 (N_12621,N_8669,N_8014);
xnor U12622 (N_12622,N_11321,N_8403);
or U12623 (N_12623,N_6449,N_8431);
nand U12624 (N_12624,N_9039,N_11969);
and U12625 (N_12625,N_7583,N_12354);
xnor U12626 (N_12626,N_9540,N_7358);
or U12627 (N_12627,N_10785,N_11225);
or U12628 (N_12628,N_11406,N_11140);
nand U12629 (N_12629,N_6672,N_6747);
or U12630 (N_12630,N_6661,N_6657);
or U12631 (N_12631,N_10838,N_8525);
nand U12632 (N_12632,N_10147,N_9582);
nand U12633 (N_12633,N_10429,N_6510);
nand U12634 (N_12634,N_12212,N_7187);
nand U12635 (N_12635,N_8809,N_6576);
nand U12636 (N_12636,N_9185,N_12353);
xor U12637 (N_12637,N_8447,N_7468);
and U12638 (N_12638,N_10983,N_8870);
or U12639 (N_12639,N_9491,N_11846);
nor U12640 (N_12640,N_7830,N_8363);
and U12641 (N_12641,N_8189,N_9115);
xor U12642 (N_12642,N_8742,N_10709);
nand U12643 (N_12643,N_6334,N_9835);
or U12644 (N_12644,N_8010,N_8341);
or U12645 (N_12645,N_8665,N_10697);
nand U12646 (N_12646,N_8410,N_10047);
xor U12647 (N_12647,N_10690,N_11429);
or U12648 (N_12648,N_9304,N_12390);
or U12649 (N_12649,N_7489,N_8948);
or U12650 (N_12650,N_10824,N_11765);
or U12651 (N_12651,N_8757,N_6324);
nor U12652 (N_12652,N_9336,N_9541);
or U12653 (N_12653,N_9924,N_11743);
or U12654 (N_12654,N_8562,N_7797);
and U12655 (N_12655,N_10091,N_9649);
and U12656 (N_12656,N_8200,N_11609);
and U12657 (N_12657,N_7336,N_9334);
nand U12658 (N_12658,N_11456,N_11282);
xor U12659 (N_12659,N_8094,N_8674);
and U12660 (N_12660,N_9340,N_12108);
nand U12661 (N_12661,N_10149,N_7701);
nor U12662 (N_12662,N_7972,N_9507);
nor U12663 (N_12663,N_7021,N_11145);
or U12664 (N_12664,N_8080,N_9598);
nor U12665 (N_12665,N_8302,N_6748);
and U12666 (N_12666,N_7684,N_8730);
nor U12667 (N_12667,N_9787,N_10787);
nand U12668 (N_12668,N_10856,N_12125);
nor U12669 (N_12669,N_6659,N_7613);
xnor U12670 (N_12670,N_7811,N_10104);
or U12671 (N_12671,N_9224,N_10554);
xnor U12672 (N_12672,N_10737,N_10401);
xor U12673 (N_12673,N_11528,N_6775);
or U12674 (N_12674,N_7341,N_10857);
and U12675 (N_12675,N_10791,N_12118);
nor U12676 (N_12676,N_9697,N_9022);
or U12677 (N_12677,N_8527,N_11614);
or U12678 (N_12678,N_11544,N_7594);
nand U12679 (N_12679,N_7624,N_7148);
or U12680 (N_12680,N_7429,N_8538);
and U12681 (N_12681,N_6814,N_7672);
xnor U12682 (N_12682,N_10625,N_11842);
xnor U12683 (N_12683,N_11588,N_11489);
or U12684 (N_12684,N_9471,N_9565);
nor U12685 (N_12685,N_9284,N_9986);
or U12686 (N_12686,N_11250,N_10382);
nand U12687 (N_12687,N_12474,N_7792);
nand U12688 (N_12688,N_7138,N_8369);
and U12689 (N_12689,N_10476,N_12106);
and U12690 (N_12690,N_11478,N_8092);
xor U12691 (N_12691,N_10107,N_6801);
nor U12692 (N_12692,N_12142,N_9655);
xor U12693 (N_12693,N_9452,N_11568);
and U12694 (N_12694,N_9497,N_11623);
and U12695 (N_12695,N_10182,N_7149);
or U12696 (N_12696,N_10497,N_7717);
or U12697 (N_12697,N_12226,N_8013);
nor U12698 (N_12698,N_7443,N_9788);
or U12699 (N_12699,N_6631,N_10272);
nand U12700 (N_12700,N_8183,N_10183);
nand U12701 (N_12701,N_6419,N_8918);
or U12702 (N_12702,N_10259,N_9338);
and U12703 (N_12703,N_10319,N_11945);
nand U12704 (N_12704,N_6438,N_8802);
nand U12705 (N_12705,N_8940,N_9803);
xor U12706 (N_12706,N_6903,N_6901);
and U12707 (N_12707,N_11423,N_11039);
or U12708 (N_12708,N_12022,N_10938);
nor U12709 (N_12709,N_6997,N_8367);
or U12710 (N_12710,N_12021,N_8329);
xor U12711 (N_12711,N_7543,N_7240);
nand U12712 (N_12712,N_8751,N_8076);
xnor U12713 (N_12713,N_8234,N_8449);
nor U12714 (N_12714,N_10716,N_12372);
and U12715 (N_12715,N_10276,N_7767);
xnor U12716 (N_12716,N_8637,N_11913);
xnor U12717 (N_12717,N_12260,N_9339);
and U12718 (N_12718,N_7427,N_8644);
xor U12719 (N_12719,N_10585,N_10993);
and U12720 (N_12720,N_10146,N_8875);
and U12721 (N_12721,N_6308,N_8472);
and U12722 (N_12722,N_12234,N_7433);
xor U12723 (N_12723,N_8317,N_12035);
and U12724 (N_12724,N_12432,N_12266);
xnor U12725 (N_12725,N_10086,N_6795);
or U12726 (N_12726,N_12381,N_10223);
and U12727 (N_12727,N_7590,N_11332);
or U12728 (N_12728,N_10155,N_7728);
or U12729 (N_12729,N_11850,N_6730);
xnor U12730 (N_12730,N_9819,N_9696);
xor U12731 (N_12731,N_11398,N_8371);
or U12732 (N_12732,N_8064,N_6926);
and U12733 (N_12733,N_8835,N_10612);
or U12734 (N_12734,N_7868,N_6793);
nor U12735 (N_12735,N_9056,N_8007);
and U12736 (N_12736,N_10718,N_7108);
and U12737 (N_12737,N_8392,N_12433);
nand U12738 (N_12738,N_7006,N_11875);
or U12739 (N_12739,N_9200,N_8677);
and U12740 (N_12740,N_11521,N_9708);
xnor U12741 (N_12741,N_6705,N_6305);
nand U12742 (N_12742,N_8554,N_12407);
or U12743 (N_12743,N_10056,N_7366);
and U12744 (N_12744,N_11112,N_7200);
or U12745 (N_12745,N_11204,N_7881);
xnor U12746 (N_12746,N_10062,N_6568);
nand U12747 (N_12747,N_9664,N_10345);
nor U12748 (N_12748,N_8764,N_10548);
and U12749 (N_12749,N_12265,N_10522);
and U12750 (N_12750,N_7141,N_9278);
or U12751 (N_12751,N_6778,N_9032);
and U12752 (N_12752,N_11055,N_7264);
nor U12753 (N_12753,N_9905,N_7362);
xnor U12754 (N_12754,N_10307,N_8962);
nand U12755 (N_12755,N_12289,N_6519);
nor U12756 (N_12756,N_9064,N_7180);
nand U12757 (N_12757,N_6952,N_8330);
nand U12758 (N_12758,N_9781,N_9233);
nor U12759 (N_12759,N_11921,N_7994);
xor U12760 (N_12760,N_8655,N_8220);
and U12761 (N_12761,N_11894,N_8480);
or U12762 (N_12762,N_12189,N_11926);
nor U12763 (N_12763,N_10914,N_9951);
nand U12764 (N_12764,N_10616,N_7247);
and U12765 (N_12765,N_10933,N_11041);
or U12766 (N_12766,N_9214,N_11812);
and U12767 (N_12767,N_9270,N_12238);
nor U12768 (N_12768,N_8615,N_8579);
xor U12769 (N_12769,N_11168,N_7421);
nor U12770 (N_12770,N_6270,N_9322);
and U12771 (N_12771,N_9782,N_8713);
and U12772 (N_12772,N_8566,N_10168);
nor U12773 (N_12773,N_12394,N_12485);
and U12774 (N_12774,N_10171,N_9152);
and U12775 (N_12775,N_7217,N_9855);
xor U12776 (N_12776,N_8771,N_8486);
nand U12777 (N_12777,N_7559,N_6643);
xnor U12778 (N_12778,N_7897,N_8571);
or U12779 (N_12779,N_7420,N_10112);
and U12780 (N_12780,N_6984,N_11075);
nand U12781 (N_12781,N_9528,N_7954);
nor U12782 (N_12782,N_12004,N_8354);
xor U12783 (N_12783,N_8158,N_7939);
xor U12784 (N_12784,N_9013,N_10389);
and U12785 (N_12785,N_6666,N_7499);
and U12786 (N_12786,N_10744,N_8182);
xor U12787 (N_12787,N_6875,N_8295);
nor U12788 (N_12788,N_9873,N_7675);
and U12789 (N_12789,N_10336,N_10855);
nor U12790 (N_12790,N_6490,N_6737);
nor U12791 (N_12791,N_7094,N_11385);
xnor U12792 (N_12792,N_6734,N_10485);
nand U12793 (N_12793,N_6725,N_8824);
and U12794 (N_12794,N_7582,N_10071);
xnor U12795 (N_12795,N_11040,N_11111);
nor U12796 (N_12796,N_9704,N_8254);
nand U12797 (N_12797,N_10041,N_9694);
nor U12798 (N_12798,N_7875,N_11497);
xor U12799 (N_12799,N_10674,N_7855);
or U12800 (N_12800,N_7623,N_6416);
and U12801 (N_12801,N_7567,N_8462);
and U12802 (N_12802,N_8790,N_8418);
nor U12803 (N_12803,N_6577,N_7644);
nand U12804 (N_12804,N_9453,N_12061);
nand U12805 (N_12805,N_6548,N_6552);
nor U12806 (N_12806,N_7930,N_11606);
xnor U12807 (N_12807,N_10053,N_12236);
nand U12808 (N_12808,N_10153,N_9573);
nand U12809 (N_12809,N_8079,N_12263);
nor U12810 (N_12810,N_9902,N_8750);
xor U12811 (N_12811,N_10205,N_10448);
and U12812 (N_12812,N_9589,N_7116);
and U12813 (N_12813,N_8336,N_11526);
nor U12814 (N_12814,N_9129,N_11392);
nor U12815 (N_12815,N_7342,N_7056);
nor U12816 (N_12816,N_11920,N_11578);
xnor U12817 (N_12817,N_9948,N_7109);
xor U12818 (N_12818,N_9747,N_8286);
nor U12819 (N_12819,N_10926,N_9219);
xor U12820 (N_12820,N_12423,N_11981);
or U12821 (N_12821,N_10958,N_8614);
nand U12822 (N_12822,N_8575,N_6298);
or U12823 (N_12823,N_9455,N_8165);
nor U12824 (N_12824,N_8512,N_12252);
xor U12825 (N_12825,N_10279,N_8053);
nand U12826 (N_12826,N_6719,N_7002);
nand U12827 (N_12827,N_12112,N_8745);
and U12828 (N_12828,N_8393,N_7584);
or U12829 (N_12829,N_11615,N_10423);
nand U12830 (N_12830,N_12080,N_9017);
and U12831 (N_12831,N_11485,N_8353);
xor U12832 (N_12832,N_6560,N_6998);
and U12833 (N_12833,N_8334,N_9907);
and U12834 (N_12834,N_11622,N_7766);
or U12835 (N_12835,N_11880,N_7378);
nand U12836 (N_12836,N_8241,N_12287);
nor U12837 (N_12837,N_7438,N_8693);
or U12838 (N_12838,N_6300,N_12038);
xnor U12839 (N_12839,N_9970,N_9207);
nor U12840 (N_12840,N_8812,N_6827);
xor U12841 (N_12841,N_8548,N_8775);
nor U12842 (N_12842,N_9363,N_9180);
or U12843 (N_12843,N_11603,N_10547);
xnor U12844 (N_12844,N_11239,N_8699);
nor U12845 (N_12845,N_9103,N_12196);
and U12846 (N_12846,N_11378,N_11661);
xnor U12847 (N_12847,N_11590,N_11209);
nor U12848 (N_12848,N_9869,N_7919);
nor U12849 (N_12849,N_10859,N_8466);
nand U12850 (N_12850,N_12169,N_11547);
nand U12851 (N_12851,N_9895,N_8303);
xnor U12852 (N_12852,N_9195,N_6936);
xor U12853 (N_12853,N_7091,N_9634);
or U12854 (N_12854,N_8652,N_7194);
nor U12855 (N_12855,N_12245,N_8881);
or U12856 (N_12856,N_7296,N_9809);
nor U12857 (N_12857,N_7970,N_7945);
nand U12858 (N_12858,N_6259,N_10328);
xor U12859 (N_12859,N_11899,N_6671);
nor U12860 (N_12860,N_8219,N_11903);
and U12861 (N_12861,N_8889,N_12043);
and U12862 (N_12862,N_9369,N_12497);
and U12863 (N_12863,N_11033,N_9347);
xor U12864 (N_12864,N_10057,N_6918);
or U12865 (N_12865,N_12357,N_12235);
nand U12866 (N_12866,N_8278,N_12200);
xor U12867 (N_12867,N_10246,N_10874);
xnor U12868 (N_12868,N_6444,N_11273);
xor U12869 (N_12869,N_10841,N_8756);
or U12870 (N_12870,N_8916,N_9742);
xnor U12871 (N_12871,N_7348,N_11820);
nor U12872 (N_12872,N_7469,N_12132);
nor U12873 (N_12873,N_11563,N_8109);
and U12874 (N_12874,N_10587,N_10528);
or U12875 (N_12875,N_12133,N_10304);
nor U12876 (N_12876,N_10293,N_11207);
xnor U12877 (N_12877,N_12389,N_8215);
nor U12878 (N_12878,N_10862,N_7066);
and U12879 (N_12879,N_9976,N_6370);
and U12880 (N_12880,N_7197,N_11410);
nand U12881 (N_12881,N_8935,N_11546);
and U12882 (N_12882,N_8149,N_9641);
and U12883 (N_12883,N_8854,N_8869);
nand U12884 (N_12884,N_11218,N_11984);
nand U12885 (N_12885,N_8719,N_10046);
nand U12886 (N_12886,N_6819,N_11421);
or U12887 (N_12887,N_9351,N_11270);
xnor U12888 (N_12888,N_9568,N_6815);
and U12889 (N_12889,N_9631,N_10706);
and U12890 (N_12890,N_8826,N_9654);
or U12891 (N_12891,N_11464,N_11954);
or U12892 (N_12892,N_9466,N_10531);
and U12893 (N_12893,N_6349,N_8990);
and U12894 (N_12894,N_6976,N_9957);
nor U12895 (N_12895,N_7226,N_11581);
nand U12896 (N_12896,N_7990,N_11147);
or U12897 (N_12897,N_11627,N_11980);
xor U12898 (N_12898,N_6554,N_10947);
nor U12899 (N_12899,N_6604,N_10130);
or U12900 (N_12900,N_12451,N_8185);
xor U12901 (N_12901,N_7621,N_12361);
nand U12902 (N_12902,N_6545,N_6787);
nand U12903 (N_12903,N_8619,N_9806);
xor U12904 (N_12904,N_7212,N_7493);
nor U12905 (N_12905,N_6258,N_12487);
nor U12906 (N_12906,N_8526,N_8148);
nor U12907 (N_12907,N_10280,N_7324);
nor U12908 (N_12908,N_7353,N_9019);
or U12909 (N_12909,N_12382,N_11038);
and U12910 (N_12910,N_7049,N_11825);
and U12911 (N_12911,N_7459,N_6514);
nand U12912 (N_12912,N_12084,N_8269);
and U12913 (N_12913,N_6880,N_6381);
or U12914 (N_12914,N_10106,N_9204);
or U12915 (N_12915,N_10294,N_7351);
nor U12916 (N_12916,N_10872,N_6335);
and U12917 (N_12917,N_11657,N_11746);
or U12918 (N_12918,N_12442,N_8202);
nand U12919 (N_12919,N_8805,N_9831);
nor U12920 (N_12920,N_12162,N_10063);
xor U12921 (N_12921,N_7512,N_8281);
nor U12922 (N_12922,N_10663,N_7064);
and U12923 (N_12923,N_10537,N_7516);
nand U12924 (N_12924,N_9712,N_12431);
and U12925 (N_12925,N_11751,N_8908);
and U12926 (N_12926,N_12116,N_8414);
nand U12927 (N_12927,N_11967,N_6260);
xor U12928 (N_12928,N_7318,N_7276);
and U12929 (N_12929,N_11745,N_10868);
xor U12930 (N_12930,N_10305,N_11821);
xnor U12931 (N_12931,N_7622,N_8957);
nand U12932 (N_12932,N_9285,N_7003);
and U12933 (N_12933,N_12015,N_9419);
nor U12934 (N_12934,N_11794,N_8905);
nor U12935 (N_12935,N_6594,N_6414);
or U12936 (N_12936,N_6731,N_10602);
and U12937 (N_12937,N_12490,N_7656);
nand U12938 (N_12938,N_8850,N_7417);
and U12939 (N_12939,N_12447,N_8791);
nor U12940 (N_12940,N_10095,N_11916);
xnor U12941 (N_12941,N_11817,N_9765);
xnor U12942 (N_12942,N_8729,N_6518);
xnor U12943 (N_12943,N_9527,N_8314);
nor U12944 (N_12944,N_7008,N_11721);
or U12945 (N_12945,N_10883,N_6376);
nand U12946 (N_12946,N_8255,N_6842);
nand U12947 (N_12947,N_7839,N_12092);
or U12948 (N_12948,N_11712,N_9893);
nor U12949 (N_12949,N_6838,N_8288);
and U12950 (N_12950,N_12445,N_9596);
nor U12951 (N_12951,N_12013,N_6826);
nand U12952 (N_12952,N_10457,N_7748);
or U12953 (N_12953,N_11407,N_12180);
xor U12954 (N_12954,N_11659,N_11937);
nor U12955 (N_12955,N_7445,N_9228);
xor U12956 (N_12956,N_12171,N_7385);
nand U12957 (N_12957,N_7770,N_8774);
and U12958 (N_12958,N_9084,N_9795);
nor U12959 (N_12959,N_8181,N_9458);
nor U12960 (N_12960,N_8271,N_7029);
xnor U12961 (N_12961,N_7805,N_10592);
nor U12962 (N_12962,N_8999,N_9237);
and U12963 (N_12963,N_10979,N_10218);
or U12964 (N_12964,N_10473,N_10264);
xnor U12965 (N_12965,N_12340,N_9894);
or U12966 (N_12966,N_8435,N_10144);
xnor U12967 (N_12967,N_10747,N_9311);
or U12968 (N_12968,N_11679,N_11572);
xnor U12969 (N_12969,N_12410,N_9814);
nor U12970 (N_12970,N_7746,N_7992);
and U12971 (N_12971,N_10055,N_10972);
and U12972 (N_12972,N_12194,N_6649);
and U12973 (N_12973,N_12262,N_9151);
and U12974 (N_12974,N_11691,N_12393);
nand U12975 (N_12975,N_10885,N_7078);
xnor U12976 (N_12976,N_10136,N_12058);
or U12977 (N_12977,N_8145,N_9389);
nand U12978 (N_12978,N_7038,N_9744);
and U12979 (N_12979,N_8504,N_9102);
and U12980 (N_12980,N_11399,N_11676);
xor U12981 (N_12981,N_6434,N_8767);
xnor U12982 (N_12982,N_11003,N_12250);
xnor U12983 (N_12983,N_8089,N_11415);
or U12984 (N_12984,N_10580,N_10179);
nor U12985 (N_12985,N_10460,N_7525);
nor U12986 (N_12986,N_9952,N_9181);
nor U12987 (N_12987,N_10776,N_9871);
nand U12988 (N_12988,N_8597,N_8996);
and U12989 (N_12989,N_8600,N_11989);
and U12990 (N_12990,N_7854,N_12375);
or U12991 (N_12991,N_10743,N_9063);
nand U12992 (N_12992,N_9688,N_9822);
nand U12993 (N_12993,N_9891,N_9316);
xor U12994 (N_12994,N_6462,N_8721);
nor U12995 (N_12995,N_7153,N_10777);
xor U12996 (N_12996,N_9569,N_7549);
nor U12997 (N_12997,N_9736,N_8636);
or U12998 (N_12998,N_11626,N_11100);
or U12999 (N_12999,N_8839,N_8638);
nor U13000 (N_13000,N_11517,N_7743);
and U13001 (N_13001,N_9731,N_11238);
and U13002 (N_13002,N_8177,N_9360);
or U13003 (N_13003,N_7418,N_8685);
and U13004 (N_13004,N_8167,N_12025);
xor U13005 (N_13005,N_9114,N_7882);
nand U13006 (N_13006,N_10772,N_10715);
xor U13007 (N_13007,N_10826,N_9239);
nand U13008 (N_13008,N_11470,N_11885);
xor U13009 (N_13009,N_6293,N_6417);
and U13010 (N_13010,N_11405,N_10245);
xnor U13011 (N_13011,N_8351,N_11923);
nand U13012 (N_13012,N_10364,N_11577);
nor U13013 (N_13013,N_12175,N_9273);
and U13014 (N_13014,N_7092,N_6517);
nor U13015 (N_13015,N_6667,N_7437);
xor U13016 (N_13016,N_11837,N_12037);
or U13017 (N_13017,N_10684,N_6250);
nand U13018 (N_13018,N_7537,N_11356);
or U13019 (N_13019,N_7471,N_9955);
and U13020 (N_13020,N_8405,N_11066);
or U13021 (N_13021,N_8929,N_6862);
xor U13022 (N_13022,N_11741,N_7759);
xnor U13023 (N_13023,N_8930,N_8104);
xor U13024 (N_13024,N_9150,N_7942);
xnor U13025 (N_13025,N_10517,N_8716);
and U13026 (N_13026,N_12183,N_8591);
nor U13027 (N_13027,N_11299,N_9121);
nand U13028 (N_13028,N_7997,N_7098);
or U13029 (N_13029,N_9909,N_6642);
nor U13030 (N_13030,N_10969,N_9140);
nor U13031 (N_13031,N_7878,N_12450);
xnor U13032 (N_13032,N_9035,N_8552);
nor U13033 (N_13033,N_10839,N_11424);
xnor U13034 (N_13034,N_8787,N_10285);
and U13035 (N_13035,N_10240,N_7504);
xor U13036 (N_13036,N_8862,N_6358);
nor U13037 (N_13037,N_6934,N_10992);
xor U13038 (N_13038,N_8506,N_9262);
nor U13039 (N_13039,N_10093,N_9973);
nor U13040 (N_13040,N_6755,N_7012);
xnor U13041 (N_13041,N_8247,N_7659);
nand U13042 (N_13042,N_9982,N_7961);
xnor U13043 (N_13043,N_6679,N_12378);
nor U13044 (N_13044,N_11261,N_10126);
and U13045 (N_13045,N_7195,N_6878);
or U13046 (N_13046,N_6751,N_6645);
nand U13047 (N_13047,N_8150,N_8130);
xor U13048 (N_13048,N_11349,N_6411);
or U13049 (N_13049,N_10335,N_7651);
nor U13050 (N_13050,N_8428,N_12281);
and U13051 (N_13051,N_10085,N_7441);
or U13052 (N_13052,N_10017,N_12309);
and U13053 (N_13053,N_9709,N_8299);
nand U13054 (N_13054,N_7851,N_8402);
or U13055 (N_13055,N_12227,N_8922);
and U13056 (N_13056,N_9133,N_11338);
xor U13057 (N_13057,N_6938,N_8136);
xor U13058 (N_13058,N_8248,N_7876);
and U13059 (N_13059,N_8235,N_8054);
nand U13060 (N_13060,N_10598,N_11739);
nand U13061 (N_13061,N_8758,N_7949);
nand U13062 (N_13062,N_10783,N_6551);
xnor U13063 (N_13063,N_12403,N_6692);
or U13064 (N_13064,N_6461,N_7952);
xnor U13065 (N_13065,N_8634,N_7973);
nor U13066 (N_13066,N_8832,N_10466);
nand U13067 (N_13067,N_9392,N_12498);
and U13068 (N_13068,N_8338,N_7669);
nand U13069 (N_13069,N_12119,N_11368);
xnor U13070 (N_13070,N_7630,N_12098);
or U13071 (N_13071,N_6987,N_7331);
and U13072 (N_13072,N_11442,N_10242);
nor U13073 (N_13073,N_8030,N_11021);
xnor U13074 (N_13074,N_11199,N_7127);
xor U13075 (N_13075,N_10374,N_8118);
nor U13076 (N_13076,N_8495,N_10896);
or U13077 (N_13077,N_8491,N_6440);
and U13078 (N_13078,N_8788,N_8069);
nand U13079 (N_13079,N_6580,N_6471);
xnor U13080 (N_13080,N_12368,N_12048);
or U13081 (N_13081,N_10799,N_12201);
and U13082 (N_13082,N_8657,N_11234);
or U13083 (N_13083,N_11683,N_9681);
nor U13084 (N_13084,N_8821,N_12371);
or U13085 (N_13085,N_8043,N_6503);
nor U13086 (N_13086,N_11694,N_7273);
nor U13087 (N_13087,N_6437,N_9268);
nor U13088 (N_13088,N_6281,N_9555);
nand U13089 (N_13089,N_10619,N_6707);
nor U13090 (N_13090,N_9689,N_8324);
and U13091 (N_13091,N_10932,N_11727);
nor U13092 (N_13092,N_9365,N_8785);
nor U13093 (N_13093,N_11089,N_7405);
and U13094 (N_13094,N_9374,N_7277);
xnor U13095 (N_13095,N_8151,N_10769);
xnor U13096 (N_13096,N_9701,N_10780);
and U13097 (N_13097,N_6763,N_8131);
nor U13098 (N_13098,N_7001,N_8063);
nand U13099 (N_13099,N_7397,N_10614);
xor U13100 (N_13100,N_9113,N_12109);
or U13101 (N_13101,N_12049,N_11166);
xnor U13102 (N_13102,N_7918,N_6922);
xor U13103 (N_13103,N_12412,N_7369);
xor U13104 (N_13104,N_9288,N_7793);
or U13105 (N_13105,N_11345,N_11358);
or U13106 (N_13106,N_7885,N_7620);
nor U13107 (N_13107,N_7236,N_10781);
nor U13108 (N_13108,N_10065,N_9988);
nor U13109 (N_13109,N_6872,N_12223);
nand U13110 (N_13110,N_9617,N_7498);
xor U13111 (N_13111,N_12232,N_7607);
or U13112 (N_13112,N_10982,N_7395);
nor U13113 (N_13113,N_9441,N_6812);
and U13114 (N_13114,N_8965,N_7023);
and U13115 (N_13115,N_8374,N_10187);
xnor U13116 (N_13116,N_8196,N_8382);
xnor U13117 (N_13117,N_9639,N_6931);
xor U13118 (N_13118,N_11902,N_11924);
xnor U13119 (N_13119,N_11795,N_9296);
xnor U13120 (N_13120,N_6288,N_10467);
and U13121 (N_13121,N_10611,N_7210);
nand U13122 (N_13122,N_7964,N_7139);
or U13123 (N_13123,N_10644,N_6791);
or U13124 (N_13124,N_8059,N_8949);
or U13125 (N_13125,N_8081,N_10202);
and U13126 (N_13126,N_11011,N_7235);
nand U13127 (N_13127,N_7455,N_7466);
xor U13128 (N_13128,N_11276,N_10924);
and U13129 (N_13129,N_8070,N_7654);
and U13130 (N_13130,N_8722,N_11524);
nor U13131 (N_13131,N_9549,N_8557);
nor U13132 (N_13132,N_6385,N_6553);
nand U13133 (N_13133,N_9944,N_10724);
nand U13134 (N_13134,N_9029,N_8328);
nor U13135 (N_13135,N_11439,N_6694);
and U13136 (N_13136,N_10621,N_7794);
xnor U13137 (N_13137,N_11069,N_12458);
or U13138 (N_13138,N_6702,N_8433);
xnor U13139 (N_13139,N_8503,N_11990);
or U13140 (N_13140,N_7531,N_7753);
xor U13141 (N_13141,N_9154,N_9227);
nand U13142 (N_13142,N_8911,N_11427);
nand U13143 (N_13143,N_8800,N_10058);
nor U13144 (N_13144,N_7747,N_11516);
xor U13145 (N_13145,N_6797,N_6467);
nand U13146 (N_13146,N_8147,N_7920);
and U13147 (N_13147,N_10301,N_11327);
and U13148 (N_13148,N_8683,N_10834);
and U13149 (N_13149,N_10311,N_11579);
nand U13150 (N_13150,N_9033,N_7173);
xnor U13151 (N_13151,N_11966,N_10764);
nor U13152 (N_13152,N_10596,N_7249);
or U13153 (N_13153,N_7400,N_9653);
nand U13154 (N_13154,N_7464,N_8819);
nor U13155 (N_13155,N_10569,N_7435);
nand U13156 (N_13156,N_9123,N_11330);
nand U13157 (N_13157,N_6965,N_7227);
and U13158 (N_13158,N_11791,N_8541);
nor U13159 (N_13159,N_8168,N_10641);
xor U13160 (N_13160,N_6448,N_7616);
or U13161 (N_13161,N_6673,N_8419);
xnor U13162 (N_13162,N_11495,N_11929);
or U13163 (N_13163,N_10077,N_6953);
nor U13164 (N_13164,N_7382,N_6299);
nand U13165 (N_13165,N_11036,N_11738);
nand U13166 (N_13166,N_10356,N_12231);
or U13167 (N_13167,N_8776,N_10990);
nor U13168 (N_13168,N_8671,N_6665);
xor U13169 (N_13169,N_9104,N_11977);
nor U13170 (N_13170,N_8842,N_7606);
nor U13171 (N_13171,N_10266,N_7311);
nor U13172 (N_13172,N_10231,N_9126);
xor U13173 (N_13173,N_10355,N_9861);
nor U13174 (N_13174,N_7332,N_9849);
nand U13175 (N_13175,N_11205,N_9485);
and U13176 (N_13176,N_9661,N_7915);
nand U13177 (N_13177,N_9718,N_12207);
nand U13178 (N_13178,N_8163,N_6392);
nor U13179 (N_13179,N_8992,N_8068);
and U13180 (N_13180,N_7515,N_6276);
xor U13181 (N_13181,N_11472,N_6764);
or U13182 (N_13182,N_8058,N_8768);
nand U13183 (N_13183,N_12352,N_12029);
xor U13184 (N_13184,N_7252,N_9906);
nand U13185 (N_13185,N_12473,N_12020);
or U13186 (N_13186,N_6502,N_11811);
xnor U13187 (N_13187,N_12154,N_8471);
or U13188 (N_13188,N_11265,N_8956);
xor U13189 (N_13189,N_7929,N_7520);
or U13190 (N_13190,N_9772,N_8062);
and U13191 (N_13191,N_11437,N_7645);
and U13192 (N_13192,N_7694,N_10950);
xor U13193 (N_13193,N_7473,N_12007);
nor U13194 (N_13194,N_8432,N_8340);
and U13195 (N_13195,N_8892,N_9840);
nor U13196 (N_13196,N_11674,N_7823);
nor U13197 (N_13197,N_11973,N_7609);
xnor U13198 (N_13198,N_9002,N_7491);
nor U13199 (N_13199,N_9610,N_9558);
xor U13200 (N_13200,N_8789,N_7733);
and U13201 (N_13201,N_10125,N_11188);
nor U13202 (N_13202,N_9959,N_11591);
and U13203 (N_13203,N_10639,N_11068);
nand U13204 (N_13204,N_8725,N_9890);
and U13205 (N_13205,N_11303,N_11198);
and U13206 (N_13206,N_10928,N_10133);
nor U13207 (N_13207,N_9752,N_10828);
nand U13208 (N_13208,N_7019,N_9067);
or U13209 (N_13209,N_6352,N_9514);
or U13210 (N_13210,N_11633,N_11670);
and U13211 (N_13211,N_11200,N_8621);
nand U13212 (N_13212,N_11797,N_9131);
nor U13213 (N_13213,N_8766,N_9095);
nor U13214 (N_13214,N_8375,N_7082);
xnor U13215 (N_13215,N_6920,N_10271);
and U13216 (N_13216,N_9174,N_9279);
nor U13217 (N_13217,N_12079,N_10786);
or U13218 (N_13218,N_10273,N_10925);
nor U13219 (N_13219,N_9647,N_6309);
xor U13220 (N_13220,N_7678,N_8451);
xnor U13221 (N_13221,N_7642,N_11030);
and U13222 (N_13222,N_10419,N_8675);
xor U13223 (N_13223,N_11027,N_7726);
nor U13224 (N_13224,N_6436,N_6961);
xnor U13225 (N_13225,N_9990,N_7199);
nor U13226 (N_13226,N_11714,N_10590);
or U13227 (N_13227,N_7365,N_9864);
and U13228 (N_13228,N_7900,N_7937);
and U13229 (N_13229,N_7463,N_8741);
xnor U13230 (N_13230,N_9832,N_12128);
and U13231 (N_13231,N_7844,N_11447);
and U13232 (N_13232,N_8702,N_11700);
and U13233 (N_13233,N_10844,N_7022);
xnor U13234 (N_13234,N_6617,N_11816);
nand U13235 (N_13235,N_7398,N_12468);
and U13236 (N_13236,N_7144,N_9954);
or U13237 (N_13237,N_6945,N_12193);
nand U13238 (N_13238,N_10848,N_11834);
xnor U13239 (N_13239,N_11096,N_8395);
nor U13240 (N_13240,N_6696,N_9345);
nor U13241 (N_13241,N_7535,N_9478);
or U13242 (N_13242,N_7279,N_6585);
xor U13243 (N_13243,N_8966,N_9760);
or U13244 (N_13244,N_9543,N_11046);
nand U13245 (N_13245,N_8140,N_7858);
and U13246 (N_13246,N_8632,N_11583);
nand U13247 (N_13247,N_8270,N_9036);
xor U13248 (N_13248,N_12421,N_12429);
or U13249 (N_13249,N_10652,N_6491);
or U13250 (N_13250,N_8474,N_9564);
nor U13251 (N_13251,N_11697,N_8006);
or U13252 (N_13252,N_9381,N_11719);
and U13253 (N_13253,N_8626,N_8696);
nand U13254 (N_13254,N_8678,N_9234);
and U13255 (N_13255,N_10066,N_6632);
and U13256 (N_13256,N_8761,N_6321);
nand U13257 (N_13257,N_9758,N_8128);
nor U13258 (N_13258,N_10720,N_9624);
nand U13259 (N_13259,N_10392,N_9510);
nand U13260 (N_13260,N_11660,N_9813);
nor U13261 (N_13261,N_11394,N_8452);
xor U13262 (N_13262,N_6728,N_12060);
xnor U13263 (N_13263,N_9935,N_9092);
and U13264 (N_13264,N_9326,N_8291);
nor U13265 (N_13265,N_12158,N_10464);
nand U13266 (N_13266,N_12302,N_10359);
or U13267 (N_13267,N_10409,N_7570);
or U13268 (N_13268,N_11859,N_7458);
nand U13269 (N_13269,N_9079,N_9111);
xor U13270 (N_13270,N_7765,N_12164);
and U13271 (N_13271,N_10515,N_6888);
or U13272 (N_13272,N_8169,N_6255);
nand U13273 (N_13273,N_8047,N_6943);
nor U13274 (N_13274,N_11316,N_9616);
and U13275 (N_13275,N_12455,N_11409);
nor U13276 (N_13276,N_7615,N_9542);
xnor U13277 (N_13277,N_8294,N_7172);
or U13278 (N_13278,N_7523,N_12233);
nand U13279 (N_13279,N_9287,N_11469);
nand U13280 (N_13280,N_11256,N_11490);
or U13281 (N_13281,N_9811,N_6521);
and U13282 (N_13282,N_6323,N_9050);
xnor U13283 (N_13283,N_11004,N_6988);
nor U13284 (N_13284,N_11049,N_11814);
xnor U13285 (N_13285,N_10478,N_9128);
nand U13286 (N_13286,N_9604,N_11584);
nand U13287 (N_13287,N_8733,N_11974);
and U13288 (N_13288,N_8620,N_7286);
xor U13289 (N_13289,N_7734,N_11451);
nor U13290 (N_13290,N_7916,N_9550);
xnor U13291 (N_13291,N_10292,N_7222);
nand U13292 (N_13292,N_10757,N_11760);
and U13293 (N_13293,N_7253,N_6595);
nor U13294 (N_13294,N_12439,N_10986);
nand U13295 (N_13295,N_8040,N_10108);
and U13296 (N_13296,N_10349,N_6829);
nor U13297 (N_13297,N_10369,N_11189);
nor U13298 (N_13298,N_11566,N_10454);
and U13299 (N_13299,N_6403,N_11689);
nand U13300 (N_13300,N_8553,N_10350);
nand U13301 (N_13301,N_9054,N_7699);
nor U13302 (N_13302,N_11611,N_6410);
and U13303 (N_13303,N_9580,N_6488);
or U13304 (N_13304,N_12184,N_6395);
nor U13305 (N_13305,N_9335,N_10850);
and U13306 (N_13306,N_10411,N_9852);
or U13307 (N_13307,N_11210,N_10991);
and U13308 (N_13308,N_9784,N_9016);
xor U13309 (N_13309,N_10227,N_7140);
and U13310 (N_13310,N_6333,N_6735);
nor U13311 (N_13311,N_9798,N_9612);
nand U13312 (N_13312,N_8460,N_10498);
nor U13313 (N_13313,N_7796,N_7036);
nand U13314 (N_13314,N_7752,N_11465);
xor U13315 (N_13315,N_11151,N_9483);
xnor U13316 (N_13316,N_10734,N_9446);
nand U13317 (N_13317,N_9281,N_7658);
nand U13318 (N_13318,N_11197,N_10995);
xor U13319 (N_13319,N_7715,N_10956);
or U13320 (N_13320,N_7781,N_10221);
xnor U13321 (N_13321,N_8646,N_7697);
and U13322 (N_13322,N_11224,N_7457);
nor U13323 (N_13323,N_9775,N_11955);
nor U13324 (N_13324,N_7202,N_11482);
nor U13325 (N_13325,N_9266,N_7596);
or U13326 (N_13326,N_11050,N_9996);
or U13327 (N_13327,N_9457,N_8251);
xnor U13328 (N_13328,N_9314,N_9025);
nand U13329 (N_13329,N_6832,N_10383);
xor U13330 (N_13330,N_7234,N_9354);
or U13331 (N_13331,N_6558,N_11170);
nor U13332 (N_13332,N_10282,N_8468);
nand U13333 (N_13333,N_9160,N_6322);
nand U13334 (N_13334,N_10503,N_9094);
nor U13335 (N_13335,N_9498,N_6973);
nand U13336 (N_13336,N_9985,N_6421);
or U13337 (N_13337,N_6777,N_11844);
and U13338 (N_13338,N_10237,N_7377);
and U13339 (N_13339,N_7995,N_8743);
nand U13340 (N_13340,N_6909,N_11278);
or U13341 (N_13341,N_7721,N_10594);
xor U13342 (N_13342,N_9677,N_6955);
or U13343 (N_13343,N_10083,N_7763);
nor U13344 (N_13344,N_10748,N_7711);
and U13345 (N_13345,N_7161,N_7806);
and U13346 (N_13346,N_9521,N_11319);
and U13347 (N_13347,N_9062,N_10243);
or U13348 (N_13348,N_6261,N_8098);
nand U13349 (N_13349,N_11462,N_7779);
or U13350 (N_13350,N_9317,N_11688);
nand U13351 (N_13351,N_7978,N_7164);
or U13352 (N_13352,N_7160,N_9073);
xnor U13353 (N_13353,N_9899,N_10818);
or U13354 (N_13354,N_12187,N_11684);
xnor U13355 (N_13355,N_6498,N_12286);
nand U13356 (N_13356,N_8963,N_8072);
nor U13357 (N_13357,N_8568,N_11770);
xor U13358 (N_13358,N_10660,N_11266);
xnor U13359 (N_13359,N_6387,N_9727);
nor U13360 (N_13360,N_9559,N_8598);
nand U13361 (N_13361,N_10094,N_10714);
nor U13362 (N_13362,N_10553,N_9229);
xor U13363 (N_13363,N_9678,N_7232);
or U13364 (N_13364,N_10858,N_6773);
and U13365 (N_13365,N_11793,N_6779);
nor U13366 (N_13366,N_10860,N_8993);
xor U13367 (N_13367,N_11778,N_8263);
and U13368 (N_13368,N_7111,N_10474);
xor U13369 (N_13369,N_7758,N_7442);
nor U13370 (N_13370,N_11263,N_12188);
xnor U13371 (N_13371,N_11852,N_10667);
nand U13372 (N_13372,N_7467,N_12271);
nand U13373 (N_13373,N_7732,N_12307);
xor U13374 (N_13374,N_9272,N_10973);
nand U13375 (N_13375,N_12185,N_11082);
and U13376 (N_13376,N_6974,N_8133);
xnor U13377 (N_13377,N_10194,N_11325);
and U13378 (N_13378,N_10816,N_9225);
or U13379 (N_13379,N_12385,N_10853);
and U13380 (N_13380,N_9099,N_12258);
or U13381 (N_13381,N_9526,N_9490);
xnor U13382 (N_13382,N_11702,N_11726);
nand U13383 (N_13383,N_10324,N_6907);
xnor U13384 (N_13384,N_9577,N_11160);
and U13385 (N_13385,N_10730,N_7333);
xor U13386 (N_13386,N_11500,N_7987);
xor U13387 (N_13387,N_7518,N_7635);
and U13388 (N_13388,N_11949,N_8806);
or U13389 (N_13389,N_6361,N_7483);
nor U13390 (N_13390,N_12489,N_7484);
nor U13391 (N_13391,N_7026,N_11766);
and U13392 (N_13392,N_10494,N_11513);
xnor U13393 (N_13393,N_6584,N_7556);
nor U13394 (N_13394,N_9937,N_8917);
nor U13395 (N_13395,N_11888,N_11217);
and U13396 (N_13396,N_9672,N_8455);
nand U13397 (N_13397,N_9828,N_11087);
or U13398 (N_13398,N_8225,N_6317);
or U13399 (N_13399,N_11971,N_10889);
or U13400 (N_13400,N_12240,N_7047);
or U13401 (N_13401,N_9821,N_12253);
or U13402 (N_13402,N_6766,N_9193);
and U13403 (N_13403,N_10193,N_6546);
xnor U13404 (N_13404,N_6315,N_8213);
and U13405 (N_13405,N_11122,N_9725);
nand U13406 (N_13406,N_10627,N_7709);
xnor U13407 (N_13407,N_6318,N_10395);
nand U13408 (N_13408,N_12273,N_6515);
nor U13409 (N_13409,N_9729,N_8509);
nand U13410 (N_13410,N_7832,N_10918);
and U13411 (N_13411,N_10137,N_6265);
xor U13412 (N_13412,N_8577,N_8273);
or U13413 (N_13413,N_10763,N_12255);
nand U13414 (N_13414,N_6754,N_8772);
and U13415 (N_13415,N_12369,N_10472);
or U13416 (N_13416,N_6635,N_6597);
and U13417 (N_13417,N_9156,N_12366);
xnor U13418 (N_13418,N_10977,N_9646);
xor U13419 (N_13419,N_10575,N_10555);
and U13420 (N_13420,N_11705,N_9201);
and U13421 (N_13421,N_7568,N_7143);
and U13422 (N_13422,N_11907,N_7534);
nor U13423 (N_13423,N_10631,N_10018);
xor U13424 (N_13424,N_10778,N_7123);
or U13425 (N_13425,N_12115,N_11313);
xnor U13426 (N_13426,N_10249,N_9342);
nor U13427 (N_13427,N_7099,N_7071);
nor U13428 (N_13428,N_10750,N_8322);
nand U13429 (N_13429,N_8349,N_6363);
nand U13430 (N_13430,N_8229,N_12288);
and U13431 (N_13431,N_6788,N_12383);
nor U13432 (N_13432,N_7863,N_7363);
nor U13433 (N_13433,N_9505,N_7852);
xor U13434 (N_13434,N_11713,N_6640);
xnor U13435 (N_13435,N_9306,N_8510);
nor U13436 (N_13436,N_7309,N_6290);
or U13437 (N_13437,N_6656,N_7600);
xnor U13438 (N_13438,N_12479,N_10483);
nand U13439 (N_13439,N_7048,N_8648);
or U13440 (N_13440,N_6536,N_9045);
xor U13441 (N_13441,N_11527,N_10197);
and U13442 (N_13442,N_10479,N_10007);
nand U13443 (N_13443,N_9364,N_9393);
or U13444 (N_13444,N_10358,N_9732);
and U13445 (N_13445,N_8786,N_8009);
and U13446 (N_13446,N_11123,N_11347);
or U13447 (N_13447,N_10213,N_10901);
and U13448 (N_13448,N_11722,N_9068);
or U13449 (N_13449,N_11120,N_6647);
xor U13450 (N_13450,N_9286,N_10910);
xnor U13451 (N_13451,N_9683,N_7722);
and U13452 (N_13452,N_8641,N_7546);
nor U13453 (N_13453,N_8236,N_8154);
nand U13454 (N_13454,N_11541,N_10045);
and U13455 (N_13455,N_11286,N_7406);
or U13456 (N_13456,N_12397,N_9908);
nand U13457 (N_13457,N_7102,N_8860);
xor U13458 (N_13458,N_11461,N_10980);
nor U13459 (N_13459,N_8549,N_7502);
xor U13460 (N_13460,N_9173,N_10898);
nor U13461 (N_13461,N_6264,N_7215);
nand U13462 (N_13462,N_11988,N_8381);
and U13463 (N_13463,N_10811,N_9774);
or U13464 (N_13464,N_7216,N_7361);
or U13465 (N_13465,N_7224,N_8034);
xor U13466 (N_13466,N_11397,N_10882);
and U13467 (N_13467,N_10604,N_11861);
xnor U13468 (N_13468,N_12144,N_10767);
nor U13469 (N_13469,N_12460,N_11843);
nand U13470 (N_13470,N_8523,N_11379);
nand U13471 (N_13471,N_10875,N_9325);
nor U13472 (N_13472,N_10698,N_9685);
nand U13473 (N_13473,N_8705,N_10725);
or U13474 (N_13474,N_7394,N_11109);
nand U13475 (N_13475,N_9815,N_6925);
nand U13476 (N_13476,N_6480,N_7856);
xnor U13477 (N_13477,N_8478,N_10584);
and U13478 (N_13478,N_7889,N_10038);
xnor U13479 (N_13479,N_10209,N_8623);
or U13480 (N_13480,N_10299,N_7104);
nor U13481 (N_13481,N_7039,N_7810);
nand U13482 (N_13482,N_10190,N_9875);
and U13483 (N_13483,N_7243,N_10427);
xor U13484 (N_13484,N_6808,N_9611);
nand U13485 (N_13485,N_10968,N_7522);
xnor U13486 (N_13486,N_6327,N_9435);
and U13487 (N_13487,N_7344,N_10260);
nand U13488 (N_13488,N_6772,N_9865);
xnor U13489 (N_13489,N_9240,N_9773);
and U13490 (N_13490,N_8681,N_11202);
nand U13491 (N_13491,N_6520,N_6418);
or U13492 (N_13492,N_8560,N_12401);
or U13493 (N_13493,N_8617,N_10103);
nor U13494 (N_13494,N_12331,N_12241);
xor U13495 (N_13495,N_7490,N_12338);
and U13496 (N_13496,N_7220,N_10525);
xor U13497 (N_13497,N_8025,N_10297);
nor U13498 (N_13498,N_7936,N_9249);
and U13499 (N_13499,N_7052,N_11156);
and U13500 (N_13500,N_9605,N_11386);
and U13501 (N_13501,N_11413,N_7756);
nand U13502 (N_13502,N_11395,N_8746);
and U13503 (N_13503,N_9139,N_10079);
or U13504 (N_13504,N_12089,N_11787);
nand U13505 (N_13505,N_8000,N_7291);
and U13506 (N_13506,N_6916,N_10054);
or U13507 (N_13507,N_7335,N_7814);
or U13508 (N_13508,N_10325,N_11621);
and U13509 (N_13509,N_7170,N_9845);
xor U13510 (N_13510,N_8603,N_10921);
and U13511 (N_13511,N_9178,N_12492);
or U13512 (N_13512,N_8188,N_8493);
and U13513 (N_13513,N_7121,N_11154);
nand U13514 (N_13514,N_10465,N_7601);
and U13515 (N_13515,N_10633,N_10987);
xor U13516 (N_13516,N_6848,N_11826);
nand U13517 (N_13517,N_9172,N_9294);
nor U13518 (N_13518,N_6409,N_10996);
nor U13519 (N_13519,N_11771,N_9987);
and U13520 (N_13520,N_6271,N_6402);
and U13521 (N_13521,N_12285,N_10845);
nor U13522 (N_13522,N_12329,N_6563);
xnor U13523 (N_13523,N_11420,N_8487);
nand U13524 (N_13524,N_12210,N_10662);
or U13525 (N_13525,N_12409,N_9627);
nor U13526 (N_13526,N_9158,N_12476);
xnor U13527 (N_13527,N_6497,N_8700);
or U13528 (N_13528,N_11881,N_10163);
or U13529 (N_13529,N_9343,N_7737);
nand U13530 (N_13530,N_10224,N_10373);
or U13531 (N_13531,N_9182,N_11149);
xnor U13532 (N_13532,N_9475,N_11494);
nand U13533 (N_13533,N_11650,N_8679);
or U13534 (N_13534,N_10352,N_8519);
nor U13535 (N_13535,N_11690,N_11419);
nand U13536 (N_13536,N_7087,N_10005);
nor U13537 (N_13537,N_7610,N_10151);
or U13538 (N_13538,N_7462,N_11201);
nand U13539 (N_13539,N_12046,N_10043);
and U13540 (N_13540,N_6944,N_6720);
or U13541 (N_13541,N_9785,N_11110);
or U13542 (N_13542,N_9733,N_9829);
nand U13543 (N_13543,N_7131,N_9297);
and U13544 (N_13544,N_9238,N_11790);
and U13545 (N_13545,N_7634,N_6579);
nand U13546 (N_13546,N_9846,N_12002);
xnor U13547 (N_13547,N_11783,N_8099);
or U13548 (N_13548,N_8115,N_8578);
or U13549 (N_13549,N_11233,N_12006);
nand U13550 (N_13550,N_10229,N_9805);
xnor U13551 (N_13551,N_9046,N_7157);
nor U13552 (N_13552,N_6646,N_7496);
nor U13553 (N_13553,N_12087,N_7864);
xor U13554 (N_13554,N_10100,N_6835);
and U13555 (N_13555,N_8342,N_6329);
xnor U13556 (N_13556,N_8376,N_12168);
nand U13557 (N_13557,N_6981,N_8714);
or U13558 (N_13558,N_10495,N_11501);
nand U13559 (N_13559,N_10562,N_7815);
xnor U13560 (N_13560,N_11802,N_11088);
nand U13561 (N_13561,N_6435,N_7695);
nand U13562 (N_13562,N_6415,N_8228);
xor U13563 (N_13563,N_11716,N_6574);
nand U13564 (N_13564,N_7129,N_11932);
xnor U13565 (N_13565,N_11035,N_8184);
and U13566 (N_13566,N_6481,N_12028);
and U13567 (N_13567,N_10940,N_11835);
nor U13568 (N_13568,N_6459,N_12488);
and U13569 (N_13569,N_8267,N_11296);
nand U13570 (N_13570,N_7412,N_10453);
xnor U13571 (N_13571,N_11017,N_7241);
xor U13572 (N_13572,N_10320,N_10384);
nand U13573 (N_13573,N_7323,N_7128);
xor U13574 (N_13574,N_6278,N_12446);
or U13575 (N_13575,N_7339,N_11534);
or U13576 (N_13576,N_10251,N_8910);
and U13577 (N_13577,N_9188,N_6959);
and U13578 (N_13578,N_7983,N_7135);
and U13579 (N_13579,N_6253,N_9076);
or U13580 (N_13580,N_7085,N_10201);
nand U13581 (N_13581,N_10541,N_9945);
nor U13582 (N_13582,N_10854,N_8627);
xor U13583 (N_13583,N_11257,N_11280);
nor U13584 (N_13584,N_8218,N_6499);
and U13585 (N_13585,N_8123,N_11435);
xor U13586 (N_13586,N_12070,N_7414);
xnor U13587 (N_13587,N_9721,N_10135);
nand U13588 (N_13588,N_8172,N_8018);
or U13589 (N_13589,N_9315,N_11215);
xor U13590 (N_13590,N_10681,N_6332);
nand U13591 (N_13591,N_7179,N_8540);
xor U13592 (N_13592,N_10312,N_12001);
xnor U13593 (N_13593,N_6319,N_10691);
or U13594 (N_13594,N_7494,N_11306);
nand U13595 (N_13595,N_9977,N_9686);
or U13596 (N_13596,N_6978,N_8613);
nor U13597 (N_13597,N_7729,N_8664);
and U13598 (N_13598,N_7740,N_10909);
nand U13599 (N_13599,N_6658,N_7267);
nand U13600 (N_13600,N_11103,N_9043);
and U13601 (N_13601,N_10723,N_12440);
or U13602 (N_13602,N_6910,N_7801);
or U13603 (N_13603,N_11762,N_10475);
and U13604 (N_13604,N_10092,N_9529);
or U13605 (N_13605,N_9058,N_9719);
and U13606 (N_13606,N_11251,N_10710);
xnor U13607 (N_13607,N_11236,N_12160);
nand U13608 (N_13608,N_6367,N_12030);
or U13609 (N_13609,N_6285,N_8396);
or U13610 (N_13610,N_11564,N_8558);
and U13611 (N_13611,N_7050,N_10372);
or U13612 (N_13612,N_7271,N_10962);
xnor U13613 (N_13613,N_6792,N_7850);
nand U13614 (N_13614,N_9007,N_10414);
xor U13615 (N_13615,N_10751,N_10313);
nand U13616 (N_13616,N_11569,N_11393);
and U13617 (N_13617,N_6993,N_7497);
and U13618 (N_13618,N_12174,N_10794);
or U13619 (N_13619,N_8814,N_9699);
nor U13620 (N_13620,N_7895,N_7218);
and U13621 (N_13621,N_7390,N_7136);
nand U13622 (N_13622,N_7495,N_7903);
nand U13623 (N_13623,N_7201,N_9161);
or U13624 (N_13624,N_6698,N_8484);
nor U13625 (N_13625,N_11991,N_6310);
nor U13626 (N_13626,N_6624,N_11115);
or U13627 (N_13627,N_6923,N_11819);
nand U13628 (N_13628,N_11221,N_12093);
xor U13629 (N_13629,N_7880,N_8203);
nor U13630 (N_13630,N_10434,N_7482);
nor U13631 (N_13631,N_8844,N_12303);
or U13632 (N_13632,N_8261,N_12122);
or U13633 (N_13633,N_8931,N_6268);
nand U13634 (N_13634,N_9003,N_6621);
or U13635 (N_13635,N_9218,N_12055);
and U13636 (N_13636,N_7908,N_8744);
nor U13637 (N_13637,N_11237,N_9197);
nand U13638 (N_13638,N_9398,N_11167);
nor U13639 (N_13639,N_9825,N_12296);
or U13640 (N_13640,N_7266,N_7176);
and U13641 (N_13641,N_9428,N_6443);
nand U13642 (N_13642,N_10431,N_11474);
xnor U13643 (N_13643,N_10064,N_8323);
nor U13644 (N_13644,N_11095,N_10482);
nand U13645 (N_13645,N_11071,N_7898);
xor U13646 (N_13646,N_11305,N_6975);
nand U13647 (N_13647,N_10175,N_10255);
nor U13648 (N_13648,N_9210,N_9692);
or U13649 (N_13649,N_9280,N_9682);
nor U13650 (N_13650,N_7660,N_9938);
xnor U13651 (N_13651,N_11999,N_7209);
or U13652 (N_13652,N_8688,N_7275);
or U13653 (N_13653,N_10742,N_7326);
xor U13654 (N_13654,N_6709,N_10694);
xor U13655 (N_13655,N_9324,N_7911);
and U13656 (N_13656,N_9656,N_12311);
nand U13657 (N_13657,N_9487,N_6354);
and U13658 (N_13658,N_7432,N_7453);
nand U13659 (N_13659,N_7325,N_11638);
xor U13660 (N_13660,N_7184,N_11449);
and U13661 (N_13661,N_11455,N_7280);
or U13662 (N_13662,N_9120,N_12477);
nor U13663 (N_13663,N_11789,N_8075);
or U13664 (N_13664,N_12053,N_6362);
and U13665 (N_13665,N_9090,N_7511);
and U13666 (N_13666,N_7306,N_11596);
nor U13667 (N_13667,N_6586,N_10268);
nand U13668 (N_13668,N_6729,N_6425);
xor U13669 (N_13669,N_10600,N_11377);
and U13670 (N_13670,N_6794,N_9789);
or U13671 (N_13671,N_11483,N_10399);
nor U13672 (N_13672,N_7166,N_9469);
and U13673 (N_13673,N_11193,N_9269);
nand U13674 (N_13674,N_9706,N_9972);
nand U13675 (N_13675,N_6776,N_11602);
xor U13676 (N_13676,N_8041,N_9700);
nor U13677 (N_13677,N_7150,N_11533);
or U13678 (N_13678,N_12355,N_8945);
nor U13679 (N_13679,N_6423,N_12333);
nand U13680 (N_13680,N_10704,N_7558);
nor U13681 (N_13681,N_12143,N_7163);
nand U13682 (N_13682,N_10330,N_10544);
nand U13683 (N_13683,N_10200,N_10899);
xor U13684 (N_13684,N_10225,N_6465);
nand U13685 (N_13685,N_9602,N_7664);
nor U13686 (N_13686,N_7755,N_7739);
or U13687 (N_13687,N_8479,N_10888);
nor U13688 (N_13688,N_6454,N_7974);
and U13689 (N_13689,N_9698,N_7401);
nand U13690 (N_13690,N_6690,N_12373);
or U13691 (N_13691,N_9330,N_11486);
and U13692 (N_13692,N_12178,N_10556);
or U13693 (N_13693,N_11828,N_12246);
nor U13694 (N_13694,N_7316,N_6610);
and U13695 (N_13695,N_6864,N_11267);
or U13696 (N_13696,N_6662,N_10568);
nand U13697 (N_13697,N_11241,N_11895);
and U13698 (N_13698,N_10738,N_12475);
nor U13699 (N_13699,N_10686,N_8701);
xnor U13700 (N_13700,N_7416,N_6614);
or U13701 (N_13701,N_7251,N_9651);
or U13702 (N_13702,N_8019,N_11573);
and U13703 (N_13703,N_12247,N_8950);
and U13704 (N_13704,N_11628,N_10798);
or U13705 (N_13705,N_11441,N_10098);
or U13706 (N_13706,N_12127,N_11507);
nand U13707 (N_13707,N_10954,N_11854);
and U13708 (N_13708,N_9072,N_6841);
and U13709 (N_13709,N_7452,N_11179);
nor U13710 (N_13710,N_9776,N_10000);
or U13711 (N_13711,N_11758,N_12337);
xor U13712 (N_13712,N_8496,N_9499);
and U13713 (N_13713,N_10740,N_6599);
or U13714 (N_13714,N_7156,N_12095);
xnor U13715 (N_13715,N_9570,N_6681);
xnor U13716 (N_13716,N_6967,N_8300);
nand U13717 (N_13717,N_11509,N_8921);
or U13718 (N_13718,N_7655,N_11874);
and U13719 (N_13719,N_8042,N_12264);
and U13720 (N_13720,N_7106,N_10188);
xor U13721 (N_13721,N_6338,N_6883);
xnor U13722 (N_13722,N_11457,N_12088);
nand U13723 (N_13723,N_8847,N_12261);
or U13724 (N_13724,N_9149,N_7114);
nand U13725 (N_13725,N_7434,N_8561);
or U13726 (N_13726,N_10034,N_12335);
xor U13727 (N_13727,N_10761,N_7680);
xor U13728 (N_13728,N_9862,N_11084);
or U13729 (N_13729,N_12202,N_10048);
nor U13730 (N_13730,N_10141,N_10265);
xor U13731 (N_13731,N_11383,N_7592);
and U13732 (N_13732,N_7749,N_10154);
nand U13733 (N_13733,N_8643,N_11542);
nand U13734 (N_13734,N_10821,N_11836);
and U13735 (N_13735,N_9480,N_8231);
and U13736 (N_13736,N_9044,N_8421);
nand U13737 (N_13737,N_11308,N_11391);
xnor U13738 (N_13738,N_11253,N_8513);
nand U13739 (N_13739,N_7551,N_9662);
nor U13740 (N_13740,N_7312,N_6760);
nand U13741 (N_13741,N_12466,N_8876);
nand U13742 (N_13742,N_9635,N_10836);
nor U13743 (N_13743,N_10236,N_8011);
or U13744 (N_13744,N_9735,N_10682);
nand U13745 (N_13745,N_12374,N_12367);
nor U13746 (N_13746,N_10582,N_10120);
nand U13747 (N_13747,N_9422,N_8088);
nor U13748 (N_13748,N_8424,N_7391);
or U13749 (N_13749,N_7088,N_9585);
xnor U13750 (N_13750,N_7632,N_6887);
nand U13751 (N_13751,N_6472,N_12254);
nand U13752 (N_13752,N_8175,N_9756);
nor U13753 (N_13753,N_6289,N_7354);
xor U13754 (N_13754,N_9621,N_6651);
or U13755 (N_13755,N_9967,N_11756);
xnor U13756 (N_13756,N_7479,N_6639);
and U13757 (N_13757,N_6655,N_12005);
xor U13758 (N_13758,N_12198,N_11641);
xor U13759 (N_13759,N_7803,N_12150);
and U13760 (N_13760,N_12219,N_12166);
and U13761 (N_13761,N_11618,N_6905);
xor U13762 (N_13762,N_10166,N_10981);
and U13763 (N_13763,N_6805,N_9394);
nor U13764 (N_13764,N_8818,N_12086);
xnor U13765 (N_13765,N_8343,N_12417);
and U13766 (N_13766,N_8587,N_9720);
xnor U13767 (N_13767,N_7819,N_11031);
nor U13768 (N_13768,N_9636,N_11133);
and U13769 (N_13769,N_6979,N_11855);
and U13770 (N_13770,N_10440,N_12215);
nor U13771 (N_13771,N_7285,N_6954);
or U13772 (N_13772,N_10936,N_9500);
xor U13773 (N_13773,N_7687,N_10080);
and U13774 (N_13774,N_9357,N_11772);
or U13775 (N_13775,N_11720,N_10518);
or U13776 (N_13776,N_6476,N_7712);
xor U13777 (N_13777,N_11872,N_8691);
nand U13778 (N_13778,N_7971,N_10167);
xor U13779 (N_13779,N_9793,N_8208);
and U13780 (N_13780,N_10655,N_9981);
nor U13781 (N_13781,N_9668,N_10070);
nor U13782 (N_13782,N_8442,N_6391);
nand U13783 (N_13783,N_11833,N_11173);
and U13784 (N_13784,N_7557,N_9401);
nand U13785 (N_13785,N_11582,N_7058);
nand U13786 (N_13786,N_6857,N_8227);
xor U13787 (N_13787,N_8164,N_9166);
xor U13788 (N_13788,N_8849,N_11302);
xor U13789 (N_13789,N_9008,N_7096);
nor U13790 (N_13790,N_10116,N_7355);
or U13791 (N_13791,N_9289,N_6485);
nor U13792 (N_13792,N_8146,N_6637);
nand U13793 (N_13793,N_11259,N_11471);
xor U13794 (N_13794,N_6407,N_9065);
and U13795 (N_13795,N_9695,N_9235);
nor U13796 (N_13796,N_9400,N_10579);
nor U13797 (N_13797,N_6877,N_8240);
or U13798 (N_13798,N_9051,N_11155);
nand U13799 (N_13799,N_7627,N_9371);
and U13800 (N_13800,N_11610,N_6958);
xor U13801 (N_13801,N_6738,N_6765);
xnor U13802 (N_13802,N_8605,N_10846);
or U13803 (N_13803,N_9431,N_7636);
nand U13804 (N_13804,N_7544,N_9108);
or U13805 (N_13805,N_10195,N_7809);
nor U13806 (N_13806,N_10309,N_8134);
nor U13807 (N_13807,N_8224,N_10184);
nand U13808 (N_13808,N_9535,N_10391);
xnor U13809 (N_13809,N_9618,N_7260);
xnor U13810 (N_13810,N_8885,N_7860);
nor U13811 (N_13811,N_6652,N_11985);
nand U13812 (N_13812,N_7327,N_10788);
or U13813 (N_13813,N_10561,N_7693);
nor U13814 (N_13814,N_8097,N_8221);
xnor U13815 (N_13815,N_8555,N_8387);
nand U13816 (N_13816,N_7628,N_10520);
or U13817 (N_13817,N_8119,N_8362);
xnor U13818 (N_13818,N_12370,N_9923);
nor U13819 (N_13819,N_9963,N_8841);
nor U13820 (N_13820,N_11285,N_6306);
nand U13821 (N_13821,N_6525,N_9405);
or U13822 (N_13822,N_10701,N_11499);
nand U13823 (N_13823,N_8983,N_11121);
or U13824 (N_13824,N_7446,N_10807);
nor U13825 (N_13825,N_9603,N_11376);
and U13826 (N_13826,N_10296,N_10239);
nand U13827 (N_13827,N_9432,N_8780);
xnor U13828 (N_13828,N_11264,N_7338);
xnor U13829 (N_13829,N_10234,N_10934);
nand U13830 (N_13830,N_12300,N_6821);
nand U13831 (N_13831,N_10099,N_11128);
xor U13832 (N_13832,N_8836,N_6871);
nand U13833 (N_13833,N_7884,N_10755);
nor U13834 (N_13834,N_7133,N_10831);
and U13835 (N_13835,N_9619,N_9168);
xnor U13836 (N_13836,N_10847,N_10861);
nor U13837 (N_13837,N_11946,N_7772);
or U13838 (N_13838,N_6351,N_7501);
and U13839 (N_13839,N_9376,N_7849);
or U13840 (N_13840,N_8926,N_10863);
or U13841 (N_13841,N_7000,N_8837);
or U13842 (N_13842,N_10026,N_6286);
and U13843 (N_13843,N_9515,N_9520);
and U13844 (N_13844,N_11901,N_9607);
nor U13845 (N_13845,N_10158,N_10997);
or U13846 (N_13846,N_10204,N_9337);
xor U13847 (N_13847,N_11484,N_6375);
and U13848 (N_13848,N_8953,N_10752);
or U13849 (N_13849,N_9260,N_8717);
nor U13850 (N_13850,N_10430,N_11938);
or U13851 (N_13851,N_11631,N_11841);
and U13852 (N_13852,N_11667,N_11294);
or U13853 (N_13853,N_8689,N_12218);
xnor U13854 (N_13854,N_8851,N_9842);
xor U13855 (N_13855,N_10814,N_9299);
nand U13856 (N_13856,N_10228,N_9936);
and U13857 (N_13857,N_7861,N_6669);
and U13858 (N_13858,N_6487,N_9533);
or U13859 (N_13859,N_8055,N_8051);
and U13860 (N_13860,N_6559,N_8724);
or U13861 (N_13861,N_10489,N_10884);
nor U13862 (N_13862,N_9308,N_10642);
xnor U13863 (N_13863,N_10766,N_9202);
xnor U13864 (N_13864,N_9368,N_10267);
nand U13865 (N_13865,N_10911,N_9693);
and U13866 (N_13866,N_9628,N_8639);
nor U13867 (N_13867,N_10291,N_6336);
xnor U13868 (N_13868,N_6269,N_8004);
or U13869 (N_13869,N_7256,N_6605);
nand U13870 (N_13870,N_7075,N_8280);
and U13871 (N_13871,N_7955,N_12398);
nand U13872 (N_13872,N_11403,N_12157);
or U13873 (N_13873,N_6509,N_6572);
or U13874 (N_13874,N_11183,N_6960);
nor U13875 (N_13875,N_11853,N_6620);
or U13876 (N_13876,N_8358,N_10250);
and U13877 (N_13877,N_11645,N_8989);
xnor U13878 (N_13878,N_11554,N_9177);
nand U13879 (N_13879,N_7027,N_10680);
nand U13880 (N_13880,N_8608,N_9509);
and U13881 (N_13881,N_6836,N_12204);
or U13882 (N_13882,N_9762,N_10851);
or U13883 (N_13883,N_8152,N_6307);
xor U13884 (N_13884,N_9594,N_10499);
or U13885 (N_13885,N_11747,N_11818);
nand U13886 (N_13886,N_8981,N_7451);
and U13887 (N_13887,N_7720,N_9810);
nor U13888 (N_13888,N_11538,N_9797);
or U13889 (N_13889,N_6464,N_7831);
or U13890 (N_13890,N_6386,N_7380);
nand U13891 (N_13891,N_11539,N_10186);
xnor U13892 (N_13892,N_7842,N_6426);
nor U13893 (N_13893,N_6275,N_7762);
nor U13894 (N_13894,N_8161,N_9232);
xnor U13895 (N_13895,N_6549,N_10540);
and U13896 (N_13896,N_10952,N_10842);
nor U13897 (N_13897,N_10949,N_11849);
nand U13898 (N_13898,N_8461,N_9531);
and U13899 (N_13899,N_10539,N_10638);
or U13900 (N_13900,N_10247,N_6263);
or U13901 (N_13901,N_9557,N_8737);
nor U13902 (N_13902,N_10052,N_7015);
xor U13903 (N_13903,N_9680,N_7472);
and U13904 (N_13904,N_8795,N_11695);
or U13905 (N_13905,N_10963,N_10685);
or U13906 (N_13906,N_6713,N_8497);
nor U13907 (N_13907,N_11580,N_9291);
xnor U13908 (N_13908,N_11593,N_8373);
nand U13909 (N_13909,N_11438,N_6937);
nand U13910 (N_13910,N_9941,N_7886);
or U13911 (N_13911,N_8676,N_8411);
and U13912 (N_13912,N_7859,N_8108);
and U13913 (N_13913,N_10852,N_9670);
nand U13914 (N_13914,N_12274,N_11194);
and U13915 (N_13915,N_9132,N_10955);
or U13916 (N_13916,N_11013,N_9418);
nor U13917 (N_13917,N_10601,N_11636);
nand U13918 (N_13918,N_8867,N_9463);
nor U13919 (N_13919,N_7364,N_9663);
xor U13920 (N_13920,N_8415,N_12137);
xnor U13921 (N_13921,N_11292,N_10756);
nand U13922 (N_13922,N_7545,N_10159);
xnor U13923 (N_13923,N_8658,N_7751);
nor U13924 (N_13924,N_8585,N_10534);
or U13925 (N_13925,N_11681,N_7046);
or U13926 (N_13926,N_12291,N_8425);
and U13927 (N_13927,N_7062,N_8173);
and U13928 (N_13928,N_11157,N_12321);
and U13929 (N_13929,N_11506,N_12438);
or U13930 (N_13930,N_12019,N_6377);
nor U13931 (N_13931,N_11549,N_10081);
and U13932 (N_13932,N_7977,N_6292);
or U13933 (N_13933,N_11710,N_6983);
nor U13934 (N_13934,N_8522,N_12224);
nor U13935 (N_13935,N_9925,N_6714);
xnor U13936 (N_13936,N_9391,N_6884);
nor U13937 (N_13937,N_12356,N_9005);
nand U13938 (N_13938,N_8573,N_9848);
nand U13939 (N_13939,N_10809,N_10795);
nand U13940 (N_13940,N_10027,N_9560);
and U13941 (N_13941,N_10538,N_8982);
nand U13942 (N_13942,N_7738,N_8954);
or U13943 (N_13943,N_9980,N_6915);
nand U13944 (N_13944,N_10020,N_8344);
nor U13945 (N_13945,N_9341,N_10588);
xnor U13946 (N_13946,N_7957,N_8142);
nand U13947 (N_13947,N_10975,N_9637);
xnor U13948 (N_13948,N_9467,N_7225);
xnor U13949 (N_13949,N_7093,N_7877);
xnor U13950 (N_13950,N_10687,N_6668);
and U13951 (N_13951,N_10502,N_10927);
nor U13952 (N_13952,N_12163,N_6394);
xnor U13953 (N_13953,N_7976,N_11656);
nor U13954 (N_13954,N_12426,N_9191);
nor U13955 (N_13955,N_9779,N_7725);
or U13956 (N_13956,N_8629,N_9926);
or U13957 (N_13957,N_10257,N_11519);
nor U13958 (N_13958,N_7181,N_10308);
nand U13959 (N_13959,N_7873,N_11318);
or U13960 (N_13960,N_11390,N_8508);
nor U13961 (N_13961,N_10649,N_6429);
or U13962 (N_13962,N_10338,N_10111);
nand U13963 (N_13963,N_8110,N_11764);
and U13964 (N_13964,N_10121,N_10840);
or U13965 (N_13965,N_12395,N_8439);
or U13966 (N_13966,N_9817,N_9711);
nand U13967 (N_13967,N_9804,N_11558);
xnor U13968 (N_13968,N_6843,N_10789);
nand U13969 (N_13969,N_9049,N_10469);
nor U13970 (N_13970,N_8257,N_6628);
nor U13971 (N_13971,N_8250,N_6294);
and U13972 (N_13972,N_7004,N_7676);
nand U13973 (N_13973,N_9613,N_10073);
xor U13974 (N_13974,N_6935,N_12197);
or U13975 (N_13975,N_11666,N_8765);
and U13976 (N_13976,N_7289,N_12452);
nor U13977 (N_13977,N_9525,N_12172);
xor U13978 (N_13978,N_7089,N_6917);
nand U13979 (N_13979,N_8955,N_11931);
and U13980 (N_13980,N_11775,N_9348);
and U13981 (N_13981,N_7883,N_11341);
and U13982 (N_13982,N_9070,N_11090);
nand U13983 (N_13983,N_10615,N_7507);
and U13984 (N_13984,N_8332,N_7988);
xor U13985 (N_13985,N_11058,N_6526);
or U13986 (N_13986,N_7283,N_6468);
nor U13987 (N_13987,N_8528,N_10564);
or U13988 (N_13988,N_10557,N_10078);
and U13989 (N_13989,N_11848,N_12459);
and U13990 (N_13990,N_10486,N_12349);
xnor U13991 (N_13991,N_8195,N_7696);
nand U13992 (N_13992,N_7171,N_11576);
or U13993 (N_13993,N_9250,N_9176);
xnor U13994 (N_13994,N_6648,N_9081);
xnor U13995 (N_13995,N_12111,N_11312);
nand U13996 (N_13996,N_10632,N_7599);
or U13997 (N_13997,N_7255,N_12279);
or U13998 (N_13998,N_10051,N_12415);
or U13999 (N_13999,N_10181,N_8533);
and U14000 (N_14000,N_7060,N_10591);
nand U14001 (N_14001,N_9918,N_9790);
or U14002 (N_14002,N_10984,N_7118);
or U14003 (N_14003,N_10344,N_9961);
and U14004 (N_14004,N_7079,N_6267);
xor U14005 (N_14005,N_7183,N_10014);
nor U14006 (N_14006,N_7706,N_9537);
nand U14007 (N_14007,N_7371,N_9040);
nor U14008 (N_14008,N_12314,N_9430);
or U14009 (N_14009,N_8429,N_6542);
nand U14010 (N_14010,N_10413,N_10784);
xnor U14011 (N_14011,N_10606,N_11680);
or U14012 (N_14012,N_12327,N_10458);
and U14013 (N_14013,N_6399,N_8065);
nand U14014 (N_14014,N_6761,N_10443);
or U14015 (N_14015,N_7800,N_7415);
or U14016 (N_14016,N_11102,N_9841);
or U14017 (N_14017,N_7389,N_12380);
and U14018 (N_14018,N_7059,N_9796);
nor U14019 (N_14019,N_6904,N_10132);
nand U14020 (N_14020,N_9863,N_9015);
nor U14021 (N_14021,N_11753,N_9093);
xor U14022 (N_14022,N_9163,N_9186);
nand U14023 (N_14023,N_10393,N_8084);
nand U14024 (N_14024,N_7835,N_12298);
nand U14025 (N_14025,N_6602,N_7152);
nor U14026 (N_14026,N_12484,N_9544);
nand U14027 (N_14027,N_11091,N_9578);
or U14028 (N_14028,N_11051,N_8583);
and U14029 (N_14029,N_8961,N_6404);
nor U14030 (N_14030,N_12216,N_12140);
or U14031 (N_14031,N_7679,N_10456);
and U14032 (N_14032,N_11277,N_12176);
nor U14033 (N_14033,N_11293,N_7101);
xnor U14034 (N_14034,N_6458,N_7478);
nor U14035 (N_14035,N_7566,N_9320);
and U14036 (N_14036,N_7999,N_9472);
and U14037 (N_14037,N_12054,N_10327);
and U14038 (N_14038,N_11703,N_9461);
xnor U14039 (N_14039,N_8483,N_11629);
xnor U14040 (N_14040,N_7818,N_10999);
xnor U14041 (N_14041,N_8882,N_7288);
nor U14042 (N_14042,N_7193,N_12310);
xor U14043 (N_14043,N_8463,N_11052);
and U14044 (N_14044,N_6523,N_8190);
nand U14045 (N_14045,N_8244,N_6769);
and U14046 (N_14046,N_8116,N_7969);
and U14047 (N_14047,N_7069,N_8347);
nor U14048 (N_14048,N_12012,N_10289);
nand U14049 (N_14049,N_10165,N_8861);
or U14050 (N_14050,N_7115,N_10471);
and U14051 (N_14051,N_9332,N_6762);
nand U14052 (N_14052,N_11935,N_8397);
nand U14053 (N_14053,N_9767,N_8871);
and U14054 (N_14054,N_10919,N_12159);
nor U14055 (N_14055,N_12141,N_7298);
xnor U14056 (N_14056,N_7688,N_9388);
or U14057 (N_14057,N_8326,N_8389);
nand U14058 (N_14058,N_7238,N_7245);
nand U14059 (N_14059,N_9425,N_7736);
nor U14060 (N_14060,N_10140,N_12444);
and U14061 (N_14061,N_8356,N_9362);
nor U14062 (N_14062,N_10916,N_6995);
and U14063 (N_14063,N_6355,N_10124);
or U14064 (N_14064,N_7119,N_8988);
nor U14065 (N_14065,N_10994,N_9060);
and U14066 (N_14066,N_10514,N_8897);
nor U14067 (N_14067,N_9934,N_12313);
xnor U14068 (N_14068,N_11922,N_10832);
nor U14069 (N_14069,N_9880,N_11389);
and U14070 (N_14070,N_12275,N_9243);
xnor U14071 (N_14071,N_6538,N_11339);
nor U14072 (N_14072,N_6701,N_8602);
nor U14073 (N_14073,N_10833,N_7637);
nand U14074 (N_14074,N_11269,N_7966);
and U14075 (N_14075,N_11043,N_9705);
nand U14076 (N_14076,N_8720,N_7454);
nand U14077 (N_14077,N_9999,N_7905);
nor U14078 (N_14078,N_9246,N_6968);
nor U14079 (N_14079,N_12418,N_9436);
nand U14080 (N_14080,N_7648,N_9109);
xnor U14081 (N_14081,N_9517,N_10894);
xor U14082 (N_14082,N_11492,N_9352);
and U14083 (N_14083,N_7492,N_10634);
nand U14084 (N_14084,N_11452,N_8045);
nand U14085 (N_14085,N_7705,N_12363);
nand U14086 (N_14086,N_11543,N_11231);
nor U14087 (N_14087,N_9900,N_11446);
and U14088 (N_14088,N_8710,N_11725);
nand U14089 (N_14089,N_7665,N_10379);
xor U14090 (N_14090,N_12295,N_8580);
nand U14091 (N_14091,N_8531,N_7244);
nor U14092 (N_14092,N_11553,N_9244);
xor U14093 (N_14093,N_10463,N_10692);
and U14094 (N_14094,N_11940,N_10617);
xor U14095 (N_14095,N_8179,N_8297);
and U14096 (N_14096,N_10558,N_9703);
xnor U14097 (N_14097,N_11918,N_7853);
or U14098 (N_14098,N_9447,N_8121);
or U14099 (N_14099,N_10749,N_9947);
or U14100 (N_14100,N_11831,N_7608);
nor U14101 (N_14101,N_9942,N_11664);
nand U14102 (N_14102,N_7509,N_7917);
and U14103 (N_14103,N_7578,N_9450);
nand U14104 (N_14104,N_11118,N_8530);
or U14105 (N_14105,N_9870,N_7045);
or U14106 (N_14106,N_8223,N_6970);
xnor U14107 (N_14107,N_8934,N_7287);
and U14108 (N_14108,N_10363,N_8998);
nor U14109 (N_14109,N_8156,N_9745);
or U14110 (N_14110,N_6583,N_10408);
or U14111 (N_14111,N_8409,N_10422);
nand U14112 (N_14112,N_8977,N_9205);
and U14113 (N_14113,N_11640,N_6912);
nand U14114 (N_14114,N_6507,N_12156);
or U14115 (N_14115,N_8913,N_10827);
and U14116 (N_14116,N_8936,N_8408);
nor U14117 (N_14117,N_7020,N_12301);
and U14118 (N_14118,N_6861,N_11634);
or U14119 (N_14119,N_7723,N_8542);
or U14120 (N_14120,N_7449,N_10565);
and U14121 (N_14121,N_8856,N_9096);
xnor U14122 (N_14122,N_12208,N_9038);
xor U14123 (N_14123,N_10567,N_8739);
nand U14124 (N_14124,N_7257,N_8499);
and U14125 (N_14125,N_11575,N_7979);
or U14126 (N_14126,N_8915,N_11062);
or U14127 (N_14127,N_11057,N_9302);
nand U14128 (N_14128,N_12350,N_8846);
or U14129 (N_14129,N_10892,N_11807);
xnor U14130 (N_14130,N_7593,N_11586);
or U14131 (N_14131,N_11956,N_10702);
or U14132 (N_14132,N_6933,N_7769);
and U14133 (N_14133,N_8680,N_12284);
and U14134 (N_14134,N_11487,N_9495);
and U14135 (N_14135,N_7334,N_7719);
and U14136 (N_14136,N_10571,N_11735);
nand U14137 (N_14137,N_7682,N_8848);
xnor U14138 (N_14138,N_6371,N_8026);
or U14139 (N_14139,N_9737,N_10089);
nand U14140 (N_14140,N_8355,N_10362);
nand U14141 (N_14141,N_7043,N_6531);
nand U14142 (N_14142,N_8753,N_6890);
or U14143 (N_14143,N_8176,N_8975);
xnor U14144 (N_14144,N_9146,N_8209);
xor U14145 (N_14145,N_8437,N_9536);
nand U14146 (N_14146,N_10248,N_11164);
nand U14147 (N_14147,N_7626,N_12408);
and U14148 (N_14148,N_10900,N_6456);
and U14149 (N_14149,N_8899,N_6396);
and U14150 (N_14150,N_11562,N_8896);
or U14151 (N_14151,N_11324,N_7602);
xnor U14152 (N_14152,N_8628,N_7374);
or U14153 (N_14153,N_7754,N_7879);
or U14154 (N_14154,N_11249,N_10198);
or U14155 (N_14155,N_8749,N_10042);
or U14156 (N_14156,N_10445,N_12011);
and U14157 (N_14157,N_10965,N_8559);
and U14158 (N_14158,N_7953,N_9791);
and U14159 (N_14159,N_6804,N_11056);
and U14160 (N_14160,N_12041,N_8684);
or U14161 (N_14161,N_7552,N_8380);
xnor U14162 (N_14162,N_10550,N_7120);
and U14163 (N_14163,N_10759,N_7589);
and U14164 (N_14164,N_8293,N_10912);
nor U14165 (N_14165,N_7393,N_12064);
xnor U14166 (N_14166,N_9145,N_11092);
and U14167 (N_14167,N_12425,N_10290);
xnor U14168 (N_14168,N_7833,N_11006);
xnor U14169 (N_14169,N_8901,N_7299);
xnor U14170 (N_14170,N_9009,N_9884);
and U14171 (N_14171,N_11065,N_11432);
nand U14172 (N_14172,N_11717,N_9995);
or U14173 (N_14173,N_8107,N_10300);
nor U14174 (N_14174,N_6474,N_8596);
nor U14175 (N_14175,N_12280,N_9098);
nor U14176 (N_14176,N_6704,N_12482);
xor U14177 (N_14177,N_10321,N_11774);
or U14178 (N_14178,N_8318,N_12225);
nor U14179 (N_14179,N_8663,N_9047);
or U14180 (N_14180,N_10765,N_10792);
xor U14181 (N_14181,N_11550,N_8912);
nor U14182 (N_14182,N_8023,N_10869);
and U14183 (N_14183,N_9889,N_9690);
and U14184 (N_14184,N_11346,N_11363);
or U14185 (N_14185,N_10035,N_6697);
nand U14186 (N_14186,N_8813,N_11646);
and U14187 (N_14187,N_6374,N_7921);
and U14188 (N_14188,N_9823,N_9503);
xor U14189 (N_14189,N_9414,N_7372);
and U14190 (N_14190,N_6397,N_9086);
xor U14191 (N_14191,N_12242,N_9722);
or U14192 (N_14192,N_10536,N_12359);
nor U14193 (N_14193,N_10873,N_7192);
xor U14194 (N_14194,N_10813,N_10076);
xnor U14195 (N_14195,N_8544,N_8370);
nor U14196 (N_14196,N_7040,N_9914);
xor U14197 (N_14197,N_11959,N_8283);
nor U14198 (N_14198,N_9991,N_10347);
and U14199 (N_14199,N_7887,N_7304);
and U14200 (N_14200,N_9818,N_6881);
nand U14201 (N_14201,N_8543,N_10069);
nand U14202 (N_14202,N_11077,N_8773);
and U14203 (N_14203,N_11522,N_9896);
or U14204 (N_14204,N_7826,N_12325);
and U14205 (N_14205,N_9192,N_8287);
and U14206 (N_14206,N_9876,N_12220);
xor U14207 (N_14207,N_9415,N_11101);
and U14208 (N_14208,N_8535,N_7647);
nor U14209 (N_14209,N_11559,N_8143);
or U14210 (N_14210,N_9519,N_9107);
xnor U14211 (N_14211,N_10340,N_7869);
nand U14212 (N_14212,N_11708,N_11214);
and U14213 (N_14213,N_9215,N_10150);
nand U14214 (N_14214,N_10804,N_11612);
nor U14215 (N_14215,N_11127,N_8670);
nand U14216 (N_14216,N_6571,N_11800);
or U14217 (N_14217,N_8995,N_11994);
or U14218 (N_14218,N_7576,N_10664);
nor U14219 (N_14219,N_6534,N_8631);
or U14220 (N_14220,N_8708,N_8404);
nor U14221 (N_14221,N_8037,N_9312);
nand U14222 (N_14222,N_9333,N_11504);
or U14223 (N_14223,N_8551,N_10566);
or U14224 (N_14224,N_11428,N_9882);
nand U14225 (N_14225,N_11174,N_8782);
and U14226 (N_14226,N_7605,N_10001);
xor U14227 (N_14227,N_7349,N_7841);
nor U14228 (N_14228,N_7686,N_9420);
and U14229 (N_14229,N_10815,N_7487);
nor U14230 (N_14230,N_9642,N_7595);
nor U14231 (N_14231,N_10805,N_9307);
or U14232 (N_14232,N_6569,N_7653);
nand U14233 (N_14233,N_8238,N_11810);
nand U14234 (N_14234,N_7204,N_10219);
or U14235 (N_14235,N_6759,N_10849);
or U14236 (N_14236,N_8192,N_11838);
nand U14237 (N_14237,N_11232,N_12328);
or U14238 (N_14238,N_9429,N_7572);
nor U14239 (N_14239,N_8038,N_12481);
xor U14240 (N_14240,N_6866,N_10496);
and U14241 (N_14241,N_9380,N_10174);
nor U14242 (N_14242,N_11729,N_9915);
xor U14243 (N_14243,N_10830,N_9028);
nor U14244 (N_14244,N_7147,N_12405);
or U14245 (N_14245,N_7611,N_8986);
nand U14246 (N_14246,N_8567,N_12097);
nand U14247 (N_14247,N_7278,N_9847);
or U14248 (N_14248,N_8878,N_9750);
or U14249 (N_14249,N_10029,N_10388);
nand U14250 (N_14250,N_9872,N_10390);
nand U14251 (N_14251,N_11788,N_8994);
or U14252 (N_14252,N_6469,N_12107);
xnor U14253 (N_14253,N_6706,N_6252);
xnor U14254 (N_14254,N_9657,N_10695);
or U14255 (N_14255,N_10117,N_9650);
or U14256 (N_14256,N_7771,N_7488);
xor U14257 (N_14257,N_8210,N_6718);
nor U14258 (N_14258,N_11625,N_11080);
nand U14259 (N_14259,N_11443,N_11925);
nand U14260 (N_14260,N_11906,N_10689);
nand U14261 (N_14261,N_10745,N_8967);
or U14262 (N_14262,N_7904,N_12277);
nand U14263 (N_14263,N_8394,N_6430);
xnor U14264 (N_14264,N_6457,N_10675);
xnor U14265 (N_14265,N_12453,N_11401);
and U14266 (N_14266,N_6711,N_11094);
and U14267 (N_14267,N_9406,N_11784);
and U14268 (N_14268,N_8859,N_9857);
nand U14269 (N_14269,N_8365,N_7577);
and U14270 (N_14270,N_10729,N_11992);
nand U14271 (N_14271,N_9562,N_11515);
xnor U14272 (N_14272,N_10683,N_11523);
xnor U14273 (N_14273,N_10707,N_10678);
or U14274 (N_14274,N_10971,N_11284);
nor U14275 (N_14275,N_6902,N_9501);
or U14276 (N_14276,N_6483,N_9715);
or U14277 (N_14277,N_6557,N_10339);
xnor U14278 (N_14278,N_11754,N_11537);
xnor U14279 (N_14279,N_8071,N_7967);
or U14280 (N_14280,N_6870,N_12494);
xnor U14281 (N_14281,N_7033,N_11763);
and U14282 (N_14282,N_7219,N_10455);
and U14283 (N_14283,N_10493,N_9723);
nand U14284 (N_14284,N_11099,N_11182);
and U14285 (N_14285,N_9826,N_10677);
and U14286 (N_14286,N_7321,N_8545);
and U14287 (N_14287,N_10754,N_11979);
nor U14288 (N_14288,N_11909,N_11755);
nand U14289 (N_14289,N_11672,N_8086);
nor U14290 (N_14290,N_11074,N_8581);
nor U14291 (N_14291,N_12471,N_10303);
nand U14292 (N_14292,N_7274,N_8536);
xnor U14293 (N_14293,N_8582,N_6911);
or U14294 (N_14294,N_8704,N_8514);
and U14295 (N_14295,N_7444,N_7162);
nand U14296 (N_14296,N_12027,N_9574);
xor U14297 (N_14297,N_12000,N_6372);
xor U14298 (N_14298,N_9106,N_7591);
xor U14299 (N_14299,N_11749,N_11510);
nand U14300 (N_14300,N_11620,N_6482);
xor U14301 (N_14301,N_9247,N_7986);
and U14302 (N_14302,N_6591,N_10404);
nand U14303 (N_14303,N_7167,N_10025);
or U14304 (N_14304,N_7533,N_8735);
or U14305 (N_14305,N_10405,N_6432);
xor U14306 (N_14306,N_11851,N_11015);
or U14307 (N_14307,N_12312,N_10316);
and U14308 (N_14308,N_7750,N_6680);
and U14309 (N_14309,N_10607,N_12146);
or U14310 (N_14310,N_7532,N_12181);
xor U14311 (N_14311,N_8001,N_8947);
or U14312 (N_14312,N_8564,N_8306);
nor U14313 (N_14313,N_10008,N_11742);
or U14314 (N_14314,N_6530,N_7821);
xor U14315 (N_14315,N_11143,N_7674);
nor U14316 (N_14316,N_8838,N_7692);
or U14317 (N_14317,N_10128,N_11796);
nand U14318 (N_14318,N_11548,N_12424);
nand U14319 (N_14319,N_9101,N_9904);
or U14320 (N_14320,N_11597,N_9929);
nor U14321 (N_14321,N_7561,N_10418);
nand U14322 (N_14322,N_9057,N_8711);
xnor U14323 (N_14323,N_12400,N_8237);
nand U14324 (N_14324,N_9257,N_11222);
xor U14325 (N_14325,N_12014,N_7485);
and U14326 (N_14326,N_8307,N_11400);
and U14327 (N_14327,N_6528,N_10501);
xnor U14328 (N_14328,N_6393,N_8834);
nor U14329 (N_14329,N_6466,N_6682);
and U14330 (N_14330,N_8350,N_8309);
nor U14331 (N_14331,N_8755,N_11488);
or U14332 (N_14332,N_6914,N_6303);
xor U14333 (N_14333,N_12152,N_8903);
nor U14334 (N_14334,N_7562,N_12267);
or U14335 (N_14335,N_9956,N_11529);
xnor U14336 (N_14336,N_9206,N_12126);
nor U14337 (N_14337,N_10488,N_9396);
and U14338 (N_14338,N_9969,N_7892);
nor U14339 (N_14339,N_6703,N_10160);
nor U14340 (N_14340,N_7560,N_6846);
xor U14341 (N_14341,N_9440,N_10768);
xor U14342 (N_14342,N_7242,N_8827);
and U14343 (N_14343,N_7402,N_6820);
xnor U14344 (N_14344,N_11139,N_7612);
nor U14345 (N_14345,N_10939,N_10907);
and U14346 (N_14346,N_6347,N_10032);
nor U14347 (N_14347,N_8925,N_8052);
xnor U14348 (N_14348,N_6693,N_11804);
and U14349 (N_14349,N_11693,N_8194);
and U14350 (N_14350,N_8337,N_10920);
or U14351 (N_14351,N_11847,N_7090);
and U14352 (N_14352,N_7347,N_7782);
xor U14353 (N_14353,N_7649,N_10618);
nor U14354 (N_14354,N_10387,N_11933);
nand U14355 (N_14355,N_7013,N_10420);
or U14356 (N_14356,N_11434,N_9885);
xnor U14357 (N_14357,N_11008,N_8868);
xor U14358 (N_14358,N_12384,N_6876);
nand U14359 (N_14359,N_9290,N_10943);
and U14360 (N_14360,N_9134,N_12248);
xor U14361 (N_14361,N_10142,N_12334);
and U14362 (N_14362,N_8166,N_11736);
or U14363 (N_14363,N_9470,N_9979);
nor U14364 (N_14364,N_8186,N_8201);
nand U14365 (N_14365,N_8843,N_9953);
xor U14366 (N_14366,N_10381,N_10636);
nor U14367 (N_14367,N_8464,N_7343);
and U14368 (N_14368,N_8864,N_8980);
nand U14369 (N_14369,N_7345,N_6422);
nand U14370 (N_14370,N_10286,N_8825);
or U14371 (N_14371,N_11730,N_10196);
and U14372 (N_14372,N_12094,N_8576);
or U14373 (N_14373,N_9932,N_10989);
xor U14374 (N_14374,N_8178,N_6251);
nor U14375 (N_14375,N_10864,N_8661);
or U14376 (N_14376,N_7529,N_11595);
nor U14377 (N_14377,N_8731,N_7519);
xor U14378 (N_14378,N_8423,N_7185);
or U14379 (N_14379,N_10504,N_7703);
nand U14380 (N_14380,N_12044,N_6897);
nand U14381 (N_14381,N_10122,N_10922);
nor U14382 (N_14382,N_8135,N_10679);
nand U14383 (N_14383,N_9749,N_8625);
nand U14384 (N_14384,N_10672,N_9213);
or U14385 (N_14385,N_6364,N_11948);
nor U14386 (N_14386,N_8111,N_8339);
or U14387 (N_14387,N_10876,N_10210);
and U14388 (N_14388,N_8379,N_11557);
or U14389 (N_14389,N_6328,N_6365);
xor U14390 (N_14390,N_7901,N_10651);
nand U14391 (N_14391,N_11314,N_10415);
and U14392 (N_14392,N_9147,N_7010);
xnor U14393 (N_14393,N_11769,N_12430);
and U14394 (N_14394,N_8667,N_9881);
nand U14395 (N_14395,N_8467,N_12315);
nand U14396 (N_14396,N_7554,N_10084);
nand U14397 (N_14397,N_7315,N_10447);
xnor U14398 (N_14398,N_11511,N_12105);
nor U14399 (N_14399,N_9755,N_11502);
and U14400 (N_14400,N_10825,N_10650);
nor U14401 (N_14401,N_9412,N_8518);
nand U14402 (N_14402,N_10310,N_8532);
and U14403 (N_14403,N_8020,N_11020);
or U14404 (N_14404,N_10269,N_11884);
xnor U14405 (N_14405,N_11290,N_6676);
xor U14406 (N_14406,N_7103,N_8877);
nor U14407 (N_14407,N_7505,N_12076);
nor U14408 (N_14408,N_11768,N_10942);
nor U14409 (N_14409,N_8475,N_6830);
and U14410 (N_14410,N_9061,N_9159);
nand U14411 (N_14411,N_8778,N_6475);
nor U14412 (N_14412,N_10532,N_10375);
and U14413 (N_14413,N_8784,N_9633);
xnor U14414 (N_14414,N_11206,N_7188);
nor U14415 (N_14415,N_7044,N_6316);
nand U14416 (N_14416,N_7284,N_6541);
and U14417 (N_14417,N_12467,N_10879);
and U14418 (N_14418,N_7430,N_8368);
xnor U14419 (N_14419,N_6582,N_11781);
and U14420 (N_14420,N_11965,N_10666);
xor U14421 (N_14421,N_6616,N_7042);
or U14422 (N_14422,N_9021,N_12155);
nand U14423 (N_14423,N_6749,N_9037);
xor U14424 (N_14424,N_10394,N_9508);
xor U14425 (N_14425,N_9175,N_11830);
nor U14426 (N_14426,N_10351,N_10843);
or U14427 (N_14427,N_8292,N_6849);
xor U14428 (N_14428,N_9451,N_11964);
nand U14429 (N_14429,N_10599,N_12362);
nand U14430 (N_14430,N_7847,N_6828);
xnor U14431 (N_14431,N_6369,N_7186);
or U14432 (N_14432,N_9761,N_11323);
nand U14433 (N_14433,N_10012,N_11466);
nand U14434 (N_14434,N_7305,N_12239);
nor U14435 (N_14435,N_11165,N_8500);
or U14436 (N_14436,N_9438,N_9812);
nand U14437 (N_14437,N_8833,N_11556);
nor U14438 (N_14438,N_6280,N_10044);
nor U14439 (N_14439,N_9566,N_7708);
xnor U14440 (N_14440,N_9768,N_12017);
nand U14441 (N_14441,N_12427,N_9066);
nand U14442 (N_14442,N_8799,N_7768);
and U14443 (N_14443,N_11678,N_11150);
xor U14444 (N_14444,N_11477,N_9251);
xnor U14445 (N_14445,N_9511,N_11295);
or U14446 (N_14446,N_7356,N_7893);
xor U14447 (N_14447,N_10274,N_10964);
and U14448 (N_14448,N_8599,N_10461);
xor U14449 (N_14449,N_6852,N_9083);
nand U14450 (N_14450,N_8783,N_9801);
or U14451 (N_14451,N_11180,N_7671);
or U14452 (N_14452,N_11010,N_6982);
xor U14453 (N_14453,N_9551,N_6431);
nor U14454 (N_14454,N_8874,N_7474);
nand U14455 (N_14455,N_8005,N_9171);
nand U14456 (N_14456,N_12317,N_9222);
and U14457 (N_14457,N_11362,N_7302);
and U14458 (N_14458,N_10480,N_9897);
nand U14459 (N_14459,N_11896,N_6477);
nand U14460 (N_14460,N_8125,N_11561);
or U14461 (N_14461,N_8984,N_11450);
nand U14462 (N_14462,N_10010,N_12270);
xnor U14463 (N_14463,N_9053,N_8942);
xnor U14464 (N_14464,N_11957,N_11001);
or U14465 (N_14465,N_10258,N_8262);
nand U14466 (N_14466,N_12136,N_9748);
xor U14467 (N_14467,N_11067,N_7677);
nor U14468 (N_14468,N_11445,N_9462);
nand U14469 (N_14469,N_11387,N_6739);
or U14470 (N_14470,N_12391,N_8604);
nor U14471 (N_14471,N_8275,N_11032);
nand U14472 (N_14472,N_11815,N_11453);
or U14473 (N_14473,N_6486,N_9122);
and U14474 (N_14474,N_7379,N_11777);
or U14475 (N_14475,N_9255,N_11119);
nor U14476 (N_14476,N_10261,N_10576);
and U14477 (N_14477,N_6654,N_8008);
nor U14478 (N_14478,N_6784,N_8096);
and U14479 (N_14479,N_9479,N_7177);
and U14480 (N_14480,N_7132,N_8622);
nand U14481 (N_14481,N_12147,N_11287);
xnor U14482 (N_14482,N_10782,N_7269);
or U14483 (N_14483,N_7989,N_7328);
nor U14484 (N_14484,N_6408,N_11137);
nor U14485 (N_14485,N_10487,N_11570);
xnor U14486 (N_14486,N_6780,N_8633);
or U14487 (N_14487,N_9921,N_10545);
nor U14488 (N_14488,N_9974,N_9669);
xnor U14489 (N_14489,N_9493,N_8308);
or U14490 (N_14490,N_8969,N_6406);
nor U14491 (N_14491,N_7189,N_6675);
nor U14492 (N_14492,N_11655,N_9248);
nand U14493 (N_14493,N_8310,N_10416);
and U14494 (N_14494,N_11718,N_9456);
nand U14495 (N_14495,N_9331,N_9626);
or U14496 (N_14496,N_9445,N_12192);
or U14497 (N_14497,N_6633,N_12297);
and U14498 (N_14498,N_11919,N_7704);
nand U14499 (N_14499,N_11359,N_7440);
xnor U14500 (N_14500,N_11047,N_12420);
or U14501 (N_14501,N_11388,N_10613);
and U14502 (N_14502,N_12316,N_8313);
xor U14503 (N_14503,N_10543,N_10905);
or U14504 (N_14504,N_10074,N_11343);
or U14505 (N_14505,N_10881,N_9010);
and U14506 (N_14506,N_7865,N_11192);
and U14507 (N_14507,N_8346,N_10377);
xnor U14508 (N_14508,N_6716,N_8656);
nand U14509 (N_14509,N_7798,N_11757);
nor U14510 (N_14510,N_8898,N_8517);
and U14511 (N_14511,N_12010,N_6908);
or U14512 (N_14512,N_10796,N_7812);
or U14513 (N_14513,N_6962,N_7938);
nor U14514 (N_14514,N_12308,N_6348);
or U14515 (N_14515,N_7874,N_6495);
nor U14516 (N_14516,N_6357,N_11662);
nand U14517 (N_14517,N_11018,N_11532);
and U14518 (N_14518,N_12283,N_8348);
nor U14519 (N_14519,N_10623,N_7614);
nand U14520 (N_14520,N_10354,N_6344);
nand U14521 (N_14521,N_12121,N_9356);
nand U14522 (N_14522,N_10699,N_9993);
or U14523 (N_14523,N_8416,N_9660);
nand U14524 (N_14524,N_9165,N_12040);
or U14525 (N_14525,N_8412,N_8997);
nand U14526 (N_14526,N_6608,N_8845);
xor U14527 (N_14527,N_10739,N_11799);
and U14528 (N_14528,N_10105,N_7396);
nand U14529 (N_14529,N_9231,N_11248);
nand U14530 (N_14530,N_12173,N_11822);
nor U14531 (N_14531,N_7925,N_8798);
and U14532 (N_14532,N_9465,N_8316);
or U14533 (N_14533,N_8840,N_10238);
xor U14534 (N_14534,N_11927,N_11934);
nand U14535 (N_14535,N_8157,N_10191);
or U14536 (N_14536,N_9962,N_8400);
and U14537 (N_14537,N_10441,N_8002);
xor U14538 (N_14538,N_7228,N_9387);
nor U14539 (N_14539,N_8258,N_9226);
xnor U14540 (N_14540,N_11696,N_6282);
nor U14541 (N_14541,N_9593,N_7250);
and U14542 (N_14542,N_11169,N_9724);
nand U14543 (N_14543,N_12123,N_10903);
xnor U14544 (N_14544,N_11887,N_10810);
xnor U14545 (N_14545,N_7948,N_10624);
xnor U14546 (N_14546,N_11514,N_11877);
and U14547 (N_14547,N_7254,N_9199);
nand U14548 (N_14548,N_12336,N_8325);
or U14549 (N_14549,N_8296,N_6500);
and U14550 (N_14550,N_12472,N_7503);
and U14551 (N_14551,N_8085,N_8320);
or U14552 (N_14552,N_8682,N_8028);
and U14553 (N_14553,N_10009,N_6556);
nand U14554 (N_14554,N_12392,N_10570);
or U14555 (N_14555,N_11042,N_6839);
xnor U14556 (N_14556,N_9883,N_8673);
and U14557 (N_14557,N_9978,N_8476);
xnor U14558 (N_14558,N_9910,N_12120);
nand U14559 (N_14559,N_9187,N_7956);
nand U14560 (N_14560,N_8640,N_7727);
and U14561 (N_14561,N_7233,N_11865);
or U14562 (N_14562,N_11404,N_7890);
nor U14563 (N_14563,N_11857,N_12117);
or U14564 (N_14564,N_9153,N_11354);
and U14565 (N_14565,N_8970,N_8174);
nor U14566 (N_14566,N_9629,N_11260);
nand U14567 (N_14567,N_11350,N_10516);
nor U14568 (N_14568,N_7586,N_9911);
nor U14569 (N_14569,N_11824,N_6859);
xnor U14570 (N_14570,N_11732,N_8126);
or U14571 (N_14571,N_6850,N_9807);
or U14572 (N_14572,N_8137,N_8357);
xnor U14573 (N_14573,N_11845,N_7934);
xnor U14574 (N_14574,N_8539,N_10173);
nor U14575 (N_14575,N_9492,N_7024);
xnor U14576 (N_14576,N_10306,N_11146);
and U14577 (N_14577,N_9327,N_6724);
and U14578 (N_14578,N_11337,N_12085);
nor U14579 (N_14579,N_11298,N_7683);
and U14580 (N_14580,N_7017,N_9777);
and U14581 (N_14581,N_10509,N_6254);
and U14582 (N_14582,N_9119,N_10177);
or U14583 (N_14583,N_6891,N_12456);
nand U14584 (N_14584,N_7731,N_6382);
or U14585 (N_14585,N_11827,N_12496);
nand U14586 (N_14586,N_11986,N_11475);
xnor U14587 (N_14587,N_7962,N_6598);
or U14588 (N_14588,N_8003,N_6380);
or U14589 (N_14589,N_10277,N_7932);
and U14590 (N_14590,N_6853,N_7834);
xor U14591 (N_14591,N_6906,N_7032);
nor U14592 (N_14592,N_8315,N_7829);
nand U14593 (N_14593,N_7061,N_12077);
nor U14594 (N_14594,N_7598,N_11737);
or U14595 (N_14595,N_11863,N_9581);
or U14596 (N_14596,N_9136,N_6816);
nand U14597 (N_14597,N_12448,N_8624);
xor U14598 (N_14598,N_7307,N_8386);
nand U14599 (N_14599,N_11498,N_10595);
xor U14600 (N_14600,N_9652,N_10546);
xnor U14601 (N_14601,N_8985,N_8113);
nand U14602 (N_14602,N_8012,N_10450);
xnor U14603 (N_14603,N_9561,N_8105);
nand U14604 (N_14604,N_7641,N_11097);
nor U14605 (N_14605,N_8444,N_11535);
and U14606 (N_14606,N_9367,N_8651);
or U14607 (N_14607,N_7965,N_8230);
xnor U14608 (N_14608,N_8590,N_7055);
and U14609 (N_14609,N_7419,N_9946);
or U14610 (N_14610,N_12138,N_10037);
or U14611 (N_14611,N_8074,N_11604);
or U14612 (N_14612,N_11571,N_8537);
and U14613 (N_14613,N_11930,N_8687);
xnor U14614 (N_14614,N_9256,N_10733);
xor U14615 (N_14615,N_7907,N_9830);
or U14616 (N_14616,N_10222,N_9927);
or U14617 (N_14617,N_11371,N_9378);
or U14618 (N_14618,N_8211,N_7041);
nor U14619 (N_14619,N_7381,N_7698);
or U14620 (N_14620,N_8489,N_11219);
nand U14621 (N_14621,N_9666,N_10331);
and U14622 (N_14622,N_9137,N_9620);
or U14623 (N_14623,N_11607,N_10696);
nand U14624 (N_14624,N_7142,N_7130);
nand U14625 (N_14625,N_7899,N_7909);
or U14626 (N_14626,N_6529,N_12462);
or U14627 (N_14627,N_9417,N_11560);
xnor U14628 (N_14628,N_9853,N_9746);
or U14629 (N_14629,N_8642,N_10705);
or U14630 (N_14630,N_8282,N_9141);
xnor U14631 (N_14631,N_11372,N_8732);
nor U14632 (N_14632,N_9477,N_7862);
or U14633 (N_14633,N_11540,N_9630);
nor U14634 (N_14634,N_11829,N_7113);
nand U14635 (N_14635,N_8448,N_10944);
nor U14636 (N_14636,N_9020,N_8572);
or U14637 (N_14637,N_10134,N_6873);
and U14638 (N_14638,N_8529,N_9221);
xor U14639 (N_14639,N_7774,N_11809);
and U14640 (N_14640,N_7968,N_10930);
or U14641 (N_14641,N_10530,N_10360);
and U14642 (N_14642,N_8417,N_9919);
or U14643 (N_14643,N_9476,N_9488);
and U14644 (N_14644,N_9739,N_11244);
nor U14645 (N_14645,N_8482,N_9006);
or U14646 (N_14646,N_7258,N_7542);
or U14647 (N_14647,N_12031,N_11113);
and U14648 (N_14648,N_11856,N_7300);
nand U14649 (N_14649,N_10039,N_7565);
and U14650 (N_14650,N_7517,N_9579);
nor U14651 (N_14651,N_10978,N_11839);
nor U14652 (N_14652,N_7716,N_10119);
xnor U14653 (N_14653,N_9640,N_11707);
xnor U14654 (N_14654,N_10870,N_8198);
and U14655 (N_14655,N_8695,N_11108);
xor U14656 (N_14656,N_10030,N_7360);
and U14657 (N_14657,N_8233,N_12324);
or U14658 (N_14658,N_9024,N_8853);
xor U14659 (N_14659,N_9097,N_11723);
and U14660 (N_14660,N_10893,N_8101);
or U14661 (N_14661,N_7790,N_7625);
nor U14662 (N_14662,N_9572,N_9264);
and U14663 (N_14663,N_9384,N_8715);
or U14664 (N_14664,N_9667,N_7689);
nand U14665 (N_14665,N_7261,N_9427);
nor U14666 (N_14666,N_7742,N_7804);
nor U14667 (N_14667,N_12469,N_8199);
and U14668 (N_14668,N_12454,N_9838);
xor U14669 (N_14669,N_11883,N_9524);
xnor U14670 (N_14670,N_7428,N_9464);
nand U14671 (N_14671,N_10180,N_12063);
nor U14672 (N_14672,N_7281,N_9856);
or U14673 (N_14673,N_10216,N_7077);
nor U14674 (N_14674,N_9645,N_7807);
and U14675 (N_14675,N_9100,N_9824);
or U14676 (N_14676,N_12449,N_12480);
or U14677 (N_14677,N_6390,N_11960);
nor U14678 (N_14678,N_8359,N_9403);
xor U14679 (N_14679,N_6930,N_12034);
nor U14680 (N_14680,N_7506,N_10605);
or U14681 (N_14681,N_9386,N_9548);
nand U14682 (N_14682,N_7787,N_11098);
or U14683 (N_14683,N_9783,N_7943);
nor U14684 (N_14684,N_12075,N_8187);
and U14685 (N_14685,N_11235,N_6710);
nor U14686 (N_14686,N_8754,N_7638);
nor U14687 (N_14687,N_8153,N_7778);
nand U14688 (N_14688,N_8672,N_12318);
nand U14689 (N_14689,N_11130,N_12237);
or U14690 (N_14690,N_8031,N_8937);
nand U14691 (N_14691,N_6964,N_12177);
or U14692 (N_14692,N_8707,N_10298);
nor U14693 (N_14693,N_7828,N_11773);
and U14694 (N_14694,N_8027,N_8858);
nor U14695 (N_14695,N_11587,N_12074);
xor U14696 (N_14696,N_11803,N_9087);
nand U14697 (N_14697,N_8331,N_8563);
nand U14698 (N_14698,N_11908,N_11203);
nand U14699 (N_14699,N_7553,N_9014);
xor U14700 (N_14700,N_12222,N_12461);
nor U14701 (N_14701,N_11223,N_10728);
nand U14702 (N_14702,N_8243,N_7117);
xnor U14703 (N_14703,N_12499,N_8565);
or U14704 (N_14704,N_8797,N_11191);
nand U14705 (N_14705,N_8057,N_9583);
nand U14706 (N_14706,N_12404,N_7639);
nor U14707 (N_14707,N_7313,N_10775);
xnor U14708 (N_14708,N_9241,N_11617);
xor U14709 (N_14709,N_6501,N_9085);
nor U14710 (N_14710,N_10096,N_11786);
xnor U14711 (N_14711,N_11878,N_7229);
nor U14712 (N_14712,N_9298,N_6451);
nand U14713 (N_14713,N_9011,N_9975);
or U14714 (N_14714,N_8611,N_9591);
and U14715 (N_14715,N_12024,N_8498);
nand U14716 (N_14716,N_7824,N_7190);
and U14717 (N_14717,N_8546,N_11531);
xnor U14718 (N_14718,N_6504,N_7526);
nor U14719 (N_14719,N_7292,N_9212);
nor U14720 (N_14720,N_11258,N_11114);
xnor U14721 (N_14721,N_6455,N_12272);
xor U14722 (N_14722,N_7213,N_9183);
xnor U14723 (N_14723,N_7165,N_9707);
nor U14724 (N_14724,N_11009,N_9443);
nand U14725 (N_14725,N_12045,N_11037);
or U14726 (N_14726,N_7016,N_8873);
xnor U14727 (N_14727,N_8024,N_7690);
xnor U14728 (N_14728,N_10152,N_8973);
nand U14729 (N_14729,N_12341,N_8093);
or U14730 (N_14730,N_7107,N_7575);
or U14731 (N_14731,N_8406,N_10428);
xor U14732 (N_14732,N_12047,N_8087);
nand U14733 (N_14733,N_6686,N_7984);
and U14734 (N_14734,N_11914,N_12052);
xnor U14735 (N_14735,N_10628,N_7500);
nor U14736 (N_14736,N_6433,N_9321);
nand U14737 (N_14737,N_10519,N_7375);
nor U14738 (N_14738,N_9710,N_6966);
xnor U14739 (N_14739,N_11682,N_9366);
and U14740 (N_14740,N_8214,N_7926);
nor U14741 (N_14741,N_10659,N_7775);
nor U14742 (N_14742,N_6947,N_7802);
nor U14743 (N_14743,N_11647,N_12365);
nor U14744 (N_14744,N_9372,N_7891);
nand U14745 (N_14745,N_9799,N_6894);
nand U14746 (N_14746,N_8927,N_6629);
xor U14747 (N_14747,N_7843,N_6537);
nand U14748 (N_14748,N_7448,N_10951);
xor U14749 (N_14749,N_7007,N_7112);
and U14750 (N_14750,N_11288,N_12348);
xnor U14751 (N_14751,N_9673,N_10208);
nand U14752 (N_14752,N_11125,N_12435);
and U14753 (N_14753,N_11106,N_11911);
nand U14754 (N_14754,N_11328,N_9922);
nand U14755 (N_14755,N_7368,N_10762);
and U14756 (N_14756,N_10797,N_9676);
nand U14757 (N_14757,N_8035,N_10346);
nand U14758 (N_14758,N_10727,N_9353);
xnor U14759 (N_14759,N_6398,N_8880);
and U14760 (N_14760,N_10444,N_8191);
or U14761 (N_14761,N_10164,N_9997);
nand U14762 (N_14762,N_9118,N_6452);
xor U14763 (N_14763,N_10337,N_7383);
nor U14764 (N_14764,N_8197,N_6575);
nor U14765 (N_14765,N_10878,N_11987);
and U14766 (N_14766,N_12082,N_9522);
or U14767 (N_14767,N_10386,N_11422);
xor U14768 (N_14768,N_12464,N_9820);
or U14769 (N_14769,N_6601,N_10022);
nand U14770 (N_14770,N_11360,N_12465);
and U14771 (N_14771,N_8390,N_7070);
and U14772 (N_14772,N_8810,N_11858);
nor U14773 (N_14773,N_9763,N_9379);
nand U14774 (N_14774,N_6732,N_8816);
nand U14775 (N_14775,N_10819,N_7436);
nand U14776 (N_14776,N_10371,N_9329);
or U14777 (N_14777,N_10937,N_10396);
and U14778 (N_14778,N_8979,N_8114);
xor U14779 (N_14779,N_7691,N_9778);
xnor U14780 (N_14780,N_7191,N_8763);
and U14781 (N_14781,N_6837,N_9194);
and U14782 (N_14782,N_7714,N_6274);
nand U14783 (N_14783,N_10511,N_10365);
xor U14784 (N_14784,N_6684,N_11212);
and U14785 (N_14785,N_10609,N_7745);
nand U14786 (N_14786,N_9410,N_11060);
xor U14787 (N_14787,N_11882,N_11480);
and U14788 (N_14788,N_7580,N_12068);
and U14789 (N_14789,N_12457,N_9563);
xor U14790 (N_14790,N_7293,N_11798);
or U14791 (N_14791,N_10793,N_6921);
or U14792 (N_14792,N_11365,N_10806);
xor U14793 (N_14793,N_8216,N_11665);
or U14794 (N_14794,N_7670,N_10610);
nand U14795 (N_14795,N_11479,N_6783);
xor U14796 (N_14796,N_10417,N_8112);
nor U14797 (N_14797,N_10669,N_12101);
nand U14798 (N_14798,N_9632,N_8589);
or U14799 (N_14799,N_11653,N_7081);
or U14800 (N_14800,N_10735,N_7034);
or U14801 (N_14801,N_9592,N_6969);
nand U14802 (N_14802,N_9358,N_10284);
or U14803 (N_14803,N_7319,N_10028);
nand U14804 (N_14804,N_11600,N_8987);
nand U14805 (N_14805,N_6896,N_7996);
nor U14806 (N_14806,N_9077,N_11247);
and U14807 (N_14807,N_9516,N_9110);
or U14808 (N_14808,N_7848,N_7407);
nand U14809 (N_14809,N_7155,N_10192);
nand U14810 (N_14810,N_10658,N_7386);
xor U14811 (N_14811,N_7268,N_8709);
nor U14812 (N_14812,N_10945,N_10059);
or U14813 (N_14813,N_12190,N_9130);
nor U14814 (N_14814,N_7657,N_8817);
and U14815 (N_14815,N_10823,N_8703);
nor U14816 (N_14816,N_10890,N_11792);
xnor U14817 (N_14817,N_6262,N_8978);
nor U14818 (N_14818,N_6699,N_9318);
or U14819 (N_14819,N_7980,N_8686);
nand U14820 (N_14820,N_8924,N_6833);
and U14821 (N_14821,N_6677,N_10988);
nand U14822 (N_14822,N_10886,N_9481);
and U14823 (N_14823,N_8481,N_11353);
xnor U14824 (N_14824,N_11116,N_9355);
or U14825 (N_14825,N_11002,N_9167);
nor U14826 (N_14826,N_6757,N_7340);
xor U14827 (N_14827,N_6796,N_9757);
xnor U14828 (N_14828,N_9080,N_9691);
nand U14829 (N_14829,N_8473,N_9091);
or U14830 (N_14830,N_6928,N_10068);
nor U14831 (N_14831,N_6484,N_10123);
nand U14832 (N_14832,N_7450,N_12463);
or U14833 (N_14833,N_12036,N_12205);
nand U14834 (N_14834,N_11780,N_12251);
nor U14835 (N_14835,N_8574,N_10622);
nand U14836 (N_14836,N_9444,N_10315);
or U14837 (N_14837,N_6741,N_12100);
nand U14838 (N_14838,N_8327,N_9917);
or U14839 (N_14839,N_12161,N_7105);
xnor U14840 (N_14840,N_10573,N_11019);
xor U14841 (N_14841,N_8301,N_7573);
nand U14842 (N_14842,N_9545,N_6723);
and U14843 (N_14843,N_11867,N_7836);
and U14844 (N_14844,N_8807,N_11252);
nand U14845 (N_14845,N_8430,N_7423);
xnor U14846 (N_14846,N_11317,N_8132);
or U14847 (N_14847,N_10966,N_8736);
or U14848 (N_14848,N_6473,N_6948);
nor U14849 (N_14849,N_11673,N_6999);
and U14850 (N_14850,N_8946,N_9674);
or U14851 (N_14851,N_6733,N_7084);
nor U14852 (N_14852,N_11138,N_11184);
nand U14853 (N_14853,N_8668,N_7051);
nand U14854 (N_14854,N_6295,N_11968);
nand U14855 (N_14855,N_9407,N_8666);
nand U14856 (N_14856,N_9042,N_12276);
nor U14857 (N_14857,N_9434,N_9770);
nand U14858 (N_14858,N_11752,N_6678);
and U14859 (N_14859,N_7239,N_10719);
and U14860 (N_14860,N_10067,N_9399);
nor U14861 (N_14861,N_10913,N_7265);
and U14862 (N_14862,N_7646,N_8129);
and U14863 (N_14863,N_9252,N_7643);
nand U14864 (N_14864,N_7574,N_11476);
nor U14865 (N_14865,N_12434,N_6858);
xor U14866 (N_14866,N_6663,N_6752);
nor U14867 (N_14867,N_11473,N_6511);
xnor U14868 (N_14868,N_6527,N_11005);
nor U14869 (N_14869,N_8139,N_10626);
nand U14870 (N_14870,N_12441,N_11240);
nor U14871 (N_14871,N_6581,N_9887);
xnor U14872 (N_14872,N_11271,N_8492);
or U14873 (N_14873,N_6700,N_8212);
nor U14874 (N_14874,N_6898,N_6860);
and U14875 (N_14875,N_8697,N_9303);
nand U14876 (N_14876,N_6356,N_7424);
nor U14877 (N_14877,N_11304,N_9597);
xnor U14878 (N_14878,N_9786,N_7262);
or U14879 (N_14879,N_10410,N_9912);
xor U14880 (N_14880,N_11512,N_9261);
xor U14881 (N_14881,N_11196,N_7837);
nand U14882 (N_14882,N_7840,N_12230);
nand U14883 (N_14883,N_12090,N_10648);
nor U14884 (N_14884,N_10721,N_9277);
or U14885 (N_14885,N_8607,N_6868);
xor U14886 (N_14886,N_9530,N_8712);
or U14887 (N_14887,N_12050,N_11291);
xor U14888 (N_14888,N_9416,N_12051);
xnor U14889 (N_14889,N_6809,N_11159);
or U14890 (N_14890,N_8226,N_7540);
or U14891 (N_14891,N_8865,N_10127);
and U14892 (N_14892,N_10985,N_7367);
nand U14893 (N_14893,N_9413,N_11776);
nand U14894 (N_14894,N_10760,N_10002);
and U14895 (N_14895,N_7317,N_12214);
or U14896 (N_14896,N_6786,N_7741);
xnor U14897 (N_14897,N_9998,N_11779);
nor U14898 (N_14898,N_12165,N_10629);
nor U14899 (N_14899,N_7666,N_11333);
xnor U14900 (N_14900,N_11978,N_10217);
or U14901 (N_14901,N_12071,N_11274);
nor U14902 (N_14902,N_9164,N_10131);
nor U14903 (N_14903,N_7388,N_9738);
nor U14904 (N_14904,N_10256,N_6412);
nor U14905 (N_14905,N_10426,N_9179);
and U14906 (N_14906,N_11029,N_8029);
nor U14907 (N_14907,N_10207,N_6401);
xor U14908 (N_14908,N_6337,N_8066);
xnor U14909 (N_14909,N_9675,N_9759);
xnor U14910 (N_14910,N_8592,N_12343);
xor U14911 (N_14911,N_6287,N_8635);
or U14912 (N_14912,N_7530,N_11481);
or U14913 (N_14913,N_10703,N_6674);
nand U14914 (N_14914,N_10559,N_10342);
xnor U14915 (N_14915,N_9713,N_6273);
nand U14916 (N_14916,N_11995,N_10837);
or U14917 (N_14917,N_6533,N_6869);
nand U14918 (N_14918,N_9211,N_9964);
nand U14919 (N_14919,N_9292,N_11608);
and U14920 (N_14920,N_6770,N_9532);
nor U14921 (N_14921,N_11644,N_6644);
or U14922 (N_14922,N_7282,N_11801);
nor U14923 (N_14923,N_7912,N_6885);
nor U14924 (N_14924,N_11518,N_6573);
nor U14925 (N_14925,N_8017,N_7538);
nand U14926 (N_14926,N_8180,N_10230);
or U14927 (N_14927,N_9878,N_8939);
nand U14928 (N_14928,N_7541,N_11124);
or U14929 (N_14929,N_10329,N_9402);
nor U14930 (N_14930,N_9538,N_12078);
nor U14931 (N_14931,N_7707,N_10572);
xor U14932 (N_14932,N_11619,N_7846);
and U14933 (N_14933,N_8383,N_10406);
or U14934 (N_14934,N_11639,N_9734);
xor U14935 (N_14935,N_10148,N_10929);
and U14936 (N_14936,N_8319,N_6353);
nand U14937 (N_14937,N_9460,N_8891);
and U14938 (N_14938,N_8245,N_10013);
or U14939 (N_14939,N_7011,N_12396);
and U14940 (N_14940,N_8090,N_9586);
and U14941 (N_14941,N_11083,N_9328);
or U14942 (N_14942,N_7461,N_8285);
nand U14943 (N_14943,N_9259,N_9916);
or U14944 (N_14944,N_6508,N_12072);
and U14945 (N_14945,N_10380,N_11172);
xnor U14946 (N_14946,N_11658,N_10322);
or U14947 (N_14947,N_10779,N_10577);
or U14948 (N_14948,N_9839,N_12221);
nor U14949 (N_14949,N_9780,N_10923);
xnor U14950 (N_14950,N_6284,N_10732);
xor U14951 (N_14951,N_8360,N_6781);
and U14952 (N_14952,N_11348,N_10803);
or U14953 (N_14953,N_6590,N_10866);
nand U14954 (N_14954,N_12124,N_6823);
and U14955 (N_14955,N_9502,N_8298);
nand U14956 (N_14956,N_11309,N_10646);
and U14957 (N_14957,N_9041,N_7035);
and U14958 (N_14958,N_10542,N_9026);
or U14959 (N_14959,N_8144,N_11307);
nor U14960 (N_14960,N_11059,N_11086);
nor U14961 (N_14961,N_9143,N_6956);
or U14962 (N_14962,N_9433,N_10302);
xnor U14963 (N_14963,N_7827,N_6803);
and U14964 (N_14964,N_7154,N_11704);
nor U14965 (N_14965,N_9622,N_6940);
nor U14966 (N_14966,N_8032,N_12268);
nor U14967 (N_14967,N_8919,N_6865);
xor U14968 (N_14968,N_10477,N_6844);
or U14969 (N_14969,N_6745,N_10620);
nor U14970 (N_14970,N_9459,N_10241);
or U14971 (N_14971,N_7392,N_7431);
and U14972 (N_14972,N_10226,N_11886);
and U14973 (N_14973,N_9989,N_10552);
nor U14974 (N_14974,N_11072,N_9300);
or U14975 (N_14975,N_7376,N_12213);
nor U14976 (N_14976,N_8222,N_7958);
nor U14977 (N_14977,N_8170,N_10361);
nor U14978 (N_14978,N_8102,N_6543);
xor U14979 (N_14979,N_11649,N_10597);
and U14980 (N_14980,N_12073,N_6615);
nor U14981 (N_14981,N_7597,N_9069);
or U14982 (N_14982,N_7168,N_9571);
nand U14983 (N_14983,N_9293,N_8511);
nor U14984 (N_14984,N_7867,N_12257);
or U14985 (N_14985,N_8521,N_10908);
or U14986 (N_14986,N_11898,N_7539);
and U14987 (N_14987,N_6489,N_12483);
xor U14988 (N_14988,N_8690,N_10143);
nand U14989 (N_14989,N_11648,N_10670);
or U14990 (N_14990,N_7025,N_7579);
nor U14991 (N_14991,N_9027,N_8159);
and U14992 (N_14992,N_9209,N_6342);
and U14993 (N_14993,N_12151,N_7935);
nor U14994 (N_14994,N_10717,N_10281);
nor U14995 (N_14995,N_6683,N_11255);
or U14996 (N_14996,N_6994,N_11262);
nor U14997 (N_14997,N_12032,N_6721);
nor U14998 (N_14998,N_9271,N_6611);
or U14999 (N_14999,N_8398,N_7124);
and U15000 (N_15000,N_10288,N_9851);
nor U15001 (N_15001,N_12342,N_8366);
and U15002 (N_15002,N_10110,N_6532);
and U15003 (N_15003,N_12319,N_11275);
nor U15004 (N_15004,N_7054,N_6895);
xnor U15005 (N_15005,N_10118,N_9267);
nand U15006 (N_15006,N_6742,N_9717);
xnor U15007 (N_15007,N_8077,N_8976);
or U15008 (N_15008,N_11320,N_10283);
nor U15009 (N_15009,N_11025,N_10820);
and U15010 (N_15010,N_8162,N_7789);
or U15011 (N_15011,N_8792,N_11444);
and U15012 (N_15012,N_8124,N_9983);
nand U15013 (N_15013,N_6600,N_10433);
and U15014 (N_15014,N_12042,N_11868);
xor U15015 (N_15015,N_12478,N_7508);
or U15016 (N_15016,N_11024,N_11178);
and U15017 (N_15017,N_9874,N_9994);
xor U15018 (N_15018,N_6893,N_6587);
or U15019 (N_15019,N_7913,N_12323);
and U15020 (N_15020,N_6963,N_7259);
and U15021 (N_15021,N_11061,N_7301);
nor U15022 (N_15022,N_10334,N_9837);
nor U15023 (N_15023,N_7357,N_9383);
or U15024 (N_15024,N_10790,N_11613);
and U15025 (N_15025,N_9601,N_7528);
xor U15026 (N_15026,N_7097,N_8958);
nand U15027 (N_15027,N_8232,N_8083);
or U15028 (N_15028,N_8779,N_8155);
or U15029 (N_15029,N_10589,N_12360);
or U15030 (N_15030,N_10508,N_8361);
xnor U15031 (N_15031,N_10774,N_10244);
or U15032 (N_15032,N_7411,N_7373);
and U15033 (N_15033,N_9474,N_7914);
nand U15034 (N_15034,N_9170,N_10484);
or U15035 (N_15035,N_9506,N_7456);
nor U15036 (N_15036,N_10113,N_6636);
and U15037 (N_15037,N_9059,N_7906);
and U15038 (N_15038,N_11525,N_8520);
nor U15039 (N_15039,N_10451,N_12411);
or U15040 (N_15040,N_6941,N_8991);
or U15041 (N_15041,N_11186,N_6256);
xor U15042 (N_15042,N_9843,N_8436);
and U15043 (N_15043,N_11228,N_9764);
xnor U15044 (N_15044,N_8960,N_10865);
nand U15045 (N_15045,N_8206,N_10897);
and U15046 (N_15046,N_11342,N_10036);
or U15047 (N_15047,N_9623,N_9283);
xor U15048 (N_15048,N_7475,N_8127);
or U15049 (N_15049,N_10254,N_8752);
and U15050 (N_15050,N_10232,N_9274);
or U15051 (N_15051,N_12003,N_9196);
and U15052 (N_15052,N_8659,N_6630);
or U15053 (N_15053,N_9658,N_10459);
xor U15054 (N_15054,N_9539,N_11246);
nor U15055 (N_15055,N_10712,N_8694);
nor U15056 (N_15056,N_7246,N_11520);
and U15057 (N_15057,N_9382,N_10887);
nor U15058 (N_15058,N_11162,N_9424);
nor U15059 (N_15059,N_9833,N_11813);
xnor U15060 (N_15060,N_12130,N_9265);
and U15061 (N_15061,N_8454,N_9892);
xor U15062 (N_15062,N_6660,N_9802);
xor U15063 (N_15063,N_9808,N_9554);
nand U15064 (N_15064,N_9943,N_9867);
xnor U15065 (N_15065,N_11187,N_12320);
and U15066 (N_15066,N_10713,N_12065);
nand U15067 (N_15067,N_8106,N_10199);
xor U15068 (N_15068,N_7618,N_10661);
or U15069 (N_15069,N_11699,N_7272);
nand U15070 (N_15070,N_10011,N_8909);
or U15071 (N_15071,N_7585,N_9454);
nor U15072 (N_15072,N_11468,N_10902);
nor U15073 (N_15073,N_7959,N_11585);
nor U15074 (N_15074,N_8470,N_12346);
nor U15075 (N_15075,N_7652,N_11601);
nand U15076 (N_15076,N_6453,N_11889);
or U15077 (N_15077,N_7902,N_7946);
xor U15078 (N_15078,N_11028,N_6625);
nor U15079 (N_15079,N_11952,N_6506);
xnor U15080 (N_15080,N_9375,N_7857);
xor U15081 (N_15081,N_8808,N_8388);
and U15082 (N_15082,N_11891,N_10976);
xor U15083 (N_15083,N_7095,N_9504);
and U15084 (N_15084,N_10449,N_11731);
nor U15085 (N_15085,N_10812,N_11496);
xor U15086 (N_15086,N_11871,N_7223);
or U15087 (N_15087,N_11686,N_10402);
or U15088 (N_15088,N_9595,N_11491);
nand U15089 (N_15089,N_12332,N_8507);
nor U15090 (N_15090,N_9888,N_9659);
nor U15091 (N_15091,N_8586,N_8952);
nor U15092 (N_15092,N_8906,N_6818);
nand U15093 (N_15093,N_10700,N_9859);
nand U15094 (N_15094,N_8777,N_8312);
xor U15095 (N_15095,N_11136,N_6847);
nand U15096 (N_15096,N_6441,N_10941);
nand U15097 (N_15097,N_8141,N_7993);
nor U15098 (N_15098,N_6727,N_10189);
nand U15099 (N_15099,N_10481,N_6612);
xor U15100 (N_15100,N_10129,N_10593);
and U15101 (N_15101,N_9769,N_7822);
or U15102 (N_15102,N_11733,N_7159);
xor U15103 (N_15103,N_11148,N_7761);
or U15104 (N_15104,N_11698,N_11599);
and U15105 (N_15105,N_11711,N_10370);
or U15106 (N_15106,N_11135,N_6726);
nor U15107 (N_15107,N_11897,N_11574);
and U15108 (N_15108,N_9344,N_9836);
nand U15109 (N_15109,N_8584,N_8803);
and U15110 (N_15110,N_8738,N_8972);
or U15111 (N_15111,N_7514,N_9148);
nor U15112 (N_15112,N_8974,N_6301);
nor U15113 (N_15113,N_6715,N_9309);
nand U15114 (N_15114,N_11279,N_12305);
nand U15115 (N_15115,N_9112,N_10468);
nor U15116 (N_15116,N_12103,N_10560);
or U15117 (N_15117,N_12096,N_6330);
or U15118 (N_15118,N_8645,N_9253);
nor U15119 (N_15119,N_11161,N_12293);
xnor U15120 (N_15120,N_10403,N_11283);
nor U15121 (N_15121,N_6882,N_7975);
or U15122 (N_15122,N_10156,N_9282);
nand U15123 (N_15123,N_10385,N_6343);
and U15124 (N_15124,N_8469,N_6996);
or U15125 (N_15125,N_7447,N_8377);
nor U15126 (N_15126,N_8441,N_7134);
or U15127 (N_15127,N_6756,N_10109);
nor U15128 (N_15128,N_6613,N_11418);
and U15129 (N_15129,N_11141,N_11943);
xnor U15130 (N_15130,N_6565,N_8256);
or U15131 (N_15131,N_9726,N_11947);
or U15132 (N_15132,N_8427,N_6272);
and U15133 (N_15133,N_7780,N_7998);
nand U15134 (N_15134,N_7422,N_7263);
nand U15135 (N_15135,N_7308,N_12306);
and U15136 (N_15136,N_12428,N_8595);
and U15137 (N_15137,N_9484,N_10726);
nand U15138 (N_15138,N_11310,N_9220);
nand U15139 (N_15139,N_8829,N_7248);
and U15140 (N_15140,N_8033,N_11671);
or U15141 (N_15141,N_7548,N_9716);
xnor U15142 (N_15142,N_8193,N_10657);
or U15143 (N_15143,N_6942,N_10090);
or U15144 (N_15144,N_11226,N_12304);
nor U15145 (N_15145,N_11093,N_9858);
or U15146 (N_15146,N_11642,N_10578);
and U15147 (N_15147,N_8311,N_6825);
nor U15148 (N_15148,N_9423,N_10708);
xor U15149 (N_15149,N_10608,N_8289);
nor U15150 (N_15150,N_9048,N_7838);
xor U15151 (N_15151,N_9920,N_6989);
nand U15152 (N_15152,N_8073,N_6320);
nor U15153 (N_15153,N_10438,N_10808);
nand U15154 (N_15154,N_6331,N_6767);
nor U15155 (N_15155,N_6378,N_10024);
or U15156 (N_15156,N_7425,N_8446);
and U15157 (N_15157,N_12056,N_11552);
xnor U15158 (N_15158,N_9217,N_7014);
xor U15159 (N_15159,N_9421,N_10323);
or U15160 (N_15160,N_8516,N_10016);
nor U15161 (N_15161,N_6774,N_11326);
and U15162 (N_15162,N_11369,N_11685);
nand U15163 (N_15163,N_11396,N_11458);
xor U15164 (N_15164,N_6340,N_11131);
nor U15165 (N_15165,N_11805,N_10368);
and U15166 (N_15166,N_11997,N_7409);
nor U15167 (N_15167,N_9714,N_7207);
and U15168 (N_15168,N_11336,N_7080);
or U15169 (N_15169,N_7872,N_10023);
nand U15170 (N_15170,N_8485,N_6688);
nor U15171 (N_15171,N_9877,N_8277);
nand U15172 (N_15172,N_6664,N_11289);
nand U15173 (N_15173,N_8630,N_8391);
or U15174 (N_15174,N_10082,N_9359);
nor U15175 (N_15175,N_10263,N_10800);
xor U15176 (N_15176,N_8959,N_8490);
and U15177 (N_15177,N_9023,N_8091);
xnor U15178 (N_15178,N_11220,N_9105);
nor U15179 (N_15179,N_6822,N_8893);
nand U15180 (N_15180,N_6424,N_11079);
xor U15181 (N_15181,N_9546,N_9728);
xor U15182 (N_15182,N_11744,N_6746);
nor U15183 (N_15183,N_6326,N_11454);
and U15184 (N_15184,N_9850,N_8272);
nand U15185 (N_15185,N_11917,N_11034);
nand U15186 (N_15186,N_6851,N_10676);
and U15187 (N_15187,N_6845,N_7631);
xor U15188 (N_15188,N_9117,N_9124);
nor U15189 (N_15189,N_9395,N_6593);
nor U15190 (N_15190,N_6867,N_10102);
or U15191 (N_15191,N_8654,N_7063);
or U15192 (N_15192,N_12243,N_11158);
nor U15193 (N_15193,N_12016,N_10446);
nand U15194 (N_15194,N_10170,N_10741);
nand U15195 (N_15195,N_7718,N_8401);
or U15196 (N_15196,N_6991,N_10491);
nand U15197 (N_15197,N_8305,N_8321);
xnor U15198 (N_15198,N_6924,N_10722);
nor U15199 (N_15199,N_9860,N_8747);
nand U15200 (N_15200,N_10432,N_8593);
or U15201 (N_15201,N_7963,N_8015);
or U15202 (N_15202,N_6360,N_10574);
or U15203 (N_15203,N_6879,N_7563);
or U15204 (N_15204,N_11012,N_10630);
nor U15205 (N_15205,N_10353,N_8056);
nor U15206 (N_15206,N_12067,N_11426);
nand U15207 (N_15207,N_12376,N_6932);
or U15208 (N_15208,N_6874,N_8266);
nand U15209 (N_15209,N_6540,N_6304);
or U15210 (N_15210,N_12388,N_10470);
nor U15211 (N_15211,N_6325,N_8290);
xor U15212 (N_15212,N_7359,N_7603);
nand U15213 (N_15213,N_8082,N_11505);
xnor U15214 (N_15214,N_12244,N_11134);
nor U15215 (N_15215,N_7571,N_10097);
or U15216 (N_15216,N_8205,N_11254);
xor U15217 (N_15217,N_7681,N_12131);
nor U15218 (N_15218,N_8692,N_7933);
or U15219 (N_15219,N_9928,N_7403);
nand U15220 (N_15220,N_10367,N_7947);
xor U15221 (N_15221,N_12414,N_10332);
and U15222 (N_15222,N_8650,N_7270);
and U15223 (N_15223,N_9992,N_11976);
xor U15224 (N_15224,N_9482,N_7065);
or U15225 (N_15225,N_10040,N_8781);
nand U15226 (N_15226,N_10462,N_7413);
xor U15227 (N_15227,N_9741,N_8502);
xnor U15228 (N_15228,N_8612,N_11382);
nor U15229 (N_15229,N_6341,N_6547);
nor U15230 (N_15230,N_6971,N_10640);
or U15231 (N_15231,N_7888,N_10931);
nor U15232 (N_15232,N_11085,N_12326);
nor U15233 (N_15233,N_6277,N_12199);
and U15234 (N_15234,N_8453,N_7158);
nor U15235 (N_15235,N_7820,N_9576);
or U15236 (N_15236,N_11352,N_6785);
or U15237 (N_15237,N_9751,N_9886);
or U15238 (N_15238,N_11904,N_9310);
nor U15239 (N_15239,N_11687,N_11910);
nand U15240 (N_15240,N_11869,N_7795);
and U15241 (N_15241,N_11078,N_7700);
and U15242 (N_15242,N_8249,N_8420);
xnor U15243 (N_15243,N_11785,N_12330);
or U15244 (N_15244,N_10526,N_11300);
nand U15245 (N_15245,N_8971,N_7477);
xor U15246 (N_15246,N_8902,N_12167);
or U15247 (N_15247,N_10169,N_7206);
nand U15248 (N_15248,N_10524,N_6522);
xor U15249 (N_15249,N_10341,N_7028);
nand U15250 (N_15250,N_6957,N_6798);
nand U15251 (N_15251,N_12358,N_8943);
and U15252 (N_15252,N_9644,N_9135);
nor U15253 (N_15253,N_10412,N_11227);
xor U15254 (N_15254,N_11366,N_9794);
nand U15255 (N_15255,N_10326,N_12379);
nand U15256 (N_15256,N_8138,N_8828);
or U15257 (N_15257,N_7073,N_8422);
or U15258 (N_15258,N_11171,N_9643);
and U15259 (N_15259,N_11436,N_11651);
nor U15260 (N_15260,N_6596,N_10513);
nand U15261 (N_15261,N_11866,N_9898);
and U15262 (N_15262,N_12339,N_9089);
or U15263 (N_15263,N_11380,N_10974);
xnor U15264 (N_15264,N_7617,N_11668);
xor U15265 (N_15265,N_9258,N_7764);
or U15266 (N_15266,N_11129,N_10829);
or U15267 (N_15267,N_11637,N_8653);
nor U15268 (N_15268,N_9390,N_11243);
and U15269 (N_15269,N_8407,N_6807);
nor U15270 (N_15270,N_11268,N_7110);
or U15271 (N_15271,N_11998,N_7399);
or U15272 (N_15272,N_11054,N_10656);
nor U15273 (N_15273,N_11936,N_10957);
nor U15274 (N_15274,N_11016,N_9600);
xor U15275 (N_15275,N_6379,N_6494);
nor U15276 (N_15276,N_10437,N_6555);
nand U15277 (N_15277,N_7297,N_6373);
and U15278 (N_15278,N_10407,N_7673);
and U15279 (N_15279,N_7295,N_7667);
xor U15280 (N_15280,N_12419,N_6986);
nand U15281 (N_15281,N_7547,N_10523);
xnor U15282 (N_15282,N_9879,N_9012);
and U15283 (N_15283,N_7067,N_10424);
nor U15284 (N_15284,N_7564,N_6512);
or U15285 (N_15285,N_9575,N_12259);
nand U15286 (N_15286,N_7068,N_7524);
or U15287 (N_15287,N_11355,N_11551);
nor U15288 (N_15288,N_10647,N_11675);
xnor U15289 (N_15289,N_6493,N_10533);
and U15290 (N_15290,N_7322,N_7072);
or U15291 (N_15291,N_12347,N_10398);
xor U15292 (N_15292,N_12422,N_10586);
nand U15293 (N_15293,N_6638,N_10688);
nand U15294 (N_15294,N_11536,N_8822);
or U15295 (N_15295,N_11361,N_9903);
and U15296 (N_15296,N_6712,N_9868);
and U15297 (N_15297,N_8762,N_9346);
xor U15298 (N_15298,N_10877,N_6470);
and U15299 (N_15299,N_6544,N_8857);
or U15300 (N_15300,N_7476,N_9771);
xor U15301 (N_15301,N_11624,N_12416);
and U15302 (N_15302,N_10333,N_8239);
xnor U15303 (N_15303,N_12249,N_8852);
and U15304 (N_15304,N_12018,N_11402);
nand U15305 (N_15305,N_9034,N_8252);
or U15306 (N_15306,N_8769,N_12294);
or U15307 (N_15307,N_7619,N_6691);
nor U15308 (N_15308,N_6578,N_9088);
nor U15309 (N_15309,N_7735,N_7816);
nor U15310 (N_15310,N_8872,N_12344);
and U15311 (N_15311,N_7169,N_11567);
nor U15312 (N_15312,N_6717,N_8445);
or U15313 (N_15313,N_6799,N_11467);
xnor U15314 (N_15314,N_7053,N_6400);
xor U15315 (N_15315,N_6311,N_10654);
xor U15316 (N_15316,N_6939,N_8364);
nor U15317 (N_15317,N_11053,N_10891);
or U15318 (N_15318,N_7924,N_9834);
or U15319 (N_15319,N_6689,N_11044);
and U15320 (N_15320,N_8928,N_12191);
xor U15321 (N_15321,N_9971,N_11912);
or U15322 (N_15322,N_10287,N_10822);
nand U15323 (N_15323,N_7581,N_12228);
and U15324 (N_15324,N_9933,N_8801);
nand U15325 (N_15325,N_8274,N_8660);
or U15326 (N_15326,N_8477,N_9144);
nor U15327 (N_15327,N_8049,N_10527);
and U15328 (N_15328,N_7018,N_6570);
nor U15329 (N_15329,N_10906,N_11351);
nand U15330 (N_15330,N_7290,N_7629);
and U15331 (N_15331,N_9323,N_7310);
or U15332 (N_15332,N_6708,N_8335);
and U15333 (N_15333,N_11508,N_6314);
and U15334 (N_15334,N_8505,N_9473);
nand U15335 (N_15335,N_11185,N_12299);
and U15336 (N_15336,N_12206,N_10376);
or U15337 (N_15337,N_11715,N_8647);
nor U15338 (N_15338,N_7588,N_11163);
or U15339 (N_15339,N_10439,N_10220);
and U15340 (N_15340,N_10506,N_7910);
and U15341 (N_15341,N_11728,N_6946);
and U15342 (N_15342,N_6607,N_10400);
and U15343 (N_15343,N_10948,N_8610);
and U15344 (N_15344,N_8120,N_8740);
nand U15345 (N_15345,N_10421,N_8811);
xor U15346 (N_15346,N_10206,N_7944);
nand U15347 (N_15347,N_8606,N_11373);
or U15348 (N_15348,N_9437,N_9030);
nor U15349 (N_15349,N_7870,N_8793);
nand U15350 (N_15350,N_7076,N_6492);
nand U15351 (N_15351,N_9730,N_7633);
nand U15352 (N_15352,N_6427,N_10967);
or U15353 (N_15353,N_6566,N_11643);
xnor U15354 (N_15354,N_10835,N_11230);
nor U15355 (N_15355,N_6359,N_12182);
xnor U15356 (N_15356,N_11893,N_6302);
nand U15357 (N_15357,N_6753,N_11117);
and U15358 (N_15358,N_11281,N_9625);
xor U15359 (N_15359,N_10946,N_11963);
nand U15360 (N_15360,N_8044,N_11064);
nand U15361 (N_15361,N_9001,N_12282);
nor U15362 (N_15362,N_11669,N_9766);
and U15363 (N_15363,N_6592,N_10935);
and U15364 (N_15364,N_10033,N_10711);
nor U15365 (N_15365,N_9127,N_7521);
nor U15366 (N_15366,N_12186,N_11594);
xor U15367 (N_15367,N_8951,N_11374);
and U15368 (N_15368,N_11322,N_9404);
nor U15369 (N_15369,N_6800,N_11335);
nor U15370 (N_15370,N_11879,N_10138);
or U15371 (N_15371,N_11993,N_8456);
and U15372 (N_15372,N_10176,N_11734);
nor U15373 (N_15373,N_7198,N_8016);
xor U15374 (N_15374,N_8264,N_12491);
or U15375 (N_15375,N_6450,N_6641);
and U15376 (N_15376,N_11652,N_12269);
nor U15377 (N_15377,N_6516,N_9082);
or U15378 (N_15378,N_6950,N_12399);
and U15379 (N_15379,N_10157,N_6283);
nor U15380 (N_15380,N_7668,N_6900);
and U15381 (N_15381,N_10436,N_7151);
nor U15382 (N_15382,N_10770,N_9638);
and U15383 (N_15383,N_6913,N_10535);
or U15384 (N_15384,N_6609,N_12345);
nor U15385 (N_15385,N_11142,N_6855);
or U15386 (N_15386,N_10521,N_8095);
nor U15387 (N_15387,N_8117,N_9125);
or U15388 (N_15388,N_7662,N_10185);
or U15389 (N_15389,N_9679,N_8217);
or U15390 (N_15390,N_11958,N_9142);
nand U15391 (N_15391,N_6567,N_10492);
xnor U15392 (N_15392,N_6750,N_12026);
nor U15393 (N_15393,N_10178,N_9448);
nand U15394 (N_15394,N_11014,N_6420);
or U15395 (N_15395,N_8895,N_9608);
nor U15396 (N_15396,N_8760,N_10668);
xnor U15397 (N_15397,N_8904,N_10253);
nand U15398 (N_15398,N_9984,N_11229);
xnor U15399 (N_15399,N_10801,N_12217);
and U15400 (N_15400,N_9169,N_6623);
nand U15401 (N_15401,N_9157,N_9075);
and U15402 (N_15402,N_6889,N_8794);
or U15403 (N_15403,N_12386,N_9552);
or U15404 (N_15404,N_11555,N_10529);
nand U15405 (N_15405,N_6736,N_6789);
xor U15406 (N_15406,N_7788,N_9743);
and U15407 (N_15407,N_11364,N_7569);
and U15408 (N_15408,N_7337,N_9512);
nor U15409 (N_15409,N_11153,N_10635);
xor U15410 (N_15410,N_7370,N_7791);
and U15411 (N_15411,N_11545,N_10953);
nor U15412 (N_15412,N_9599,N_8253);
or U15413 (N_15413,N_10172,N_8260);
or U15414 (N_15414,N_6817,N_7384);
nand U15415 (N_15415,N_7866,N_7205);
or U15416 (N_15416,N_6524,N_7981);
and U15417 (N_15417,N_9665,N_10087);
nand U15418 (N_15418,N_9950,N_8060);
xor U15419 (N_15419,N_12364,N_10003);
and U15420 (N_15420,N_10490,N_8914);
nand U15421 (N_15421,N_12179,N_7928);
or U15422 (N_15422,N_7486,N_9486);
xnor U15423 (N_15423,N_12470,N_9553);
or U15424 (N_15424,N_10101,N_11000);
nand U15425 (N_15425,N_9753,N_8616);
nor U15426 (N_15426,N_9000,N_6413);
nand U15427 (N_15427,N_11975,N_12145);
xnor U15428 (N_15428,N_8078,N_6291);
and U15429 (N_15429,N_11663,N_9349);
nand U15430 (N_15430,N_7174,N_11105);
or U15431 (N_15431,N_8036,N_9518);
or U15432 (N_15432,N_7126,N_12486);
xnor U15433 (N_15433,N_10075,N_8265);
nor U15434 (N_15434,N_11782,N_10671);
and U15435 (N_15435,N_8067,N_7650);
nor U15436 (N_15436,N_10917,N_11242);
nor U15437 (N_15437,N_12083,N_11430);
xnor U15438 (N_15438,N_10758,N_12292);
xor U15439 (N_15439,N_7146,N_7214);
nand U15440 (N_15440,N_6350,N_9496);
and U15441 (N_15441,N_9198,N_7685);
nand U15442 (N_15442,N_8890,N_11761);
nand U15443 (N_15443,N_9590,N_11107);
and U15444 (N_15444,N_6447,N_6366);
nor U15445 (N_15445,N_7871,N_8594);
xor U15446 (N_15446,N_6886,N_12057);
xnor U15447 (N_15447,N_6439,N_9827);
nor U15448 (N_15448,N_12148,N_7784);
nand U15449 (N_15449,N_11081,N_8728);
nand U15450 (N_15450,N_9513,N_9614);
nand U15451 (N_15451,N_8863,N_10115);
and U15452 (N_15452,N_11905,N_8333);
or U15453 (N_15453,N_9615,N_10880);
or U15454 (N_15454,N_9966,N_7122);
nor U15455 (N_15455,N_9854,N_12203);
or U15456 (N_15456,N_11982,N_8061);
nand U15457 (N_15457,N_11195,N_12104);
or U15458 (N_15458,N_6634,N_11213);
or U15459 (N_15459,N_7510,N_7783);
xor U15460 (N_15460,N_6539,N_7480);
nor U15461 (N_15461,N_12493,N_7960);
nor U15462 (N_15462,N_9494,N_8804);
nand U15463 (N_15463,N_11026,N_6463);
or U15464 (N_15464,N_10551,N_6479);
or U15465 (N_15465,N_9208,N_8831);
or U15466 (N_15466,N_6606,N_7661);
and U15467 (N_15467,N_9409,N_12008);
nand U15468 (N_15468,N_11412,N_10771);
nor U15469 (N_15469,N_12436,N_11767);
xor U15470 (N_15470,N_11892,N_8618);
nand U15471 (N_15471,N_7237,N_6951);
and U15472 (N_15472,N_11048,N_8046);
or U15473 (N_15473,N_8938,N_6977);
xnor U15474 (N_15474,N_11750,N_6927);
xnor U15475 (N_15475,N_9534,N_8550);
xor U15476 (N_15476,N_9189,N_9968);
or U15477 (N_15477,N_11177,N_11073);
xnor U15478 (N_15478,N_7587,N_11996);
and U15479 (N_15479,N_11962,N_7845);
or U15480 (N_15480,N_6929,N_11864);
xor U15481 (N_15481,N_11493,N_7757);
or U15482 (N_15482,N_6722,N_11301);
or U15483 (N_15483,N_9606,N_7005);
or U15484 (N_15484,N_11944,N_6949);
and U15485 (N_15485,N_7352,N_7813);
and U15486 (N_15486,N_7951,N_9305);
nand U15487 (N_15487,N_7175,N_8022);
nor U15488 (N_15488,N_9489,N_6383);
nor U15489 (N_15489,N_7536,N_11344);
or U15490 (N_15490,N_11862,N_8932);
nand U15491 (N_15491,N_9740,N_8385);
and U15492 (N_15492,N_8855,N_6618);
nand U15493 (N_15493,N_11329,N_8601);
nand U15494 (N_15494,N_10959,N_9913);
xnor U15495 (N_15495,N_9584,N_8465);
nor U15496 (N_15496,N_11951,N_7663);
or U15497 (N_15497,N_7100,N_7799);
xnor U15498 (N_15498,N_9184,N_10442);
nor U15499 (N_15499,N_7346,N_8968);
xnor U15500 (N_15500,N_6442,N_6985);
and U15501 (N_15501,N_10961,N_10318);
xor U15502 (N_15502,N_11939,N_11126);
or U15503 (N_15503,N_9567,N_6990);
nand U15504 (N_15504,N_7460,N_11076);
or U15505 (N_15505,N_10693,N_10583);
and U15506 (N_15506,N_7940,N_6345);
nand U15507 (N_15507,N_7555,N_6790);
or U15508 (N_15508,N_10317,N_8207);
xor U15509 (N_15509,N_8866,N_11654);
or U15510 (N_15510,N_6744,N_10802);
and U15511 (N_15511,N_9931,N_6588);
and U15512 (N_15512,N_11007,N_9275);
xor U15513 (N_15513,N_8718,N_11942);
nor U15514 (N_15514,N_11357,N_7777);
xor U15515 (N_15515,N_8698,N_6279);
nor U15516 (N_15516,N_7294,N_8588);
xor U15517 (N_15517,N_11832,N_9190);
nor U15518 (N_15518,N_11503,N_9648);
xnor U15519 (N_15519,N_9960,N_9031);
and U15520 (N_15520,N_9203,N_10060);
nor U15521 (N_15521,N_8440,N_9313);
or U15522 (N_15522,N_7086,N_9350);
and U15523 (N_15523,N_7182,N_8458);
and U15524 (N_15524,N_11416,N_9866);
nor U15525 (N_15525,N_7760,N_9442);
and U15526 (N_15526,N_8501,N_8494);
xor U15527 (N_15527,N_8352,N_8021);
and U15528 (N_15528,N_8279,N_11022);
nor U15529 (N_15529,N_6564,N_9295);
or U15530 (N_15530,N_10603,N_10343);
xnor U15531 (N_15531,N_7894,N_10581);
nand U15532 (N_15532,N_8399,N_7927);
nor U15533 (N_15533,N_11616,N_7320);
and U15534 (N_15534,N_10295,N_9816);
nor U15535 (N_15535,N_7710,N_6831);
xnor U15536 (N_15536,N_12134,N_7330);
xnor U15537 (N_15537,N_11941,N_6627);
or U15538 (N_15538,N_11459,N_6561);
nor U15539 (N_15539,N_6445,N_6992);
and U15540 (N_15540,N_8649,N_9116);
nor U15541 (N_15541,N_7776,N_11181);
nand U15542 (N_15542,N_9319,N_12135);
nand U15543 (N_15543,N_10235,N_6297);
or U15544 (N_15544,N_7773,N_8488);
nand U15545 (N_15545,N_10998,N_11045);
or U15546 (N_15546,N_8515,N_6685);
nand U15547 (N_15547,N_6856,N_9671);
nand U15548 (N_15548,N_9609,N_8888);
and U15549 (N_15549,N_7922,N_11190);
or U15550 (N_15550,N_8438,N_7896);
or U15551 (N_15551,N_11152,N_11070);
or U15552 (N_15552,N_11104,N_11592);
nand U15553 (N_15553,N_11840,N_12110);
nor U15554 (N_15554,N_11311,N_6687);
or U15555 (N_15555,N_10019,N_11740);
nor U15556 (N_15556,N_9426,N_9373);
nor U15557 (N_15557,N_9449,N_10203);
nand U15558 (N_15558,N_10867,N_9230);
xor U15559 (N_15559,N_10262,N_6980);
nand U15560 (N_15560,N_6603,N_7030);
or U15561 (N_15561,N_9556,N_8103);
or U15562 (N_15562,N_8726,N_6346);
or U15563 (N_15563,N_10645,N_6496);
xnor U15564 (N_15564,N_7808,N_7074);
and U15565 (N_15565,N_11431,N_6810);
xnor U15566 (N_15566,N_9004,N_10378);
or U15567 (N_15567,N_9965,N_9687);
and U15568 (N_15568,N_11208,N_8276);
nor U15569 (N_15569,N_11890,N_10050);
nand U15570 (N_15570,N_8246,N_6854);
or U15571 (N_15571,N_8886,N_11023);
nor U15572 (N_15572,N_11440,N_9377);
nand U15573 (N_15573,N_12229,N_12102);
nor U15574 (N_15574,N_9439,N_7203);
xnor U15575 (N_15575,N_12406,N_7230);
or U15576 (N_15576,N_8122,N_8570);
nand U15577 (N_15577,N_9370,N_8920);
or U15578 (N_15578,N_11460,N_8413);
nor U15579 (N_15579,N_6899,N_7329);
and U15580 (N_15580,N_10006,N_12413);
and U15581 (N_15581,N_10072,N_6813);
xnor U15582 (N_15582,N_10114,N_7785);
nor U15583 (N_15583,N_11808,N_11408);
nand U15584 (N_15584,N_11709,N_9702);
xnor U15585 (N_15585,N_12377,N_8434);
or U15586 (N_15586,N_11245,N_7817);
nand U15587 (N_15587,N_7009,N_12114);
nand U15588 (N_15588,N_7481,N_9242);
or U15589 (N_15589,N_8759,N_8304);
nand U15590 (N_15590,N_8964,N_12402);
and U15591 (N_15591,N_7145,N_11915);
nor U15592 (N_15592,N_10061,N_9078);
nor U15593 (N_15593,N_11961,N_9587);
or U15594 (N_15594,N_12351,N_8378);
and U15595 (N_15595,N_6405,N_7439);
nand U15596 (N_15596,N_7985,N_7037);
nor U15597 (N_15597,N_10348,N_10653);
nand U15598 (N_15598,N_9162,N_10215);
nor U15599 (N_15599,N_12099,N_9411);
or U15600 (N_15600,N_12069,N_10211);
nor U15601 (N_15601,N_6368,N_10673);
nand U15602 (N_15602,N_9254,N_6972);
xnor U15603 (N_15603,N_6834,N_6339);
xor U15604 (N_15604,N_10397,N_7303);
nor U15605 (N_15605,N_6562,N_9901);
xnor U15606 (N_15606,N_7991,N_12129);
nor U15607 (N_15607,N_7031,N_8923);
nor U15608 (N_15608,N_8933,N_11748);
and U15609 (N_15609,N_11175,N_12290);
and U15610 (N_15610,N_10512,N_6743);
and U15611 (N_15611,N_7550,N_10871);
nor U15612 (N_15612,N_9074,N_8457);
nand U15613 (N_15613,N_7931,N_8887);
nor U15614 (N_15614,N_8426,N_8443);
or U15615 (N_15615,N_11565,N_11873);
xor U15616 (N_15616,N_10233,N_12059);
or U15617 (N_15617,N_11340,N_8815);
and U15618 (N_15618,N_12278,N_6758);
nand U15619 (N_15619,N_6446,N_9263);
or U15620 (N_15620,N_10161,N_6622);
and U15621 (N_15621,N_10505,N_11216);
nor U15622 (N_15622,N_12170,N_8941);
and U15623 (N_15623,N_7527,N_6460);
nand U15624 (N_15624,N_12387,N_11272);
xor U15625 (N_15625,N_6718,N_8997);
and U15626 (N_15626,N_10913,N_11732);
or U15627 (N_15627,N_10666,N_9759);
or U15628 (N_15628,N_6774,N_12236);
nand U15629 (N_15629,N_11200,N_8223);
or U15630 (N_15630,N_6980,N_11449);
nand U15631 (N_15631,N_12460,N_9082);
xnor U15632 (N_15632,N_10959,N_7625);
nor U15633 (N_15633,N_7644,N_8387);
xor U15634 (N_15634,N_10803,N_12256);
nand U15635 (N_15635,N_8490,N_11636);
and U15636 (N_15636,N_9935,N_8691);
nor U15637 (N_15637,N_6578,N_9465);
and U15638 (N_15638,N_11378,N_9487);
and U15639 (N_15639,N_6516,N_11418);
nand U15640 (N_15640,N_8180,N_6742);
nor U15641 (N_15641,N_10100,N_11336);
or U15642 (N_15642,N_7708,N_7644);
nand U15643 (N_15643,N_8532,N_12341);
xnor U15644 (N_15644,N_7466,N_7024);
or U15645 (N_15645,N_11914,N_8584);
and U15646 (N_15646,N_12179,N_10131);
nand U15647 (N_15647,N_9961,N_6378);
or U15648 (N_15648,N_10474,N_11005);
and U15649 (N_15649,N_11228,N_7423);
nand U15650 (N_15650,N_10215,N_7824);
nand U15651 (N_15651,N_8328,N_7569);
and U15652 (N_15652,N_6612,N_7913);
nor U15653 (N_15653,N_8659,N_7555);
or U15654 (N_15654,N_12339,N_11269);
xnor U15655 (N_15655,N_7570,N_11401);
and U15656 (N_15656,N_9850,N_7270);
nor U15657 (N_15657,N_9569,N_12303);
and U15658 (N_15658,N_11279,N_7468);
xor U15659 (N_15659,N_9989,N_12224);
xor U15660 (N_15660,N_12331,N_10319);
or U15661 (N_15661,N_8538,N_10790);
nand U15662 (N_15662,N_7292,N_7676);
nand U15663 (N_15663,N_7562,N_11447);
nand U15664 (N_15664,N_11065,N_12487);
or U15665 (N_15665,N_8896,N_9090);
xnor U15666 (N_15666,N_10641,N_11338);
and U15667 (N_15667,N_7243,N_9383);
or U15668 (N_15668,N_7818,N_11875);
xnor U15669 (N_15669,N_9995,N_7421);
nor U15670 (N_15670,N_7486,N_6882);
xnor U15671 (N_15671,N_11230,N_11298);
or U15672 (N_15672,N_9655,N_12170);
and U15673 (N_15673,N_10275,N_6650);
xor U15674 (N_15674,N_10335,N_11960);
nor U15675 (N_15675,N_9516,N_8284);
or U15676 (N_15676,N_9716,N_9379);
nand U15677 (N_15677,N_8735,N_9646);
nand U15678 (N_15678,N_6746,N_9344);
nor U15679 (N_15679,N_10661,N_12187);
and U15680 (N_15680,N_8476,N_10099);
xor U15681 (N_15681,N_6396,N_7713);
nand U15682 (N_15682,N_7400,N_10643);
nor U15683 (N_15683,N_11466,N_9950);
and U15684 (N_15684,N_9659,N_11918);
xor U15685 (N_15685,N_6290,N_8646);
or U15686 (N_15686,N_8898,N_10243);
nand U15687 (N_15687,N_6744,N_6479);
xor U15688 (N_15688,N_10863,N_9819);
nand U15689 (N_15689,N_9623,N_6822);
nand U15690 (N_15690,N_10941,N_7279);
and U15691 (N_15691,N_9955,N_9718);
xnor U15692 (N_15692,N_11686,N_6397);
or U15693 (N_15693,N_11431,N_9643);
xor U15694 (N_15694,N_11971,N_8441);
xnor U15695 (N_15695,N_9662,N_12320);
xnor U15696 (N_15696,N_6737,N_6561);
nand U15697 (N_15697,N_6258,N_11803);
xor U15698 (N_15698,N_8881,N_8358);
or U15699 (N_15699,N_7191,N_6656);
nor U15700 (N_15700,N_12253,N_12002);
nand U15701 (N_15701,N_6668,N_7929);
nor U15702 (N_15702,N_9374,N_9238);
and U15703 (N_15703,N_10721,N_6736);
nand U15704 (N_15704,N_9094,N_8459);
and U15705 (N_15705,N_7492,N_10467);
or U15706 (N_15706,N_6529,N_11283);
and U15707 (N_15707,N_7497,N_8366);
nand U15708 (N_15708,N_6914,N_11464);
nand U15709 (N_15709,N_8195,N_6660);
xnor U15710 (N_15710,N_8025,N_8428);
and U15711 (N_15711,N_7735,N_7917);
or U15712 (N_15712,N_10088,N_11823);
and U15713 (N_15713,N_10941,N_7088);
and U15714 (N_15714,N_6864,N_8352);
nor U15715 (N_15715,N_11784,N_11365);
or U15716 (N_15716,N_6949,N_9477);
or U15717 (N_15717,N_9197,N_7762);
xnor U15718 (N_15718,N_9097,N_7986);
nor U15719 (N_15719,N_7686,N_6339);
nand U15720 (N_15720,N_8237,N_6504);
nor U15721 (N_15721,N_7468,N_6844);
xnor U15722 (N_15722,N_6754,N_9460);
and U15723 (N_15723,N_7414,N_7453);
nor U15724 (N_15724,N_9400,N_8721);
and U15725 (N_15725,N_10524,N_9404);
nor U15726 (N_15726,N_8552,N_7676);
and U15727 (N_15727,N_7495,N_10256);
xnor U15728 (N_15728,N_9558,N_8426);
and U15729 (N_15729,N_6373,N_11247);
xnor U15730 (N_15730,N_10189,N_10000);
nand U15731 (N_15731,N_10739,N_8277);
xnor U15732 (N_15732,N_7048,N_8326);
nor U15733 (N_15733,N_9137,N_10050);
and U15734 (N_15734,N_12268,N_10778);
nor U15735 (N_15735,N_6374,N_6616);
nor U15736 (N_15736,N_11059,N_8638);
and U15737 (N_15737,N_7444,N_10981);
nand U15738 (N_15738,N_9236,N_10367);
nor U15739 (N_15739,N_6474,N_11727);
xnor U15740 (N_15740,N_11181,N_10153);
nand U15741 (N_15741,N_10230,N_9469);
nor U15742 (N_15742,N_11988,N_8716);
xor U15743 (N_15743,N_9095,N_11609);
nand U15744 (N_15744,N_10411,N_10375);
nor U15745 (N_15745,N_8014,N_7751);
or U15746 (N_15746,N_8326,N_8641);
or U15747 (N_15747,N_8785,N_12287);
nand U15748 (N_15748,N_7851,N_9872);
xor U15749 (N_15749,N_7421,N_6254);
or U15750 (N_15750,N_10633,N_8105);
and U15751 (N_15751,N_8415,N_11461);
nor U15752 (N_15752,N_9834,N_6568);
or U15753 (N_15753,N_9462,N_8422);
and U15754 (N_15754,N_7081,N_10880);
nor U15755 (N_15755,N_11896,N_11269);
nand U15756 (N_15756,N_12175,N_7279);
xnor U15757 (N_15757,N_8273,N_12075);
nor U15758 (N_15758,N_8648,N_8628);
xnor U15759 (N_15759,N_7572,N_9838);
nand U15760 (N_15760,N_6594,N_9603);
or U15761 (N_15761,N_6852,N_10291);
or U15762 (N_15762,N_6828,N_6976);
nor U15763 (N_15763,N_9569,N_10286);
nand U15764 (N_15764,N_6549,N_6606);
xnor U15765 (N_15765,N_9581,N_7992);
nor U15766 (N_15766,N_8632,N_7501);
xor U15767 (N_15767,N_10804,N_7490);
nand U15768 (N_15768,N_11284,N_10130);
and U15769 (N_15769,N_9675,N_11968);
nand U15770 (N_15770,N_8051,N_10296);
and U15771 (N_15771,N_10819,N_11228);
xor U15772 (N_15772,N_9523,N_7708);
nor U15773 (N_15773,N_7274,N_11962);
nand U15774 (N_15774,N_8508,N_10641);
xor U15775 (N_15775,N_8670,N_8416);
or U15776 (N_15776,N_10544,N_6340);
or U15777 (N_15777,N_10578,N_7211);
nand U15778 (N_15778,N_6395,N_7406);
xnor U15779 (N_15779,N_8700,N_7178);
and U15780 (N_15780,N_9346,N_7472);
nand U15781 (N_15781,N_10369,N_8330);
or U15782 (N_15782,N_8630,N_9443);
xnor U15783 (N_15783,N_7101,N_6293);
xnor U15784 (N_15784,N_12327,N_11271);
or U15785 (N_15785,N_6495,N_12222);
nor U15786 (N_15786,N_10831,N_11263);
xor U15787 (N_15787,N_10283,N_9952);
nand U15788 (N_15788,N_12412,N_6898);
xor U15789 (N_15789,N_9048,N_7365);
and U15790 (N_15790,N_9488,N_8023);
nor U15791 (N_15791,N_8289,N_7037);
and U15792 (N_15792,N_8156,N_10035);
and U15793 (N_15793,N_10124,N_12393);
xnor U15794 (N_15794,N_7010,N_11198);
nor U15795 (N_15795,N_6845,N_6807);
nor U15796 (N_15796,N_7769,N_9357);
nand U15797 (N_15797,N_9694,N_11795);
and U15798 (N_15798,N_10004,N_6725);
xor U15799 (N_15799,N_6289,N_12073);
nand U15800 (N_15800,N_8131,N_8865);
nor U15801 (N_15801,N_9793,N_8073);
xor U15802 (N_15802,N_6964,N_11864);
nand U15803 (N_15803,N_7893,N_7934);
and U15804 (N_15804,N_12039,N_10636);
nand U15805 (N_15805,N_7119,N_8295);
nand U15806 (N_15806,N_12111,N_9209);
xnor U15807 (N_15807,N_10030,N_11164);
nand U15808 (N_15808,N_8159,N_8638);
xnor U15809 (N_15809,N_8748,N_7863);
and U15810 (N_15810,N_11840,N_12123);
and U15811 (N_15811,N_8511,N_8331);
or U15812 (N_15812,N_11914,N_11680);
nor U15813 (N_15813,N_12357,N_10635);
or U15814 (N_15814,N_11093,N_8400);
nor U15815 (N_15815,N_7256,N_11452);
and U15816 (N_15816,N_12372,N_6983);
nor U15817 (N_15817,N_7713,N_12321);
and U15818 (N_15818,N_11650,N_8510);
and U15819 (N_15819,N_9225,N_6566);
xor U15820 (N_15820,N_7104,N_6454);
or U15821 (N_15821,N_11673,N_7760);
or U15822 (N_15822,N_11194,N_10771);
nand U15823 (N_15823,N_10215,N_10510);
nor U15824 (N_15824,N_9756,N_9903);
or U15825 (N_15825,N_8860,N_10261);
nor U15826 (N_15826,N_9296,N_11592);
nand U15827 (N_15827,N_10250,N_12322);
and U15828 (N_15828,N_8152,N_7990);
xnor U15829 (N_15829,N_10501,N_10421);
or U15830 (N_15830,N_12146,N_7588);
and U15831 (N_15831,N_9622,N_6586);
nand U15832 (N_15832,N_12111,N_8784);
xnor U15833 (N_15833,N_11886,N_9199);
and U15834 (N_15834,N_11710,N_12090);
nor U15835 (N_15835,N_11171,N_7179);
nor U15836 (N_15836,N_11910,N_7461);
or U15837 (N_15837,N_12374,N_12236);
nand U15838 (N_15838,N_7605,N_8073);
and U15839 (N_15839,N_7087,N_6265);
nand U15840 (N_15840,N_6494,N_6988);
nor U15841 (N_15841,N_11561,N_12131);
xor U15842 (N_15842,N_11733,N_10624);
xor U15843 (N_15843,N_12333,N_7599);
nand U15844 (N_15844,N_6616,N_11254);
xnor U15845 (N_15845,N_7154,N_6507);
nor U15846 (N_15846,N_8183,N_6926);
and U15847 (N_15847,N_10354,N_9088);
nor U15848 (N_15848,N_11504,N_11908);
nor U15849 (N_15849,N_7175,N_9075);
and U15850 (N_15850,N_8856,N_8358);
and U15851 (N_15851,N_9482,N_9716);
and U15852 (N_15852,N_10540,N_10061);
nor U15853 (N_15853,N_11783,N_6711);
xor U15854 (N_15854,N_9801,N_9446);
xnor U15855 (N_15855,N_10018,N_11642);
or U15856 (N_15856,N_6675,N_9462);
nand U15857 (N_15857,N_8689,N_12143);
nor U15858 (N_15858,N_7692,N_11979);
nor U15859 (N_15859,N_10650,N_8279);
nor U15860 (N_15860,N_9504,N_8260);
nor U15861 (N_15861,N_8804,N_8340);
or U15862 (N_15862,N_9108,N_10183);
xor U15863 (N_15863,N_10021,N_6716);
xor U15864 (N_15864,N_8867,N_8785);
and U15865 (N_15865,N_7935,N_8489);
nand U15866 (N_15866,N_6992,N_10918);
xnor U15867 (N_15867,N_10870,N_11505);
and U15868 (N_15868,N_10358,N_8918);
nor U15869 (N_15869,N_11358,N_10986);
xor U15870 (N_15870,N_6650,N_7273);
and U15871 (N_15871,N_10139,N_7771);
and U15872 (N_15872,N_7457,N_6251);
and U15873 (N_15873,N_9130,N_10363);
nand U15874 (N_15874,N_6546,N_8248);
xnor U15875 (N_15875,N_12469,N_9398);
or U15876 (N_15876,N_9225,N_11340);
and U15877 (N_15877,N_10129,N_10270);
or U15878 (N_15878,N_9896,N_7700);
nand U15879 (N_15879,N_6903,N_8134);
nand U15880 (N_15880,N_7809,N_9393);
and U15881 (N_15881,N_9412,N_9585);
nor U15882 (N_15882,N_12471,N_12328);
or U15883 (N_15883,N_9305,N_11444);
or U15884 (N_15884,N_8000,N_8270);
xnor U15885 (N_15885,N_8112,N_9189);
or U15886 (N_15886,N_6252,N_7544);
or U15887 (N_15887,N_11036,N_6395);
nand U15888 (N_15888,N_6934,N_9101);
and U15889 (N_15889,N_8469,N_10772);
or U15890 (N_15890,N_8321,N_7073);
and U15891 (N_15891,N_10788,N_8082);
nand U15892 (N_15892,N_11347,N_6952);
or U15893 (N_15893,N_7716,N_10410);
and U15894 (N_15894,N_11587,N_11742);
or U15895 (N_15895,N_7421,N_10029);
or U15896 (N_15896,N_8104,N_8650);
or U15897 (N_15897,N_6734,N_11699);
or U15898 (N_15898,N_6854,N_11685);
and U15899 (N_15899,N_6874,N_6498);
nand U15900 (N_15900,N_6745,N_8366);
nand U15901 (N_15901,N_8841,N_6923);
nand U15902 (N_15902,N_12322,N_7948);
nand U15903 (N_15903,N_6846,N_10553);
nor U15904 (N_15904,N_7129,N_6537);
nand U15905 (N_15905,N_6627,N_11898);
nand U15906 (N_15906,N_10666,N_6434);
and U15907 (N_15907,N_10537,N_9453);
xor U15908 (N_15908,N_8873,N_12021);
xnor U15909 (N_15909,N_6883,N_6910);
or U15910 (N_15910,N_7497,N_10445);
or U15911 (N_15911,N_7682,N_11251);
nor U15912 (N_15912,N_11439,N_9989);
and U15913 (N_15913,N_11341,N_10673);
nor U15914 (N_15914,N_11370,N_8064);
or U15915 (N_15915,N_12445,N_8726);
xnor U15916 (N_15916,N_11405,N_9346);
nor U15917 (N_15917,N_11380,N_10887);
xor U15918 (N_15918,N_7944,N_6274);
nor U15919 (N_15919,N_8144,N_10026);
nor U15920 (N_15920,N_9961,N_12101);
and U15921 (N_15921,N_6273,N_9287);
nor U15922 (N_15922,N_8873,N_7718);
nor U15923 (N_15923,N_8143,N_11298);
nor U15924 (N_15924,N_9552,N_11706);
or U15925 (N_15925,N_11574,N_11718);
or U15926 (N_15926,N_9130,N_9994);
and U15927 (N_15927,N_11103,N_9339);
xnor U15928 (N_15928,N_7196,N_11157);
nand U15929 (N_15929,N_11275,N_7671);
nand U15930 (N_15930,N_11383,N_12450);
or U15931 (N_15931,N_10090,N_6340);
xor U15932 (N_15932,N_10318,N_12281);
nand U15933 (N_15933,N_7621,N_12179);
and U15934 (N_15934,N_7530,N_8858);
and U15935 (N_15935,N_7486,N_7264);
or U15936 (N_15936,N_8361,N_7209);
nand U15937 (N_15937,N_9836,N_8603);
xnor U15938 (N_15938,N_6714,N_12359);
nor U15939 (N_15939,N_10590,N_8900);
or U15940 (N_15940,N_6523,N_7430);
or U15941 (N_15941,N_10751,N_11259);
xor U15942 (N_15942,N_10035,N_11874);
or U15943 (N_15943,N_7618,N_11413);
nand U15944 (N_15944,N_7275,N_6864);
and U15945 (N_15945,N_11694,N_7623);
xor U15946 (N_15946,N_7155,N_9849);
or U15947 (N_15947,N_8320,N_9417);
nor U15948 (N_15948,N_11899,N_7105);
or U15949 (N_15949,N_8201,N_7736);
nand U15950 (N_15950,N_11772,N_10114);
nand U15951 (N_15951,N_11746,N_8655);
and U15952 (N_15952,N_8114,N_8082);
and U15953 (N_15953,N_7658,N_7420);
nor U15954 (N_15954,N_8249,N_7766);
nand U15955 (N_15955,N_10820,N_8962);
or U15956 (N_15956,N_12241,N_7284);
nor U15957 (N_15957,N_6947,N_9438);
nand U15958 (N_15958,N_10759,N_9083);
nand U15959 (N_15959,N_10764,N_10086);
nand U15960 (N_15960,N_6298,N_9394);
or U15961 (N_15961,N_6723,N_10311);
xnor U15962 (N_15962,N_8672,N_7353);
xor U15963 (N_15963,N_11483,N_11402);
nor U15964 (N_15964,N_10921,N_9895);
nor U15965 (N_15965,N_12313,N_12123);
nand U15966 (N_15966,N_10208,N_11979);
nor U15967 (N_15967,N_6531,N_9158);
or U15968 (N_15968,N_10699,N_12177);
or U15969 (N_15969,N_6450,N_11925);
and U15970 (N_15970,N_10709,N_9629);
nor U15971 (N_15971,N_10533,N_11577);
and U15972 (N_15972,N_9198,N_7120);
nor U15973 (N_15973,N_12085,N_10335);
nand U15974 (N_15974,N_10631,N_6794);
or U15975 (N_15975,N_7558,N_7418);
nor U15976 (N_15976,N_7791,N_9504);
nor U15977 (N_15977,N_12250,N_7952);
or U15978 (N_15978,N_7958,N_9975);
or U15979 (N_15979,N_8937,N_12184);
xor U15980 (N_15980,N_10201,N_6615);
or U15981 (N_15981,N_10572,N_11089);
and U15982 (N_15982,N_11793,N_7921);
nand U15983 (N_15983,N_10834,N_10385);
xor U15984 (N_15984,N_10726,N_9349);
nand U15985 (N_15985,N_11812,N_11572);
xor U15986 (N_15986,N_10318,N_6591);
or U15987 (N_15987,N_9984,N_10325);
or U15988 (N_15988,N_9601,N_11303);
nand U15989 (N_15989,N_9012,N_11728);
xnor U15990 (N_15990,N_12408,N_10395);
and U15991 (N_15991,N_8360,N_6543);
nand U15992 (N_15992,N_8574,N_6385);
nand U15993 (N_15993,N_8762,N_11561);
nor U15994 (N_15994,N_9403,N_7169);
nor U15995 (N_15995,N_9218,N_6924);
nor U15996 (N_15996,N_11003,N_6916);
xor U15997 (N_15997,N_7779,N_10008);
nor U15998 (N_15998,N_8246,N_11747);
and U15999 (N_15999,N_7780,N_9290);
and U16000 (N_16000,N_7771,N_9766);
and U16001 (N_16001,N_8467,N_7598);
xor U16002 (N_16002,N_8028,N_10055);
nor U16003 (N_16003,N_11006,N_9823);
and U16004 (N_16004,N_7007,N_11581);
or U16005 (N_16005,N_9717,N_11433);
and U16006 (N_16006,N_12432,N_11259);
xor U16007 (N_16007,N_7573,N_6849);
and U16008 (N_16008,N_12223,N_7651);
nand U16009 (N_16009,N_8625,N_6509);
and U16010 (N_16010,N_12446,N_10927);
and U16011 (N_16011,N_8770,N_11242);
or U16012 (N_16012,N_11933,N_6866);
nor U16013 (N_16013,N_9282,N_8370);
or U16014 (N_16014,N_6402,N_7760);
nand U16015 (N_16015,N_8965,N_8423);
nor U16016 (N_16016,N_9279,N_10520);
xor U16017 (N_16017,N_10572,N_8327);
nor U16018 (N_16018,N_6513,N_11180);
nand U16019 (N_16019,N_9239,N_12432);
nand U16020 (N_16020,N_9780,N_10539);
nor U16021 (N_16021,N_9942,N_12146);
nand U16022 (N_16022,N_9444,N_7618);
nand U16023 (N_16023,N_7268,N_9496);
nand U16024 (N_16024,N_8723,N_7045);
xnor U16025 (N_16025,N_11118,N_6978);
nand U16026 (N_16026,N_7094,N_7134);
and U16027 (N_16027,N_10928,N_12038);
and U16028 (N_16028,N_7797,N_10872);
xor U16029 (N_16029,N_8548,N_12139);
nand U16030 (N_16030,N_9962,N_11906);
or U16031 (N_16031,N_7679,N_6545);
nand U16032 (N_16032,N_6627,N_7869);
or U16033 (N_16033,N_9548,N_6934);
or U16034 (N_16034,N_11355,N_12474);
nand U16035 (N_16035,N_6591,N_12214);
nand U16036 (N_16036,N_10768,N_7579);
or U16037 (N_16037,N_6292,N_8299);
nand U16038 (N_16038,N_9410,N_8570);
nand U16039 (N_16039,N_10939,N_12311);
and U16040 (N_16040,N_9317,N_12069);
and U16041 (N_16041,N_8220,N_10862);
nor U16042 (N_16042,N_8521,N_8811);
or U16043 (N_16043,N_7829,N_10671);
and U16044 (N_16044,N_6378,N_12161);
or U16045 (N_16045,N_7679,N_9348);
xor U16046 (N_16046,N_10259,N_7103);
nand U16047 (N_16047,N_9810,N_6860);
nand U16048 (N_16048,N_12103,N_11249);
and U16049 (N_16049,N_8548,N_6911);
nor U16050 (N_16050,N_10420,N_7953);
or U16051 (N_16051,N_10901,N_6481);
nand U16052 (N_16052,N_9532,N_10714);
nand U16053 (N_16053,N_11918,N_9635);
nand U16054 (N_16054,N_12462,N_12100);
xnor U16055 (N_16055,N_7535,N_7141);
and U16056 (N_16056,N_6574,N_11192);
nor U16057 (N_16057,N_7240,N_7730);
nor U16058 (N_16058,N_8997,N_8917);
or U16059 (N_16059,N_10830,N_10629);
or U16060 (N_16060,N_9739,N_7265);
xor U16061 (N_16061,N_6915,N_11129);
or U16062 (N_16062,N_10000,N_10773);
nand U16063 (N_16063,N_11990,N_9905);
and U16064 (N_16064,N_9705,N_7413);
or U16065 (N_16065,N_8473,N_9325);
and U16066 (N_16066,N_11747,N_9594);
and U16067 (N_16067,N_7473,N_9348);
nand U16068 (N_16068,N_10449,N_8516);
and U16069 (N_16069,N_11101,N_6738);
and U16070 (N_16070,N_7106,N_11052);
and U16071 (N_16071,N_10195,N_12150);
nor U16072 (N_16072,N_7411,N_10107);
or U16073 (N_16073,N_7584,N_11876);
and U16074 (N_16074,N_11300,N_12260);
xnor U16075 (N_16075,N_9846,N_11495);
nor U16076 (N_16076,N_10233,N_7836);
or U16077 (N_16077,N_10088,N_7771);
and U16078 (N_16078,N_10218,N_10626);
or U16079 (N_16079,N_11005,N_9639);
and U16080 (N_16080,N_7205,N_11176);
and U16081 (N_16081,N_10790,N_6658);
or U16082 (N_16082,N_10710,N_11830);
or U16083 (N_16083,N_9546,N_8839);
nand U16084 (N_16084,N_7941,N_11614);
and U16085 (N_16085,N_7585,N_11043);
nand U16086 (N_16086,N_8072,N_7828);
nor U16087 (N_16087,N_10268,N_11638);
or U16088 (N_16088,N_10652,N_11647);
xnor U16089 (N_16089,N_12300,N_11692);
nor U16090 (N_16090,N_9440,N_7482);
nor U16091 (N_16091,N_9606,N_7571);
xnor U16092 (N_16092,N_6982,N_10860);
or U16093 (N_16093,N_11993,N_8565);
nor U16094 (N_16094,N_11665,N_7185);
and U16095 (N_16095,N_6519,N_7933);
nand U16096 (N_16096,N_6968,N_9878);
nand U16097 (N_16097,N_8871,N_8488);
and U16098 (N_16098,N_11281,N_11094);
xnor U16099 (N_16099,N_9914,N_11631);
or U16100 (N_16100,N_11144,N_11962);
nor U16101 (N_16101,N_10874,N_11485);
nor U16102 (N_16102,N_9269,N_8383);
and U16103 (N_16103,N_11251,N_11606);
nand U16104 (N_16104,N_6642,N_11627);
and U16105 (N_16105,N_10023,N_10981);
nand U16106 (N_16106,N_11732,N_11420);
nor U16107 (N_16107,N_6954,N_8485);
or U16108 (N_16108,N_8130,N_9958);
or U16109 (N_16109,N_7505,N_10526);
xor U16110 (N_16110,N_9281,N_7330);
nor U16111 (N_16111,N_8864,N_10915);
and U16112 (N_16112,N_10331,N_7546);
nand U16113 (N_16113,N_10742,N_11190);
and U16114 (N_16114,N_11748,N_9412);
xor U16115 (N_16115,N_7464,N_8538);
and U16116 (N_16116,N_11761,N_7393);
nor U16117 (N_16117,N_7524,N_9150);
nor U16118 (N_16118,N_8699,N_10323);
xor U16119 (N_16119,N_7038,N_10408);
nor U16120 (N_16120,N_8617,N_11672);
nand U16121 (N_16121,N_6452,N_9983);
nor U16122 (N_16122,N_8787,N_11189);
xnor U16123 (N_16123,N_10310,N_11487);
or U16124 (N_16124,N_11220,N_9892);
xor U16125 (N_16125,N_7886,N_7436);
nor U16126 (N_16126,N_6501,N_9802);
or U16127 (N_16127,N_6279,N_11734);
xnor U16128 (N_16128,N_8589,N_10770);
nand U16129 (N_16129,N_10614,N_8719);
nor U16130 (N_16130,N_10702,N_12127);
or U16131 (N_16131,N_8227,N_12287);
nor U16132 (N_16132,N_7589,N_6368);
xnor U16133 (N_16133,N_7200,N_7036);
and U16134 (N_16134,N_11111,N_8485);
nand U16135 (N_16135,N_10982,N_10167);
nand U16136 (N_16136,N_8244,N_7832);
nor U16137 (N_16137,N_9034,N_11054);
and U16138 (N_16138,N_7531,N_8445);
or U16139 (N_16139,N_9108,N_9063);
xnor U16140 (N_16140,N_10544,N_6558);
nor U16141 (N_16141,N_11634,N_6758);
xor U16142 (N_16142,N_9059,N_7364);
xnor U16143 (N_16143,N_9026,N_12145);
nor U16144 (N_16144,N_7153,N_11594);
nand U16145 (N_16145,N_8349,N_6924);
or U16146 (N_16146,N_10697,N_8258);
or U16147 (N_16147,N_6469,N_6917);
xor U16148 (N_16148,N_8074,N_10484);
nor U16149 (N_16149,N_9678,N_10922);
xor U16150 (N_16150,N_10201,N_7838);
xnor U16151 (N_16151,N_8710,N_8227);
nand U16152 (N_16152,N_10876,N_9158);
nand U16153 (N_16153,N_11159,N_10965);
nand U16154 (N_16154,N_7921,N_6424);
xor U16155 (N_16155,N_11915,N_9862);
nand U16156 (N_16156,N_8975,N_8672);
xor U16157 (N_16157,N_10338,N_8037);
xnor U16158 (N_16158,N_7034,N_9654);
and U16159 (N_16159,N_8689,N_12376);
nor U16160 (N_16160,N_11737,N_8980);
xor U16161 (N_16161,N_7571,N_10018);
or U16162 (N_16162,N_10628,N_6648);
nand U16163 (N_16163,N_9382,N_7147);
and U16164 (N_16164,N_10633,N_6806);
nand U16165 (N_16165,N_8885,N_10896);
and U16166 (N_16166,N_10299,N_9944);
xnor U16167 (N_16167,N_7968,N_9003);
nor U16168 (N_16168,N_9354,N_9335);
and U16169 (N_16169,N_12024,N_9443);
xnor U16170 (N_16170,N_8355,N_9376);
and U16171 (N_16171,N_9650,N_6403);
and U16172 (N_16172,N_10600,N_10347);
and U16173 (N_16173,N_10389,N_7792);
nand U16174 (N_16174,N_12445,N_9081);
nor U16175 (N_16175,N_8636,N_7216);
nor U16176 (N_16176,N_10371,N_8859);
nor U16177 (N_16177,N_11116,N_6943);
nor U16178 (N_16178,N_10688,N_8620);
and U16179 (N_16179,N_9097,N_9141);
and U16180 (N_16180,N_11119,N_12446);
nand U16181 (N_16181,N_7460,N_7718);
or U16182 (N_16182,N_10837,N_9448);
xnor U16183 (N_16183,N_8297,N_12331);
xor U16184 (N_16184,N_9520,N_6375);
nand U16185 (N_16185,N_9219,N_9018);
nor U16186 (N_16186,N_8631,N_9050);
and U16187 (N_16187,N_12252,N_7042);
or U16188 (N_16188,N_7102,N_9518);
or U16189 (N_16189,N_7569,N_11099);
nor U16190 (N_16190,N_12492,N_10039);
nor U16191 (N_16191,N_11889,N_7795);
nand U16192 (N_16192,N_8524,N_7802);
xor U16193 (N_16193,N_7923,N_12064);
or U16194 (N_16194,N_6988,N_10151);
nor U16195 (N_16195,N_8764,N_9623);
and U16196 (N_16196,N_10569,N_10239);
nor U16197 (N_16197,N_7036,N_7196);
and U16198 (N_16198,N_12194,N_9202);
nor U16199 (N_16199,N_8920,N_11589);
nand U16200 (N_16200,N_10979,N_6416);
nand U16201 (N_16201,N_10250,N_10678);
xor U16202 (N_16202,N_11167,N_7141);
and U16203 (N_16203,N_11898,N_7587);
and U16204 (N_16204,N_8230,N_10789);
nand U16205 (N_16205,N_7373,N_11485);
nand U16206 (N_16206,N_10708,N_12217);
xnor U16207 (N_16207,N_9815,N_6938);
and U16208 (N_16208,N_12048,N_10867);
or U16209 (N_16209,N_12494,N_6628);
nor U16210 (N_16210,N_7349,N_9652);
or U16211 (N_16211,N_8743,N_10933);
nor U16212 (N_16212,N_11570,N_7747);
or U16213 (N_16213,N_6846,N_10837);
and U16214 (N_16214,N_7842,N_6768);
nand U16215 (N_16215,N_9094,N_9208);
nand U16216 (N_16216,N_10294,N_10526);
xor U16217 (N_16217,N_6847,N_8609);
or U16218 (N_16218,N_6967,N_12321);
and U16219 (N_16219,N_9516,N_9566);
xnor U16220 (N_16220,N_11683,N_11424);
nand U16221 (N_16221,N_10786,N_11838);
nor U16222 (N_16222,N_7598,N_11091);
xnor U16223 (N_16223,N_9574,N_12244);
and U16224 (N_16224,N_11397,N_10800);
xnor U16225 (N_16225,N_9214,N_9964);
or U16226 (N_16226,N_8029,N_9981);
and U16227 (N_16227,N_9172,N_11858);
xor U16228 (N_16228,N_7962,N_8290);
and U16229 (N_16229,N_10040,N_11593);
xnor U16230 (N_16230,N_8150,N_10132);
or U16231 (N_16231,N_11647,N_8536);
and U16232 (N_16232,N_11624,N_12287);
xor U16233 (N_16233,N_9638,N_8848);
nor U16234 (N_16234,N_7994,N_9768);
or U16235 (N_16235,N_6904,N_9518);
nand U16236 (N_16236,N_9904,N_8963);
or U16237 (N_16237,N_10943,N_9257);
or U16238 (N_16238,N_11257,N_6918);
or U16239 (N_16239,N_6847,N_11011);
and U16240 (N_16240,N_11234,N_10400);
nand U16241 (N_16241,N_10982,N_9803);
and U16242 (N_16242,N_10002,N_8973);
and U16243 (N_16243,N_7674,N_8102);
nor U16244 (N_16244,N_6802,N_11299);
or U16245 (N_16245,N_11227,N_9956);
or U16246 (N_16246,N_11644,N_6528);
xor U16247 (N_16247,N_10896,N_8961);
nor U16248 (N_16248,N_11506,N_10317);
and U16249 (N_16249,N_8894,N_11015);
and U16250 (N_16250,N_10811,N_6252);
nor U16251 (N_16251,N_6807,N_10797);
nor U16252 (N_16252,N_10968,N_12087);
and U16253 (N_16253,N_6258,N_10468);
nand U16254 (N_16254,N_8618,N_8655);
nor U16255 (N_16255,N_8420,N_12284);
or U16256 (N_16256,N_9462,N_10404);
nor U16257 (N_16257,N_9223,N_9997);
nor U16258 (N_16258,N_10659,N_11355);
xnor U16259 (N_16259,N_6739,N_12320);
xor U16260 (N_16260,N_7424,N_6859);
and U16261 (N_16261,N_11213,N_11712);
or U16262 (N_16262,N_6442,N_11682);
xor U16263 (N_16263,N_12026,N_8890);
and U16264 (N_16264,N_8289,N_10795);
and U16265 (N_16265,N_8640,N_7001);
nand U16266 (N_16266,N_12426,N_7472);
xnor U16267 (N_16267,N_6343,N_6757);
nand U16268 (N_16268,N_8681,N_11874);
xor U16269 (N_16269,N_6494,N_11378);
and U16270 (N_16270,N_6481,N_7544);
nand U16271 (N_16271,N_9988,N_6421);
or U16272 (N_16272,N_11842,N_7796);
and U16273 (N_16273,N_7356,N_8854);
nor U16274 (N_16274,N_12460,N_11857);
xor U16275 (N_16275,N_10069,N_10408);
xor U16276 (N_16276,N_6719,N_7007);
nor U16277 (N_16277,N_6622,N_7650);
or U16278 (N_16278,N_7322,N_10753);
nand U16279 (N_16279,N_7032,N_9409);
nor U16280 (N_16280,N_7659,N_8496);
nand U16281 (N_16281,N_12357,N_9061);
xor U16282 (N_16282,N_9414,N_11210);
and U16283 (N_16283,N_6748,N_7902);
or U16284 (N_16284,N_11075,N_8971);
or U16285 (N_16285,N_8008,N_11087);
xnor U16286 (N_16286,N_11552,N_9581);
or U16287 (N_16287,N_7013,N_9549);
and U16288 (N_16288,N_8294,N_7560);
nor U16289 (N_16289,N_11089,N_10190);
nand U16290 (N_16290,N_9417,N_7420);
nand U16291 (N_16291,N_6714,N_7887);
nand U16292 (N_16292,N_11904,N_8033);
xor U16293 (N_16293,N_8807,N_10423);
xnor U16294 (N_16294,N_7198,N_8974);
xnor U16295 (N_16295,N_9070,N_7221);
xnor U16296 (N_16296,N_11262,N_9417);
nor U16297 (N_16297,N_6674,N_11681);
nor U16298 (N_16298,N_6425,N_9195);
nor U16299 (N_16299,N_6267,N_12043);
or U16300 (N_16300,N_7888,N_8313);
or U16301 (N_16301,N_11442,N_9763);
or U16302 (N_16302,N_11732,N_7139);
xnor U16303 (N_16303,N_10580,N_8859);
nand U16304 (N_16304,N_7892,N_10744);
nor U16305 (N_16305,N_10795,N_8733);
and U16306 (N_16306,N_9425,N_12488);
and U16307 (N_16307,N_9817,N_8125);
or U16308 (N_16308,N_7318,N_12417);
and U16309 (N_16309,N_8433,N_9132);
and U16310 (N_16310,N_6561,N_10017);
xnor U16311 (N_16311,N_8287,N_7817);
nor U16312 (N_16312,N_9475,N_6349);
nand U16313 (N_16313,N_6723,N_8479);
nor U16314 (N_16314,N_10882,N_6626);
nand U16315 (N_16315,N_12158,N_7482);
nand U16316 (N_16316,N_8655,N_11310);
nor U16317 (N_16317,N_9458,N_11802);
and U16318 (N_16318,N_11824,N_11959);
nand U16319 (N_16319,N_11129,N_7032);
or U16320 (N_16320,N_8439,N_9820);
xor U16321 (N_16321,N_8919,N_8254);
nand U16322 (N_16322,N_8955,N_10202);
nor U16323 (N_16323,N_12251,N_12131);
nand U16324 (N_16324,N_8793,N_11395);
or U16325 (N_16325,N_11750,N_7606);
nor U16326 (N_16326,N_10358,N_11728);
nor U16327 (N_16327,N_8807,N_6984);
and U16328 (N_16328,N_8858,N_12107);
or U16329 (N_16329,N_9341,N_6815);
xnor U16330 (N_16330,N_10504,N_9954);
nand U16331 (N_16331,N_9788,N_9341);
xor U16332 (N_16332,N_7308,N_7965);
nand U16333 (N_16333,N_12483,N_11495);
nand U16334 (N_16334,N_8226,N_7928);
and U16335 (N_16335,N_7944,N_10018);
or U16336 (N_16336,N_6408,N_7657);
nand U16337 (N_16337,N_10060,N_11106);
and U16338 (N_16338,N_11723,N_8704);
nor U16339 (N_16339,N_8575,N_9051);
nor U16340 (N_16340,N_9566,N_6492);
nor U16341 (N_16341,N_9510,N_6962);
nor U16342 (N_16342,N_10475,N_8693);
nand U16343 (N_16343,N_9564,N_6560);
and U16344 (N_16344,N_12217,N_11681);
nand U16345 (N_16345,N_12187,N_11288);
nand U16346 (N_16346,N_8146,N_10332);
xnor U16347 (N_16347,N_8384,N_12168);
and U16348 (N_16348,N_6378,N_11527);
and U16349 (N_16349,N_12146,N_9545);
nand U16350 (N_16350,N_9069,N_6827);
nand U16351 (N_16351,N_9719,N_10532);
nor U16352 (N_16352,N_8685,N_10202);
and U16353 (N_16353,N_7058,N_9468);
nor U16354 (N_16354,N_7640,N_9060);
xor U16355 (N_16355,N_12133,N_11381);
and U16356 (N_16356,N_7429,N_11363);
xor U16357 (N_16357,N_9423,N_12276);
and U16358 (N_16358,N_9287,N_9526);
nor U16359 (N_16359,N_11886,N_10040);
and U16360 (N_16360,N_6737,N_7325);
or U16361 (N_16361,N_12371,N_10542);
xnor U16362 (N_16362,N_8333,N_9656);
nor U16363 (N_16363,N_6558,N_6723);
xnor U16364 (N_16364,N_11178,N_8710);
xor U16365 (N_16365,N_11910,N_10437);
nand U16366 (N_16366,N_8472,N_7923);
and U16367 (N_16367,N_10642,N_8534);
and U16368 (N_16368,N_6936,N_11653);
xor U16369 (N_16369,N_9757,N_7284);
nand U16370 (N_16370,N_9618,N_11657);
or U16371 (N_16371,N_12105,N_8352);
xor U16372 (N_16372,N_10494,N_6573);
xor U16373 (N_16373,N_10050,N_11611);
or U16374 (N_16374,N_6276,N_10399);
and U16375 (N_16375,N_6471,N_10092);
or U16376 (N_16376,N_9533,N_11823);
nand U16377 (N_16377,N_9775,N_10696);
nor U16378 (N_16378,N_9220,N_6967);
nor U16379 (N_16379,N_8438,N_6873);
and U16380 (N_16380,N_10453,N_6301);
nand U16381 (N_16381,N_10947,N_7559);
nor U16382 (N_16382,N_6511,N_6678);
or U16383 (N_16383,N_7395,N_8160);
and U16384 (N_16384,N_9318,N_9201);
or U16385 (N_16385,N_12034,N_8716);
nand U16386 (N_16386,N_10827,N_10796);
nor U16387 (N_16387,N_10613,N_9393);
nor U16388 (N_16388,N_7027,N_7548);
or U16389 (N_16389,N_8045,N_7059);
nor U16390 (N_16390,N_9301,N_7060);
xor U16391 (N_16391,N_9105,N_10500);
xor U16392 (N_16392,N_9906,N_10102);
xnor U16393 (N_16393,N_10521,N_7823);
nor U16394 (N_16394,N_9150,N_8648);
xor U16395 (N_16395,N_9453,N_7285);
nor U16396 (N_16396,N_11456,N_8475);
nand U16397 (N_16397,N_11876,N_7916);
nand U16398 (N_16398,N_10665,N_9887);
nand U16399 (N_16399,N_9234,N_10060);
xnor U16400 (N_16400,N_7128,N_11091);
nor U16401 (N_16401,N_12262,N_7936);
nand U16402 (N_16402,N_11140,N_10991);
nor U16403 (N_16403,N_9084,N_8179);
or U16404 (N_16404,N_12411,N_11755);
xnor U16405 (N_16405,N_6571,N_12375);
nor U16406 (N_16406,N_7550,N_10508);
nor U16407 (N_16407,N_8804,N_8482);
and U16408 (N_16408,N_10133,N_12412);
xor U16409 (N_16409,N_7111,N_12213);
nor U16410 (N_16410,N_6313,N_10015);
nand U16411 (N_16411,N_8784,N_12343);
nor U16412 (N_16412,N_11299,N_10847);
and U16413 (N_16413,N_7807,N_12483);
or U16414 (N_16414,N_9691,N_12389);
and U16415 (N_16415,N_11671,N_9462);
nand U16416 (N_16416,N_11838,N_10887);
xnor U16417 (N_16417,N_7523,N_9039);
or U16418 (N_16418,N_9334,N_8474);
nor U16419 (N_16419,N_9625,N_8018);
nand U16420 (N_16420,N_7946,N_10313);
and U16421 (N_16421,N_11963,N_9533);
xnor U16422 (N_16422,N_9905,N_8918);
xnor U16423 (N_16423,N_7521,N_12077);
nand U16424 (N_16424,N_8947,N_10663);
nand U16425 (N_16425,N_9866,N_7935);
or U16426 (N_16426,N_6765,N_10440);
nand U16427 (N_16427,N_11654,N_11956);
or U16428 (N_16428,N_7420,N_11733);
or U16429 (N_16429,N_7301,N_11679);
nor U16430 (N_16430,N_6869,N_9059);
xor U16431 (N_16431,N_11513,N_7280);
nor U16432 (N_16432,N_10972,N_6504);
or U16433 (N_16433,N_10193,N_9756);
xor U16434 (N_16434,N_8442,N_10314);
nor U16435 (N_16435,N_11489,N_8709);
and U16436 (N_16436,N_8698,N_6614);
xnor U16437 (N_16437,N_9275,N_10378);
nand U16438 (N_16438,N_8691,N_9768);
or U16439 (N_16439,N_12039,N_9395);
nor U16440 (N_16440,N_10132,N_11550);
and U16441 (N_16441,N_9338,N_6380);
nor U16442 (N_16442,N_8919,N_10659);
xor U16443 (N_16443,N_8339,N_6562);
or U16444 (N_16444,N_11418,N_10254);
or U16445 (N_16445,N_6294,N_7145);
or U16446 (N_16446,N_7179,N_6477);
or U16447 (N_16447,N_10599,N_12439);
or U16448 (N_16448,N_8316,N_9299);
nand U16449 (N_16449,N_9885,N_9334);
nand U16450 (N_16450,N_11732,N_12338);
or U16451 (N_16451,N_10434,N_8488);
nand U16452 (N_16452,N_11090,N_10300);
nor U16453 (N_16453,N_10406,N_6480);
and U16454 (N_16454,N_12438,N_10111);
and U16455 (N_16455,N_12190,N_11609);
xnor U16456 (N_16456,N_9880,N_7887);
nor U16457 (N_16457,N_12356,N_10155);
or U16458 (N_16458,N_9203,N_10355);
and U16459 (N_16459,N_7218,N_6387);
nor U16460 (N_16460,N_10784,N_11873);
nand U16461 (N_16461,N_10352,N_8188);
nand U16462 (N_16462,N_7609,N_11657);
nor U16463 (N_16463,N_8770,N_6872);
and U16464 (N_16464,N_11474,N_9346);
or U16465 (N_16465,N_7367,N_7116);
nor U16466 (N_16466,N_9239,N_9063);
nand U16467 (N_16467,N_10834,N_8896);
or U16468 (N_16468,N_8634,N_11039);
and U16469 (N_16469,N_10346,N_10321);
nor U16470 (N_16470,N_8416,N_7293);
and U16471 (N_16471,N_7024,N_9234);
and U16472 (N_16472,N_9088,N_10961);
xor U16473 (N_16473,N_8893,N_8815);
nand U16474 (N_16474,N_6453,N_8424);
nand U16475 (N_16475,N_7832,N_10343);
xnor U16476 (N_16476,N_8105,N_12263);
nand U16477 (N_16477,N_7494,N_7272);
or U16478 (N_16478,N_7794,N_12000);
or U16479 (N_16479,N_12262,N_7040);
or U16480 (N_16480,N_11473,N_7076);
or U16481 (N_16481,N_7879,N_7843);
or U16482 (N_16482,N_7708,N_6946);
and U16483 (N_16483,N_7147,N_10304);
or U16484 (N_16484,N_9301,N_10757);
and U16485 (N_16485,N_7411,N_7315);
xor U16486 (N_16486,N_11927,N_8083);
and U16487 (N_16487,N_9402,N_8395);
nor U16488 (N_16488,N_7294,N_8040);
nand U16489 (N_16489,N_9103,N_11432);
xnor U16490 (N_16490,N_11412,N_11200);
and U16491 (N_16491,N_8758,N_10741);
nand U16492 (N_16492,N_9356,N_9413);
nand U16493 (N_16493,N_9820,N_11893);
nand U16494 (N_16494,N_12042,N_10109);
nand U16495 (N_16495,N_10643,N_8833);
nand U16496 (N_16496,N_7910,N_6717);
xor U16497 (N_16497,N_11595,N_7964);
and U16498 (N_16498,N_11610,N_9074);
nor U16499 (N_16499,N_11606,N_7078);
or U16500 (N_16500,N_9899,N_10688);
nand U16501 (N_16501,N_10928,N_11489);
or U16502 (N_16502,N_8803,N_8888);
xor U16503 (N_16503,N_6921,N_12310);
and U16504 (N_16504,N_11299,N_12015);
xnor U16505 (N_16505,N_9405,N_7781);
and U16506 (N_16506,N_12227,N_6252);
nor U16507 (N_16507,N_6752,N_12376);
and U16508 (N_16508,N_10909,N_7837);
nor U16509 (N_16509,N_12165,N_9453);
nor U16510 (N_16510,N_8010,N_7527);
nor U16511 (N_16511,N_10894,N_9752);
or U16512 (N_16512,N_9657,N_9538);
nor U16513 (N_16513,N_10011,N_7197);
nor U16514 (N_16514,N_7718,N_7006);
and U16515 (N_16515,N_11986,N_11028);
and U16516 (N_16516,N_7197,N_10676);
or U16517 (N_16517,N_10982,N_7381);
nor U16518 (N_16518,N_9930,N_7727);
nand U16519 (N_16519,N_10482,N_10997);
nand U16520 (N_16520,N_7900,N_9976);
nor U16521 (N_16521,N_7804,N_11249);
xnor U16522 (N_16522,N_10736,N_11587);
and U16523 (N_16523,N_6955,N_8411);
nand U16524 (N_16524,N_10332,N_10956);
or U16525 (N_16525,N_10385,N_7345);
or U16526 (N_16526,N_12065,N_7495);
or U16527 (N_16527,N_8992,N_8120);
nor U16528 (N_16528,N_10791,N_7485);
nand U16529 (N_16529,N_9639,N_9116);
nand U16530 (N_16530,N_11442,N_11202);
nand U16531 (N_16531,N_8521,N_9667);
or U16532 (N_16532,N_6642,N_6718);
xor U16533 (N_16533,N_8341,N_12019);
nor U16534 (N_16534,N_8335,N_8097);
xnor U16535 (N_16535,N_10735,N_10237);
or U16536 (N_16536,N_6956,N_10133);
xnor U16537 (N_16537,N_8368,N_10344);
or U16538 (N_16538,N_7156,N_8117);
or U16539 (N_16539,N_6807,N_11831);
xnor U16540 (N_16540,N_7891,N_9453);
nand U16541 (N_16541,N_12247,N_10272);
xnor U16542 (N_16542,N_10065,N_9907);
nand U16543 (N_16543,N_8497,N_12074);
nand U16544 (N_16544,N_9682,N_11046);
nand U16545 (N_16545,N_12278,N_11574);
nand U16546 (N_16546,N_8936,N_9555);
nor U16547 (N_16547,N_10530,N_8057);
nand U16548 (N_16548,N_6932,N_8631);
nand U16549 (N_16549,N_12332,N_7444);
nor U16550 (N_16550,N_11894,N_10907);
or U16551 (N_16551,N_12386,N_8611);
nor U16552 (N_16552,N_10053,N_10126);
xnor U16553 (N_16553,N_11724,N_7826);
nand U16554 (N_16554,N_12188,N_12287);
nand U16555 (N_16555,N_6429,N_9137);
nand U16556 (N_16556,N_7792,N_9075);
or U16557 (N_16557,N_6424,N_10077);
xnor U16558 (N_16558,N_11898,N_7924);
and U16559 (N_16559,N_7842,N_9077);
xor U16560 (N_16560,N_8213,N_11185);
or U16561 (N_16561,N_8039,N_7416);
nand U16562 (N_16562,N_9741,N_6875);
and U16563 (N_16563,N_11954,N_10701);
nand U16564 (N_16564,N_7972,N_8257);
nand U16565 (N_16565,N_9542,N_6413);
and U16566 (N_16566,N_9892,N_11490);
or U16567 (N_16567,N_9792,N_10121);
and U16568 (N_16568,N_12096,N_7776);
xnor U16569 (N_16569,N_9620,N_7450);
nor U16570 (N_16570,N_9581,N_7649);
nand U16571 (N_16571,N_12200,N_10889);
xnor U16572 (N_16572,N_7696,N_10302);
nor U16573 (N_16573,N_11775,N_8193);
nand U16574 (N_16574,N_7213,N_12201);
or U16575 (N_16575,N_12396,N_10326);
and U16576 (N_16576,N_10660,N_12274);
nor U16577 (N_16577,N_11981,N_10273);
nor U16578 (N_16578,N_6913,N_8006);
and U16579 (N_16579,N_6959,N_7516);
nand U16580 (N_16580,N_8363,N_9695);
nor U16581 (N_16581,N_7685,N_7063);
or U16582 (N_16582,N_7152,N_11094);
and U16583 (N_16583,N_6369,N_8770);
or U16584 (N_16584,N_8137,N_7988);
and U16585 (N_16585,N_8465,N_11658);
nor U16586 (N_16586,N_10970,N_11170);
or U16587 (N_16587,N_10041,N_10461);
nand U16588 (N_16588,N_8439,N_11858);
xnor U16589 (N_16589,N_7461,N_6938);
nand U16590 (N_16590,N_9056,N_11275);
nand U16591 (N_16591,N_11267,N_7103);
nand U16592 (N_16592,N_9767,N_7931);
and U16593 (N_16593,N_7613,N_9398);
nor U16594 (N_16594,N_7513,N_11087);
xnor U16595 (N_16595,N_11358,N_10179);
and U16596 (N_16596,N_8577,N_9701);
nor U16597 (N_16597,N_9163,N_8040);
and U16598 (N_16598,N_6658,N_12171);
nand U16599 (N_16599,N_8632,N_9607);
or U16600 (N_16600,N_11358,N_6866);
xor U16601 (N_16601,N_10213,N_7258);
nand U16602 (N_16602,N_8514,N_11043);
xnor U16603 (N_16603,N_8113,N_6843);
xnor U16604 (N_16604,N_10688,N_9867);
or U16605 (N_16605,N_12234,N_8702);
nand U16606 (N_16606,N_7608,N_7227);
and U16607 (N_16607,N_10746,N_10889);
or U16608 (N_16608,N_10288,N_8473);
xor U16609 (N_16609,N_6811,N_11331);
or U16610 (N_16610,N_8697,N_12281);
or U16611 (N_16611,N_8806,N_8369);
nor U16612 (N_16612,N_7190,N_11686);
nor U16613 (N_16613,N_7972,N_9905);
nor U16614 (N_16614,N_8705,N_6426);
nor U16615 (N_16615,N_9473,N_7522);
and U16616 (N_16616,N_9886,N_10156);
and U16617 (N_16617,N_11948,N_11989);
nand U16618 (N_16618,N_11552,N_9853);
nor U16619 (N_16619,N_6650,N_8225);
xnor U16620 (N_16620,N_6497,N_11222);
nor U16621 (N_16621,N_11365,N_7910);
nor U16622 (N_16622,N_6299,N_7856);
xor U16623 (N_16623,N_11966,N_11090);
nor U16624 (N_16624,N_11983,N_10130);
and U16625 (N_16625,N_9073,N_10994);
or U16626 (N_16626,N_9105,N_10633);
xor U16627 (N_16627,N_7315,N_10190);
xor U16628 (N_16628,N_10888,N_11696);
or U16629 (N_16629,N_8857,N_6750);
xnor U16630 (N_16630,N_11640,N_7694);
nand U16631 (N_16631,N_7521,N_7421);
and U16632 (N_16632,N_10573,N_11546);
nor U16633 (N_16633,N_9104,N_6647);
nand U16634 (N_16634,N_10903,N_11115);
nand U16635 (N_16635,N_11875,N_8664);
and U16636 (N_16636,N_11236,N_10238);
nor U16637 (N_16637,N_6957,N_11130);
nand U16638 (N_16638,N_11585,N_6293);
xnor U16639 (N_16639,N_10574,N_8790);
nand U16640 (N_16640,N_12218,N_7944);
nor U16641 (N_16641,N_9626,N_7739);
nor U16642 (N_16642,N_8121,N_10577);
and U16643 (N_16643,N_9305,N_7744);
or U16644 (N_16644,N_9340,N_8634);
and U16645 (N_16645,N_6812,N_6783);
or U16646 (N_16646,N_8658,N_7308);
xor U16647 (N_16647,N_11123,N_6640);
nand U16648 (N_16648,N_8236,N_10646);
xnor U16649 (N_16649,N_11904,N_10641);
or U16650 (N_16650,N_6536,N_8019);
nor U16651 (N_16651,N_11699,N_9088);
nor U16652 (N_16652,N_7954,N_9133);
nand U16653 (N_16653,N_6658,N_9937);
nand U16654 (N_16654,N_11386,N_7742);
nand U16655 (N_16655,N_12039,N_6296);
or U16656 (N_16656,N_10673,N_11407);
xor U16657 (N_16657,N_10611,N_11961);
xnor U16658 (N_16658,N_11847,N_12350);
nand U16659 (N_16659,N_10087,N_7097);
and U16660 (N_16660,N_8406,N_9580);
or U16661 (N_16661,N_11839,N_8200);
and U16662 (N_16662,N_10588,N_6607);
or U16663 (N_16663,N_9383,N_12146);
or U16664 (N_16664,N_7006,N_10188);
xor U16665 (N_16665,N_8514,N_12283);
nor U16666 (N_16666,N_7637,N_6593);
or U16667 (N_16667,N_7488,N_7138);
nor U16668 (N_16668,N_7130,N_6934);
nor U16669 (N_16669,N_12409,N_9962);
xor U16670 (N_16670,N_10062,N_8131);
nor U16671 (N_16671,N_7463,N_11392);
nor U16672 (N_16672,N_9788,N_9039);
nand U16673 (N_16673,N_9945,N_7739);
nand U16674 (N_16674,N_7794,N_8933);
or U16675 (N_16675,N_11837,N_7524);
or U16676 (N_16676,N_7745,N_11454);
and U16677 (N_16677,N_12190,N_9858);
nor U16678 (N_16678,N_9881,N_7280);
xor U16679 (N_16679,N_7020,N_8557);
nand U16680 (N_16680,N_11816,N_9391);
or U16681 (N_16681,N_12311,N_7741);
nor U16682 (N_16682,N_12329,N_6511);
nor U16683 (N_16683,N_6856,N_10258);
nand U16684 (N_16684,N_9906,N_6507);
and U16685 (N_16685,N_7742,N_9635);
and U16686 (N_16686,N_8102,N_8938);
nor U16687 (N_16687,N_8780,N_10192);
and U16688 (N_16688,N_6300,N_11921);
nand U16689 (N_16689,N_9673,N_9570);
and U16690 (N_16690,N_6717,N_9692);
and U16691 (N_16691,N_12008,N_11767);
nor U16692 (N_16692,N_12332,N_7722);
nor U16693 (N_16693,N_6527,N_7291);
or U16694 (N_16694,N_7817,N_11802);
xnor U16695 (N_16695,N_10678,N_9058);
nand U16696 (N_16696,N_10379,N_6849);
and U16697 (N_16697,N_10376,N_11216);
nor U16698 (N_16698,N_7704,N_7090);
or U16699 (N_16699,N_10495,N_9735);
and U16700 (N_16700,N_6956,N_7037);
xor U16701 (N_16701,N_8460,N_9662);
nand U16702 (N_16702,N_12116,N_12361);
xnor U16703 (N_16703,N_6469,N_7782);
xor U16704 (N_16704,N_7015,N_11066);
or U16705 (N_16705,N_7633,N_7556);
nor U16706 (N_16706,N_7157,N_7426);
nand U16707 (N_16707,N_8334,N_8889);
nand U16708 (N_16708,N_7678,N_12473);
and U16709 (N_16709,N_8425,N_9411);
nor U16710 (N_16710,N_9116,N_9393);
or U16711 (N_16711,N_8695,N_9255);
and U16712 (N_16712,N_9092,N_8592);
nor U16713 (N_16713,N_6730,N_12034);
nor U16714 (N_16714,N_8017,N_10175);
nand U16715 (N_16715,N_7725,N_10006);
xor U16716 (N_16716,N_6647,N_9864);
xor U16717 (N_16717,N_9036,N_10885);
and U16718 (N_16718,N_7917,N_10908);
nor U16719 (N_16719,N_7948,N_10187);
or U16720 (N_16720,N_11974,N_12173);
and U16721 (N_16721,N_7545,N_10252);
nand U16722 (N_16722,N_10345,N_12281);
xor U16723 (N_16723,N_9858,N_8419);
nand U16724 (N_16724,N_11424,N_12219);
nor U16725 (N_16725,N_11095,N_10403);
nor U16726 (N_16726,N_12353,N_8944);
or U16727 (N_16727,N_11157,N_6833);
and U16728 (N_16728,N_8065,N_11351);
or U16729 (N_16729,N_11336,N_9476);
nand U16730 (N_16730,N_7446,N_12345);
and U16731 (N_16731,N_9440,N_9704);
nor U16732 (N_16732,N_7202,N_8784);
nand U16733 (N_16733,N_6708,N_10442);
nand U16734 (N_16734,N_9143,N_11950);
nand U16735 (N_16735,N_9881,N_11129);
nor U16736 (N_16736,N_11686,N_6547);
or U16737 (N_16737,N_10266,N_6981);
xnor U16738 (N_16738,N_8573,N_7049);
and U16739 (N_16739,N_10417,N_8759);
nand U16740 (N_16740,N_8054,N_10122);
nand U16741 (N_16741,N_10727,N_11458);
and U16742 (N_16742,N_6286,N_7901);
nor U16743 (N_16743,N_11853,N_9386);
xor U16744 (N_16744,N_12115,N_8904);
nor U16745 (N_16745,N_11084,N_9253);
or U16746 (N_16746,N_9074,N_6631);
or U16747 (N_16747,N_8223,N_11697);
or U16748 (N_16748,N_7569,N_10582);
or U16749 (N_16749,N_8647,N_12313);
nand U16750 (N_16750,N_9949,N_11579);
or U16751 (N_16751,N_12075,N_8185);
xnor U16752 (N_16752,N_12047,N_10505);
and U16753 (N_16753,N_7161,N_6854);
and U16754 (N_16754,N_10425,N_10501);
nor U16755 (N_16755,N_9994,N_7128);
nor U16756 (N_16756,N_9689,N_7783);
nand U16757 (N_16757,N_6331,N_6676);
or U16758 (N_16758,N_10218,N_8871);
nor U16759 (N_16759,N_11060,N_8440);
nor U16760 (N_16760,N_12482,N_6415);
or U16761 (N_16761,N_7373,N_7519);
or U16762 (N_16762,N_10160,N_10243);
or U16763 (N_16763,N_8991,N_7978);
nand U16764 (N_16764,N_8514,N_8539);
xor U16765 (N_16765,N_11162,N_11327);
nor U16766 (N_16766,N_9678,N_8734);
xor U16767 (N_16767,N_8667,N_7426);
nand U16768 (N_16768,N_7444,N_8588);
nand U16769 (N_16769,N_11005,N_8739);
nand U16770 (N_16770,N_10877,N_8382);
xor U16771 (N_16771,N_7593,N_8647);
and U16772 (N_16772,N_9140,N_6382);
and U16773 (N_16773,N_10237,N_7424);
or U16774 (N_16774,N_6820,N_8028);
or U16775 (N_16775,N_8981,N_10093);
and U16776 (N_16776,N_10905,N_11905);
nor U16777 (N_16777,N_7670,N_11325);
nor U16778 (N_16778,N_12131,N_6265);
or U16779 (N_16779,N_11827,N_7346);
or U16780 (N_16780,N_10664,N_7116);
nor U16781 (N_16781,N_11680,N_12180);
nor U16782 (N_16782,N_11088,N_7706);
xor U16783 (N_16783,N_11852,N_12078);
xor U16784 (N_16784,N_9744,N_11134);
nor U16785 (N_16785,N_8998,N_7387);
xnor U16786 (N_16786,N_8901,N_10341);
or U16787 (N_16787,N_11693,N_8799);
nand U16788 (N_16788,N_12028,N_7968);
or U16789 (N_16789,N_9812,N_11714);
xor U16790 (N_16790,N_8975,N_8373);
nand U16791 (N_16791,N_11944,N_11491);
nand U16792 (N_16792,N_8801,N_12194);
and U16793 (N_16793,N_9977,N_8102);
nand U16794 (N_16794,N_9576,N_7575);
and U16795 (N_16795,N_9702,N_10562);
or U16796 (N_16796,N_12046,N_8208);
or U16797 (N_16797,N_9379,N_9868);
nor U16798 (N_16798,N_7551,N_9899);
nor U16799 (N_16799,N_8651,N_11702);
and U16800 (N_16800,N_8981,N_8824);
nor U16801 (N_16801,N_8761,N_8308);
nand U16802 (N_16802,N_9119,N_7841);
xnor U16803 (N_16803,N_11309,N_10211);
and U16804 (N_16804,N_8192,N_10721);
nor U16805 (N_16805,N_7789,N_10137);
and U16806 (N_16806,N_10779,N_9586);
xor U16807 (N_16807,N_9790,N_8897);
nor U16808 (N_16808,N_7053,N_11263);
nand U16809 (N_16809,N_12407,N_7561);
or U16810 (N_16810,N_7989,N_6710);
nor U16811 (N_16811,N_8595,N_11499);
and U16812 (N_16812,N_9735,N_9171);
and U16813 (N_16813,N_10200,N_11471);
nand U16814 (N_16814,N_8676,N_12167);
nand U16815 (N_16815,N_8568,N_11714);
and U16816 (N_16816,N_11531,N_11172);
or U16817 (N_16817,N_10282,N_7475);
xor U16818 (N_16818,N_8577,N_9512);
or U16819 (N_16819,N_8057,N_9051);
or U16820 (N_16820,N_7785,N_6933);
and U16821 (N_16821,N_10271,N_11235);
xor U16822 (N_16822,N_6935,N_7260);
and U16823 (N_16823,N_11276,N_8244);
or U16824 (N_16824,N_9089,N_12346);
xor U16825 (N_16825,N_8887,N_8490);
or U16826 (N_16826,N_10190,N_8443);
and U16827 (N_16827,N_11221,N_8436);
and U16828 (N_16828,N_11080,N_7835);
or U16829 (N_16829,N_10173,N_11347);
nor U16830 (N_16830,N_6767,N_10345);
or U16831 (N_16831,N_12484,N_10383);
or U16832 (N_16832,N_9468,N_8209);
and U16833 (N_16833,N_6590,N_9804);
nand U16834 (N_16834,N_10574,N_9051);
or U16835 (N_16835,N_9596,N_11928);
nor U16836 (N_16836,N_9399,N_8713);
and U16837 (N_16837,N_6927,N_7622);
xor U16838 (N_16838,N_11253,N_11687);
nand U16839 (N_16839,N_6541,N_12218);
and U16840 (N_16840,N_8838,N_12424);
nor U16841 (N_16841,N_7042,N_10621);
and U16842 (N_16842,N_8349,N_12314);
nor U16843 (N_16843,N_8621,N_7080);
or U16844 (N_16844,N_6759,N_8070);
nor U16845 (N_16845,N_12152,N_11602);
or U16846 (N_16846,N_12281,N_12172);
nand U16847 (N_16847,N_9970,N_8249);
or U16848 (N_16848,N_10367,N_8638);
nand U16849 (N_16849,N_10839,N_10700);
or U16850 (N_16850,N_7576,N_8474);
nor U16851 (N_16851,N_9308,N_12333);
and U16852 (N_16852,N_6729,N_9768);
nand U16853 (N_16853,N_12314,N_11089);
nor U16854 (N_16854,N_11722,N_12195);
and U16855 (N_16855,N_6439,N_7197);
nand U16856 (N_16856,N_6898,N_9917);
and U16857 (N_16857,N_8075,N_9294);
nor U16858 (N_16858,N_6877,N_7192);
and U16859 (N_16859,N_8305,N_6525);
or U16860 (N_16860,N_12483,N_10654);
xor U16861 (N_16861,N_8001,N_9357);
and U16862 (N_16862,N_11916,N_10189);
and U16863 (N_16863,N_8511,N_8520);
xor U16864 (N_16864,N_9001,N_8811);
xnor U16865 (N_16865,N_9560,N_10114);
or U16866 (N_16866,N_7168,N_9597);
and U16867 (N_16867,N_6664,N_8159);
or U16868 (N_16868,N_11332,N_8909);
nand U16869 (N_16869,N_11200,N_12296);
and U16870 (N_16870,N_9210,N_11827);
nand U16871 (N_16871,N_11590,N_9251);
nor U16872 (N_16872,N_8370,N_11038);
nand U16873 (N_16873,N_6488,N_12338);
nor U16874 (N_16874,N_6554,N_11303);
or U16875 (N_16875,N_12312,N_10184);
nand U16876 (N_16876,N_7956,N_6463);
and U16877 (N_16877,N_10542,N_9886);
nand U16878 (N_16878,N_11710,N_11550);
nor U16879 (N_16879,N_6425,N_9406);
or U16880 (N_16880,N_9547,N_10208);
or U16881 (N_16881,N_6967,N_11793);
or U16882 (N_16882,N_9753,N_12374);
or U16883 (N_16883,N_8950,N_10175);
nand U16884 (N_16884,N_11396,N_8020);
nor U16885 (N_16885,N_7918,N_7334);
or U16886 (N_16886,N_7362,N_10699);
nand U16887 (N_16887,N_11835,N_8055);
or U16888 (N_16888,N_8563,N_7696);
nand U16889 (N_16889,N_12475,N_9561);
and U16890 (N_16890,N_12109,N_6629);
nand U16891 (N_16891,N_6821,N_12462);
and U16892 (N_16892,N_8119,N_6499);
and U16893 (N_16893,N_9781,N_9272);
or U16894 (N_16894,N_10958,N_9831);
nor U16895 (N_16895,N_6422,N_10635);
xnor U16896 (N_16896,N_8271,N_8379);
or U16897 (N_16897,N_12392,N_6882);
or U16898 (N_16898,N_12210,N_9095);
nand U16899 (N_16899,N_9767,N_9661);
or U16900 (N_16900,N_6364,N_7094);
nand U16901 (N_16901,N_11470,N_11210);
nand U16902 (N_16902,N_7453,N_10048);
and U16903 (N_16903,N_11000,N_10992);
and U16904 (N_16904,N_8327,N_7873);
xor U16905 (N_16905,N_6543,N_7268);
and U16906 (N_16906,N_11760,N_9078);
and U16907 (N_16907,N_11312,N_7382);
and U16908 (N_16908,N_6382,N_9549);
and U16909 (N_16909,N_10693,N_8367);
nand U16910 (N_16910,N_10912,N_9483);
nand U16911 (N_16911,N_6710,N_7613);
xnor U16912 (N_16912,N_7497,N_6953);
xor U16913 (N_16913,N_8194,N_11779);
nand U16914 (N_16914,N_8404,N_8170);
and U16915 (N_16915,N_6476,N_12446);
nand U16916 (N_16916,N_11003,N_6300);
and U16917 (N_16917,N_10669,N_11903);
and U16918 (N_16918,N_10846,N_11001);
nor U16919 (N_16919,N_10534,N_10688);
nand U16920 (N_16920,N_8525,N_9915);
nor U16921 (N_16921,N_7973,N_12141);
nand U16922 (N_16922,N_7710,N_8131);
or U16923 (N_16923,N_6420,N_8148);
nor U16924 (N_16924,N_8023,N_11691);
xnor U16925 (N_16925,N_10143,N_10088);
xnor U16926 (N_16926,N_7372,N_6537);
nand U16927 (N_16927,N_10478,N_6514);
and U16928 (N_16928,N_8795,N_9506);
and U16929 (N_16929,N_11422,N_11551);
or U16930 (N_16930,N_9369,N_6630);
and U16931 (N_16931,N_11692,N_11943);
nor U16932 (N_16932,N_10386,N_10858);
and U16933 (N_16933,N_11509,N_6770);
and U16934 (N_16934,N_8094,N_6387);
nor U16935 (N_16935,N_8837,N_7494);
or U16936 (N_16936,N_11785,N_11438);
nor U16937 (N_16937,N_10258,N_6441);
nand U16938 (N_16938,N_8932,N_7144);
nor U16939 (N_16939,N_8234,N_10985);
nand U16940 (N_16940,N_9486,N_9765);
nand U16941 (N_16941,N_7904,N_11295);
or U16942 (N_16942,N_6618,N_9430);
or U16943 (N_16943,N_10099,N_6554);
and U16944 (N_16944,N_9494,N_9956);
or U16945 (N_16945,N_10845,N_11784);
xor U16946 (N_16946,N_9476,N_7045);
nand U16947 (N_16947,N_11054,N_7695);
nor U16948 (N_16948,N_7093,N_8553);
or U16949 (N_16949,N_8446,N_10967);
and U16950 (N_16950,N_11847,N_10225);
nand U16951 (N_16951,N_7988,N_9114);
or U16952 (N_16952,N_6793,N_9572);
or U16953 (N_16953,N_12428,N_6264);
nor U16954 (N_16954,N_10754,N_11047);
and U16955 (N_16955,N_9901,N_7754);
and U16956 (N_16956,N_12065,N_12253);
nor U16957 (N_16957,N_11020,N_12407);
xor U16958 (N_16958,N_9656,N_7361);
nor U16959 (N_16959,N_8298,N_8599);
xnor U16960 (N_16960,N_8741,N_9349);
nor U16961 (N_16961,N_12054,N_10277);
nand U16962 (N_16962,N_11639,N_10128);
nand U16963 (N_16963,N_12399,N_7446);
nand U16964 (N_16964,N_8776,N_8208);
xnor U16965 (N_16965,N_10319,N_9700);
or U16966 (N_16966,N_7638,N_7265);
or U16967 (N_16967,N_8330,N_9716);
nand U16968 (N_16968,N_6469,N_6985);
or U16969 (N_16969,N_11675,N_10767);
xnor U16970 (N_16970,N_11526,N_10716);
or U16971 (N_16971,N_6591,N_9722);
nand U16972 (N_16972,N_9962,N_6385);
xnor U16973 (N_16973,N_9595,N_10603);
nand U16974 (N_16974,N_8341,N_11321);
or U16975 (N_16975,N_8615,N_7899);
and U16976 (N_16976,N_6371,N_8853);
nand U16977 (N_16977,N_6310,N_9846);
and U16978 (N_16978,N_9201,N_11144);
and U16979 (N_16979,N_8889,N_8697);
and U16980 (N_16980,N_12055,N_8874);
and U16981 (N_16981,N_11497,N_10178);
and U16982 (N_16982,N_11694,N_6954);
or U16983 (N_16983,N_10999,N_9459);
nor U16984 (N_16984,N_7941,N_8943);
nand U16985 (N_16985,N_10419,N_12419);
nor U16986 (N_16986,N_8607,N_10763);
xor U16987 (N_16987,N_8353,N_7549);
nand U16988 (N_16988,N_10636,N_8082);
nor U16989 (N_16989,N_11103,N_10861);
nor U16990 (N_16990,N_11730,N_6347);
xnor U16991 (N_16991,N_8348,N_8095);
and U16992 (N_16992,N_8701,N_7113);
xnor U16993 (N_16993,N_9517,N_12091);
and U16994 (N_16994,N_7305,N_10151);
and U16995 (N_16995,N_11191,N_7108);
nor U16996 (N_16996,N_10588,N_11963);
nor U16997 (N_16997,N_11874,N_11124);
or U16998 (N_16998,N_7997,N_8541);
nor U16999 (N_16999,N_10155,N_10552);
nor U17000 (N_17000,N_9715,N_11550);
and U17001 (N_17001,N_11726,N_8690);
nor U17002 (N_17002,N_10318,N_10114);
or U17003 (N_17003,N_8862,N_10216);
or U17004 (N_17004,N_9463,N_9064);
nand U17005 (N_17005,N_10655,N_10560);
or U17006 (N_17006,N_8859,N_9017);
or U17007 (N_17007,N_9188,N_8632);
or U17008 (N_17008,N_11552,N_8313);
xor U17009 (N_17009,N_11105,N_9215);
nor U17010 (N_17010,N_10424,N_9314);
xor U17011 (N_17011,N_7552,N_6841);
or U17012 (N_17012,N_7622,N_7083);
and U17013 (N_17013,N_9371,N_7322);
xnor U17014 (N_17014,N_8108,N_8845);
and U17015 (N_17015,N_10888,N_6713);
xor U17016 (N_17016,N_7071,N_9361);
and U17017 (N_17017,N_9021,N_7972);
nand U17018 (N_17018,N_6867,N_11333);
and U17019 (N_17019,N_9286,N_6511);
and U17020 (N_17020,N_11620,N_6960);
or U17021 (N_17021,N_12221,N_6677);
or U17022 (N_17022,N_9609,N_9695);
nand U17023 (N_17023,N_7434,N_8823);
or U17024 (N_17024,N_8993,N_9500);
nor U17025 (N_17025,N_10513,N_9361);
nor U17026 (N_17026,N_8515,N_6327);
and U17027 (N_17027,N_12391,N_9844);
xor U17028 (N_17028,N_11524,N_11586);
and U17029 (N_17029,N_10190,N_8349);
and U17030 (N_17030,N_10107,N_6757);
and U17031 (N_17031,N_8474,N_12437);
nor U17032 (N_17032,N_8318,N_10688);
xor U17033 (N_17033,N_7090,N_9476);
nand U17034 (N_17034,N_11951,N_9011);
nand U17035 (N_17035,N_9154,N_9132);
or U17036 (N_17036,N_8326,N_8978);
xor U17037 (N_17037,N_11728,N_6505);
or U17038 (N_17038,N_7080,N_12081);
nand U17039 (N_17039,N_7249,N_7393);
or U17040 (N_17040,N_10498,N_11016);
xor U17041 (N_17041,N_9064,N_7145);
and U17042 (N_17042,N_8852,N_6825);
or U17043 (N_17043,N_6813,N_8288);
nor U17044 (N_17044,N_6807,N_10690);
xnor U17045 (N_17045,N_11757,N_9010);
nand U17046 (N_17046,N_7423,N_12317);
and U17047 (N_17047,N_10317,N_9550);
and U17048 (N_17048,N_8307,N_9717);
nand U17049 (N_17049,N_10258,N_8933);
and U17050 (N_17050,N_8706,N_8441);
and U17051 (N_17051,N_10217,N_6458);
and U17052 (N_17052,N_10888,N_12270);
nor U17053 (N_17053,N_9998,N_6812);
xor U17054 (N_17054,N_11266,N_11806);
nand U17055 (N_17055,N_10456,N_8211);
nor U17056 (N_17056,N_9880,N_11170);
xnor U17057 (N_17057,N_11052,N_6431);
or U17058 (N_17058,N_12315,N_11253);
xor U17059 (N_17059,N_8108,N_6861);
xnor U17060 (N_17060,N_9433,N_11155);
and U17061 (N_17061,N_9145,N_11713);
or U17062 (N_17062,N_11967,N_10368);
nand U17063 (N_17063,N_8023,N_11932);
or U17064 (N_17064,N_8510,N_7411);
and U17065 (N_17065,N_6358,N_8830);
nand U17066 (N_17066,N_6346,N_11804);
or U17067 (N_17067,N_9606,N_7783);
nor U17068 (N_17068,N_7739,N_9911);
nor U17069 (N_17069,N_8501,N_10720);
xor U17070 (N_17070,N_11613,N_12194);
nand U17071 (N_17071,N_10927,N_12496);
nor U17072 (N_17072,N_9880,N_10788);
nand U17073 (N_17073,N_7477,N_10824);
or U17074 (N_17074,N_9635,N_8889);
and U17075 (N_17075,N_9948,N_9992);
nand U17076 (N_17076,N_7628,N_7673);
nand U17077 (N_17077,N_10991,N_12136);
nand U17078 (N_17078,N_9912,N_7148);
xor U17079 (N_17079,N_8900,N_7607);
nor U17080 (N_17080,N_11768,N_7239);
nand U17081 (N_17081,N_11408,N_8890);
and U17082 (N_17082,N_11751,N_11086);
nand U17083 (N_17083,N_6665,N_12106);
and U17084 (N_17084,N_8636,N_9006);
or U17085 (N_17085,N_10570,N_9974);
or U17086 (N_17086,N_11814,N_9930);
xnor U17087 (N_17087,N_11981,N_11735);
or U17088 (N_17088,N_10446,N_7028);
xor U17089 (N_17089,N_9025,N_9150);
nand U17090 (N_17090,N_10465,N_9836);
and U17091 (N_17091,N_6912,N_9315);
and U17092 (N_17092,N_8094,N_7756);
nand U17093 (N_17093,N_7593,N_6385);
or U17094 (N_17094,N_6727,N_7461);
and U17095 (N_17095,N_7613,N_10974);
nor U17096 (N_17096,N_11315,N_7388);
nand U17097 (N_17097,N_9718,N_9431);
nor U17098 (N_17098,N_10844,N_11819);
or U17099 (N_17099,N_9030,N_8346);
nand U17100 (N_17100,N_7968,N_11922);
or U17101 (N_17101,N_7257,N_6573);
or U17102 (N_17102,N_6334,N_10625);
and U17103 (N_17103,N_6544,N_9725);
nor U17104 (N_17104,N_6976,N_11307);
nand U17105 (N_17105,N_9709,N_12361);
and U17106 (N_17106,N_10700,N_10862);
and U17107 (N_17107,N_7216,N_7034);
nand U17108 (N_17108,N_6924,N_11122);
xor U17109 (N_17109,N_9962,N_8180);
xnor U17110 (N_17110,N_7974,N_10086);
and U17111 (N_17111,N_11265,N_7617);
and U17112 (N_17112,N_8066,N_9366);
nor U17113 (N_17113,N_8681,N_11321);
or U17114 (N_17114,N_6863,N_10663);
xor U17115 (N_17115,N_8446,N_9429);
and U17116 (N_17116,N_7150,N_12099);
or U17117 (N_17117,N_7669,N_9598);
or U17118 (N_17118,N_12248,N_8666);
xor U17119 (N_17119,N_8490,N_8061);
xnor U17120 (N_17120,N_10640,N_7694);
or U17121 (N_17121,N_7683,N_9469);
nor U17122 (N_17122,N_9119,N_10413);
nand U17123 (N_17123,N_9652,N_6929);
xor U17124 (N_17124,N_7169,N_11063);
and U17125 (N_17125,N_6397,N_9732);
nor U17126 (N_17126,N_10527,N_12450);
nand U17127 (N_17127,N_12304,N_8983);
nand U17128 (N_17128,N_7903,N_10813);
xor U17129 (N_17129,N_9271,N_7178);
or U17130 (N_17130,N_10438,N_7987);
xnor U17131 (N_17131,N_10067,N_9833);
nor U17132 (N_17132,N_8128,N_10715);
xor U17133 (N_17133,N_8198,N_10780);
xor U17134 (N_17134,N_7382,N_7545);
nor U17135 (N_17135,N_7988,N_8102);
and U17136 (N_17136,N_9397,N_10552);
nand U17137 (N_17137,N_8688,N_12104);
nand U17138 (N_17138,N_9481,N_6769);
nand U17139 (N_17139,N_11304,N_8847);
and U17140 (N_17140,N_6803,N_12137);
xor U17141 (N_17141,N_7997,N_11984);
nand U17142 (N_17142,N_12373,N_11845);
nand U17143 (N_17143,N_6274,N_9900);
nand U17144 (N_17144,N_11353,N_11338);
xor U17145 (N_17145,N_6594,N_10531);
and U17146 (N_17146,N_6870,N_10163);
xnor U17147 (N_17147,N_7912,N_8287);
or U17148 (N_17148,N_7984,N_6467);
or U17149 (N_17149,N_9901,N_11405);
nand U17150 (N_17150,N_9692,N_10306);
nand U17151 (N_17151,N_6921,N_9675);
and U17152 (N_17152,N_11888,N_8001);
and U17153 (N_17153,N_7454,N_12400);
or U17154 (N_17154,N_12357,N_7797);
nand U17155 (N_17155,N_7826,N_10304);
nand U17156 (N_17156,N_11567,N_12325);
xnor U17157 (N_17157,N_9076,N_9411);
or U17158 (N_17158,N_8234,N_10843);
xor U17159 (N_17159,N_9954,N_6939);
nor U17160 (N_17160,N_8834,N_9439);
and U17161 (N_17161,N_11281,N_11384);
nor U17162 (N_17162,N_11173,N_9519);
nand U17163 (N_17163,N_10863,N_12249);
nand U17164 (N_17164,N_11434,N_7269);
nand U17165 (N_17165,N_11930,N_7257);
nor U17166 (N_17166,N_10340,N_12382);
nor U17167 (N_17167,N_10849,N_8389);
nor U17168 (N_17168,N_9889,N_9380);
nor U17169 (N_17169,N_10442,N_11906);
nand U17170 (N_17170,N_6753,N_9008);
and U17171 (N_17171,N_9887,N_7215);
xnor U17172 (N_17172,N_11098,N_8880);
nand U17173 (N_17173,N_7984,N_9629);
and U17174 (N_17174,N_7130,N_7451);
and U17175 (N_17175,N_11618,N_6507);
or U17176 (N_17176,N_9248,N_10385);
xor U17177 (N_17177,N_10702,N_10032);
and U17178 (N_17178,N_7474,N_10107);
and U17179 (N_17179,N_11285,N_11425);
xor U17180 (N_17180,N_9826,N_9897);
nand U17181 (N_17181,N_9632,N_10060);
nand U17182 (N_17182,N_7221,N_11302);
or U17183 (N_17183,N_10208,N_12153);
or U17184 (N_17184,N_9003,N_7946);
nand U17185 (N_17185,N_8351,N_6485);
and U17186 (N_17186,N_9083,N_9367);
xor U17187 (N_17187,N_11266,N_8536);
nor U17188 (N_17188,N_11263,N_8305);
nand U17189 (N_17189,N_10025,N_6422);
and U17190 (N_17190,N_11516,N_12088);
nor U17191 (N_17191,N_8032,N_11254);
xnor U17192 (N_17192,N_8602,N_7589);
nand U17193 (N_17193,N_10987,N_9221);
nor U17194 (N_17194,N_6287,N_10247);
and U17195 (N_17195,N_11427,N_8291);
xnor U17196 (N_17196,N_8500,N_6366);
and U17197 (N_17197,N_6920,N_11961);
xnor U17198 (N_17198,N_10949,N_7545);
xor U17199 (N_17199,N_10966,N_6718);
nand U17200 (N_17200,N_11597,N_9651);
or U17201 (N_17201,N_8001,N_9882);
and U17202 (N_17202,N_6704,N_9107);
xor U17203 (N_17203,N_10695,N_8496);
nor U17204 (N_17204,N_11999,N_10247);
or U17205 (N_17205,N_11682,N_10573);
nor U17206 (N_17206,N_10956,N_9674);
xnor U17207 (N_17207,N_6757,N_8106);
xnor U17208 (N_17208,N_10287,N_9848);
and U17209 (N_17209,N_12139,N_7171);
or U17210 (N_17210,N_11636,N_6877);
nand U17211 (N_17211,N_7131,N_11932);
and U17212 (N_17212,N_6644,N_10450);
xnor U17213 (N_17213,N_10039,N_7331);
or U17214 (N_17214,N_8150,N_6626);
nand U17215 (N_17215,N_6297,N_12211);
nand U17216 (N_17216,N_8093,N_7840);
xnor U17217 (N_17217,N_7427,N_11968);
nand U17218 (N_17218,N_8144,N_9704);
nand U17219 (N_17219,N_11988,N_8803);
and U17220 (N_17220,N_10406,N_7625);
nand U17221 (N_17221,N_8760,N_9839);
nand U17222 (N_17222,N_9951,N_8618);
and U17223 (N_17223,N_8819,N_9796);
or U17224 (N_17224,N_8591,N_10947);
nor U17225 (N_17225,N_8341,N_6320);
xor U17226 (N_17226,N_11070,N_9223);
xor U17227 (N_17227,N_7626,N_12100);
nand U17228 (N_17228,N_12295,N_10871);
and U17229 (N_17229,N_7217,N_6461);
or U17230 (N_17230,N_7812,N_11620);
nor U17231 (N_17231,N_9261,N_7428);
nand U17232 (N_17232,N_11581,N_8749);
nand U17233 (N_17233,N_11516,N_12450);
and U17234 (N_17234,N_7873,N_8516);
and U17235 (N_17235,N_12489,N_11053);
nand U17236 (N_17236,N_8395,N_11487);
and U17237 (N_17237,N_8655,N_11987);
xnor U17238 (N_17238,N_8922,N_10173);
nand U17239 (N_17239,N_11454,N_12132);
or U17240 (N_17240,N_12321,N_12203);
nor U17241 (N_17241,N_7527,N_8462);
or U17242 (N_17242,N_7512,N_9574);
or U17243 (N_17243,N_8964,N_7610);
nand U17244 (N_17244,N_6586,N_11867);
nor U17245 (N_17245,N_11253,N_9616);
nor U17246 (N_17246,N_7290,N_10695);
or U17247 (N_17247,N_7973,N_9691);
or U17248 (N_17248,N_7242,N_12428);
nor U17249 (N_17249,N_8936,N_10046);
and U17250 (N_17250,N_7938,N_7658);
xor U17251 (N_17251,N_9584,N_7098);
xnor U17252 (N_17252,N_12256,N_11831);
nor U17253 (N_17253,N_6485,N_9903);
or U17254 (N_17254,N_7775,N_6619);
xor U17255 (N_17255,N_11406,N_7989);
and U17256 (N_17256,N_7121,N_7376);
or U17257 (N_17257,N_9065,N_11798);
and U17258 (N_17258,N_12345,N_9033);
xor U17259 (N_17259,N_10776,N_9328);
and U17260 (N_17260,N_9898,N_8545);
or U17261 (N_17261,N_9217,N_8072);
xnor U17262 (N_17262,N_12049,N_10712);
xnor U17263 (N_17263,N_11049,N_6670);
xor U17264 (N_17264,N_8452,N_12044);
nand U17265 (N_17265,N_10746,N_8861);
or U17266 (N_17266,N_10791,N_6264);
or U17267 (N_17267,N_12010,N_12259);
nand U17268 (N_17268,N_6881,N_11298);
and U17269 (N_17269,N_10510,N_8208);
nand U17270 (N_17270,N_11867,N_12299);
nor U17271 (N_17271,N_7724,N_8008);
nor U17272 (N_17272,N_9768,N_9750);
or U17273 (N_17273,N_11886,N_11152);
xnor U17274 (N_17274,N_11331,N_10129);
or U17275 (N_17275,N_7562,N_12045);
nor U17276 (N_17276,N_11053,N_10086);
xor U17277 (N_17277,N_9838,N_7495);
or U17278 (N_17278,N_9654,N_7045);
xnor U17279 (N_17279,N_6731,N_11642);
or U17280 (N_17280,N_8314,N_9592);
nand U17281 (N_17281,N_7254,N_11289);
xnor U17282 (N_17282,N_11712,N_6396);
xnor U17283 (N_17283,N_12336,N_11725);
nor U17284 (N_17284,N_10794,N_9420);
xnor U17285 (N_17285,N_11102,N_10001);
nor U17286 (N_17286,N_12095,N_9320);
and U17287 (N_17287,N_7985,N_9578);
or U17288 (N_17288,N_11306,N_10234);
xnor U17289 (N_17289,N_9898,N_8488);
xnor U17290 (N_17290,N_8382,N_6505);
nand U17291 (N_17291,N_11426,N_11239);
xnor U17292 (N_17292,N_6926,N_11422);
and U17293 (N_17293,N_10930,N_8552);
xor U17294 (N_17294,N_6278,N_6848);
or U17295 (N_17295,N_7989,N_9384);
nor U17296 (N_17296,N_7159,N_8992);
and U17297 (N_17297,N_11011,N_9862);
nand U17298 (N_17298,N_11621,N_6989);
or U17299 (N_17299,N_8654,N_8320);
xor U17300 (N_17300,N_10785,N_7593);
and U17301 (N_17301,N_11193,N_11576);
xor U17302 (N_17302,N_9406,N_6550);
nor U17303 (N_17303,N_10421,N_8601);
and U17304 (N_17304,N_11499,N_11988);
nand U17305 (N_17305,N_7427,N_7212);
xnor U17306 (N_17306,N_9398,N_12098);
or U17307 (N_17307,N_10541,N_7367);
nand U17308 (N_17308,N_12028,N_10415);
and U17309 (N_17309,N_9013,N_11991);
or U17310 (N_17310,N_11765,N_10884);
nor U17311 (N_17311,N_7343,N_7336);
and U17312 (N_17312,N_8566,N_6545);
or U17313 (N_17313,N_11416,N_11537);
or U17314 (N_17314,N_10481,N_9331);
and U17315 (N_17315,N_7887,N_12473);
or U17316 (N_17316,N_6359,N_7426);
and U17317 (N_17317,N_10519,N_8057);
nor U17318 (N_17318,N_10482,N_11328);
xor U17319 (N_17319,N_7658,N_12490);
or U17320 (N_17320,N_10043,N_7757);
or U17321 (N_17321,N_6487,N_11328);
nand U17322 (N_17322,N_9602,N_11107);
xnor U17323 (N_17323,N_9311,N_8183);
or U17324 (N_17324,N_8137,N_7837);
xnor U17325 (N_17325,N_11955,N_11289);
nand U17326 (N_17326,N_8150,N_7573);
or U17327 (N_17327,N_8921,N_8325);
xor U17328 (N_17328,N_10466,N_9214);
nor U17329 (N_17329,N_7432,N_11370);
nor U17330 (N_17330,N_9758,N_7754);
nand U17331 (N_17331,N_11564,N_8559);
xnor U17332 (N_17332,N_8101,N_11487);
and U17333 (N_17333,N_10040,N_7109);
and U17334 (N_17334,N_10445,N_11890);
nor U17335 (N_17335,N_8236,N_9909);
nor U17336 (N_17336,N_8193,N_8180);
and U17337 (N_17337,N_12292,N_11176);
nand U17338 (N_17338,N_10325,N_10541);
and U17339 (N_17339,N_6479,N_11288);
nand U17340 (N_17340,N_10492,N_10839);
nor U17341 (N_17341,N_10463,N_8393);
or U17342 (N_17342,N_11319,N_11600);
nor U17343 (N_17343,N_11065,N_7750);
xor U17344 (N_17344,N_12088,N_9380);
nor U17345 (N_17345,N_8864,N_10128);
nor U17346 (N_17346,N_7818,N_6581);
nor U17347 (N_17347,N_9954,N_6277);
or U17348 (N_17348,N_12016,N_10178);
nand U17349 (N_17349,N_10030,N_11281);
and U17350 (N_17350,N_8094,N_9154);
xor U17351 (N_17351,N_6379,N_10888);
nor U17352 (N_17352,N_8380,N_11223);
and U17353 (N_17353,N_7018,N_11467);
xnor U17354 (N_17354,N_9926,N_9397);
or U17355 (N_17355,N_7556,N_7249);
xor U17356 (N_17356,N_11500,N_11974);
and U17357 (N_17357,N_10563,N_6849);
and U17358 (N_17358,N_6717,N_9898);
and U17359 (N_17359,N_10514,N_7154);
and U17360 (N_17360,N_12279,N_11514);
and U17361 (N_17361,N_8421,N_12440);
and U17362 (N_17362,N_12108,N_11771);
nand U17363 (N_17363,N_11808,N_8281);
nor U17364 (N_17364,N_9972,N_9384);
nand U17365 (N_17365,N_11044,N_6878);
xnor U17366 (N_17366,N_7535,N_11780);
and U17367 (N_17367,N_11720,N_9624);
xor U17368 (N_17368,N_11806,N_11987);
nand U17369 (N_17369,N_8975,N_9058);
nand U17370 (N_17370,N_10295,N_7073);
and U17371 (N_17371,N_6910,N_6392);
nand U17372 (N_17372,N_10178,N_10348);
nor U17373 (N_17373,N_11508,N_6521);
xnor U17374 (N_17374,N_9685,N_7490);
nor U17375 (N_17375,N_11952,N_10078);
nor U17376 (N_17376,N_7139,N_8254);
or U17377 (N_17377,N_12483,N_9230);
or U17378 (N_17378,N_12015,N_10719);
or U17379 (N_17379,N_11637,N_7018);
and U17380 (N_17380,N_9513,N_10106);
xnor U17381 (N_17381,N_6922,N_9730);
or U17382 (N_17382,N_9661,N_9127);
nand U17383 (N_17383,N_7781,N_9705);
nor U17384 (N_17384,N_11991,N_11127);
xnor U17385 (N_17385,N_7487,N_10953);
nor U17386 (N_17386,N_9937,N_9304);
nand U17387 (N_17387,N_9734,N_7995);
or U17388 (N_17388,N_6893,N_6953);
nand U17389 (N_17389,N_6795,N_6437);
or U17390 (N_17390,N_8973,N_9480);
nor U17391 (N_17391,N_10791,N_8412);
nand U17392 (N_17392,N_9534,N_11098);
or U17393 (N_17393,N_7610,N_11528);
nor U17394 (N_17394,N_11879,N_6804);
nor U17395 (N_17395,N_11784,N_7607);
nor U17396 (N_17396,N_12372,N_8984);
nand U17397 (N_17397,N_9146,N_11728);
nand U17398 (N_17398,N_11291,N_8652);
and U17399 (N_17399,N_9332,N_9542);
nand U17400 (N_17400,N_10597,N_10353);
xnor U17401 (N_17401,N_6335,N_8430);
or U17402 (N_17402,N_9416,N_10812);
and U17403 (N_17403,N_7412,N_6798);
xnor U17404 (N_17404,N_9902,N_7192);
or U17405 (N_17405,N_7727,N_6662);
xor U17406 (N_17406,N_11392,N_11421);
nor U17407 (N_17407,N_6497,N_10133);
and U17408 (N_17408,N_12026,N_8046);
and U17409 (N_17409,N_9519,N_7232);
nand U17410 (N_17410,N_10451,N_6995);
or U17411 (N_17411,N_11146,N_7164);
xor U17412 (N_17412,N_7831,N_6842);
xnor U17413 (N_17413,N_10769,N_10011);
and U17414 (N_17414,N_6541,N_6639);
nand U17415 (N_17415,N_6571,N_9562);
nor U17416 (N_17416,N_7788,N_7756);
nand U17417 (N_17417,N_11843,N_8951);
and U17418 (N_17418,N_6453,N_10026);
or U17419 (N_17419,N_10821,N_9265);
nand U17420 (N_17420,N_8123,N_12384);
xnor U17421 (N_17421,N_10407,N_10328);
xnor U17422 (N_17422,N_11246,N_8763);
nor U17423 (N_17423,N_8926,N_12322);
xor U17424 (N_17424,N_10225,N_8267);
nand U17425 (N_17425,N_8459,N_8022);
and U17426 (N_17426,N_11760,N_9444);
nor U17427 (N_17427,N_6886,N_6949);
and U17428 (N_17428,N_9028,N_12371);
nor U17429 (N_17429,N_10861,N_9937);
or U17430 (N_17430,N_7585,N_8301);
and U17431 (N_17431,N_12011,N_11470);
or U17432 (N_17432,N_11704,N_11748);
nor U17433 (N_17433,N_8497,N_8130);
nand U17434 (N_17434,N_9868,N_9161);
nor U17435 (N_17435,N_6690,N_11832);
xor U17436 (N_17436,N_12356,N_10701);
or U17437 (N_17437,N_11504,N_11860);
and U17438 (N_17438,N_7783,N_9653);
nor U17439 (N_17439,N_6642,N_9664);
nand U17440 (N_17440,N_6475,N_10543);
or U17441 (N_17441,N_8040,N_11427);
or U17442 (N_17442,N_11030,N_10139);
and U17443 (N_17443,N_8512,N_12256);
and U17444 (N_17444,N_9444,N_6486);
nand U17445 (N_17445,N_8686,N_11548);
and U17446 (N_17446,N_10652,N_10343);
xnor U17447 (N_17447,N_10195,N_8203);
xnor U17448 (N_17448,N_12158,N_10143);
or U17449 (N_17449,N_10332,N_11439);
xor U17450 (N_17450,N_9621,N_11882);
nand U17451 (N_17451,N_10469,N_11909);
or U17452 (N_17452,N_9663,N_11944);
nor U17453 (N_17453,N_8277,N_7151);
xnor U17454 (N_17454,N_11470,N_10623);
or U17455 (N_17455,N_9085,N_9460);
and U17456 (N_17456,N_10129,N_9958);
and U17457 (N_17457,N_12356,N_7121);
nand U17458 (N_17458,N_11955,N_8671);
or U17459 (N_17459,N_9522,N_7702);
and U17460 (N_17460,N_11463,N_9589);
or U17461 (N_17461,N_11492,N_11428);
and U17462 (N_17462,N_6334,N_6811);
nor U17463 (N_17463,N_12478,N_10424);
xor U17464 (N_17464,N_7937,N_8723);
nor U17465 (N_17465,N_7456,N_8773);
xor U17466 (N_17466,N_10538,N_10306);
nor U17467 (N_17467,N_7214,N_7866);
nand U17468 (N_17468,N_7137,N_12086);
nor U17469 (N_17469,N_8760,N_6865);
and U17470 (N_17470,N_7562,N_9374);
and U17471 (N_17471,N_6472,N_8496);
or U17472 (N_17472,N_8769,N_7722);
xor U17473 (N_17473,N_8458,N_10498);
xor U17474 (N_17474,N_8655,N_7760);
xor U17475 (N_17475,N_7242,N_9793);
nand U17476 (N_17476,N_8914,N_9895);
and U17477 (N_17477,N_10924,N_9701);
xnor U17478 (N_17478,N_10899,N_12396);
xnor U17479 (N_17479,N_8193,N_7935);
nand U17480 (N_17480,N_9224,N_7749);
nor U17481 (N_17481,N_9536,N_7500);
xnor U17482 (N_17482,N_8037,N_8990);
nor U17483 (N_17483,N_11314,N_8775);
and U17484 (N_17484,N_7114,N_8050);
xor U17485 (N_17485,N_12197,N_6448);
nand U17486 (N_17486,N_8125,N_6391);
or U17487 (N_17487,N_9981,N_9060);
nand U17488 (N_17488,N_6299,N_11378);
xnor U17489 (N_17489,N_11184,N_6993);
nand U17490 (N_17490,N_9084,N_8507);
and U17491 (N_17491,N_12164,N_12197);
and U17492 (N_17492,N_6561,N_6604);
xnor U17493 (N_17493,N_9730,N_7108);
nand U17494 (N_17494,N_7532,N_12471);
or U17495 (N_17495,N_10641,N_8690);
or U17496 (N_17496,N_10972,N_8150);
xor U17497 (N_17497,N_9312,N_7093);
or U17498 (N_17498,N_10044,N_7290);
and U17499 (N_17499,N_7371,N_9618);
or U17500 (N_17500,N_9915,N_10238);
or U17501 (N_17501,N_6367,N_10581);
nor U17502 (N_17502,N_7324,N_6648);
or U17503 (N_17503,N_11729,N_12024);
xnor U17504 (N_17504,N_7716,N_11308);
nor U17505 (N_17505,N_6708,N_9775);
nand U17506 (N_17506,N_11163,N_7388);
xor U17507 (N_17507,N_7862,N_10843);
nand U17508 (N_17508,N_7939,N_8556);
xnor U17509 (N_17509,N_12034,N_11516);
or U17510 (N_17510,N_6298,N_7437);
nor U17511 (N_17511,N_9076,N_10410);
xor U17512 (N_17512,N_9403,N_11919);
xor U17513 (N_17513,N_11975,N_12016);
xnor U17514 (N_17514,N_10770,N_9307);
xor U17515 (N_17515,N_7730,N_10983);
or U17516 (N_17516,N_10391,N_12269);
or U17517 (N_17517,N_10067,N_8152);
nor U17518 (N_17518,N_10883,N_10704);
nor U17519 (N_17519,N_10184,N_6652);
and U17520 (N_17520,N_6816,N_10176);
xor U17521 (N_17521,N_9253,N_11291);
or U17522 (N_17522,N_10836,N_11594);
xnor U17523 (N_17523,N_8684,N_12307);
nor U17524 (N_17524,N_9467,N_10170);
nor U17525 (N_17525,N_8395,N_9015);
nand U17526 (N_17526,N_8385,N_9150);
nor U17527 (N_17527,N_7999,N_10206);
nand U17528 (N_17528,N_9567,N_9688);
nor U17529 (N_17529,N_10353,N_9348);
xnor U17530 (N_17530,N_11714,N_10033);
or U17531 (N_17531,N_11162,N_10347);
and U17532 (N_17532,N_9232,N_6948);
nand U17533 (N_17533,N_10794,N_11617);
nor U17534 (N_17534,N_8700,N_7625);
nor U17535 (N_17535,N_8783,N_10577);
xnor U17536 (N_17536,N_8761,N_9746);
or U17537 (N_17537,N_9341,N_9739);
xor U17538 (N_17538,N_11515,N_8162);
or U17539 (N_17539,N_8915,N_10543);
nor U17540 (N_17540,N_6268,N_7161);
nand U17541 (N_17541,N_7568,N_11660);
nor U17542 (N_17542,N_12253,N_8442);
or U17543 (N_17543,N_10468,N_8653);
and U17544 (N_17544,N_10341,N_10105);
nor U17545 (N_17545,N_8597,N_9650);
xor U17546 (N_17546,N_12497,N_9511);
and U17547 (N_17547,N_7119,N_10907);
nor U17548 (N_17548,N_7625,N_10182);
nor U17549 (N_17549,N_7273,N_8443);
nand U17550 (N_17550,N_11226,N_7845);
nand U17551 (N_17551,N_8426,N_9752);
nand U17552 (N_17552,N_11063,N_11696);
xnor U17553 (N_17553,N_9448,N_8560);
nand U17554 (N_17554,N_11075,N_8617);
nor U17555 (N_17555,N_11921,N_12355);
nor U17556 (N_17556,N_6500,N_8789);
and U17557 (N_17557,N_11958,N_10636);
nand U17558 (N_17558,N_9223,N_9438);
and U17559 (N_17559,N_8096,N_10559);
xor U17560 (N_17560,N_8293,N_9896);
nand U17561 (N_17561,N_11218,N_11748);
or U17562 (N_17562,N_10649,N_8303);
nand U17563 (N_17563,N_6956,N_10416);
nor U17564 (N_17564,N_7805,N_7526);
nor U17565 (N_17565,N_6993,N_7494);
or U17566 (N_17566,N_11900,N_6269);
nor U17567 (N_17567,N_6489,N_6863);
or U17568 (N_17568,N_11270,N_11670);
nand U17569 (N_17569,N_6538,N_12122);
or U17570 (N_17570,N_6712,N_10912);
and U17571 (N_17571,N_7169,N_12382);
nor U17572 (N_17572,N_9399,N_12249);
xnor U17573 (N_17573,N_11931,N_9204);
nand U17574 (N_17574,N_12301,N_7143);
or U17575 (N_17575,N_8767,N_7737);
nand U17576 (N_17576,N_11096,N_7094);
xnor U17577 (N_17577,N_9861,N_11060);
nand U17578 (N_17578,N_10289,N_7648);
nor U17579 (N_17579,N_12249,N_6719);
nand U17580 (N_17580,N_12007,N_9217);
xnor U17581 (N_17581,N_7222,N_6678);
and U17582 (N_17582,N_11946,N_11934);
nand U17583 (N_17583,N_8289,N_7600);
or U17584 (N_17584,N_11544,N_9360);
nand U17585 (N_17585,N_10061,N_11210);
xor U17586 (N_17586,N_9413,N_10631);
nor U17587 (N_17587,N_12207,N_7086);
nand U17588 (N_17588,N_9796,N_11827);
or U17589 (N_17589,N_7340,N_7255);
nor U17590 (N_17590,N_7089,N_10882);
nor U17591 (N_17591,N_11686,N_12139);
or U17592 (N_17592,N_8350,N_12326);
and U17593 (N_17593,N_9866,N_9270);
or U17594 (N_17594,N_11805,N_11315);
xnor U17595 (N_17595,N_7250,N_11458);
or U17596 (N_17596,N_10164,N_11951);
nor U17597 (N_17597,N_9850,N_10389);
or U17598 (N_17598,N_9628,N_12283);
or U17599 (N_17599,N_8041,N_8584);
and U17600 (N_17600,N_9504,N_8396);
or U17601 (N_17601,N_7620,N_9685);
nor U17602 (N_17602,N_10213,N_8489);
xnor U17603 (N_17603,N_7519,N_9837);
and U17604 (N_17604,N_8341,N_8854);
and U17605 (N_17605,N_7503,N_9496);
or U17606 (N_17606,N_6286,N_9913);
xnor U17607 (N_17607,N_6332,N_10871);
or U17608 (N_17608,N_12323,N_8029);
nand U17609 (N_17609,N_10304,N_11802);
and U17610 (N_17610,N_9469,N_7738);
or U17611 (N_17611,N_11459,N_11647);
nand U17612 (N_17612,N_9080,N_11749);
and U17613 (N_17613,N_9678,N_10266);
or U17614 (N_17614,N_7127,N_11916);
and U17615 (N_17615,N_7386,N_9398);
or U17616 (N_17616,N_11363,N_8364);
or U17617 (N_17617,N_7759,N_7597);
nor U17618 (N_17618,N_12174,N_11234);
nor U17619 (N_17619,N_6371,N_8032);
xnor U17620 (N_17620,N_8074,N_7016);
and U17621 (N_17621,N_12322,N_11505);
or U17622 (N_17622,N_8268,N_11603);
nor U17623 (N_17623,N_6293,N_11507);
nand U17624 (N_17624,N_12490,N_6865);
or U17625 (N_17625,N_6384,N_7450);
or U17626 (N_17626,N_9819,N_6681);
nand U17627 (N_17627,N_7129,N_11837);
nor U17628 (N_17628,N_12005,N_7771);
nor U17629 (N_17629,N_9664,N_8390);
nand U17630 (N_17630,N_7154,N_6903);
and U17631 (N_17631,N_6256,N_11513);
nand U17632 (N_17632,N_6908,N_9827);
nor U17633 (N_17633,N_11503,N_9367);
nor U17634 (N_17634,N_7926,N_12149);
or U17635 (N_17635,N_11326,N_8689);
nor U17636 (N_17636,N_7327,N_6979);
nand U17637 (N_17637,N_9486,N_9258);
xnor U17638 (N_17638,N_9095,N_10988);
and U17639 (N_17639,N_9349,N_6757);
or U17640 (N_17640,N_11910,N_9707);
or U17641 (N_17641,N_8370,N_6967);
nand U17642 (N_17642,N_6956,N_9523);
and U17643 (N_17643,N_7183,N_9528);
and U17644 (N_17644,N_9615,N_10278);
and U17645 (N_17645,N_7690,N_8652);
and U17646 (N_17646,N_11966,N_8842);
nor U17647 (N_17647,N_6745,N_11784);
nand U17648 (N_17648,N_9806,N_10585);
xor U17649 (N_17649,N_7803,N_8843);
xnor U17650 (N_17650,N_9794,N_7684);
or U17651 (N_17651,N_6646,N_7031);
and U17652 (N_17652,N_10418,N_11974);
nand U17653 (N_17653,N_7360,N_7504);
and U17654 (N_17654,N_9875,N_10206);
or U17655 (N_17655,N_9108,N_8730);
nand U17656 (N_17656,N_11177,N_11120);
nand U17657 (N_17657,N_9859,N_9391);
xnor U17658 (N_17658,N_8182,N_10937);
xnor U17659 (N_17659,N_9789,N_9412);
xnor U17660 (N_17660,N_11841,N_7699);
or U17661 (N_17661,N_10511,N_8800);
and U17662 (N_17662,N_9295,N_9776);
xor U17663 (N_17663,N_6486,N_7550);
xor U17664 (N_17664,N_11403,N_11191);
nand U17665 (N_17665,N_11561,N_11386);
xor U17666 (N_17666,N_9307,N_6285);
and U17667 (N_17667,N_12343,N_7408);
nor U17668 (N_17668,N_10128,N_11021);
xor U17669 (N_17669,N_9378,N_12138);
or U17670 (N_17670,N_6608,N_11649);
or U17671 (N_17671,N_10576,N_12124);
or U17672 (N_17672,N_7887,N_7318);
xnor U17673 (N_17673,N_9921,N_10731);
or U17674 (N_17674,N_9066,N_9574);
or U17675 (N_17675,N_6629,N_9080);
and U17676 (N_17676,N_11446,N_10060);
and U17677 (N_17677,N_9586,N_9738);
and U17678 (N_17678,N_9929,N_8761);
and U17679 (N_17679,N_7382,N_6854);
nor U17680 (N_17680,N_6270,N_8810);
and U17681 (N_17681,N_9222,N_9485);
xnor U17682 (N_17682,N_10719,N_12156);
nand U17683 (N_17683,N_8974,N_11718);
and U17684 (N_17684,N_7441,N_8230);
and U17685 (N_17685,N_7234,N_12238);
nand U17686 (N_17686,N_11607,N_7818);
xnor U17687 (N_17687,N_11984,N_8610);
xor U17688 (N_17688,N_6921,N_11525);
and U17689 (N_17689,N_9540,N_10953);
xor U17690 (N_17690,N_12265,N_10355);
and U17691 (N_17691,N_7532,N_9268);
nand U17692 (N_17692,N_6426,N_11791);
or U17693 (N_17693,N_7928,N_12269);
and U17694 (N_17694,N_12244,N_6600);
or U17695 (N_17695,N_11552,N_9123);
and U17696 (N_17696,N_12280,N_12424);
or U17697 (N_17697,N_11212,N_11140);
or U17698 (N_17698,N_7532,N_9757);
nand U17699 (N_17699,N_11194,N_12279);
xor U17700 (N_17700,N_7019,N_12081);
xor U17701 (N_17701,N_10403,N_7906);
nand U17702 (N_17702,N_10701,N_7999);
nor U17703 (N_17703,N_9795,N_10455);
xnor U17704 (N_17704,N_10996,N_7441);
nor U17705 (N_17705,N_11913,N_11923);
xnor U17706 (N_17706,N_7316,N_6706);
and U17707 (N_17707,N_8174,N_8213);
or U17708 (N_17708,N_9798,N_11833);
and U17709 (N_17709,N_6956,N_10462);
xor U17710 (N_17710,N_10337,N_10519);
and U17711 (N_17711,N_6535,N_11685);
xor U17712 (N_17712,N_8716,N_8527);
nand U17713 (N_17713,N_11201,N_12199);
xnor U17714 (N_17714,N_9593,N_12242);
nand U17715 (N_17715,N_7756,N_6946);
and U17716 (N_17716,N_10266,N_7036);
or U17717 (N_17717,N_11095,N_11129);
nor U17718 (N_17718,N_8893,N_9220);
nor U17719 (N_17719,N_8822,N_10787);
nor U17720 (N_17720,N_10915,N_6988);
nor U17721 (N_17721,N_8138,N_10778);
nand U17722 (N_17722,N_11133,N_8309);
or U17723 (N_17723,N_9247,N_10191);
nor U17724 (N_17724,N_10218,N_7337);
and U17725 (N_17725,N_10906,N_9617);
or U17726 (N_17726,N_7421,N_8883);
and U17727 (N_17727,N_9525,N_8187);
or U17728 (N_17728,N_11257,N_11005);
nor U17729 (N_17729,N_12265,N_11709);
and U17730 (N_17730,N_6520,N_10164);
and U17731 (N_17731,N_9125,N_9006);
nand U17732 (N_17732,N_11663,N_6369);
nor U17733 (N_17733,N_9449,N_6906);
nand U17734 (N_17734,N_6609,N_7507);
nor U17735 (N_17735,N_11256,N_9140);
nor U17736 (N_17736,N_8017,N_11780);
or U17737 (N_17737,N_8723,N_8920);
nor U17738 (N_17738,N_11005,N_11376);
and U17739 (N_17739,N_7928,N_8390);
xor U17740 (N_17740,N_10824,N_9747);
or U17741 (N_17741,N_8678,N_11356);
or U17742 (N_17742,N_8812,N_10842);
xor U17743 (N_17743,N_10496,N_12358);
and U17744 (N_17744,N_9206,N_7050);
nand U17745 (N_17745,N_10502,N_9002);
nand U17746 (N_17746,N_8266,N_8542);
nand U17747 (N_17747,N_6656,N_8323);
nand U17748 (N_17748,N_12273,N_10057);
xnor U17749 (N_17749,N_7266,N_12459);
xnor U17750 (N_17750,N_8970,N_12468);
and U17751 (N_17751,N_10203,N_6914);
xnor U17752 (N_17752,N_10500,N_6960);
nand U17753 (N_17753,N_7989,N_8757);
and U17754 (N_17754,N_7664,N_6913);
or U17755 (N_17755,N_10117,N_8653);
and U17756 (N_17756,N_10676,N_8252);
nand U17757 (N_17757,N_6348,N_8585);
and U17758 (N_17758,N_6359,N_12079);
xor U17759 (N_17759,N_11919,N_6463);
or U17760 (N_17760,N_8200,N_10942);
nor U17761 (N_17761,N_11235,N_7954);
and U17762 (N_17762,N_7693,N_6475);
or U17763 (N_17763,N_6903,N_6952);
xor U17764 (N_17764,N_10429,N_11294);
nor U17765 (N_17765,N_11610,N_9735);
xor U17766 (N_17766,N_9935,N_8610);
nor U17767 (N_17767,N_8589,N_10098);
nor U17768 (N_17768,N_10453,N_9415);
xnor U17769 (N_17769,N_12425,N_11524);
nor U17770 (N_17770,N_10514,N_11707);
xnor U17771 (N_17771,N_9768,N_8572);
and U17772 (N_17772,N_12256,N_7007);
nor U17773 (N_17773,N_6830,N_7323);
or U17774 (N_17774,N_6410,N_8738);
or U17775 (N_17775,N_6534,N_12324);
and U17776 (N_17776,N_7292,N_8701);
or U17777 (N_17777,N_10450,N_7711);
xor U17778 (N_17778,N_8985,N_7616);
nor U17779 (N_17779,N_11066,N_7007);
nand U17780 (N_17780,N_9027,N_10877);
nand U17781 (N_17781,N_9125,N_12120);
nor U17782 (N_17782,N_10031,N_9743);
or U17783 (N_17783,N_12005,N_9303);
nand U17784 (N_17784,N_12222,N_7485);
xor U17785 (N_17785,N_12182,N_7575);
and U17786 (N_17786,N_6733,N_8701);
and U17787 (N_17787,N_11854,N_11244);
or U17788 (N_17788,N_6965,N_10999);
and U17789 (N_17789,N_12042,N_8782);
and U17790 (N_17790,N_6838,N_8066);
nor U17791 (N_17791,N_7848,N_11359);
nand U17792 (N_17792,N_7426,N_9538);
and U17793 (N_17793,N_7536,N_9275);
xnor U17794 (N_17794,N_11454,N_10206);
nor U17795 (N_17795,N_9030,N_10551);
nor U17796 (N_17796,N_8049,N_6931);
xnor U17797 (N_17797,N_9384,N_8088);
and U17798 (N_17798,N_9701,N_9310);
and U17799 (N_17799,N_11455,N_7963);
or U17800 (N_17800,N_7058,N_8801);
xnor U17801 (N_17801,N_8201,N_10790);
xor U17802 (N_17802,N_7381,N_6527);
and U17803 (N_17803,N_7285,N_7665);
and U17804 (N_17804,N_9957,N_11738);
and U17805 (N_17805,N_9371,N_8944);
nor U17806 (N_17806,N_6884,N_10506);
or U17807 (N_17807,N_11742,N_7360);
nand U17808 (N_17808,N_8889,N_9296);
and U17809 (N_17809,N_9605,N_7431);
nor U17810 (N_17810,N_11802,N_7865);
nor U17811 (N_17811,N_12324,N_8612);
nor U17812 (N_17812,N_9854,N_7638);
nand U17813 (N_17813,N_10368,N_10615);
nand U17814 (N_17814,N_10553,N_8883);
nand U17815 (N_17815,N_11886,N_12137);
nor U17816 (N_17816,N_11517,N_6404);
nor U17817 (N_17817,N_7100,N_10331);
nor U17818 (N_17818,N_11235,N_9535);
and U17819 (N_17819,N_12477,N_11320);
nor U17820 (N_17820,N_8669,N_8655);
and U17821 (N_17821,N_7547,N_10734);
and U17822 (N_17822,N_9233,N_11379);
xnor U17823 (N_17823,N_7280,N_11115);
xnor U17824 (N_17824,N_11763,N_10817);
nand U17825 (N_17825,N_9130,N_11184);
nand U17826 (N_17826,N_11020,N_7953);
and U17827 (N_17827,N_12308,N_8845);
nor U17828 (N_17828,N_6992,N_11753);
and U17829 (N_17829,N_11579,N_9295);
nor U17830 (N_17830,N_10897,N_9682);
or U17831 (N_17831,N_12204,N_11197);
or U17832 (N_17832,N_10187,N_7993);
nand U17833 (N_17833,N_7356,N_8754);
nor U17834 (N_17834,N_11511,N_11876);
nor U17835 (N_17835,N_11990,N_10308);
nor U17836 (N_17836,N_7704,N_9182);
and U17837 (N_17837,N_8760,N_11405);
and U17838 (N_17838,N_7711,N_12158);
nand U17839 (N_17839,N_8759,N_11820);
or U17840 (N_17840,N_11303,N_12202);
nand U17841 (N_17841,N_6505,N_6846);
xor U17842 (N_17842,N_11481,N_10362);
nor U17843 (N_17843,N_9335,N_6588);
nor U17844 (N_17844,N_12051,N_8952);
nor U17845 (N_17845,N_12266,N_10628);
xnor U17846 (N_17846,N_11679,N_11849);
and U17847 (N_17847,N_7233,N_9120);
nand U17848 (N_17848,N_11307,N_6450);
xnor U17849 (N_17849,N_10900,N_6866);
or U17850 (N_17850,N_6690,N_7557);
or U17851 (N_17851,N_12071,N_6884);
and U17852 (N_17852,N_7529,N_8218);
xnor U17853 (N_17853,N_9222,N_9053);
and U17854 (N_17854,N_11046,N_8337);
or U17855 (N_17855,N_8408,N_11827);
and U17856 (N_17856,N_11739,N_8962);
or U17857 (N_17857,N_6609,N_11446);
and U17858 (N_17858,N_7141,N_8458);
xnor U17859 (N_17859,N_11074,N_10045);
xor U17860 (N_17860,N_8077,N_7306);
nand U17861 (N_17861,N_9106,N_9681);
xor U17862 (N_17862,N_10654,N_10329);
nor U17863 (N_17863,N_9243,N_9966);
or U17864 (N_17864,N_12346,N_8597);
nor U17865 (N_17865,N_8729,N_12313);
xnor U17866 (N_17866,N_9569,N_10983);
xnor U17867 (N_17867,N_7819,N_7494);
or U17868 (N_17868,N_8977,N_6678);
nor U17869 (N_17869,N_10322,N_6951);
or U17870 (N_17870,N_10744,N_6532);
nand U17871 (N_17871,N_9873,N_8152);
nand U17872 (N_17872,N_9977,N_6418);
nand U17873 (N_17873,N_8300,N_7996);
nand U17874 (N_17874,N_10613,N_6756);
xor U17875 (N_17875,N_7549,N_9047);
nand U17876 (N_17876,N_11530,N_10482);
nand U17877 (N_17877,N_11473,N_6443);
nor U17878 (N_17878,N_10723,N_9496);
nor U17879 (N_17879,N_9550,N_7315);
and U17880 (N_17880,N_7528,N_11826);
nand U17881 (N_17881,N_7996,N_8921);
and U17882 (N_17882,N_11748,N_10502);
and U17883 (N_17883,N_6710,N_7850);
and U17884 (N_17884,N_11946,N_10961);
nand U17885 (N_17885,N_7803,N_7225);
or U17886 (N_17886,N_8671,N_6943);
xnor U17887 (N_17887,N_10641,N_9237);
nor U17888 (N_17888,N_8067,N_9542);
xnor U17889 (N_17889,N_9738,N_10809);
xor U17890 (N_17890,N_9717,N_9848);
nor U17891 (N_17891,N_8113,N_7227);
and U17892 (N_17892,N_8828,N_10717);
nor U17893 (N_17893,N_9917,N_8740);
nand U17894 (N_17894,N_9085,N_7787);
nand U17895 (N_17895,N_8352,N_11919);
nor U17896 (N_17896,N_8197,N_8584);
and U17897 (N_17897,N_10993,N_7907);
nor U17898 (N_17898,N_11839,N_9295);
nand U17899 (N_17899,N_6682,N_11961);
nor U17900 (N_17900,N_9032,N_11611);
nor U17901 (N_17901,N_12482,N_10088);
and U17902 (N_17902,N_12475,N_7209);
nor U17903 (N_17903,N_7845,N_7119);
nand U17904 (N_17904,N_7187,N_11326);
nor U17905 (N_17905,N_9709,N_10447);
nor U17906 (N_17906,N_8506,N_10602);
and U17907 (N_17907,N_10613,N_8573);
nand U17908 (N_17908,N_11256,N_7691);
or U17909 (N_17909,N_7038,N_10078);
xor U17910 (N_17910,N_10258,N_9839);
xnor U17911 (N_17911,N_12324,N_10084);
nor U17912 (N_17912,N_12495,N_7590);
and U17913 (N_17913,N_11708,N_11469);
and U17914 (N_17914,N_6749,N_10288);
xnor U17915 (N_17915,N_11402,N_11611);
xnor U17916 (N_17916,N_8592,N_9322);
and U17917 (N_17917,N_9744,N_6291);
nand U17918 (N_17918,N_12281,N_10596);
xor U17919 (N_17919,N_9917,N_8269);
xnor U17920 (N_17920,N_11626,N_8403);
nand U17921 (N_17921,N_7924,N_10278);
nor U17922 (N_17922,N_12020,N_9987);
xor U17923 (N_17923,N_7434,N_6825);
xnor U17924 (N_17924,N_8696,N_8400);
nand U17925 (N_17925,N_9668,N_10044);
or U17926 (N_17926,N_11035,N_8030);
xor U17927 (N_17927,N_10115,N_6982);
xor U17928 (N_17928,N_6528,N_12159);
xnor U17929 (N_17929,N_12163,N_7011);
nor U17930 (N_17930,N_7758,N_7595);
or U17931 (N_17931,N_7802,N_8693);
or U17932 (N_17932,N_12466,N_8941);
and U17933 (N_17933,N_7460,N_10952);
or U17934 (N_17934,N_8728,N_10054);
and U17935 (N_17935,N_8775,N_11735);
or U17936 (N_17936,N_8663,N_8480);
nand U17937 (N_17937,N_10601,N_10526);
nand U17938 (N_17938,N_7889,N_11666);
and U17939 (N_17939,N_11158,N_10607);
or U17940 (N_17940,N_10150,N_7333);
and U17941 (N_17941,N_10211,N_6981);
nand U17942 (N_17942,N_8928,N_11385);
nor U17943 (N_17943,N_10672,N_9955);
nand U17944 (N_17944,N_9881,N_8794);
and U17945 (N_17945,N_10769,N_8924);
nor U17946 (N_17946,N_9186,N_7006);
and U17947 (N_17947,N_10485,N_9944);
and U17948 (N_17948,N_9538,N_7873);
xnor U17949 (N_17949,N_7861,N_9843);
and U17950 (N_17950,N_7076,N_8787);
or U17951 (N_17951,N_12231,N_11000);
nand U17952 (N_17952,N_10630,N_8634);
nand U17953 (N_17953,N_7886,N_11143);
xnor U17954 (N_17954,N_9726,N_12055);
nand U17955 (N_17955,N_10795,N_9759);
xnor U17956 (N_17956,N_8487,N_12349);
nand U17957 (N_17957,N_8287,N_9869);
nand U17958 (N_17958,N_12066,N_8471);
xor U17959 (N_17959,N_12168,N_8838);
nor U17960 (N_17960,N_8422,N_11911);
xnor U17961 (N_17961,N_9603,N_12092);
xor U17962 (N_17962,N_10676,N_11743);
nand U17963 (N_17963,N_12374,N_8160);
xor U17964 (N_17964,N_11468,N_7633);
xnor U17965 (N_17965,N_6319,N_7701);
and U17966 (N_17966,N_7976,N_10489);
and U17967 (N_17967,N_11472,N_6814);
and U17968 (N_17968,N_9399,N_8732);
nand U17969 (N_17969,N_8472,N_11745);
or U17970 (N_17970,N_9346,N_9912);
and U17971 (N_17971,N_11778,N_9138);
nor U17972 (N_17972,N_10237,N_8906);
or U17973 (N_17973,N_7312,N_9686);
or U17974 (N_17974,N_7395,N_11252);
and U17975 (N_17975,N_9337,N_9946);
and U17976 (N_17976,N_6323,N_10746);
nand U17977 (N_17977,N_8874,N_11852);
or U17978 (N_17978,N_11731,N_8284);
xor U17979 (N_17979,N_9826,N_7410);
and U17980 (N_17980,N_11322,N_9925);
xor U17981 (N_17981,N_7996,N_11768);
and U17982 (N_17982,N_10203,N_6426);
or U17983 (N_17983,N_9687,N_7037);
and U17984 (N_17984,N_8453,N_7425);
and U17985 (N_17985,N_7338,N_7249);
nand U17986 (N_17986,N_9950,N_8706);
xnor U17987 (N_17987,N_10754,N_8014);
xnor U17988 (N_17988,N_7655,N_11427);
or U17989 (N_17989,N_6546,N_8275);
xnor U17990 (N_17990,N_9120,N_6876);
or U17991 (N_17991,N_9978,N_9920);
or U17992 (N_17992,N_8934,N_8371);
xnor U17993 (N_17993,N_11640,N_7332);
and U17994 (N_17994,N_11015,N_10400);
or U17995 (N_17995,N_10999,N_8369);
nand U17996 (N_17996,N_9635,N_12030);
and U17997 (N_17997,N_6320,N_9648);
and U17998 (N_17998,N_8936,N_9947);
nand U17999 (N_17999,N_6421,N_6889);
or U18000 (N_18000,N_11994,N_11964);
nor U18001 (N_18001,N_7976,N_7129);
nand U18002 (N_18002,N_9340,N_7179);
xnor U18003 (N_18003,N_9558,N_7122);
or U18004 (N_18004,N_8564,N_9802);
nor U18005 (N_18005,N_12189,N_12145);
nand U18006 (N_18006,N_7113,N_11882);
and U18007 (N_18007,N_8456,N_7717);
nor U18008 (N_18008,N_9395,N_9945);
nor U18009 (N_18009,N_7523,N_9749);
nand U18010 (N_18010,N_10756,N_12328);
xnor U18011 (N_18011,N_8394,N_10918);
and U18012 (N_18012,N_9148,N_12346);
nand U18013 (N_18013,N_11605,N_12441);
xnor U18014 (N_18014,N_6776,N_9096);
and U18015 (N_18015,N_7281,N_6320);
or U18016 (N_18016,N_7529,N_8222);
and U18017 (N_18017,N_6355,N_11513);
nand U18018 (N_18018,N_9135,N_9438);
nand U18019 (N_18019,N_11178,N_7176);
xnor U18020 (N_18020,N_7282,N_6522);
or U18021 (N_18021,N_8199,N_9032);
nor U18022 (N_18022,N_12211,N_6419);
and U18023 (N_18023,N_6724,N_11549);
and U18024 (N_18024,N_7793,N_11491);
xor U18025 (N_18025,N_8262,N_9285);
and U18026 (N_18026,N_8520,N_11216);
nand U18027 (N_18027,N_8199,N_10940);
nor U18028 (N_18028,N_6565,N_7609);
and U18029 (N_18029,N_6506,N_9643);
nor U18030 (N_18030,N_7089,N_11602);
and U18031 (N_18031,N_9787,N_7503);
and U18032 (N_18032,N_7816,N_9120);
nor U18033 (N_18033,N_6468,N_11672);
or U18034 (N_18034,N_6253,N_9337);
nand U18035 (N_18035,N_8155,N_12457);
and U18036 (N_18036,N_9541,N_8755);
xor U18037 (N_18037,N_11372,N_10166);
nor U18038 (N_18038,N_8819,N_6688);
nor U18039 (N_18039,N_6384,N_7317);
nand U18040 (N_18040,N_9301,N_11564);
nand U18041 (N_18041,N_8458,N_9742);
nand U18042 (N_18042,N_9834,N_9149);
or U18043 (N_18043,N_6527,N_10582);
or U18044 (N_18044,N_12147,N_6520);
and U18045 (N_18045,N_10683,N_12448);
nand U18046 (N_18046,N_6770,N_6732);
nand U18047 (N_18047,N_7813,N_7822);
nor U18048 (N_18048,N_11972,N_10947);
or U18049 (N_18049,N_7705,N_12267);
nor U18050 (N_18050,N_10913,N_9489);
xnor U18051 (N_18051,N_8545,N_11921);
nand U18052 (N_18052,N_9400,N_8118);
nor U18053 (N_18053,N_10289,N_10460);
nand U18054 (N_18054,N_11602,N_10001);
xnor U18055 (N_18055,N_11459,N_12154);
xnor U18056 (N_18056,N_9773,N_10884);
or U18057 (N_18057,N_11358,N_9669);
nor U18058 (N_18058,N_7732,N_6908);
nand U18059 (N_18059,N_8565,N_12228);
and U18060 (N_18060,N_10325,N_11988);
or U18061 (N_18061,N_8833,N_12023);
xor U18062 (N_18062,N_10190,N_10302);
or U18063 (N_18063,N_11716,N_6696);
nand U18064 (N_18064,N_9639,N_12147);
and U18065 (N_18065,N_9094,N_11422);
xnor U18066 (N_18066,N_6764,N_6981);
xor U18067 (N_18067,N_7697,N_8459);
xor U18068 (N_18068,N_11485,N_10779);
nand U18069 (N_18069,N_10536,N_11178);
xor U18070 (N_18070,N_7319,N_8590);
xor U18071 (N_18071,N_8049,N_7172);
nand U18072 (N_18072,N_11558,N_8791);
and U18073 (N_18073,N_10917,N_9176);
or U18074 (N_18074,N_8746,N_8532);
xor U18075 (N_18075,N_12163,N_9843);
xnor U18076 (N_18076,N_8494,N_7775);
xor U18077 (N_18077,N_7410,N_10540);
or U18078 (N_18078,N_10078,N_11227);
xnor U18079 (N_18079,N_9116,N_6427);
xnor U18080 (N_18080,N_10907,N_6661);
and U18081 (N_18081,N_10298,N_11769);
xor U18082 (N_18082,N_11591,N_11605);
nor U18083 (N_18083,N_11172,N_11133);
xnor U18084 (N_18084,N_8740,N_6910);
nor U18085 (N_18085,N_6693,N_11763);
and U18086 (N_18086,N_6886,N_7106);
xnor U18087 (N_18087,N_10085,N_9495);
or U18088 (N_18088,N_8701,N_11664);
nor U18089 (N_18089,N_10404,N_8735);
xnor U18090 (N_18090,N_8708,N_12371);
or U18091 (N_18091,N_10380,N_11203);
nor U18092 (N_18092,N_9196,N_6360);
nand U18093 (N_18093,N_7117,N_9571);
or U18094 (N_18094,N_9725,N_12197);
or U18095 (N_18095,N_11082,N_11446);
nor U18096 (N_18096,N_11414,N_12299);
and U18097 (N_18097,N_11167,N_7498);
nor U18098 (N_18098,N_11781,N_6798);
and U18099 (N_18099,N_11340,N_6500);
nor U18100 (N_18100,N_6992,N_6578);
nor U18101 (N_18101,N_10596,N_8775);
xor U18102 (N_18102,N_10886,N_12354);
nor U18103 (N_18103,N_10572,N_10989);
nor U18104 (N_18104,N_7977,N_10496);
nand U18105 (N_18105,N_9185,N_11562);
xnor U18106 (N_18106,N_7137,N_6478);
xor U18107 (N_18107,N_6643,N_8290);
nand U18108 (N_18108,N_11146,N_9857);
xnor U18109 (N_18109,N_9940,N_8485);
or U18110 (N_18110,N_7602,N_10199);
nor U18111 (N_18111,N_7989,N_9808);
nor U18112 (N_18112,N_8494,N_11611);
or U18113 (N_18113,N_11892,N_10916);
and U18114 (N_18114,N_7060,N_9639);
or U18115 (N_18115,N_9423,N_6772);
xor U18116 (N_18116,N_9682,N_10942);
nor U18117 (N_18117,N_8413,N_9416);
nand U18118 (N_18118,N_11240,N_8595);
or U18119 (N_18119,N_7363,N_11650);
nor U18120 (N_18120,N_8237,N_11663);
or U18121 (N_18121,N_10174,N_11124);
nand U18122 (N_18122,N_9834,N_12178);
or U18123 (N_18123,N_8111,N_10624);
nand U18124 (N_18124,N_10468,N_10075);
or U18125 (N_18125,N_11230,N_6363);
and U18126 (N_18126,N_11766,N_8020);
nor U18127 (N_18127,N_8173,N_11464);
nand U18128 (N_18128,N_9420,N_7259);
nor U18129 (N_18129,N_7734,N_7093);
or U18130 (N_18130,N_11017,N_6466);
xnor U18131 (N_18131,N_9023,N_10504);
nand U18132 (N_18132,N_9378,N_7380);
and U18133 (N_18133,N_6684,N_11290);
nor U18134 (N_18134,N_11209,N_7986);
xor U18135 (N_18135,N_7183,N_11997);
xnor U18136 (N_18136,N_11149,N_9715);
xnor U18137 (N_18137,N_7044,N_10593);
nand U18138 (N_18138,N_7755,N_11328);
nand U18139 (N_18139,N_9299,N_9372);
or U18140 (N_18140,N_9761,N_9507);
or U18141 (N_18141,N_8552,N_7308);
and U18142 (N_18142,N_12283,N_7016);
nand U18143 (N_18143,N_8898,N_10966);
or U18144 (N_18144,N_8700,N_8266);
and U18145 (N_18145,N_11943,N_7247);
nor U18146 (N_18146,N_12260,N_7715);
or U18147 (N_18147,N_10958,N_8536);
nor U18148 (N_18148,N_7195,N_8348);
and U18149 (N_18149,N_8829,N_6858);
or U18150 (N_18150,N_9458,N_9978);
and U18151 (N_18151,N_11339,N_6476);
xnor U18152 (N_18152,N_6585,N_8364);
or U18153 (N_18153,N_10515,N_9696);
xor U18154 (N_18154,N_11908,N_9608);
nand U18155 (N_18155,N_9465,N_11012);
nand U18156 (N_18156,N_11763,N_10568);
nand U18157 (N_18157,N_10075,N_8232);
nand U18158 (N_18158,N_11842,N_8128);
xnor U18159 (N_18159,N_9188,N_10527);
and U18160 (N_18160,N_9583,N_11415);
nand U18161 (N_18161,N_9061,N_10973);
nand U18162 (N_18162,N_10333,N_12370);
nand U18163 (N_18163,N_12127,N_9121);
nand U18164 (N_18164,N_11824,N_11072);
and U18165 (N_18165,N_10903,N_9888);
nand U18166 (N_18166,N_8499,N_9914);
nand U18167 (N_18167,N_6601,N_9186);
nor U18168 (N_18168,N_10297,N_11863);
nand U18169 (N_18169,N_10859,N_12381);
nand U18170 (N_18170,N_12091,N_11333);
or U18171 (N_18171,N_10996,N_7049);
xnor U18172 (N_18172,N_9841,N_7845);
or U18173 (N_18173,N_9334,N_12153);
xnor U18174 (N_18174,N_8289,N_12390);
nor U18175 (N_18175,N_8652,N_9382);
xor U18176 (N_18176,N_11590,N_12192);
and U18177 (N_18177,N_8008,N_7990);
xnor U18178 (N_18178,N_8005,N_11675);
xor U18179 (N_18179,N_10024,N_8784);
or U18180 (N_18180,N_7519,N_6793);
xnor U18181 (N_18181,N_6399,N_10309);
nand U18182 (N_18182,N_7933,N_8098);
nor U18183 (N_18183,N_7019,N_11270);
xor U18184 (N_18184,N_8723,N_7443);
nor U18185 (N_18185,N_6502,N_11816);
or U18186 (N_18186,N_7932,N_6621);
and U18187 (N_18187,N_9424,N_12386);
or U18188 (N_18188,N_7927,N_9235);
nand U18189 (N_18189,N_10247,N_9922);
nor U18190 (N_18190,N_12435,N_11830);
or U18191 (N_18191,N_6653,N_11077);
xor U18192 (N_18192,N_8968,N_6942);
or U18193 (N_18193,N_12427,N_9344);
or U18194 (N_18194,N_10876,N_12306);
nand U18195 (N_18195,N_6752,N_8892);
nand U18196 (N_18196,N_10241,N_10482);
xnor U18197 (N_18197,N_9987,N_12234);
xnor U18198 (N_18198,N_9518,N_6392);
nand U18199 (N_18199,N_8652,N_10758);
xnor U18200 (N_18200,N_8611,N_7699);
xnor U18201 (N_18201,N_7736,N_10684);
xnor U18202 (N_18202,N_9287,N_11760);
and U18203 (N_18203,N_10582,N_9440);
nor U18204 (N_18204,N_12160,N_7606);
nand U18205 (N_18205,N_11135,N_6304);
nand U18206 (N_18206,N_11754,N_10787);
xnor U18207 (N_18207,N_11090,N_9294);
nand U18208 (N_18208,N_11113,N_9816);
and U18209 (N_18209,N_11643,N_7127);
nand U18210 (N_18210,N_9160,N_11096);
and U18211 (N_18211,N_8549,N_11903);
or U18212 (N_18212,N_8173,N_6270);
or U18213 (N_18213,N_6723,N_11872);
and U18214 (N_18214,N_11358,N_10594);
nand U18215 (N_18215,N_9598,N_10363);
xnor U18216 (N_18216,N_7506,N_7731);
or U18217 (N_18217,N_6324,N_7522);
nand U18218 (N_18218,N_10572,N_10812);
and U18219 (N_18219,N_7271,N_9449);
and U18220 (N_18220,N_6691,N_9524);
and U18221 (N_18221,N_7382,N_10048);
nand U18222 (N_18222,N_9479,N_8239);
or U18223 (N_18223,N_11698,N_10876);
nor U18224 (N_18224,N_10631,N_7508);
nand U18225 (N_18225,N_7896,N_10551);
nand U18226 (N_18226,N_12248,N_12025);
xnor U18227 (N_18227,N_12092,N_9619);
or U18228 (N_18228,N_12126,N_8414);
or U18229 (N_18229,N_11109,N_8754);
nand U18230 (N_18230,N_7110,N_10989);
nand U18231 (N_18231,N_10893,N_12304);
nor U18232 (N_18232,N_8318,N_8374);
nor U18233 (N_18233,N_6371,N_8829);
and U18234 (N_18234,N_9021,N_10217);
nand U18235 (N_18235,N_11284,N_9160);
or U18236 (N_18236,N_7109,N_12303);
and U18237 (N_18237,N_9276,N_8635);
or U18238 (N_18238,N_10581,N_10607);
or U18239 (N_18239,N_8553,N_11952);
nor U18240 (N_18240,N_6827,N_10316);
and U18241 (N_18241,N_8331,N_10324);
xor U18242 (N_18242,N_12391,N_10582);
nand U18243 (N_18243,N_10613,N_9605);
nand U18244 (N_18244,N_12446,N_7012);
nor U18245 (N_18245,N_6388,N_6646);
xnor U18246 (N_18246,N_10568,N_6405);
or U18247 (N_18247,N_10701,N_12431);
nand U18248 (N_18248,N_7632,N_11123);
and U18249 (N_18249,N_10288,N_10212);
nor U18250 (N_18250,N_10785,N_11086);
nor U18251 (N_18251,N_7595,N_12034);
or U18252 (N_18252,N_10380,N_10021);
nor U18253 (N_18253,N_9921,N_7627);
xnor U18254 (N_18254,N_8024,N_9823);
xnor U18255 (N_18255,N_8156,N_8553);
or U18256 (N_18256,N_7853,N_7741);
nor U18257 (N_18257,N_8087,N_10021);
nor U18258 (N_18258,N_10304,N_7537);
nor U18259 (N_18259,N_10152,N_10291);
and U18260 (N_18260,N_11261,N_8391);
nor U18261 (N_18261,N_9002,N_6593);
and U18262 (N_18262,N_7082,N_12232);
or U18263 (N_18263,N_7696,N_9960);
nand U18264 (N_18264,N_11053,N_7054);
nand U18265 (N_18265,N_9363,N_7308);
nor U18266 (N_18266,N_9728,N_10874);
xor U18267 (N_18267,N_7397,N_6471);
or U18268 (N_18268,N_7344,N_8966);
nand U18269 (N_18269,N_7794,N_9122);
nor U18270 (N_18270,N_8620,N_10437);
nand U18271 (N_18271,N_8061,N_9298);
or U18272 (N_18272,N_11403,N_10931);
or U18273 (N_18273,N_7705,N_10812);
and U18274 (N_18274,N_10817,N_11676);
nor U18275 (N_18275,N_8754,N_12341);
xnor U18276 (N_18276,N_10441,N_9266);
or U18277 (N_18277,N_9095,N_7155);
nor U18278 (N_18278,N_9523,N_11172);
and U18279 (N_18279,N_8431,N_7343);
xor U18280 (N_18280,N_10009,N_10784);
nand U18281 (N_18281,N_8329,N_6286);
nand U18282 (N_18282,N_10843,N_9115);
nand U18283 (N_18283,N_11472,N_12257);
nand U18284 (N_18284,N_11232,N_11264);
nand U18285 (N_18285,N_7784,N_12185);
or U18286 (N_18286,N_7936,N_11132);
nand U18287 (N_18287,N_6386,N_7667);
xor U18288 (N_18288,N_6411,N_12172);
xnor U18289 (N_18289,N_10343,N_8087);
nand U18290 (N_18290,N_7295,N_11999);
nor U18291 (N_18291,N_11378,N_10200);
and U18292 (N_18292,N_9821,N_11998);
and U18293 (N_18293,N_11226,N_9899);
xnor U18294 (N_18294,N_9657,N_11208);
nor U18295 (N_18295,N_8887,N_8131);
and U18296 (N_18296,N_7516,N_7145);
nand U18297 (N_18297,N_9464,N_11408);
or U18298 (N_18298,N_7270,N_11689);
xor U18299 (N_18299,N_12460,N_6522);
nand U18300 (N_18300,N_8267,N_12364);
or U18301 (N_18301,N_11671,N_8074);
nor U18302 (N_18302,N_6755,N_11836);
nand U18303 (N_18303,N_11039,N_11018);
nor U18304 (N_18304,N_9345,N_11568);
xor U18305 (N_18305,N_6324,N_9952);
and U18306 (N_18306,N_10925,N_9945);
nor U18307 (N_18307,N_9101,N_9343);
xnor U18308 (N_18308,N_10143,N_8020);
nand U18309 (N_18309,N_8937,N_6299);
xor U18310 (N_18310,N_6326,N_10553);
nor U18311 (N_18311,N_8720,N_10823);
and U18312 (N_18312,N_10835,N_7139);
xnor U18313 (N_18313,N_11577,N_9842);
nor U18314 (N_18314,N_6622,N_6608);
or U18315 (N_18315,N_8309,N_11010);
xnor U18316 (N_18316,N_10846,N_11515);
xor U18317 (N_18317,N_8579,N_7459);
nand U18318 (N_18318,N_9612,N_9608);
and U18319 (N_18319,N_11265,N_6704);
nand U18320 (N_18320,N_6803,N_7195);
nand U18321 (N_18321,N_8446,N_8055);
xnor U18322 (N_18322,N_12498,N_7057);
nor U18323 (N_18323,N_10730,N_7244);
xor U18324 (N_18324,N_11198,N_11604);
or U18325 (N_18325,N_9172,N_11575);
nor U18326 (N_18326,N_7441,N_7651);
nor U18327 (N_18327,N_9556,N_9234);
xnor U18328 (N_18328,N_9233,N_12357);
nand U18329 (N_18329,N_9439,N_9596);
xnor U18330 (N_18330,N_9767,N_9854);
xor U18331 (N_18331,N_11601,N_10767);
nor U18332 (N_18332,N_6476,N_10933);
and U18333 (N_18333,N_10515,N_11746);
and U18334 (N_18334,N_11305,N_7764);
nand U18335 (N_18335,N_9132,N_11400);
nor U18336 (N_18336,N_12231,N_7777);
or U18337 (N_18337,N_12238,N_9320);
nand U18338 (N_18338,N_6972,N_11722);
xnor U18339 (N_18339,N_7153,N_8090);
xnor U18340 (N_18340,N_7265,N_10703);
nand U18341 (N_18341,N_9625,N_11183);
and U18342 (N_18342,N_7975,N_10787);
xnor U18343 (N_18343,N_7102,N_6318);
nand U18344 (N_18344,N_12285,N_6876);
xor U18345 (N_18345,N_10062,N_12052);
nor U18346 (N_18346,N_6688,N_10861);
nand U18347 (N_18347,N_8326,N_8599);
nand U18348 (N_18348,N_9095,N_7130);
xnor U18349 (N_18349,N_10891,N_7867);
and U18350 (N_18350,N_6872,N_6297);
nand U18351 (N_18351,N_12400,N_12464);
xor U18352 (N_18352,N_10867,N_8159);
nor U18353 (N_18353,N_8419,N_7640);
nand U18354 (N_18354,N_9490,N_8782);
and U18355 (N_18355,N_7731,N_11429);
nand U18356 (N_18356,N_6835,N_9830);
and U18357 (N_18357,N_10270,N_6595);
nand U18358 (N_18358,N_10046,N_8206);
nand U18359 (N_18359,N_11289,N_6549);
nand U18360 (N_18360,N_10050,N_8440);
nand U18361 (N_18361,N_7121,N_12078);
nor U18362 (N_18362,N_8843,N_8846);
xnor U18363 (N_18363,N_6978,N_10874);
nand U18364 (N_18364,N_7639,N_9573);
xnor U18365 (N_18365,N_7058,N_12148);
xnor U18366 (N_18366,N_10790,N_6322);
and U18367 (N_18367,N_12256,N_6443);
xor U18368 (N_18368,N_12141,N_9200);
and U18369 (N_18369,N_12182,N_11938);
or U18370 (N_18370,N_6883,N_10576);
nor U18371 (N_18371,N_7278,N_8212);
nand U18372 (N_18372,N_7898,N_8287);
xor U18373 (N_18373,N_6679,N_9981);
nor U18374 (N_18374,N_6521,N_7042);
nand U18375 (N_18375,N_10654,N_6449);
xnor U18376 (N_18376,N_11442,N_10105);
and U18377 (N_18377,N_9245,N_8690);
nor U18378 (N_18378,N_6528,N_7086);
and U18379 (N_18379,N_6538,N_10186);
xor U18380 (N_18380,N_6336,N_7238);
nor U18381 (N_18381,N_8597,N_9956);
or U18382 (N_18382,N_12439,N_8254);
and U18383 (N_18383,N_6408,N_10631);
or U18384 (N_18384,N_12277,N_7101);
nand U18385 (N_18385,N_10297,N_8090);
xnor U18386 (N_18386,N_11592,N_9927);
nand U18387 (N_18387,N_6330,N_6515);
nand U18388 (N_18388,N_9703,N_9249);
xnor U18389 (N_18389,N_8156,N_6396);
xnor U18390 (N_18390,N_7315,N_9164);
and U18391 (N_18391,N_11367,N_9113);
and U18392 (N_18392,N_12343,N_11764);
xnor U18393 (N_18393,N_6342,N_11484);
nor U18394 (N_18394,N_8000,N_6481);
or U18395 (N_18395,N_7733,N_8538);
nor U18396 (N_18396,N_12370,N_7211);
nand U18397 (N_18397,N_9035,N_9205);
nor U18398 (N_18398,N_7941,N_9745);
xor U18399 (N_18399,N_9418,N_7372);
xor U18400 (N_18400,N_7583,N_7310);
and U18401 (N_18401,N_11557,N_11818);
nor U18402 (N_18402,N_11583,N_6327);
nor U18403 (N_18403,N_7573,N_11509);
xnor U18404 (N_18404,N_10150,N_12469);
nand U18405 (N_18405,N_9009,N_9825);
and U18406 (N_18406,N_10397,N_6609);
or U18407 (N_18407,N_7103,N_12177);
or U18408 (N_18408,N_8811,N_6834);
xor U18409 (N_18409,N_7402,N_8636);
and U18410 (N_18410,N_10792,N_11565);
nand U18411 (N_18411,N_12441,N_10720);
nor U18412 (N_18412,N_12002,N_6489);
nor U18413 (N_18413,N_11779,N_6446);
nor U18414 (N_18414,N_11470,N_7494);
nand U18415 (N_18415,N_11611,N_12418);
nor U18416 (N_18416,N_6807,N_11991);
or U18417 (N_18417,N_10786,N_12149);
or U18418 (N_18418,N_7699,N_12078);
nand U18419 (N_18419,N_7150,N_7122);
and U18420 (N_18420,N_10123,N_11398);
nor U18421 (N_18421,N_10697,N_9933);
or U18422 (N_18422,N_12086,N_11537);
nand U18423 (N_18423,N_8861,N_10512);
and U18424 (N_18424,N_11705,N_7968);
or U18425 (N_18425,N_9748,N_8030);
xor U18426 (N_18426,N_10554,N_6624);
xor U18427 (N_18427,N_6327,N_9154);
nand U18428 (N_18428,N_10347,N_11782);
and U18429 (N_18429,N_11924,N_10052);
nand U18430 (N_18430,N_6831,N_10278);
nand U18431 (N_18431,N_8991,N_10590);
nor U18432 (N_18432,N_7166,N_10317);
nor U18433 (N_18433,N_8103,N_7834);
nor U18434 (N_18434,N_7083,N_9030);
and U18435 (N_18435,N_9484,N_9446);
xor U18436 (N_18436,N_9486,N_11355);
and U18437 (N_18437,N_8926,N_9440);
nor U18438 (N_18438,N_10796,N_12261);
or U18439 (N_18439,N_6725,N_6890);
nor U18440 (N_18440,N_7938,N_8090);
and U18441 (N_18441,N_11523,N_10930);
or U18442 (N_18442,N_8248,N_6894);
or U18443 (N_18443,N_7204,N_8291);
xnor U18444 (N_18444,N_8241,N_6790);
xor U18445 (N_18445,N_8560,N_11338);
nand U18446 (N_18446,N_6526,N_11784);
nor U18447 (N_18447,N_9945,N_10494);
or U18448 (N_18448,N_10059,N_8509);
xnor U18449 (N_18449,N_8898,N_7572);
nand U18450 (N_18450,N_12148,N_8681);
nand U18451 (N_18451,N_9152,N_9716);
and U18452 (N_18452,N_11611,N_7913);
xnor U18453 (N_18453,N_6615,N_11358);
or U18454 (N_18454,N_7326,N_7517);
nand U18455 (N_18455,N_9194,N_10394);
nor U18456 (N_18456,N_11521,N_9932);
nand U18457 (N_18457,N_7876,N_7711);
nor U18458 (N_18458,N_9485,N_11440);
nor U18459 (N_18459,N_12461,N_9537);
nand U18460 (N_18460,N_7752,N_10130);
nor U18461 (N_18461,N_9728,N_7744);
nor U18462 (N_18462,N_7067,N_11502);
or U18463 (N_18463,N_10349,N_8096);
xnor U18464 (N_18464,N_10815,N_6361);
nor U18465 (N_18465,N_6362,N_12353);
and U18466 (N_18466,N_8707,N_8027);
and U18467 (N_18467,N_10702,N_6830);
xor U18468 (N_18468,N_11780,N_10901);
xor U18469 (N_18469,N_10528,N_8970);
or U18470 (N_18470,N_8679,N_10415);
nand U18471 (N_18471,N_11396,N_11238);
nor U18472 (N_18472,N_9544,N_8031);
or U18473 (N_18473,N_9922,N_6339);
or U18474 (N_18474,N_6479,N_9721);
nor U18475 (N_18475,N_6561,N_8048);
xor U18476 (N_18476,N_7634,N_8750);
nand U18477 (N_18477,N_6270,N_10957);
and U18478 (N_18478,N_12189,N_7314);
xor U18479 (N_18479,N_7496,N_10986);
nand U18480 (N_18480,N_6329,N_12439);
or U18481 (N_18481,N_8358,N_12210);
or U18482 (N_18482,N_8583,N_11297);
nand U18483 (N_18483,N_9418,N_10620);
or U18484 (N_18484,N_12298,N_11583);
xnor U18485 (N_18485,N_12153,N_6257);
and U18486 (N_18486,N_10215,N_8994);
nand U18487 (N_18487,N_8177,N_8907);
and U18488 (N_18488,N_8612,N_8055);
and U18489 (N_18489,N_8560,N_10478);
and U18490 (N_18490,N_9425,N_7884);
xnor U18491 (N_18491,N_11520,N_12147);
nor U18492 (N_18492,N_6439,N_6495);
xor U18493 (N_18493,N_9405,N_9890);
or U18494 (N_18494,N_9669,N_8483);
and U18495 (N_18495,N_11645,N_11327);
nor U18496 (N_18496,N_10217,N_8868);
or U18497 (N_18497,N_11001,N_6698);
nor U18498 (N_18498,N_6599,N_12322);
nor U18499 (N_18499,N_12133,N_9670);
nand U18500 (N_18500,N_6411,N_8169);
xnor U18501 (N_18501,N_6726,N_11698);
or U18502 (N_18502,N_9986,N_8234);
and U18503 (N_18503,N_8689,N_10073);
nor U18504 (N_18504,N_10943,N_6351);
and U18505 (N_18505,N_6549,N_7906);
xnor U18506 (N_18506,N_12367,N_7260);
or U18507 (N_18507,N_6795,N_7944);
nor U18508 (N_18508,N_7482,N_9635);
xor U18509 (N_18509,N_7679,N_8055);
and U18510 (N_18510,N_10978,N_10399);
nor U18511 (N_18511,N_11046,N_7869);
nand U18512 (N_18512,N_9544,N_8367);
nor U18513 (N_18513,N_11812,N_9488);
or U18514 (N_18514,N_7630,N_6419);
nand U18515 (N_18515,N_9074,N_7642);
xnor U18516 (N_18516,N_6944,N_9478);
xnor U18517 (N_18517,N_10886,N_8637);
and U18518 (N_18518,N_7610,N_6899);
nand U18519 (N_18519,N_10511,N_11530);
and U18520 (N_18520,N_11263,N_7836);
nand U18521 (N_18521,N_12402,N_12256);
or U18522 (N_18522,N_10504,N_7529);
nor U18523 (N_18523,N_12094,N_7611);
xor U18524 (N_18524,N_8355,N_9310);
and U18525 (N_18525,N_10206,N_8326);
xor U18526 (N_18526,N_8989,N_8181);
or U18527 (N_18527,N_7693,N_11634);
nor U18528 (N_18528,N_8697,N_10315);
nand U18529 (N_18529,N_9558,N_10709);
and U18530 (N_18530,N_10792,N_9609);
or U18531 (N_18531,N_8983,N_10697);
xor U18532 (N_18532,N_10966,N_11862);
xnor U18533 (N_18533,N_9459,N_7636);
nand U18534 (N_18534,N_9070,N_11476);
and U18535 (N_18535,N_11472,N_9192);
xnor U18536 (N_18536,N_8604,N_8301);
or U18537 (N_18537,N_8512,N_6576);
or U18538 (N_18538,N_11194,N_8452);
or U18539 (N_18539,N_9571,N_7493);
and U18540 (N_18540,N_6436,N_6296);
nand U18541 (N_18541,N_11438,N_9173);
or U18542 (N_18542,N_12482,N_8728);
nor U18543 (N_18543,N_8249,N_6535);
xnor U18544 (N_18544,N_8560,N_10162);
nor U18545 (N_18545,N_6870,N_11145);
and U18546 (N_18546,N_11468,N_6867);
nor U18547 (N_18547,N_8653,N_7100);
nor U18548 (N_18548,N_10195,N_10878);
or U18549 (N_18549,N_7012,N_7484);
and U18550 (N_18550,N_8804,N_6732);
and U18551 (N_18551,N_7938,N_9237);
or U18552 (N_18552,N_8174,N_10564);
and U18553 (N_18553,N_10056,N_8088);
nand U18554 (N_18554,N_8166,N_7544);
nor U18555 (N_18555,N_8722,N_8443);
nor U18556 (N_18556,N_12347,N_6379);
xor U18557 (N_18557,N_7417,N_6817);
nor U18558 (N_18558,N_10291,N_12241);
and U18559 (N_18559,N_7009,N_6274);
nor U18560 (N_18560,N_11397,N_10103);
nor U18561 (N_18561,N_11325,N_12293);
nor U18562 (N_18562,N_12117,N_8989);
xor U18563 (N_18563,N_12439,N_7996);
nor U18564 (N_18564,N_10554,N_10206);
and U18565 (N_18565,N_11963,N_10669);
or U18566 (N_18566,N_12441,N_6588);
nand U18567 (N_18567,N_7490,N_8368);
xor U18568 (N_18568,N_6407,N_9350);
or U18569 (N_18569,N_7680,N_9245);
and U18570 (N_18570,N_7653,N_9927);
and U18571 (N_18571,N_9877,N_8767);
nor U18572 (N_18572,N_10046,N_7498);
xnor U18573 (N_18573,N_9808,N_11014);
or U18574 (N_18574,N_7259,N_6758);
or U18575 (N_18575,N_12104,N_11245);
xnor U18576 (N_18576,N_12139,N_7863);
and U18577 (N_18577,N_12153,N_8959);
nor U18578 (N_18578,N_11129,N_8307);
nor U18579 (N_18579,N_11949,N_11357);
xor U18580 (N_18580,N_9481,N_6411);
or U18581 (N_18581,N_6613,N_10752);
or U18582 (N_18582,N_12287,N_11169);
nand U18583 (N_18583,N_12130,N_8492);
and U18584 (N_18584,N_6787,N_11210);
and U18585 (N_18585,N_8837,N_6309);
nand U18586 (N_18586,N_6321,N_11484);
nor U18587 (N_18587,N_6432,N_11169);
nor U18588 (N_18588,N_12387,N_12401);
nor U18589 (N_18589,N_7145,N_8034);
nor U18590 (N_18590,N_7576,N_7448);
and U18591 (N_18591,N_10472,N_11053);
xor U18592 (N_18592,N_7279,N_9352);
or U18593 (N_18593,N_12129,N_6523);
nor U18594 (N_18594,N_7729,N_11246);
nand U18595 (N_18595,N_9121,N_7655);
nand U18596 (N_18596,N_10130,N_12418);
and U18597 (N_18597,N_11409,N_8429);
or U18598 (N_18598,N_6427,N_7170);
or U18599 (N_18599,N_11012,N_10667);
nor U18600 (N_18600,N_9275,N_8426);
or U18601 (N_18601,N_7157,N_6937);
xnor U18602 (N_18602,N_11473,N_8889);
and U18603 (N_18603,N_10238,N_9262);
xnor U18604 (N_18604,N_6393,N_6400);
or U18605 (N_18605,N_10957,N_10660);
nand U18606 (N_18606,N_6860,N_8804);
nor U18607 (N_18607,N_8581,N_9505);
and U18608 (N_18608,N_6291,N_6904);
and U18609 (N_18609,N_11479,N_8072);
or U18610 (N_18610,N_11836,N_6605);
and U18611 (N_18611,N_11118,N_12015);
and U18612 (N_18612,N_7400,N_7499);
nor U18613 (N_18613,N_12407,N_10125);
nand U18614 (N_18614,N_10652,N_11042);
xnor U18615 (N_18615,N_10597,N_11589);
nor U18616 (N_18616,N_8470,N_6612);
nor U18617 (N_18617,N_6440,N_6766);
or U18618 (N_18618,N_11636,N_10436);
and U18619 (N_18619,N_10057,N_8252);
nand U18620 (N_18620,N_8956,N_9737);
xor U18621 (N_18621,N_6400,N_8638);
and U18622 (N_18622,N_12220,N_6714);
nor U18623 (N_18623,N_7328,N_10154);
xor U18624 (N_18624,N_9199,N_11973);
nor U18625 (N_18625,N_7505,N_11249);
or U18626 (N_18626,N_10554,N_10241);
xnor U18627 (N_18627,N_11408,N_10684);
and U18628 (N_18628,N_11105,N_11534);
nand U18629 (N_18629,N_10217,N_7692);
xnor U18630 (N_18630,N_9620,N_12484);
xor U18631 (N_18631,N_9015,N_7817);
and U18632 (N_18632,N_12286,N_7115);
or U18633 (N_18633,N_10431,N_9335);
and U18634 (N_18634,N_9261,N_12377);
nor U18635 (N_18635,N_7267,N_8866);
xnor U18636 (N_18636,N_11305,N_8755);
and U18637 (N_18637,N_9381,N_11710);
nand U18638 (N_18638,N_8119,N_11953);
nor U18639 (N_18639,N_11459,N_10512);
xor U18640 (N_18640,N_6835,N_6356);
nand U18641 (N_18641,N_7978,N_12071);
nor U18642 (N_18642,N_10862,N_10620);
nor U18643 (N_18643,N_7951,N_6309);
xnor U18644 (N_18644,N_8644,N_7727);
nor U18645 (N_18645,N_8850,N_7772);
or U18646 (N_18646,N_9724,N_12075);
or U18647 (N_18647,N_9617,N_10388);
and U18648 (N_18648,N_8154,N_8176);
nor U18649 (N_18649,N_9963,N_10600);
nand U18650 (N_18650,N_6762,N_10704);
xor U18651 (N_18651,N_7266,N_9949);
nor U18652 (N_18652,N_6413,N_9656);
and U18653 (N_18653,N_9527,N_8574);
or U18654 (N_18654,N_8946,N_6605);
nor U18655 (N_18655,N_7720,N_7904);
nand U18656 (N_18656,N_10139,N_11166);
nand U18657 (N_18657,N_8904,N_8926);
and U18658 (N_18658,N_10392,N_7740);
nand U18659 (N_18659,N_9833,N_8487);
and U18660 (N_18660,N_9319,N_10315);
nor U18661 (N_18661,N_9142,N_8805);
nand U18662 (N_18662,N_8381,N_11427);
or U18663 (N_18663,N_8376,N_7456);
or U18664 (N_18664,N_6385,N_11729);
nor U18665 (N_18665,N_7817,N_10452);
nand U18666 (N_18666,N_11490,N_7287);
and U18667 (N_18667,N_8496,N_7299);
and U18668 (N_18668,N_8271,N_8478);
or U18669 (N_18669,N_6427,N_8250);
nand U18670 (N_18670,N_8963,N_11434);
or U18671 (N_18671,N_12198,N_8422);
xor U18672 (N_18672,N_9260,N_9898);
nand U18673 (N_18673,N_7090,N_7707);
and U18674 (N_18674,N_6425,N_11870);
or U18675 (N_18675,N_11544,N_11390);
nand U18676 (N_18676,N_11340,N_7821);
xor U18677 (N_18677,N_8327,N_11141);
and U18678 (N_18678,N_8329,N_11638);
and U18679 (N_18679,N_6665,N_11050);
and U18680 (N_18680,N_7435,N_11371);
nor U18681 (N_18681,N_10735,N_8972);
and U18682 (N_18682,N_12188,N_7327);
or U18683 (N_18683,N_9451,N_12153);
xor U18684 (N_18684,N_9714,N_7629);
or U18685 (N_18685,N_11030,N_9892);
xnor U18686 (N_18686,N_7933,N_7296);
xor U18687 (N_18687,N_12249,N_10439);
nor U18688 (N_18688,N_8838,N_6706);
or U18689 (N_18689,N_6737,N_8896);
or U18690 (N_18690,N_9584,N_8013);
and U18691 (N_18691,N_8030,N_6677);
nor U18692 (N_18692,N_9333,N_11967);
or U18693 (N_18693,N_9078,N_8773);
or U18694 (N_18694,N_10928,N_9767);
or U18695 (N_18695,N_9373,N_7376);
and U18696 (N_18696,N_7613,N_12072);
nand U18697 (N_18697,N_12183,N_7792);
xor U18698 (N_18698,N_10886,N_10347);
nor U18699 (N_18699,N_8012,N_9821);
nand U18700 (N_18700,N_6801,N_6626);
nor U18701 (N_18701,N_9697,N_10611);
and U18702 (N_18702,N_8530,N_7011);
xor U18703 (N_18703,N_9407,N_7972);
nor U18704 (N_18704,N_9337,N_12047);
or U18705 (N_18705,N_8761,N_6255);
or U18706 (N_18706,N_8476,N_8747);
nor U18707 (N_18707,N_10752,N_9498);
nand U18708 (N_18708,N_8298,N_9826);
nand U18709 (N_18709,N_10101,N_10724);
nand U18710 (N_18710,N_10404,N_10917);
nand U18711 (N_18711,N_10547,N_10932);
nor U18712 (N_18712,N_12181,N_6549);
and U18713 (N_18713,N_6387,N_8487);
and U18714 (N_18714,N_10555,N_7457);
nand U18715 (N_18715,N_8798,N_12440);
nor U18716 (N_18716,N_10857,N_12000);
or U18717 (N_18717,N_12006,N_7706);
or U18718 (N_18718,N_7704,N_7946);
and U18719 (N_18719,N_6660,N_11500);
xnor U18720 (N_18720,N_10847,N_7610);
xnor U18721 (N_18721,N_11860,N_10605);
nor U18722 (N_18722,N_8838,N_10197);
nor U18723 (N_18723,N_10803,N_9373);
xor U18724 (N_18724,N_6340,N_8047);
xnor U18725 (N_18725,N_10092,N_8941);
nor U18726 (N_18726,N_7762,N_9294);
and U18727 (N_18727,N_12211,N_9128);
or U18728 (N_18728,N_7355,N_11789);
nor U18729 (N_18729,N_8635,N_6525);
xnor U18730 (N_18730,N_7057,N_11418);
xnor U18731 (N_18731,N_9977,N_7014);
nand U18732 (N_18732,N_10316,N_9726);
nand U18733 (N_18733,N_12116,N_7513);
or U18734 (N_18734,N_10397,N_8448);
nand U18735 (N_18735,N_9428,N_11109);
or U18736 (N_18736,N_6387,N_6867);
and U18737 (N_18737,N_12135,N_6542);
or U18738 (N_18738,N_7251,N_8186);
or U18739 (N_18739,N_9634,N_11038);
and U18740 (N_18740,N_9778,N_8950);
nand U18741 (N_18741,N_10051,N_6681);
nand U18742 (N_18742,N_11949,N_11200);
and U18743 (N_18743,N_10059,N_11488);
nor U18744 (N_18744,N_9697,N_8529);
and U18745 (N_18745,N_11815,N_6932);
xnor U18746 (N_18746,N_10017,N_9320);
nor U18747 (N_18747,N_10213,N_6439);
xor U18748 (N_18748,N_11558,N_12131);
nand U18749 (N_18749,N_7512,N_8969);
nand U18750 (N_18750,N_17088,N_16979);
xor U18751 (N_18751,N_14939,N_15129);
nand U18752 (N_18752,N_16398,N_18112);
nor U18753 (N_18753,N_14624,N_17729);
xor U18754 (N_18754,N_17249,N_17252);
or U18755 (N_18755,N_14107,N_15196);
xor U18756 (N_18756,N_13226,N_14923);
xnor U18757 (N_18757,N_16717,N_17938);
nor U18758 (N_18758,N_13670,N_14253);
or U18759 (N_18759,N_15654,N_16213);
and U18760 (N_18760,N_15607,N_14728);
nor U18761 (N_18761,N_14057,N_12759);
nor U18762 (N_18762,N_17797,N_16957);
xnor U18763 (N_18763,N_16329,N_18736);
xor U18764 (N_18764,N_18268,N_17479);
and U18765 (N_18765,N_17773,N_18175);
and U18766 (N_18766,N_16987,N_17518);
nand U18767 (N_18767,N_18407,N_14128);
or U18768 (N_18768,N_17258,N_14602);
or U18769 (N_18769,N_12790,N_13002);
nor U18770 (N_18770,N_17863,N_12646);
and U18771 (N_18771,N_14342,N_17717);
xnor U18772 (N_18772,N_13339,N_12730);
nor U18773 (N_18773,N_17512,N_12742);
and U18774 (N_18774,N_12532,N_14955);
nor U18775 (N_18775,N_17255,N_17861);
xnor U18776 (N_18776,N_15232,N_15724);
and U18777 (N_18777,N_12628,N_14269);
nor U18778 (N_18778,N_15145,N_13520);
xnor U18779 (N_18779,N_17668,N_16027);
xor U18780 (N_18780,N_17999,N_14983);
and U18781 (N_18781,N_18267,N_15161);
nand U18782 (N_18782,N_14320,N_13535);
nor U18783 (N_18783,N_16395,N_16931);
xor U18784 (N_18784,N_13634,N_13692);
and U18785 (N_18785,N_14291,N_15311);
nand U18786 (N_18786,N_17800,N_17403);
xnor U18787 (N_18787,N_13401,N_16089);
nor U18788 (N_18788,N_16558,N_16664);
or U18789 (N_18789,N_17264,N_15316);
and U18790 (N_18790,N_16454,N_15868);
nand U18791 (N_18791,N_17596,N_17468);
nor U18792 (N_18792,N_18490,N_14875);
nor U18793 (N_18793,N_18003,N_12666);
or U18794 (N_18794,N_13583,N_12756);
or U18795 (N_18795,N_17884,N_12729);
or U18796 (N_18796,N_13764,N_18563);
xnor U18797 (N_18797,N_15584,N_18403);
nand U18798 (N_18798,N_14447,N_13828);
nor U18799 (N_18799,N_13126,N_18091);
nor U18800 (N_18800,N_17948,N_18246);
nor U18801 (N_18801,N_15136,N_13526);
and U18802 (N_18802,N_14858,N_13131);
xnor U18803 (N_18803,N_17516,N_17913);
and U18804 (N_18804,N_14750,N_12866);
xor U18805 (N_18805,N_17080,N_18012);
xnor U18806 (N_18806,N_13539,N_13079);
nor U18807 (N_18807,N_17296,N_13537);
nor U18808 (N_18808,N_14257,N_16673);
or U18809 (N_18809,N_15665,N_18644);
xor U18810 (N_18810,N_13811,N_14483);
nor U18811 (N_18811,N_15670,N_14190);
or U18812 (N_18812,N_16981,N_17779);
xnor U18813 (N_18813,N_14941,N_15380);
xor U18814 (N_18814,N_13358,N_16726);
xnor U18815 (N_18815,N_16426,N_18000);
and U18816 (N_18816,N_13864,N_15237);
or U18817 (N_18817,N_12837,N_17290);
or U18818 (N_18818,N_13902,N_16016);
nand U18819 (N_18819,N_15191,N_16070);
xnor U18820 (N_18820,N_14663,N_15532);
xnor U18821 (N_18821,N_13708,N_13296);
nor U18822 (N_18822,N_16382,N_12961);
or U18823 (N_18823,N_13819,N_18711);
or U18824 (N_18824,N_13375,N_14244);
xnor U18825 (N_18825,N_13865,N_14432);
nor U18826 (N_18826,N_16134,N_17337);
and U18827 (N_18827,N_13672,N_13363);
xnor U18828 (N_18828,N_16668,N_15011);
or U18829 (N_18829,N_18600,N_15771);
xor U18830 (N_18830,N_14300,N_13356);
and U18831 (N_18831,N_16391,N_12537);
or U18832 (N_18832,N_13313,N_16681);
nor U18833 (N_18833,N_16674,N_13372);
nor U18834 (N_18834,N_14702,N_18180);
and U18835 (N_18835,N_14917,N_13745);
nor U18836 (N_18836,N_17905,N_13561);
and U18837 (N_18837,N_12772,N_18245);
and U18838 (N_18838,N_18052,N_15101);
and U18839 (N_18839,N_15408,N_15583);
nand U18840 (N_18840,N_17236,N_16119);
nand U18841 (N_18841,N_13306,N_14112);
and U18842 (N_18842,N_14333,N_15080);
xor U18843 (N_18843,N_18122,N_18241);
and U18844 (N_18844,N_15546,N_15928);
and U18845 (N_18845,N_17679,N_14593);
nand U18846 (N_18846,N_18418,N_12768);
or U18847 (N_18847,N_15178,N_12873);
nor U18848 (N_18848,N_15201,N_18040);
xnor U18849 (N_18849,N_17416,N_16340);
and U18850 (N_18850,N_12807,N_14867);
nand U18851 (N_18851,N_17650,N_16909);
nor U18852 (N_18852,N_18062,N_18461);
nor U18853 (N_18853,N_13582,N_13014);
nor U18854 (N_18854,N_17764,N_13281);
and U18855 (N_18855,N_14589,N_15609);
xor U18856 (N_18856,N_13930,N_16706);
and U18857 (N_18857,N_14059,N_13450);
and U18858 (N_18858,N_14938,N_12500);
nand U18859 (N_18859,N_18748,N_17231);
or U18860 (N_18860,N_15705,N_18692);
xnor U18861 (N_18861,N_15298,N_13996);
nand U18862 (N_18862,N_17825,N_12641);
nor U18863 (N_18863,N_12891,N_14101);
and U18864 (N_18864,N_12607,N_17611);
nor U18865 (N_18865,N_18088,N_17995);
and U18866 (N_18866,N_12985,N_15171);
or U18867 (N_18867,N_12561,N_18255);
xnor U18868 (N_18868,N_13743,N_16182);
xor U18869 (N_18869,N_18445,N_18363);
xor U18870 (N_18870,N_12517,N_14007);
or U18871 (N_18871,N_17306,N_17633);
nand U18872 (N_18872,N_13758,N_17034);
or U18873 (N_18873,N_15776,N_12982);
nand U18874 (N_18874,N_18610,N_14371);
and U18875 (N_18875,N_16373,N_12906);
or U18876 (N_18876,N_18511,N_13509);
nand U18877 (N_18877,N_18683,N_17918);
xnor U18878 (N_18878,N_18675,N_14000);
xnor U18879 (N_18879,N_15401,N_12962);
and U18880 (N_18880,N_14523,N_16015);
nor U18881 (N_18881,N_17104,N_14228);
xnor U18882 (N_18882,N_16460,N_14977);
nor U18883 (N_18883,N_16291,N_15498);
nand U18884 (N_18884,N_14123,N_13525);
nor U18885 (N_18885,N_14219,N_18450);
or U18886 (N_18886,N_16445,N_18048);
or U18887 (N_18887,N_15436,N_17666);
or U18888 (N_18888,N_15787,N_15400);
or U18889 (N_18889,N_16366,N_17720);
nand U18890 (N_18890,N_14175,N_14402);
and U18891 (N_18891,N_13760,N_17979);
and U18892 (N_18892,N_14405,N_13072);
nor U18893 (N_18893,N_13353,N_17068);
xor U18894 (N_18894,N_15122,N_17838);
or U18895 (N_18895,N_17911,N_17124);
xor U18896 (N_18896,N_13705,N_18194);
nand U18897 (N_18897,N_12663,N_13010);
nor U18898 (N_18898,N_12806,N_14408);
xor U18899 (N_18899,N_16954,N_16171);
or U18900 (N_18900,N_17853,N_17239);
or U18901 (N_18901,N_16453,N_15327);
and U18902 (N_18902,N_14064,N_14301);
xnor U18903 (N_18903,N_15313,N_14726);
and U18904 (N_18904,N_15393,N_14278);
or U18905 (N_18905,N_18617,N_13156);
xor U18906 (N_18906,N_15961,N_18107);
xnor U18907 (N_18907,N_14613,N_17365);
nand U18908 (N_18908,N_13510,N_12907);
or U18909 (N_18909,N_18611,N_13975);
nor U18910 (N_18910,N_14611,N_14361);
or U18911 (N_18911,N_12626,N_17826);
or U18912 (N_18912,N_13646,N_15992);
nor U18913 (N_18913,N_16850,N_15679);
xnor U18914 (N_18914,N_13457,N_15369);
xnor U18915 (N_18915,N_13447,N_17303);
xor U18916 (N_18916,N_17547,N_16776);
nor U18917 (N_18917,N_17311,N_15000);
nand U18918 (N_18918,N_14028,N_15385);
and U18919 (N_18919,N_14559,N_18275);
nand U18920 (N_18920,N_17546,N_17366);
nand U18921 (N_18921,N_12645,N_15518);
and U18922 (N_18922,N_16962,N_16569);
or U18923 (N_18923,N_12547,N_18599);
and U18924 (N_18924,N_12920,N_16998);
nor U18925 (N_18925,N_18090,N_14554);
nor U18926 (N_18926,N_16273,N_13045);
nand U18927 (N_18927,N_17307,N_16517);
or U18928 (N_18928,N_13790,N_16055);
nor U18929 (N_18929,N_15788,N_14162);
nor U18930 (N_18930,N_13032,N_18467);
or U18931 (N_18931,N_15035,N_14073);
nor U18932 (N_18932,N_16500,N_17506);
nor U18933 (N_18933,N_13972,N_17453);
nor U18934 (N_18934,N_14988,N_16547);
nor U18935 (N_18935,N_14088,N_17660);
and U18936 (N_18936,N_13664,N_13267);
or U18937 (N_18937,N_13444,N_14086);
xor U18938 (N_18938,N_13486,N_15454);
nand U18939 (N_18939,N_16052,N_16508);
and U18940 (N_18940,N_14699,N_14286);
nor U18941 (N_18941,N_15277,N_16039);
nand U18942 (N_18942,N_14400,N_16729);
or U18943 (N_18943,N_18651,N_13603);
xnor U18944 (N_18944,N_15195,N_16184);
or U18945 (N_18945,N_14594,N_16908);
xnor U18946 (N_18946,N_13320,N_18685);
or U18947 (N_18947,N_18316,N_12928);
and U18948 (N_18948,N_14231,N_17081);
nand U18949 (N_18949,N_13049,N_18127);
nand U18950 (N_18950,N_14713,N_13903);
nand U18951 (N_18951,N_15226,N_15224);
nor U18952 (N_18952,N_15392,N_16014);
and U18953 (N_18953,N_13058,N_15878);
xor U18954 (N_18954,N_18402,N_13794);
or U18955 (N_18955,N_15124,N_14982);
and U18956 (N_18956,N_12736,N_18655);
nor U18957 (N_18957,N_13448,N_16946);
nor U18958 (N_18958,N_15605,N_12978);
xnor U18959 (N_18959,N_13658,N_14159);
nor U18960 (N_18960,N_17789,N_17493);
and U18961 (N_18961,N_13605,N_17484);
and U18962 (N_18962,N_14129,N_17606);
and U18963 (N_18963,N_14695,N_16128);
or U18964 (N_18964,N_18388,N_17051);
nand U18965 (N_18965,N_15519,N_13173);
nand U18966 (N_18966,N_16731,N_12583);
or U18967 (N_18967,N_13879,N_16821);
or U18968 (N_18968,N_16930,N_14310);
nor U18969 (N_18969,N_18050,N_15090);
nor U18970 (N_18970,N_16375,N_16073);
nor U18971 (N_18971,N_13142,N_15796);
and U18972 (N_18972,N_15044,N_18022);
nand U18973 (N_18973,N_17994,N_15434);
nor U18974 (N_18974,N_14058,N_12851);
xor U18975 (N_18975,N_17703,N_16141);
xor U18976 (N_18976,N_17697,N_15775);
or U18977 (N_18977,N_14810,N_17165);
and U18978 (N_18978,N_18193,N_13995);
nor U18979 (N_18979,N_13169,N_17009);
nand U18980 (N_18980,N_13039,N_15940);
or U18981 (N_18981,N_13266,N_12610);
xor U18982 (N_18982,N_15113,N_18576);
and U18983 (N_18983,N_17610,N_15744);
xor U18984 (N_18984,N_14326,N_18042);
nor U18985 (N_18985,N_13850,N_12556);
nor U18986 (N_18986,N_15105,N_14715);
and U18987 (N_18987,N_17709,N_16921);
nor U18988 (N_18988,N_14808,N_17730);
xor U18989 (N_18989,N_13549,N_18295);
xor U18990 (N_18990,N_16648,N_15246);
nand U18991 (N_18991,N_16314,N_14953);
nand U18992 (N_18992,N_12676,N_18059);
or U18993 (N_18993,N_16805,N_17375);
xor U18994 (N_18994,N_16788,N_16863);
nand U18995 (N_18995,N_15506,N_14732);
nor U18996 (N_18996,N_17500,N_18548);
and U18997 (N_18997,N_13709,N_13084);
and U18998 (N_18998,N_13229,N_17732);
nor U18999 (N_18999,N_13683,N_17976);
or U19000 (N_19000,N_16640,N_13748);
nand U19001 (N_19001,N_17794,N_16552);
or U19002 (N_19002,N_14377,N_15347);
and U19003 (N_19003,N_13633,N_16029);
and U19004 (N_19004,N_16684,N_16306);
xor U19005 (N_19005,N_13984,N_15710);
or U19006 (N_19006,N_16732,N_18176);
nor U19007 (N_19007,N_15926,N_12872);
nand U19008 (N_19008,N_13262,N_18328);
nand U19009 (N_19009,N_18741,N_14452);
and U19010 (N_19010,N_18277,N_18594);
xor U19011 (N_19011,N_16905,N_14209);
nor U19012 (N_19012,N_18452,N_16406);
nor U19013 (N_19013,N_15736,N_17818);
xnor U19014 (N_19014,N_17588,N_18478);
nor U19015 (N_19015,N_18115,N_12582);
xnor U19016 (N_19016,N_17459,N_17445);
xnor U19017 (N_19017,N_16614,N_14974);
and U19018 (N_19018,N_18013,N_14185);
xor U19019 (N_19019,N_17919,N_14106);
nand U19020 (N_19020,N_14583,N_15364);
xnor U19021 (N_19021,N_13224,N_17056);
or U19022 (N_19022,N_18263,N_14772);
nand U19023 (N_19023,N_14677,N_16549);
or U19024 (N_19024,N_12546,N_18266);
nand U19025 (N_19025,N_16363,N_17584);
nand U19026 (N_19026,N_12634,N_13590);
nand U19027 (N_19027,N_14218,N_17632);
nand U19028 (N_19028,N_12588,N_12566);
or U19029 (N_19029,N_15989,N_16299);
xnor U19030 (N_19030,N_13104,N_15322);
nor U19031 (N_19031,N_12799,N_17599);
nand U19032 (N_19032,N_16818,N_17939);
or U19033 (N_19033,N_14413,N_17333);
nand U19034 (N_19034,N_14020,N_15995);
nor U19035 (N_19035,N_17001,N_12611);
or U19036 (N_19036,N_14662,N_15648);
and U19037 (N_19037,N_13698,N_15990);
nand U19038 (N_19038,N_16992,N_13671);
and U19039 (N_19039,N_15138,N_13556);
and U19040 (N_19040,N_17684,N_14633);
nand U19041 (N_19041,N_15714,N_17628);
nor U19042 (N_19042,N_13435,N_12908);
and U19043 (N_19043,N_16478,N_17969);
or U19044 (N_19044,N_17889,N_18498);
xor U19045 (N_19045,N_16539,N_17049);
nor U19046 (N_19046,N_15779,N_15001);
nand U19047 (N_19047,N_17966,N_18141);
nand U19048 (N_19048,N_14896,N_12889);
nand U19049 (N_19049,N_16572,N_17601);
and U19050 (N_19050,N_15869,N_14091);
xor U19051 (N_19051,N_16896,N_12927);
nor U19052 (N_19052,N_13766,N_14477);
and U19053 (N_19053,N_16310,N_16078);
nand U19054 (N_19054,N_16289,N_15484);
and U19055 (N_19055,N_17289,N_17345);
or U19056 (N_19056,N_16487,N_18453);
and U19057 (N_19057,N_17997,N_18162);
nand U19058 (N_19058,N_16711,N_12892);
and U19059 (N_19059,N_16615,N_14227);
nor U19060 (N_19060,N_14587,N_17381);
nor U19061 (N_19061,N_16165,N_16189);
nor U19062 (N_19062,N_17204,N_15447);
or U19063 (N_19063,N_12817,N_15855);
xor U19064 (N_19064,N_12827,N_17869);
nor U19065 (N_19065,N_17291,N_16510);
nor U19066 (N_19066,N_17943,N_16503);
xnor U19067 (N_19067,N_12980,N_17321);
nand U19068 (N_19068,N_13547,N_15650);
and U19069 (N_19069,N_17952,N_13472);
nand U19070 (N_19070,N_13280,N_12791);
nor U19071 (N_19071,N_18739,N_13754);
or U19072 (N_19072,N_15167,N_16149);
nor U19073 (N_19073,N_15244,N_16111);
and U19074 (N_19074,N_14744,N_16103);
or U19075 (N_19075,N_13710,N_15960);
or U19076 (N_19076,N_17431,N_12848);
nor U19077 (N_19077,N_14443,N_13715);
and U19078 (N_19078,N_17698,N_15697);
nand U19079 (N_19079,N_12722,N_14548);
nand U19080 (N_19080,N_13842,N_12670);
nor U19081 (N_19081,N_15398,N_15932);
xor U19082 (N_19082,N_17523,N_15482);
nor U19083 (N_19083,N_16974,N_15287);
nor U19084 (N_19084,N_16768,N_18561);
xor U19085 (N_19085,N_12876,N_17669);
nor U19086 (N_19086,N_17949,N_13133);
xor U19087 (N_19087,N_14290,N_16178);
xor U19088 (N_19088,N_17141,N_16744);
and U19089 (N_19089,N_14618,N_17674);
nor U19090 (N_19090,N_17614,N_16831);
nand U19091 (N_19091,N_14098,N_15358);
nand U19092 (N_19092,N_15691,N_12865);
or U19093 (N_19093,N_17274,N_17125);
and U19094 (N_19094,N_15896,N_15439);
nand U19095 (N_19095,N_14832,N_13005);
nor U19096 (N_19096,N_17787,N_16439);
or U19097 (N_19097,N_15264,N_17560);
or U19098 (N_19098,N_13347,N_16769);
and U19099 (N_19099,N_17786,N_14918);
xnor U19100 (N_19100,N_18497,N_14516);
nand U19101 (N_19101,N_16385,N_16745);
or U19102 (N_19102,N_14370,N_15923);
and U19103 (N_19103,N_15712,N_17180);
nor U19104 (N_19104,N_12959,N_15554);
nand U19105 (N_19105,N_16535,N_16056);
nor U19106 (N_19106,N_13137,N_13211);
and U19107 (N_19107,N_15967,N_13947);
nor U19108 (N_19108,N_13225,N_16362);
nor U19109 (N_19109,N_15805,N_16241);
or U19110 (N_19110,N_15108,N_14132);
and U19111 (N_19111,N_14048,N_16163);
nor U19112 (N_19112,N_18367,N_14187);
nor U19113 (N_19113,N_14962,N_16442);
nor U19114 (N_19114,N_15726,N_15953);
nor U19115 (N_19115,N_18355,N_17676);
and U19116 (N_19116,N_17076,N_16457);
and U19117 (N_19117,N_13430,N_14099);
xnor U19118 (N_19118,N_15437,N_18416);
nor U19119 (N_19119,N_13082,N_16042);
or U19120 (N_19120,N_13086,N_18188);
and U19121 (N_19121,N_13382,N_16413);
and U19122 (N_19122,N_18058,N_15361);
nor U19123 (N_19123,N_14202,N_12625);
or U19124 (N_19124,N_16735,N_17670);
and U19125 (N_19125,N_17817,N_17718);
and U19126 (N_19126,N_18656,N_13064);
nand U19127 (N_19127,N_14283,N_18103);
or U19128 (N_19128,N_16809,N_13034);
or U19129 (N_19129,N_16807,N_17624);
nand U19130 (N_19130,N_15107,N_15689);
nand U19131 (N_19131,N_17578,N_13431);
nor U19132 (N_19132,N_14070,N_15041);
nand U19133 (N_19133,N_12926,N_18647);
or U19134 (N_19134,N_12945,N_16026);
nor U19135 (N_19135,N_13544,N_17065);
nor U19136 (N_19136,N_16701,N_12691);
nand U19137 (N_19137,N_14480,N_12895);
xor U19138 (N_19138,N_13852,N_13380);
nand U19139 (N_19139,N_15324,N_17002);
nor U19140 (N_19140,N_15221,N_17197);
xor U19141 (N_19141,N_14894,N_12751);
xor U19142 (N_19142,N_15680,N_13451);
xnor U19143 (N_19143,N_13836,N_16512);
and U19144 (N_19144,N_16815,N_15418);
nand U19145 (N_19145,N_16245,N_16579);
or U19146 (N_19146,N_12574,N_17540);
nand U19147 (N_19147,N_16839,N_15150);
or U19148 (N_19148,N_16166,N_14169);
and U19149 (N_19149,N_12699,N_13061);
or U19150 (N_19150,N_13127,N_14444);
xnor U19151 (N_19151,N_17330,N_14501);
or U19152 (N_19152,N_13685,N_14276);
nand U19153 (N_19153,N_14509,N_15891);
or U19154 (N_19154,N_16079,N_14619);
nand U19155 (N_19155,N_17388,N_15292);
and U19156 (N_19156,N_16064,N_14579);
nand U19157 (N_19157,N_17151,N_15898);
and U19158 (N_19158,N_18354,N_15631);
or U19159 (N_19159,N_17912,N_12897);
nand U19160 (N_19160,N_13198,N_13914);
or U19161 (N_19161,N_13323,N_17349);
nor U19162 (N_19162,N_18337,N_17206);
and U19163 (N_19163,N_16789,N_15471);
xnor U19164 (N_19164,N_14024,N_17182);
and U19165 (N_19165,N_14857,N_16311);
and U19166 (N_19166,N_15033,N_17917);
nor U19167 (N_19167,N_18029,N_17605);
xor U19168 (N_19168,N_18426,N_13812);
or U19169 (N_19169,N_14534,N_14538);
nor U19170 (N_19170,N_14497,N_14814);
nor U19171 (N_19171,N_15661,N_17383);
nand U19172 (N_19172,N_16309,N_16326);
or U19173 (N_19173,N_17285,N_12792);
xor U19174 (N_19174,N_18150,N_13492);
and U19175 (N_19175,N_17749,N_13179);
nand U19176 (N_19176,N_18339,N_13487);
nor U19177 (N_19177,N_15157,N_13376);
nor U19178 (N_19178,N_16050,N_18442);
nand U19179 (N_19179,N_14313,N_14386);
or U19180 (N_19180,N_13562,N_14936);
xor U19181 (N_19181,N_18242,N_13138);
or U19182 (N_19182,N_14920,N_12538);
or U19183 (N_19183,N_17758,N_15789);
or U19184 (N_19184,N_16197,N_14463);
nor U19185 (N_19185,N_12916,N_13884);
nand U19186 (N_19186,N_16990,N_13707);
nor U19187 (N_19187,N_18466,N_17327);
nand U19188 (N_19188,N_13939,N_14348);
xor U19189 (N_19189,N_14019,N_17017);
xnor U19190 (N_19190,N_12562,N_13333);
nand U19191 (N_19191,N_14803,N_16301);
nand U19192 (N_19192,N_14359,N_14552);
nand U19193 (N_19193,N_14036,N_17347);
or U19194 (N_19194,N_16335,N_13019);
or U19195 (N_19195,N_14349,N_14621);
nand U19196 (N_19196,N_13774,N_16242);
nor U19197 (N_19197,N_16760,N_13305);
nand U19198 (N_19198,N_16881,N_13967);
or U19199 (N_19199,N_16519,N_16794);
or U19200 (N_19200,N_14758,N_14863);
and U19201 (N_19201,N_18051,N_17675);
xor U19202 (N_19202,N_13147,N_15480);
xnor U19203 (N_19203,N_16754,N_12784);
and U19204 (N_19204,N_16867,N_16995);
or U19205 (N_19205,N_16853,N_12619);
nand U19206 (N_19206,N_15873,N_17183);
xnor U19207 (N_19207,N_13324,N_15184);
or U19208 (N_19208,N_16620,N_16793);
xor U19209 (N_19209,N_15809,N_12795);
xnor U19210 (N_19210,N_14610,N_17185);
xnor U19211 (N_19211,N_16228,N_16922);
xnor U19212 (N_19212,N_15207,N_16396);
xnor U19213 (N_19213,N_17565,N_18201);
nor U19214 (N_19214,N_17087,N_17243);
xnor U19215 (N_19215,N_16953,N_16376);
or U19216 (N_19216,N_14229,N_12942);
and U19217 (N_19217,N_13394,N_13857);
nand U19218 (N_19218,N_15653,N_17972);
and U19219 (N_19219,N_14395,N_13017);
nor U19220 (N_19220,N_12777,N_15582);
and U19221 (N_19221,N_18182,N_13721);
xor U19222 (N_19222,N_12918,N_15758);
xnor U19223 (N_19223,N_14499,N_18132);
and U19224 (N_19224,N_16890,N_14986);
nand U19225 (N_19225,N_12675,N_16332);
nand U19226 (N_19226,N_18134,N_14161);
or U19227 (N_19227,N_14753,N_13135);
or U19228 (N_19228,N_17816,N_15981);
xor U19229 (N_19229,N_15993,N_12738);
and U19230 (N_19230,N_15045,N_13570);
xnor U19231 (N_19231,N_15096,N_15078);
nand U19232 (N_19232,N_17831,N_15667);
xor U19233 (N_19233,N_18098,N_12651);
or U19234 (N_19234,N_15334,N_18494);
and U19235 (N_19235,N_13007,N_18488);
and U19236 (N_19236,N_13300,N_13065);
and U19237 (N_19237,N_13063,N_16557);
nor U19238 (N_19238,N_14755,N_13691);
nand U19239 (N_19239,N_15552,N_18158);
nor U19240 (N_19240,N_13531,N_13110);
nor U19241 (N_19241,N_18582,N_14394);
and U19242 (N_19242,N_18186,N_16341);
nand U19243 (N_19243,N_14717,N_14127);
and U19244 (N_19244,N_13704,N_14267);
xnor U19245 (N_19245,N_13613,N_14249);
nand U19246 (N_19246,N_17485,N_16824);
or U19247 (N_19247,N_16619,N_12869);
nor U19248 (N_19248,N_12708,N_18744);
or U19249 (N_19249,N_14047,N_14493);
or U19250 (N_19250,N_18626,N_17881);
xor U19251 (N_19251,N_13588,N_15912);
or U19252 (N_19252,N_17112,N_15611);
xor U19253 (N_19253,N_14887,N_17150);
or U19254 (N_19254,N_13003,N_13755);
and U19255 (N_19255,N_13795,N_16887);
or U19256 (N_19256,N_18219,N_12854);
xor U19257 (N_19257,N_13591,N_17122);
xor U19258 (N_19258,N_14236,N_15381);
nor U19259 (N_19259,N_14770,N_12861);
xor U19260 (N_19260,N_13379,N_17423);
or U19261 (N_19261,N_15701,N_15880);
and U19262 (N_19262,N_16499,N_18521);
xnor U19263 (N_19263,N_14737,N_15297);
nor U19264 (N_19264,N_15352,N_18379);
and U19265 (N_19265,N_13330,N_14551);
nor U19266 (N_19266,N_17907,N_13724);
nor U19267 (N_19267,N_12637,N_14550);
and U19268 (N_19268,N_14830,N_17731);
or U19269 (N_19269,N_13665,N_14145);
and U19270 (N_19270,N_13901,N_18319);
nand U19271 (N_19271,N_17354,N_14951);
or U19272 (N_19272,N_15382,N_14971);
xnor U19273 (N_19273,N_18077,N_13674);
and U19274 (N_19274,N_18615,N_16468);
nor U19275 (N_19275,N_14629,N_13490);
and U19276 (N_19276,N_13627,N_14696);
or U19277 (N_19277,N_15618,N_14911);
xor U19278 (N_19278,N_17154,N_14492);
and U19279 (N_19279,N_17951,N_17279);
or U19280 (N_19280,N_12787,N_12821);
nand U19281 (N_19281,N_13511,N_13364);
nand U19282 (N_19282,N_18455,N_16327);
xnor U19283 (N_19283,N_15010,N_12614);
nand U19284 (N_19284,N_15093,N_18740);
or U19285 (N_19285,N_14163,N_17040);
xnor U19286 (N_19286,N_17086,N_16004);
and U19287 (N_19287,N_14353,N_13572);
xnor U19288 (N_19288,N_14496,N_12852);
and U19289 (N_19289,N_18312,N_16520);
nor U19290 (N_19290,N_15116,N_17741);
xnor U19291 (N_19291,N_14933,N_14396);
or U19292 (N_19292,N_12800,N_18100);
nor U19293 (N_19293,N_16806,N_18113);
nand U19294 (N_19294,N_17957,N_17248);
xnor U19295 (N_19295,N_14448,N_13833);
xnor U19296 (N_19296,N_15363,N_13546);
or U19297 (N_19297,N_15935,N_18369);
xnor U19298 (N_19298,N_17740,N_16982);
and U19299 (N_19299,N_16034,N_18119);
or U19300 (N_19300,N_16531,N_15592);
and U19301 (N_19301,N_16688,N_17558);
nor U19302 (N_19302,N_12874,N_14844);
nor U19303 (N_19303,N_13679,N_13092);
xor U19304 (N_19304,N_12868,N_16848);
or U19305 (N_19305,N_14719,N_13093);
xor U19306 (N_19306,N_13782,N_13501);
and U19307 (N_19307,N_14060,N_18749);
nand U19308 (N_19308,N_16011,N_14531);
xor U19309 (N_19309,N_15114,N_12616);
nand U19310 (N_19310,N_12903,N_15664);
and U19311 (N_19311,N_16915,N_14688);
xor U19312 (N_19312,N_15766,N_13611);
nand U19313 (N_19313,N_17815,N_12687);
or U19314 (N_19314,N_16338,N_14110);
or U19315 (N_19315,N_18424,N_17380);
nand U19316 (N_19316,N_16903,N_14646);
nor U19317 (N_19317,N_18589,N_14200);
xor U19318 (N_19318,N_17178,N_16507);
or U19319 (N_19319,N_17678,N_15417);
xnor U19320 (N_19320,N_16970,N_16624);
nor U19321 (N_19321,N_15784,N_12686);
nand U19322 (N_19322,N_15100,N_13029);
nor U19323 (N_19323,N_13423,N_14730);
xnor U19324 (N_19324,N_13642,N_14597);
xnor U19325 (N_19325,N_17896,N_12909);
and U19326 (N_19326,N_13038,N_17677);
nor U19327 (N_19327,N_13771,N_14768);
xnor U19328 (N_19328,N_15902,N_13283);
nand U19329 (N_19329,N_13113,N_17314);
or U19330 (N_19330,N_15072,N_15922);
xnor U19331 (N_19331,N_18730,N_15020);
nor U19332 (N_19332,N_17210,N_16246);
and U19333 (N_19333,N_16389,N_14756);
nand U19334 (N_19334,N_15153,N_15288);
nor U19335 (N_19335,N_15602,N_15021);
xnor U19336 (N_19336,N_13797,N_13445);
nor U19337 (N_19337,N_18673,N_17862);
or U19338 (N_19338,N_15979,N_12771);
or U19339 (N_19339,N_17320,N_18217);
nor U19340 (N_19340,N_15780,N_14963);
or U19341 (N_19341,N_15310,N_14886);
or U19342 (N_19342,N_16109,N_15885);
xor U19343 (N_19343,N_15306,N_14412);
and U19344 (N_19344,N_17412,N_16069);
xor U19345 (N_19345,N_14030,N_13609);
nand U19346 (N_19346,N_13233,N_17983);
or U19347 (N_19347,N_17735,N_13731);
and U19348 (N_19348,N_15972,N_13247);
xor U19349 (N_19349,N_17572,N_13678);
nand U19350 (N_19350,N_14735,N_17164);
and U19351 (N_19351,N_16756,N_12890);
or U19352 (N_19352,N_14957,N_17724);
and U19353 (N_19353,N_14238,N_13270);
xnor U19354 (N_19354,N_12822,N_18049);
or U19355 (N_19355,N_15182,N_16402);
xor U19356 (N_19356,N_18094,N_13365);
xnor U19357 (N_19357,N_14822,N_14801);
xor U19358 (N_19358,N_15344,N_15414);
or U19359 (N_19359,N_14627,N_17808);
nor U19360 (N_19360,N_14711,N_13328);
nor U19361 (N_19361,N_14346,N_16748);
xnor U19362 (N_19362,N_13303,N_18340);
nand U19363 (N_19363,N_12818,N_13338);
nand U19364 (N_19364,N_14005,N_14222);
and U19365 (N_19365,N_18653,N_14027);
nand U19366 (N_19366,N_13700,N_15228);
nand U19367 (N_19367,N_15820,N_12721);
or U19368 (N_19368,N_15455,N_13604);
nor U19369 (N_19369,N_15867,N_14158);
xnor U19370 (N_19370,N_15508,N_14905);
or U19371 (N_19371,N_14450,N_12630);
and U19372 (N_19372,N_14557,N_16955);
nand U19373 (N_19373,N_13341,N_15106);
and U19374 (N_19374,N_14519,N_13703);
nand U19375 (N_19375,N_15175,N_14258);
or U19376 (N_19376,N_18415,N_18409);
or U19377 (N_19377,N_13589,N_15920);
nor U19378 (N_19378,N_14472,N_13015);
and U19379 (N_19379,N_13566,N_13826);
or U19380 (N_19380,N_17444,N_15423);
and U19381 (N_19381,N_17251,N_13391);
or U19382 (N_19382,N_15890,N_15346);
xnor U19383 (N_19383,N_16901,N_16354);
xnor U19384 (N_19384,N_18118,N_16437);
nor U19385 (N_19385,N_17096,N_18131);
and U19386 (N_19386,N_13097,N_14384);
or U19387 (N_19387,N_14095,N_15829);
nand U19388 (N_19388,N_15842,N_14842);
xor U19389 (N_19389,N_13600,N_15256);
nor U19390 (N_19390,N_15786,N_13111);
or U19391 (N_19391,N_17595,N_18624);
nor U19392 (N_19392,N_15349,N_16501);
or U19393 (N_19393,N_17664,N_18564);
nor U19394 (N_19394,N_12508,N_16830);
xnor U19395 (N_19395,N_17766,N_15925);
xnor U19396 (N_19396,N_16912,N_12503);
or U19397 (N_19397,N_12977,N_13223);
xor U19398 (N_19398,N_15539,N_15091);
nand U19399 (N_19399,N_15411,N_15555);
or U19400 (N_19400,N_16699,N_17401);
xor U19401 (N_19401,N_13175,N_17544);
and U19402 (N_19402,N_18715,N_14490);
or U19403 (N_19403,N_15765,N_15768);
nor U19404 (N_19404,N_17213,N_18074);
and U19405 (N_19405,N_12682,N_12783);
nor U19406 (N_19406,N_16835,N_13374);
or U19407 (N_19407,N_16734,N_16838);
nand U19408 (N_19408,N_17155,N_12545);
xor U19409 (N_19409,N_12911,N_12688);
nor U19410 (N_19410,N_17438,N_17870);
and U19411 (N_19411,N_15973,N_12602);
and U19412 (N_19412,N_12893,N_14362);
and U19413 (N_19413,N_16906,N_15939);
nand U19414 (N_19414,N_17247,N_15949);
or U19415 (N_19415,N_13349,N_16691);
or U19416 (N_19416,N_16804,N_16260);
nand U19417 (N_19417,N_13926,N_18476);
and U19418 (N_19418,N_15267,N_17663);
and U19419 (N_19419,N_14345,N_17673);
or U19420 (N_19420,N_18657,N_13461);
or U19421 (N_19421,N_14331,N_17745);
or U19422 (N_19422,N_16891,N_14025);
xnor U19423 (N_19423,N_17280,N_13426);
nor U19424 (N_19424,N_15492,N_13377);
or U19425 (N_19425,N_18019,N_14578);
nor U19426 (N_19426,N_14328,N_16261);
and U19427 (N_19427,N_12725,N_16177);
or U19428 (N_19428,N_17836,N_17507);
and U19429 (N_19429,N_14545,N_13834);
xor U19430 (N_19430,N_17571,N_14707);
xnor U19431 (N_19431,N_13208,N_15082);
nand U19432 (N_19432,N_15586,N_18037);
or U19433 (N_19433,N_14817,N_17564);
and U19434 (N_19434,N_13414,N_12677);
nor U19435 (N_19435,N_12674,N_13524);
and U19436 (N_19436,N_13718,N_15137);
xor U19437 (N_19437,N_17704,N_13610);
or U19438 (N_19438,N_14773,N_14174);
xnor U19439 (N_19439,N_14100,N_15389);
nor U19440 (N_19440,N_15832,N_15284);
nor U19441 (N_19441,N_15763,N_14877);
nand U19442 (N_19442,N_16522,N_14125);
and U19443 (N_19443,N_17511,N_16131);
or U19444 (N_19444,N_17405,N_15985);
nor U19445 (N_19445,N_12951,N_16490);
nor U19446 (N_19446,N_17570,N_16554);
nor U19447 (N_19447,N_18030,N_16840);
and U19448 (N_19448,N_18699,N_17465);
nor U19449 (N_19449,N_14398,N_14507);
and U19450 (N_19450,N_18025,N_13657);
nor U19451 (N_19451,N_14874,N_17946);
nand U19452 (N_19452,N_18039,N_13484);
and U19453 (N_19453,N_18283,N_14080);
nor U19454 (N_19454,N_16404,N_16108);
or U19455 (N_19455,N_17639,N_16359);
xor U19456 (N_19456,N_16337,N_18258);
xor U19457 (N_19457,N_14504,N_16191);
or U19458 (N_19458,N_15696,N_13593);
or U19459 (N_19459,N_16144,N_13845);
nor U19460 (N_19460,N_17487,N_17083);
or U19461 (N_19461,N_17348,N_14087);
xor U19462 (N_19462,N_17941,N_14149);
xor U19463 (N_19463,N_18221,N_18400);
nor U19464 (N_19464,N_16796,N_13936);
or U19465 (N_19465,N_13738,N_14113);
or U19466 (N_19466,N_16929,N_12530);
xnor U19467 (N_19467,N_14152,N_17263);
xnor U19468 (N_19468,N_18362,N_17466);
nand U19469 (N_19469,N_13352,N_14102);
or U19470 (N_19470,N_16018,N_14414);
and U19471 (N_19471,N_18265,N_15741);
and U19472 (N_19472,N_16698,N_15378);
nor U19473 (N_19473,N_15916,N_18648);
or U19474 (N_19474,N_16045,N_18506);
nor U19475 (N_19475,N_13390,N_17121);
or U19476 (N_19476,N_18578,N_18583);
xnor U19477 (N_19477,N_18505,N_12695);
and U19478 (N_19478,N_15693,N_16773);
nor U19479 (N_19479,N_13800,N_17374);
nand U19480 (N_19480,N_16973,N_14883);
nand U19481 (N_19481,N_18390,N_14804);
nand U19482 (N_19482,N_14895,N_17501);
and U19483 (N_19483,N_13785,N_14915);
or U19484 (N_19484,N_12701,N_13053);
or U19485 (N_19485,N_16139,N_15956);
or U19486 (N_19486,N_14568,N_16360);
and U19487 (N_19487,N_14601,N_18540);
and U19488 (N_19488,N_16904,N_15088);
nor U19489 (N_19489,N_12859,N_14002);
nor U19490 (N_19490,N_15881,N_15849);
and U19491 (N_19491,N_16114,N_16635);
nand U19492 (N_19492,N_17364,N_13961);
xnor U19493 (N_19493,N_17179,N_18634);
or U19494 (N_19494,N_18464,N_16044);
nor U19495 (N_19495,N_18250,N_16586);
and U19496 (N_19496,N_16157,N_17010);
nand U19497 (N_19497,N_13059,N_16160);
and U19498 (N_19498,N_18060,N_17657);
nand U19499 (N_19499,N_16036,N_15887);
and U19500 (N_19500,N_13197,N_12589);
nand U19501 (N_19501,N_13485,N_15007);
xnor U19502 (N_19502,N_17813,N_14280);
or U19503 (N_19503,N_13499,N_15075);
xor U19504 (N_19504,N_17620,N_15473);
or U19505 (N_19505,N_14004,N_13909);
nor U19506 (N_19506,N_18069,N_15499);
nand U19507 (N_19507,N_18609,N_12933);
or U19508 (N_19508,N_16743,N_14925);
and U19509 (N_19509,N_17561,N_16696);
or U19510 (N_19510,N_13596,N_18305);
nor U19511 (N_19511,N_16466,N_17385);
and U19512 (N_19512,N_15646,N_17888);
or U19513 (N_19513,N_14771,N_14284);
or U19514 (N_19514,N_18620,N_17341);
or U19515 (N_19515,N_16345,N_16592);
or U19516 (N_19516,N_15144,N_16296);
and U19517 (N_19517,N_17654,N_16669);
and U19518 (N_19518,N_13628,N_13859);
xor U19519 (N_19519,N_16917,N_14969);
nor U19520 (N_19520,N_13929,N_14316);
or U19521 (N_19521,N_14419,N_17221);
or U19522 (N_19522,N_15146,N_12655);
or U19523 (N_19523,N_18318,N_15535);
nor U19524 (N_19524,N_17761,N_18070);
nor U19525 (N_19525,N_18413,N_15735);
xnor U19526 (N_19526,N_17433,N_18041);
and U19527 (N_19527,N_18274,N_18352);
or U19528 (N_19528,N_16482,N_18111);
or U19529 (N_19529,N_13157,N_13459);
nor U19530 (N_19530,N_14805,N_15038);
nand U19531 (N_19531,N_17904,N_13035);
nand U19532 (N_19532,N_16766,N_15258);
or U19533 (N_19533,N_17782,N_15730);
nor U19534 (N_19534,N_13207,N_15904);
nand U19535 (N_19535,N_13454,N_17089);
nor U19536 (N_19536,N_16952,N_14524);
and U19537 (N_19537,N_12653,N_15071);
nor U19538 (N_19538,N_15469,N_12502);
nand U19539 (N_19539,N_15792,N_13442);
or U19540 (N_19540,N_12785,N_14074);
nor U19541 (N_19541,N_17075,N_13740);
nand U19542 (N_19542,N_17326,N_15843);
and U19543 (N_19543,N_17618,N_14263);
nor U19544 (N_19544,N_12608,N_18543);
xor U19545 (N_19545,N_17215,N_16676);
or U19546 (N_19546,N_18737,N_12702);
and U19547 (N_19547,N_16174,N_16623);
nor U19548 (N_19548,N_16136,N_15963);
xnor U19549 (N_19549,N_15651,N_17579);
xnor U19550 (N_19550,N_17621,N_15225);
nor U19551 (N_19551,N_16416,N_17146);
and U19552 (N_19552,N_13946,N_13235);
nand U19553 (N_19553,N_15280,N_17419);
xnor U19554 (N_19554,N_13067,N_14606);
or U19555 (N_19555,N_15276,N_14826);
or U19556 (N_19556,N_16607,N_14144);
and U19557 (N_19557,N_14094,N_17389);
and U19558 (N_19558,N_18562,N_16209);
or U19559 (N_19559,N_15913,N_15991);
xnor U19560 (N_19560,N_17886,N_18604);
or U19561 (N_19561,N_12689,N_12841);
xor U19562 (N_19562,N_15756,N_12842);
or U19563 (N_19563,N_13584,N_17880);
xnor U19564 (N_19564,N_16013,N_17970);
nor U19565 (N_19565,N_16902,N_13318);
nor U19566 (N_19566,N_18336,N_14862);
or U19567 (N_19567,N_15797,N_13060);
nor U19568 (N_19568,N_17013,N_15301);
nor U19569 (N_19569,N_17426,N_15527);
nand U19570 (N_19570,N_18710,N_15104);
or U19571 (N_19571,N_14470,N_13890);
nand U19572 (N_19572,N_16565,N_13987);
and U19573 (N_19573,N_14675,N_17954);
nor U19574 (N_19574,N_18565,N_17909);
and U19575 (N_19575,N_13513,N_18495);
and U19576 (N_19576,N_17335,N_13615);
nor U19577 (N_19577,N_18429,N_16455);
nor U19578 (N_19578,N_13277,N_16515);
nor U19579 (N_19579,N_14273,N_12992);
or U19580 (N_19580,N_16300,N_13777);
xnor U19581 (N_19581,N_16637,N_14809);
nand U19582 (N_19582,N_17491,N_14706);
nand U19583 (N_19583,N_17450,N_14403);
and U19584 (N_19584,N_18230,N_13730);
and U19585 (N_19585,N_15254,N_16074);
nor U19586 (N_19586,N_16256,N_17368);
and U19587 (N_19587,N_16243,N_17701);
nand U19588 (N_19588,N_15173,N_15601);
xor U19589 (N_19589,N_16714,N_17722);
nor U19590 (N_19590,N_18658,N_14843);
xor U19591 (N_19591,N_12705,N_14254);
or U19592 (N_19592,N_14793,N_18366);
and U19593 (N_19593,N_18550,N_16293);
nor U19594 (N_19594,N_18174,N_15537);
and U19595 (N_19595,N_17014,N_15544);
xnor U19596 (N_19596,N_16790,N_16130);
nor U19597 (N_19597,N_14525,N_17792);
or U19598 (N_19598,N_13470,N_13954);
nand U19599 (N_19599,N_14738,N_13693);
and U19600 (N_19600,N_13594,N_13136);
nand U19601 (N_19601,N_12744,N_12860);
nand U19602 (N_19602,N_12564,N_17845);
xnor U19603 (N_19603,N_13162,N_14664);
xnor U19604 (N_19604,N_16403,N_15641);
nand U19605 (N_19605,N_18727,N_14766);
or U19606 (N_19606,N_16528,N_17464);
or U19607 (N_19607,N_15800,N_16934);
xor U19608 (N_19608,N_15966,N_17379);
or U19609 (N_19609,N_12570,N_16324);
nor U19610 (N_19610,N_12750,N_18704);
or U19611 (N_19611,N_16994,N_17623);
nor U19612 (N_19612,N_16193,N_15318);
xnor U19613 (N_19613,N_13817,N_14434);
and U19614 (N_19614,N_15465,N_14837);
nor U19615 (N_19615,N_18717,N_17295);
nor U19616 (N_19616,N_17842,N_14834);
and U19617 (N_19617,N_18140,N_17101);
xor U19618 (N_19618,N_16646,N_17169);
nand U19619 (N_19619,N_12618,N_14368);
xor U19620 (N_19620,N_12986,N_16588);
nor U19621 (N_19621,N_16318,N_13355);
nand U19622 (N_19622,N_13234,N_13945);
xor U19623 (N_19623,N_12555,N_18567);
or U19624 (N_19624,N_15707,N_15864);
xnor U19625 (N_19625,N_16871,N_15983);
nand U19626 (N_19626,N_15372,N_15767);
nor U19627 (N_19627,N_12864,N_15626);
xor U19628 (N_19628,N_18079,N_16791);
xor U19629 (N_19629,N_12525,N_16603);
and U19630 (N_19630,N_13100,N_18167);
nor U19631 (N_19631,N_13411,N_15917);
xnor U19632 (N_19632,N_12635,N_15571);
nand U19633 (N_19633,N_17655,N_16285);
nand U19634 (N_19634,N_16784,N_13216);
nor U19635 (N_19635,N_14314,N_18249);
nand U19636 (N_19636,N_15563,N_14051);
nor U19637 (N_19637,N_17768,N_13763);
xor U19638 (N_19638,N_16852,N_13950);
or U19639 (N_19639,N_15699,N_15086);
nand U19640 (N_19640,N_17298,N_12824);
or U19641 (N_19641,N_14090,N_13630);
xnor U19642 (N_19642,N_12600,N_18347);
or U19643 (N_19643,N_17113,N_15405);
and U19644 (N_19644,N_13143,N_17604);
nand U19645 (N_19645,N_15037,N_14177);
and U19646 (N_19646,N_15386,N_14708);
and U19647 (N_19647,N_17839,N_17188);
nand U19648 (N_19648,N_15561,N_18499);
and U19649 (N_19649,N_18256,N_16948);
and U19650 (N_19650,N_13319,N_17830);
or U19651 (N_19651,N_15627,N_16092);
or U19652 (N_19652,N_13523,N_18650);
xor U19653 (N_19653,N_17981,N_13696);
and U19654 (N_19654,N_16452,N_15062);
nand U19655 (N_19655,N_17360,N_18235);
xnor U19656 (N_19656,N_16526,N_14416);
nand U19657 (N_19657,N_17801,N_14126);
xor U19658 (N_19658,N_17471,N_15039);
or U19659 (N_19659,N_16628,N_15954);
and U19660 (N_19660,N_16216,N_18076);
xnor U19661 (N_19661,N_16988,N_16718);
nor U19662 (N_19662,N_14453,N_12990);
and U19663 (N_19663,N_15969,N_15299);
and U19664 (N_19664,N_15073,N_15478);
and U19665 (N_19665,N_18210,N_17755);
or U19666 (N_19666,N_17085,N_12780);
nor U19667 (N_19667,N_18451,N_18192);
xor U19668 (N_19668,N_17332,N_15823);
nor U19669 (N_19669,N_15305,N_14653);
and U19670 (N_19670,N_16087,N_13134);
nand U19671 (N_19671,N_16493,N_18386);
and U19672 (N_19672,N_18223,N_18577);
or U19673 (N_19673,N_13437,N_15295);
nor U19674 (N_19674,N_13301,N_17653);
xnor U19675 (N_19675,N_14654,N_16444);
xnor U19676 (N_19676,N_13074,N_12878);
and U19677 (N_19677,N_15791,N_18144);
and U19678 (N_19678,N_12578,N_12809);
and U19679 (N_19679,N_17963,N_16320);
xnor U19680 (N_19680,N_17199,N_16655);
nor U19681 (N_19681,N_13949,N_14595);
and U19682 (N_19682,N_18213,N_14246);
xnor U19683 (N_19683,N_12930,N_12605);
or U19684 (N_19684,N_12741,N_18682);
nand U19685 (N_19685,N_16135,N_16720);
nand U19686 (N_19686,N_17746,N_16206);
and U19687 (N_19687,N_17042,N_15118);
xor U19688 (N_19688,N_17129,N_13070);
nor U19689 (N_19689,N_16800,N_12849);
xnor U19690 (N_19690,N_13952,N_12514);
nor U19691 (N_19691,N_16975,N_17686);
nor U19692 (N_19692,N_16513,N_17149);
and U19693 (N_19693,N_15247,N_18716);
nand U19694 (N_19694,N_16844,N_16132);
and U19695 (N_19695,N_18269,N_12946);
nand U19696 (N_19696,N_15886,N_18197);
nor U19697 (N_19697,N_17331,N_18376);
and U19698 (N_19698,N_14555,N_13676);
and U19699 (N_19699,N_13361,N_16845);
nand U19700 (N_19700,N_14319,N_18726);
nor U19701 (N_19701,N_14186,N_13897);
nor U19702 (N_19702,N_13076,N_17641);
or U19703 (N_19703,N_12506,N_15818);
nand U19704 (N_19704,N_17171,N_18722);
nor U19705 (N_19705,N_17550,N_14323);
nand U19706 (N_19706,N_14553,N_17973);
xnor U19707 (N_19707,N_16084,N_16798);
nand U19708 (N_19708,N_15353,N_16305);
and U19709 (N_19709,N_18446,N_17361);
and U19710 (N_19710,N_13805,N_14562);
or U19711 (N_19711,N_18190,N_15850);
or U19712 (N_19712,N_14764,N_13006);
nor U19713 (N_19713,N_13493,N_16062);
xnor U19714 (N_19714,N_16420,N_15642);
nor U19715 (N_19715,N_15092,N_18212);
xor U19716 (N_19716,N_13001,N_14642);
nor U19717 (N_19717,N_15452,N_16504);
nand U19718 (N_19718,N_14816,N_13181);
or U19719 (N_19719,N_12770,N_17168);
and U19720 (N_19720,N_18703,N_18630);
nand U19721 (N_19721,N_13576,N_16834);
nand U19722 (N_19722,N_13030,N_17424);
and U19723 (N_19723,N_14369,N_17780);
nand U19724 (N_19724,N_14679,N_15483);
nand U19725 (N_19725,N_13123,N_18687);
and U19726 (N_19726,N_13054,N_14813);
nand U19727 (N_19727,N_14820,N_14865);
xor U19728 (N_19728,N_13908,N_15472);
nand U19729 (N_19729,N_15813,N_14937);
nor U19730 (N_19730,N_16692,N_17543);
xnor U19731 (N_19731,N_14217,N_17162);
or U19732 (N_19732,N_15188,N_15409);
xnor U19733 (N_19733,N_15024,N_17893);
and U19734 (N_19734,N_17947,N_18149);
or U19735 (N_19735,N_14906,N_13416);
nand U19736 (N_19736,N_16386,N_14164);
and U19737 (N_19737,N_14010,N_15166);
and U19738 (N_19738,N_13240,N_15871);
or U19739 (N_19739,N_13383,N_13155);
xor U19740 (N_19740,N_18440,N_15790);
nor U19741 (N_19741,N_16485,N_14315);
or U19742 (N_19742,N_13746,N_14833);
or U19743 (N_19743,N_15534,N_18660);
xor U19744 (N_19744,N_13218,N_15929);
nor U19745 (N_19745,N_14054,N_17661);
nand U19746 (N_19746,N_18248,N_15686);
xnor U19747 (N_19747,N_13081,N_17580);
xor U19748 (N_19748,N_13094,N_16898);
nor U19749 (N_19749,N_14372,N_17760);
nand U19750 (N_19750,N_13965,N_17489);
nand U19751 (N_19751,N_14723,N_14191);
or U19752 (N_19752,N_18106,N_13802);
nor U19753 (N_19753,N_16577,N_18718);
nor U19754 (N_19754,N_15270,N_12623);
or U19755 (N_19755,N_15222,N_15525);
or U19756 (N_19756,N_17187,N_14176);
nor U19757 (N_19757,N_14260,N_14056);
xor U19758 (N_19758,N_18203,N_16632);
xnor U19759 (N_19759,N_17134,N_14807);
or U19760 (N_19760,N_13273,N_12644);
xnor U19761 (N_19761,N_12997,N_15050);
or U19762 (N_19762,N_16582,N_18483);
nand U19763 (N_19763,N_15831,N_13542);
xnor U19764 (N_19764,N_16587,N_13823);
xnor U19765 (N_19765,N_14948,N_16322);
nand U19766 (N_19766,N_13505,N_16330);
or U19767 (N_19767,N_17235,N_17696);
nand U19768 (N_19768,N_18099,N_18293);
nand U19769 (N_19769,N_17238,N_15879);
xnor U19770 (N_19770,N_13840,N_13140);
nor U19771 (N_19771,N_13960,N_14388);
nand U19772 (N_19772,N_13784,N_14824);
or U19773 (N_19773,N_16900,N_15220);
xnor U19774 (N_19774,N_16893,N_13873);
nand U19775 (N_19775,N_15536,N_17848);
nor U19776 (N_19776,N_15877,N_13168);
or U19777 (N_19777,N_15435,N_13757);
nand U19778 (N_19778,N_18697,N_14682);
or U19779 (N_19779,N_12719,N_18646);
and U19780 (N_19780,N_13188,N_14017);
nand U19781 (N_19781,N_16497,N_17455);
xor U19782 (N_19782,N_17855,N_16219);
or U19783 (N_19783,N_17430,N_14989);
and U19784 (N_19784,N_13130,N_13684);
and U19785 (N_19785,N_15899,N_17753);
or U19786 (N_19786,N_16440,N_18472);
nor U19787 (N_19787,N_15219,N_17460);
nor U19788 (N_19788,N_16000,N_14199);
and U19789 (N_19789,N_17378,N_14173);
nand U19790 (N_19790,N_17300,N_16855);
nand U19791 (N_19791,N_18397,N_14966);
or U19792 (N_19792,N_13159,N_14673);
nor U19793 (N_19793,N_17646,N_13171);
xor U19794 (N_19794,N_13571,N_17462);
nor U19795 (N_19795,N_13722,N_15210);
and U19796 (N_19796,N_14118,N_17095);
xnor U19797 (N_19797,N_17733,N_12976);
and U19798 (N_19798,N_13469,N_18239);
or U19799 (N_19799,N_15497,N_17860);
xor U19800 (N_19800,N_17396,N_13752);
nand U19801 (N_19801,N_13883,N_16412);
nor U19802 (N_19802,N_15892,N_12579);
xor U19803 (N_19803,N_14835,N_13616);
nand U19804 (N_19804,N_12552,N_14022);
nand U19805 (N_19805,N_16259,N_14774);
nor U19806 (N_19806,N_14942,N_15341);
nand U19807 (N_19807,N_14742,N_12987);
or U19808 (N_19808,N_12577,N_17651);
or U19809 (N_19809,N_16081,N_15016);
and U19810 (N_19810,N_18285,N_12505);
nor U19811 (N_19811,N_13807,N_16860);
or U19812 (N_19812,N_16202,N_16146);
xor U19813 (N_19813,N_13392,N_15845);
or U19814 (N_19814,N_12647,N_16423);
nand U19815 (N_19815,N_16584,N_12853);
nand U19816 (N_19816,N_13419,N_17982);
and U19817 (N_19817,N_17194,N_17685);
or U19818 (N_19818,N_13992,N_15066);
xor U19819 (N_19819,N_16498,N_13243);
or U19820 (N_19820,N_13668,N_14620);
or U19821 (N_19821,N_17245,N_18385);
and U19822 (N_19822,N_13787,N_18343);
nor U19823 (N_19823,N_15215,N_16250);
nor U19824 (N_19824,N_15742,N_17928);
nand U19825 (N_19825,N_15275,N_14769);
or U19826 (N_19826,N_13681,N_17315);
and U19827 (N_19827,N_18121,N_16231);
xor U19828 (N_19828,N_14926,N_13624);
or U19829 (N_19829,N_17229,N_13866);
xor U19830 (N_19830,N_12652,N_16608);
nor U19831 (N_19831,N_14997,N_16611);
or U19832 (N_19832,N_16947,N_15857);
nand U19833 (N_19833,N_14193,N_13906);
or U19834 (N_19834,N_18300,N_15263);
or U19835 (N_19835,N_16679,N_18706);
nand U19836 (N_19836,N_14539,N_16284);
or U19837 (N_19837,N_16443,N_13212);
and U19838 (N_19838,N_14312,N_17190);
and U19839 (N_19839,N_14433,N_15143);
nor U19840 (N_19840,N_18535,N_15575);
and U19841 (N_19841,N_16662,N_15248);
and U19842 (N_19842,N_14856,N_12749);
or U19843 (N_19843,N_15481,N_15359);
nand U19844 (N_19844,N_14479,N_14860);
nor U19845 (N_19845,N_16474,N_18470);
or U19846 (N_19846,N_15747,N_12802);
and U19847 (N_19847,N_12972,N_16210);
nor U19848 (N_19848,N_12929,N_14473);
and U19849 (N_19849,N_14727,N_16618);
xnor U19850 (N_19850,N_18108,N_12828);
nand U19851 (N_19851,N_18240,N_14297);
nand U19852 (N_19852,N_13792,N_12955);
xor U19853 (N_19853,N_17470,N_17968);
nand U19854 (N_19854,N_15580,N_16255);
nand U19855 (N_19855,N_13727,N_16458);
and U19856 (N_19856,N_17805,N_18504);
and U19857 (N_19857,N_13368,N_13299);
nor U19858 (N_19858,N_12794,N_14591);
nor U19859 (N_19859,N_16019,N_13068);
xor U19860 (N_19860,N_13644,N_16099);
nor U19861 (N_19861,N_17898,N_17476);
or U19862 (N_19862,N_15656,N_14082);
and U19863 (N_19863,N_15074,N_17637);
or U19864 (N_19864,N_14198,N_14763);
or U19865 (N_19865,N_15115,N_12681);
or U19866 (N_19866,N_16738,N_13204);
xnor U19867 (N_19867,N_16093,N_15682);
or U19868 (N_19868,N_16660,N_18428);
nand U19869 (N_19869,N_13653,N_16786);
xor U19870 (N_19870,N_14670,N_18196);
nand U19871 (N_19871,N_15729,N_16675);
or U19872 (N_19872,N_12840,N_18471);
nor U19873 (N_19873,N_15049,N_16841);
nor U19874 (N_19874,N_16347,N_13287);
nand U19875 (N_19875,N_15241,N_14693);
nand U19876 (N_19876,N_14437,N_17458);
and U19877 (N_19877,N_15177,N_17705);
and U19878 (N_19878,N_13626,N_14882);
xor U19879 (N_19879,N_18170,N_13983);
nand U19880 (N_19880,N_12940,N_18232);
and U19881 (N_19881,N_18031,N_15728);
and U19882 (N_19882,N_17854,N_13793);
or U19883 (N_19883,N_18138,N_18262);
xnor U19884 (N_19884,N_16377,N_13112);
nand U19885 (N_19885,N_17008,N_16469);
xor U19886 (N_19886,N_18668,N_15415);
nor U19887 (N_19887,N_13298,N_12767);
and U19888 (N_19888,N_16568,N_15462);
and U19889 (N_19889,N_12856,N_18663);
nand U19890 (N_19890,N_13601,N_15711);
nand U19891 (N_19891,N_15209,N_14289);
or U19892 (N_19892,N_13592,N_14008);
nand U19893 (N_19893,N_15749,N_16433);
nand U19894 (N_19894,N_16185,N_13095);
or U19895 (N_19895,N_18514,N_14489);
nand U19896 (N_19896,N_13652,N_17929);
nand U19897 (N_19897,N_18252,N_15968);
or U19898 (N_19898,N_15987,N_14155);
nand U19899 (N_19899,N_16622,N_14612);
xor U19900 (N_19900,N_13560,N_16546);
xor U19901 (N_19901,N_15420,N_16351);
xor U19902 (N_19902,N_15669,N_12658);
nand U19903 (N_19903,N_16810,N_12969);
or U19904 (N_19904,N_12758,N_16749);
nand U19905 (N_19905,N_13761,N_16094);
nor U19906 (N_19906,N_16367,N_18086);
nand U19907 (N_19907,N_15357,N_13872);
and U19908 (N_19908,N_16551,N_13314);
nor U19909 (N_19909,N_17820,N_17092);
xor U19910 (N_19910,N_16448,N_12639);
or U19911 (N_19911,N_16685,N_16126);
and U19912 (N_19912,N_14340,N_18592);
and U19913 (N_19913,N_17914,N_14237);
and U19914 (N_19914,N_17172,N_14272);
and U19915 (N_19915,N_14488,N_12581);
xor U19916 (N_19916,N_12934,N_18189);
and U19917 (N_19917,N_14495,N_16462);
or U19918 (N_19918,N_14884,N_17865);
nor U19919 (N_19919,N_13105,N_13425);
and U19920 (N_19920,N_18357,N_18596);
or U19921 (N_19921,N_17875,N_16407);
or U19922 (N_19922,N_18544,N_16964);
or U19923 (N_19923,N_13378,N_12587);
nand U19924 (N_19924,N_18016,N_17174);
or U19925 (N_19925,N_13291,N_13206);
or U19926 (N_19926,N_15013,N_17811);
xor U19927 (N_19927,N_14139,N_12617);
nor U19928 (N_19928,N_17959,N_13222);
nor U19929 (N_19929,N_16278,N_13744);
xnor U19930 (N_19930,N_17276,N_12629);
nand U19931 (N_19931,N_16449,N_14890);
nor U19932 (N_19932,N_16529,N_16941);
nand U19933 (N_19933,N_14748,N_14042);
xnor U19934 (N_19934,N_13228,N_15431);
nand U19935 (N_19935,N_16007,N_15198);
and U19936 (N_19936,N_16612,N_16451);
xor U19937 (N_19937,N_15205,N_18214);
or U19938 (N_19938,N_18528,N_15853);
xor U19939 (N_19939,N_13268,N_13479);
or U19940 (N_19940,N_14680,N_14285);
nand U19941 (N_19941,N_16188,N_18430);
nor U19942 (N_19942,N_16104,N_12615);
xnor U19943 (N_19943,N_18032,N_12991);
and U19944 (N_19944,N_13217,N_14011);
and U19945 (N_19945,N_17189,N_16023);
and U19946 (N_19946,N_13178,N_15058);
or U19947 (N_19947,N_13250,N_14248);
and U19948 (N_19948,N_16158,N_13021);
nand U19949 (N_19949,N_15192,N_16304);
or U19950 (N_19950,N_16544,N_17138);
xor U19951 (N_19951,N_14546,N_13765);
or U19952 (N_19952,N_14678,N_13346);
xor U19953 (N_19953,N_14385,N_18485);
xnor U19954 (N_19954,N_15562,N_12764);
nand U19955 (N_19955,N_16969,N_15057);
and U19956 (N_19956,N_17514,N_15542);
xnor U19957 (N_19957,N_14093,N_15051);
and U19958 (N_19958,N_14921,N_13528);
xnor U19959 (N_19959,N_14356,N_17061);
nand U19960 (N_19960,N_17338,N_16227);
nand U19961 (N_19961,N_16506,N_16864);
xor U19962 (N_19962,N_15370,N_14998);
xor U19963 (N_19963,N_12833,N_12518);
or U19964 (N_19964,N_18092,N_15154);
or U19965 (N_19965,N_15399,N_18169);
nand U19966 (N_19966,N_15242,N_14836);
and U19967 (N_19967,N_12941,N_18619);
or U19968 (N_19968,N_13139,N_18166);
and U19969 (N_19969,N_13489,N_18373);
and U19970 (N_19970,N_12549,N_13832);
or U19971 (N_19971,N_16985,N_13799);
nor U19972 (N_19972,N_16511,N_16847);
nand U19973 (N_19973,N_14754,N_14900);
and U19974 (N_19974,N_13979,N_14105);
xor U19975 (N_19975,N_15690,N_18156);
and U19976 (N_19976,N_17806,N_17849);
xnor U19977 (N_19977,N_16049,N_14135);
and U19978 (N_19978,N_14484,N_18087);
nand U19979 (N_19979,N_18396,N_13335);
nor U19980 (N_19980,N_14827,N_18447);
or U19981 (N_19981,N_17071,N_15466);
or U19982 (N_19982,N_15671,N_14338);
and U19983 (N_19983,N_13512,N_17407);
nand U19984 (N_19984,N_14471,N_17967);
nor U19985 (N_19985,N_17492,N_18566);
xor U19986 (N_19986,N_16400,N_12524);
nor U19987 (N_19987,N_15814,N_14847);
or U19988 (N_19988,N_13245,N_16606);
and U19989 (N_19989,N_13012,N_17443);
xnor U19990 (N_19990,N_14603,N_14628);
xor U19991 (N_19991,N_18234,N_16865);
nand U19992 (N_19992,N_17352,N_16771);
or U19993 (N_19993,N_17890,N_16200);
xor U19994 (N_19994,N_16115,N_13031);
nor U19995 (N_19995,N_18593,N_18512);
nor U19996 (N_19996,N_17775,N_17342);
xnor U19997 (N_19997,N_16060,N_17953);
or U19998 (N_19998,N_17858,N_14637);
nor U19999 (N_19999,N_18689,N_12964);
nor U20000 (N_20000,N_16812,N_15156);
nand U20001 (N_20001,N_18462,N_14840);
nor U20002 (N_20002,N_15448,N_17804);
xor U20003 (N_20003,N_14275,N_16374);
nor U20004 (N_20004,N_14304,N_18044);
nand U20005 (N_20005,N_17627,N_13773);
and U20006 (N_20006,N_14062,N_17681);
xnor U20007 (N_20007,N_17435,N_18046);
nand U20008 (N_20008,N_18420,N_16705);
nor U20009 (N_20009,N_17906,N_15419);
nor U20010 (N_20010,N_13261,N_13008);
nor U20011 (N_20011,N_15500,N_16894);
or U20012 (N_20012,N_18742,N_14718);
and U20013 (N_20013,N_15894,N_14171);
and U20014 (N_20014,N_15594,N_16657);
nor U20015 (N_20015,N_13887,N_16591);
nand U20016 (N_20016,N_15296,N_16058);
nand U20017 (N_20017,N_16148,N_17566);
nor U20018 (N_20018,N_14829,N_17776);
nor U20019 (N_20019,N_16658,N_17821);
and U20020 (N_20020,N_18225,N_14873);
nor U20021 (N_20021,N_16173,N_17195);
xor U20022 (N_20022,N_12717,N_15731);
nor U20023 (N_20023,N_14456,N_18116);
xnor U20024 (N_20024,N_13695,N_18579);
nand U20025 (N_20025,N_15303,N_14914);
or U20026 (N_20026,N_13530,N_14038);
and U20027 (N_20027,N_18104,N_18665);
nand U20028 (N_20028,N_16849,N_14387);
or U20029 (N_20029,N_13820,N_15443);
xor U20030 (N_20030,N_18177,N_15951);
nand U20031 (N_20031,N_18281,N_14466);
nor U20032 (N_20032,N_17795,N_16100);
xor U20033 (N_20033,N_17305,N_13366);
nand U20034 (N_20034,N_17586,N_17937);
nand U20035 (N_20035,N_15234,N_14478);
and U20036 (N_20036,N_12839,N_16417);
nor U20037 (N_20037,N_18348,N_12726);
and U20038 (N_20038,N_15836,N_17286);
nor U20039 (N_20039,N_16155,N_13636);
nand U20040 (N_20040,N_15901,N_15543);
xnor U20041 (N_20041,N_14069,N_17059);
xnor U20042 (N_20042,N_14050,N_17955);
nor U20043 (N_20043,N_15846,N_18436);
nand U20044 (N_20044,N_16054,N_15623);
xnor U20045 (N_20045,N_17170,N_15064);
xor U20046 (N_20046,N_17781,N_13406);
nand U20047 (N_20047,N_17989,N_16911);
and U20048 (N_20048,N_17328,N_12938);
or U20049 (N_20049,N_16597,N_15366);
nand U20050 (N_20050,N_16334,N_16590);
nor U20051 (N_20051,N_18602,N_17241);
nor U20052 (N_20052,N_13978,N_15668);
nand U20053 (N_20053,N_13317,N_18007);
nand U20054 (N_20054,N_17488,N_15649);
or U20055 (N_20055,N_17272,N_14160);
nor U20056 (N_20056,N_12529,N_15433);
nor U20057 (N_20057,N_15345,N_15944);
or U20058 (N_20058,N_16695,N_15463);
or U20059 (N_20059,N_16430,N_15304);
nor U20060 (N_20060,N_12596,N_15865);
nor U20061 (N_20061,N_15468,N_15638);
or U20062 (N_20062,N_18057,N_14993);
xnor U20063 (N_20063,N_14424,N_18224);
nand U20064 (N_20064,N_14281,N_15514);
and U20065 (N_20065,N_15218,N_14893);
or U20066 (N_20066,N_18621,N_16972);
xor U20067 (N_20067,N_15629,N_16933);
xor U20068 (N_20068,N_18344,N_17441);
nor U20069 (N_20069,N_17362,N_13449);
xor U20070 (N_20070,N_15633,N_15524);
nand U20071 (N_20071,N_14422,N_16825);
nand U20072 (N_20072,N_15307,N_15774);
or U20073 (N_20073,N_13158,N_17721);
xor U20074 (N_20074,N_16763,N_15223);
nand U20075 (N_20075,N_15986,N_14614);
or U20076 (N_20076,N_17769,N_13272);
or U20077 (N_20077,N_13279,N_12844);
xor U20078 (N_20078,N_16761,N_13729);
xnor U20079 (N_20079,N_17726,N_17743);
and U20080 (N_20080,N_12886,N_17393);
nor U20081 (N_20081,N_12612,N_18475);
nor U20082 (N_20082,N_16212,N_17118);
nor U20083 (N_20083,N_17757,N_13847);
xor U20084 (N_20084,N_17203,N_18531);
nand U20085 (N_20085,N_18261,N_16596);
and U20086 (N_20086,N_18114,N_13517);
nand U20087 (N_20087,N_15637,N_14787);
nor U20088 (N_20088,N_12936,N_12779);
and U20089 (N_20089,N_14292,N_12597);
or U20090 (N_20090,N_15099,N_12883);
or U20091 (N_20091,N_13656,N_13170);
nor U20092 (N_20092,N_13251,N_15351);
xor U20093 (N_20093,N_17410,N_15147);
xor U20094 (N_20094,N_15164,N_12531);
nor U20095 (N_20095,N_13429,N_17032);
or U20096 (N_20096,N_12665,N_18231);
xor U20097 (N_20097,N_17522,N_17103);
or U20098 (N_20098,N_13290,N_15998);
nor U20099 (N_20099,N_18199,N_12752);
or U20100 (N_20100,N_16599,N_18638);
and U20101 (N_20101,N_16105,N_15547);
nor U20102 (N_20102,N_13567,N_12621);
nor U20103 (N_20103,N_14114,N_13779);
xor U20104 (N_20104,N_16082,N_15734);
nand U20105 (N_20105,N_18061,N_16926);
nand U20106 (N_20106,N_18661,N_15936);
xnor U20107 (N_20107,N_16617,N_14308);
nor U20108 (N_20108,N_16350,N_16072);
or U20109 (N_20109,N_16358,N_14790);
nand U20110 (N_20110,N_16916,N_16492);
or U20111 (N_20111,N_18089,N_15959);
and U20112 (N_20112,N_17823,N_15570);
xor U20113 (N_20113,N_16258,N_17427);
xor U20114 (N_20114,N_18552,N_14430);
nor U20115 (N_20115,N_16813,N_15065);
and U20116 (N_20116,N_12683,N_17556);
nor U20117 (N_20117,N_13620,N_16287);
xor U20118 (N_20118,N_15593,N_17828);
and U20119 (N_20119,N_15320,N_17278);
and U20120 (N_20120,N_14541,N_17110);
or U20121 (N_20121,N_18341,N_16161);
and U20122 (N_20122,N_16207,N_15416);
xor U20123 (N_20123,N_13042,N_13427);
nand U20124 (N_20124,N_17971,N_13825);
and U20125 (N_20125,N_16066,N_13309);
or U20126 (N_20126,N_15801,N_15268);
xor U20127 (N_20127,N_15474,N_12573);
nand U20128 (N_20128,N_12875,N_18097);
xnor U20129 (N_20129,N_12512,N_17397);
and U20130 (N_20130,N_16409,N_18469);
and U20131 (N_20131,N_12762,N_18304);
xnor U20132 (N_20132,N_13141,N_13734);
xnor U20133 (N_20133,N_14089,N_16071);
and U20134 (N_20134,N_17559,N_18439);
or U20135 (N_20135,N_13917,N_16940);
xor U20136 (N_20136,N_16491,N_16829);
nor U20137 (N_20137,N_17737,N_13855);
or U20138 (N_20138,N_15467,N_17844);
and U20139 (N_20139,N_17871,N_15395);
and U20140 (N_20140,N_15233,N_12884);
and U20141 (N_20141,N_17923,N_14517);
xor U20142 (N_20142,N_16886,N_13483);
or U20143 (N_20143,N_14655,N_15924);
or U20144 (N_20144,N_14293,N_15772);
and U20145 (N_20145,N_17613,N_17232);
and U20146 (N_20146,N_16224,N_16244);
or U20147 (N_20147,N_12712,N_13000);
xnor U20148 (N_20148,N_16959,N_16383);
nor U20149 (N_20149,N_17322,N_16249);
xnor U20150 (N_20150,N_16387,N_16397);
nand U20151 (N_20151,N_17529,N_12584);
or U20152 (N_20152,N_15190,N_16598);
nor U20153 (N_20153,N_18570,N_14608);
or U20154 (N_20154,N_15589,N_17617);
or U20155 (N_20155,N_14460,N_17744);
or U20156 (N_20156,N_18154,N_16047);
nor U20157 (N_20157,N_13575,N_17602);
xor U20158 (N_20158,N_16248,N_14792);
xor U20159 (N_20159,N_14530,N_16951);
nor U20160 (N_20160,N_16098,N_13220);
nor U20161 (N_20161,N_17414,N_13638);
xnor U20162 (N_20162,N_14459,N_13384);
xor U20163 (N_20163,N_17626,N_17960);
and U20164 (N_20164,N_16257,N_16043);
and U20165 (N_20165,N_14441,N_16694);
nor U20166 (N_20166,N_13161,N_15718);
xnor U20167 (N_20167,N_15907,N_17446);
or U20168 (N_20168,N_17930,N_14751);
nand U20169 (N_20169,N_16740,N_16269);
and U20170 (N_20170,N_18332,N_15870);
nor U20171 (N_20171,N_15186,N_18251);
or U20172 (N_20172,N_18731,N_18686);
and U20173 (N_20173,N_15269,N_14337);
xor U20174 (N_20174,N_13911,N_14213);
or U20175 (N_20175,N_17874,N_13688);
nor U20176 (N_20176,N_13548,N_14053);
nand U20177 (N_20177,N_17984,N_13495);
or U20178 (N_20178,N_18674,N_13438);
nor U20179 (N_20179,N_14828,N_15083);
nor U20180 (N_20180,N_13602,N_18693);
xor U20181 (N_20181,N_17908,N_15895);
nor U20182 (N_20182,N_16843,N_15528);
and U20183 (N_20183,N_13085,N_15172);
or U20184 (N_20184,N_14854,N_17642);
nor U20185 (N_20185,N_17074,N_13726);
or U20186 (N_20186,N_14239,N_18503);
xor U20187 (N_20187,N_18489,N_15048);
xnor U20188 (N_20188,N_14503,N_17145);
nor U20189 (N_20189,N_15702,N_13749);
nand U20190 (N_20190,N_17882,N_15828);
or U20191 (N_20191,N_14170,N_12829);
nand U20192 (N_20192,N_17425,N_17091);
and U20193 (N_20193,N_14697,N_13236);
nor U20194 (N_20194,N_13434,N_14812);
xnor U20195 (N_20195,N_18028,N_17585);
nand U20196 (N_20196,N_18500,N_13088);
or U20197 (N_20197,N_12766,N_14001);
nand U20198 (N_20198,N_17390,N_16583);
xnor U20199 (N_20199,N_17499,N_17041);
nor U20200 (N_20200,N_16540,N_16575);
and U20201 (N_20201,N_17903,N_15825);
xor U20202 (N_20202,N_12914,N_17344);
nand U20203 (N_20203,N_14457,N_12543);
nand U20204 (N_20204,N_18371,N_13963);
nor U20205 (N_20205,N_15189,N_16308);
and U20206 (N_20206,N_16918,N_18468);
xor U20207 (N_20207,N_12560,N_12944);
nor U20208 (N_20208,N_12703,N_18406);
and U20209 (N_20209,N_14560,N_15289);
or U20210 (N_20210,N_14845,N_14615);
or U20211 (N_20211,N_17202,N_16295);
nor U20212 (N_20212,N_17700,N_18627);
nand U20213 (N_20213,N_13502,N_13096);
nor U20214 (N_20214,N_15918,N_15458);
nand U20215 (N_20215,N_14180,N_18185);
and U20216 (N_20216,N_15666,N_17394);
nor U20217 (N_20217,N_16636,N_13637);
or U20218 (N_20218,N_13835,N_14165);
nor U20219 (N_20219,N_16986,N_13476);
or U20220 (N_20220,N_14104,N_14739);
nor U20221 (N_20221,N_17475,N_12680);
xnor U20222 (N_20222,N_13265,N_18301);
or U20223 (N_20223,N_17067,N_13433);
nand U20224 (N_20224,N_18434,N_16280);
or U20225 (N_20225,N_15407,N_16782);
nand U20226 (N_20226,N_16214,N_13249);
xor U20227 (N_20227,N_18708,N_18329);
xor U20228 (N_20228,N_16059,N_13875);
xor U20229 (N_20229,N_15616,N_17254);
or U20230 (N_20230,N_12924,N_18743);
nand U20231 (N_20231,N_12657,N_16343);
or U20232 (N_20232,N_17810,N_12898);
or U20233 (N_20233,N_16518,N_12789);
or U20234 (N_20234,N_17612,N_16700);
nand U20235 (N_20235,N_14785,N_14026);
xor U20236 (N_20236,N_12793,N_14881);
and U20237 (N_20237,N_13264,N_16888);
nor U20238 (N_20238,N_14949,N_14892);
nand U20239 (N_20239,N_14075,N_12515);
and U20240 (N_20240,N_13322,N_15012);
xnor U20241 (N_20241,N_16467,N_18501);
nand U20242 (N_20242,N_18229,N_13399);
xor U20243 (N_20243,N_13398,N_13108);
nor U20244 (N_20244,N_13870,N_16321);
xor U20245 (N_20245,N_17719,N_18546);
and U20246 (N_20246,N_17557,N_15685);
and U20247 (N_20247,N_17137,N_13342);
nor U20248 (N_20248,N_17372,N_17750);
or U20249 (N_20249,N_12812,N_15029);
or U20250 (N_20250,N_16626,N_13851);
or U20251 (N_20251,N_14179,N_14442);
or U20252 (N_20252,N_16152,N_16709);
or U20253 (N_20253,N_14476,N_13532);
xnor U20254 (N_20254,N_15490,N_15291);
nand U20255 (N_20255,N_16876,N_18309);
nand U20256 (N_20256,N_14616,N_14327);
or U20257 (N_20257,N_14354,N_13116);
nor U20258 (N_20258,N_17574,N_17494);
nor U20259 (N_20259,N_16689,N_12935);
xnor U20260 (N_20260,N_15461,N_14709);
nor U20261 (N_20261,N_17652,N_17035);
or U20262 (N_20262,N_16379,N_13418);
or U20263 (N_20263,N_18676,N_17748);
nor U20264 (N_20264,N_12754,N_13998);
nand U20265 (N_20265,N_15315,N_14733);
xor U20266 (N_20266,N_17029,N_16851);
xor U20267 (N_20267,N_16112,N_16868);
xor U20268 (N_20268,N_17767,N_13690);
nor U20269 (N_20269,N_15581,N_17658);
xor U20270 (N_20270,N_13360,N_15511);
or U20271 (N_20271,N_14919,N_17783);
or U20272 (N_20272,N_12826,N_17350);
nor U20273 (N_20273,N_18159,N_15148);
xnor U20274 (N_20274,N_15957,N_16907);
nand U20275 (N_20275,N_15819,N_13331);
nand U20276 (N_20276,N_15336,N_17940);
xnor U20277 (N_20277,N_16764,N_18129);
or U20278 (N_20278,N_18273,N_14241);
xor U20279 (N_20279,N_15840,N_14137);
and U20280 (N_20280,N_12513,N_13957);
nand U20281 (N_20281,N_15281,N_18383);
or U20282 (N_20282,N_13446,N_14461);
or U20283 (N_20283,N_16017,N_13432);
nand U20284 (N_20284,N_16124,N_13913);
nand U20285 (N_20285,N_13973,N_16096);
or U20286 (N_20286,N_16505,N_12788);
or U20287 (N_20287,N_14264,N_15445);
or U20288 (N_20288,N_14201,N_16095);
nor U20289 (N_20289,N_14721,N_14167);
nor U20290 (N_20290,N_13959,N_14013);
nand U20291 (N_20291,N_12672,N_12966);
or U20292 (N_20292,N_16704,N_16581);
and U20293 (N_20293,N_16484,N_15884);
nand U20294 (N_20294,N_16666,N_18474);
xor U20295 (N_20295,N_12569,N_12899);
and U20296 (N_20296,N_16370,N_15974);
or U20297 (N_20297,N_13373,N_13519);
nand U20298 (N_20298,N_16240,N_14224);
or U20299 (N_20299,N_13403,N_13073);
or U20300 (N_20300,N_17990,N_15860);
and U20301 (N_20301,N_15456,N_13989);
or U20302 (N_20302,N_14924,N_12958);
or U20303 (N_20303,N_14046,N_14358);
or U20304 (N_20304,N_14749,N_16977);
xor U20305 (N_20305,N_15134,N_15491);
xor U20306 (N_20306,N_14427,N_18672);
nand U20307 (N_20307,N_18522,N_17868);
nor U20308 (N_20308,N_14954,N_17224);
nand U20309 (N_20309,N_18172,N_18616);
or U20310 (N_20310,N_14757,N_13410);
nor U20311 (N_20311,N_18419,N_13697);
nor U20312 (N_20312,N_16077,N_12622);
and U20313 (N_20313,N_15155,N_18247);
nand U20314 (N_20314,N_12797,N_13464);
xor U20315 (N_20315,N_14212,N_16496);
xnor U20316 (N_20316,N_13463,N_12763);
and U20317 (N_20317,N_12989,N_18649);
xor U20318 (N_20318,N_17152,N_14685);
nor U20319 (N_20319,N_15042,N_17702);
nand U20320 (N_20320,N_12921,N_14802);
nand U20321 (N_20321,N_17117,N_16441);
nor U20322 (N_20322,N_18734,N_15300);
and U20323 (N_20323,N_15723,N_16687);
nor U20324 (N_20324,N_12896,N_14520);
nand U20325 (N_20325,N_14009,N_14762);
xnor U20326 (N_20326,N_12755,N_17070);
nor U20327 (N_20327,N_15056,N_14197);
nor U20328 (N_20328,N_12715,N_15937);
or U20329 (N_20329,N_18530,N_12656);
xnor U20330 (N_20330,N_13938,N_12723);
xnor U20331 (N_20331,N_17060,N_18286);
or U20332 (N_20332,N_15513,N_17016);
and U20333 (N_20333,N_14096,N_14990);
nor U20334 (N_20334,N_12803,N_14343);
nor U20335 (N_20335,N_15622,N_17978);
and U20336 (N_20336,N_12882,N_17457);
nor U20337 (N_20337,N_17962,N_13165);
and U20338 (N_20338,N_14959,N_12563);
nand U20339 (N_20339,N_18640,N_18207);
xor U20340 (N_20340,N_13455,N_14068);
and U20341 (N_20341,N_13215,N_17803);
and U20342 (N_20342,N_18545,N_12690);
and U20343 (N_20343,N_17552,N_13407);
and U20344 (N_20344,N_15485,N_18542);
and U20345 (N_20345,N_15397,N_15332);
nor U20346 (N_20346,N_17807,N_13953);
and U20347 (N_20347,N_17977,N_14781);
xnor U20348 (N_20348,N_17031,N_13889);
nand U20349 (N_20349,N_14904,N_13737);
nand U20350 (N_20350,N_17833,N_13815);
xor U20351 (N_20351,N_14776,N_13801);
or U20352 (N_20352,N_14468,N_14124);
nand U20353 (N_20353,N_12835,N_14577);
and U20354 (N_20354,N_15330,N_16716);
or U20355 (N_20355,N_15556,N_18389);
and U20356 (N_20356,N_15888,N_16724);
nand U20357 (N_20357,N_17964,N_15095);
or U20358 (N_20358,N_13467,N_17038);
nor U20359 (N_20359,N_14397,N_17371);
nand U20360 (N_20360,N_15212,N_17829);
and U20361 (N_20361,N_14797,N_14294);
or U20362 (N_20362,N_16040,N_15515);
and U20363 (N_20363,N_18595,N_16357);
and U20364 (N_20364,N_14420,N_18387);
nand U20365 (N_20365,N_17747,N_17921);
and U20366 (N_20366,N_16880,N_13924);
nand U20367 (N_20367,N_17738,N_14196);
xor U20368 (N_20368,N_17822,N_17160);
and U20369 (N_20369,N_16576,N_15271);
xnor U20370 (N_20370,N_16041,N_13896);
and U20371 (N_20371,N_16253,N_12862);
nor U20372 (N_20372,N_14287,N_13809);
and U20373 (N_20373,N_16991,N_15777);
xor U20374 (N_20374,N_18723,N_15807);
nand U20375 (N_20375,N_13846,N_15952);
nand U20376 (N_20376,N_16262,N_14740);
and U20377 (N_20377,N_15568,N_14410);
or U20378 (N_20378,N_18005,N_16147);
nor U20379 (N_20379,N_12664,N_17725);
nand U20380 (N_20380,N_12757,N_17945);
and U20381 (N_20381,N_12575,N_17473);
xor U20382 (N_20382,N_13816,N_16792);
nand U20383 (N_20383,N_13677,N_12994);
nand U20384 (N_20384,N_14381,N_13907);
and U20385 (N_20385,N_13160,N_15319);
nor U20386 (N_20386,N_14657,N_15183);
or U20387 (N_20387,N_17589,N_16190);
nand U20388 (N_20388,N_13508,N_17126);
nor U20389 (N_20389,N_17409,N_15947);
or U20390 (N_20390,N_18160,N_15732);
nand U20391 (N_20391,N_13284,N_15312);
xor U20392 (N_20392,N_17123,N_12692);
nand U20393 (N_20393,N_12697,N_16303);
nand U20394 (N_20394,N_14945,N_15751);
and U20395 (N_20395,N_17950,N_13422);
xor U20396 (N_20396,N_18278,N_18065);
or U20397 (N_20397,N_18534,N_16201);
xnor U20398 (N_20398,N_17218,N_16604);
or U20399 (N_20399,N_18233,N_13315);
nand U20400 (N_20400,N_14641,N_13937);
or U20401 (N_20401,N_17323,N_12568);
and U20402 (N_20402,N_16203,N_16063);
nand U20403 (N_20403,N_17956,N_16555);
nor U20404 (N_20404,N_14850,N_13892);
nand U20405 (N_20405,N_13238,N_14037);
nand U20406 (N_20406,N_12718,N_13369);
nand U20407 (N_20407,N_17451,N_16751);
xnor U20408 (N_20408,N_13271,N_16475);
xnor U20409 (N_20409,N_16488,N_18670);
nor U20410 (N_20410,N_15778,N_17233);
nor U20411 (N_20411,N_17598,N_14576);
xor U20412 (N_20412,N_15804,N_15883);
nor U20413 (N_20413,N_15502,N_18636);
and U20414 (N_20414,N_14147,N_16461);
or U20415 (N_20415,N_17230,N_16481);
and U20416 (N_20416,N_13651,N_17153);
nand U20417 (N_20417,N_14329,N_15798);
nor U20418 (N_20418,N_15503,N_17339);
nor U20419 (N_20419,N_13163,N_18253);
xnor U20420 (N_20420,N_18068,N_15541);
nand U20421 (N_20421,N_16654,N_14194);
xor U20422 (N_20422,N_14544,N_14299);
xnor U20423 (N_20423,N_18608,N_14151);
xor U20424 (N_20424,N_18572,N_16641);
nand U20425 (N_20425,N_17708,N_15214);
xor U20426 (N_20426,N_13089,N_14440);
nand U20427 (N_20427,N_13818,N_12888);
xor U20428 (N_20428,N_12879,N_15158);
xnor U20429 (N_20429,N_15087,N_13036);
and U20430 (N_20430,N_13595,N_15905);
nor U20431 (N_20431,N_14571,N_18055);
and U20432 (N_20432,N_13044,N_18575);
nand U20433 (N_20433,N_18297,N_12609);
and U20434 (N_20434,N_14547,N_15687);
nor U20435 (N_20435,N_18720,N_14274);
nor U20436 (N_20436,N_13424,N_15488);
xnor U20437 (N_20437,N_17363,N_17147);
nor U20438 (N_20438,N_18299,N_18056);
or U20439 (N_20439,N_15965,N_17319);
nor U20440 (N_20440,N_15402,N_15329);
nor U20441 (N_20441,N_15459,N_13798);
xnor U20442 (N_20442,N_16961,N_17988);
nor U20443 (N_20443,N_13371,N_13009);
or U20444 (N_20444,N_17662,N_15279);
nor U20445 (N_20445,N_18733,N_17318);
xnor U20446 (N_20446,N_18391,N_15373);
xor U20447 (N_20447,N_18072,N_16361);
or U20448 (N_20448,N_13351,N_18084);
and U20449 (N_20449,N_13488,N_13172);
nand U20450 (N_20450,N_18161,N_18358);
nor U20451 (N_20451,N_16175,N_18287);
nand U20452 (N_20452,N_17796,N_12567);
nand U20453 (N_20453,N_14692,N_13912);
nand U20454 (N_20454,N_13742,N_16811);
or U20455 (N_20455,N_14898,N_13231);
or U20456 (N_20456,N_16215,N_12669);
nor U20457 (N_20457,N_17288,N_14012);
nand U20458 (N_20458,N_14039,N_13043);
xor U20459 (N_20459,N_16282,N_12963);
xor U20460 (N_20460,N_18110,N_15132);
or U20461 (N_20461,N_16428,N_15317);
or U20462 (N_20462,N_13016,N_13415);
nand U20463 (N_20463,N_14761,N_14487);
or U20464 (N_20464,N_12731,N_16937);
nand U20465 (N_20465,N_17434,N_18695);
nand U20466 (N_20466,N_18314,N_15262);
or U20467 (N_20467,N_12804,N_13263);
and U20468 (N_20468,N_18587,N_14034);
nor U20469 (N_20469,N_14765,N_15128);
or U20470 (N_20470,N_16180,N_15126);
nand U20471 (N_20471,N_15333,N_15558);
xor U20472 (N_20472,N_16846,N_18553);
nor U20473 (N_20473,N_16348,N_15486);
nor U20474 (N_20474,N_15549,N_17253);
nor U20475 (N_20475,N_15769,N_13278);
nand U20476 (N_20476,N_15047,N_13047);
xnor U20477 (N_20477,N_13496,N_17293);
xnor U20478 (N_20478,N_13117,N_16723);
nand U20479 (N_20479,N_16802,N_18709);
nand U20480 (N_20480,N_14454,N_13538);
or U20481 (N_20481,N_16086,N_17265);
nor U20482 (N_20482,N_15910,N_18654);
or U20483 (N_20483,N_15882,N_16633);
or U20484 (N_20484,N_12696,N_15285);
or U20485 (N_20485,N_16388,N_13164);
nand U20486 (N_20486,N_16298,N_12693);
and U20487 (N_20487,N_17411,N_12649);
or U20488 (N_20488,N_14411,N_14233);
or U20489 (N_20489,N_16179,N_15521);
or U20490 (N_20490,N_12522,N_16795);
nand U20491 (N_20491,N_14085,N_15217);
xnor U20492 (N_20492,N_16524,N_18664);
xor U20493 (N_20493,N_18021,N_13711);
nor U20494 (N_20494,N_18395,N_14903);
nor U20495 (N_20495,N_18520,N_13103);
nor U20496 (N_20496,N_14666,N_16667);
or U20497 (N_20497,N_16816,N_13732);
or U20498 (N_20498,N_16483,N_14759);
nor U20499 (N_20499,N_13869,N_15757);
and U20500 (N_20500,N_13806,N_18538);
or U20501 (N_20501,N_15942,N_18054);
nor U20502 (N_20502,N_14976,N_15838);
nor U20503 (N_20503,N_12671,N_15231);
xor U20504 (N_20504,N_18539,N_16884);
xor U20505 (N_20505,N_14947,N_18669);
or U20506 (N_20506,N_17778,N_16920);
nor U20507 (N_20507,N_15140,N_14536);
xnor U20508 (N_20508,N_18024,N_18523);
and U20509 (N_20509,N_18688,N_18026);
xnor U20510 (N_20510,N_14245,N_16993);
and U20511 (N_20511,N_17012,N_16644);
nor U20512 (N_20512,N_14672,N_18342);
and U20513 (N_20513,N_14344,N_16032);
nor U20514 (N_20514,N_18508,N_16942);
nand U20515 (N_20515,N_17109,N_13210);
nor U20516 (N_20516,N_15639,N_18408);
or U20517 (N_20517,N_15008,N_14282);
nand U20518 (N_20518,N_14690,N_15493);
nor U20519 (N_20519,N_15737,N_16331);
nand U20520 (N_20520,N_18574,N_17277);
xor U20521 (N_20521,N_14055,N_14189);
nor U20522 (N_20522,N_15692,N_14262);
or U20523 (N_20523,N_16826,N_16138);
and U20524 (N_20524,N_16854,N_16842);
nor U20525 (N_20525,N_17643,N_17131);
and U20526 (N_20526,N_13336,N_13023);
xor U20527 (N_20527,N_17275,N_13848);
nor U20528 (N_20528,N_15578,N_13808);
or U20529 (N_20529,N_15014,N_12786);
nand U20530 (N_20530,N_12776,N_12527);
or U20531 (N_20531,N_17987,N_15577);
nand U20532 (N_20532,N_13246,N_14821);
nor U20533 (N_20533,N_17133,N_13255);
nand U20534 (N_20534,N_13918,N_14529);
or U20535 (N_20535,N_15342,N_18435);
nand U20536 (N_20536,N_18334,N_13294);
xnor U20537 (N_20537,N_17734,N_17944);
nand U20538 (N_20538,N_17727,N_16542);
nor U20539 (N_20539,N_18083,N_12855);
or U20540 (N_20540,N_15612,N_17376);
nor U20541 (N_20541,N_18701,N_17594);
and U20542 (N_20542,N_17157,N_16822);
nand U20543 (N_20543,N_16033,N_17894);
nand U20544 (N_20544,N_15412,N_16708);
and U20545 (N_20545,N_13326,N_13192);
or U20546 (N_20546,N_15945,N_17593);
nand U20547 (N_20547,N_15424,N_14686);
xor U20548 (N_20548,N_17439,N_14234);
xor U20549 (N_20549,N_15745,N_16145);
or U20550 (N_20550,N_14033,N_14482);
xor U20551 (N_20551,N_15130,N_16819);
and U20552 (N_20552,N_15245,N_16328);
and U20553 (N_20553,N_13332,N_16264);
nand U20554 (N_20554,N_17689,N_16384);
nand U20555 (N_20555,N_13087,N_14296);
nor U20556 (N_20556,N_16778,N_17292);
and U20557 (N_20557,N_18085,N_17841);
or U20558 (N_20558,N_17413,N_17069);
and U20559 (N_20559,N_15102,N_15383);
or U20560 (N_20560,N_13244,N_15121);
nand U20561 (N_20561,N_14799,N_15444);
nor U20562 (N_20562,N_15139,N_13128);
nor U20563 (N_20563,N_17036,N_16814);
or U20564 (N_20564,N_17301,N_18690);
nand U20565 (N_20565,N_13340,N_13650);
nand U20566 (N_20566,N_16989,N_16181);
nor U20567 (N_20567,N_17106,N_13150);
or U20568 (N_20568,N_13899,N_15326);
nor U20569 (N_20569,N_14223,N_16463);
or U20570 (N_20570,N_14825,N_18282);
and U20571 (N_20571,N_17809,N_15604);
or U20572 (N_20572,N_17714,N_12814);
or U20573 (N_20573,N_12660,N_16294);
and U20574 (N_20574,N_13862,N_16877);
nand U20575 (N_20575,N_17791,N_17130);
nand U20576 (N_20576,N_18307,N_12592);
xor U20577 (N_20577,N_13166,N_13719);
nand U20578 (N_20578,N_14563,N_18652);
nand U20579 (N_20579,N_13606,N_18707);
nor U20580 (N_20580,N_12516,N_16339);
or U20581 (N_20581,N_15553,N_17055);
nor U20582 (N_20582,N_16647,N_14944);
nand U20583 (N_20583,N_18205,N_15230);
nand U20584 (N_20584,N_18364,N_15438);
xnor U20585 (N_20585,N_14916,N_18351);
xnor U20586 (N_20586,N_18353,N_13214);
or U20587 (N_20587,N_17054,N_14140);
and U20588 (N_20588,N_14378,N_12823);
nand U20589 (N_20589,N_16817,N_13529);
nor U20590 (N_20590,N_16183,N_16956);
or U20591 (N_20591,N_13167,N_14973);
nand U20592 (N_20592,N_17478,N_17432);
and U20593 (N_20593,N_17053,N_16712);
and U20594 (N_20594,N_13673,N_16005);
nand U20595 (N_20595,N_13404,N_16625);
nand U20596 (N_20596,N_12648,N_13694);
and U20597 (N_20597,N_12968,N_14117);
or U20598 (N_20598,N_18320,N_15839);
nor U20599 (N_20599,N_15354,N_13289);
nor U20600 (N_20600,N_17772,N_14644);
and U20601 (N_20601,N_12850,N_15043);
or U20602 (N_20602,N_13421,N_16663);
xnor U20603 (N_20603,N_18684,N_15340);
nor U20604 (N_20604,N_14210,N_16631);
nor U20605 (N_20605,N_18667,N_18361);
or U20606 (N_20606,N_12778,N_13849);
or U20607 (N_20607,N_14341,N_17798);
xnor U20608 (N_20608,N_16967,N_17649);
nor U20609 (N_20609,N_18331,N_12948);
nor U20610 (N_20610,N_17496,N_17039);
xnor U20611 (N_20611,N_15197,N_14455);
nor U20612 (N_20612,N_16639,N_13518);
nand U20613 (N_20613,N_18591,N_18746);
xor U20614 (N_20614,N_14382,N_12534);
nor U20615 (N_20615,N_14066,N_17763);
and U20616 (N_20616,N_17325,N_15564);
xnor U20617 (N_20617,N_16198,N_13258);
xor U20618 (N_20618,N_15984,N_17201);
and U20619 (N_20619,N_17837,N_16102);
xnor U20620 (N_20620,N_13232,N_12727);
or U20621 (N_20621,N_13736,N_16414);
nor U20622 (N_20622,N_14148,N_14747);
and U20623 (N_20623,N_14600,N_17771);
nand U20624 (N_20624,N_14775,N_16678);
xnor U20625 (N_20625,N_17625,N_16275);
xnor U20626 (N_20626,N_18517,N_16697);
nand U20627 (N_20627,N_14043,N_13617);
nand U20628 (N_20628,N_12509,N_17824);
or U20629 (N_20629,N_13783,N_18313);
or U20630 (N_20630,N_13048,N_13788);
nor U20631 (N_20631,N_15559,N_16823);
nor U20632 (N_20632,N_14421,N_14467);
nand U20633 (N_20633,N_14256,N_14743);
nand U20634 (N_20634,N_17926,N_12923);
nand U20635 (N_20635,N_18515,N_15208);
or U20636 (N_20636,N_12746,N_17021);
nor U20637 (N_20637,N_14864,N_18368);
and U20638 (N_20638,N_12919,N_17136);
or U20639 (N_20639,N_15376,N_15239);
nor U20640 (N_20640,N_15866,N_15429);
nor U20641 (N_20641,N_16319,N_13942);
or U20642 (N_20642,N_17119,N_13558);
xor U20643 (N_20643,N_15743,N_16653);
or U20644 (N_20644,N_17835,N_17619);
nor U20645 (N_20645,N_17504,N_15068);
nor U20646 (N_20646,N_15822,N_18211);
nor U20647 (N_20647,N_16757,N_16910);
nor U20648 (N_20648,N_16767,N_17284);
or U20649 (N_20649,N_14965,N_16601);
nor U20650 (N_20650,N_15628,N_16450);
nand U20651 (N_20651,N_14498,N_12867);
nand U20652 (N_20652,N_16564,N_13471);
or U20653 (N_20653,N_14540,N_17856);
nand U20654 (N_20654,N_12998,N_17629);
xnor U20655 (N_20655,N_13304,N_17417);
xor U20656 (N_20656,N_18135,N_18519);
nand U20657 (N_20657,N_16832,N_15328);
nor U20658 (N_20658,N_15632,N_13635);
nand U20659 (N_20659,N_14815,N_13932);
nand U20660 (N_20660,N_16288,N_16425);
xnor U20661 (N_20661,N_18433,N_18136);
nand U20662 (N_20662,N_13933,N_13789);
and U20663 (N_20663,N_14392,N_17480);
or U20664 (N_20664,N_14819,N_16958);
or U20665 (N_20665,N_13124,N_13239);
or U20666 (N_20666,N_15470,N_14522);
nand U20667 (N_20667,N_17502,N_16602);
and U20668 (N_20668,N_16502,N_18008);
nand U20669 (N_20669,N_18480,N_18333);
and U20670 (N_20670,N_14537,N_14791);
nand U20671 (N_20671,N_12554,N_13951);
xor U20672 (N_20672,N_18586,N_17562);
nor U20673 (N_20673,N_13409,N_15111);
nor U20674 (N_20674,N_15717,N_18378);
xnor U20675 (N_20675,N_12937,N_14604);
or U20676 (N_20676,N_13286,N_15273);
xnor U20677 (N_20677,N_12904,N_18033);
xnor U20678 (N_20678,N_14515,N_16168);
nand U20679 (N_20679,N_17257,N_15889);
nor U20680 (N_20680,N_15475,N_13190);
xnor U20681 (N_20681,N_17751,N_13420);
and U20682 (N_20682,N_13184,N_13791);
or U20683 (N_20683,N_14083,N_15606);
nor U20684 (N_20684,N_17454,N_18208);
nor U20685 (N_20685,N_14511,N_13106);
xor U20686 (N_20686,N_14581,N_15427);
or U20687 (N_20687,N_17924,N_18292);
nand U20688 (N_20688,N_16533,N_13129);
and U20689 (N_20689,N_16024,N_13359);
nor U20690 (N_20690,N_16775,N_12711);
and U20691 (N_20691,N_15815,N_17695);
and U20692 (N_20692,N_13796,N_17047);
or U20693 (N_20693,N_14996,N_13312);
or U20694 (N_20694,N_16746,N_18427);
nand U20695 (N_20695,N_18093,N_12947);
nand U20696 (N_20696,N_16878,N_16353);
xor U20697 (N_20697,N_13209,N_15587);
and U20698 (N_20698,N_15530,N_13569);
and U20699 (N_20699,N_17266,N_14950);
nor U20700 (N_20700,N_17128,N_16758);
nor U20701 (N_20701,N_17846,N_16233);
xnor U20702 (N_20702,N_14798,N_17208);
or U20703 (N_20703,N_18643,N_14339);
nor U20704 (N_20704,N_18073,N_17219);
and U20705 (N_20705,N_14518,N_14115);
and U20706 (N_20706,N_16030,N_15005);
nor U20707 (N_20707,N_17242,N_14255);
and U20708 (N_20708,N_14510,N_12774);
nand U20709 (N_20709,N_13838,N_13991);
nand U20710 (N_20710,N_15187,N_16464);
and U20711 (N_20711,N_13920,N_14879);
or U20712 (N_20712,N_17980,N_13878);
and U20713 (N_20713,N_15688,N_17634);
nand U20714 (N_20714,N_16123,N_15658);
nor U20715 (N_20715,N_16997,N_15085);
xnor U20716 (N_20716,N_16471,N_13252);
or U20717 (N_20717,N_17899,N_17472);
nand U20718 (N_20718,N_14528,N_12894);
nor U20719 (N_20719,N_15125,N_14888);
nand U20720 (N_20720,N_13248,N_16983);
or U20721 (N_20721,N_17739,N_18580);
or U20722 (N_20722,N_16266,N_18454);
or U20723 (N_20723,N_14380,N_18569);
xnor U20724 (N_20724,N_14355,N_15858);
and U20725 (N_20725,N_13682,N_13115);
nor U20726 (N_20726,N_16538,N_18377);
and U20727 (N_20727,N_16561,N_17260);
or U20728 (N_20728,N_14978,N_12820);
and U20729 (N_20729,N_18606,N_17832);
nand U20730 (N_20730,N_13102,N_17541);
or U20731 (N_20731,N_17135,N_15761);
nand U20732 (N_20732,N_18425,N_14076);
nand U20733 (N_20733,N_13316,N_13554);
nor U20734 (N_20734,N_13659,N_16965);
xnor U20735 (N_20735,N_13904,N_18350);
xor U20736 (N_20736,N_15597,N_13098);
or U20737 (N_20737,N_18335,N_15203);
nor U20738 (N_20738,N_14660,N_15595);
xnor U20739 (N_20739,N_12576,N_17037);
or U20740 (N_20740,N_17942,N_16759);
nand U20741 (N_20741,N_16235,N_16925);
xor U20742 (N_20742,N_13741,N_16509);
nand U20743 (N_20743,N_16302,N_15338);
xnor U20744 (N_20744,N_13756,N_18721);
and U20745 (N_20745,N_14084,N_16323);
nand U20746 (N_20746,N_18133,N_18728);
nor U20747 (N_20747,N_13735,N_15799);
nand U20748 (N_20748,N_17699,N_14401);
or U20749 (N_20749,N_13040,N_14435);
nor U20750 (N_20750,N_12620,N_16781);
nand U20751 (N_20751,N_13201,N_14458);
and U20752 (N_20752,N_13020,N_17974);
nor U20753 (N_20753,N_16271,N_15403);
and U20754 (N_20754,N_17958,N_14192);
and U20755 (N_20755,N_13822,N_15464);
or U20756 (N_20756,N_12631,N_17992);
and U20757 (N_20757,N_13056,N_17509);
nor U20758 (N_20758,N_17400,N_14701);
xor U20759 (N_20759,N_13274,N_15479);
or U20760 (N_20760,N_15709,N_17548);
or U20761 (N_20761,N_15517,N_15487);
nand U20762 (N_20762,N_15421,N_15720);
xnor U20763 (N_20763,N_18507,N_18678);
xnor U20764 (N_20764,N_16733,N_16595);
or U20765 (N_20765,N_14741,N_17115);
nand U20766 (N_20766,N_15450,N_12650);
xnor U20767 (N_20767,N_18370,N_15170);
nand U20768 (N_20768,N_15978,N_14991);
or U20769 (N_20769,N_12825,N_12917);
nor U20770 (N_20770,N_16525,N_14449);
nand U20771 (N_20771,N_13988,N_13468);
xor U20772 (N_20772,N_15323,N_15425);
and U20773 (N_20773,N_13080,N_17638);
nor U20774 (N_20774,N_15509,N_13259);
nor U20775 (N_20775,N_16472,N_18315);
xnor U20776 (N_20776,N_12957,N_12580);
xnor U20777 (N_20777,N_16971,N_14872);
xnor U20778 (N_20778,N_13686,N_15168);
or U20779 (N_20779,N_18601,N_14848);
xnor U20780 (N_20780,N_17901,N_17690);
nand U20781 (N_20781,N_17166,N_17993);
xnor U20782 (N_20782,N_17111,N_14505);
nor U20783 (N_20783,N_12939,N_14298);
or U20784 (N_20784,N_18178,N_16008);
and U20785 (N_20785,N_14389,N_15844);
and U20786 (N_20786,N_16106,N_16566);
and U20787 (N_20787,N_15608,N_17933);
xnor U20788 (N_20788,N_18284,N_12943);
nor U20789 (N_20789,N_18324,N_12858);
xnor U20790 (N_20790,N_16532,N_15531);
nand U20791 (N_20791,N_17539,N_12902);
and U20792 (N_20792,N_18414,N_17600);
and U20793 (N_20793,N_13985,N_12846);
and U20794 (N_20794,N_16186,N_16035);
nor U20795 (N_20795,N_16621,N_16650);
or U20796 (N_20796,N_13871,N_17167);
xor U20797 (N_20797,N_14006,N_15034);
nand U20798 (N_20798,N_18015,N_15523);
xnor U20799 (N_20799,N_15662,N_12960);
xnor U20800 (N_20800,N_17536,N_15908);
or U20801 (N_20801,N_15684,N_17752);
xor U20802 (N_20802,N_18421,N_18010);
and U20803 (N_20803,N_17902,N_17576);
xnor U20804 (N_20804,N_17351,N_12775);
and U20805 (N_20805,N_14306,N_15854);
xnor U20806 (N_20806,N_17609,N_17020);
and U20807 (N_20807,N_18724,N_16665);
nand U20808 (N_20808,N_13687,N_18002);
nand U20809 (N_20809,N_14605,N_14780);
xor U20810 (N_20810,N_13970,N_17834);
nor U20811 (N_20811,N_18662,N_17027);
nand U20812 (N_20812,N_15934,N_14015);
and U20813 (N_20813,N_17597,N_12550);
or U20814 (N_20814,N_14796,N_12965);
or U20815 (N_20815,N_18745,N_16061);
and U20816 (N_20816,N_16563,N_12624);
or U20817 (N_20817,N_18481,N_17004);
nand U20818 (N_20818,N_12713,N_14195);
and U20819 (N_20819,N_13481,N_14561);
nand U20820 (N_20820,N_16580,N_18641);
xnor U20821 (N_20821,N_15746,N_17227);
and U20822 (N_20822,N_13011,N_14133);
nand U20823 (N_20823,N_18486,N_15812);
nor U20824 (N_20824,N_18496,N_17421);
nor U20825 (N_20825,N_17139,N_17582);
or U20826 (N_20826,N_16980,N_14207);
or U20827 (N_20827,N_17802,N_17108);
nand U20828 (N_20828,N_17711,N_12521);
or U20829 (N_20829,N_18622,N_16142);
nand U20830 (N_20830,N_13935,N_14376);
nor U20831 (N_20831,N_18125,N_15675);
xor U20832 (N_20832,N_15512,N_13543);
and U20833 (N_20833,N_15019,N_14322);
nand U20834 (N_20834,N_12559,N_14065);
xnor U20835 (N_20835,N_13717,N_13854);
nor U20836 (N_20836,N_18168,N_13387);
xnor U20837 (N_20837,N_13362,N_12709);
or U20838 (N_20838,N_17244,N_16446);
or U20839 (N_20839,N_12983,N_17936);
nor U20840 (N_20840,N_15971,N_17876);
and U20841 (N_20841,N_15457,N_15152);
or U20842 (N_20842,N_14183,N_15569);
or U20843 (N_20843,N_16808,N_16352);
nor U20844 (N_20844,N_13516,N_17148);
xnor U20845 (N_20845,N_13119,N_14722);
or U20846 (N_20846,N_14508,N_15390);
xor U20847 (N_20847,N_13830,N_14889);
nor U20848 (N_20848,N_18541,N_12901);
nor U20849 (N_20849,N_13024,N_18560);
and U20850 (N_20850,N_15826,N_14647);
nand U20851 (N_20851,N_15997,N_18271);
and U20852 (N_20852,N_15621,N_13534);
nor U20853 (N_20853,N_14078,N_18372);
and U20854 (N_20854,N_13868,N_15432);
xor U20855 (N_20855,N_15835,N_18102);
nand U20856 (N_20856,N_16283,N_18259);
and U20857 (N_20857,N_18551,N_14097);
or U20858 (N_20858,N_18380,N_18124);
or U20859 (N_20859,N_14119,N_13462);
xnor U20860 (N_20860,N_13182,N_13396);
or U20861 (N_20861,N_13148,N_18128);
nor U20862 (N_20862,N_15339,N_17370);
nand U20863 (N_20863,N_14003,N_12732);
nand U20864 (N_20864,N_15600,N_14573);
nor U20865 (N_20865,N_18555,N_16167);
and U20866 (N_20866,N_13491,N_18236);
nand U20867 (N_20867,N_16415,N_18411);
xor U20868 (N_20868,N_15727,N_12636);
nand U20869 (N_20869,N_18308,N_14081);
and U20870 (N_20870,N_14891,N_13078);
and U20871 (N_20871,N_16652,N_13013);
and U20872 (N_20872,N_15950,N_18153);
and U20873 (N_20873,N_17161,N_17545);
and U20874 (N_20874,N_14650,N_14651);
or U20875 (N_20875,N_14016,N_16002);
and U20876 (N_20876,N_15516,N_14652);
nor U20877 (N_20877,N_14181,N_14691);
nand U20878 (N_20878,N_15574,N_14981);
nor U20879 (N_20879,N_16589,N_14428);
or U20880 (N_20880,N_18280,N_17282);
or U20881 (N_20881,N_13910,N_16627);
and U20882 (N_20882,N_17045,N_12748);
nand U20883 (N_20883,N_17023,N_14622);
xor U20884 (N_20884,N_16536,N_17181);
or U20885 (N_20885,N_16750,N_17710);
xnor U20886 (N_20886,N_13521,N_13837);
nand U20887 (N_20887,N_15165,N_15760);
xor U20888 (N_20888,N_17058,N_17538);
nor U20889 (N_20889,N_12603,N_14156);
nand U20890 (N_20890,N_16737,N_17217);
and U20891 (N_20891,N_18163,N_16076);
nand U20892 (N_20892,N_14445,N_14767);
or U20893 (N_20893,N_13203,N_13977);
or U20894 (N_20894,N_15290,N_15566);
nor U20895 (N_20895,N_17367,N_12520);
nor U20896 (N_20896,N_12970,N_15003);
nand U20897 (N_20897,N_15119,N_13666);
or U20898 (N_20898,N_13663,N_16274);
nor U20899 (N_20899,N_13608,N_17225);
or U20900 (N_20900,N_17986,N_18346);
nand U20901 (N_20901,N_12781,N_14897);
xor U20902 (N_20902,N_13916,N_15755);
xnor U20903 (N_20903,N_16393,N_14869);
and U20904 (N_20904,N_12504,N_17851);
nor U20905 (N_20905,N_18349,N_13275);
and U20906 (N_20906,N_18027,N_12863);
nor U20907 (N_20907,N_18637,N_13337);
nand U20908 (N_20908,N_13839,N_17712);
nand U20909 (N_20909,N_15243,N_13919);
and U20910 (N_20910,N_15018,N_14999);
xnor U20911 (N_20911,N_13702,N_18412);
nand U20912 (N_20912,N_16966,N_15811);
or U20913 (N_20913,N_15557,N_13482);
nor U20914 (N_20914,N_17186,N_18200);
nand U20915 (N_20915,N_17531,N_16785);
or U20916 (N_20916,N_15251,N_12507);
and U20917 (N_20917,N_17723,N_13720);
xor U20918 (N_20918,N_15169,N_16121);
and U20919 (N_20919,N_16162,N_15142);
or U20920 (N_20920,N_14325,N_15206);
and U20921 (N_20921,N_16392,N_14138);
or U20922 (N_20922,N_13153,N_12551);
nand U20923 (N_20923,N_13943,N_18392);
or U20924 (N_20924,N_18700,N_15906);
or U20925 (N_20925,N_18738,N_17793);
or U20926 (N_20926,N_17935,N_17583);
xnor U20927 (N_20927,N_17283,N_13775);
and U20928 (N_20928,N_15919,N_14632);
nand U20929 (N_20929,N_16787,N_18066);
nand U20930 (N_20930,N_12739,N_15368);
or U20931 (N_20931,N_16927,N_12925);
or U20932 (N_20932,N_15921,N_13293);
nand U20933 (N_20933,N_13071,N_17072);
and U20934 (N_20934,N_13574,N_18448);
or U20935 (N_20935,N_13329,N_16559);
and U20936 (N_20936,N_13579,N_16239);
and U20937 (N_20937,N_15900,N_17234);
nand U20938 (N_20938,N_14032,N_13814);
xnor U20939 (N_20939,N_16537,N_17456);
xor U20940 (N_20940,N_15715,N_14899);
and U20941 (N_20941,N_17382,N_14731);
or U20942 (N_20942,N_18713,N_12604);
nand U20943 (N_20943,N_13827,N_13762);
nor U20944 (N_20944,N_18465,N_18423);
nand U20945 (N_20945,N_18359,N_16325);
xor U20946 (N_20946,N_13772,N_17132);
or U20947 (N_20947,N_18204,N_16736);
and U20948 (N_20948,N_16914,N_14648);
and U20949 (N_20949,N_14415,N_14649);
nor U20950 (N_20950,N_12900,N_13619);
nor U20951 (N_20951,N_12761,N_13680);
or U20952 (N_20952,N_13466,N_14178);
and U20953 (N_20953,N_17028,N_15391);
and U20954 (N_20954,N_14585,N_15660);
nor U20955 (N_20955,N_12526,N_12857);
or U20956 (N_20956,N_15911,N_18216);
and U20957 (N_20957,N_15356,N_12661);
xnor U20958 (N_20958,N_12601,N_14383);
or U20959 (N_20959,N_16879,N_14855);
nor U20960 (N_20960,N_17120,N_18404);
nand U20961 (N_20961,N_14556,N_15856);
xnor U20962 (N_20962,N_15379,N_17062);
and U20963 (N_20963,N_15522,N_16753);
nand U20964 (N_20964,N_17127,N_13295);
xor U20965 (N_20965,N_16560,N_16645);
or U20966 (N_20966,N_14252,N_15238);
or U20967 (N_20967,N_17392,N_13177);
xor U20968 (N_20968,N_16858,N_13618);
nand U20969 (N_20969,N_14956,N_15782);
nor U20970 (N_20970,N_13507,N_18382);
and U20971 (N_20971,N_13881,N_13176);
or U20972 (N_20972,N_15620,N_13716);
nand U20973 (N_20973,N_13968,N_13230);
and U20974 (N_20974,N_14375,N_17469);
nor U20975 (N_20975,N_17513,N_14061);
or U20976 (N_20976,N_17592,N_15674);
and U20977 (N_20977,N_17398,N_18460);
nand U20978 (N_20978,N_12662,N_18457);
nor U20979 (N_20979,N_15430,N_17607);
or U20980 (N_20980,N_15501,N_17073);
xnor U20981 (N_20981,N_14103,N_14871);
and U20982 (N_20982,N_16129,N_16935);
and U20983 (N_20983,N_16205,N_14566);
and U20984 (N_20984,N_13553,N_15560);
xor U20985 (N_20985,N_15591,N_16944);
and U20986 (N_20986,N_14141,N_15933);
nand U20987 (N_20987,N_16091,N_15229);
and U20988 (N_20988,N_12819,N_17812);
nor U20989 (N_20989,N_16470,N_18294);
or U20990 (N_20990,N_17765,N_17915);
and U20991 (N_20991,N_18036,N_15174);
or U20992 (N_20992,N_15579,N_17404);
xnor U20993 (N_20993,N_15994,N_15540);
nand U20994 (N_20994,N_14712,N_16859);
and U20995 (N_20995,N_14232,N_13282);
xnor U20996 (N_20996,N_17622,N_15272);
xnor U20997 (N_20997,N_16550,N_18581);
xor U20998 (N_20998,N_13146,N_13654);
nor U20999 (N_20999,N_14242,N_15097);
or U21000 (N_21000,N_17877,N_13631);
nor U21001 (N_21001,N_18272,N_14436);
or U21002 (N_21002,N_18559,N_15673);
nor U21003 (N_21003,N_14393,N_17483);
nand U21004 (N_21004,N_16777,N_13027);
and U21005 (N_21005,N_13861,N_18557);
xnor U21006 (N_21006,N_16770,N_13955);
nand U21007 (N_21007,N_14668,N_15194);
nand U21008 (N_21008,N_17090,N_16779);
xor U21009 (N_21009,N_17267,N_18191);
xor U21010 (N_21010,N_17299,N_17467);
nand U21011 (N_21011,N_15975,N_14689);
or U21012 (N_21012,N_15040,N_12668);
or U21013 (N_21013,N_18635,N_13120);
nand U21014 (N_21014,N_17048,N_13090);
and U21015 (N_21015,N_15282,N_14261);
or U21016 (N_21016,N_15348,N_13625);
or U21017 (N_21017,N_14752,N_15293);
and U21018 (N_21018,N_17542,N_18681);
xor U21019 (N_21019,N_14168,N_15176);
or U21020 (N_21020,N_16133,N_14268);
or U21021 (N_21021,N_16869,N_13514);
nor U21022 (N_21022,N_14984,N_17474);
nand U21023 (N_21023,N_16021,N_13931);
nor U21024 (N_21024,N_13856,N_13781);
nor U21025 (N_21025,N_14674,N_17173);
xor U21026 (N_21026,N_15941,N_18053);
nor U21027 (N_21027,N_15903,N_17693);
nand U21028 (N_21028,N_15733,N_13189);
nor U21029 (N_21029,N_13689,N_14687);
nor U21030 (N_21030,N_17530,N_15872);
and U21031 (N_21031,N_18698,N_16556);
or U21032 (N_21032,N_16368,N_14676);
xor U21033 (N_21033,N_13614,N_14788);
or U21034 (N_21034,N_17098,N_14251);
or U21035 (N_21035,N_15652,N_17644);
or U21036 (N_21036,N_13874,N_14311);
and U21037 (N_21037,N_16418,N_18666);
and U21038 (N_21038,N_17387,N_15211);
or U21039 (N_21039,N_15002,N_15236);
nand U21040 (N_21040,N_17635,N_15428);
and U21041 (N_21041,N_12539,N_15695);
xor U21042 (N_21042,N_17447,N_18399);
and U21043 (N_21043,N_12769,N_15948);
nor U21044 (N_21044,N_14818,N_16254);
and U21045 (N_21045,N_12975,N_14868);
xnor U21046 (N_21046,N_15053,N_15131);
nand U21047 (N_21047,N_15762,N_14122);
or U21048 (N_21048,N_15257,N_17024);
xnor U21049 (N_21049,N_18547,N_13706);
nand U21050 (N_21050,N_15278,N_14215);
xnor U21051 (N_21051,N_15946,N_17519);
or U21052 (N_21052,N_14961,N_13066);
or U21053 (N_21053,N_15999,N_15859);
nor U21054 (N_21054,N_18590,N_18456);
or U21055 (N_21055,N_18573,N_18137);
nor U21056 (N_21056,N_13563,N_14205);
nor U21057 (N_21057,N_17358,N_12949);
nand U21058 (N_21058,N_14852,N_17269);
and U21059 (N_21059,N_17343,N_15495);
and U21060 (N_21060,N_17003,N_18527);
nand U21061 (N_21061,N_13257,N_15657);
and U21062 (N_21062,N_17630,N_13269);
or U21063 (N_21063,N_18011,N_17715);
nand U21064 (N_21064,N_12996,N_17891);
nand U21065 (N_21065,N_14206,N_13180);
nor U21066 (N_21066,N_17384,N_13894);
nand U21067 (N_21067,N_14521,N_12590);
nand U21068 (N_21068,N_17391,N_14870);
nand U21069 (N_21069,N_14716,N_14332);
and U21070 (N_21070,N_13701,N_15120);
and U21071 (N_21071,N_15031,N_16435);
xnor U21072 (N_21072,N_18034,N_16543);
or U21073 (N_21073,N_13395,N_12956);
xnor U21074 (N_21074,N_14357,N_12747);
nor U21075 (N_21075,N_13639,N_14811);
nand U21076 (N_21076,N_16225,N_13969);
and U21077 (N_21077,N_14572,N_13964);
and U21078 (N_21078,N_12511,N_12528);
and U21079 (N_21079,N_16221,N_16659);
and U21080 (N_21080,N_14330,N_15640);
nor U21081 (N_21081,N_16199,N_13025);
or U21082 (N_21082,N_13551,N_18095);
nand U21083 (N_21083,N_15159,N_17879);
xnor U21084 (N_21084,N_16682,N_17052);
or U21085 (N_21085,N_16828,N_15834);
nor U21086 (N_21086,N_16431,N_16465);
nand U21087 (N_21087,N_16677,N_15255);
nand U21088 (N_21088,N_13923,N_17011);
nor U21089 (N_21089,N_13122,N_16075);
and U21090 (N_21090,N_13125,N_17567);
xnor U21091 (N_21091,N_12698,N_15127);
xor U21092 (N_21092,N_15302,N_15619);
nand U21093 (N_21093,N_15893,N_14684);
and U21094 (N_21094,N_12548,N_17211);
or U21095 (N_21095,N_15630,N_14366);
nor U21096 (N_21096,N_18220,N_13971);
xnor U21097 (N_21097,N_18441,N_17355);
or U21098 (N_21098,N_18729,N_15089);
nor U21099 (N_21099,N_16010,N_18222);
nor U21100 (N_21100,N_14902,N_13195);
nor U21101 (N_21101,N_13253,N_16833);
nor U21102 (N_21102,N_16516,N_18184);
and U21103 (N_21103,N_14407,N_16783);
nor U21104 (N_21104,N_14760,N_13256);
xor U21105 (N_21105,N_18529,N_13297);
xor U21106 (N_21106,N_14913,N_16799);
or U21107 (N_21107,N_16372,N_17920);
nand U21108 (N_21108,N_16192,N_17616);
nand U21109 (N_21109,N_15036,N_15716);
nor U21110 (N_21110,N_18045,N_12593);
nand U21111 (N_21111,N_13641,N_17079);
xnor U21112 (N_21112,N_13075,N_15061);
nor U21113 (N_21113,N_13400,N_17046);
xnor U21114 (N_21114,N_18375,N_14592);
nand U21115 (N_21115,N_14109,N_16355);
or U21116 (N_21116,N_13927,N_13453);
xor U21117 (N_21117,N_16634,N_18443);
and U21118 (N_21118,N_13860,N_14014);
xor U21119 (N_21119,N_14617,N_15613);
nand U21120 (N_21120,N_14746,N_13101);
nor U21121 (N_21121,N_13780,N_18410);
nor U21122 (N_21122,N_16862,N_17525);
and U21123 (N_21123,N_18323,N_18613);
and U21124 (N_21124,N_14464,N_17866);
nand U21125 (N_21125,N_13728,N_12880);
or U21126 (N_21126,N_16232,N_15117);
and U21127 (N_21127,N_16651,N_14305);
and U21128 (N_21128,N_13460,N_14131);
nand U21129 (N_21129,N_13999,N_14789);
or U21130 (N_21130,N_17294,N_14067);
xor U21131 (N_21131,N_18155,N_15590);
nor U21132 (N_21132,N_15476,N_13405);
nor U21133 (N_21133,N_17346,N_12753);
nand U21134 (N_21134,N_14533,N_16272);
and U21135 (N_21135,N_17268,N_13477);
nor U21136 (N_21136,N_13713,N_14108);
xnor U21137 (N_21137,N_17209,N_12760);
or U21138 (N_21138,N_13500,N_13944);
xnor U21139 (N_21139,N_13585,N_18173);
and U21140 (N_21140,N_12838,N_16217);
and U21141 (N_21141,N_13402,N_16530);
xor U21142 (N_21142,N_16661,N_16151);
xnor U21143 (N_21143,N_14063,N_14302);
xnor U21144 (N_21144,N_13480,N_18179);
nor U21145 (N_21145,N_13747,N_15496);
xor U21146 (N_21146,N_15384,N_13753);
and U21147 (N_21147,N_16486,N_18645);
and U21148 (N_21148,N_15199,N_16292);
nand U21149 (N_21149,N_18302,N_18198);
nor U21150 (N_21150,N_15030,N_18327);
xnor U21151 (N_21151,N_16222,N_14265);
xnor U21152 (N_21152,N_16371,N_18712);
or U21153 (N_21153,N_18477,N_13876);
and U21154 (N_21154,N_15009,N_15781);
and U21155 (N_21155,N_12831,N_15529);
or U21156 (N_21156,N_17672,N_14035);
nand U21157 (N_21157,N_17099,N_16356);
and U21158 (N_21158,N_15545,N_16456);
or U21159 (N_21159,N_13498,N_17408);
nand U21160 (N_21160,N_18237,N_18549);
nand U21161 (N_21161,N_18009,N_17287);
nor U21162 (N_21162,N_14934,N_17799);
xnor U21163 (N_21163,N_17640,N_18078);
nand U21164 (N_21164,N_16110,N_15538);
xor U21165 (N_21165,N_15343,N_12638);
nand U21166 (N_21166,N_17449,N_13886);
or U21167 (N_21167,N_15810,N_17916);
nor U21168 (N_21168,N_12594,N_15803);
and U21169 (N_21169,N_16268,N_15202);
nor U21170 (N_21170,N_12808,N_17406);
xnor U21171 (N_21171,N_18181,N_16573);
nor U21172 (N_21172,N_12572,N_16521);
nand U21173 (N_21173,N_17859,N_18714);
nand U21174 (N_21174,N_13647,N_18458);
nor U21175 (N_21175,N_12679,N_17066);
nor U21176 (N_21176,N_12952,N_12995);
nor U21177 (N_21177,N_14574,N_13714);
nand U21178 (N_21178,N_13976,N_16609);
nor U21179 (N_21179,N_17510,N_16118);
or U21180 (N_21180,N_12805,N_16680);
xnor U21181 (N_21181,N_12811,N_14694);
nor U21182 (N_21182,N_14040,N_16534);
xnor U21183 (N_21183,N_17399,N_15180);
xor U21184 (N_21184,N_17175,N_13829);
nand U21185 (N_21185,N_15754,N_17329);
nor U21186 (N_21186,N_12984,N_15505);
xor U21187 (N_21187,N_17900,N_13370);
nand U21188 (N_21188,N_12654,N_13381);
nor U21189 (N_21189,N_15185,N_18438);
xor U21190 (N_21190,N_15163,N_14876);
or U21191 (N_21191,N_17429,N_14321);
nor U21192 (N_21192,N_16025,N_17084);
nor U21193 (N_21193,N_17563,N_13254);
and U21194 (N_21194,N_18597,N_12745);
and U21195 (N_21195,N_13478,N_16315);
nor U21196 (N_21196,N_16747,N_12599);
or U21197 (N_21197,N_15308,N_13655);
nor U21198 (N_21198,N_16297,N_15958);
or U21199 (N_21199,N_16459,N_15103);
nand U21200 (N_21200,N_14318,N_14045);
nor U21201 (N_21201,N_14130,N_15625);
or U21202 (N_21202,N_14214,N_13974);
and U21203 (N_21203,N_18279,N_13327);
or U21204 (N_21204,N_12905,N_15235);
or U21205 (N_21205,N_12678,N_16307);
nand U21206 (N_21206,N_18671,N_14532);
or U21207 (N_21207,N_15015,N_18493);
and U21208 (N_21208,N_16693,N_15706);
xor U21209 (N_21209,N_12773,N_13581);
xor U21210 (N_21210,N_17094,N_13186);
nor U21211 (N_21211,N_15598,N_16057);
nor U21212 (N_21212,N_15063,N_15753);
xor U21213 (N_21213,N_15565,N_17840);
or U21214 (N_21214,N_15759,N_13145);
xnor U21215 (N_21215,N_15149,N_12881);
or U21216 (N_21216,N_17910,N_14502);
or U21217 (N_21217,N_15672,N_17353);
xnor U21218 (N_21218,N_16012,N_14783);
and U21219 (N_21219,N_17026,N_14526);
and U21220 (N_21220,N_17742,N_13660);
and U21221 (N_21221,N_13564,N_14607);
or U21222 (N_21222,N_17030,N_17044);
nand U21223 (N_21223,N_13393,N_12954);
or U21224 (N_21224,N_17843,N_14590);
and U21225 (N_21225,N_12728,N_18571);
nand U21226 (N_21226,N_14681,N_14157);
or U21227 (N_21227,N_16276,N_13439);
nand U21228 (N_21228,N_15025,N_14623);
or U21229 (N_21229,N_18524,N_13863);
nor U21230 (N_21230,N_17814,N_15704);
and U21231 (N_21231,N_18603,N_12915);
nand U21232 (N_21232,N_14786,N_15266);
xor U21233 (N_21233,N_14975,N_14838);
nand U21234 (N_21234,N_18195,N_17608);
or U21235 (N_21235,N_16892,N_14425);
and U21236 (N_21236,N_16230,N_18218);
nand U21237 (N_21237,N_18510,N_15841);
and U21238 (N_21238,N_15283,N_18130);
and U21239 (N_21239,N_17770,N_12740);
xnor U21240 (N_21240,N_16153,N_16752);
and U21241 (N_21241,N_13241,N_16476);
and U21242 (N_21242,N_17097,N_18612);
and U21243 (N_21243,N_12953,N_13302);
nand U21244 (N_21244,N_18004,N_13649);
or U21245 (N_21245,N_14777,N_18071);
and U21246 (N_21246,N_14710,N_18264);
nor U21247 (N_21247,N_17018,N_15996);
and U21248 (N_21248,N_13385,N_17340);
and U21249 (N_21249,N_12700,N_17688);
nand U21250 (N_21250,N_12836,N_17590);
or U21251 (N_21251,N_18254,N_15824);
or U21252 (N_21252,N_16600,N_18096);
nand U21253 (N_21253,N_16380,N_15927);
nand U21254 (N_21254,N_15477,N_13597);
or U21255 (N_21255,N_15794,N_12627);
nor U21256 (N_21256,N_18444,N_18705);
xor U21257 (N_21257,N_16053,N_17309);
and U21258 (N_21258,N_12815,N_15750);
nor U21259 (N_21259,N_15261,N_12950);
nor U21260 (N_21260,N_16150,N_17756);
nor U21261 (N_21261,N_17645,N_16277);
or U21262 (N_21262,N_17357,N_17495);
or U21263 (N_21263,N_16489,N_16137);
and U21264 (N_21264,N_16936,N_12519);
and U21265 (N_21265,N_18509,N_17019);
or U21266 (N_21266,N_13880,N_14390);
and U21267 (N_21267,N_18276,N_12973);
or U21268 (N_21268,N_13640,N_18109);
or U21269 (N_21269,N_14704,N_14542);
or U21270 (N_21270,N_15748,N_14071);
nor U21271 (N_21271,N_15785,N_14220);
xnor U21272 (N_21272,N_16364,N_17256);
nand U21273 (N_21273,N_13237,N_15719);
nor U21274 (N_21274,N_12743,N_16897);
xnor U21275 (N_21275,N_12871,N_14928);
and U21276 (N_21276,N_16218,N_14958);
nand U21277 (N_21277,N_14985,N_18148);
nor U21278 (N_21278,N_18322,N_18325);
or U21279 (N_21279,N_14580,N_18075);
xor U21280 (N_21280,N_12706,N_12643);
or U21281 (N_21281,N_17706,N_18607);
nand U21282 (N_21282,N_17373,N_14494);
nor U21283 (N_21283,N_18394,N_15387);
and U21284 (N_21284,N_17336,N_16780);
and U21285 (N_21285,N_13441,N_17575);
and U21286 (N_21286,N_16710,N_13069);
or U21287 (N_21287,N_17005,N_15388);
xor U21288 (N_21288,N_15252,N_14745);
and U21289 (N_21289,N_16827,N_16703);
or U21290 (N_21290,N_13956,N_12877);
or U21291 (N_21291,N_14558,N_14347);
xor U21292 (N_21292,N_18677,N_17535);
and U21293 (N_21293,N_16837,N_13199);
xor U21294 (N_21294,N_14230,N_15955);
or U21295 (N_21295,N_16690,N_13154);
nand U21296 (N_21296,N_17415,N_18260);
and U21297 (N_21297,N_12981,N_15678);
xnor U21298 (N_21298,N_12735,N_13905);
nand U21299 (N_21299,N_18401,N_12510);
nand U21300 (N_21300,N_14363,N_17063);
nand U21301 (N_21301,N_13004,N_13769);
nor U21302 (N_21302,N_14527,N_17428);
or U21303 (N_21303,N_14404,N_14153);
and U21304 (N_21304,N_14072,N_14079);
and U21305 (N_21305,N_15204,N_15494);
nor U21306 (N_21306,N_15617,N_13921);
xor U21307 (N_21307,N_13219,N_14166);
and U21308 (N_21308,N_17222,N_15526);
xor U21309 (N_21309,N_15510,N_14960);
xnor U21310 (N_21310,N_13522,N_14567);
nand U21311 (N_21311,N_18537,N_16739);
or U21312 (N_21312,N_17932,N_18270);
nor U21313 (N_21313,N_16772,N_14226);
nor U21314 (N_21314,N_12684,N_17927);
nand U21315 (N_21315,N_14120,N_14683);
and U21316 (N_21316,N_13934,N_15783);
or U21317 (N_21317,N_14846,N_15725);
and U21318 (N_21318,N_15863,N_18209);
and U21319 (N_21319,N_14927,N_15325);
and U21320 (N_21320,N_18459,N_18018);
xnor U21321 (N_21321,N_15449,N_16562);
or U21322 (N_21322,N_15708,N_14150);
xor U21323 (N_21323,N_13545,N_14446);
or U21324 (N_21324,N_13057,N_18696);
xnor U21325 (N_21325,N_14851,N_13055);
nand U21326 (N_21326,N_15643,N_13121);
xnor U21327 (N_21327,N_17498,N_14806);
nor U21328 (N_21328,N_15355,N_16938);
xnor U21329 (N_21329,N_18064,N_15681);
nand U21330 (N_21330,N_15624,N_13221);
or U21331 (N_21331,N_16154,N_16670);
xnor U21332 (N_21332,N_17261,N_16585);
nand U21333 (N_21333,N_16195,N_13898);
nand U21334 (N_21334,N_12847,N_13540);
xnor U21335 (N_21335,N_16410,N_16642);
nand U21336 (N_21336,N_14021,N_13893);
nor U21337 (N_21337,N_18043,N_12979);
or U21338 (N_21338,N_14839,N_14643);
xor U21339 (N_21339,N_15377,N_13723);
nand U21340 (N_21340,N_14952,N_15453);
and U21341 (N_21341,N_16945,N_16122);
and U21342 (N_21342,N_17271,N_13308);
nand U21343 (N_21343,N_14564,N_15394);
nor U21344 (N_21344,N_18618,N_18482);
nor U21345 (N_21345,N_16797,N_13993);
and U21346 (N_21346,N_14588,N_17785);
xor U21347 (N_21347,N_13804,N_15265);
xor U21348 (N_21348,N_16996,N_14049);
and U21349 (N_21349,N_13750,N_18306);
and U21350 (N_21350,N_13813,N_15722);
xnor U21351 (N_21351,N_16755,N_14295);
xor U21352 (N_21352,N_14724,N_13598);
nand U21353 (N_21353,N_14317,N_14782);
or U21354 (N_21354,N_15852,N_17440);
nand U21355 (N_21355,N_13882,N_13503);
or U21356 (N_21356,N_14940,N_13357);
xnor U21357 (N_21357,N_17631,N_16238);
and U21358 (N_21358,N_14266,N_18384);
xor U21359 (N_21359,N_17887,N_16872);
nor U21360 (N_21360,N_18202,N_15962);
xor U21361 (N_21361,N_16046,N_13114);
xnor U21362 (N_21362,N_15309,N_15022);
and U21363 (N_21363,N_14970,N_18298);
or U21364 (N_21364,N_14143,N_13174);
and U21365 (N_21365,N_16187,N_14667);
and U21366 (N_21366,N_14374,N_15551);
and U21367 (N_21367,N_13958,N_17105);
and U21368 (N_21368,N_15588,N_15442);
nand U21369 (N_21369,N_13109,N_14725);
nor U21370 (N_21370,N_16028,N_17537);
nor U21371 (N_21371,N_14334,N_16702);
or U21372 (N_21372,N_15160,N_18117);
xnor U21373 (N_21373,N_18023,N_13599);
xor U21374 (N_21374,N_14270,N_17102);
or U21375 (N_21375,N_18631,N_13824);
or U21376 (N_21376,N_15599,N_13099);
or U21377 (N_21377,N_16514,N_14661);
xnor U21378 (N_21378,N_13041,N_17297);
or U21379 (N_21379,N_18063,N_17461);
and U21380 (N_21380,N_17395,N_15294);
xnor U21381 (N_21381,N_18536,N_15909);
and U21382 (N_21382,N_14188,N_17961);
or U21383 (N_21383,N_15874,N_17228);
nor U21384 (N_21384,N_13940,N_16265);
xnor U21385 (N_21385,N_14543,N_17310);
and U21386 (N_21386,N_17212,N_16605);
xnor U21387 (N_21387,N_18625,N_18598);
xor U21388 (N_21388,N_15110,N_18680);
nand U21389 (N_21389,N_12685,N_13980);
xor U21390 (N_21390,N_12834,N_16978);
nor U21391 (N_21391,N_14582,N_12541);
and U21392 (N_21392,N_13191,N_15081);
xor U21393 (N_21393,N_13354,N_13712);
or U21394 (N_21394,N_13213,N_12810);
and U21395 (N_21395,N_16080,N_12536);
or U21396 (N_21396,N_16725,N_15943);
nand U21397 (N_21397,N_17647,N_15422);
and U21398 (N_21398,N_17033,N_16140);
xor U21399 (N_21399,N_15572,N_16290);
nor U21400 (N_21400,N_18145,N_13458);
and U21401 (N_21401,N_16237,N_15055);
and U21402 (N_21402,N_17223,N_13632);
nand U21403 (N_21403,N_16349,N_18584);
nor U21404 (N_21404,N_14462,N_17377);
or U21405 (N_21405,N_17553,N_16932);
xor U21406 (N_21406,N_13465,N_14052);
and U21407 (N_21407,N_17922,N_16885);
nor U21408 (N_21408,N_13900,N_14565);
and U21409 (N_21409,N_18556,N_17591);
nor U21410 (N_21410,N_17420,N_17872);
or U21411 (N_21411,N_14935,N_17022);
nand U21412 (N_21412,N_18014,N_14154);
and U21413 (N_21413,N_13928,N_16031);
nor U21414 (N_21414,N_17636,N_17648);
nor U21415 (N_21415,N_16422,N_13321);
nand U21416 (N_21416,N_16317,N_13776);
and U21417 (N_21417,N_18215,N_15610);
nor U21418 (N_21418,N_16424,N_13895);
nor U21419 (N_21419,N_18303,N_18143);
nand U21420 (N_21420,N_17226,N_16875);
nor U21421 (N_21421,N_17925,N_14669);
and U21422 (N_21422,N_15964,N_16765);
nand U21423 (N_21423,N_12544,N_14335);
nand U21424 (N_21424,N_17250,N_14703);
xnor U21425 (N_21425,N_13622,N_13925);
xnor U21426 (N_21426,N_16085,N_14216);
nand U21427 (N_21427,N_17975,N_18405);
xor U21428 (N_21428,N_17521,N_17692);
nand U21429 (N_21429,N_12595,N_13966);
nor U21430 (N_21430,N_16610,N_18311);
nor U21431 (N_21431,N_17694,N_18479);
or U21432 (N_21432,N_14409,N_15644);
xor U21433 (N_21433,N_14665,N_14625);
nand U21434 (N_21434,N_16820,N_17885);
and U21435 (N_21435,N_16861,N_13107);
or U21436 (N_21436,N_13725,N_14203);
xor U21437 (N_21437,N_17324,N_17246);
and U21438 (N_21438,N_16523,N_15683);
xnor U21439 (N_21439,N_14350,N_16194);
and U21440 (N_21440,N_16143,N_14575);
and U21441 (N_21441,N_18047,N_18463);
nor U21442 (N_21442,N_15321,N_18568);
nand U21443 (N_21443,N_17847,N_16976);
and U21444 (N_21444,N_18330,N_16672);
nor U21445 (N_21445,N_14859,N_14964);
and U21446 (N_21446,N_16857,N_13436);
and U21447 (N_21447,N_14841,N_17603);
xnor U21448 (N_21448,N_16401,N_17532);
xor U21449 (N_21449,N_16719,N_16545);
or U21450 (N_21450,N_17192,N_13474);
xnor U21451 (N_21451,N_15141,N_13052);
nor U21452 (N_21452,N_16638,N_16643);
or U21453 (N_21453,N_13587,N_16172);
and U21454 (N_21454,N_16037,N_18642);
nand U21455 (N_21455,N_12801,N_17482);
or U21456 (N_21456,N_17007,N_13994);
and U21457 (N_21457,N_14598,N_13345);
xnor U21458 (N_21458,N_13661,N_18628);
nor U21459 (N_21459,N_18165,N_12870);
nand U21460 (N_21460,N_18157,N_14431);
and U21461 (N_21461,N_13091,N_16715);
nor U21462 (N_21462,N_16527,N_18633);
xnor U21463 (N_21463,N_13440,N_13408);
or U21464 (N_21464,N_17503,N_17505);
and U21465 (N_21465,N_17895,N_16742);
nor U21466 (N_21466,N_13497,N_13196);
and U21467 (N_21467,N_13557,N_17312);
or U21468 (N_21468,N_14994,N_13037);
nor U21469 (N_21469,N_15635,N_18321);
or U21470 (N_21470,N_12613,N_12535);
or U21471 (N_21471,N_16365,N_17857);
xor U21472 (N_21472,N_18006,N_16616);
and U21473 (N_21473,N_13022,N_14645);
nor U21474 (N_21474,N_14853,N_18101);
nand U21475 (N_21475,N_12542,N_13565);
nor U21476 (N_21476,N_14469,N_12988);
nor U21477 (N_21477,N_15028,N_13885);
or U21478 (N_21478,N_13573,N_14426);
nor U21479 (N_21479,N_13144,N_16963);
or U21480 (N_21480,N_13051,N_15084);
nor U21481 (N_21481,N_17656,N_14247);
and U21482 (N_21482,N_17184,N_13202);
and U21483 (N_21483,N_18082,N_13515);
xnor U21484 (N_21484,N_12912,N_16346);
and U21485 (N_21485,N_14943,N_14379);
or U21486 (N_21486,N_15585,N_18356);
or U21487 (N_21487,N_15931,N_17497);
nor U21488 (N_21488,N_14908,N_16571);
or U21489 (N_21489,N_14931,N_15533);
and U21490 (N_21490,N_15698,N_15094);
xor U21491 (N_21491,N_13149,N_18525);
nand U21492 (N_21492,N_16116,N_16574);
nand U21493 (N_21493,N_12845,N_16088);
or U21494 (N_21494,N_15249,N_18588);
or U21495 (N_21495,N_16164,N_16369);
nand U21496 (N_21496,N_13389,N_15059);
or U21497 (N_21497,N_17965,N_15615);
or U21498 (N_21498,N_18151,N_17883);
nor U21499 (N_21499,N_14609,N_17402);
or U21500 (N_21500,N_16427,N_13348);
nor U21501 (N_21501,N_16247,N_15077);
nand U21502 (N_21502,N_13821,N_15636);
or U21503 (N_21503,N_16722,N_17713);
xor U21504 (N_21504,N_14418,N_13841);
nor U21505 (N_21505,N_15659,N_12585);
xor U21506 (N_21506,N_12796,N_12832);
xor U21507 (N_21507,N_16159,N_17143);
nor U21508 (N_21508,N_17025,N_14486);
nand U21509 (N_21509,N_15375,N_17317);
and U21510 (N_21510,N_16882,N_15133);
nand U21511 (N_21511,N_14946,N_16866);
and U21512 (N_21512,N_17205,N_17707);
and U21513 (N_21513,N_13413,N_16949);
nor U21514 (N_21514,N_16999,N_15410);
nor U21515 (N_21515,N_18146,N_17308);
nand U21516 (N_21516,N_13559,N_18487);
xnor U21517 (N_21517,N_16553,N_17517);
and U21518 (N_21518,N_12710,N_17573);
or U21519 (N_21519,N_13831,N_16801);
nand U21520 (N_21520,N_17931,N_18120);
nor U21521 (N_21521,N_16234,N_13667);
xnor U21522 (N_21522,N_16279,N_18492);
nand U21523 (N_21523,N_15337,N_17386);
xor U21524 (N_21524,N_15773,N_15603);
or U21525 (N_21525,N_15655,N_16419);
and U21526 (N_21526,N_14142,N_17527);
nand U21527 (N_21527,N_16683,N_13185);
nand U21528 (N_21528,N_13552,N_15634);
or U21529 (N_21529,N_16578,N_14658);
and U21530 (N_21530,N_13733,N_15027);
nor U21531 (N_21531,N_12910,N_15833);
or U21532 (N_21532,N_15067,N_16630);
xnor U21533 (N_21533,N_12974,N_14259);
nor U21534 (N_21534,N_14930,N_18432);
xnor U21535 (N_21535,N_18502,N_17437);
nand U21536 (N_21536,N_16629,N_16263);
xor U21537 (N_21537,N_12993,N_14029);
nand U21538 (N_21538,N_14077,N_16874);
nand U21539 (N_21539,N_13310,N_12971);
nor U21540 (N_21540,N_14221,N_18227);
nor U21541 (N_21541,N_16686,N_17156);
nor U21542 (N_21542,N_13292,N_14569);
nor U21543 (N_21543,N_16051,N_12565);
nand U21544 (N_21544,N_14823,N_18417);
or U21545 (N_21545,N_17774,N_14979);
nand U21546 (N_21546,N_14795,N_15004);
nor U21547 (N_21547,N_15314,N_13568);
and U21548 (N_21548,N_18381,N_18123);
and U21549 (N_21549,N_14309,N_15193);
nand U21550 (N_21550,N_12967,N_16120);
nand U21551 (N_21551,N_13193,N_17777);
nor U21552 (N_21552,N_14172,N_18719);
xnor U21553 (N_21553,N_17082,N_13386);
xnor U21554 (N_21554,N_16251,N_16211);
nor U21555 (N_21555,N_13050,N_17892);
and U21556 (N_21556,N_13062,N_16541);
nand U21557 (N_21557,N_16836,N_18080);
nand U21558 (N_21558,N_13888,N_13018);
nand U21559 (N_21559,N_17728,N_16048);
xnor U21560 (N_21560,N_14922,N_15830);
and U21561 (N_21561,N_14705,N_16960);
nand U21562 (N_21562,N_15700,N_15614);
nor U21563 (N_21563,N_18437,N_16156);
xnor U21564 (N_21564,N_13456,N_16336);
and U21565 (N_21565,N_14849,N_14967);
nor U21566 (N_21566,N_18518,N_13643);
and U21567 (N_21567,N_13648,N_15026);
nor U21568 (N_21568,N_17486,N_16429);
nor U21569 (N_21569,N_16873,N_18629);
and U21570 (N_21570,N_18691,N_13494);
and U21571 (N_21571,N_15396,N_15404);
and U21572 (N_21572,N_15054,N_16097);
xnor U21573 (N_21573,N_14831,N_13325);
nand U21574 (N_21574,N_14225,N_17214);
nor U21575 (N_21575,N_17452,N_17356);
xnor U21576 (N_21576,N_14351,N_17000);
nand U21577 (N_21577,N_14352,N_12553);
nor U21578 (N_21578,N_18747,N_14121);
nand U21579 (N_21579,N_18257,N_18310);
nor U21580 (N_21580,N_14630,N_18164);
and U21581 (N_21581,N_15740,N_15703);
or U21582 (N_21582,N_18639,N_12887);
and U21583 (N_21583,N_18147,N_15162);
xor U21584 (N_21584,N_12673,N_17524);
xor U21585 (N_21585,N_14208,N_17515);
nand U21586 (N_21586,N_18289,N_18365);
nand U21587 (N_21587,N_17050,N_14636);
or U21588 (N_21588,N_13768,N_13770);
and U21589 (N_21589,N_17682,N_15806);
or U21590 (N_21590,N_15216,N_18398);
xnor U21591 (N_21591,N_17043,N_18296);
xor U21592 (N_21592,N_13853,N_14373);
nor U21593 (N_21593,N_16381,N_15441);
and U21594 (N_21594,N_16065,N_17273);
nand U21595 (N_21595,N_14736,N_17270);
or U21596 (N_21596,N_17827,N_14929);
nand U21597 (N_21597,N_12640,N_16009);
nand U21598 (N_21598,N_17551,N_17534);
xnor U21599 (N_21599,N_17158,N_13194);
nor U21600 (N_21600,N_17262,N_16447);
or U21601 (N_21601,N_14018,N_15752);
or U21602 (N_21602,N_17788,N_15851);
xor U21603 (N_21603,N_15764,N_14535);
and U21604 (N_21604,N_17680,N_16236);
nand U21605 (N_21605,N_13612,N_17207);
xor U21606 (N_21606,N_15816,N_14909);
nor U21607 (N_21607,N_16727,N_17991);
nand U21608 (N_21608,N_13891,N_15793);
or U21609 (N_21609,N_13877,N_14980);
nand U21610 (N_21610,N_17220,N_16594);
xor U21611 (N_21611,N_18067,N_16006);
xor U21612 (N_21612,N_16730,N_14136);
xnor U21613 (N_21613,N_14506,N_18659);
nand U21614 (N_21614,N_15504,N_16477);
and U21615 (N_21615,N_17691,N_14031);
and U21616 (N_21616,N_16204,N_16889);
xor U21617 (N_21617,N_13580,N_13533);
or U21618 (N_21618,N_15897,N_15069);
nand U21619 (N_21619,N_17334,N_16928);
xor U21620 (N_21620,N_13645,N_17477);
nand U21621 (N_21621,N_17191,N_17316);
xor U21622 (N_21622,N_14626,N_17015);
and U21623 (N_21623,N_17683,N_12667);
nand U21624 (N_21624,N_14307,N_17716);
or U21625 (N_21625,N_15647,N_17985);
xnor U21626 (N_21626,N_17481,N_13675);
and U21627 (N_21627,N_18533,N_12714);
xor U21628 (N_21628,N_17302,N_17163);
nor U21629 (N_21629,N_13786,N_18374);
nor U21630 (N_21630,N_16870,N_16494);
nor U21631 (N_21631,N_15426,N_15848);
xnor U21632 (N_21632,N_18694,N_18725);
and U21633 (N_21633,N_14640,N_15676);
or U21634 (N_21634,N_12885,N_13662);
and U21635 (N_21635,N_18105,N_14700);
nor U21636 (N_21636,N_14729,N_14417);
nor U21637 (N_21637,N_17259,N_18422);
or U21638 (N_21638,N_14475,N_15795);
xnor U21639 (N_21639,N_15576,N_16312);
and U21640 (N_21640,N_14714,N_17144);
or U21641 (N_21641,N_15406,N_18585);
xnor U21642 (N_21642,N_15982,N_16270);
nor U21643 (N_21643,N_15694,N_12704);
nor U21644 (N_21644,N_14992,N_14599);
nand U21645 (N_21645,N_18473,N_16378);
nor U21646 (N_21646,N_16984,N_17159);
nand U21647 (N_21647,N_13536,N_13452);
or U21648 (N_21648,N_18326,N_14481);
nand U21649 (N_21649,N_15367,N_13350);
xor U21650 (N_21650,N_16593,N_16803);
xor U21651 (N_21651,N_13739,N_13922);
nand U21652 (N_21652,N_15362,N_16567);
and U21653 (N_21653,N_15914,N_13260);
and U21654 (N_21654,N_13026,N_12598);
or U21655 (N_21655,N_15259,N_15770);
or U21656 (N_21656,N_15286,N_18554);
or U21657 (N_21657,N_18139,N_16286);
xor U21658 (N_21658,N_16762,N_14514);
and U21659 (N_21659,N_15938,N_17114);
or U21660 (N_21660,N_13311,N_15109);
xor U21661 (N_21661,N_17193,N_14240);
nor U21662 (N_21662,N_18126,N_15123);
and U21663 (N_21663,N_17784,N_13187);
or U21664 (N_21664,N_18288,N_12782);
and U21665 (N_21665,N_12999,N_15520);
and U21666 (N_21666,N_13751,N_13397);
nand U21667 (N_21667,N_17819,N_18614);
nor U21668 (N_21668,N_17418,N_16394);
or U21669 (N_21669,N_15915,N_18183);
xnor U21670 (N_21670,N_17577,N_15032);
xnor U21671 (N_21671,N_16707,N_18491);
xnor U21672 (N_21672,N_18243,N_13227);
and U21673 (N_21673,N_15663,N_16479);
and U21674 (N_21674,N_13412,N_16316);
nand U21675 (N_21675,N_16170,N_14656);
nand U21676 (N_21676,N_15980,N_13285);
nor U21677 (N_21677,N_16107,N_17369);
nand U21678 (N_21678,N_13083,N_17177);
nand U21679 (N_21679,N_14367,N_13118);
nor U21680 (N_21680,N_18623,N_17093);
and U21681 (N_21681,N_17107,N_14972);
nor U21682 (N_21682,N_14474,N_18001);
xnor U21683 (N_21683,N_13033,N_18142);
nand U21684 (N_21684,N_12843,N_13132);
or U21685 (N_21685,N_17304,N_13506);
nor U21686 (N_21686,N_18732,N_12558);
or U21687 (N_21687,N_14698,N_12720);
xor U21688 (N_21688,N_16223,N_14634);
xor U21689 (N_21689,N_13288,N_15135);
xor U21690 (N_21690,N_14465,N_12913);
nand U21691 (N_21691,N_12733,N_16127);
and U21692 (N_21692,N_12557,N_15371);
nor U21693 (N_21693,N_15802,N_17057);
xnor U21694 (N_21694,N_14324,N_15365);
nand U21695 (N_21695,N_17526,N_17850);
nor U21696 (N_21696,N_17196,N_18228);
xnor U21697 (N_21697,N_12707,N_14570);
nor U21698 (N_21698,N_17528,N_16656);
nand U21699 (N_21699,N_12591,N_14720);
nand U21700 (N_21700,N_14639,N_13344);
or U21701 (N_21701,N_13151,N_18345);
nor U21702 (N_21702,N_14092,N_17448);
and U21703 (N_21703,N_15331,N_16713);
or U21704 (N_21704,N_17463,N_14901);
xor U21705 (N_21705,N_17998,N_12586);
nand U21706 (N_21706,N_17520,N_17142);
or U21707 (N_21707,N_12642,N_15451);
nor U21708 (N_21708,N_15213,N_15260);
or U21709 (N_21709,N_14512,N_16408);
and U21710 (N_21710,N_15988,N_15713);
or U21711 (N_21711,N_15023,N_16473);
xnor U21712 (N_21712,N_17934,N_16267);
and U21713 (N_21713,N_16421,N_14303);
or U21714 (N_21714,N_13475,N_13443);
and U21715 (N_21715,N_14491,N_14659);
nor U21716 (N_21716,N_15006,N_14794);
xnor U21717 (N_21717,N_18679,N_16570);
and U21718 (N_21718,N_18516,N_17436);
nand U21719 (N_21719,N_12501,N_14596);
and U21720 (N_21720,N_14041,N_18338);
and U21721 (N_21721,N_16226,N_13778);
and U21722 (N_21722,N_18038,N_15112);
xnor U21723 (N_21723,N_16895,N_18735);
nor U21724 (N_21724,N_15930,N_15227);
or U21725 (N_21725,N_15181,N_15446);
or U21726 (N_21726,N_17422,N_15738);
nand U21727 (N_21727,N_13982,N_12830);
xor U21728 (N_21728,N_13334,N_16939);
nand U21729 (N_21729,N_14360,N_16434);
or U21730 (N_21730,N_13367,N_17240);
and U21731 (N_21731,N_17687,N_15070);
xor U21732 (N_21732,N_17852,N_14912);
xnor U21733 (N_21733,N_15440,N_17006);
and U21734 (N_21734,N_16438,N_13077);
xor U21735 (N_21735,N_15253,N_13183);
nor U21736 (N_21736,N_17568,N_15060);
xnor U21737 (N_21737,N_17313,N_13843);
and U21738 (N_21738,N_14800,N_14880);
xnor U21739 (N_21739,N_18532,N_17176);
or U21740 (N_21740,N_18484,N_15079);
and U21741 (N_21741,N_14671,N_14631);
nor U21742 (N_21742,N_13997,N_16883);
nor U21743 (N_21743,N_15240,N_16856);
and U21744 (N_21744,N_13915,N_13046);
nand U21745 (N_21745,N_14277,N_16117);
or U21746 (N_21746,N_17754,N_14866);
xor U21747 (N_21747,N_13428,N_14451);
xor U21748 (N_21748,N_14406,N_18187);
nand U21749 (N_21749,N_15808,N_18290);
nor U21750 (N_21750,N_18513,N_14635);
and U21751 (N_21751,N_15862,N_13417);
nor U21752 (N_21752,N_14995,N_17665);
or U21753 (N_21753,N_18558,N_14116);
or U21754 (N_21754,N_13200,N_13541);
xor U21755 (N_21755,N_17897,N_16919);
nor U21756 (N_21756,N_15017,N_17078);
nor U21757 (N_21757,N_13473,N_13527);
nand U21758 (N_21758,N_13577,N_17659);
nand U21759 (N_21759,N_17216,N_12632);
or U21760 (N_21760,N_17549,N_17077);
nor U21761 (N_21761,N_14638,N_15739);
xnor U21762 (N_21762,N_14878,N_14111);
nand U21763 (N_21763,N_15179,N_13767);
xnor U21764 (N_21764,N_14485,N_13941);
and U21765 (N_21765,N_15489,N_14399);
nor U21766 (N_21766,N_17237,N_16613);
xnor U21767 (N_21767,N_17878,N_16649);
and U21768 (N_21768,N_16721,N_13867);
xor U21769 (N_21769,N_12694,N_18605);
and U21770 (N_21770,N_17762,N_13242);
nand U21771 (N_21771,N_17759,N_16001);
or U21772 (N_21772,N_13550,N_14271);
or U21773 (N_21773,N_12571,N_18226);
nand U21774 (N_21774,N_16968,N_18244);
and U21775 (N_21775,N_15374,N_15573);
or U21776 (N_21776,N_15413,N_17996);
nor U21777 (N_21777,N_18291,N_15335);
and U21778 (N_21778,N_14584,N_17064);
or U21779 (N_21779,N_14861,N_17736);
nand U21780 (N_21780,N_17615,N_16125);
or U21781 (N_21781,N_12816,N_14235);
nor U21782 (N_21782,N_12523,N_14734);
and U21783 (N_21783,N_15596,N_15151);
nor U21784 (N_21784,N_13699,N_15360);
nand U21785 (N_21785,N_16020,N_13205);
and U21786 (N_21786,N_15098,N_15507);
and U21787 (N_21787,N_17867,N_17587);
nand U21788 (N_21788,N_17490,N_13607);
nor U21789 (N_21789,N_18632,N_16436);
xnor U21790 (N_21790,N_15847,N_13759);
and U21791 (N_21791,N_16741,N_15721);
and U21792 (N_21792,N_17554,N_16774);
nor U21793 (N_21793,N_15827,N_16090);
nor U21794 (N_21794,N_14513,N_16252);
nand U21795 (N_21795,N_17200,N_15817);
xor U21796 (N_21796,N_14279,N_14439);
xnor U21797 (N_21797,N_13621,N_16281);
xor U21798 (N_21798,N_18035,N_12724);
nor U21799 (N_21799,N_15837,N_13578);
nand U21800 (N_21800,N_13276,N_15970);
nor U21801 (N_21801,N_16405,N_18206);
and U21802 (N_21802,N_18449,N_15821);
xor U21803 (N_21803,N_14423,N_16176);
nor U21804 (N_21804,N_16899,N_15976);
xor U21805 (N_21805,N_15200,N_15875);
nand U21806 (N_21806,N_15861,N_17442);
nand U21807 (N_21807,N_15548,N_14146);
and U21808 (N_21808,N_16342,N_14182);
xnor U21809 (N_21809,N_14932,N_14910);
and U21810 (N_21810,N_18526,N_16208);
xnor U21811 (N_21811,N_17873,N_16068);
nor U21812 (N_21812,N_13152,N_13986);
or U21813 (N_21813,N_17864,N_16333);
or U21814 (N_21814,N_15274,N_14134);
nor U21815 (N_21815,N_13990,N_16083);
xnor U21816 (N_21816,N_17281,N_14365);
or U21817 (N_21817,N_12922,N_12606);
nand U21818 (N_21818,N_13962,N_16113);
nand U21819 (N_21819,N_16943,N_15550);
nand U21820 (N_21820,N_16548,N_15977);
xnor U21821 (N_21821,N_13586,N_16495);
or U21822 (N_21822,N_13858,N_13388);
nor U21823 (N_21823,N_17359,N_12533);
and U21824 (N_21824,N_18393,N_15052);
or U21825 (N_21825,N_14987,N_14250);
nor U21826 (N_21826,N_14023,N_18081);
or U21827 (N_21827,N_13803,N_16924);
nor U21828 (N_21828,N_16411,N_16913);
nand U21829 (N_21829,N_13504,N_13028);
nand U21830 (N_21830,N_13948,N_17667);
nor U21831 (N_21831,N_16313,N_13981);
or U21832 (N_21832,N_16169,N_16022);
or U21833 (N_21833,N_17508,N_15460);
or U21834 (N_21834,N_13669,N_14500);
xnor U21835 (N_21835,N_12734,N_18017);
nand U21836 (N_21836,N_17581,N_15876);
xnor U21837 (N_21837,N_18702,N_17100);
or U21838 (N_21838,N_12540,N_18317);
nand U21839 (N_21839,N_15677,N_15076);
and U21840 (N_21840,N_16671,N_17555);
nor U21841 (N_21841,N_14211,N_14288);
and U21842 (N_21842,N_16923,N_16480);
xnor U21843 (N_21843,N_14549,N_16432);
xor U21844 (N_21844,N_12633,N_17790);
and U21845 (N_21845,N_12813,N_16399);
or U21846 (N_21846,N_12765,N_12798);
or U21847 (N_21847,N_14778,N_12659);
nor U21848 (N_21848,N_17671,N_14184);
nand U21849 (N_21849,N_18152,N_14204);
and U21850 (N_21850,N_16038,N_14968);
nand U21851 (N_21851,N_15350,N_14586);
nand U21852 (N_21852,N_13844,N_13623);
xnor U21853 (N_21853,N_13555,N_13629);
and U21854 (N_21854,N_15645,N_14885);
nor U21855 (N_21855,N_12716,N_14438);
or U21856 (N_21856,N_17140,N_13307);
nor U21857 (N_21857,N_14784,N_14336);
xor U21858 (N_21858,N_17198,N_16950);
or U21859 (N_21859,N_12931,N_15250);
xnor U21860 (N_21860,N_14364,N_14044);
or U21861 (N_21861,N_15567,N_17116);
nand U21862 (N_21862,N_14243,N_12932);
xnor U21863 (N_21863,N_17569,N_12737);
nor U21864 (N_21864,N_13810,N_14907);
and U21865 (N_21865,N_16229,N_14779);
and U21866 (N_21866,N_16067,N_18431);
xnor U21867 (N_21867,N_15046,N_16390);
nand U21868 (N_21868,N_17533,N_14391);
nor U21869 (N_21869,N_13343,N_16003);
xor U21870 (N_21870,N_14429,N_18238);
nor U21871 (N_21871,N_16344,N_16196);
xnor U21872 (N_21872,N_18020,N_16220);
xor U21873 (N_21873,N_18360,N_16101);
or U21874 (N_21874,N_18171,N_16728);
xnor U21875 (N_21875,N_18261,N_17915);
nor U21876 (N_21876,N_18575,N_16807);
nor U21877 (N_21877,N_16582,N_13026);
or U21878 (N_21878,N_16344,N_16074);
nand U21879 (N_21879,N_18538,N_14544);
xor U21880 (N_21880,N_16476,N_16863);
or U21881 (N_21881,N_14039,N_14400);
nand U21882 (N_21882,N_16642,N_13615);
or U21883 (N_21883,N_16022,N_14177);
and U21884 (N_21884,N_17303,N_15130);
and U21885 (N_21885,N_14629,N_13409);
and U21886 (N_21886,N_15891,N_17601);
nand U21887 (N_21887,N_13877,N_17000);
and U21888 (N_21888,N_17288,N_18174);
or U21889 (N_21889,N_13895,N_14632);
or U21890 (N_21890,N_15923,N_15664);
and U21891 (N_21891,N_15682,N_16937);
or U21892 (N_21892,N_12975,N_16203);
and U21893 (N_21893,N_18740,N_13945);
or U21894 (N_21894,N_14288,N_16972);
and U21895 (N_21895,N_13928,N_17832);
nor U21896 (N_21896,N_12850,N_17375);
nand U21897 (N_21897,N_17448,N_18378);
and U21898 (N_21898,N_16743,N_14996);
nor U21899 (N_21899,N_14498,N_16629);
nand U21900 (N_21900,N_16178,N_16079);
or U21901 (N_21901,N_15459,N_15119);
xnor U21902 (N_21902,N_17501,N_14980);
nand U21903 (N_21903,N_15587,N_18587);
or U21904 (N_21904,N_12551,N_13857);
nor U21905 (N_21905,N_16322,N_16091);
nor U21906 (N_21906,N_14938,N_17206);
or U21907 (N_21907,N_13129,N_16300);
or U21908 (N_21908,N_13504,N_13110);
or U21909 (N_21909,N_15594,N_15612);
and U21910 (N_21910,N_18594,N_14817);
nor U21911 (N_21911,N_14929,N_15677);
xor U21912 (N_21912,N_16469,N_16222);
and U21913 (N_21913,N_17713,N_15676);
nor U21914 (N_21914,N_15673,N_15883);
and U21915 (N_21915,N_16530,N_16111);
and U21916 (N_21916,N_12825,N_13818);
nor U21917 (N_21917,N_16537,N_18558);
and U21918 (N_21918,N_13210,N_15689);
nand U21919 (N_21919,N_14163,N_18617);
or U21920 (N_21920,N_16274,N_13589);
and U21921 (N_21921,N_13047,N_14684);
or U21922 (N_21922,N_17128,N_16305);
nor U21923 (N_21923,N_15468,N_13606);
or U21924 (N_21924,N_17848,N_16373);
nand U21925 (N_21925,N_13642,N_13205);
nand U21926 (N_21926,N_16671,N_12947);
xnor U21927 (N_21927,N_12784,N_13157);
nor U21928 (N_21928,N_14903,N_18372);
or U21929 (N_21929,N_18089,N_18700);
and U21930 (N_21930,N_15142,N_14025);
or U21931 (N_21931,N_15803,N_18263);
or U21932 (N_21932,N_15838,N_16778);
xnor U21933 (N_21933,N_13742,N_17572);
xor U21934 (N_21934,N_13251,N_17609);
or U21935 (N_21935,N_12504,N_14100);
and U21936 (N_21936,N_17048,N_12627);
nor U21937 (N_21937,N_15816,N_12650);
xnor U21938 (N_21938,N_13445,N_14335);
and U21939 (N_21939,N_13706,N_16204);
nor U21940 (N_21940,N_18022,N_14840);
xor U21941 (N_21941,N_15329,N_16052);
xnor U21942 (N_21942,N_18064,N_17225);
or U21943 (N_21943,N_18497,N_16026);
xor U21944 (N_21944,N_14391,N_12578);
nor U21945 (N_21945,N_17400,N_13933);
nand U21946 (N_21946,N_18028,N_16956);
nand U21947 (N_21947,N_17741,N_14469);
or U21948 (N_21948,N_17056,N_12738);
and U21949 (N_21949,N_13713,N_15594);
nand U21950 (N_21950,N_16369,N_15144);
and U21951 (N_21951,N_15149,N_17450);
xor U21952 (N_21952,N_14902,N_15960);
nand U21953 (N_21953,N_13261,N_17024);
nand U21954 (N_21954,N_16065,N_13523);
nor U21955 (N_21955,N_15084,N_18179);
nand U21956 (N_21956,N_15575,N_18735);
nand U21957 (N_21957,N_14495,N_16990);
and U21958 (N_21958,N_16541,N_16873);
or U21959 (N_21959,N_16104,N_17353);
xnor U21960 (N_21960,N_16545,N_16243);
nand U21961 (N_21961,N_16663,N_18025);
nor U21962 (N_21962,N_17942,N_17983);
nor U21963 (N_21963,N_16500,N_13385);
and U21964 (N_21964,N_17143,N_18282);
or U21965 (N_21965,N_12502,N_12668);
xor U21966 (N_21966,N_13316,N_18475);
and U21967 (N_21967,N_18645,N_18284);
nor U21968 (N_21968,N_13126,N_15440);
xnor U21969 (N_21969,N_18088,N_13027);
xor U21970 (N_21970,N_14338,N_16576);
nand U21971 (N_21971,N_12645,N_15150);
nor U21972 (N_21972,N_16668,N_15810);
nor U21973 (N_21973,N_15787,N_15171);
nor U21974 (N_21974,N_14875,N_17181);
xnor U21975 (N_21975,N_15667,N_15571);
and U21976 (N_21976,N_15383,N_13224);
xor U21977 (N_21977,N_12600,N_16770);
nor U21978 (N_21978,N_12873,N_15777);
nand U21979 (N_21979,N_13488,N_13678);
or U21980 (N_21980,N_12823,N_14045);
or U21981 (N_21981,N_14210,N_15006);
xnor U21982 (N_21982,N_18209,N_16163);
xor U21983 (N_21983,N_18060,N_17768);
xnor U21984 (N_21984,N_13451,N_13703);
and U21985 (N_21985,N_13306,N_14235);
nand U21986 (N_21986,N_13786,N_14920);
and U21987 (N_21987,N_14620,N_14606);
and U21988 (N_21988,N_15023,N_14604);
xor U21989 (N_21989,N_14436,N_13987);
xor U21990 (N_21990,N_14653,N_13689);
and U21991 (N_21991,N_14945,N_18348);
nor U21992 (N_21992,N_18124,N_13812);
and U21993 (N_21993,N_13160,N_17903);
or U21994 (N_21994,N_18078,N_15346);
nand U21995 (N_21995,N_16365,N_13477);
nor U21996 (N_21996,N_12533,N_16278);
and U21997 (N_21997,N_18055,N_12517);
or U21998 (N_21998,N_16005,N_17789);
or U21999 (N_21999,N_13561,N_13637);
xnor U22000 (N_22000,N_15893,N_15248);
nand U22001 (N_22001,N_13178,N_14289);
or U22002 (N_22002,N_15518,N_16659);
nor U22003 (N_22003,N_13745,N_14660);
and U22004 (N_22004,N_15807,N_18530);
xor U22005 (N_22005,N_16429,N_14204);
and U22006 (N_22006,N_12881,N_13373);
nand U22007 (N_22007,N_16015,N_14216);
nand U22008 (N_22008,N_18747,N_14186);
or U22009 (N_22009,N_17273,N_16561);
or U22010 (N_22010,N_15257,N_13312);
nand U22011 (N_22011,N_16918,N_15004);
xor U22012 (N_22012,N_12582,N_16806);
nor U22013 (N_22013,N_18664,N_15052);
or U22014 (N_22014,N_12506,N_15600);
nand U22015 (N_22015,N_16126,N_18223);
nand U22016 (N_22016,N_14316,N_16842);
nor U22017 (N_22017,N_16190,N_14265);
or U22018 (N_22018,N_15152,N_12704);
or U22019 (N_22019,N_14262,N_18210);
or U22020 (N_22020,N_15094,N_14268);
nor U22021 (N_22021,N_15455,N_18093);
xor U22022 (N_22022,N_16942,N_14501);
or U22023 (N_22023,N_16268,N_13132);
and U22024 (N_22024,N_18292,N_16966);
nor U22025 (N_22025,N_12568,N_13234);
nand U22026 (N_22026,N_14335,N_12808);
nand U22027 (N_22027,N_16559,N_15338);
or U22028 (N_22028,N_12633,N_13898);
nand U22029 (N_22029,N_13895,N_13283);
or U22030 (N_22030,N_13128,N_12751);
nor U22031 (N_22031,N_16726,N_17570);
xnor U22032 (N_22032,N_18085,N_16427);
nor U22033 (N_22033,N_18725,N_16667);
or U22034 (N_22034,N_16901,N_12557);
nor U22035 (N_22035,N_18123,N_16225);
nor U22036 (N_22036,N_15067,N_14959);
nand U22037 (N_22037,N_17054,N_14637);
or U22038 (N_22038,N_14768,N_17490);
or U22039 (N_22039,N_17088,N_17369);
nand U22040 (N_22040,N_15024,N_15459);
and U22041 (N_22041,N_15909,N_18082);
xor U22042 (N_22042,N_15928,N_17751);
and U22043 (N_22043,N_18119,N_18298);
and U22044 (N_22044,N_15663,N_17508);
or U22045 (N_22045,N_15302,N_18139);
xor U22046 (N_22046,N_16126,N_17913);
nor U22047 (N_22047,N_13070,N_16591);
and U22048 (N_22048,N_16289,N_16535);
and U22049 (N_22049,N_13103,N_17209);
xor U22050 (N_22050,N_17098,N_14491);
xor U22051 (N_22051,N_15085,N_13338);
nand U22052 (N_22052,N_12767,N_13737);
and U22053 (N_22053,N_12631,N_15999);
nor U22054 (N_22054,N_18156,N_18465);
xor U22055 (N_22055,N_13691,N_16991);
nand U22056 (N_22056,N_14816,N_15490);
and U22057 (N_22057,N_16061,N_18448);
or U22058 (N_22058,N_14565,N_13349);
xor U22059 (N_22059,N_12972,N_14794);
nor U22060 (N_22060,N_13473,N_16346);
xnor U22061 (N_22061,N_18379,N_15931);
nor U22062 (N_22062,N_12764,N_17734);
nor U22063 (N_22063,N_14232,N_12575);
nand U22064 (N_22064,N_17585,N_14770);
nor U22065 (N_22065,N_14694,N_12501);
xnor U22066 (N_22066,N_18681,N_18420);
nor U22067 (N_22067,N_17170,N_18672);
xnor U22068 (N_22068,N_14641,N_16246);
xnor U22069 (N_22069,N_16673,N_17487);
or U22070 (N_22070,N_13959,N_13038);
xnor U22071 (N_22071,N_17278,N_16222);
xor U22072 (N_22072,N_16190,N_18735);
xnor U22073 (N_22073,N_14399,N_13024);
nand U22074 (N_22074,N_14421,N_18019);
xnor U22075 (N_22075,N_17638,N_16567);
and U22076 (N_22076,N_17744,N_12855);
or U22077 (N_22077,N_17356,N_13493);
or U22078 (N_22078,N_14962,N_15927);
nand U22079 (N_22079,N_15599,N_16246);
xnor U22080 (N_22080,N_15113,N_18685);
nor U22081 (N_22081,N_17415,N_15752);
and U22082 (N_22082,N_13060,N_18023);
xnor U22083 (N_22083,N_13372,N_13125);
and U22084 (N_22084,N_13238,N_13195);
xnor U22085 (N_22085,N_17960,N_13839);
nand U22086 (N_22086,N_18452,N_14072);
nor U22087 (N_22087,N_14170,N_12755);
nand U22088 (N_22088,N_13712,N_13314);
or U22089 (N_22089,N_15140,N_13926);
or U22090 (N_22090,N_13177,N_13017);
and U22091 (N_22091,N_18116,N_15530);
xor U22092 (N_22092,N_13876,N_13812);
and U22093 (N_22093,N_12667,N_16367);
nand U22094 (N_22094,N_14281,N_14296);
and U22095 (N_22095,N_13108,N_14613);
and U22096 (N_22096,N_14298,N_18191);
nor U22097 (N_22097,N_12500,N_12657);
xor U22098 (N_22098,N_16364,N_15892);
and U22099 (N_22099,N_17139,N_18035);
nand U22100 (N_22100,N_17154,N_12891);
nor U22101 (N_22101,N_13075,N_16196);
or U22102 (N_22102,N_15496,N_17546);
or U22103 (N_22103,N_14627,N_16340);
nor U22104 (N_22104,N_13948,N_14818);
and U22105 (N_22105,N_15850,N_15694);
nor U22106 (N_22106,N_14872,N_17778);
xor U22107 (N_22107,N_15819,N_18633);
or U22108 (N_22108,N_17021,N_16475);
and U22109 (N_22109,N_18118,N_15059);
nand U22110 (N_22110,N_14485,N_14575);
or U22111 (N_22111,N_15989,N_17667);
xor U22112 (N_22112,N_13270,N_16061);
or U22113 (N_22113,N_15342,N_16809);
nand U22114 (N_22114,N_14526,N_12945);
nand U22115 (N_22115,N_15971,N_14489);
nor U22116 (N_22116,N_16383,N_14012);
nor U22117 (N_22117,N_16905,N_15978);
nor U22118 (N_22118,N_17061,N_12620);
nor U22119 (N_22119,N_14193,N_17862);
or U22120 (N_22120,N_14553,N_12604);
xnor U22121 (N_22121,N_13867,N_17972);
nand U22122 (N_22122,N_15246,N_17512);
or U22123 (N_22123,N_16531,N_13190);
xor U22124 (N_22124,N_15101,N_15948);
or U22125 (N_22125,N_12962,N_18713);
xnor U22126 (N_22126,N_15271,N_15185);
and U22127 (N_22127,N_16782,N_12620);
nor U22128 (N_22128,N_14062,N_15995);
or U22129 (N_22129,N_17459,N_17817);
or U22130 (N_22130,N_18213,N_18131);
xnor U22131 (N_22131,N_14268,N_15280);
xor U22132 (N_22132,N_12572,N_12996);
nand U22133 (N_22133,N_18482,N_15031);
nor U22134 (N_22134,N_16987,N_13019);
nor U22135 (N_22135,N_17190,N_15667);
nor U22136 (N_22136,N_17315,N_13327);
or U22137 (N_22137,N_13004,N_18460);
or U22138 (N_22138,N_16439,N_17929);
or U22139 (N_22139,N_16896,N_16009);
and U22140 (N_22140,N_16014,N_16643);
and U22141 (N_22141,N_15345,N_18308);
and U22142 (N_22142,N_16460,N_14549);
or U22143 (N_22143,N_16911,N_13257);
xor U22144 (N_22144,N_15696,N_15497);
or U22145 (N_22145,N_18463,N_14850);
or U22146 (N_22146,N_18343,N_14338);
or U22147 (N_22147,N_18291,N_14946);
xor U22148 (N_22148,N_14526,N_13916);
or U22149 (N_22149,N_15019,N_16406);
xnor U22150 (N_22150,N_13864,N_15809);
or U22151 (N_22151,N_14708,N_14363);
nor U22152 (N_22152,N_17649,N_16093);
or U22153 (N_22153,N_14728,N_13844);
or U22154 (N_22154,N_14466,N_13884);
nand U22155 (N_22155,N_17465,N_16625);
xnor U22156 (N_22156,N_15768,N_15442);
xnor U22157 (N_22157,N_18746,N_14172);
and U22158 (N_22158,N_13644,N_18280);
or U22159 (N_22159,N_16546,N_13496);
nor U22160 (N_22160,N_15222,N_15211);
nor U22161 (N_22161,N_13310,N_16339);
nor U22162 (N_22162,N_13172,N_16287);
xor U22163 (N_22163,N_15450,N_18476);
xor U22164 (N_22164,N_12958,N_16423);
nand U22165 (N_22165,N_14809,N_15556);
nor U22166 (N_22166,N_16900,N_14614);
and U22167 (N_22167,N_18731,N_17386);
or U22168 (N_22168,N_12980,N_17225);
nor U22169 (N_22169,N_18615,N_17799);
nor U22170 (N_22170,N_16227,N_18101);
xor U22171 (N_22171,N_13148,N_18464);
nor U22172 (N_22172,N_15129,N_17446);
and U22173 (N_22173,N_18043,N_16539);
or U22174 (N_22174,N_15023,N_16700);
nor U22175 (N_22175,N_17125,N_17588);
nor U22176 (N_22176,N_16620,N_12842);
and U22177 (N_22177,N_17146,N_15321);
or U22178 (N_22178,N_14271,N_18480);
nand U22179 (N_22179,N_13389,N_18531);
xnor U22180 (N_22180,N_15419,N_16032);
nand U22181 (N_22181,N_14876,N_17557);
nor U22182 (N_22182,N_15006,N_14147);
and U22183 (N_22183,N_16165,N_16735);
xnor U22184 (N_22184,N_17088,N_18521);
nand U22185 (N_22185,N_16957,N_18456);
nor U22186 (N_22186,N_14293,N_14446);
or U22187 (N_22187,N_13279,N_12860);
xor U22188 (N_22188,N_16686,N_15217);
xor U22189 (N_22189,N_17207,N_17882);
nand U22190 (N_22190,N_13727,N_13556);
and U22191 (N_22191,N_13002,N_13057);
xnor U22192 (N_22192,N_13216,N_12664);
xor U22193 (N_22193,N_16707,N_17443);
nor U22194 (N_22194,N_16940,N_17174);
nand U22195 (N_22195,N_14716,N_18532);
and U22196 (N_22196,N_13290,N_18016);
xor U22197 (N_22197,N_12578,N_13325);
or U22198 (N_22198,N_13503,N_13828);
or U22199 (N_22199,N_15102,N_13999);
and U22200 (N_22200,N_16045,N_12707);
nor U22201 (N_22201,N_12841,N_17055);
nor U22202 (N_22202,N_15978,N_18165);
nor U22203 (N_22203,N_13612,N_17524);
and U22204 (N_22204,N_17659,N_17392);
nor U22205 (N_22205,N_12811,N_14182);
and U22206 (N_22206,N_15421,N_15981);
and U22207 (N_22207,N_16421,N_14884);
xnor U22208 (N_22208,N_18461,N_18206);
nand U22209 (N_22209,N_14593,N_13511);
or U22210 (N_22210,N_17202,N_14478);
nor U22211 (N_22211,N_13051,N_15058);
or U22212 (N_22212,N_15379,N_16087);
xnor U22213 (N_22213,N_15193,N_18416);
nand U22214 (N_22214,N_15004,N_13343);
nor U22215 (N_22215,N_14393,N_15971);
nor U22216 (N_22216,N_14047,N_17643);
nor U22217 (N_22217,N_18424,N_12602);
nor U22218 (N_22218,N_14738,N_13554);
or U22219 (N_22219,N_14752,N_15656);
and U22220 (N_22220,N_14678,N_13567);
or U22221 (N_22221,N_18492,N_14723);
nor U22222 (N_22222,N_18616,N_13466);
or U22223 (N_22223,N_16356,N_17351);
xor U22224 (N_22224,N_14471,N_15610);
xnor U22225 (N_22225,N_18412,N_14387);
nand U22226 (N_22226,N_13084,N_13209);
and U22227 (N_22227,N_15254,N_18248);
nand U22228 (N_22228,N_18648,N_12560);
nor U22229 (N_22229,N_15068,N_16491);
nor U22230 (N_22230,N_15377,N_15826);
nor U22231 (N_22231,N_16745,N_18196);
xnor U22232 (N_22232,N_12916,N_16104);
or U22233 (N_22233,N_17751,N_17804);
and U22234 (N_22234,N_15766,N_15617);
nor U22235 (N_22235,N_13952,N_15146);
and U22236 (N_22236,N_12724,N_15046);
nor U22237 (N_22237,N_16379,N_14094);
xor U22238 (N_22238,N_16979,N_15333);
nand U22239 (N_22239,N_18341,N_17774);
xor U22240 (N_22240,N_18373,N_15230);
xor U22241 (N_22241,N_18631,N_17420);
xor U22242 (N_22242,N_18509,N_13506);
or U22243 (N_22243,N_16160,N_17044);
nor U22244 (N_22244,N_12633,N_16564);
xnor U22245 (N_22245,N_16301,N_13154);
and U22246 (N_22246,N_14331,N_13485);
xnor U22247 (N_22247,N_12925,N_14570);
nand U22248 (N_22248,N_16852,N_12939);
or U22249 (N_22249,N_13761,N_17014);
nor U22250 (N_22250,N_14712,N_18505);
xor U22251 (N_22251,N_14502,N_17473);
xnor U22252 (N_22252,N_18492,N_18079);
nand U22253 (N_22253,N_17661,N_18234);
nor U22254 (N_22254,N_14388,N_18185);
xnor U22255 (N_22255,N_18341,N_12966);
and U22256 (N_22256,N_14093,N_14370);
nand U22257 (N_22257,N_15360,N_14953);
or U22258 (N_22258,N_14939,N_14874);
xnor U22259 (N_22259,N_18293,N_16414);
xnor U22260 (N_22260,N_12650,N_15252);
and U22261 (N_22261,N_18288,N_17748);
nor U22262 (N_22262,N_18715,N_14096);
nor U22263 (N_22263,N_13551,N_15389);
nor U22264 (N_22264,N_17987,N_17584);
and U22265 (N_22265,N_12787,N_15956);
and U22266 (N_22266,N_12881,N_17061);
or U22267 (N_22267,N_13949,N_13322);
or U22268 (N_22268,N_14480,N_16015);
nor U22269 (N_22269,N_12713,N_14503);
and U22270 (N_22270,N_16295,N_18710);
nor U22271 (N_22271,N_16873,N_13012);
nand U22272 (N_22272,N_13784,N_15093);
nor U22273 (N_22273,N_14809,N_12872);
or U22274 (N_22274,N_13367,N_17985);
and U22275 (N_22275,N_14321,N_18212);
and U22276 (N_22276,N_18583,N_16965);
and U22277 (N_22277,N_13847,N_14153);
and U22278 (N_22278,N_14284,N_15404);
or U22279 (N_22279,N_16033,N_14912);
and U22280 (N_22280,N_16120,N_12618);
xor U22281 (N_22281,N_14244,N_13566);
nor U22282 (N_22282,N_12971,N_17017);
nand U22283 (N_22283,N_18217,N_17689);
nor U22284 (N_22284,N_17319,N_16637);
xor U22285 (N_22285,N_13012,N_18102);
or U22286 (N_22286,N_16862,N_12786);
or U22287 (N_22287,N_12961,N_15157);
nand U22288 (N_22288,N_15646,N_15659);
xnor U22289 (N_22289,N_17044,N_18641);
nor U22290 (N_22290,N_12771,N_13722);
and U22291 (N_22291,N_15238,N_17105);
nand U22292 (N_22292,N_14453,N_16402);
nor U22293 (N_22293,N_16671,N_17234);
xnor U22294 (N_22294,N_17970,N_13670);
nand U22295 (N_22295,N_17551,N_16044);
or U22296 (N_22296,N_18600,N_17434);
nor U22297 (N_22297,N_12743,N_15526);
or U22298 (N_22298,N_13632,N_13207);
xnor U22299 (N_22299,N_12787,N_15083);
or U22300 (N_22300,N_13157,N_14014);
nand U22301 (N_22301,N_13838,N_12922);
nor U22302 (N_22302,N_16436,N_16827);
xnor U22303 (N_22303,N_17963,N_13931);
nor U22304 (N_22304,N_17285,N_14303);
or U22305 (N_22305,N_12630,N_13682);
xnor U22306 (N_22306,N_13404,N_13173);
or U22307 (N_22307,N_17294,N_13248);
and U22308 (N_22308,N_17283,N_18267);
or U22309 (N_22309,N_13395,N_17298);
and U22310 (N_22310,N_17271,N_18440);
and U22311 (N_22311,N_14829,N_16532);
nor U22312 (N_22312,N_14035,N_16943);
nand U22313 (N_22313,N_14438,N_14373);
and U22314 (N_22314,N_18675,N_18183);
or U22315 (N_22315,N_17715,N_14440);
xnor U22316 (N_22316,N_16243,N_17584);
xnor U22317 (N_22317,N_13532,N_18192);
nor U22318 (N_22318,N_14376,N_15271);
or U22319 (N_22319,N_16455,N_17179);
xnor U22320 (N_22320,N_14063,N_14132);
nor U22321 (N_22321,N_13892,N_14793);
and U22322 (N_22322,N_17520,N_14331);
or U22323 (N_22323,N_15167,N_15165);
nor U22324 (N_22324,N_14712,N_17782);
or U22325 (N_22325,N_17433,N_14382);
xor U22326 (N_22326,N_16367,N_17581);
or U22327 (N_22327,N_15200,N_15252);
nand U22328 (N_22328,N_15768,N_17869);
nand U22329 (N_22329,N_14680,N_18137);
and U22330 (N_22330,N_13019,N_14705);
nor U22331 (N_22331,N_16609,N_13027);
nand U22332 (N_22332,N_16228,N_18420);
nand U22333 (N_22333,N_15604,N_15979);
nand U22334 (N_22334,N_18055,N_16042);
nand U22335 (N_22335,N_17725,N_18452);
or U22336 (N_22336,N_15565,N_18516);
or U22337 (N_22337,N_16348,N_14661);
and U22338 (N_22338,N_16300,N_15753);
or U22339 (N_22339,N_15748,N_15092);
or U22340 (N_22340,N_13017,N_12551);
or U22341 (N_22341,N_14017,N_15284);
xor U22342 (N_22342,N_13104,N_15681);
and U22343 (N_22343,N_15986,N_17904);
or U22344 (N_22344,N_18249,N_15951);
nand U22345 (N_22345,N_13993,N_14580);
nand U22346 (N_22346,N_16377,N_17153);
or U22347 (N_22347,N_16778,N_12736);
nand U22348 (N_22348,N_15067,N_18242);
and U22349 (N_22349,N_13325,N_15950);
or U22350 (N_22350,N_16333,N_17707);
xor U22351 (N_22351,N_18486,N_13077);
nand U22352 (N_22352,N_15592,N_13790);
and U22353 (N_22353,N_15550,N_14168);
nand U22354 (N_22354,N_14209,N_13843);
xnor U22355 (N_22355,N_17228,N_18078);
nand U22356 (N_22356,N_12913,N_16197);
and U22357 (N_22357,N_14378,N_17629);
xor U22358 (N_22358,N_18407,N_14314);
or U22359 (N_22359,N_15591,N_16709);
or U22360 (N_22360,N_13224,N_12792);
or U22361 (N_22361,N_17560,N_14734);
nor U22362 (N_22362,N_15696,N_14698);
or U22363 (N_22363,N_15080,N_18627);
xor U22364 (N_22364,N_17791,N_14200);
or U22365 (N_22365,N_12756,N_16995);
nor U22366 (N_22366,N_18083,N_12905);
nand U22367 (N_22367,N_12889,N_16299);
and U22368 (N_22368,N_18512,N_18574);
or U22369 (N_22369,N_18746,N_14582);
and U22370 (N_22370,N_14842,N_14237);
nand U22371 (N_22371,N_16033,N_16693);
xor U22372 (N_22372,N_14718,N_18259);
or U22373 (N_22373,N_14177,N_14973);
nand U22374 (N_22374,N_13075,N_13676);
or U22375 (N_22375,N_13027,N_15211);
and U22376 (N_22376,N_15446,N_17555);
xor U22377 (N_22377,N_15026,N_15629);
and U22378 (N_22378,N_13326,N_14860);
nand U22379 (N_22379,N_14129,N_17087);
nand U22380 (N_22380,N_15278,N_17160);
or U22381 (N_22381,N_18404,N_17252);
nor U22382 (N_22382,N_16698,N_16308);
and U22383 (N_22383,N_12539,N_15060);
nand U22384 (N_22384,N_15479,N_16455);
nand U22385 (N_22385,N_13674,N_18726);
or U22386 (N_22386,N_16306,N_14463);
nor U22387 (N_22387,N_13289,N_14454);
and U22388 (N_22388,N_17445,N_14182);
nor U22389 (N_22389,N_18562,N_13182);
or U22390 (N_22390,N_16765,N_16846);
nor U22391 (N_22391,N_16964,N_16254);
nand U22392 (N_22392,N_15320,N_16951);
and U22393 (N_22393,N_14657,N_18009);
xor U22394 (N_22394,N_18494,N_13746);
xnor U22395 (N_22395,N_13545,N_16445);
nor U22396 (N_22396,N_18547,N_13744);
nor U22397 (N_22397,N_16155,N_17831);
nor U22398 (N_22398,N_14339,N_12530);
and U22399 (N_22399,N_16223,N_12625);
nor U22400 (N_22400,N_16781,N_13877);
or U22401 (N_22401,N_18423,N_16930);
nand U22402 (N_22402,N_14785,N_14606);
and U22403 (N_22403,N_13800,N_17574);
xor U22404 (N_22404,N_17425,N_15526);
xnor U22405 (N_22405,N_18108,N_14278);
nand U22406 (N_22406,N_17340,N_12869);
or U22407 (N_22407,N_17606,N_17588);
and U22408 (N_22408,N_18419,N_17602);
nor U22409 (N_22409,N_12726,N_14394);
or U22410 (N_22410,N_17124,N_16033);
xor U22411 (N_22411,N_12893,N_17779);
nor U22412 (N_22412,N_15132,N_17610);
or U22413 (N_22413,N_14486,N_12802);
nand U22414 (N_22414,N_15410,N_16477);
nor U22415 (N_22415,N_13964,N_13896);
nand U22416 (N_22416,N_16485,N_12815);
xor U22417 (N_22417,N_13987,N_16530);
xor U22418 (N_22418,N_16979,N_13347);
and U22419 (N_22419,N_17797,N_14737);
nand U22420 (N_22420,N_15180,N_12838);
nor U22421 (N_22421,N_18221,N_18491);
xnor U22422 (N_22422,N_15899,N_18487);
or U22423 (N_22423,N_18127,N_13601);
xor U22424 (N_22424,N_13588,N_17144);
xor U22425 (N_22425,N_14198,N_17038);
and U22426 (N_22426,N_13365,N_13696);
nor U22427 (N_22427,N_17562,N_16574);
and U22428 (N_22428,N_17175,N_12914);
xor U22429 (N_22429,N_18227,N_13212);
nor U22430 (N_22430,N_18600,N_18695);
or U22431 (N_22431,N_16660,N_16204);
nor U22432 (N_22432,N_17492,N_12666);
xor U22433 (N_22433,N_17266,N_14664);
or U22434 (N_22434,N_18652,N_12994);
or U22435 (N_22435,N_15794,N_17688);
nand U22436 (N_22436,N_18072,N_17017);
nor U22437 (N_22437,N_15536,N_14176);
or U22438 (N_22438,N_13457,N_14311);
and U22439 (N_22439,N_15021,N_17119);
xnor U22440 (N_22440,N_16577,N_16593);
nor U22441 (N_22441,N_12907,N_15040);
nand U22442 (N_22442,N_13419,N_14027);
or U22443 (N_22443,N_15165,N_15114);
nand U22444 (N_22444,N_14228,N_17124);
and U22445 (N_22445,N_18058,N_13798);
nand U22446 (N_22446,N_14218,N_12585);
or U22447 (N_22447,N_14689,N_15283);
nor U22448 (N_22448,N_15299,N_12697);
or U22449 (N_22449,N_13856,N_15660);
xnor U22450 (N_22450,N_16409,N_13285);
and U22451 (N_22451,N_12814,N_16555);
xnor U22452 (N_22452,N_16437,N_15194);
nor U22453 (N_22453,N_15676,N_16831);
nor U22454 (N_22454,N_13053,N_14982);
or U22455 (N_22455,N_13776,N_16164);
nand U22456 (N_22456,N_17224,N_12896);
and U22457 (N_22457,N_12680,N_13176);
xor U22458 (N_22458,N_16983,N_13714);
nor U22459 (N_22459,N_12862,N_18488);
and U22460 (N_22460,N_14288,N_13782);
or U22461 (N_22461,N_16857,N_17107);
or U22462 (N_22462,N_17434,N_13113);
nand U22463 (N_22463,N_16559,N_13563);
or U22464 (N_22464,N_18592,N_15780);
xnor U22465 (N_22465,N_17989,N_16285);
and U22466 (N_22466,N_15748,N_17799);
xnor U22467 (N_22467,N_16034,N_17534);
or U22468 (N_22468,N_17344,N_15678);
nor U22469 (N_22469,N_17049,N_16139);
and U22470 (N_22470,N_15539,N_17650);
nand U22471 (N_22471,N_15538,N_14696);
nor U22472 (N_22472,N_14365,N_17472);
nor U22473 (N_22473,N_18492,N_18344);
xor U22474 (N_22474,N_14776,N_17959);
nand U22475 (N_22475,N_17125,N_12606);
nand U22476 (N_22476,N_14678,N_15778);
nor U22477 (N_22477,N_16954,N_13823);
nand U22478 (N_22478,N_14826,N_13519);
nor U22479 (N_22479,N_13812,N_17278);
or U22480 (N_22480,N_12926,N_14722);
nand U22481 (N_22481,N_18027,N_18060);
xnor U22482 (N_22482,N_18131,N_17827);
nor U22483 (N_22483,N_14858,N_13775);
nor U22484 (N_22484,N_15199,N_13694);
nor U22485 (N_22485,N_15224,N_14331);
or U22486 (N_22486,N_13785,N_12994);
xnor U22487 (N_22487,N_16569,N_16359);
or U22488 (N_22488,N_16126,N_13118);
or U22489 (N_22489,N_17783,N_15424);
nor U22490 (N_22490,N_14414,N_18510);
or U22491 (N_22491,N_16028,N_16171);
and U22492 (N_22492,N_13258,N_16667);
nor U22493 (N_22493,N_17776,N_13886);
xnor U22494 (N_22494,N_18532,N_16597);
nand U22495 (N_22495,N_18568,N_12863);
nand U22496 (N_22496,N_18657,N_14127);
nand U22497 (N_22497,N_15992,N_15909);
and U22498 (N_22498,N_14407,N_16903);
and U22499 (N_22499,N_18469,N_14210);
and U22500 (N_22500,N_18041,N_15281);
and U22501 (N_22501,N_17452,N_13593);
and U22502 (N_22502,N_16352,N_18583);
nand U22503 (N_22503,N_13192,N_16827);
nor U22504 (N_22504,N_18187,N_12646);
nor U22505 (N_22505,N_18486,N_18548);
or U22506 (N_22506,N_16421,N_18385);
xnor U22507 (N_22507,N_16903,N_15428);
and U22508 (N_22508,N_18513,N_14034);
nand U22509 (N_22509,N_12970,N_12810);
nor U22510 (N_22510,N_15681,N_17593);
and U22511 (N_22511,N_14576,N_12906);
and U22512 (N_22512,N_16087,N_17389);
nor U22513 (N_22513,N_13654,N_14251);
or U22514 (N_22514,N_18559,N_16357);
and U22515 (N_22515,N_14426,N_16550);
nand U22516 (N_22516,N_14336,N_16599);
xnor U22517 (N_22517,N_13834,N_17986);
xnor U22518 (N_22518,N_17585,N_17473);
or U22519 (N_22519,N_16612,N_17227);
nand U22520 (N_22520,N_17969,N_16758);
or U22521 (N_22521,N_14639,N_18330);
nand U22522 (N_22522,N_16057,N_18484);
and U22523 (N_22523,N_13495,N_15316);
or U22524 (N_22524,N_14832,N_14775);
nor U22525 (N_22525,N_15433,N_17715);
and U22526 (N_22526,N_14760,N_14683);
nor U22527 (N_22527,N_17173,N_17897);
xor U22528 (N_22528,N_13363,N_16961);
nand U22529 (N_22529,N_13727,N_18334);
or U22530 (N_22530,N_17627,N_14801);
and U22531 (N_22531,N_12523,N_16441);
and U22532 (N_22532,N_17738,N_14119);
nor U22533 (N_22533,N_13375,N_13452);
nand U22534 (N_22534,N_15860,N_14142);
nor U22535 (N_22535,N_18220,N_13131);
nor U22536 (N_22536,N_16587,N_18423);
nor U22537 (N_22537,N_16382,N_12915);
xor U22538 (N_22538,N_16696,N_16205);
nor U22539 (N_22539,N_14837,N_16308);
nand U22540 (N_22540,N_16051,N_13660);
or U22541 (N_22541,N_12778,N_13746);
nand U22542 (N_22542,N_13732,N_16966);
and U22543 (N_22543,N_14585,N_18468);
or U22544 (N_22544,N_13390,N_13230);
nor U22545 (N_22545,N_16824,N_16157);
or U22546 (N_22546,N_13003,N_14083);
or U22547 (N_22547,N_12531,N_14375);
xor U22548 (N_22548,N_14321,N_16427);
nor U22549 (N_22549,N_14412,N_17765);
or U22550 (N_22550,N_16153,N_17259);
and U22551 (N_22551,N_12644,N_16692);
xor U22552 (N_22552,N_16037,N_13716);
nand U22553 (N_22553,N_14093,N_14048);
or U22554 (N_22554,N_13206,N_12882);
nand U22555 (N_22555,N_17354,N_13247);
and U22556 (N_22556,N_16625,N_13283);
xnor U22557 (N_22557,N_18515,N_15663);
or U22558 (N_22558,N_18109,N_17719);
nor U22559 (N_22559,N_18744,N_14648);
nor U22560 (N_22560,N_18534,N_16673);
or U22561 (N_22561,N_17702,N_14351);
xnor U22562 (N_22562,N_15515,N_12670);
nand U22563 (N_22563,N_13229,N_13015);
nor U22564 (N_22564,N_13657,N_15246);
and U22565 (N_22565,N_17111,N_16834);
nor U22566 (N_22566,N_16423,N_17300);
and U22567 (N_22567,N_14564,N_17855);
or U22568 (N_22568,N_14385,N_12917);
nand U22569 (N_22569,N_15737,N_13147);
nand U22570 (N_22570,N_18053,N_16433);
nand U22571 (N_22571,N_15443,N_13809);
nor U22572 (N_22572,N_17173,N_16408);
nand U22573 (N_22573,N_17891,N_16009);
nand U22574 (N_22574,N_16205,N_16508);
or U22575 (N_22575,N_16681,N_13995);
or U22576 (N_22576,N_13623,N_16977);
nand U22577 (N_22577,N_17053,N_14591);
nand U22578 (N_22578,N_12746,N_14945);
xor U22579 (N_22579,N_13173,N_18251);
or U22580 (N_22580,N_14938,N_14401);
nor U22581 (N_22581,N_12703,N_18692);
and U22582 (N_22582,N_15117,N_15710);
xnor U22583 (N_22583,N_14500,N_15697);
and U22584 (N_22584,N_17952,N_12900);
nand U22585 (N_22585,N_17988,N_18649);
nor U22586 (N_22586,N_12989,N_16320);
and U22587 (N_22587,N_15289,N_13722);
and U22588 (N_22588,N_14073,N_17496);
or U22589 (N_22589,N_13744,N_15099);
xnor U22590 (N_22590,N_12848,N_15755);
nor U22591 (N_22591,N_14209,N_12725);
xor U22592 (N_22592,N_16161,N_18159);
nor U22593 (N_22593,N_17660,N_17598);
and U22594 (N_22594,N_14042,N_18468);
nand U22595 (N_22595,N_18012,N_16159);
nor U22596 (N_22596,N_14776,N_16988);
or U22597 (N_22597,N_17867,N_15639);
or U22598 (N_22598,N_15581,N_13727);
nand U22599 (N_22599,N_14260,N_17355);
nor U22600 (N_22600,N_12641,N_17494);
xor U22601 (N_22601,N_18341,N_18403);
xnor U22602 (N_22602,N_14153,N_15874);
nor U22603 (N_22603,N_18177,N_16072);
xor U22604 (N_22604,N_17831,N_12729);
nor U22605 (N_22605,N_14416,N_14820);
nor U22606 (N_22606,N_16260,N_14965);
nand U22607 (N_22607,N_12918,N_17567);
xor U22608 (N_22608,N_14426,N_15915);
xor U22609 (N_22609,N_17981,N_15391);
and U22610 (N_22610,N_12622,N_18129);
nand U22611 (N_22611,N_17590,N_14100);
xnor U22612 (N_22612,N_13183,N_17159);
nand U22613 (N_22613,N_14936,N_12509);
xor U22614 (N_22614,N_18733,N_14842);
and U22615 (N_22615,N_16320,N_14300);
and U22616 (N_22616,N_16681,N_13708);
and U22617 (N_22617,N_13978,N_17751);
nor U22618 (N_22618,N_14552,N_13669);
or U22619 (N_22619,N_14048,N_16317);
nor U22620 (N_22620,N_17341,N_16828);
xnor U22621 (N_22621,N_16349,N_18535);
xor U22622 (N_22622,N_15995,N_18673);
or U22623 (N_22623,N_13359,N_16148);
nand U22624 (N_22624,N_17333,N_18381);
nand U22625 (N_22625,N_17556,N_12966);
xnor U22626 (N_22626,N_17482,N_18176);
and U22627 (N_22627,N_14286,N_17128);
nor U22628 (N_22628,N_14939,N_14440);
or U22629 (N_22629,N_13955,N_16706);
and U22630 (N_22630,N_15836,N_15052);
and U22631 (N_22631,N_17657,N_17640);
or U22632 (N_22632,N_16861,N_14818);
nand U22633 (N_22633,N_17905,N_17063);
or U22634 (N_22634,N_17630,N_16870);
and U22635 (N_22635,N_15257,N_16718);
nand U22636 (N_22636,N_16558,N_17786);
nor U22637 (N_22637,N_18211,N_15429);
xor U22638 (N_22638,N_18593,N_14372);
or U22639 (N_22639,N_17599,N_18627);
nand U22640 (N_22640,N_13427,N_16078);
and U22641 (N_22641,N_14673,N_12894);
nand U22642 (N_22642,N_18683,N_18235);
nand U22643 (N_22643,N_18269,N_17194);
or U22644 (N_22644,N_17753,N_18127);
and U22645 (N_22645,N_12722,N_13526);
nand U22646 (N_22646,N_16324,N_18502);
xnor U22647 (N_22647,N_15067,N_13025);
and U22648 (N_22648,N_18425,N_12659);
nor U22649 (N_22649,N_18008,N_17280);
and U22650 (N_22650,N_13836,N_15345);
nor U22651 (N_22651,N_13205,N_13316);
or U22652 (N_22652,N_14767,N_17611);
nand U22653 (N_22653,N_15690,N_17297);
and U22654 (N_22654,N_15324,N_13820);
or U22655 (N_22655,N_15019,N_18202);
or U22656 (N_22656,N_14652,N_13199);
or U22657 (N_22657,N_13005,N_16417);
nor U22658 (N_22658,N_17516,N_16366);
nand U22659 (N_22659,N_13523,N_14719);
and U22660 (N_22660,N_15217,N_16730);
or U22661 (N_22661,N_17675,N_13477);
or U22662 (N_22662,N_18474,N_17074);
xnor U22663 (N_22663,N_16987,N_12938);
xnor U22664 (N_22664,N_13670,N_18174);
xor U22665 (N_22665,N_14630,N_14806);
nand U22666 (N_22666,N_17512,N_15459);
nor U22667 (N_22667,N_16240,N_13702);
nor U22668 (N_22668,N_17422,N_14156);
nand U22669 (N_22669,N_14182,N_15113);
or U22670 (N_22670,N_17145,N_18313);
nor U22671 (N_22671,N_14150,N_13594);
or U22672 (N_22672,N_17015,N_14498);
xor U22673 (N_22673,N_15348,N_15482);
nand U22674 (N_22674,N_15227,N_17894);
and U22675 (N_22675,N_14849,N_13669);
xnor U22676 (N_22676,N_12766,N_15806);
nor U22677 (N_22677,N_17137,N_13554);
and U22678 (N_22678,N_14831,N_17322);
xnor U22679 (N_22679,N_15768,N_13641);
xnor U22680 (N_22680,N_18379,N_15046);
or U22681 (N_22681,N_15920,N_16050);
and U22682 (N_22682,N_14698,N_16535);
and U22683 (N_22683,N_16667,N_16201);
and U22684 (N_22684,N_15841,N_17927);
nor U22685 (N_22685,N_18617,N_12629);
nor U22686 (N_22686,N_15926,N_14502);
and U22687 (N_22687,N_16924,N_18237);
or U22688 (N_22688,N_12960,N_15972);
xor U22689 (N_22689,N_17389,N_17578);
nand U22690 (N_22690,N_17911,N_18259);
nand U22691 (N_22691,N_14619,N_17404);
and U22692 (N_22692,N_13663,N_14280);
nor U22693 (N_22693,N_14037,N_14426);
or U22694 (N_22694,N_13856,N_14953);
or U22695 (N_22695,N_17224,N_18189);
nand U22696 (N_22696,N_16818,N_12782);
xor U22697 (N_22697,N_16452,N_12989);
nand U22698 (N_22698,N_14321,N_17841);
xnor U22699 (N_22699,N_15136,N_15750);
and U22700 (N_22700,N_16998,N_16893);
and U22701 (N_22701,N_13402,N_18197);
and U22702 (N_22702,N_17088,N_16803);
and U22703 (N_22703,N_14031,N_15772);
nand U22704 (N_22704,N_18442,N_17415);
xor U22705 (N_22705,N_15005,N_18212);
nand U22706 (N_22706,N_16046,N_15706);
nand U22707 (N_22707,N_14366,N_14470);
nand U22708 (N_22708,N_13661,N_18454);
or U22709 (N_22709,N_14909,N_13871);
nand U22710 (N_22710,N_18413,N_14570);
or U22711 (N_22711,N_16275,N_14620);
or U22712 (N_22712,N_13168,N_13061);
nor U22713 (N_22713,N_18055,N_14945);
or U22714 (N_22714,N_14396,N_17504);
or U22715 (N_22715,N_13103,N_13538);
and U22716 (N_22716,N_17157,N_14357);
nand U22717 (N_22717,N_15607,N_13182);
nand U22718 (N_22718,N_16518,N_18725);
nand U22719 (N_22719,N_14629,N_14898);
nand U22720 (N_22720,N_17772,N_14395);
xor U22721 (N_22721,N_16298,N_12897);
and U22722 (N_22722,N_14411,N_16818);
xnor U22723 (N_22723,N_12860,N_18320);
and U22724 (N_22724,N_18580,N_16572);
and U22725 (N_22725,N_14962,N_16188);
xor U22726 (N_22726,N_13338,N_16802);
nand U22727 (N_22727,N_12539,N_17152);
xor U22728 (N_22728,N_15643,N_17856);
nor U22729 (N_22729,N_17616,N_17594);
and U22730 (N_22730,N_17632,N_18259);
nor U22731 (N_22731,N_15014,N_17028);
and U22732 (N_22732,N_18272,N_14218);
nor U22733 (N_22733,N_12596,N_13799);
nand U22734 (N_22734,N_14900,N_12742);
xnor U22735 (N_22735,N_15481,N_16922);
or U22736 (N_22736,N_16386,N_12996);
and U22737 (N_22737,N_15000,N_16398);
or U22738 (N_22738,N_15358,N_13083);
or U22739 (N_22739,N_16794,N_17166);
nor U22740 (N_22740,N_13769,N_17143);
nor U22741 (N_22741,N_13697,N_18478);
nand U22742 (N_22742,N_18722,N_13342);
and U22743 (N_22743,N_15822,N_16367);
nor U22744 (N_22744,N_17724,N_13403);
or U22745 (N_22745,N_12795,N_15552);
and U22746 (N_22746,N_13124,N_14064);
and U22747 (N_22747,N_15124,N_12545);
or U22748 (N_22748,N_16188,N_18250);
nor U22749 (N_22749,N_17723,N_13878);
nand U22750 (N_22750,N_12566,N_12778);
nor U22751 (N_22751,N_17294,N_14596);
nor U22752 (N_22752,N_17963,N_17722);
or U22753 (N_22753,N_12614,N_13406);
nand U22754 (N_22754,N_12740,N_14175);
or U22755 (N_22755,N_14110,N_14132);
nand U22756 (N_22756,N_13841,N_14389);
nor U22757 (N_22757,N_15254,N_13653);
xnor U22758 (N_22758,N_14004,N_13224);
nand U22759 (N_22759,N_13706,N_15481);
or U22760 (N_22760,N_13371,N_17565);
nor U22761 (N_22761,N_17616,N_16313);
nand U22762 (N_22762,N_12705,N_17076);
or U22763 (N_22763,N_13854,N_13019);
nand U22764 (N_22764,N_15438,N_17983);
nor U22765 (N_22765,N_16617,N_18146);
nor U22766 (N_22766,N_15944,N_12554);
xnor U22767 (N_22767,N_14319,N_16982);
and U22768 (N_22768,N_15836,N_14451);
xnor U22769 (N_22769,N_17661,N_13644);
nor U22770 (N_22770,N_18549,N_18625);
nand U22771 (N_22771,N_13228,N_15840);
or U22772 (N_22772,N_18630,N_18671);
nand U22773 (N_22773,N_12601,N_15656);
nor U22774 (N_22774,N_14426,N_15653);
xor U22775 (N_22775,N_13903,N_12675);
and U22776 (N_22776,N_15231,N_17660);
xnor U22777 (N_22777,N_14872,N_15117);
xor U22778 (N_22778,N_13430,N_17209);
or U22779 (N_22779,N_16631,N_17422);
nor U22780 (N_22780,N_17658,N_18541);
or U22781 (N_22781,N_14214,N_16015);
xor U22782 (N_22782,N_14831,N_18050);
nor U22783 (N_22783,N_14057,N_16176);
or U22784 (N_22784,N_15846,N_13684);
nand U22785 (N_22785,N_16505,N_18712);
and U22786 (N_22786,N_13523,N_16781);
or U22787 (N_22787,N_18256,N_15414);
and U22788 (N_22788,N_13555,N_17624);
and U22789 (N_22789,N_15584,N_15367);
or U22790 (N_22790,N_18178,N_13934);
or U22791 (N_22791,N_15102,N_17281);
nand U22792 (N_22792,N_17098,N_12757);
xnor U22793 (N_22793,N_14949,N_14163);
or U22794 (N_22794,N_16235,N_13290);
and U22795 (N_22795,N_17112,N_16777);
xnor U22796 (N_22796,N_16001,N_16300);
nand U22797 (N_22797,N_15414,N_14229);
nor U22798 (N_22798,N_14241,N_14970);
or U22799 (N_22799,N_15134,N_16898);
or U22800 (N_22800,N_16774,N_14332);
nor U22801 (N_22801,N_14763,N_16647);
nand U22802 (N_22802,N_13224,N_17637);
and U22803 (N_22803,N_16772,N_13680);
and U22804 (N_22804,N_16262,N_13402);
nand U22805 (N_22805,N_16061,N_16695);
or U22806 (N_22806,N_12761,N_17747);
or U22807 (N_22807,N_15636,N_14280);
or U22808 (N_22808,N_16989,N_15412);
and U22809 (N_22809,N_13018,N_16743);
nand U22810 (N_22810,N_14779,N_16754);
or U22811 (N_22811,N_17969,N_17314);
or U22812 (N_22812,N_15751,N_12724);
xnor U22813 (N_22813,N_18026,N_15648);
and U22814 (N_22814,N_13936,N_17437);
xnor U22815 (N_22815,N_13218,N_15242);
nand U22816 (N_22816,N_16668,N_17960);
nand U22817 (N_22817,N_14044,N_12538);
or U22818 (N_22818,N_18726,N_13058);
and U22819 (N_22819,N_13069,N_16294);
and U22820 (N_22820,N_15450,N_15077);
and U22821 (N_22821,N_16694,N_15941);
xnor U22822 (N_22822,N_15634,N_15800);
and U22823 (N_22823,N_12800,N_16506);
and U22824 (N_22824,N_17349,N_15350);
and U22825 (N_22825,N_17807,N_15708);
xor U22826 (N_22826,N_16748,N_12860);
xnor U22827 (N_22827,N_16079,N_14250);
nor U22828 (N_22828,N_18695,N_12584);
nor U22829 (N_22829,N_18355,N_16976);
nand U22830 (N_22830,N_18504,N_17759);
nor U22831 (N_22831,N_16962,N_12970);
nand U22832 (N_22832,N_13612,N_18514);
nor U22833 (N_22833,N_17320,N_17300);
xor U22834 (N_22834,N_16095,N_17807);
or U22835 (N_22835,N_12948,N_17706);
or U22836 (N_22836,N_12739,N_14494);
nand U22837 (N_22837,N_12879,N_16706);
and U22838 (N_22838,N_18375,N_13901);
nor U22839 (N_22839,N_17783,N_18303);
nand U22840 (N_22840,N_18400,N_18325);
and U22841 (N_22841,N_13130,N_18650);
nand U22842 (N_22842,N_17538,N_16768);
nand U22843 (N_22843,N_16748,N_17360);
nand U22844 (N_22844,N_17225,N_14218);
xnor U22845 (N_22845,N_18103,N_18180);
and U22846 (N_22846,N_14526,N_18109);
and U22847 (N_22847,N_18370,N_13924);
and U22848 (N_22848,N_18357,N_17397);
nor U22849 (N_22849,N_18121,N_13912);
nor U22850 (N_22850,N_18492,N_12791);
or U22851 (N_22851,N_17183,N_16293);
or U22852 (N_22852,N_14909,N_15364);
nor U22853 (N_22853,N_16777,N_16393);
nor U22854 (N_22854,N_18229,N_14376);
and U22855 (N_22855,N_16661,N_15956);
or U22856 (N_22856,N_13216,N_15727);
and U22857 (N_22857,N_13990,N_12848);
and U22858 (N_22858,N_15948,N_14545);
xnor U22859 (N_22859,N_16702,N_18312);
nor U22860 (N_22860,N_16725,N_18052);
and U22861 (N_22861,N_18532,N_15049);
or U22862 (N_22862,N_14383,N_13749);
xor U22863 (N_22863,N_13784,N_12654);
or U22864 (N_22864,N_13171,N_17643);
or U22865 (N_22865,N_15202,N_18274);
nand U22866 (N_22866,N_16143,N_15667);
and U22867 (N_22867,N_15336,N_13070);
xnor U22868 (N_22868,N_13153,N_12958);
or U22869 (N_22869,N_15113,N_17729);
nor U22870 (N_22870,N_17520,N_16431);
xor U22871 (N_22871,N_14191,N_18177);
xnor U22872 (N_22872,N_15243,N_13637);
and U22873 (N_22873,N_14746,N_12843);
or U22874 (N_22874,N_13824,N_15196);
or U22875 (N_22875,N_13274,N_17482);
and U22876 (N_22876,N_16527,N_16522);
nor U22877 (N_22877,N_13877,N_16964);
nand U22878 (N_22878,N_17326,N_17899);
or U22879 (N_22879,N_18358,N_17667);
nand U22880 (N_22880,N_16333,N_16030);
or U22881 (N_22881,N_14356,N_18340);
nor U22882 (N_22882,N_12613,N_16851);
xor U22883 (N_22883,N_12660,N_14450);
and U22884 (N_22884,N_12761,N_14650);
xnor U22885 (N_22885,N_15668,N_14018);
nor U22886 (N_22886,N_15233,N_18689);
or U22887 (N_22887,N_17911,N_15302);
nor U22888 (N_22888,N_16305,N_12794);
and U22889 (N_22889,N_17990,N_18129);
xor U22890 (N_22890,N_14527,N_18468);
and U22891 (N_22891,N_13305,N_12897);
xnor U22892 (N_22892,N_18267,N_13731);
and U22893 (N_22893,N_13766,N_13830);
xor U22894 (N_22894,N_18570,N_15767);
nand U22895 (N_22895,N_13059,N_15066);
nand U22896 (N_22896,N_13104,N_14188);
xnor U22897 (N_22897,N_14025,N_16727);
and U22898 (N_22898,N_13265,N_14297);
nand U22899 (N_22899,N_16161,N_13511);
nand U22900 (N_22900,N_16898,N_15936);
and U22901 (N_22901,N_16785,N_17100);
nand U22902 (N_22902,N_15096,N_18196);
nor U22903 (N_22903,N_18499,N_14686);
xnor U22904 (N_22904,N_16096,N_16332);
or U22905 (N_22905,N_14686,N_17484);
nor U22906 (N_22906,N_17737,N_14627);
and U22907 (N_22907,N_17652,N_15122);
xnor U22908 (N_22908,N_17530,N_13617);
xnor U22909 (N_22909,N_17860,N_17173);
and U22910 (N_22910,N_16928,N_15297);
and U22911 (N_22911,N_16420,N_18557);
xor U22912 (N_22912,N_16067,N_13842);
nor U22913 (N_22913,N_15980,N_17236);
xor U22914 (N_22914,N_17810,N_12551);
nor U22915 (N_22915,N_17127,N_13904);
nand U22916 (N_22916,N_18665,N_17816);
nor U22917 (N_22917,N_16012,N_15411);
or U22918 (N_22918,N_14662,N_16108);
nor U22919 (N_22919,N_14969,N_16440);
nor U22920 (N_22920,N_12924,N_14249);
or U22921 (N_22921,N_14708,N_13173);
nor U22922 (N_22922,N_16884,N_18719);
or U22923 (N_22923,N_13819,N_13946);
xor U22924 (N_22924,N_17252,N_12790);
and U22925 (N_22925,N_16091,N_12520);
nor U22926 (N_22926,N_14760,N_12541);
and U22927 (N_22927,N_18183,N_14216);
or U22928 (N_22928,N_17596,N_17501);
nand U22929 (N_22929,N_16248,N_18658);
and U22930 (N_22930,N_12906,N_16337);
nand U22931 (N_22931,N_13833,N_14423);
nand U22932 (N_22932,N_17330,N_18211);
nor U22933 (N_22933,N_14716,N_14212);
nor U22934 (N_22934,N_18056,N_16938);
nor U22935 (N_22935,N_13142,N_14001);
nand U22936 (N_22936,N_15986,N_14804);
or U22937 (N_22937,N_16660,N_17615);
nor U22938 (N_22938,N_16574,N_13765);
nor U22939 (N_22939,N_17726,N_18345);
or U22940 (N_22940,N_13457,N_16087);
nand U22941 (N_22941,N_14343,N_15955);
nand U22942 (N_22942,N_16581,N_15459);
or U22943 (N_22943,N_13642,N_17998);
nand U22944 (N_22944,N_15188,N_14197);
nor U22945 (N_22945,N_15837,N_15933);
and U22946 (N_22946,N_17540,N_17095);
nand U22947 (N_22947,N_12825,N_17817);
and U22948 (N_22948,N_13095,N_13740);
nand U22949 (N_22949,N_15043,N_15270);
nand U22950 (N_22950,N_16383,N_18723);
xor U22951 (N_22951,N_17219,N_13240);
xor U22952 (N_22952,N_17893,N_16857);
or U22953 (N_22953,N_13299,N_15642);
nand U22954 (N_22954,N_14592,N_13286);
xnor U22955 (N_22955,N_15898,N_15742);
nand U22956 (N_22956,N_14968,N_14483);
nand U22957 (N_22957,N_13858,N_16200);
xnor U22958 (N_22958,N_16903,N_16681);
or U22959 (N_22959,N_12547,N_14322);
nand U22960 (N_22960,N_16362,N_17713);
or U22961 (N_22961,N_17260,N_14019);
nand U22962 (N_22962,N_17889,N_17996);
or U22963 (N_22963,N_16866,N_14662);
and U22964 (N_22964,N_13503,N_13228);
and U22965 (N_22965,N_16961,N_13084);
or U22966 (N_22966,N_14375,N_13499);
and U22967 (N_22967,N_16118,N_17763);
nand U22968 (N_22968,N_13594,N_15796);
nand U22969 (N_22969,N_16506,N_17567);
nand U22970 (N_22970,N_16281,N_14948);
xnor U22971 (N_22971,N_15810,N_16266);
or U22972 (N_22972,N_12870,N_12645);
or U22973 (N_22973,N_12617,N_14556);
and U22974 (N_22974,N_14644,N_16760);
xor U22975 (N_22975,N_17802,N_13631);
and U22976 (N_22976,N_13621,N_13477);
xnor U22977 (N_22977,N_16712,N_15621);
nor U22978 (N_22978,N_17323,N_12709);
or U22979 (N_22979,N_18734,N_15265);
nor U22980 (N_22980,N_15903,N_16044);
or U22981 (N_22981,N_14948,N_15521);
xnor U22982 (N_22982,N_15879,N_15989);
nor U22983 (N_22983,N_13330,N_18227);
nand U22984 (N_22984,N_13960,N_13702);
or U22985 (N_22985,N_18088,N_15952);
and U22986 (N_22986,N_18350,N_16918);
and U22987 (N_22987,N_18547,N_18518);
xnor U22988 (N_22988,N_14828,N_13148);
nand U22989 (N_22989,N_12563,N_16351);
or U22990 (N_22990,N_16931,N_17884);
xnor U22991 (N_22991,N_15692,N_15320);
nor U22992 (N_22992,N_12946,N_13052);
or U22993 (N_22993,N_17591,N_18315);
or U22994 (N_22994,N_12552,N_18321);
and U22995 (N_22995,N_18270,N_16038);
nor U22996 (N_22996,N_18523,N_14663);
xnor U22997 (N_22997,N_17982,N_14314);
xnor U22998 (N_22998,N_12789,N_13463);
xor U22999 (N_22999,N_17535,N_14643);
or U23000 (N_23000,N_17572,N_13932);
and U23001 (N_23001,N_16495,N_17242);
nor U23002 (N_23002,N_14081,N_15351);
nand U23003 (N_23003,N_12784,N_18029);
or U23004 (N_23004,N_17632,N_12792);
or U23005 (N_23005,N_12826,N_13910);
or U23006 (N_23006,N_16370,N_16185);
nand U23007 (N_23007,N_16624,N_13668);
xnor U23008 (N_23008,N_15032,N_15107);
nand U23009 (N_23009,N_15660,N_15046);
nor U23010 (N_23010,N_14126,N_12987);
or U23011 (N_23011,N_18273,N_14147);
xor U23012 (N_23012,N_15524,N_12586);
nor U23013 (N_23013,N_15040,N_17801);
nand U23014 (N_23014,N_18317,N_13906);
nor U23015 (N_23015,N_15399,N_18292);
and U23016 (N_23016,N_13471,N_18248);
nand U23017 (N_23017,N_16618,N_15547);
nor U23018 (N_23018,N_13991,N_13197);
nand U23019 (N_23019,N_16173,N_13346);
or U23020 (N_23020,N_14707,N_13190);
xnor U23021 (N_23021,N_16073,N_13135);
and U23022 (N_23022,N_18702,N_17009);
and U23023 (N_23023,N_12850,N_15446);
nand U23024 (N_23024,N_13516,N_18301);
xnor U23025 (N_23025,N_15365,N_13509);
nor U23026 (N_23026,N_14505,N_13578);
nor U23027 (N_23027,N_18407,N_16092);
xnor U23028 (N_23028,N_12679,N_14852);
nor U23029 (N_23029,N_16423,N_14157);
nor U23030 (N_23030,N_15255,N_17185);
nand U23031 (N_23031,N_14671,N_17427);
nor U23032 (N_23032,N_16507,N_18380);
nor U23033 (N_23033,N_13004,N_17321);
nand U23034 (N_23034,N_15756,N_17315);
and U23035 (N_23035,N_13787,N_13803);
xor U23036 (N_23036,N_14868,N_16317);
and U23037 (N_23037,N_18695,N_16339);
or U23038 (N_23038,N_13070,N_16878);
and U23039 (N_23039,N_16793,N_17752);
nand U23040 (N_23040,N_13472,N_13971);
and U23041 (N_23041,N_15026,N_18636);
xnor U23042 (N_23042,N_17971,N_12513);
and U23043 (N_23043,N_16757,N_17573);
and U23044 (N_23044,N_12912,N_13702);
nor U23045 (N_23045,N_12662,N_15483);
xnor U23046 (N_23046,N_14529,N_13319);
or U23047 (N_23047,N_17825,N_14986);
and U23048 (N_23048,N_15050,N_17271);
xnor U23049 (N_23049,N_12774,N_18098);
and U23050 (N_23050,N_14864,N_15223);
or U23051 (N_23051,N_17587,N_13579);
or U23052 (N_23052,N_14452,N_15665);
or U23053 (N_23053,N_12661,N_12789);
and U23054 (N_23054,N_18298,N_12527);
xor U23055 (N_23055,N_13830,N_14255);
or U23056 (N_23056,N_13215,N_15152);
xnor U23057 (N_23057,N_16208,N_16652);
nand U23058 (N_23058,N_18739,N_16919);
xnor U23059 (N_23059,N_14039,N_15238);
xnor U23060 (N_23060,N_14390,N_13348);
nand U23061 (N_23061,N_12945,N_13572);
nor U23062 (N_23062,N_18171,N_14079);
nand U23063 (N_23063,N_16517,N_15674);
nand U23064 (N_23064,N_15866,N_13009);
nor U23065 (N_23065,N_14748,N_15770);
nor U23066 (N_23066,N_18422,N_14348);
nor U23067 (N_23067,N_14519,N_17433);
nor U23068 (N_23068,N_16088,N_17979);
xor U23069 (N_23069,N_18113,N_13601);
nor U23070 (N_23070,N_14936,N_16862);
nand U23071 (N_23071,N_13073,N_14678);
nor U23072 (N_23072,N_17372,N_13467);
nor U23073 (N_23073,N_14703,N_16195);
nor U23074 (N_23074,N_16660,N_13514);
or U23075 (N_23075,N_13413,N_17194);
nand U23076 (N_23076,N_12511,N_16341);
xnor U23077 (N_23077,N_16575,N_13690);
and U23078 (N_23078,N_13100,N_17701);
nor U23079 (N_23079,N_15364,N_15523);
xnor U23080 (N_23080,N_15216,N_13036);
or U23081 (N_23081,N_18176,N_15670);
nand U23082 (N_23082,N_17302,N_16832);
xnor U23083 (N_23083,N_15231,N_14744);
and U23084 (N_23084,N_17660,N_13943);
xor U23085 (N_23085,N_15850,N_18637);
xor U23086 (N_23086,N_14261,N_18384);
nor U23087 (N_23087,N_15392,N_14421);
and U23088 (N_23088,N_13717,N_13810);
nand U23089 (N_23089,N_12791,N_16197);
nor U23090 (N_23090,N_15219,N_16525);
and U23091 (N_23091,N_15397,N_17777);
nand U23092 (N_23092,N_17666,N_18518);
nor U23093 (N_23093,N_17001,N_14648);
or U23094 (N_23094,N_16493,N_18422);
nor U23095 (N_23095,N_13824,N_15270);
xor U23096 (N_23096,N_17578,N_15051);
and U23097 (N_23097,N_17853,N_17963);
or U23098 (N_23098,N_14818,N_14661);
nand U23099 (N_23099,N_14166,N_16463);
nand U23100 (N_23100,N_12911,N_12731);
nor U23101 (N_23101,N_14692,N_15506);
or U23102 (N_23102,N_15484,N_13173);
or U23103 (N_23103,N_14898,N_17748);
xor U23104 (N_23104,N_12845,N_13974);
or U23105 (N_23105,N_16609,N_15259);
nand U23106 (N_23106,N_13593,N_13999);
xor U23107 (N_23107,N_13342,N_15910);
nor U23108 (N_23108,N_15714,N_15725);
nand U23109 (N_23109,N_13752,N_15530);
nor U23110 (N_23110,N_13599,N_18149);
nor U23111 (N_23111,N_17920,N_14906);
nor U23112 (N_23112,N_13472,N_17966);
and U23113 (N_23113,N_17545,N_15818);
or U23114 (N_23114,N_15839,N_13331);
nor U23115 (N_23115,N_18267,N_12877);
or U23116 (N_23116,N_16042,N_18163);
nor U23117 (N_23117,N_17489,N_13255);
or U23118 (N_23118,N_13854,N_15402);
nor U23119 (N_23119,N_17161,N_15324);
and U23120 (N_23120,N_15641,N_12731);
nor U23121 (N_23121,N_14295,N_15694);
and U23122 (N_23122,N_12871,N_15765);
xor U23123 (N_23123,N_15878,N_13418);
nand U23124 (N_23124,N_12754,N_18718);
nand U23125 (N_23125,N_14113,N_14472);
nor U23126 (N_23126,N_12903,N_17374);
or U23127 (N_23127,N_16974,N_17716);
or U23128 (N_23128,N_12610,N_14647);
or U23129 (N_23129,N_13617,N_17604);
xor U23130 (N_23130,N_14361,N_14534);
xnor U23131 (N_23131,N_16867,N_15764);
nand U23132 (N_23132,N_15797,N_13361);
nor U23133 (N_23133,N_14952,N_17284);
nand U23134 (N_23134,N_14485,N_17984);
nor U23135 (N_23135,N_17243,N_13021);
nor U23136 (N_23136,N_12639,N_16368);
and U23137 (N_23137,N_12555,N_15878);
or U23138 (N_23138,N_18248,N_16410);
or U23139 (N_23139,N_16560,N_13666);
or U23140 (N_23140,N_14752,N_14584);
nor U23141 (N_23141,N_14153,N_14121);
and U23142 (N_23142,N_15674,N_15363);
or U23143 (N_23143,N_17016,N_15259);
nand U23144 (N_23144,N_17177,N_15150);
nor U23145 (N_23145,N_15634,N_14779);
and U23146 (N_23146,N_16861,N_14738);
nor U23147 (N_23147,N_14242,N_13332);
or U23148 (N_23148,N_16673,N_15306);
nor U23149 (N_23149,N_16511,N_18031);
nor U23150 (N_23150,N_12998,N_17382);
nand U23151 (N_23151,N_16765,N_14338);
nor U23152 (N_23152,N_15614,N_12834);
nand U23153 (N_23153,N_14448,N_18682);
and U23154 (N_23154,N_18155,N_17544);
or U23155 (N_23155,N_14683,N_12520);
nor U23156 (N_23156,N_18070,N_18113);
and U23157 (N_23157,N_13703,N_12647);
and U23158 (N_23158,N_14252,N_13953);
and U23159 (N_23159,N_12914,N_12761);
and U23160 (N_23160,N_13336,N_15126);
or U23161 (N_23161,N_17897,N_17179);
nand U23162 (N_23162,N_18696,N_17456);
and U23163 (N_23163,N_16212,N_16209);
and U23164 (N_23164,N_14393,N_15653);
or U23165 (N_23165,N_16259,N_14891);
or U23166 (N_23166,N_18149,N_18134);
xor U23167 (N_23167,N_15093,N_16042);
and U23168 (N_23168,N_14302,N_12868);
or U23169 (N_23169,N_17258,N_18157);
xnor U23170 (N_23170,N_15839,N_14077);
or U23171 (N_23171,N_14595,N_13384);
xor U23172 (N_23172,N_13032,N_17768);
and U23173 (N_23173,N_17724,N_17741);
and U23174 (N_23174,N_13968,N_13674);
nand U23175 (N_23175,N_13427,N_15265);
or U23176 (N_23176,N_16822,N_15905);
and U23177 (N_23177,N_18529,N_13214);
nand U23178 (N_23178,N_17685,N_14316);
and U23179 (N_23179,N_16850,N_13842);
nor U23180 (N_23180,N_14354,N_16452);
nand U23181 (N_23181,N_16850,N_14943);
nand U23182 (N_23182,N_18012,N_16703);
and U23183 (N_23183,N_14407,N_17073);
or U23184 (N_23184,N_14204,N_13226);
and U23185 (N_23185,N_14040,N_15027);
xor U23186 (N_23186,N_17559,N_17179);
nand U23187 (N_23187,N_14221,N_18149);
xor U23188 (N_23188,N_16237,N_16069);
nor U23189 (N_23189,N_15416,N_16811);
nand U23190 (N_23190,N_14788,N_13475);
xor U23191 (N_23191,N_16777,N_12585);
nor U23192 (N_23192,N_17983,N_18420);
nor U23193 (N_23193,N_13286,N_17811);
nor U23194 (N_23194,N_17813,N_13891);
or U23195 (N_23195,N_18702,N_14771);
nor U23196 (N_23196,N_14467,N_17964);
nand U23197 (N_23197,N_17787,N_13334);
nand U23198 (N_23198,N_18630,N_13253);
xor U23199 (N_23199,N_13514,N_18247);
or U23200 (N_23200,N_14602,N_15960);
or U23201 (N_23201,N_14164,N_12982);
nand U23202 (N_23202,N_12951,N_15130);
nor U23203 (N_23203,N_14047,N_17119);
nor U23204 (N_23204,N_15485,N_13343);
and U23205 (N_23205,N_14297,N_15508);
nor U23206 (N_23206,N_15302,N_14312);
xor U23207 (N_23207,N_17055,N_13720);
nand U23208 (N_23208,N_15719,N_16121);
nand U23209 (N_23209,N_14824,N_12733);
nor U23210 (N_23210,N_13901,N_15158);
nand U23211 (N_23211,N_14539,N_16509);
or U23212 (N_23212,N_14029,N_17804);
nand U23213 (N_23213,N_13591,N_14323);
or U23214 (N_23214,N_18025,N_12617);
or U23215 (N_23215,N_12751,N_14275);
or U23216 (N_23216,N_17362,N_13615);
xnor U23217 (N_23217,N_16908,N_14277);
nor U23218 (N_23218,N_18415,N_14093);
nor U23219 (N_23219,N_13867,N_14458);
nor U23220 (N_23220,N_17203,N_18543);
and U23221 (N_23221,N_14758,N_14581);
nand U23222 (N_23222,N_17519,N_16209);
and U23223 (N_23223,N_15009,N_13822);
nor U23224 (N_23224,N_14713,N_13454);
nand U23225 (N_23225,N_16681,N_16736);
xor U23226 (N_23226,N_17166,N_16932);
nor U23227 (N_23227,N_13303,N_18681);
and U23228 (N_23228,N_15700,N_18218);
nor U23229 (N_23229,N_16179,N_14793);
and U23230 (N_23230,N_18132,N_13457);
xnor U23231 (N_23231,N_18036,N_13714);
nand U23232 (N_23232,N_16883,N_13096);
nor U23233 (N_23233,N_15814,N_13867);
xnor U23234 (N_23234,N_14002,N_18033);
or U23235 (N_23235,N_13711,N_15033);
xnor U23236 (N_23236,N_18562,N_14128);
and U23237 (N_23237,N_12989,N_14110);
nor U23238 (N_23238,N_13972,N_14407);
nor U23239 (N_23239,N_13119,N_13884);
and U23240 (N_23240,N_15547,N_14997);
nor U23241 (N_23241,N_15613,N_15342);
or U23242 (N_23242,N_17993,N_13619);
xnor U23243 (N_23243,N_17029,N_15111);
or U23244 (N_23244,N_18549,N_14621);
xnor U23245 (N_23245,N_16785,N_17974);
or U23246 (N_23246,N_12823,N_16868);
nor U23247 (N_23247,N_17981,N_18286);
and U23248 (N_23248,N_18169,N_18652);
or U23249 (N_23249,N_15632,N_16402);
and U23250 (N_23250,N_16312,N_17704);
or U23251 (N_23251,N_17911,N_12842);
or U23252 (N_23252,N_16673,N_13649);
xor U23253 (N_23253,N_18310,N_15175);
nor U23254 (N_23254,N_16094,N_18448);
nand U23255 (N_23255,N_14417,N_15007);
xor U23256 (N_23256,N_14529,N_13794);
and U23257 (N_23257,N_14132,N_16049);
xnor U23258 (N_23258,N_13980,N_16543);
or U23259 (N_23259,N_18660,N_13191);
xor U23260 (N_23260,N_15867,N_15415);
and U23261 (N_23261,N_18500,N_18494);
xnor U23262 (N_23262,N_14851,N_15011);
nand U23263 (N_23263,N_14534,N_15538);
and U23264 (N_23264,N_15911,N_13363);
or U23265 (N_23265,N_14747,N_17809);
or U23266 (N_23266,N_17281,N_16573);
and U23267 (N_23267,N_18705,N_12739);
xnor U23268 (N_23268,N_12776,N_15909);
nand U23269 (N_23269,N_16388,N_14474);
nor U23270 (N_23270,N_16690,N_15356);
and U23271 (N_23271,N_14143,N_17492);
xnor U23272 (N_23272,N_16754,N_17182);
or U23273 (N_23273,N_15037,N_13281);
and U23274 (N_23274,N_14592,N_15844);
nand U23275 (N_23275,N_15909,N_15336);
nor U23276 (N_23276,N_12785,N_18237);
or U23277 (N_23277,N_15418,N_17016);
xor U23278 (N_23278,N_13341,N_12716);
and U23279 (N_23279,N_13372,N_18474);
and U23280 (N_23280,N_14421,N_18701);
xor U23281 (N_23281,N_17124,N_15209);
nand U23282 (N_23282,N_17076,N_18309);
nor U23283 (N_23283,N_18744,N_18339);
nor U23284 (N_23284,N_14217,N_15410);
or U23285 (N_23285,N_18065,N_13931);
xnor U23286 (N_23286,N_18274,N_15673);
nand U23287 (N_23287,N_13518,N_13770);
nor U23288 (N_23288,N_14339,N_18205);
nor U23289 (N_23289,N_14344,N_14336);
xnor U23290 (N_23290,N_17821,N_16935);
and U23291 (N_23291,N_12948,N_16974);
nand U23292 (N_23292,N_16539,N_13104);
xnor U23293 (N_23293,N_16722,N_13277);
and U23294 (N_23294,N_15278,N_12710);
or U23295 (N_23295,N_13146,N_16125);
xnor U23296 (N_23296,N_12809,N_13080);
nand U23297 (N_23297,N_17152,N_17238);
nor U23298 (N_23298,N_14002,N_18678);
and U23299 (N_23299,N_14500,N_17025);
nor U23300 (N_23300,N_16499,N_18396);
nand U23301 (N_23301,N_18122,N_17502);
and U23302 (N_23302,N_16585,N_18183);
nor U23303 (N_23303,N_16949,N_13458);
and U23304 (N_23304,N_17597,N_17866);
nor U23305 (N_23305,N_15152,N_14074);
xnor U23306 (N_23306,N_17631,N_16212);
xnor U23307 (N_23307,N_15857,N_17054);
or U23308 (N_23308,N_17842,N_15214);
nor U23309 (N_23309,N_16097,N_13398);
nand U23310 (N_23310,N_13483,N_18490);
nand U23311 (N_23311,N_14570,N_15859);
and U23312 (N_23312,N_13809,N_18225);
nand U23313 (N_23313,N_16978,N_15197);
xnor U23314 (N_23314,N_16992,N_12907);
and U23315 (N_23315,N_14187,N_17902);
xor U23316 (N_23316,N_17516,N_15373);
nand U23317 (N_23317,N_13177,N_18234);
or U23318 (N_23318,N_17769,N_13171);
and U23319 (N_23319,N_16432,N_17296);
and U23320 (N_23320,N_14565,N_17492);
or U23321 (N_23321,N_12890,N_17241);
or U23322 (N_23322,N_16975,N_17220);
nand U23323 (N_23323,N_12653,N_16946);
nor U23324 (N_23324,N_12854,N_12872);
nand U23325 (N_23325,N_18365,N_15690);
nor U23326 (N_23326,N_14172,N_16963);
and U23327 (N_23327,N_14386,N_18488);
nor U23328 (N_23328,N_17151,N_13775);
nor U23329 (N_23329,N_12808,N_13251);
xor U23330 (N_23330,N_13689,N_18182);
nor U23331 (N_23331,N_15686,N_13548);
nand U23332 (N_23332,N_18116,N_17591);
and U23333 (N_23333,N_16955,N_12554);
or U23334 (N_23334,N_17280,N_14915);
xor U23335 (N_23335,N_12662,N_18498);
and U23336 (N_23336,N_17371,N_16874);
nor U23337 (N_23337,N_18552,N_16321);
or U23338 (N_23338,N_14163,N_17062);
nor U23339 (N_23339,N_18323,N_16128);
and U23340 (N_23340,N_15839,N_17681);
xnor U23341 (N_23341,N_15859,N_16368);
and U23342 (N_23342,N_15684,N_13695);
and U23343 (N_23343,N_13055,N_15905);
or U23344 (N_23344,N_16384,N_16450);
nand U23345 (N_23345,N_16421,N_13893);
and U23346 (N_23346,N_14091,N_16435);
nor U23347 (N_23347,N_13404,N_14009);
or U23348 (N_23348,N_18655,N_13009);
and U23349 (N_23349,N_13152,N_16368);
nor U23350 (N_23350,N_15647,N_13798);
nor U23351 (N_23351,N_16594,N_17918);
nor U23352 (N_23352,N_17346,N_12648);
nor U23353 (N_23353,N_15531,N_13974);
or U23354 (N_23354,N_18518,N_12506);
or U23355 (N_23355,N_14230,N_16624);
nor U23356 (N_23356,N_15703,N_16524);
and U23357 (N_23357,N_15931,N_15121);
and U23358 (N_23358,N_16875,N_12978);
nor U23359 (N_23359,N_16737,N_17209);
xnor U23360 (N_23360,N_15476,N_12780);
nand U23361 (N_23361,N_18482,N_15232);
and U23362 (N_23362,N_15702,N_17029);
nor U23363 (N_23363,N_16570,N_15179);
and U23364 (N_23364,N_18246,N_14485);
xor U23365 (N_23365,N_13645,N_17573);
and U23366 (N_23366,N_12877,N_14836);
or U23367 (N_23367,N_12930,N_15088);
or U23368 (N_23368,N_12588,N_14408);
and U23369 (N_23369,N_16157,N_14840);
nand U23370 (N_23370,N_13595,N_16503);
xor U23371 (N_23371,N_16781,N_12663);
nor U23372 (N_23372,N_15162,N_15486);
xor U23373 (N_23373,N_14171,N_15754);
nand U23374 (N_23374,N_17836,N_13866);
nand U23375 (N_23375,N_12867,N_16735);
nand U23376 (N_23376,N_12694,N_18679);
and U23377 (N_23377,N_12518,N_13802);
or U23378 (N_23378,N_16248,N_14123);
xor U23379 (N_23379,N_16671,N_15718);
or U23380 (N_23380,N_16787,N_12874);
nand U23381 (N_23381,N_16658,N_12935);
or U23382 (N_23382,N_13622,N_17283);
nor U23383 (N_23383,N_12944,N_16417);
or U23384 (N_23384,N_17906,N_12665);
and U23385 (N_23385,N_14736,N_14103);
nand U23386 (N_23386,N_15117,N_13604);
xnor U23387 (N_23387,N_14899,N_17133);
nand U23388 (N_23388,N_14813,N_16262);
nand U23389 (N_23389,N_16245,N_12732);
xor U23390 (N_23390,N_15918,N_17559);
nand U23391 (N_23391,N_15520,N_16008);
nor U23392 (N_23392,N_15870,N_13447);
nand U23393 (N_23393,N_14026,N_18602);
or U23394 (N_23394,N_13621,N_15547);
nor U23395 (N_23395,N_17958,N_13308);
xnor U23396 (N_23396,N_14048,N_18483);
or U23397 (N_23397,N_17427,N_16021);
xnor U23398 (N_23398,N_12616,N_13807);
or U23399 (N_23399,N_17379,N_14859);
nor U23400 (N_23400,N_17021,N_18580);
or U23401 (N_23401,N_13725,N_16755);
and U23402 (N_23402,N_16300,N_18614);
nor U23403 (N_23403,N_15036,N_14548);
xnor U23404 (N_23404,N_15758,N_14952);
nor U23405 (N_23405,N_13497,N_15092);
xor U23406 (N_23406,N_13129,N_15010);
and U23407 (N_23407,N_13835,N_15505);
or U23408 (N_23408,N_14452,N_18399);
nand U23409 (N_23409,N_18235,N_14944);
nor U23410 (N_23410,N_15986,N_18215);
or U23411 (N_23411,N_16196,N_16600);
or U23412 (N_23412,N_16423,N_14873);
nand U23413 (N_23413,N_16589,N_12870);
and U23414 (N_23414,N_14231,N_17413);
xor U23415 (N_23415,N_13393,N_18643);
and U23416 (N_23416,N_13997,N_17117);
and U23417 (N_23417,N_18490,N_16923);
xor U23418 (N_23418,N_15252,N_14708);
xnor U23419 (N_23419,N_13583,N_17055);
or U23420 (N_23420,N_13047,N_13028);
and U23421 (N_23421,N_16279,N_15814);
xnor U23422 (N_23422,N_17871,N_14196);
nor U23423 (N_23423,N_18443,N_15671);
and U23424 (N_23424,N_14286,N_14410);
xnor U23425 (N_23425,N_14240,N_15920);
or U23426 (N_23426,N_16378,N_15471);
and U23427 (N_23427,N_16274,N_18574);
xnor U23428 (N_23428,N_16080,N_15736);
xor U23429 (N_23429,N_14663,N_12929);
nor U23430 (N_23430,N_15372,N_12829);
nor U23431 (N_23431,N_13361,N_16487);
and U23432 (N_23432,N_13266,N_15186);
nand U23433 (N_23433,N_16985,N_13151);
nand U23434 (N_23434,N_12503,N_16014);
nand U23435 (N_23435,N_16387,N_17789);
xnor U23436 (N_23436,N_16203,N_16855);
nor U23437 (N_23437,N_13924,N_13750);
and U23438 (N_23438,N_13305,N_14296);
xnor U23439 (N_23439,N_17301,N_13800);
xnor U23440 (N_23440,N_18689,N_16145);
xor U23441 (N_23441,N_18418,N_13224);
nand U23442 (N_23442,N_16415,N_16764);
and U23443 (N_23443,N_14997,N_18044);
and U23444 (N_23444,N_18721,N_18289);
and U23445 (N_23445,N_17822,N_14184);
nand U23446 (N_23446,N_16145,N_13980);
nand U23447 (N_23447,N_12990,N_15076);
nand U23448 (N_23448,N_15307,N_18512);
nand U23449 (N_23449,N_13217,N_16106);
or U23450 (N_23450,N_16090,N_17478);
and U23451 (N_23451,N_16247,N_17958);
and U23452 (N_23452,N_15599,N_17161);
nand U23453 (N_23453,N_18492,N_16024);
nand U23454 (N_23454,N_15185,N_17265);
nand U23455 (N_23455,N_18589,N_14834);
nand U23456 (N_23456,N_16668,N_17378);
xor U23457 (N_23457,N_17070,N_16598);
and U23458 (N_23458,N_16598,N_14997);
or U23459 (N_23459,N_14005,N_16759);
xnor U23460 (N_23460,N_17848,N_18379);
xor U23461 (N_23461,N_13221,N_12904);
or U23462 (N_23462,N_16715,N_13691);
nor U23463 (N_23463,N_13600,N_15675);
nor U23464 (N_23464,N_14670,N_15425);
nor U23465 (N_23465,N_16395,N_16783);
and U23466 (N_23466,N_13039,N_14676);
nor U23467 (N_23467,N_13632,N_17572);
nand U23468 (N_23468,N_16536,N_14503);
xnor U23469 (N_23469,N_16211,N_18192);
nand U23470 (N_23470,N_12959,N_12655);
nand U23471 (N_23471,N_13294,N_17704);
or U23472 (N_23472,N_15305,N_16959);
nor U23473 (N_23473,N_14162,N_13413);
or U23474 (N_23474,N_17319,N_16697);
and U23475 (N_23475,N_18307,N_14397);
or U23476 (N_23476,N_15782,N_14802);
or U23477 (N_23477,N_17194,N_17023);
or U23478 (N_23478,N_16040,N_16437);
xnor U23479 (N_23479,N_15115,N_13505);
and U23480 (N_23480,N_13718,N_17967);
or U23481 (N_23481,N_14613,N_15648);
nand U23482 (N_23482,N_12769,N_16105);
xnor U23483 (N_23483,N_14379,N_16042);
nor U23484 (N_23484,N_12796,N_17527);
xnor U23485 (N_23485,N_13446,N_12647);
and U23486 (N_23486,N_16866,N_16274);
and U23487 (N_23487,N_18317,N_18637);
and U23488 (N_23488,N_15521,N_16836);
or U23489 (N_23489,N_12728,N_18704);
nor U23490 (N_23490,N_15767,N_13901);
or U23491 (N_23491,N_13195,N_12835);
or U23492 (N_23492,N_18226,N_12654);
or U23493 (N_23493,N_16965,N_12806);
nor U23494 (N_23494,N_14174,N_18712);
and U23495 (N_23495,N_14218,N_16462);
and U23496 (N_23496,N_17941,N_15901);
nor U23497 (N_23497,N_13843,N_14671);
nand U23498 (N_23498,N_17272,N_12509);
or U23499 (N_23499,N_14060,N_18312);
and U23500 (N_23500,N_13782,N_15058);
xnor U23501 (N_23501,N_16386,N_16929);
nand U23502 (N_23502,N_14703,N_18485);
and U23503 (N_23503,N_14710,N_12746);
nor U23504 (N_23504,N_15465,N_16124);
and U23505 (N_23505,N_16289,N_12522);
nand U23506 (N_23506,N_13499,N_17848);
nand U23507 (N_23507,N_18378,N_14040);
nand U23508 (N_23508,N_14148,N_14625);
nand U23509 (N_23509,N_17925,N_17455);
nor U23510 (N_23510,N_15540,N_13239);
nor U23511 (N_23511,N_18285,N_17219);
nand U23512 (N_23512,N_17062,N_17638);
nand U23513 (N_23513,N_14111,N_18687);
or U23514 (N_23514,N_14285,N_12905);
or U23515 (N_23515,N_15741,N_12528);
or U23516 (N_23516,N_12913,N_13576);
nand U23517 (N_23517,N_15101,N_16922);
nand U23518 (N_23518,N_14435,N_12645);
nand U23519 (N_23519,N_17256,N_13162);
or U23520 (N_23520,N_14831,N_12866);
or U23521 (N_23521,N_13401,N_13744);
nand U23522 (N_23522,N_17589,N_12754);
nand U23523 (N_23523,N_16831,N_13953);
nand U23524 (N_23524,N_14515,N_17589);
xnor U23525 (N_23525,N_14589,N_15316);
or U23526 (N_23526,N_13012,N_18450);
or U23527 (N_23527,N_16005,N_18292);
nand U23528 (N_23528,N_17122,N_15043);
nand U23529 (N_23529,N_17527,N_12974);
nor U23530 (N_23530,N_12724,N_14345);
nand U23531 (N_23531,N_17295,N_14568);
nand U23532 (N_23532,N_15749,N_18266);
or U23533 (N_23533,N_17037,N_14521);
and U23534 (N_23534,N_14275,N_13357);
and U23535 (N_23535,N_13422,N_15150);
nor U23536 (N_23536,N_17682,N_12947);
or U23537 (N_23537,N_13160,N_16624);
xor U23538 (N_23538,N_12775,N_16413);
or U23539 (N_23539,N_14544,N_18536);
nand U23540 (N_23540,N_18132,N_15702);
or U23541 (N_23541,N_13323,N_15485);
nor U23542 (N_23542,N_18187,N_16465);
nand U23543 (N_23543,N_18743,N_18616);
and U23544 (N_23544,N_17448,N_13754);
and U23545 (N_23545,N_15877,N_15271);
nand U23546 (N_23546,N_12683,N_18400);
and U23547 (N_23547,N_13364,N_17348);
or U23548 (N_23548,N_16882,N_16950);
nor U23549 (N_23549,N_12775,N_15371);
and U23550 (N_23550,N_14158,N_15377);
or U23551 (N_23551,N_16595,N_14409);
or U23552 (N_23552,N_13299,N_15358);
and U23553 (N_23553,N_13295,N_18715);
nor U23554 (N_23554,N_13694,N_14441);
and U23555 (N_23555,N_14634,N_14674);
or U23556 (N_23556,N_15263,N_15603);
and U23557 (N_23557,N_13643,N_14367);
nand U23558 (N_23558,N_15289,N_16843);
nand U23559 (N_23559,N_17970,N_13343);
xnor U23560 (N_23560,N_14203,N_14144);
and U23561 (N_23561,N_18061,N_13526);
xnor U23562 (N_23562,N_16280,N_16333);
and U23563 (N_23563,N_14689,N_18702);
xnor U23564 (N_23564,N_13404,N_14486);
nand U23565 (N_23565,N_14239,N_18405);
nand U23566 (N_23566,N_18464,N_16635);
xnor U23567 (N_23567,N_14071,N_17121);
nand U23568 (N_23568,N_16015,N_14439);
and U23569 (N_23569,N_14127,N_14039);
or U23570 (N_23570,N_15471,N_13853);
nor U23571 (N_23571,N_15879,N_15950);
xor U23572 (N_23572,N_18225,N_14454);
nand U23573 (N_23573,N_13851,N_16908);
nor U23574 (N_23574,N_18646,N_12766);
nor U23575 (N_23575,N_18001,N_15180);
and U23576 (N_23576,N_15594,N_14825);
xor U23577 (N_23577,N_14461,N_16294);
nor U23578 (N_23578,N_15114,N_15820);
xor U23579 (N_23579,N_17236,N_14396);
xor U23580 (N_23580,N_16506,N_16220);
xnor U23581 (N_23581,N_17601,N_16389);
nand U23582 (N_23582,N_17585,N_18392);
nor U23583 (N_23583,N_15196,N_15982);
or U23584 (N_23584,N_13218,N_17887);
or U23585 (N_23585,N_15131,N_16338);
nand U23586 (N_23586,N_16555,N_12694);
or U23587 (N_23587,N_17459,N_14409);
and U23588 (N_23588,N_16818,N_13280);
and U23589 (N_23589,N_16515,N_17633);
or U23590 (N_23590,N_13520,N_18643);
and U23591 (N_23591,N_16240,N_15502);
xnor U23592 (N_23592,N_12787,N_17770);
nor U23593 (N_23593,N_15645,N_17372);
nand U23594 (N_23594,N_16878,N_15082);
or U23595 (N_23595,N_14327,N_18159);
and U23596 (N_23596,N_16807,N_17152);
xor U23597 (N_23597,N_17197,N_14887);
or U23598 (N_23598,N_17399,N_15014);
and U23599 (N_23599,N_18266,N_14253);
or U23600 (N_23600,N_16244,N_16952);
xnor U23601 (N_23601,N_13981,N_15037);
nand U23602 (N_23602,N_14963,N_15914);
xor U23603 (N_23603,N_15347,N_17808);
xor U23604 (N_23604,N_16161,N_17087);
nor U23605 (N_23605,N_12793,N_13244);
and U23606 (N_23606,N_16370,N_13243);
xor U23607 (N_23607,N_15079,N_12879);
nand U23608 (N_23608,N_16014,N_18324);
and U23609 (N_23609,N_15834,N_14736);
and U23610 (N_23610,N_12568,N_14976);
nand U23611 (N_23611,N_15477,N_16325);
xor U23612 (N_23612,N_14632,N_13751);
and U23613 (N_23613,N_16598,N_13384);
xnor U23614 (N_23614,N_14579,N_17739);
nand U23615 (N_23615,N_16387,N_13148);
xnor U23616 (N_23616,N_14222,N_17961);
or U23617 (N_23617,N_15606,N_17764);
or U23618 (N_23618,N_13944,N_18736);
and U23619 (N_23619,N_16314,N_14626);
nand U23620 (N_23620,N_13501,N_13548);
nor U23621 (N_23621,N_16004,N_17623);
nor U23622 (N_23622,N_15564,N_13336);
nor U23623 (N_23623,N_16366,N_16550);
xor U23624 (N_23624,N_18587,N_17306);
or U23625 (N_23625,N_15867,N_13968);
xor U23626 (N_23626,N_15155,N_15006);
xor U23627 (N_23627,N_18057,N_17760);
nand U23628 (N_23628,N_17110,N_16777);
nor U23629 (N_23629,N_14211,N_16296);
nor U23630 (N_23630,N_18617,N_13474);
nand U23631 (N_23631,N_12678,N_17493);
xor U23632 (N_23632,N_15644,N_18425);
or U23633 (N_23633,N_15282,N_14929);
and U23634 (N_23634,N_18652,N_17706);
nor U23635 (N_23635,N_17614,N_16333);
xor U23636 (N_23636,N_18199,N_15458);
nor U23637 (N_23637,N_15228,N_12997);
or U23638 (N_23638,N_14140,N_14253);
nand U23639 (N_23639,N_14374,N_14255);
or U23640 (N_23640,N_16628,N_15916);
or U23641 (N_23641,N_15369,N_14980);
nor U23642 (N_23642,N_13559,N_14310);
or U23643 (N_23643,N_13696,N_14102);
and U23644 (N_23644,N_14554,N_18536);
or U23645 (N_23645,N_12523,N_13072);
xnor U23646 (N_23646,N_15490,N_13297);
and U23647 (N_23647,N_17693,N_16613);
or U23648 (N_23648,N_17892,N_18391);
and U23649 (N_23649,N_16263,N_13806);
and U23650 (N_23650,N_18436,N_18273);
nand U23651 (N_23651,N_13682,N_15991);
or U23652 (N_23652,N_17527,N_16245);
nand U23653 (N_23653,N_14474,N_16386);
nor U23654 (N_23654,N_12932,N_12711);
or U23655 (N_23655,N_17689,N_18423);
nand U23656 (N_23656,N_18072,N_17753);
nand U23657 (N_23657,N_12995,N_16432);
nand U23658 (N_23658,N_13535,N_17327);
and U23659 (N_23659,N_12563,N_14841);
xor U23660 (N_23660,N_16383,N_15817);
xor U23661 (N_23661,N_17389,N_13579);
or U23662 (N_23662,N_13129,N_18565);
or U23663 (N_23663,N_13802,N_13470);
and U23664 (N_23664,N_17568,N_12557);
nor U23665 (N_23665,N_18029,N_17934);
nor U23666 (N_23666,N_13673,N_16945);
nand U23667 (N_23667,N_14583,N_14661);
or U23668 (N_23668,N_13530,N_16950);
or U23669 (N_23669,N_17715,N_12917);
xnor U23670 (N_23670,N_14699,N_14334);
nand U23671 (N_23671,N_14942,N_15579);
xor U23672 (N_23672,N_16913,N_17058);
xnor U23673 (N_23673,N_16964,N_17418);
nor U23674 (N_23674,N_16208,N_16356);
xor U23675 (N_23675,N_17233,N_15439);
nor U23676 (N_23676,N_18160,N_17298);
nor U23677 (N_23677,N_13729,N_12703);
nor U23678 (N_23678,N_13480,N_13710);
and U23679 (N_23679,N_13061,N_14242);
nand U23680 (N_23680,N_12701,N_13887);
nor U23681 (N_23681,N_17642,N_14184);
xnor U23682 (N_23682,N_16111,N_15709);
or U23683 (N_23683,N_13535,N_14753);
nand U23684 (N_23684,N_17894,N_17838);
xnor U23685 (N_23685,N_18162,N_13829);
nand U23686 (N_23686,N_16349,N_14580);
nor U23687 (N_23687,N_17114,N_15733);
nor U23688 (N_23688,N_16528,N_15857);
or U23689 (N_23689,N_13034,N_13315);
or U23690 (N_23690,N_15397,N_17597);
and U23691 (N_23691,N_17908,N_13008);
or U23692 (N_23692,N_17832,N_13984);
nand U23693 (N_23693,N_13475,N_16599);
nor U23694 (N_23694,N_15094,N_15401);
nand U23695 (N_23695,N_15663,N_14263);
and U23696 (N_23696,N_12695,N_13557);
xor U23697 (N_23697,N_13710,N_17701);
nor U23698 (N_23698,N_18452,N_16237);
nor U23699 (N_23699,N_18471,N_18443);
or U23700 (N_23700,N_17136,N_18641);
or U23701 (N_23701,N_17858,N_15207);
nor U23702 (N_23702,N_17660,N_17630);
or U23703 (N_23703,N_14766,N_13393);
and U23704 (N_23704,N_14052,N_12873);
xor U23705 (N_23705,N_12608,N_13743);
nand U23706 (N_23706,N_16294,N_15608);
nand U23707 (N_23707,N_17239,N_13481);
nand U23708 (N_23708,N_15051,N_14708);
nor U23709 (N_23709,N_18171,N_18388);
xnor U23710 (N_23710,N_16535,N_16861);
xor U23711 (N_23711,N_17967,N_14576);
and U23712 (N_23712,N_17451,N_18606);
nand U23713 (N_23713,N_13612,N_18422);
and U23714 (N_23714,N_13839,N_13309);
nand U23715 (N_23715,N_18102,N_13252);
and U23716 (N_23716,N_17671,N_17835);
or U23717 (N_23717,N_14153,N_15607);
xnor U23718 (N_23718,N_17194,N_16847);
nand U23719 (N_23719,N_13247,N_13554);
nor U23720 (N_23720,N_15816,N_17660);
and U23721 (N_23721,N_16470,N_13372);
xor U23722 (N_23722,N_16465,N_13343);
nor U23723 (N_23723,N_14317,N_13881);
nor U23724 (N_23724,N_18160,N_13562);
or U23725 (N_23725,N_15784,N_17756);
and U23726 (N_23726,N_17867,N_17903);
xnor U23727 (N_23727,N_13297,N_16445);
xor U23728 (N_23728,N_15083,N_12875);
nor U23729 (N_23729,N_15711,N_15104);
nor U23730 (N_23730,N_13733,N_15239);
and U23731 (N_23731,N_15715,N_13454);
and U23732 (N_23732,N_16352,N_13429);
xnor U23733 (N_23733,N_13829,N_16272);
or U23734 (N_23734,N_13106,N_17240);
nand U23735 (N_23735,N_14964,N_18563);
and U23736 (N_23736,N_15938,N_12909);
or U23737 (N_23737,N_16664,N_16668);
and U23738 (N_23738,N_14412,N_18510);
and U23739 (N_23739,N_17292,N_13926);
xor U23740 (N_23740,N_15953,N_17879);
or U23741 (N_23741,N_17586,N_17109);
nor U23742 (N_23742,N_18636,N_15644);
xnor U23743 (N_23743,N_14847,N_14902);
xor U23744 (N_23744,N_14276,N_18723);
xor U23745 (N_23745,N_17707,N_12902);
or U23746 (N_23746,N_13147,N_14165);
and U23747 (N_23747,N_15621,N_14655);
xor U23748 (N_23748,N_17148,N_13950);
nand U23749 (N_23749,N_14956,N_14523);
nor U23750 (N_23750,N_18428,N_13203);
nor U23751 (N_23751,N_13894,N_16724);
or U23752 (N_23752,N_13377,N_17300);
nand U23753 (N_23753,N_15590,N_18329);
nor U23754 (N_23754,N_18732,N_14264);
or U23755 (N_23755,N_17613,N_16610);
and U23756 (N_23756,N_17999,N_17024);
or U23757 (N_23757,N_15707,N_16964);
nor U23758 (N_23758,N_12804,N_17167);
nor U23759 (N_23759,N_14555,N_14901);
nor U23760 (N_23760,N_14651,N_17816);
or U23761 (N_23761,N_18626,N_12758);
xnor U23762 (N_23762,N_15358,N_13368);
or U23763 (N_23763,N_13026,N_12741);
or U23764 (N_23764,N_14889,N_15896);
nand U23765 (N_23765,N_13781,N_16520);
xnor U23766 (N_23766,N_13669,N_17850);
xor U23767 (N_23767,N_13996,N_18000);
xnor U23768 (N_23768,N_18278,N_15498);
nand U23769 (N_23769,N_13817,N_17177);
nand U23770 (N_23770,N_15092,N_17898);
xor U23771 (N_23771,N_14381,N_12517);
xor U23772 (N_23772,N_17987,N_14795);
or U23773 (N_23773,N_13378,N_15010);
nor U23774 (N_23774,N_14024,N_14402);
nor U23775 (N_23775,N_17403,N_16546);
nor U23776 (N_23776,N_16176,N_14807);
and U23777 (N_23777,N_14534,N_18297);
or U23778 (N_23778,N_15632,N_12791);
or U23779 (N_23779,N_14684,N_17088);
xor U23780 (N_23780,N_15854,N_17723);
nand U23781 (N_23781,N_14880,N_13790);
nor U23782 (N_23782,N_16171,N_14626);
nand U23783 (N_23783,N_13602,N_15385);
xnor U23784 (N_23784,N_14906,N_17743);
and U23785 (N_23785,N_15187,N_12877);
nor U23786 (N_23786,N_12578,N_13378);
nand U23787 (N_23787,N_17276,N_16383);
xor U23788 (N_23788,N_15179,N_14596);
or U23789 (N_23789,N_15580,N_18659);
nor U23790 (N_23790,N_13805,N_15181);
and U23791 (N_23791,N_16210,N_17194);
nor U23792 (N_23792,N_18495,N_13557);
nand U23793 (N_23793,N_18728,N_14587);
nor U23794 (N_23794,N_18460,N_15544);
nor U23795 (N_23795,N_15411,N_15868);
or U23796 (N_23796,N_18582,N_15905);
nand U23797 (N_23797,N_17662,N_16174);
and U23798 (N_23798,N_15130,N_15236);
and U23799 (N_23799,N_18200,N_14262);
and U23800 (N_23800,N_13869,N_18266);
nand U23801 (N_23801,N_15177,N_15381);
nor U23802 (N_23802,N_15623,N_13449);
nand U23803 (N_23803,N_18073,N_14680);
or U23804 (N_23804,N_14765,N_18018);
xnor U23805 (N_23805,N_17748,N_14355);
xnor U23806 (N_23806,N_12598,N_15164);
nor U23807 (N_23807,N_17632,N_16436);
nor U23808 (N_23808,N_16673,N_16777);
xnor U23809 (N_23809,N_16047,N_14580);
xor U23810 (N_23810,N_13285,N_17730);
or U23811 (N_23811,N_17206,N_16636);
nand U23812 (N_23812,N_16161,N_18186);
nand U23813 (N_23813,N_17626,N_14516);
xor U23814 (N_23814,N_13322,N_14372);
xnor U23815 (N_23815,N_18438,N_14414);
nor U23816 (N_23816,N_17051,N_13394);
and U23817 (N_23817,N_18570,N_18096);
xnor U23818 (N_23818,N_13920,N_16504);
nor U23819 (N_23819,N_17917,N_13470);
nand U23820 (N_23820,N_12836,N_13443);
xnor U23821 (N_23821,N_13340,N_18093);
and U23822 (N_23822,N_14593,N_14440);
nand U23823 (N_23823,N_17668,N_16081);
or U23824 (N_23824,N_18414,N_15072);
nor U23825 (N_23825,N_14604,N_15865);
nand U23826 (N_23826,N_18336,N_15966);
nand U23827 (N_23827,N_17733,N_17839);
nor U23828 (N_23828,N_14232,N_14066);
xor U23829 (N_23829,N_15350,N_17820);
and U23830 (N_23830,N_13184,N_13705);
or U23831 (N_23831,N_12594,N_15910);
nand U23832 (N_23832,N_17522,N_14147);
nor U23833 (N_23833,N_16559,N_12614);
and U23834 (N_23834,N_15141,N_14026);
nand U23835 (N_23835,N_15351,N_17254);
nand U23836 (N_23836,N_12605,N_15032);
or U23837 (N_23837,N_16484,N_14338);
and U23838 (N_23838,N_14733,N_18563);
or U23839 (N_23839,N_16447,N_16124);
xnor U23840 (N_23840,N_17337,N_14550);
xor U23841 (N_23841,N_12609,N_17098);
or U23842 (N_23842,N_15561,N_14384);
and U23843 (N_23843,N_15810,N_14723);
nor U23844 (N_23844,N_14227,N_17355);
xor U23845 (N_23845,N_18444,N_14437);
or U23846 (N_23846,N_18085,N_15502);
xor U23847 (N_23847,N_14902,N_18654);
and U23848 (N_23848,N_16554,N_14011);
nand U23849 (N_23849,N_13849,N_18666);
or U23850 (N_23850,N_14053,N_12786);
nand U23851 (N_23851,N_14253,N_15742);
nand U23852 (N_23852,N_17272,N_17198);
nor U23853 (N_23853,N_14954,N_16336);
nand U23854 (N_23854,N_17542,N_17129);
and U23855 (N_23855,N_12506,N_15502);
nand U23856 (N_23856,N_15967,N_17416);
or U23857 (N_23857,N_15928,N_17493);
xnor U23858 (N_23858,N_14161,N_16047);
nor U23859 (N_23859,N_16755,N_14726);
or U23860 (N_23860,N_16797,N_13543);
nor U23861 (N_23861,N_18200,N_12842);
or U23862 (N_23862,N_13855,N_14980);
or U23863 (N_23863,N_17568,N_18018);
nor U23864 (N_23864,N_18312,N_13191);
nor U23865 (N_23865,N_14866,N_15901);
xnor U23866 (N_23866,N_16698,N_15502);
nor U23867 (N_23867,N_16278,N_13494);
or U23868 (N_23868,N_13594,N_17883);
nor U23869 (N_23869,N_17212,N_12848);
or U23870 (N_23870,N_18344,N_14783);
nand U23871 (N_23871,N_15737,N_18485);
nand U23872 (N_23872,N_13086,N_14535);
or U23873 (N_23873,N_15502,N_15872);
xor U23874 (N_23874,N_15429,N_18637);
nor U23875 (N_23875,N_17208,N_16876);
or U23876 (N_23876,N_14510,N_18657);
nor U23877 (N_23877,N_16271,N_13970);
or U23878 (N_23878,N_14765,N_14251);
xnor U23879 (N_23879,N_15128,N_15512);
nor U23880 (N_23880,N_16100,N_14933);
and U23881 (N_23881,N_18341,N_13536);
and U23882 (N_23882,N_13704,N_16757);
nand U23883 (N_23883,N_13278,N_18662);
xor U23884 (N_23884,N_17259,N_14399);
nand U23885 (N_23885,N_17737,N_15083);
nor U23886 (N_23886,N_16204,N_16845);
nor U23887 (N_23887,N_13858,N_18545);
nor U23888 (N_23888,N_15517,N_14209);
or U23889 (N_23889,N_15737,N_14137);
or U23890 (N_23890,N_15675,N_17210);
and U23891 (N_23891,N_12757,N_14373);
nor U23892 (N_23892,N_16132,N_16432);
nor U23893 (N_23893,N_13392,N_17947);
nand U23894 (N_23894,N_16136,N_15633);
or U23895 (N_23895,N_13988,N_15053);
xor U23896 (N_23896,N_15226,N_14810);
and U23897 (N_23897,N_13005,N_13084);
nor U23898 (N_23898,N_14886,N_14239);
xor U23899 (N_23899,N_15127,N_13481);
or U23900 (N_23900,N_15349,N_13857);
nor U23901 (N_23901,N_15415,N_12695);
nand U23902 (N_23902,N_16717,N_18037);
or U23903 (N_23903,N_15223,N_16894);
nand U23904 (N_23904,N_14678,N_18177);
nand U23905 (N_23905,N_16584,N_15624);
nand U23906 (N_23906,N_16067,N_14137);
xnor U23907 (N_23907,N_14172,N_12926);
nor U23908 (N_23908,N_16426,N_17434);
nand U23909 (N_23909,N_14709,N_17831);
and U23910 (N_23910,N_13604,N_13206);
nor U23911 (N_23911,N_18118,N_16423);
xor U23912 (N_23912,N_13993,N_15712);
nand U23913 (N_23913,N_14207,N_14304);
nand U23914 (N_23914,N_15209,N_16537);
xnor U23915 (N_23915,N_13370,N_16824);
xnor U23916 (N_23916,N_17914,N_14300);
and U23917 (N_23917,N_12745,N_15575);
nor U23918 (N_23918,N_13582,N_16815);
nor U23919 (N_23919,N_18174,N_17282);
nand U23920 (N_23920,N_16244,N_14474);
or U23921 (N_23921,N_15611,N_14008);
nand U23922 (N_23922,N_15860,N_17974);
nand U23923 (N_23923,N_13469,N_15953);
xor U23924 (N_23924,N_14423,N_15152);
nor U23925 (N_23925,N_14385,N_16372);
xnor U23926 (N_23926,N_14423,N_15998);
nand U23927 (N_23927,N_15398,N_18700);
nor U23928 (N_23928,N_17640,N_17406);
and U23929 (N_23929,N_17550,N_18586);
nor U23930 (N_23930,N_15067,N_18690);
and U23931 (N_23931,N_18723,N_16765);
xnor U23932 (N_23932,N_12938,N_15309);
nor U23933 (N_23933,N_14736,N_14563);
or U23934 (N_23934,N_13943,N_17297);
nand U23935 (N_23935,N_18196,N_13630);
or U23936 (N_23936,N_13864,N_14365);
nand U23937 (N_23937,N_15332,N_18177);
nand U23938 (N_23938,N_17267,N_18402);
or U23939 (N_23939,N_13237,N_18120);
xnor U23940 (N_23940,N_14558,N_14877);
or U23941 (N_23941,N_17183,N_14561);
nand U23942 (N_23942,N_17741,N_15896);
and U23943 (N_23943,N_16154,N_16021);
xnor U23944 (N_23944,N_13591,N_14843);
nor U23945 (N_23945,N_15402,N_17853);
nor U23946 (N_23946,N_14279,N_17350);
or U23947 (N_23947,N_15174,N_16395);
nand U23948 (N_23948,N_17346,N_17689);
and U23949 (N_23949,N_14639,N_16778);
nor U23950 (N_23950,N_18357,N_16131);
nand U23951 (N_23951,N_15921,N_16733);
or U23952 (N_23952,N_15281,N_12917);
nand U23953 (N_23953,N_17876,N_13162);
and U23954 (N_23954,N_18012,N_18330);
or U23955 (N_23955,N_15165,N_15229);
xnor U23956 (N_23956,N_13732,N_17106);
or U23957 (N_23957,N_14242,N_15220);
xor U23958 (N_23958,N_17431,N_17399);
and U23959 (N_23959,N_16675,N_17571);
nor U23960 (N_23960,N_16265,N_14542);
or U23961 (N_23961,N_15405,N_13039);
or U23962 (N_23962,N_13566,N_14283);
nor U23963 (N_23963,N_12768,N_17856);
or U23964 (N_23964,N_14136,N_17777);
nand U23965 (N_23965,N_18253,N_12898);
xor U23966 (N_23966,N_16549,N_12897);
or U23967 (N_23967,N_17019,N_15304);
nor U23968 (N_23968,N_12767,N_16178);
and U23969 (N_23969,N_17151,N_15825);
and U23970 (N_23970,N_13494,N_15100);
or U23971 (N_23971,N_15553,N_13609);
xor U23972 (N_23972,N_16566,N_12745);
nor U23973 (N_23973,N_14532,N_13935);
nand U23974 (N_23974,N_14104,N_13896);
nand U23975 (N_23975,N_14942,N_14179);
xnor U23976 (N_23976,N_15176,N_16418);
or U23977 (N_23977,N_17799,N_14229);
or U23978 (N_23978,N_18741,N_14117);
and U23979 (N_23979,N_18657,N_13713);
or U23980 (N_23980,N_16931,N_17363);
nor U23981 (N_23981,N_15162,N_18494);
xor U23982 (N_23982,N_16082,N_13501);
or U23983 (N_23983,N_15978,N_14254);
and U23984 (N_23984,N_18360,N_13271);
nand U23985 (N_23985,N_18264,N_13949);
and U23986 (N_23986,N_16094,N_13459);
nand U23987 (N_23987,N_13582,N_14221);
or U23988 (N_23988,N_15913,N_14936);
xor U23989 (N_23989,N_17567,N_14453);
nand U23990 (N_23990,N_17411,N_14364);
xnor U23991 (N_23991,N_15127,N_16154);
and U23992 (N_23992,N_15693,N_17178);
nor U23993 (N_23993,N_16976,N_12517);
or U23994 (N_23994,N_16354,N_15281);
nand U23995 (N_23995,N_12753,N_18125);
nand U23996 (N_23996,N_16502,N_14026);
or U23997 (N_23997,N_13124,N_15107);
nand U23998 (N_23998,N_15178,N_17911);
and U23999 (N_23999,N_16924,N_13080);
nand U24000 (N_24000,N_15269,N_18116);
nor U24001 (N_24001,N_13105,N_12923);
xor U24002 (N_24002,N_12519,N_17736);
and U24003 (N_24003,N_15181,N_15001);
nand U24004 (N_24004,N_12619,N_15073);
and U24005 (N_24005,N_15225,N_17108);
nor U24006 (N_24006,N_16312,N_18442);
or U24007 (N_24007,N_17742,N_18491);
xnor U24008 (N_24008,N_15175,N_12514);
nor U24009 (N_24009,N_14446,N_18242);
xor U24010 (N_24010,N_15272,N_12773);
xor U24011 (N_24011,N_14548,N_16463);
xor U24012 (N_24012,N_17014,N_14621);
and U24013 (N_24013,N_17910,N_16397);
and U24014 (N_24014,N_15173,N_14120);
nand U24015 (N_24015,N_17462,N_18565);
nor U24016 (N_24016,N_12829,N_15065);
nand U24017 (N_24017,N_16360,N_18606);
or U24018 (N_24018,N_15726,N_15766);
xor U24019 (N_24019,N_13584,N_13322);
and U24020 (N_24020,N_17827,N_17160);
nor U24021 (N_24021,N_16828,N_17134);
or U24022 (N_24022,N_14369,N_12953);
or U24023 (N_24023,N_18270,N_12633);
and U24024 (N_24024,N_13498,N_13878);
xor U24025 (N_24025,N_12540,N_15063);
and U24026 (N_24026,N_14055,N_14948);
xor U24027 (N_24027,N_13205,N_16477);
nand U24028 (N_24028,N_15330,N_17731);
xnor U24029 (N_24029,N_16935,N_13366);
nand U24030 (N_24030,N_15531,N_18374);
nand U24031 (N_24031,N_17832,N_18006);
or U24032 (N_24032,N_15748,N_14811);
or U24033 (N_24033,N_18223,N_13375);
xor U24034 (N_24034,N_17240,N_14725);
and U24035 (N_24035,N_13500,N_13040);
nor U24036 (N_24036,N_18402,N_18020);
nor U24037 (N_24037,N_16033,N_17224);
nand U24038 (N_24038,N_14211,N_16342);
and U24039 (N_24039,N_18019,N_14237);
nand U24040 (N_24040,N_13039,N_18147);
or U24041 (N_24041,N_13654,N_16751);
and U24042 (N_24042,N_13123,N_13726);
nand U24043 (N_24043,N_14179,N_17957);
nand U24044 (N_24044,N_15826,N_13279);
nor U24045 (N_24045,N_14508,N_16979);
nand U24046 (N_24046,N_17745,N_18196);
xnor U24047 (N_24047,N_17357,N_16033);
or U24048 (N_24048,N_16619,N_15601);
or U24049 (N_24049,N_15754,N_16609);
and U24050 (N_24050,N_15115,N_15578);
xor U24051 (N_24051,N_14773,N_18482);
nand U24052 (N_24052,N_15126,N_17634);
or U24053 (N_24053,N_12613,N_13400);
xnor U24054 (N_24054,N_16081,N_12873);
and U24055 (N_24055,N_13605,N_14646);
nor U24056 (N_24056,N_14640,N_15281);
nand U24057 (N_24057,N_17453,N_14102);
xor U24058 (N_24058,N_14877,N_14705);
nor U24059 (N_24059,N_18535,N_15480);
and U24060 (N_24060,N_13009,N_16771);
xor U24061 (N_24061,N_16862,N_15922);
xor U24062 (N_24062,N_17940,N_17115);
or U24063 (N_24063,N_15481,N_16628);
xnor U24064 (N_24064,N_14747,N_13003);
xor U24065 (N_24065,N_14484,N_15810);
nand U24066 (N_24066,N_15173,N_14381);
nor U24067 (N_24067,N_15182,N_17100);
nand U24068 (N_24068,N_14629,N_17755);
nand U24069 (N_24069,N_12983,N_14104);
nand U24070 (N_24070,N_14502,N_13543);
nor U24071 (N_24071,N_18609,N_13011);
or U24072 (N_24072,N_16903,N_17940);
nand U24073 (N_24073,N_13693,N_12632);
and U24074 (N_24074,N_16785,N_14765);
and U24075 (N_24075,N_18689,N_18513);
xnor U24076 (N_24076,N_18044,N_14491);
and U24077 (N_24077,N_16289,N_15167);
nand U24078 (N_24078,N_14477,N_18236);
and U24079 (N_24079,N_15602,N_18642);
or U24080 (N_24080,N_15345,N_12957);
xor U24081 (N_24081,N_18542,N_15410);
nand U24082 (N_24082,N_15121,N_13279);
or U24083 (N_24083,N_16596,N_15983);
and U24084 (N_24084,N_14135,N_14431);
nor U24085 (N_24085,N_17401,N_18583);
nand U24086 (N_24086,N_16721,N_18229);
nand U24087 (N_24087,N_18671,N_13832);
and U24088 (N_24088,N_16004,N_17409);
xor U24089 (N_24089,N_14904,N_15844);
or U24090 (N_24090,N_15848,N_14136);
or U24091 (N_24091,N_14266,N_17444);
nand U24092 (N_24092,N_13131,N_14971);
xnor U24093 (N_24093,N_13474,N_16930);
and U24094 (N_24094,N_15755,N_16370);
nor U24095 (N_24095,N_18075,N_16640);
xor U24096 (N_24096,N_16421,N_18019);
nor U24097 (N_24097,N_16062,N_14791);
or U24098 (N_24098,N_18616,N_12922);
nor U24099 (N_24099,N_18049,N_18611);
nor U24100 (N_24100,N_13116,N_17102);
xnor U24101 (N_24101,N_13820,N_13390);
and U24102 (N_24102,N_15737,N_15399);
nor U24103 (N_24103,N_14548,N_14917);
xnor U24104 (N_24104,N_16239,N_15928);
nor U24105 (N_24105,N_13389,N_16041);
or U24106 (N_24106,N_14915,N_15569);
or U24107 (N_24107,N_15115,N_17482);
nand U24108 (N_24108,N_17476,N_12829);
xor U24109 (N_24109,N_17429,N_12677);
xor U24110 (N_24110,N_18439,N_13393);
or U24111 (N_24111,N_13904,N_13814);
and U24112 (N_24112,N_15760,N_12986);
and U24113 (N_24113,N_15986,N_14907);
nand U24114 (N_24114,N_13806,N_16723);
or U24115 (N_24115,N_17103,N_16947);
nand U24116 (N_24116,N_17688,N_17603);
or U24117 (N_24117,N_17147,N_16877);
xor U24118 (N_24118,N_12974,N_17741);
and U24119 (N_24119,N_16277,N_14061);
nand U24120 (N_24120,N_18174,N_15684);
nand U24121 (N_24121,N_16430,N_18634);
and U24122 (N_24122,N_17533,N_14889);
xor U24123 (N_24123,N_14226,N_12850);
and U24124 (N_24124,N_13111,N_13146);
nor U24125 (N_24125,N_15379,N_17672);
or U24126 (N_24126,N_15533,N_16590);
xnor U24127 (N_24127,N_12768,N_15742);
nor U24128 (N_24128,N_13922,N_14432);
or U24129 (N_24129,N_13199,N_16512);
or U24130 (N_24130,N_12532,N_17950);
nand U24131 (N_24131,N_13717,N_15926);
or U24132 (N_24132,N_18092,N_15393);
nand U24133 (N_24133,N_13056,N_16065);
nor U24134 (N_24134,N_18563,N_18396);
nand U24135 (N_24135,N_16950,N_13962);
or U24136 (N_24136,N_14209,N_17974);
nor U24137 (N_24137,N_18747,N_14231);
xor U24138 (N_24138,N_16684,N_17919);
or U24139 (N_24139,N_16406,N_15862);
xnor U24140 (N_24140,N_13972,N_12631);
xnor U24141 (N_24141,N_13654,N_15694);
or U24142 (N_24142,N_13092,N_16954);
and U24143 (N_24143,N_14098,N_13339);
and U24144 (N_24144,N_16110,N_13914);
or U24145 (N_24145,N_15464,N_16371);
and U24146 (N_24146,N_15303,N_13261);
and U24147 (N_24147,N_12912,N_14476);
nor U24148 (N_24148,N_15250,N_18327);
nand U24149 (N_24149,N_16616,N_14576);
and U24150 (N_24150,N_15797,N_16604);
or U24151 (N_24151,N_16244,N_17829);
or U24152 (N_24152,N_17044,N_14397);
nor U24153 (N_24153,N_15152,N_14903);
and U24154 (N_24154,N_12777,N_17954);
xor U24155 (N_24155,N_12744,N_12545);
nand U24156 (N_24156,N_14319,N_18674);
nand U24157 (N_24157,N_13935,N_13959);
and U24158 (N_24158,N_12970,N_15278);
nand U24159 (N_24159,N_17044,N_15357);
nand U24160 (N_24160,N_13388,N_16865);
xnor U24161 (N_24161,N_18600,N_13699);
nor U24162 (N_24162,N_18581,N_16809);
nor U24163 (N_24163,N_16209,N_18280);
xor U24164 (N_24164,N_14872,N_17371);
nand U24165 (N_24165,N_14758,N_12853);
and U24166 (N_24166,N_16663,N_14851);
xnor U24167 (N_24167,N_16863,N_17408);
xnor U24168 (N_24168,N_15595,N_13576);
nand U24169 (N_24169,N_13590,N_16643);
nor U24170 (N_24170,N_16381,N_12873);
nand U24171 (N_24171,N_16954,N_13119);
nand U24172 (N_24172,N_17602,N_14199);
nand U24173 (N_24173,N_17970,N_18074);
or U24174 (N_24174,N_12828,N_14897);
or U24175 (N_24175,N_17634,N_12518);
nand U24176 (N_24176,N_15966,N_14653);
and U24177 (N_24177,N_13868,N_17959);
and U24178 (N_24178,N_12558,N_14115);
and U24179 (N_24179,N_15780,N_16120);
nand U24180 (N_24180,N_13188,N_17279);
nand U24181 (N_24181,N_17938,N_14134);
and U24182 (N_24182,N_13609,N_12583);
nor U24183 (N_24183,N_13107,N_13587);
or U24184 (N_24184,N_16591,N_16774);
nor U24185 (N_24185,N_12760,N_12884);
xor U24186 (N_24186,N_17314,N_17063);
xor U24187 (N_24187,N_17209,N_18613);
and U24188 (N_24188,N_17033,N_13519);
nor U24189 (N_24189,N_15232,N_13069);
nand U24190 (N_24190,N_17404,N_13275);
nor U24191 (N_24191,N_17487,N_13101);
nand U24192 (N_24192,N_14680,N_16190);
and U24193 (N_24193,N_17033,N_13490);
or U24194 (N_24194,N_14087,N_18104);
and U24195 (N_24195,N_17281,N_13739);
and U24196 (N_24196,N_13973,N_17026);
xnor U24197 (N_24197,N_17160,N_12565);
or U24198 (N_24198,N_17611,N_18519);
nor U24199 (N_24199,N_17960,N_15598);
and U24200 (N_24200,N_15070,N_15900);
xor U24201 (N_24201,N_16195,N_13040);
or U24202 (N_24202,N_12696,N_17090);
xnor U24203 (N_24203,N_13153,N_16530);
or U24204 (N_24204,N_17723,N_17622);
xnor U24205 (N_24205,N_18646,N_13553);
xor U24206 (N_24206,N_13865,N_13165);
nand U24207 (N_24207,N_13841,N_15900);
xor U24208 (N_24208,N_14334,N_14588);
and U24209 (N_24209,N_14541,N_17511);
nor U24210 (N_24210,N_13322,N_14662);
nand U24211 (N_24211,N_13002,N_17636);
or U24212 (N_24212,N_17252,N_15401);
nor U24213 (N_24213,N_16630,N_15542);
nand U24214 (N_24214,N_15447,N_16854);
xnor U24215 (N_24215,N_14207,N_12782);
xor U24216 (N_24216,N_15426,N_17588);
nor U24217 (N_24217,N_17982,N_13670);
nand U24218 (N_24218,N_17936,N_16100);
and U24219 (N_24219,N_15381,N_17275);
nand U24220 (N_24220,N_14352,N_15657);
nand U24221 (N_24221,N_12765,N_16615);
or U24222 (N_24222,N_16656,N_17675);
or U24223 (N_24223,N_14675,N_15398);
or U24224 (N_24224,N_15225,N_13340);
nand U24225 (N_24225,N_15325,N_12989);
xnor U24226 (N_24226,N_15498,N_14501);
nor U24227 (N_24227,N_16166,N_15300);
nand U24228 (N_24228,N_18592,N_18653);
or U24229 (N_24229,N_15556,N_15899);
nor U24230 (N_24230,N_13800,N_12791);
nand U24231 (N_24231,N_16854,N_17515);
nand U24232 (N_24232,N_14396,N_17152);
and U24233 (N_24233,N_17633,N_16006);
nand U24234 (N_24234,N_13183,N_16848);
and U24235 (N_24235,N_16808,N_12645);
nor U24236 (N_24236,N_16772,N_15082);
xor U24237 (N_24237,N_14242,N_18557);
or U24238 (N_24238,N_18095,N_13634);
nor U24239 (N_24239,N_13425,N_14813);
nand U24240 (N_24240,N_13298,N_18043);
or U24241 (N_24241,N_15335,N_16813);
or U24242 (N_24242,N_18190,N_15248);
and U24243 (N_24243,N_16043,N_15936);
and U24244 (N_24244,N_15711,N_16790);
xnor U24245 (N_24245,N_13812,N_18644);
nand U24246 (N_24246,N_14242,N_14721);
or U24247 (N_24247,N_14883,N_16887);
or U24248 (N_24248,N_16725,N_14406);
or U24249 (N_24249,N_17082,N_13381);
or U24250 (N_24250,N_17195,N_17476);
nor U24251 (N_24251,N_13374,N_14825);
nor U24252 (N_24252,N_16307,N_16934);
or U24253 (N_24253,N_13131,N_16695);
xor U24254 (N_24254,N_16041,N_14158);
xnor U24255 (N_24255,N_14426,N_12927);
or U24256 (N_24256,N_14180,N_15254);
and U24257 (N_24257,N_14960,N_18741);
or U24258 (N_24258,N_12815,N_13896);
nor U24259 (N_24259,N_18600,N_16408);
xor U24260 (N_24260,N_12577,N_15137);
xnor U24261 (N_24261,N_15916,N_17501);
and U24262 (N_24262,N_14198,N_13940);
or U24263 (N_24263,N_14388,N_13798);
and U24264 (N_24264,N_12585,N_12562);
xnor U24265 (N_24265,N_12744,N_15444);
and U24266 (N_24266,N_14447,N_18176);
and U24267 (N_24267,N_17007,N_16985);
nor U24268 (N_24268,N_17233,N_13261);
xor U24269 (N_24269,N_14376,N_16855);
or U24270 (N_24270,N_15712,N_13496);
xor U24271 (N_24271,N_15014,N_13120);
nor U24272 (N_24272,N_16065,N_15056);
and U24273 (N_24273,N_14001,N_16618);
and U24274 (N_24274,N_14344,N_17831);
or U24275 (N_24275,N_13699,N_18404);
xor U24276 (N_24276,N_13788,N_16795);
or U24277 (N_24277,N_16258,N_17201);
nor U24278 (N_24278,N_13975,N_15110);
or U24279 (N_24279,N_17233,N_15671);
nand U24280 (N_24280,N_17289,N_16462);
nand U24281 (N_24281,N_16320,N_18254);
or U24282 (N_24282,N_14595,N_17097);
or U24283 (N_24283,N_13392,N_16792);
or U24284 (N_24284,N_17800,N_18114);
xor U24285 (N_24285,N_17579,N_15306);
and U24286 (N_24286,N_13652,N_12582);
and U24287 (N_24287,N_15009,N_15932);
nor U24288 (N_24288,N_16109,N_14484);
xor U24289 (N_24289,N_15572,N_15540);
xor U24290 (N_24290,N_17687,N_12656);
nor U24291 (N_24291,N_18439,N_17063);
or U24292 (N_24292,N_17760,N_12638);
nor U24293 (N_24293,N_16727,N_15352);
and U24294 (N_24294,N_15787,N_17381);
xnor U24295 (N_24295,N_12525,N_16384);
or U24296 (N_24296,N_13341,N_17140);
nor U24297 (N_24297,N_14878,N_17094);
and U24298 (N_24298,N_17950,N_14798);
or U24299 (N_24299,N_15961,N_15832);
nor U24300 (N_24300,N_14141,N_14842);
or U24301 (N_24301,N_17662,N_14247);
and U24302 (N_24302,N_17087,N_17605);
xor U24303 (N_24303,N_13333,N_18555);
or U24304 (N_24304,N_17656,N_14051);
nor U24305 (N_24305,N_14947,N_16215);
or U24306 (N_24306,N_17936,N_17106);
and U24307 (N_24307,N_17543,N_13053);
nand U24308 (N_24308,N_18331,N_15099);
nand U24309 (N_24309,N_17364,N_18674);
nor U24310 (N_24310,N_14471,N_15123);
xor U24311 (N_24311,N_16860,N_14330);
xor U24312 (N_24312,N_16169,N_14889);
or U24313 (N_24313,N_17317,N_15495);
nor U24314 (N_24314,N_13609,N_16151);
xnor U24315 (N_24315,N_17588,N_16043);
nand U24316 (N_24316,N_13925,N_15525);
nor U24317 (N_24317,N_13752,N_16693);
nand U24318 (N_24318,N_18351,N_13488);
nand U24319 (N_24319,N_15400,N_14824);
nor U24320 (N_24320,N_13399,N_14800);
xnor U24321 (N_24321,N_15577,N_12811);
or U24322 (N_24322,N_12823,N_15536);
nor U24323 (N_24323,N_12802,N_12901);
nor U24324 (N_24324,N_14021,N_17261);
and U24325 (N_24325,N_14378,N_18414);
nand U24326 (N_24326,N_13621,N_17418);
xor U24327 (N_24327,N_16397,N_14068);
or U24328 (N_24328,N_14923,N_17727);
xnor U24329 (N_24329,N_16811,N_17524);
xnor U24330 (N_24330,N_13312,N_13504);
xnor U24331 (N_24331,N_15162,N_13188);
nor U24332 (N_24332,N_14659,N_16837);
xor U24333 (N_24333,N_14611,N_13901);
and U24334 (N_24334,N_15758,N_13663);
nand U24335 (N_24335,N_17339,N_18429);
xnor U24336 (N_24336,N_16304,N_14072);
and U24337 (N_24337,N_15252,N_16333);
nand U24338 (N_24338,N_17024,N_16786);
or U24339 (N_24339,N_17168,N_13760);
nor U24340 (N_24340,N_12970,N_14208);
xor U24341 (N_24341,N_13616,N_14670);
xnor U24342 (N_24342,N_13807,N_14584);
or U24343 (N_24343,N_15105,N_14598);
and U24344 (N_24344,N_16761,N_17029);
nand U24345 (N_24345,N_14644,N_14154);
xnor U24346 (N_24346,N_16248,N_17810);
nor U24347 (N_24347,N_18612,N_17819);
nor U24348 (N_24348,N_12811,N_16429);
and U24349 (N_24349,N_13987,N_13777);
and U24350 (N_24350,N_12867,N_16722);
nand U24351 (N_24351,N_14729,N_15227);
nor U24352 (N_24352,N_13117,N_17295);
xnor U24353 (N_24353,N_16314,N_16478);
nand U24354 (N_24354,N_14775,N_13284);
nor U24355 (N_24355,N_16702,N_18421);
xor U24356 (N_24356,N_16052,N_18304);
nor U24357 (N_24357,N_18169,N_16944);
or U24358 (N_24358,N_13739,N_15410);
xnor U24359 (N_24359,N_14145,N_16294);
nand U24360 (N_24360,N_15026,N_14174);
nand U24361 (N_24361,N_15544,N_17870);
nand U24362 (N_24362,N_16745,N_13272);
nor U24363 (N_24363,N_15276,N_14588);
nand U24364 (N_24364,N_16075,N_13067);
or U24365 (N_24365,N_13352,N_18711);
or U24366 (N_24366,N_12538,N_14591);
xnor U24367 (N_24367,N_17545,N_15655);
xnor U24368 (N_24368,N_18516,N_17316);
or U24369 (N_24369,N_14684,N_17762);
and U24370 (N_24370,N_13885,N_18584);
and U24371 (N_24371,N_15510,N_14099);
xnor U24372 (N_24372,N_17702,N_18563);
xor U24373 (N_24373,N_12897,N_18472);
xor U24374 (N_24374,N_18218,N_13989);
nor U24375 (N_24375,N_14788,N_15579);
nand U24376 (N_24376,N_17859,N_17930);
xor U24377 (N_24377,N_17381,N_14040);
xor U24378 (N_24378,N_12830,N_15091);
xor U24379 (N_24379,N_12637,N_17917);
and U24380 (N_24380,N_14681,N_18058);
nor U24381 (N_24381,N_16729,N_16085);
nor U24382 (N_24382,N_16185,N_12730);
and U24383 (N_24383,N_16219,N_14653);
and U24384 (N_24384,N_12950,N_14512);
nand U24385 (N_24385,N_14610,N_17370);
or U24386 (N_24386,N_13989,N_14356);
and U24387 (N_24387,N_15511,N_15667);
or U24388 (N_24388,N_13740,N_15530);
nand U24389 (N_24389,N_17541,N_15167);
nor U24390 (N_24390,N_16768,N_16549);
and U24391 (N_24391,N_12951,N_16932);
xor U24392 (N_24392,N_17741,N_17487);
nor U24393 (N_24393,N_16215,N_12653);
and U24394 (N_24394,N_16080,N_17605);
or U24395 (N_24395,N_17007,N_12618);
and U24396 (N_24396,N_13319,N_16315);
or U24397 (N_24397,N_17777,N_12508);
or U24398 (N_24398,N_16795,N_15367);
and U24399 (N_24399,N_12772,N_15328);
nand U24400 (N_24400,N_16968,N_15324);
nand U24401 (N_24401,N_18409,N_16130);
and U24402 (N_24402,N_13693,N_14155);
nand U24403 (N_24403,N_16628,N_13128);
or U24404 (N_24404,N_17010,N_12973);
and U24405 (N_24405,N_14725,N_13148);
xor U24406 (N_24406,N_16727,N_17058);
and U24407 (N_24407,N_17698,N_14878);
xnor U24408 (N_24408,N_14245,N_16602);
nor U24409 (N_24409,N_14841,N_12884);
xnor U24410 (N_24410,N_16152,N_16671);
and U24411 (N_24411,N_14232,N_15382);
nand U24412 (N_24412,N_18334,N_15064);
nor U24413 (N_24413,N_17718,N_14021);
nand U24414 (N_24414,N_15685,N_14467);
and U24415 (N_24415,N_13919,N_17068);
nor U24416 (N_24416,N_15337,N_13098);
or U24417 (N_24417,N_13800,N_13083);
nor U24418 (N_24418,N_13165,N_13373);
nand U24419 (N_24419,N_15413,N_17672);
xor U24420 (N_24420,N_14331,N_17623);
nor U24421 (N_24421,N_15452,N_14687);
and U24422 (N_24422,N_17411,N_14108);
nor U24423 (N_24423,N_14507,N_14088);
xor U24424 (N_24424,N_14254,N_16138);
nand U24425 (N_24425,N_18526,N_14244);
nand U24426 (N_24426,N_14400,N_13577);
nor U24427 (N_24427,N_17695,N_12944);
nor U24428 (N_24428,N_17720,N_13887);
nor U24429 (N_24429,N_16941,N_14699);
or U24430 (N_24430,N_18497,N_15848);
nor U24431 (N_24431,N_15038,N_18632);
nor U24432 (N_24432,N_18489,N_14071);
xor U24433 (N_24433,N_18532,N_17693);
or U24434 (N_24434,N_18669,N_18385);
nor U24435 (N_24435,N_13869,N_16180);
nor U24436 (N_24436,N_17300,N_14219);
nor U24437 (N_24437,N_13149,N_16396);
nand U24438 (N_24438,N_12613,N_16001);
nand U24439 (N_24439,N_15966,N_15381);
nor U24440 (N_24440,N_13532,N_15442);
xnor U24441 (N_24441,N_17538,N_17566);
nand U24442 (N_24442,N_16767,N_16861);
and U24443 (N_24443,N_17004,N_12798);
nor U24444 (N_24444,N_12762,N_18521);
nand U24445 (N_24445,N_15441,N_13438);
xor U24446 (N_24446,N_13880,N_15706);
nand U24447 (N_24447,N_14084,N_17224);
or U24448 (N_24448,N_17121,N_12957);
and U24449 (N_24449,N_14686,N_17911);
nor U24450 (N_24450,N_13312,N_15300);
nor U24451 (N_24451,N_16194,N_15776);
xor U24452 (N_24452,N_17335,N_18710);
nand U24453 (N_24453,N_17106,N_14982);
nor U24454 (N_24454,N_17759,N_15388);
nor U24455 (N_24455,N_13838,N_15710);
or U24456 (N_24456,N_16301,N_16626);
nor U24457 (N_24457,N_15534,N_13757);
xnor U24458 (N_24458,N_17563,N_13616);
xor U24459 (N_24459,N_17295,N_16824);
nor U24460 (N_24460,N_17341,N_16542);
and U24461 (N_24461,N_14331,N_15891);
nor U24462 (N_24462,N_13412,N_14244);
or U24463 (N_24463,N_12597,N_16302);
or U24464 (N_24464,N_15014,N_13481);
and U24465 (N_24465,N_14673,N_18558);
nor U24466 (N_24466,N_17918,N_16677);
nand U24467 (N_24467,N_13430,N_15393);
nor U24468 (N_24468,N_18204,N_14204);
nand U24469 (N_24469,N_17886,N_17652);
and U24470 (N_24470,N_13128,N_14886);
nand U24471 (N_24471,N_18632,N_14688);
xor U24472 (N_24472,N_17700,N_16561);
xor U24473 (N_24473,N_13697,N_18230);
nor U24474 (N_24474,N_18273,N_17003);
xnor U24475 (N_24475,N_16518,N_14166);
nor U24476 (N_24476,N_13510,N_14802);
xor U24477 (N_24477,N_17610,N_15980);
xnor U24478 (N_24478,N_18124,N_16605);
and U24479 (N_24479,N_14585,N_12599);
or U24480 (N_24480,N_14598,N_17922);
or U24481 (N_24481,N_18490,N_13291);
nand U24482 (N_24482,N_17280,N_16954);
xnor U24483 (N_24483,N_15353,N_12677);
xor U24484 (N_24484,N_16538,N_15518);
nand U24485 (N_24485,N_16294,N_13754);
nor U24486 (N_24486,N_18533,N_17555);
nor U24487 (N_24487,N_13271,N_15068);
and U24488 (N_24488,N_12736,N_14882);
nand U24489 (N_24489,N_13707,N_18487);
xnor U24490 (N_24490,N_14838,N_12805);
nand U24491 (N_24491,N_16389,N_16442);
nor U24492 (N_24492,N_13286,N_14805);
nand U24493 (N_24493,N_18017,N_15540);
and U24494 (N_24494,N_16264,N_18334);
or U24495 (N_24495,N_17949,N_16919);
nor U24496 (N_24496,N_16608,N_18718);
or U24497 (N_24497,N_17860,N_13035);
nor U24498 (N_24498,N_17935,N_15528);
nand U24499 (N_24499,N_15145,N_17649);
nor U24500 (N_24500,N_16471,N_13154);
xnor U24501 (N_24501,N_13550,N_15611);
or U24502 (N_24502,N_17761,N_15505);
or U24503 (N_24503,N_16576,N_16080);
and U24504 (N_24504,N_13297,N_13524);
and U24505 (N_24505,N_17300,N_13540);
nand U24506 (N_24506,N_16590,N_18171);
xnor U24507 (N_24507,N_14101,N_13039);
nor U24508 (N_24508,N_14261,N_17784);
and U24509 (N_24509,N_16090,N_14135);
xor U24510 (N_24510,N_18297,N_17767);
nand U24511 (N_24511,N_15990,N_16709);
and U24512 (N_24512,N_18186,N_18613);
and U24513 (N_24513,N_17569,N_18287);
or U24514 (N_24514,N_14488,N_16453);
xnor U24515 (N_24515,N_14997,N_13822);
or U24516 (N_24516,N_12540,N_15995);
xnor U24517 (N_24517,N_15555,N_14545);
xnor U24518 (N_24518,N_14063,N_17393);
nor U24519 (N_24519,N_17095,N_16221);
nor U24520 (N_24520,N_17003,N_17568);
nand U24521 (N_24521,N_15162,N_13921);
or U24522 (N_24522,N_14059,N_18117);
nand U24523 (N_24523,N_15868,N_13783);
or U24524 (N_24524,N_16327,N_15003);
and U24525 (N_24525,N_13067,N_17161);
and U24526 (N_24526,N_16480,N_13459);
nand U24527 (N_24527,N_16279,N_13170);
xor U24528 (N_24528,N_18719,N_15235);
nor U24529 (N_24529,N_14658,N_15875);
nand U24530 (N_24530,N_18219,N_12921);
nand U24531 (N_24531,N_12686,N_18466);
xnor U24532 (N_24532,N_16308,N_15432);
xor U24533 (N_24533,N_18080,N_14376);
and U24534 (N_24534,N_18677,N_15739);
nand U24535 (N_24535,N_14316,N_15265);
nor U24536 (N_24536,N_15827,N_15447);
nand U24537 (N_24537,N_13066,N_16836);
and U24538 (N_24538,N_12998,N_17607);
and U24539 (N_24539,N_15102,N_13941);
nor U24540 (N_24540,N_15599,N_17869);
and U24541 (N_24541,N_18570,N_13201);
and U24542 (N_24542,N_12628,N_17069);
nand U24543 (N_24543,N_14484,N_14530);
xnor U24544 (N_24544,N_16059,N_18683);
or U24545 (N_24545,N_13509,N_12988);
or U24546 (N_24546,N_17512,N_15975);
nor U24547 (N_24547,N_15961,N_18389);
nand U24548 (N_24548,N_16813,N_13155);
nor U24549 (N_24549,N_12590,N_17093);
or U24550 (N_24550,N_13107,N_13720);
xor U24551 (N_24551,N_16422,N_16373);
xnor U24552 (N_24552,N_16384,N_13971);
and U24553 (N_24553,N_14611,N_17273);
xor U24554 (N_24554,N_13772,N_16879);
or U24555 (N_24555,N_16597,N_13934);
xnor U24556 (N_24556,N_16779,N_15028);
and U24557 (N_24557,N_18568,N_16300);
or U24558 (N_24558,N_17039,N_16516);
or U24559 (N_24559,N_14767,N_16101);
xor U24560 (N_24560,N_12753,N_13892);
or U24561 (N_24561,N_15261,N_13356);
or U24562 (N_24562,N_12603,N_15137);
or U24563 (N_24563,N_13027,N_17746);
and U24564 (N_24564,N_17000,N_15589);
xor U24565 (N_24565,N_13779,N_14390);
nor U24566 (N_24566,N_12544,N_14529);
nor U24567 (N_24567,N_18079,N_17316);
nand U24568 (N_24568,N_14347,N_13008);
nor U24569 (N_24569,N_18417,N_13247);
nor U24570 (N_24570,N_14544,N_12703);
xor U24571 (N_24571,N_13581,N_15461);
nand U24572 (N_24572,N_16178,N_18518);
xor U24573 (N_24573,N_13628,N_18645);
nor U24574 (N_24574,N_18372,N_18555);
xnor U24575 (N_24575,N_17603,N_17248);
and U24576 (N_24576,N_14053,N_13052);
nor U24577 (N_24577,N_15367,N_16171);
or U24578 (N_24578,N_17373,N_13214);
xor U24579 (N_24579,N_17165,N_16806);
xnor U24580 (N_24580,N_16041,N_18151);
nand U24581 (N_24581,N_18010,N_17244);
xnor U24582 (N_24582,N_12697,N_13300);
or U24583 (N_24583,N_13453,N_18257);
xor U24584 (N_24584,N_18721,N_17688);
or U24585 (N_24585,N_18691,N_15393);
nand U24586 (N_24586,N_13348,N_16176);
nor U24587 (N_24587,N_14074,N_15001);
and U24588 (N_24588,N_18256,N_13747);
or U24589 (N_24589,N_17215,N_15314);
xor U24590 (N_24590,N_15569,N_13523);
or U24591 (N_24591,N_13875,N_16664);
and U24592 (N_24592,N_15036,N_16601);
xnor U24593 (N_24593,N_13891,N_17763);
nand U24594 (N_24594,N_15737,N_13909);
and U24595 (N_24595,N_17160,N_14527);
or U24596 (N_24596,N_15024,N_18175);
nor U24597 (N_24597,N_17660,N_13455);
or U24598 (N_24598,N_15248,N_14657);
nand U24599 (N_24599,N_16436,N_18123);
nand U24600 (N_24600,N_14172,N_13380);
or U24601 (N_24601,N_16921,N_12827);
nor U24602 (N_24602,N_16666,N_14828);
xnor U24603 (N_24603,N_18608,N_12511);
nor U24604 (N_24604,N_16794,N_18277);
nand U24605 (N_24605,N_15984,N_14688);
nor U24606 (N_24606,N_13943,N_17648);
and U24607 (N_24607,N_13323,N_13898);
xor U24608 (N_24608,N_17784,N_18391);
xor U24609 (N_24609,N_16817,N_14989);
nand U24610 (N_24610,N_16135,N_17843);
nand U24611 (N_24611,N_13629,N_15667);
nand U24612 (N_24612,N_13810,N_15047);
nand U24613 (N_24613,N_18679,N_13590);
xnor U24614 (N_24614,N_14227,N_15708);
nand U24615 (N_24615,N_17059,N_17737);
nor U24616 (N_24616,N_15140,N_15238);
and U24617 (N_24617,N_13219,N_17171);
nand U24618 (N_24618,N_17314,N_13811);
nand U24619 (N_24619,N_18270,N_12830);
and U24620 (N_24620,N_13584,N_16227);
or U24621 (N_24621,N_15525,N_13168);
nor U24622 (N_24622,N_18240,N_17606);
nor U24623 (N_24623,N_17201,N_17564);
and U24624 (N_24624,N_14160,N_13140);
or U24625 (N_24625,N_15347,N_16434);
or U24626 (N_24626,N_14146,N_14143);
nand U24627 (N_24627,N_16541,N_13951);
or U24628 (N_24628,N_18410,N_13272);
nor U24629 (N_24629,N_13211,N_16146);
xnor U24630 (N_24630,N_14140,N_13306);
or U24631 (N_24631,N_13022,N_16392);
nand U24632 (N_24632,N_13194,N_14870);
nor U24633 (N_24633,N_18180,N_16480);
or U24634 (N_24634,N_12617,N_17931);
and U24635 (N_24635,N_17454,N_13007);
xor U24636 (N_24636,N_15257,N_14186);
nor U24637 (N_24637,N_18420,N_14203);
xor U24638 (N_24638,N_17652,N_15237);
or U24639 (N_24639,N_15134,N_18253);
or U24640 (N_24640,N_15866,N_16755);
or U24641 (N_24641,N_12561,N_18172);
xnor U24642 (N_24642,N_15121,N_15247);
nand U24643 (N_24643,N_15547,N_17693);
nor U24644 (N_24644,N_17194,N_15665);
xor U24645 (N_24645,N_16256,N_12675);
xor U24646 (N_24646,N_17021,N_17736);
nand U24647 (N_24647,N_18299,N_12892);
and U24648 (N_24648,N_13015,N_17492);
or U24649 (N_24649,N_14128,N_17086);
nor U24650 (N_24650,N_15833,N_17949);
nor U24651 (N_24651,N_15636,N_17147);
xnor U24652 (N_24652,N_14483,N_14752);
xor U24653 (N_24653,N_18544,N_12614);
and U24654 (N_24654,N_18170,N_14330);
xnor U24655 (N_24655,N_15215,N_13550);
and U24656 (N_24656,N_14287,N_14653);
xnor U24657 (N_24657,N_15200,N_17903);
nor U24658 (N_24658,N_14716,N_14771);
nor U24659 (N_24659,N_15758,N_17197);
or U24660 (N_24660,N_14489,N_17100);
or U24661 (N_24661,N_15150,N_16604);
nand U24662 (N_24662,N_15246,N_18072);
xor U24663 (N_24663,N_18597,N_18447);
or U24664 (N_24664,N_16381,N_16800);
or U24665 (N_24665,N_15775,N_13718);
nand U24666 (N_24666,N_14161,N_18560);
xor U24667 (N_24667,N_17152,N_17424);
or U24668 (N_24668,N_18701,N_15481);
and U24669 (N_24669,N_13441,N_18227);
xnor U24670 (N_24670,N_17585,N_14543);
nand U24671 (N_24671,N_14450,N_13348);
or U24672 (N_24672,N_15452,N_12621);
nor U24673 (N_24673,N_12634,N_16335);
nand U24674 (N_24674,N_17776,N_18394);
nand U24675 (N_24675,N_16306,N_18243);
nand U24676 (N_24676,N_15545,N_14778);
and U24677 (N_24677,N_18570,N_16842);
xnor U24678 (N_24678,N_18111,N_15449);
and U24679 (N_24679,N_15539,N_15357);
and U24680 (N_24680,N_17164,N_14170);
or U24681 (N_24681,N_17913,N_17898);
or U24682 (N_24682,N_16796,N_18357);
xor U24683 (N_24683,N_14560,N_13661);
xnor U24684 (N_24684,N_14199,N_17401);
nand U24685 (N_24685,N_18237,N_14256);
nand U24686 (N_24686,N_16667,N_17507);
nand U24687 (N_24687,N_17822,N_13973);
xnor U24688 (N_24688,N_12695,N_15218);
or U24689 (N_24689,N_14186,N_17160);
or U24690 (N_24690,N_15947,N_16278);
nor U24691 (N_24691,N_17576,N_13932);
nor U24692 (N_24692,N_18532,N_15870);
xnor U24693 (N_24693,N_13059,N_17237);
nand U24694 (N_24694,N_14707,N_15648);
xor U24695 (N_24695,N_13178,N_13233);
or U24696 (N_24696,N_14699,N_16762);
xnor U24697 (N_24697,N_16554,N_14753);
nand U24698 (N_24698,N_17861,N_12726);
nand U24699 (N_24699,N_13573,N_13579);
or U24700 (N_24700,N_18378,N_12714);
nand U24701 (N_24701,N_18045,N_16298);
nor U24702 (N_24702,N_17331,N_18445);
nand U24703 (N_24703,N_16297,N_14727);
or U24704 (N_24704,N_13827,N_16566);
xnor U24705 (N_24705,N_16347,N_18581);
nand U24706 (N_24706,N_14623,N_12817);
or U24707 (N_24707,N_15293,N_16120);
nand U24708 (N_24708,N_17639,N_14057);
nand U24709 (N_24709,N_17498,N_18201);
and U24710 (N_24710,N_14309,N_18188);
nand U24711 (N_24711,N_16153,N_14594);
or U24712 (N_24712,N_15476,N_16958);
or U24713 (N_24713,N_13538,N_13095);
nor U24714 (N_24714,N_13804,N_18369);
or U24715 (N_24715,N_16992,N_12671);
and U24716 (N_24716,N_13284,N_13340);
nor U24717 (N_24717,N_13866,N_16846);
nor U24718 (N_24718,N_14793,N_17555);
or U24719 (N_24719,N_12964,N_13062);
or U24720 (N_24720,N_17895,N_17632);
nand U24721 (N_24721,N_17345,N_15285);
or U24722 (N_24722,N_14185,N_16847);
nor U24723 (N_24723,N_17109,N_14808);
nor U24724 (N_24724,N_14343,N_18373);
and U24725 (N_24725,N_16522,N_18114);
nand U24726 (N_24726,N_13591,N_13430);
and U24727 (N_24727,N_18075,N_17879);
xor U24728 (N_24728,N_18342,N_14379);
xor U24729 (N_24729,N_17335,N_14038);
nor U24730 (N_24730,N_14855,N_15204);
or U24731 (N_24731,N_13933,N_12508);
xnor U24732 (N_24732,N_18610,N_16272);
nand U24733 (N_24733,N_17570,N_13404);
nor U24734 (N_24734,N_17604,N_17434);
nor U24735 (N_24735,N_18650,N_16077);
nand U24736 (N_24736,N_17593,N_13848);
xnor U24737 (N_24737,N_16022,N_16883);
xor U24738 (N_24738,N_13553,N_16365);
or U24739 (N_24739,N_18288,N_14756);
nand U24740 (N_24740,N_16292,N_16869);
and U24741 (N_24741,N_13031,N_14896);
or U24742 (N_24742,N_16517,N_12840);
or U24743 (N_24743,N_14103,N_13809);
xnor U24744 (N_24744,N_16961,N_17023);
and U24745 (N_24745,N_15829,N_13417);
nand U24746 (N_24746,N_12600,N_14766);
or U24747 (N_24747,N_13824,N_12536);
xor U24748 (N_24748,N_15939,N_14535);
xor U24749 (N_24749,N_12669,N_17735);
and U24750 (N_24750,N_18103,N_16519);
or U24751 (N_24751,N_17631,N_17544);
and U24752 (N_24752,N_18265,N_14096);
nor U24753 (N_24753,N_12502,N_15134);
or U24754 (N_24754,N_15963,N_17420);
nand U24755 (N_24755,N_13180,N_13632);
or U24756 (N_24756,N_13832,N_16203);
nand U24757 (N_24757,N_15487,N_13826);
and U24758 (N_24758,N_17581,N_16835);
nor U24759 (N_24759,N_16749,N_14267);
nand U24760 (N_24760,N_17455,N_12980);
xor U24761 (N_24761,N_12836,N_15661);
or U24762 (N_24762,N_12612,N_13167);
or U24763 (N_24763,N_18358,N_12823);
xnor U24764 (N_24764,N_17677,N_14421);
and U24765 (N_24765,N_16327,N_13980);
xnor U24766 (N_24766,N_15987,N_18485);
xnor U24767 (N_24767,N_14876,N_14288);
nand U24768 (N_24768,N_18338,N_16772);
and U24769 (N_24769,N_16757,N_14469);
nand U24770 (N_24770,N_13633,N_17571);
nand U24771 (N_24771,N_13319,N_14485);
or U24772 (N_24772,N_14859,N_12688);
xor U24773 (N_24773,N_16714,N_16806);
and U24774 (N_24774,N_17570,N_12689);
nand U24775 (N_24775,N_14566,N_13813);
xnor U24776 (N_24776,N_18648,N_18076);
nand U24777 (N_24777,N_14369,N_16244);
and U24778 (N_24778,N_17709,N_14256);
nor U24779 (N_24779,N_15995,N_16076);
and U24780 (N_24780,N_14010,N_16430);
nor U24781 (N_24781,N_13839,N_18592);
nor U24782 (N_24782,N_18198,N_14900);
nor U24783 (N_24783,N_14169,N_12968);
xor U24784 (N_24784,N_15281,N_17126);
nand U24785 (N_24785,N_14660,N_13492);
xor U24786 (N_24786,N_18636,N_15798);
and U24787 (N_24787,N_14427,N_16259);
nand U24788 (N_24788,N_15477,N_14516);
nand U24789 (N_24789,N_16338,N_12631);
xor U24790 (N_24790,N_18182,N_12820);
or U24791 (N_24791,N_12943,N_18611);
nand U24792 (N_24792,N_15250,N_15231);
and U24793 (N_24793,N_17182,N_16036);
or U24794 (N_24794,N_14795,N_15109);
nor U24795 (N_24795,N_17288,N_17192);
and U24796 (N_24796,N_13601,N_16425);
nor U24797 (N_24797,N_16827,N_15550);
nand U24798 (N_24798,N_14435,N_15603);
and U24799 (N_24799,N_16696,N_14852);
or U24800 (N_24800,N_13369,N_14203);
and U24801 (N_24801,N_17381,N_13513);
xor U24802 (N_24802,N_16471,N_15401);
or U24803 (N_24803,N_18269,N_17795);
xnor U24804 (N_24804,N_16346,N_18677);
xor U24805 (N_24805,N_18524,N_14250);
or U24806 (N_24806,N_14160,N_12943);
nand U24807 (N_24807,N_14288,N_14684);
and U24808 (N_24808,N_18237,N_13829);
and U24809 (N_24809,N_12995,N_14905);
nor U24810 (N_24810,N_18689,N_17172);
xnor U24811 (N_24811,N_15700,N_17148);
and U24812 (N_24812,N_17370,N_18475);
nor U24813 (N_24813,N_14214,N_18061);
xor U24814 (N_24814,N_17168,N_16204);
or U24815 (N_24815,N_16777,N_15595);
and U24816 (N_24816,N_12630,N_14377);
or U24817 (N_24817,N_16327,N_16631);
or U24818 (N_24818,N_13220,N_18396);
xnor U24819 (N_24819,N_18724,N_17111);
and U24820 (N_24820,N_13513,N_12518);
and U24821 (N_24821,N_18094,N_12579);
or U24822 (N_24822,N_18037,N_15468);
and U24823 (N_24823,N_13083,N_18528);
nand U24824 (N_24824,N_13606,N_14207);
nor U24825 (N_24825,N_14195,N_12664);
and U24826 (N_24826,N_16050,N_17454);
nand U24827 (N_24827,N_15873,N_18699);
xor U24828 (N_24828,N_18384,N_17961);
or U24829 (N_24829,N_15298,N_13816);
nand U24830 (N_24830,N_13070,N_15040);
and U24831 (N_24831,N_17909,N_15530);
nor U24832 (N_24832,N_16671,N_14857);
or U24833 (N_24833,N_17723,N_14123);
nor U24834 (N_24834,N_17912,N_17492);
and U24835 (N_24835,N_15029,N_17707);
nand U24836 (N_24836,N_16465,N_14278);
or U24837 (N_24837,N_12568,N_16218);
nand U24838 (N_24838,N_17221,N_16031);
nand U24839 (N_24839,N_12630,N_17945);
nor U24840 (N_24840,N_17666,N_12562);
or U24841 (N_24841,N_13641,N_15401);
nand U24842 (N_24842,N_13413,N_14266);
and U24843 (N_24843,N_12608,N_15589);
and U24844 (N_24844,N_13046,N_14507);
nand U24845 (N_24845,N_17314,N_14564);
nand U24846 (N_24846,N_16102,N_16220);
xor U24847 (N_24847,N_12867,N_13964);
and U24848 (N_24848,N_15743,N_13320);
or U24849 (N_24849,N_16770,N_15825);
and U24850 (N_24850,N_14009,N_17912);
nor U24851 (N_24851,N_12790,N_15373);
and U24852 (N_24852,N_14557,N_14280);
or U24853 (N_24853,N_18610,N_16434);
and U24854 (N_24854,N_13309,N_18051);
or U24855 (N_24855,N_13404,N_15943);
nand U24856 (N_24856,N_18133,N_15909);
and U24857 (N_24857,N_13589,N_13186);
nor U24858 (N_24858,N_12736,N_15952);
and U24859 (N_24859,N_17667,N_16306);
nand U24860 (N_24860,N_14117,N_18021);
or U24861 (N_24861,N_17138,N_13219);
or U24862 (N_24862,N_14921,N_17087);
nor U24863 (N_24863,N_17817,N_15071);
or U24864 (N_24864,N_17705,N_18631);
or U24865 (N_24865,N_18336,N_13511);
or U24866 (N_24866,N_18255,N_15600);
xor U24867 (N_24867,N_12871,N_13115);
nand U24868 (N_24868,N_12564,N_15820);
nor U24869 (N_24869,N_12885,N_14436);
xnor U24870 (N_24870,N_16027,N_12522);
or U24871 (N_24871,N_15412,N_18654);
nand U24872 (N_24872,N_17623,N_15881);
xor U24873 (N_24873,N_13650,N_17704);
or U24874 (N_24874,N_18384,N_17807);
and U24875 (N_24875,N_18248,N_14333);
nor U24876 (N_24876,N_12722,N_17723);
or U24877 (N_24877,N_13522,N_17557);
nand U24878 (N_24878,N_15372,N_16587);
and U24879 (N_24879,N_16770,N_16362);
xor U24880 (N_24880,N_12871,N_13068);
or U24881 (N_24881,N_14765,N_14349);
and U24882 (N_24882,N_14992,N_13574);
nor U24883 (N_24883,N_15321,N_15798);
xnor U24884 (N_24884,N_17063,N_16796);
xor U24885 (N_24885,N_12918,N_15703);
nor U24886 (N_24886,N_14627,N_14332);
nor U24887 (N_24887,N_17049,N_17520);
and U24888 (N_24888,N_12916,N_12990);
nand U24889 (N_24889,N_17245,N_18034);
xor U24890 (N_24890,N_17153,N_16054);
and U24891 (N_24891,N_16960,N_16508);
nand U24892 (N_24892,N_17577,N_15889);
nor U24893 (N_24893,N_14166,N_18143);
and U24894 (N_24894,N_15081,N_16179);
nand U24895 (N_24895,N_17012,N_12632);
nand U24896 (N_24896,N_14491,N_14405);
nor U24897 (N_24897,N_13160,N_14825);
nor U24898 (N_24898,N_18205,N_16520);
xor U24899 (N_24899,N_15024,N_17668);
xor U24900 (N_24900,N_13909,N_18417);
and U24901 (N_24901,N_15211,N_15607);
xor U24902 (N_24902,N_18658,N_13442);
xor U24903 (N_24903,N_15176,N_14564);
xor U24904 (N_24904,N_15620,N_13766);
xnor U24905 (N_24905,N_13365,N_12874);
nand U24906 (N_24906,N_13625,N_12580);
nand U24907 (N_24907,N_18508,N_18467);
nand U24908 (N_24908,N_16962,N_14446);
xor U24909 (N_24909,N_15036,N_17907);
xnor U24910 (N_24910,N_18033,N_14118);
or U24911 (N_24911,N_17687,N_13820);
and U24912 (N_24912,N_18659,N_14250);
and U24913 (N_24913,N_12691,N_17368);
or U24914 (N_24914,N_14963,N_17725);
nand U24915 (N_24915,N_16987,N_18179);
xnor U24916 (N_24916,N_15959,N_16655);
nand U24917 (N_24917,N_15223,N_12844);
or U24918 (N_24918,N_14622,N_18338);
xnor U24919 (N_24919,N_18451,N_17812);
and U24920 (N_24920,N_14758,N_16628);
nor U24921 (N_24921,N_14195,N_15880);
or U24922 (N_24922,N_15654,N_15863);
nor U24923 (N_24923,N_14410,N_12604);
nor U24924 (N_24924,N_13552,N_12804);
or U24925 (N_24925,N_17578,N_12957);
nand U24926 (N_24926,N_13656,N_15618);
and U24927 (N_24927,N_12982,N_17662);
nand U24928 (N_24928,N_13443,N_16184);
nand U24929 (N_24929,N_14923,N_18407);
nor U24930 (N_24930,N_15680,N_17476);
nor U24931 (N_24931,N_18087,N_16701);
or U24932 (N_24932,N_15117,N_13747);
nand U24933 (N_24933,N_12689,N_13752);
or U24934 (N_24934,N_18431,N_16836);
nand U24935 (N_24935,N_16887,N_15561);
or U24936 (N_24936,N_12856,N_18213);
or U24937 (N_24937,N_13824,N_12634);
nor U24938 (N_24938,N_13800,N_16169);
nor U24939 (N_24939,N_18506,N_18645);
nor U24940 (N_24940,N_17863,N_13789);
nand U24941 (N_24941,N_16330,N_16574);
or U24942 (N_24942,N_13378,N_13301);
nor U24943 (N_24943,N_17669,N_17105);
nor U24944 (N_24944,N_15998,N_15657);
xor U24945 (N_24945,N_16200,N_16265);
and U24946 (N_24946,N_15744,N_12617);
nand U24947 (N_24947,N_16706,N_12914);
and U24948 (N_24948,N_16693,N_14288);
nor U24949 (N_24949,N_18724,N_15418);
nand U24950 (N_24950,N_13556,N_14364);
or U24951 (N_24951,N_16330,N_13506);
or U24952 (N_24952,N_17127,N_14047);
or U24953 (N_24953,N_17110,N_15149);
nor U24954 (N_24954,N_18483,N_15061);
xor U24955 (N_24955,N_16024,N_15856);
and U24956 (N_24956,N_15972,N_15957);
nand U24957 (N_24957,N_17216,N_17238);
nor U24958 (N_24958,N_12830,N_17267);
xnor U24959 (N_24959,N_16470,N_15398);
nor U24960 (N_24960,N_13554,N_17365);
and U24961 (N_24961,N_15850,N_17448);
xor U24962 (N_24962,N_17735,N_14180);
xnor U24963 (N_24963,N_15860,N_14240);
or U24964 (N_24964,N_12620,N_15420);
or U24965 (N_24965,N_16728,N_13114);
nor U24966 (N_24966,N_14451,N_16910);
or U24967 (N_24967,N_17610,N_14932);
nor U24968 (N_24968,N_14395,N_14953);
and U24969 (N_24969,N_15417,N_15759);
nand U24970 (N_24970,N_18744,N_15679);
nand U24971 (N_24971,N_17331,N_18326);
nand U24972 (N_24972,N_18384,N_13477);
and U24973 (N_24973,N_17391,N_15029);
or U24974 (N_24974,N_13758,N_14744);
xor U24975 (N_24975,N_13989,N_14983);
and U24976 (N_24976,N_18609,N_18695);
xor U24977 (N_24977,N_18141,N_18284);
or U24978 (N_24978,N_17110,N_13903);
xnor U24979 (N_24979,N_15369,N_12710);
or U24980 (N_24980,N_14669,N_16570);
and U24981 (N_24981,N_16620,N_15209);
nand U24982 (N_24982,N_13854,N_14444);
nand U24983 (N_24983,N_15530,N_17925);
and U24984 (N_24984,N_13633,N_16975);
or U24985 (N_24985,N_12776,N_16672);
nor U24986 (N_24986,N_14999,N_14372);
and U24987 (N_24987,N_13867,N_16514);
and U24988 (N_24988,N_13063,N_17487);
or U24989 (N_24989,N_18470,N_17141);
or U24990 (N_24990,N_14333,N_12749);
and U24991 (N_24991,N_18654,N_16209);
and U24992 (N_24992,N_16404,N_14719);
or U24993 (N_24993,N_13930,N_12994);
or U24994 (N_24994,N_16588,N_17426);
xor U24995 (N_24995,N_16919,N_16100);
nand U24996 (N_24996,N_14641,N_18575);
xor U24997 (N_24997,N_13411,N_17519);
nor U24998 (N_24998,N_18372,N_12868);
xor U24999 (N_24999,N_17329,N_14240);
nor UO_0 (O_0,N_18899,N_19697);
and UO_1 (O_1,N_24135,N_24277);
or UO_2 (O_2,N_23625,N_20290);
nand UO_3 (O_3,N_24006,N_24464);
or UO_4 (O_4,N_21937,N_20191);
or UO_5 (O_5,N_22191,N_24700);
nand UO_6 (O_6,N_23236,N_20014);
nor UO_7 (O_7,N_23753,N_18851);
xnor UO_8 (O_8,N_24812,N_23423);
xor UO_9 (O_9,N_22316,N_19734);
or UO_10 (O_10,N_23481,N_20761);
nor UO_11 (O_11,N_19528,N_22313);
nor UO_12 (O_12,N_19279,N_24578);
or UO_13 (O_13,N_24462,N_20617);
xnor UO_14 (O_14,N_24182,N_23885);
nor UO_15 (O_15,N_23595,N_21971);
nand UO_16 (O_16,N_24386,N_23091);
nor UO_17 (O_17,N_21489,N_20385);
xor UO_18 (O_18,N_19945,N_19406);
or UO_19 (O_19,N_23063,N_23280);
or UO_20 (O_20,N_23429,N_19491);
nor UO_21 (O_21,N_22854,N_23095);
and UO_22 (O_22,N_24769,N_20540);
nor UO_23 (O_23,N_19300,N_23331);
nand UO_24 (O_24,N_24230,N_24664);
nor UO_25 (O_25,N_22539,N_23802);
xnor UO_26 (O_26,N_20409,N_24860);
or UO_27 (O_27,N_21618,N_19322);
xnor UO_28 (O_28,N_18768,N_22711);
nor UO_29 (O_29,N_19329,N_23231);
nor UO_30 (O_30,N_20543,N_22591);
nand UO_31 (O_31,N_21554,N_20247);
or UO_32 (O_32,N_20489,N_21347);
nor UO_33 (O_33,N_24511,N_22922);
nor UO_34 (O_34,N_23448,N_22701);
nor UO_35 (O_35,N_24702,N_19567);
or UO_36 (O_36,N_21686,N_23165);
xor UO_37 (O_37,N_21607,N_22174);
xor UO_38 (O_38,N_23703,N_20101);
or UO_39 (O_39,N_18809,N_20765);
nand UO_40 (O_40,N_20737,N_21533);
nor UO_41 (O_41,N_22203,N_19564);
xnor UO_42 (O_42,N_19484,N_24460);
xnor UO_43 (O_43,N_23384,N_23870);
nand UO_44 (O_44,N_21332,N_19824);
xor UO_45 (O_45,N_22958,N_19664);
or UO_46 (O_46,N_22261,N_22264);
and UO_47 (O_47,N_24121,N_19969);
or UO_48 (O_48,N_22382,N_23037);
nor UO_49 (O_49,N_22433,N_21890);
nor UO_50 (O_50,N_22252,N_22153);
nor UO_51 (O_51,N_19580,N_23195);
and UO_52 (O_52,N_21737,N_24184);
and UO_53 (O_53,N_24770,N_20573);
and UO_54 (O_54,N_19098,N_20837);
or UO_55 (O_55,N_21804,N_23895);
xor UO_56 (O_56,N_19961,N_22414);
nor UO_57 (O_57,N_22534,N_20299);
xnor UO_58 (O_58,N_21628,N_19285);
or UO_59 (O_59,N_24715,N_19317);
xor UO_60 (O_60,N_22108,N_19554);
xnor UO_61 (O_61,N_24328,N_21519);
nor UO_62 (O_62,N_19553,N_24589);
or UO_63 (O_63,N_20957,N_22005);
xor UO_64 (O_64,N_21190,N_21078);
or UO_65 (O_65,N_19611,N_24630);
or UO_66 (O_66,N_22358,N_20240);
nor UO_67 (O_67,N_20411,N_21830);
nand UO_68 (O_68,N_18909,N_23103);
or UO_69 (O_69,N_19102,N_23270);
or UO_70 (O_70,N_20195,N_21598);
nor UO_71 (O_71,N_20781,N_22717);
xor UO_72 (O_72,N_23957,N_24965);
and UO_73 (O_73,N_20393,N_24424);
and UO_74 (O_74,N_24795,N_21179);
and UO_75 (O_75,N_21558,N_24943);
nand UO_76 (O_76,N_23377,N_24818);
nand UO_77 (O_77,N_24270,N_24895);
nor UO_78 (O_78,N_20924,N_24111);
nor UO_79 (O_79,N_22848,N_20034);
nor UO_80 (O_80,N_23849,N_24572);
and UO_81 (O_81,N_20580,N_19988);
and UO_82 (O_82,N_23482,N_24783);
xnor UO_83 (O_83,N_24995,N_23706);
nor UO_84 (O_84,N_19655,N_18763);
nand UO_85 (O_85,N_22975,N_19231);
nor UO_86 (O_86,N_24670,N_22079);
nor UO_87 (O_87,N_21876,N_19077);
nand UO_88 (O_88,N_21739,N_20357);
nand UO_89 (O_89,N_19157,N_24763);
nand UO_90 (O_90,N_22648,N_21509);
and UO_91 (O_91,N_23690,N_24740);
xor UO_92 (O_92,N_20990,N_23646);
nand UO_93 (O_93,N_19025,N_22175);
nand UO_94 (O_94,N_24421,N_21163);
nand UO_95 (O_95,N_21772,N_22551);
or UO_96 (O_96,N_20770,N_21637);
nor UO_97 (O_97,N_20007,N_23139);
and UO_98 (O_98,N_20552,N_22101);
xnor UO_99 (O_99,N_19042,N_21416);
nor UO_100 (O_100,N_19617,N_24312);
or UO_101 (O_101,N_24505,N_23055);
nand UO_102 (O_102,N_23830,N_19423);
nor UO_103 (O_103,N_19462,N_24202);
nor UO_104 (O_104,N_22051,N_20318);
nand UO_105 (O_105,N_24799,N_19134);
or UO_106 (O_106,N_20639,N_19670);
nand UO_107 (O_107,N_23379,N_21107);
xnor UO_108 (O_108,N_20287,N_22185);
nand UO_109 (O_109,N_21382,N_22508);
nand UO_110 (O_110,N_21999,N_24010);
nand UO_111 (O_111,N_19416,N_23712);
xor UO_112 (O_112,N_20129,N_22860);
and UO_113 (O_113,N_20105,N_23532);
nand UO_114 (O_114,N_19411,N_19514);
or UO_115 (O_115,N_19118,N_19414);
or UO_116 (O_116,N_21317,N_23577);
nand UO_117 (O_117,N_21459,N_22959);
nand UO_118 (O_118,N_21645,N_24959);
and UO_119 (O_119,N_24363,N_21353);
and UO_120 (O_120,N_18806,N_23921);
or UO_121 (O_121,N_19819,N_24502);
or UO_122 (O_122,N_24084,N_24128);
nand UO_123 (O_123,N_20584,N_20421);
xor UO_124 (O_124,N_20220,N_20766);
or UO_125 (O_125,N_19537,N_23940);
xor UO_126 (O_126,N_20417,N_20139);
xnor UO_127 (O_127,N_19494,N_19344);
or UO_128 (O_128,N_19777,N_23639);
and UO_129 (O_129,N_23111,N_24913);
xor UO_130 (O_130,N_18876,N_23444);
xnor UO_131 (O_131,N_20131,N_21716);
nand UO_132 (O_132,N_24489,N_22281);
or UO_133 (O_133,N_21540,N_21866);
or UO_134 (O_134,N_24908,N_20371);
xor UO_135 (O_135,N_19725,N_20301);
nand UO_136 (O_136,N_20069,N_20642);
or UO_137 (O_137,N_21206,N_20738);
xnor UO_138 (O_138,N_21796,N_23442);
and UO_139 (O_139,N_22920,N_23981);
nand UO_140 (O_140,N_21947,N_24169);
and UO_141 (O_141,N_19667,N_19066);
nand UO_142 (O_142,N_19064,N_23016);
and UO_143 (O_143,N_24894,N_23689);
or UO_144 (O_144,N_24619,N_22912);
nand UO_145 (O_145,N_22110,N_19804);
xnor UO_146 (O_146,N_24286,N_23651);
or UO_147 (O_147,N_24551,N_20078);
or UO_148 (O_148,N_24005,N_24017);
or UO_149 (O_149,N_20412,N_19900);
nor UO_150 (O_150,N_19361,N_21215);
nor UO_151 (O_151,N_21221,N_21478);
nand UO_152 (O_152,N_24416,N_20810);
and UO_153 (O_153,N_20051,N_22077);
xnor UO_154 (O_154,N_24170,N_24099);
nand UO_155 (O_155,N_20029,N_22790);
nand UO_156 (O_156,N_24532,N_22574);
or UO_157 (O_157,N_23036,N_21114);
nand UO_158 (O_158,N_24899,N_21004);
xnor UO_159 (O_159,N_23268,N_19549);
or UO_160 (O_160,N_20204,N_19366);
or UO_161 (O_161,N_20067,N_22291);
or UO_162 (O_162,N_22986,N_24616);
nand UO_163 (O_163,N_21100,N_23949);
xnor UO_164 (O_164,N_20481,N_23815);
nand UO_165 (O_165,N_22863,N_19103);
nor UO_166 (O_166,N_20043,N_19660);
nor UO_167 (O_167,N_24242,N_22978);
xor UO_168 (O_168,N_23796,N_20381);
or UO_169 (O_169,N_24023,N_22442);
and UO_170 (O_170,N_24678,N_21798);
xor UO_171 (O_171,N_20423,N_19793);
nand UO_172 (O_172,N_22159,N_23800);
or UO_173 (O_173,N_20877,N_19674);
nand UO_174 (O_174,N_19562,N_21160);
nor UO_175 (O_175,N_19033,N_22156);
xnor UO_176 (O_176,N_22980,N_21481);
nor UO_177 (O_177,N_24889,N_19812);
xor UO_178 (O_178,N_21968,N_24711);
nand UO_179 (O_179,N_20082,N_22049);
xor UO_180 (O_180,N_21122,N_22544);
xor UO_181 (O_181,N_22310,N_23627);
and UO_182 (O_182,N_23529,N_22803);
nand UO_183 (O_183,N_19270,N_18881);
and UO_184 (O_184,N_19653,N_21121);
xnor UO_185 (O_185,N_20668,N_21523);
nor UO_186 (O_186,N_22495,N_21886);
xor UO_187 (O_187,N_22248,N_19682);
xnor UO_188 (O_188,N_20510,N_24922);
xor UO_189 (O_189,N_20075,N_20901);
nand UO_190 (O_190,N_24669,N_24226);
nor UO_191 (O_191,N_19844,N_22541);
nand UO_192 (O_192,N_23265,N_19792);
and UO_193 (O_193,N_21172,N_20074);
nor UO_194 (O_194,N_20377,N_24171);
xnor UO_195 (O_195,N_20133,N_22670);
nand UO_196 (O_196,N_20793,N_21531);
xnor UO_197 (O_197,N_23929,N_21068);
xnor UO_198 (O_198,N_22964,N_21965);
nand UO_199 (O_199,N_18891,N_20464);
and UO_200 (O_200,N_23294,N_21434);
or UO_201 (O_201,N_21859,N_24928);
nand UO_202 (O_202,N_23705,N_19437);
or UO_203 (O_203,N_19364,N_19055);
nand UO_204 (O_204,N_24082,N_23147);
and UO_205 (O_205,N_23344,N_23758);
and UO_206 (O_206,N_20618,N_23022);
nand UO_207 (O_207,N_20647,N_23917);
nand UO_208 (O_208,N_19908,N_21015);
and UO_209 (O_209,N_23329,N_19786);
and UO_210 (O_210,N_19913,N_23743);
nand UO_211 (O_211,N_23585,N_24788);
xnor UO_212 (O_212,N_21575,N_24074);
and UO_213 (O_213,N_21504,N_19343);
and UO_214 (O_214,N_19519,N_23506);
or UO_215 (O_215,N_19629,N_24035);
nand UO_216 (O_216,N_19436,N_23660);
nand UO_217 (O_217,N_22205,N_24457);
nand UO_218 (O_218,N_19114,N_24317);
xnor UO_219 (O_219,N_22199,N_19807);
or UO_220 (O_220,N_24794,N_24036);
nor UO_221 (O_221,N_21195,N_20092);
and UO_222 (O_222,N_23029,N_24966);
and UO_223 (O_223,N_20307,N_22081);
or UO_224 (O_224,N_22809,N_19086);
xnor UO_225 (O_225,N_23163,N_20719);
or UO_226 (O_226,N_19937,N_20439);
and UO_227 (O_227,N_20872,N_20408);
or UO_228 (O_228,N_19334,N_21132);
or UO_229 (O_229,N_21211,N_20923);
and UO_230 (O_230,N_20685,N_24583);
or UO_231 (O_231,N_20081,N_23823);
nand UO_232 (O_232,N_22739,N_20087);
or UO_233 (O_233,N_22330,N_22145);
or UO_234 (O_234,N_19823,N_23552);
and UO_235 (O_235,N_22862,N_22475);
nor UO_236 (O_236,N_21367,N_22989);
and UO_237 (O_237,N_24797,N_20211);
and UO_238 (O_238,N_24584,N_22836);
xor UO_239 (O_239,N_21116,N_19142);
nand UO_240 (O_240,N_21566,N_20805);
nor UO_241 (O_241,N_22503,N_19376);
nor UO_242 (O_242,N_21874,N_21824);
xnor UO_243 (O_243,N_24150,N_19072);
or UO_244 (O_244,N_19596,N_20951);
nand UO_245 (O_245,N_18829,N_23038);
nor UO_246 (O_246,N_22824,N_21024);
nor UO_247 (O_247,N_18939,N_24166);
and UO_248 (O_248,N_24628,N_24605);
nand UO_249 (O_249,N_24696,N_18925);
or UO_250 (O_250,N_20525,N_23638);
xnor UO_251 (O_251,N_22143,N_23395);
or UO_252 (O_252,N_21082,N_20746);
xor UO_253 (O_253,N_22131,N_22280);
nor UO_254 (O_254,N_18785,N_19798);
nand UO_255 (O_255,N_23749,N_19885);
or UO_256 (O_256,N_24534,N_19840);
nand UO_257 (O_257,N_24806,N_19613);
or UO_258 (O_258,N_20223,N_24701);
xnor UO_259 (O_259,N_21563,N_20836);
xnor UO_260 (O_260,N_23900,N_21774);
nand UO_261 (O_261,N_20742,N_23459);
or UO_262 (O_262,N_21003,N_19910);
or UO_263 (O_263,N_23581,N_23297);
nand UO_264 (O_264,N_24050,N_24634);
xor UO_265 (O_265,N_23347,N_21544);
nor UO_266 (O_266,N_24064,N_20401);
nor UO_267 (O_267,N_20148,N_19453);
nand UO_268 (O_268,N_20531,N_24427);
or UO_269 (O_269,N_22764,N_21105);
and UO_270 (O_270,N_24767,N_19310);
or UO_271 (O_271,N_23741,N_18874);
or UO_272 (O_272,N_22543,N_20415);
nor UO_273 (O_273,N_20042,N_21313);
or UO_274 (O_274,N_20047,N_19480);
or UO_275 (O_275,N_23164,N_22781);
nor UO_276 (O_276,N_21421,N_21695);
or UO_277 (O_277,N_20689,N_24494);
xnor UO_278 (O_278,N_21721,N_24436);
xnor UO_279 (O_279,N_22309,N_19545);
xnor UO_280 (O_280,N_18865,N_21401);
nor UO_281 (O_281,N_19417,N_18797);
or UO_282 (O_282,N_21460,N_21209);
xor UO_283 (O_283,N_20270,N_24401);
xor UO_284 (O_284,N_23953,N_20600);
nand UO_285 (O_285,N_23228,N_21461);
nand UO_286 (O_286,N_24495,N_24685);
or UO_287 (O_287,N_22103,N_21120);
nor UO_288 (O_288,N_22664,N_18779);
or UO_289 (O_289,N_18811,N_23669);
and UO_290 (O_290,N_21011,N_23736);
and UO_291 (O_291,N_24964,N_23338);
nor UO_292 (O_292,N_23093,N_18992);
nor UO_293 (O_293,N_21560,N_20355);
nand UO_294 (O_294,N_24252,N_20593);
nor UO_295 (O_295,N_23237,N_20795);
nand UO_296 (O_296,N_18756,N_20545);
and UO_297 (O_297,N_19335,N_22961);
and UO_298 (O_298,N_22142,N_20321);
xnor UO_299 (O_299,N_19022,N_20595);
and UO_300 (O_300,N_21660,N_22882);
nor UO_301 (O_301,N_19657,N_19162);
nor UO_302 (O_302,N_22260,N_18833);
nor UO_303 (O_303,N_21166,N_24469);
or UO_304 (O_304,N_22188,N_19923);
or UO_305 (O_305,N_23845,N_19760);
or UO_306 (O_306,N_19618,N_23335);
nor UO_307 (O_307,N_22467,N_23304);
nor UO_308 (O_308,N_23558,N_19280);
or UO_309 (O_309,N_22925,N_19772);
nor UO_310 (O_310,N_24233,N_18772);
and UO_311 (O_311,N_23198,N_20504);
nor UO_312 (O_312,N_21222,N_21070);
xor UO_313 (O_313,N_23871,N_24671);
nor UO_314 (O_314,N_21827,N_20019);
xnor UO_315 (O_315,N_21779,N_23194);
nand UO_316 (O_316,N_24138,N_20285);
xnor UO_317 (O_317,N_21091,N_24380);
or UO_318 (O_318,N_19836,N_24565);
nor UO_319 (O_319,N_21281,N_21298);
nor UO_320 (O_320,N_19112,N_20707);
nor UO_321 (O_321,N_19048,N_21699);
nor UO_322 (O_322,N_23186,N_20035);
or UO_323 (O_323,N_20676,N_19707);
nand UO_324 (O_324,N_18751,N_19152);
xnor UO_325 (O_325,N_24249,N_23526);
and UO_326 (O_326,N_22597,N_19950);
xor UO_327 (O_327,N_24823,N_21917);
nor UO_328 (O_328,N_22094,N_24553);
xor UO_329 (O_329,N_23708,N_19234);
and UO_330 (O_330,N_19499,N_22960);
or UO_331 (O_331,N_21199,N_22001);
xnor UO_332 (O_332,N_20296,N_20609);
nor UO_333 (O_333,N_21549,N_21342);
or UO_334 (O_334,N_21735,N_24548);
nand UO_335 (O_335,N_21914,N_21200);
nor UO_336 (O_336,N_23618,N_20115);
xnor UO_337 (O_337,N_23601,N_20232);
xor UO_338 (O_338,N_23589,N_19828);
and UO_339 (O_339,N_23279,N_20369);
nor UO_340 (O_340,N_22259,N_21335);
xnor UO_341 (O_341,N_21500,N_20396);
or UO_342 (O_342,N_21996,N_23977);
or UO_343 (O_343,N_19225,N_24311);
nor UO_344 (O_344,N_19123,N_19337);
or UO_345 (O_345,N_21064,N_22977);
or UO_346 (O_346,N_19432,N_18770);
nor UO_347 (O_347,N_20340,N_22704);
and UO_348 (O_348,N_23383,N_20216);
nor UO_349 (O_349,N_24159,N_19435);
xor UO_350 (O_350,N_18917,N_20945);
nand UO_351 (O_351,N_21662,N_24835);
nand UO_352 (O_352,N_19294,N_20127);
nand UO_353 (O_353,N_22378,N_22288);
or UO_354 (O_354,N_23407,N_19221);
xor UO_355 (O_355,N_20845,N_19825);
and UO_356 (O_356,N_19919,N_23006);
xnor UO_357 (O_357,N_23653,N_21256);
nand UO_358 (O_358,N_20454,N_18802);
or UO_359 (O_359,N_18952,N_20027);
or UO_360 (O_360,N_20677,N_22913);
and UO_361 (O_361,N_22522,N_21633);
nand UO_362 (O_362,N_18974,N_22839);
nor UO_363 (O_363,N_19744,N_20244);
nor UO_364 (O_364,N_22010,N_22741);
and UO_365 (O_365,N_20063,N_23611);
xor UO_366 (O_366,N_21128,N_20817);
and UO_367 (O_367,N_23762,N_21518);
and UO_368 (O_368,N_23969,N_21168);
nand UO_369 (O_369,N_20851,N_20869);
nand UO_370 (O_370,N_20266,N_22660);
nor UO_371 (O_371,N_24007,N_18813);
and UO_372 (O_372,N_19560,N_19496);
nand UO_373 (O_373,N_22738,N_24383);
nor UO_374 (O_374,N_23746,N_23243);
xnor UO_375 (O_375,N_19403,N_20346);
xor UO_376 (O_376,N_19184,N_22691);
xor UO_377 (O_377,N_20205,N_24869);
and UO_378 (O_378,N_21980,N_24490);
nand UO_379 (O_379,N_20784,N_23944);
and UO_380 (O_380,N_23851,N_19522);
or UO_381 (O_381,N_24622,N_22111);
or UO_382 (O_382,N_21058,N_19626);
nor UO_383 (O_383,N_22472,N_21276);
xnor UO_384 (O_384,N_19196,N_20916);
or UO_385 (O_385,N_23542,N_23978);
and UO_386 (O_386,N_24420,N_24463);
or UO_387 (O_387,N_20966,N_19565);
nand UO_388 (O_388,N_24732,N_19952);
xor UO_389 (O_389,N_22679,N_23783);
nor UO_390 (O_390,N_21698,N_19358);
xor UO_391 (O_391,N_23230,N_22161);
or UO_392 (O_392,N_23426,N_22416);
and UO_393 (O_393,N_22407,N_21530);
nor UO_394 (O_394,N_23816,N_21701);
nor UO_395 (O_395,N_18987,N_20124);
xnor UO_396 (O_396,N_20878,N_22703);
and UO_397 (O_397,N_24103,N_20790);
nor UO_398 (O_398,N_19701,N_22976);
nand UO_399 (O_399,N_18774,N_22903);
and UO_400 (O_400,N_19547,N_22804);
nor UO_401 (O_401,N_21205,N_23089);
or UO_402 (O_402,N_23214,N_21189);
and UO_403 (O_403,N_21978,N_20335);
nor UO_404 (O_404,N_22215,N_21738);
nor UO_405 (O_405,N_22319,N_20432);
and UO_406 (O_406,N_19085,N_20775);
or UO_407 (O_407,N_19419,N_21600);
and UO_408 (O_408,N_23599,N_22088);
nor UO_409 (O_409,N_20233,N_22087);
xnor UO_410 (O_410,N_24196,N_23531);
or UO_411 (O_411,N_23702,N_20777);
and UO_412 (O_412,N_23612,N_20449);
or UO_413 (O_413,N_22604,N_24115);
nand UO_414 (O_414,N_24178,N_23342);
nor UO_415 (O_415,N_20820,N_23242);
xor UO_416 (O_416,N_24606,N_21878);
nand UO_417 (O_417,N_19281,N_23856);
or UO_418 (O_418,N_20606,N_18857);
nand UO_419 (O_419,N_21821,N_19446);
xnor UO_420 (O_420,N_23614,N_21788);
nor UO_421 (O_421,N_23797,N_19780);
nor UO_422 (O_422,N_21644,N_18830);
or UO_423 (O_423,N_24626,N_19986);
nor UO_424 (O_424,N_24602,N_22428);
nor UO_425 (O_425,N_21767,N_20583);
or UO_426 (O_426,N_20164,N_21057);
nor UO_427 (O_427,N_23927,N_21895);
and UO_428 (O_428,N_23670,N_19972);
or UO_429 (O_429,N_20895,N_20814);
and UO_430 (O_430,N_19014,N_24917);
nor UO_431 (O_431,N_22355,N_19267);
xor UO_432 (O_432,N_20275,N_23789);
and UO_433 (O_433,N_23661,N_22929);
and UO_434 (O_434,N_23854,N_20844);
xor UO_435 (O_435,N_23245,N_21696);
xnor UO_436 (O_436,N_19286,N_19607);
and UO_437 (O_437,N_24435,N_22201);
nand UO_438 (O_438,N_21594,N_21568);
nand UO_439 (O_439,N_19845,N_20918);
or UO_440 (O_440,N_21173,N_19313);
or UO_441 (O_441,N_22083,N_23617);
or UO_442 (O_442,N_23697,N_19365);
xor UO_443 (O_443,N_20280,N_19409);
nand UO_444 (O_444,N_21253,N_21389);
xnor UO_445 (O_445,N_24681,N_24815);
and UO_446 (O_446,N_22939,N_22012);
nor UO_447 (O_447,N_23907,N_20203);
nand UO_448 (O_448,N_18805,N_23381);
nand UO_449 (O_449,N_19594,N_23945);
nor UO_450 (O_450,N_24322,N_22021);
and UO_451 (O_451,N_23346,N_18877);
nor UO_452 (O_452,N_22745,N_20711);
or UO_453 (O_453,N_21156,N_19268);
and UO_454 (O_454,N_20626,N_21994);
or UO_455 (O_455,N_20054,N_22471);
nor UO_456 (O_456,N_19951,N_22099);
or UO_457 (O_457,N_21169,N_19255);
xor UO_458 (O_458,N_20947,N_18873);
xor UO_459 (O_459,N_22155,N_20477);
nand UO_460 (O_460,N_20208,N_22726);
nor UO_461 (O_461,N_22511,N_18823);
or UO_462 (O_462,N_22890,N_20537);
or UO_463 (O_463,N_23368,N_23579);
xor UO_464 (O_464,N_24225,N_21577);
nor UO_465 (O_465,N_23152,N_20554);
nor UO_466 (O_466,N_19752,N_19478);
nor UO_467 (O_467,N_24388,N_19941);
nand UO_468 (O_468,N_22454,N_24570);
xor UO_469 (O_469,N_20031,N_22942);
xor UO_470 (O_470,N_19485,N_23389);
or UO_471 (O_471,N_22512,N_23414);
or UO_472 (O_472,N_22399,N_24198);
xnor UO_473 (O_473,N_22200,N_23416);
nand UO_474 (O_474,N_24391,N_23366);
or UO_475 (O_475,N_19367,N_20843);
or UO_476 (O_476,N_22292,N_20444);
nor UO_477 (O_477,N_19604,N_19608);
and UO_478 (O_478,N_18965,N_18982);
nor UO_479 (O_479,N_19016,N_19766);
xor UO_480 (O_480,N_20474,N_20722);
xor UO_481 (O_481,N_19850,N_18961);
and UO_482 (O_482,N_19727,N_24747);
nand UO_483 (O_483,N_18815,N_19301);
and UO_484 (O_484,N_23999,N_24656);
nand UO_485 (O_485,N_22908,N_20659);
and UO_486 (O_486,N_21148,N_19330);
or UO_487 (O_487,N_24524,N_20037);
or UO_488 (O_488,N_20492,N_22400);
nor UO_489 (O_489,N_21274,N_24560);
nor UO_490 (O_490,N_18926,N_20395);
and UO_491 (O_491,N_19465,N_24620);
and UO_492 (O_492,N_21073,N_24264);
nand UO_493 (O_493,N_20892,N_19694);
xnor UO_494 (O_494,N_22889,N_24774);
xor UO_495 (O_495,N_19771,N_20509);
nor UO_496 (O_496,N_21555,N_21809);
nor UO_497 (O_497,N_19190,N_21901);
nor UO_498 (O_498,N_18783,N_20565);
xnor UO_499 (O_499,N_23880,N_19810);
xnor UO_500 (O_500,N_22232,N_22130);
and UO_501 (O_501,N_19930,N_20846);
nand UO_502 (O_502,N_23225,N_19800);
or UO_503 (O_503,N_19838,N_24720);
xnor UO_504 (O_504,N_20832,N_18973);
nand UO_505 (O_505,N_20438,N_20100);
nor UO_506 (O_506,N_24831,N_19525);
nand UO_507 (O_507,N_21028,N_19314);
nand UO_508 (O_508,N_22444,N_19628);
nor UO_509 (O_509,N_21605,N_22253);
nand UO_510 (O_510,N_24481,N_19139);
nor UO_511 (O_511,N_20995,N_19614);
or UO_512 (O_512,N_24885,N_24475);
or UO_513 (O_513,N_23457,N_19402);
and UO_514 (O_514,N_23431,N_20182);
and UO_515 (O_515,N_21063,N_20468);
and UO_516 (O_516,N_23108,N_23396);
or UO_517 (O_517,N_24223,N_23803);
xnor UO_518 (O_518,N_22752,N_24297);
xor UO_519 (O_519,N_20094,N_24652);
xor UO_520 (O_520,N_24951,N_22709);
and UO_521 (O_521,N_20267,N_19161);
or UO_522 (O_522,N_23156,N_20006);
or UO_523 (O_523,N_23151,N_21470);
nand UO_524 (O_524,N_21921,N_22579);
nand UO_525 (O_525,N_24131,N_20348);
xor UO_526 (O_526,N_20522,N_23348);
nand UO_527 (O_527,N_19336,N_22783);
or UO_528 (O_528,N_24011,N_19678);
nor UO_529 (O_529,N_24786,N_22538);
and UO_530 (O_530,N_19665,N_22505);
and UO_531 (O_531,N_22056,N_18990);
nand UO_532 (O_532,N_21235,N_21458);
xor UO_533 (O_533,N_19718,N_21280);
xnor UO_534 (O_534,N_19524,N_22880);
and UO_535 (O_535,N_19349,N_24404);
nor UO_536 (O_536,N_24629,N_22693);
or UO_537 (O_537,N_18921,N_24938);
or UO_538 (O_538,N_23040,N_18755);
nor UO_539 (O_539,N_23308,N_20715);
and UO_540 (O_540,N_21376,N_23591);
or UO_541 (O_541,N_23148,N_19814);
xor UO_542 (O_542,N_23436,N_23382);
xor UO_543 (O_543,N_19263,N_23085);
xnor UO_544 (O_544,N_23105,N_24520);
nand UO_545 (O_545,N_22173,N_22016);
nand UO_546 (O_546,N_24221,N_22931);
or UO_547 (O_547,N_20091,N_24648);
nor UO_548 (O_548,N_24516,N_21888);
or UO_549 (O_549,N_21037,N_22446);
nor UO_550 (O_550,N_24549,N_22861);
and UO_551 (O_551,N_19650,N_23309);
or UO_552 (O_552,N_22676,N_20987);
or UO_553 (O_553,N_24948,N_21268);
nand UO_554 (O_554,N_21547,N_24079);
or UO_555 (O_555,N_20062,N_21728);
nand UO_556 (O_556,N_22314,N_20978);
nor UO_557 (O_557,N_22024,N_19782);
nor UO_558 (O_558,N_19037,N_19641);
xnor UO_559 (O_559,N_19477,N_23810);
nand UO_560 (O_560,N_21957,N_21718);
xnor UO_561 (O_561,N_23136,N_24210);
or UO_562 (O_562,N_20708,N_20733);
nor UO_563 (O_563,N_20762,N_23087);
or UO_564 (O_564,N_23932,N_21186);
xnor UO_565 (O_565,N_21218,N_20483);
or UO_566 (O_566,N_24144,N_20494);
nor UO_567 (O_567,N_24576,N_20842);
nor UO_568 (O_568,N_22778,N_22523);
or UO_569 (O_569,N_23315,N_24741);
nor UO_570 (O_570,N_19443,N_21527);
and UO_571 (O_571,N_18765,N_19668);
xnor UO_572 (O_572,N_24423,N_22699);
or UO_573 (O_573,N_18986,N_24186);
or UO_574 (O_574,N_24174,N_19895);
nor UO_575 (O_575,N_23826,N_19254);
nor UO_576 (O_576,N_21087,N_22146);
or UO_577 (O_577,N_18962,N_24092);
or UO_578 (O_578,N_24827,N_24308);
or UO_579 (O_579,N_20496,N_20404);
and UO_580 (O_580,N_24603,N_19296);
xnor UO_581 (O_581,N_19981,N_24353);
or UO_582 (O_582,N_21203,N_20425);
and UO_583 (O_583,N_20759,N_24029);
or UO_584 (O_584,N_20931,N_19993);
nand UO_585 (O_585,N_21278,N_21141);
nor UO_586 (O_586,N_20379,N_24923);
or UO_587 (O_587,N_22702,N_21867);
xnor UO_588 (O_588,N_19976,N_23915);
nand UO_589 (O_589,N_24290,N_19606);
nor UO_590 (O_590,N_24803,N_22426);
xnor UO_591 (O_591,N_23356,N_18795);
or UO_592 (O_592,N_19773,N_23805);
xor UO_593 (O_593,N_22638,N_24704);
xnor UO_594 (O_594,N_23972,N_19968);
xor UO_595 (O_595,N_22509,N_19346);
nand UO_596 (O_596,N_21476,N_19622);
xnor UO_597 (O_597,N_24980,N_19983);
xnor UO_598 (O_598,N_18953,N_21007);
nor UO_599 (O_599,N_20693,N_21623);
nor UO_600 (O_600,N_22468,N_23290);
and UO_601 (O_601,N_19404,N_20327);
xor UO_602 (O_602,N_18787,N_20839);
or UO_603 (O_603,N_20002,N_23551);
and UO_604 (O_604,N_23123,N_19681);
nand UO_605 (O_605,N_20134,N_21842);
nand UO_606 (O_606,N_20607,N_19898);
or UO_607 (O_607,N_22068,N_19872);
nor UO_608 (O_608,N_21768,N_21778);
nand UO_609 (O_609,N_24478,N_20801);
xor UO_610 (O_610,N_23954,N_21426);
nand UO_611 (O_611,N_23947,N_24726);
nand UO_612 (O_612,N_21170,N_24283);
or UO_613 (O_613,N_24239,N_21440);
xnor UO_614 (O_614,N_24850,N_19345);
nand UO_615 (O_615,N_24047,N_20611);
xnor UO_616 (O_616,N_24585,N_21296);
nand UO_617 (O_617,N_19692,N_22402);
xnor UO_618 (O_618,N_21498,N_21366);
nor UO_619 (O_619,N_23973,N_21746);
nor UO_620 (O_620,N_22125,N_22045);
xor UO_621 (O_621,N_21732,N_20827);
xor UO_622 (O_622,N_21129,N_23633);
nand UO_623 (O_623,N_22194,N_23820);
or UO_624 (O_624,N_22570,N_24122);
nor UO_625 (O_625,N_19095,N_20085);
nor UO_626 (O_626,N_22169,N_19307);
nand UO_627 (O_627,N_19218,N_19174);
nand UO_628 (O_628,N_21651,N_19362);
nand UO_629 (O_629,N_19011,N_22213);
and UO_630 (O_630,N_24461,N_19532);
xnor UO_631 (O_631,N_21625,N_19967);
and UO_632 (O_632,N_23145,N_20643);
xor UO_633 (O_633,N_23761,N_23545);
or UO_634 (O_634,N_21766,N_24257);
xnor UO_635 (O_635,N_23686,N_24915);
nor UO_636 (O_636,N_19866,N_23597);
xnor UO_637 (O_637,N_20748,N_19561);
or UO_638 (O_638,N_20960,N_24412);
or UO_639 (O_639,N_19520,N_22469);
nand UO_640 (O_640,N_19839,N_24327);
nor UO_641 (O_641,N_22189,N_24352);
nor UO_642 (O_642,N_20942,N_22246);
and UO_643 (O_643,N_22616,N_22568);
or UO_644 (O_644,N_22226,N_18866);
or UO_645 (O_645,N_19568,N_19570);
xnor UO_646 (O_646,N_22282,N_24789);
and UO_647 (O_647,N_24861,N_19258);
nor UO_648 (O_648,N_24146,N_23306);
or UO_649 (O_649,N_20880,N_22518);
nor UO_650 (O_650,N_20214,N_21387);
nand UO_651 (O_651,N_24708,N_22899);
xor UO_652 (O_652,N_24484,N_24642);
xnor UO_653 (O_653,N_21945,N_24623);
nand UO_654 (O_654,N_19687,N_22949);
and UO_655 (O_655,N_20390,N_19487);
and UO_656 (O_656,N_21485,N_18972);
and UO_657 (O_657,N_18946,N_20602);
xor UO_658 (O_658,N_20117,N_24838);
or UO_659 (O_659,N_21339,N_23154);
or UO_660 (O_660,N_20156,N_21334);
and UO_661 (O_661,N_23053,N_19204);
nand UO_662 (O_662,N_19309,N_20479);
nor UO_663 (O_663,N_21524,N_21959);
and UO_664 (O_664,N_20658,N_20910);
nor UO_665 (O_665,N_20819,N_23118);
or UO_666 (O_666,N_23667,N_24102);
or UO_667 (O_667,N_22995,N_19616);
or UO_668 (O_668,N_21720,N_21970);
or UO_669 (O_669,N_21055,N_22046);
or UO_670 (O_670,N_22716,N_20723);
nand UO_671 (O_671,N_19027,N_22540);
and UO_672 (O_672,N_20912,N_21176);
and UO_673 (O_673,N_19452,N_18750);
xor UO_674 (O_674,N_21667,N_20300);
and UO_675 (O_675,N_19779,N_23460);
nor UO_676 (O_676,N_19505,N_19220);
and UO_677 (O_677,N_23435,N_20077);
and UO_678 (O_678,N_22553,N_20589);
or UO_679 (O_679,N_20768,N_19169);
xnor UO_680 (O_680,N_20705,N_23520);
and UO_681 (O_681,N_22090,N_19956);
or UO_682 (O_682,N_24668,N_23750);
and UO_683 (O_683,N_23124,N_21158);
xnor UO_684 (O_684,N_19451,N_18859);
nand UO_685 (O_685,N_21741,N_22178);
or UO_686 (O_686,N_19106,N_23258);
or UO_687 (O_687,N_19706,N_24052);
nor UO_688 (O_688,N_21657,N_19936);
or UO_689 (O_689,N_22067,N_21583);
and UO_690 (O_690,N_22439,N_21032);
xnor UO_691 (O_691,N_23131,N_19428);
xnor UO_692 (O_692,N_21153,N_22601);
xnor UO_693 (O_693,N_19156,N_22004);
or UO_694 (O_694,N_20886,N_23068);
nand UO_695 (O_695,N_19046,N_24607);
or UO_696 (O_696,N_20785,N_23391);
and UO_697 (O_697,N_19517,N_24057);
xnor UO_698 (O_698,N_23310,N_24745);
and UO_699 (O_699,N_19501,N_18766);
or UO_700 (O_700,N_22578,N_19045);
nand UO_701 (O_701,N_21567,N_23684);
or UO_702 (O_702,N_22562,N_24033);
xnor UO_703 (O_703,N_23887,N_22774);
and UO_704 (O_704,N_24698,N_23696);
xnor UO_705 (O_705,N_19243,N_22748);
or UO_706 (O_706,N_24887,N_20553);
nand UO_707 (O_707,N_19536,N_24961);
and UO_708 (O_708,N_20958,N_21041);
nor UO_709 (O_709,N_22369,N_23413);
and UO_710 (O_710,N_22437,N_23319);
nor UO_711 (O_711,N_20349,N_24654);
nor UO_712 (O_712,N_21428,N_22583);
nor UO_713 (O_713,N_19412,N_19401);
nor UO_714 (O_714,N_23719,N_24213);
xor UO_715 (O_715,N_21025,N_24139);
xor UO_716 (O_716,N_24062,N_23266);
and UO_717 (O_717,N_21963,N_22760);
nand UO_718 (O_718,N_24862,N_20265);
nor UO_719 (O_719,N_22035,N_22674);
and UO_720 (O_720,N_18754,N_22869);
or UO_721 (O_721,N_20591,N_20818);
nor UO_722 (O_722,N_24714,N_22897);
nor UO_723 (O_723,N_19305,N_21761);
nor UO_724 (O_724,N_20567,N_23418);
nor UO_725 (O_725,N_21704,N_24293);
or UO_726 (O_726,N_23043,N_22661);
or UO_727 (O_727,N_18762,N_24373);
nor UO_728 (O_728,N_23971,N_20376);
nor UO_729 (O_729,N_22209,N_24991);
nand UO_730 (O_730,N_23233,N_19259);
and UO_731 (O_731,N_23187,N_21294);
nor UO_732 (O_732,N_24378,N_21378);
nor UO_733 (O_733,N_24000,N_23676);
and UO_734 (O_734,N_19041,N_24268);
nand UO_735 (O_735,N_22731,N_20888);
or UO_736 (O_736,N_24758,N_21410);
and UO_737 (O_737,N_20008,N_22847);
nand UO_738 (O_738,N_22195,N_21709);
nand UO_739 (O_739,N_22491,N_19880);
or UO_740 (O_740,N_22356,N_21252);
nand UO_741 (O_741,N_19963,N_18933);
nor UO_742 (O_742,N_20368,N_21136);
nand UO_743 (O_743,N_19149,N_24425);
nor UO_744 (O_744,N_20823,N_21400);
or UO_745 (O_745,N_22032,N_21552);
and UO_746 (O_746,N_23275,N_19017);
nor UO_747 (O_747,N_20048,N_21765);
nor UO_748 (O_748,N_20585,N_18927);
and UO_749 (O_749,N_21497,N_19380);
or UO_750 (O_750,N_21038,N_20992);
nor UO_751 (O_751,N_19460,N_20086);
nor UO_752 (O_752,N_23212,N_19110);
nor UO_753 (O_753,N_24867,N_20515);
or UO_754 (O_754,N_21331,N_22332);
or UO_755 (O_755,N_24989,N_21414);
or UO_756 (O_756,N_23465,N_24660);
xor UO_757 (O_757,N_23411,N_21033);
or UO_758 (O_758,N_22096,N_23564);
nand UO_759 (O_759,N_19938,N_24755);
or UO_760 (O_760,N_23031,N_22576);
and UO_761 (O_761,N_21269,N_24937);
or UO_762 (O_762,N_20058,N_24232);
and UO_763 (O_763,N_19504,N_22479);
nand UO_764 (O_764,N_24389,N_19949);
xnor UO_765 (O_765,N_19381,N_21084);
nor UO_766 (O_766,N_24112,N_20551);
nand UO_767 (O_767,N_23643,N_23125);
nor UO_768 (O_768,N_23787,N_23496);
nor UO_769 (O_769,N_21814,N_22230);
nand UO_770 (O_770,N_22381,N_24280);
and UO_771 (O_771,N_22458,N_19588);
nor UO_772 (O_772,N_23897,N_18903);
nor UO_773 (O_773,N_22613,N_19889);
or UO_774 (O_774,N_18814,N_21675);
nor UO_775 (O_775,N_20443,N_22746);
and UO_776 (O_776,N_20498,N_19662);
nor UO_777 (O_777,N_23084,N_24976);
nand UO_778 (O_778,N_24890,N_24394);
nor UO_779 (O_779,N_19595,N_19224);
or UO_780 (O_780,N_24271,N_19197);
or UO_781 (O_781,N_22044,N_23571);
and UO_782 (O_782,N_24218,N_23664);
or UO_783 (O_783,N_23838,N_19150);
nand UO_784 (O_784,N_23458,N_23734);
xnor UO_785 (O_785,N_19047,N_21514);
or UO_786 (O_786,N_21840,N_19722);
nand UO_787 (O_787,N_23862,N_22573);
and UO_788 (O_788,N_23863,N_20353);
nor UO_789 (O_789,N_24956,N_24821);
xnor UO_790 (O_790,N_19928,N_22968);
xnor UO_791 (O_791,N_20215,N_19846);
nand UO_792 (O_792,N_18989,N_23725);
nand UO_793 (O_793,N_20773,N_19023);
and UO_794 (O_794,N_22640,N_24151);
nor UO_795 (O_795,N_22901,N_20936);
nand UO_796 (O_796,N_24931,N_21792);
and UO_797 (O_797,N_19998,N_21455);
and UO_798 (O_798,N_19082,N_24365);
xnor UO_799 (O_799,N_21629,N_24724);
and UO_800 (O_800,N_19940,N_20125);
and UO_801 (O_801,N_19921,N_23493);
or UO_802 (O_802,N_23982,N_20587);
or UO_803 (O_803,N_24739,N_24651);
nor UO_804 (O_804,N_21356,N_19842);
and UO_805 (O_805,N_19698,N_23914);
xnor UO_806 (O_806,N_20882,N_23942);
nor UO_807 (O_807,N_19148,N_22128);
and UO_808 (O_808,N_21787,N_24080);
nand UO_809 (O_809,N_24089,N_20171);
xor UO_810 (O_810,N_24907,N_22936);
or UO_811 (O_811,N_22318,N_19637);
nand UO_812 (O_812,N_24819,N_22418);
and UO_813 (O_813,N_23341,N_19492);
or UO_814 (O_814,N_24282,N_21697);
xnor UO_815 (O_815,N_23284,N_24409);
nor UO_816 (O_816,N_21981,N_20578);
nand UO_817 (O_817,N_21602,N_24345);
and UO_818 (O_818,N_20044,N_23846);
nor UO_819 (O_819,N_24665,N_21397);
nor UO_820 (O_820,N_22821,N_21692);
nor UO_821 (O_821,N_20151,N_24229);
or UO_822 (O_822,N_20506,N_22240);
or UO_823 (O_823,N_24191,N_21147);
or UO_824 (O_824,N_24571,N_20116);
nand UO_825 (O_825,N_24893,N_23146);
nor UO_826 (O_826,N_21318,N_24716);
or UO_827 (O_827,N_22982,N_22953);
or UO_828 (O_828,N_24393,N_24026);
or UO_829 (O_829,N_24405,N_23825);
or UO_830 (O_830,N_24430,N_22210);
nor UO_831 (O_831,N_21591,N_23650);
and UO_832 (O_832,N_23119,N_21702);
nand UO_833 (O_833,N_22168,N_21952);
and UO_834 (O_834,N_24145,N_23326);
xor UO_835 (O_835,N_20045,N_24095);
nor UO_836 (O_836,N_21301,N_23586);
xnor UO_837 (O_837,N_22000,N_19442);
and UO_838 (O_838,N_24537,N_19841);
nor UO_839 (O_839,N_20791,N_20261);
nor UO_840 (O_840,N_22038,N_19019);
and UO_841 (O_841,N_23698,N_23724);
or UO_842 (O_842,N_24563,N_19621);
xor UO_843 (O_843,N_21040,N_23066);
xnor UO_844 (O_844,N_21928,N_22300);
nand UO_845 (O_845,N_21919,N_24344);
or UO_846 (O_846,N_24153,N_20022);
nand UO_847 (O_847,N_21330,N_24746);
xor UO_848 (O_848,N_20152,N_22271);
nor UO_849 (O_849,N_22610,N_23648);
or UO_850 (O_850,N_22299,N_20351);
or UO_851 (O_851,N_24857,N_22207);
or UO_852 (O_852,N_20808,N_22725);
nor UO_853 (O_853,N_20779,N_23193);
and UO_854 (O_854,N_21706,N_24552);
nand UO_855 (O_855,N_20114,N_24718);
nand UO_856 (O_856,N_22080,N_21797);
and UO_857 (O_857,N_19677,N_21361);
or UO_858 (O_858,N_24968,N_20467);
xnor UO_859 (O_859,N_21902,N_20604);
xor UO_860 (O_860,N_24658,N_20315);
nor UO_861 (O_861,N_23011,N_24599);
xor UO_862 (O_862,N_20539,N_21822);
or UO_863 (O_863,N_23106,N_24542);
xnor UO_864 (O_864,N_24243,N_22114);
nand UO_865 (O_865,N_18985,N_19398);
and UO_866 (O_866,N_23997,N_21539);
nor UO_867 (O_867,N_23114,N_20776);
nand UO_868 (O_868,N_21546,N_19579);
xnor UO_869 (O_869,N_22797,N_21422);
nand UO_870 (O_870,N_19195,N_19180);
xor UO_871 (O_871,N_21677,N_20359);
and UO_872 (O_872,N_23604,N_24418);
nand UO_873 (O_873,N_22617,N_21395);
and UO_874 (O_874,N_24279,N_23072);
xnor UO_875 (O_875,N_24813,N_23975);
nand UO_876 (O_876,N_20876,N_24053);
nor UO_877 (O_877,N_20999,N_21522);
nor UO_878 (O_878,N_21918,N_21894);
and UO_879 (O_879,N_23056,N_21327);
xor UO_880 (O_880,N_20490,N_19105);
xnor UO_881 (O_881,N_21433,N_19146);
nor UO_882 (O_882,N_23654,N_22815);
or UO_883 (O_883,N_20436,N_22867);
xnor UO_884 (O_884,N_20168,N_20835);
and UO_885 (O_885,N_23926,N_22047);
and UO_886 (O_886,N_23715,N_24038);
nor UO_887 (O_887,N_22376,N_18991);
nand UO_888 (O_888,N_22868,N_21238);
xnor UO_889 (O_889,N_24847,N_24780);
nand UO_890 (O_890,N_21835,N_21873);
or UO_891 (O_891,N_23933,N_24269);
xor UO_892 (O_892,N_21364,N_24212);
or UO_893 (O_893,N_21595,N_22519);
nor UO_894 (O_894,N_21494,N_22435);
and UO_895 (O_895,N_22078,N_20613);
and UO_896 (O_896,N_19052,N_24919);
or UO_897 (O_897,N_23918,N_24507);
nor UO_898 (O_898,N_21251,N_23182);
nand UO_899 (O_899,N_23378,N_21181);
xnor UO_900 (O_900,N_23047,N_24065);
nor UO_901 (O_901,N_24137,N_21425);
nor UO_902 (O_902,N_24916,N_21622);
nand UO_903 (O_903,N_19997,N_18850);
nor UO_904 (O_904,N_20534,N_21543);
xnor UO_905 (O_905,N_24925,N_19236);
nor UO_906 (O_906,N_24999,N_20885);
or UO_907 (O_907,N_24167,N_23065);
and UO_908 (O_908,N_23543,N_23350);
xnor UO_909 (O_909,N_20503,N_21626);
nor UO_910 (O_910,N_19371,N_22455);
and UO_911 (O_911,N_19977,N_24142);
and UO_912 (O_912,N_24278,N_21755);
and UO_913 (O_913,N_19566,N_21810);
nor UO_914 (O_914,N_19434,N_22290);
xnor UO_915 (O_915,N_23726,N_20243);
xnor UO_916 (O_916,N_18889,N_21399);
nor UO_917 (O_917,N_22135,N_20841);
and UO_918 (O_918,N_22687,N_21550);
xnor UO_919 (O_919,N_20416,N_20356);
xor UO_920 (O_920,N_22673,N_19003);
and UO_921 (O_921,N_23178,N_24307);
and UO_922 (O_922,N_24777,N_22339);
and UO_923 (O_923,N_24653,N_19223);
nor UO_924 (O_924,N_22097,N_23960);
xnor UO_925 (O_925,N_21415,N_21689);
nor UO_926 (O_926,N_19876,N_20850);
and UO_927 (O_927,N_20813,N_21230);
nor UO_928 (O_928,N_23695,N_24143);
and UO_929 (O_929,N_24941,N_23064);
xnor UO_930 (O_930,N_19153,N_23181);
or UO_931 (O_931,N_22463,N_23196);
or UO_932 (O_932,N_22526,N_23375);
nor UO_933 (O_933,N_19587,N_23561);
and UO_934 (O_934,N_22677,N_20889);
xor UO_935 (O_935,N_22695,N_21027);
nor UO_936 (O_936,N_23051,N_19248);
xor UO_937 (O_937,N_24206,N_23781);
and UO_938 (O_938,N_24055,N_23866);
nand UO_939 (O_939,N_23438,N_19516);
or UO_940 (O_940,N_23645,N_19392);
nand UO_941 (O_941,N_23905,N_19732);
nor UO_942 (O_942,N_24969,N_21288);
nand UO_943 (O_943,N_22654,N_19338);
xnor UO_944 (O_944,N_19253,N_23790);
xor UO_945 (O_945,N_19929,N_19497);
nor UO_946 (O_946,N_24119,N_18819);
and UO_947 (O_947,N_22900,N_19982);
xnor UO_948 (O_948,N_24864,N_20375);
and UO_949 (O_949,N_20512,N_24640);
xnor UO_950 (O_950,N_19207,N_22218);
xnor UO_951 (O_951,N_24193,N_19630);
xor UO_952 (O_952,N_22053,N_24508);
nor UO_953 (O_953,N_19717,N_19374);
or UO_954 (O_954,N_22132,N_23330);
nor UO_955 (O_955,N_20309,N_20730);
xor UO_956 (O_956,N_22362,N_20704);
and UO_957 (O_957,N_21799,N_21303);
and UO_958 (O_958,N_23216,N_24855);
and UO_959 (O_959,N_20691,N_24785);
nor UO_960 (O_960,N_20806,N_24160);
nor UO_961 (O_961,N_21652,N_21828);
xnor UO_962 (O_962,N_20354,N_23647);
nor UO_963 (O_963,N_24403,N_24967);
and UO_964 (O_964,N_20605,N_23222);
nor UO_965 (O_965,N_22833,N_22747);
and UO_966 (O_966,N_22287,N_23410);
nor UO_967 (O_967,N_21435,N_22546);
xor UO_968 (O_968,N_23269,N_19576);
nand UO_969 (O_969,N_23213,N_21490);
nor UO_970 (O_970,N_20372,N_23688);
and UO_971 (O_971,N_19360,N_20397);
and UO_972 (O_972,N_24124,N_24545);
or UO_973 (O_973,N_23891,N_23523);
and UO_974 (O_974,N_21468,N_20169);
nand UO_975 (O_975,N_19074,N_19265);
nor UO_976 (O_976,N_19445,N_23323);
nor UO_977 (O_977,N_22243,N_21777);
nor UO_978 (O_978,N_22793,N_18943);
nor UO_979 (O_979,N_20387,N_22572);
nand UO_980 (O_980,N_20698,N_20856);
or UO_981 (O_981,N_23562,N_19385);
nand UO_982 (O_982,N_23721,N_19535);
xnor UO_983 (O_983,N_21962,N_24974);
and UO_984 (O_984,N_20521,N_20967);
or UO_985 (O_985,N_21370,N_20021);
and UO_986 (O_986,N_21844,N_23628);
and UO_987 (O_987,N_21412,N_24672);
and UO_988 (O_988,N_24214,N_19119);
and UO_989 (O_989,N_18831,N_19573);
or UO_990 (O_990,N_23764,N_19502);
and UO_991 (O_991,N_20165,N_21794);
or UO_992 (O_992,N_20953,N_19315);
and UO_993 (O_993,N_19143,N_23112);
nor UO_994 (O_994,N_19213,N_21022);
nor UO_995 (O_995,N_19743,N_20968);
nand UO_996 (O_996,N_20258,N_21983);
or UO_997 (O_997,N_20084,N_22380);
and UO_998 (O_998,N_24318,N_22750);
nand UO_999 (O_999,N_24675,N_24261);
and UO_1000 (O_1000,N_24802,N_21358);
and UO_1001 (O_1001,N_19778,N_24379);
xor UO_1002 (O_1002,N_19151,N_19509);
nor UO_1003 (O_1003,N_23640,N_22312);
xnor UO_1004 (O_1004,N_24426,N_22532);
nor UO_1005 (O_1005,N_23965,N_22224);
xor UO_1006 (O_1006,N_21586,N_21687);
or UO_1007 (O_1007,N_24643,N_23533);
or UO_1008 (O_1008,N_22969,N_23538);
nand UO_1009 (O_1009,N_24314,N_24814);
or UO_1010 (O_1010,N_22060,N_23005);
and UO_1011 (O_1011,N_21134,N_24450);
and UO_1012 (O_1012,N_21929,N_20829);
xor UO_1013 (O_1013,N_23565,N_24313);
xnor UO_1014 (O_1014,N_22657,N_20227);
xor UO_1015 (O_1015,N_21931,N_22043);
nor UO_1016 (O_1016,N_20344,N_22521);
nor UO_1017 (O_1017,N_21020,N_20582);
nand UO_1018 (O_1018,N_22866,N_21515);
nand UO_1019 (O_1019,N_20024,N_23567);
or UO_1020 (O_1020,N_23337,N_19030);
xnor UO_1021 (O_1021,N_20292,N_22678);
or UO_1022 (O_1022,N_20098,N_22501);
or UO_1023 (O_1023,N_23422,N_21759);
nor UO_1024 (O_1024,N_22594,N_22008);
xor UO_1025 (O_1025,N_20213,N_22127);
nor UO_1026 (O_1026,N_23030,N_18870);
nor UO_1027 (O_1027,N_22320,N_20638);
and UO_1028 (O_1028,N_24377,N_19574);
or UO_1029 (O_1029,N_24004,N_21477);
nand UO_1030 (O_1030,N_21151,N_20666);
xnor UO_1031 (O_1031,N_23509,N_20484);
and UO_1032 (O_1032,N_19890,N_22222);
or UO_1033 (O_1033,N_24486,N_22782);
nand UO_1034 (O_1034,N_20144,N_21679);
nand UO_1035 (O_1035,N_24493,N_23025);
xor UO_1036 (O_1036,N_20109,N_20986);
and UO_1037 (O_1037,N_19581,N_23991);
nor UO_1038 (O_1038,N_20137,N_22593);
nor UO_1039 (O_1039,N_20495,N_24808);
or UO_1040 (O_1040,N_23858,N_23613);
and UO_1041 (O_1041,N_20974,N_20736);
and UO_1042 (O_1042,N_19884,N_24983);
nor UO_1043 (O_1043,N_20943,N_23936);
and UO_1044 (O_1044,N_23241,N_18799);
xor UO_1045 (O_1045,N_22971,N_24577);
xnor UO_1046 (O_1046,N_20150,N_24509);
and UO_1047 (O_1047,N_23678,N_20700);
and UO_1048 (O_1048,N_21182,N_22966);
nand UO_1049 (O_1049,N_21811,N_19591);
and UO_1050 (O_1050,N_19820,N_20026);
nand UO_1051 (O_1051,N_18794,N_21905);
xor UO_1052 (O_1052,N_23129,N_20068);
or UO_1053 (O_1053,N_19246,N_21212);
and UO_1054 (O_1054,N_23723,N_24738);
nand UO_1055 (O_1055,N_24533,N_20472);
xnor UO_1056 (O_1056,N_24498,N_20302);
or UO_1057 (O_1057,N_19489,N_20816);
and UO_1058 (O_1058,N_19586,N_21616);
nor UO_1059 (O_1059,N_21711,N_24561);
xnor UO_1060 (O_1060,N_24960,N_24987);
or UO_1061 (O_1061,N_23456,N_21044);
or UO_1062 (O_1062,N_24949,N_18869);
and UO_1063 (O_1063,N_22401,N_21693);
nor UO_1064 (O_1064,N_21304,N_24072);
nand UO_1065 (O_1065,N_24811,N_21752);
nor UO_1066 (O_1066,N_20870,N_23328);
nor UO_1067 (O_1067,N_21059,N_21231);
or UO_1068 (O_1068,N_24621,N_24782);
nor UO_1069 (O_1069,N_22323,N_20189);
or UO_1070 (O_1070,N_19523,N_23393);
xnor UO_1071 (O_1071,N_23767,N_18988);
or UO_1072 (O_1072,N_20329,N_24086);
or UO_1073 (O_1073,N_22791,N_19135);
or UO_1074 (O_1074,N_20601,N_20160);
nand UO_1075 (O_1075,N_19690,N_20879);
and UO_1076 (O_1076,N_19383,N_20491);
xor UO_1077 (O_1077,N_22700,N_23874);
xor UO_1078 (O_1078,N_21352,N_20971);
xor UO_1079 (O_1079,N_18983,N_24012);
and UO_1080 (O_1080,N_22516,N_20234);
nand UO_1081 (O_1081,N_23607,N_20932);
xnor UO_1082 (O_1082,N_24932,N_19122);
nor UO_1083 (O_1083,N_19932,N_22250);
or UO_1084 (O_1084,N_22876,N_19831);
nor UO_1085 (O_1085,N_23305,N_20648);
nand UO_1086 (O_1086,N_19355,N_24141);
nand UO_1087 (O_1087,N_23619,N_22697);
xnor UO_1088 (O_1088,N_22924,N_20456);
nand UO_1089 (O_1089,N_19351,N_23126);
nor UO_1090 (O_1090,N_22637,N_19410);
or UO_1091 (O_1091,N_23677,N_24263);
nand UO_1092 (O_1092,N_22837,N_19421);
nand UO_1093 (O_1093,N_19925,N_20641);
nand UO_1094 (O_1094,N_21295,N_20848);
nor UO_1095 (O_1095,N_22884,N_22061);
nand UO_1096 (O_1096,N_23229,N_20221);
or UO_1097 (O_1097,N_21715,N_20709);
xnor UO_1098 (O_1098,N_22649,N_24348);
or UO_1099 (O_1099,N_20130,N_22365);
or UO_1100 (O_1100,N_24368,N_19483);
nor UO_1101 (O_1101,N_19251,N_20238);
nor UO_1102 (O_1102,N_24025,N_23217);
or UO_1103 (O_1103,N_19835,N_21159);
xnor UO_1104 (O_1104,N_23017,N_20462);
nand UO_1105 (O_1105,N_19173,N_22877);
xnor UO_1106 (O_1106,N_22951,N_24691);
nor UO_1107 (O_1107,N_21557,N_19264);
nand UO_1108 (O_1108,N_22263,N_19901);
or UO_1109 (O_1109,N_20669,N_19601);
and UO_1110 (O_1110,N_19137,N_20861);
or UO_1111 (O_1111,N_21656,N_20049);
and UO_1112 (O_1112,N_21941,N_21302);
or UO_1113 (O_1113,N_20295,N_19865);
nor UO_1114 (O_1114,N_22022,N_24281);
xor UO_1115 (O_1115,N_24291,N_21795);
or UO_1116 (O_1116,N_23737,N_23860);
or UO_1117 (O_1117,N_21260,N_23408);
or UO_1118 (O_1118,N_23177,N_22829);
and UO_1119 (O_1119,N_19768,N_24071);
or UO_1120 (O_1120,N_24132,N_23861);
xor UO_1121 (O_1121,N_20010,N_23799);
and UO_1122 (O_1122,N_24657,N_20294);
xor UO_1123 (O_1123,N_24562,N_24341);
or UO_1124 (O_1124,N_22865,N_23488);
nor UO_1125 (O_1125,N_21448,N_23809);
nand UO_1126 (O_1126,N_22559,N_19028);
nand UO_1127 (O_1127,N_23898,N_23109);
nand UO_1128 (O_1128,N_20016,N_20052);
nor UO_1129 (O_1129,N_24635,N_21137);
or UO_1130 (O_1130,N_18769,N_22013);
or UO_1131 (O_1131,N_22507,N_19897);
nand UO_1132 (O_1132,N_24310,N_22595);
or UO_1133 (O_1133,N_19955,N_23405);
nand UO_1134 (O_1134,N_20431,N_21620);
and UO_1135 (O_1135,N_22336,N_24667);
and UO_1136 (O_1136,N_22375,N_24518);
and UO_1137 (O_1137,N_24911,N_23082);
xor UO_1138 (O_1138,N_24434,N_21526);
and UO_1139 (O_1139,N_18844,N_24772);
nor UO_1140 (O_1140,N_19803,N_20563);
and UO_1141 (O_1141,N_19912,N_24458);
and UO_1142 (O_1142,N_22204,N_20985);
nor UO_1143 (O_1143,N_23425,N_20361);
xnor UO_1144 (O_1144,N_19896,N_23259);
nand UO_1145 (O_1145,N_19104,N_21851);
nand UO_1146 (O_1146,N_22520,N_24564);
and UO_1147 (O_1147,N_23432,N_24963);
nand UO_1148 (O_1148,N_24866,N_19795);
xor UO_1149 (O_1149,N_20113,N_22321);
nor UO_1150 (O_1150,N_20352,N_23760);
or UO_1151 (O_1151,N_22301,N_19359);
nor UO_1152 (O_1152,N_19761,N_23535);
or UO_1153 (O_1153,N_24433,N_21733);
xnor UO_1154 (O_1154,N_20222,N_21747);
and UO_1155 (O_1155,N_22533,N_20104);
xor UO_1156 (O_1156,N_19632,N_21807);
nor UO_1157 (O_1157,N_19394,N_24189);
nand UO_1158 (O_1158,N_21245,N_21275);
xor UO_1159 (O_1159,N_18892,N_23792);
or UO_1160 (O_1160,N_21646,N_21885);
xnor UO_1161 (O_1161,N_22198,N_23039);
xor UO_1162 (O_1162,N_23644,N_22727);
and UO_1163 (O_1163,N_19021,N_22421);
xor UO_1164 (O_1164,N_20518,N_24957);
and UO_1165 (O_1165,N_24896,N_23188);
or UO_1166 (O_1166,N_22171,N_22408);
or UO_1167 (O_1167,N_21185,N_20030);
or UO_1168 (O_1168,N_20755,N_21973);
xnor UO_1169 (O_1169,N_23950,N_24168);
xnor UO_1170 (O_1170,N_19117,N_23622);
nand UO_1171 (O_1171,N_24944,N_19431);
nand UO_1172 (O_1172,N_24094,N_19312);
nand UO_1173 (O_1173,N_22550,N_20963);
or UO_1174 (O_1174,N_19084,N_22555);
and UO_1175 (O_1175,N_21464,N_19531);
and UO_1176 (O_1176,N_21009,N_24305);
nor UO_1177 (O_1177,N_22902,N_23603);
and UO_1178 (O_1178,N_23621,N_20649);
and UO_1179 (O_1179,N_21392,N_19731);
xor UO_1180 (O_1180,N_19356,N_19794);
nor UO_1181 (O_1181,N_22117,N_23808);
or UO_1182 (O_1182,N_20975,N_21753);
or UO_1183 (O_1183,N_19855,N_19441);
nor UO_1184 (O_1184,N_20830,N_19088);
nand UO_1185 (O_1185,N_19282,N_21805);
nor UO_1186 (O_1186,N_21574,N_21045);
and UO_1187 (O_1187,N_24300,N_24467);
nor UO_1188 (O_1188,N_23394,N_22347);
and UO_1189 (O_1189,N_20254,N_23584);
nor UO_1190 (O_1190,N_24699,N_19926);
and UO_1191 (O_1191,N_20009,N_21441);
xnor UO_1192 (O_1192,N_21350,N_20145);
nor UO_1193 (O_1193,N_22962,N_19715);
and UO_1194 (O_1194,N_23560,N_23203);
and UO_1195 (O_1195,N_20657,N_21098);
and UO_1196 (O_1196,N_19764,N_21989);
and UO_1197 (O_1197,N_21634,N_23122);
nand UO_1198 (O_1198,N_23901,N_20631);
xnor UO_1199 (O_1199,N_24164,N_23287);
and UO_1200 (O_1200,N_22120,N_24309);
xnor UO_1201 (O_1201,N_24088,N_20530);
nor UO_1202 (O_1202,N_21021,N_23334);
xnor UO_1203 (O_1203,N_19886,N_22950);
nand UO_1204 (O_1204,N_20983,N_24194);
nor UO_1205 (O_1205,N_19721,N_18775);
nor UO_1206 (O_1206,N_19471,N_20038);
xor UO_1207 (O_1207,N_24877,N_24452);
nand UO_1208 (O_1208,N_19271,N_23077);
nor UO_1209 (O_1209,N_24107,N_19861);
xnor UO_1210 (O_1210,N_24487,N_20997);
nand UO_1211 (O_1211,N_21849,N_19059);
or UO_1212 (O_1212,N_23073,N_22415);
nor UO_1213 (O_1213,N_20192,N_24594);
nor UO_1214 (O_1214,N_19958,N_21621);
nor UO_1215 (O_1215,N_24742,N_19219);
and UO_1216 (O_1216,N_19132,N_24287);
nand UO_1217 (O_1217,N_22587,N_24538);
and UO_1218 (O_1218,N_24536,N_20180);
and UO_1219 (O_1219,N_24836,N_18849);
xnor UO_1220 (O_1220,N_19318,N_24203);
and UO_1221 (O_1221,N_23293,N_23902);
and UO_1222 (O_1222,N_20328,N_23102);
xnor UO_1223 (O_1223,N_21161,N_19856);
xnor UO_1224 (O_1224,N_19530,N_19450);
or UO_1225 (O_1225,N_23867,N_23028);
or UO_1226 (O_1226,N_18897,N_20731);
xnor UO_1227 (O_1227,N_19796,N_22431);
xor UO_1228 (O_1228,N_19277,N_21803);
nand UO_1229 (O_1229,N_19093,N_23821);
xnor UO_1230 (O_1230,N_21884,N_19755);
xnor UO_1231 (O_1231,N_23020,N_22148);
nor UO_1232 (O_1232,N_22488,N_19288);
nand UO_1233 (O_1233,N_20362,N_22548);
xnor UO_1234 (O_1234,N_24638,N_23903);
or UO_1235 (O_1235,N_23768,N_22799);
and UO_1236 (O_1236,N_21250,N_23086);
and UO_1237 (O_1237,N_23819,N_20590);
and UO_1238 (O_1238,N_20083,N_18871);
or UO_1239 (O_1239,N_24574,N_21986);
and UO_1240 (O_1240,N_21613,N_19763);
or UO_1241 (O_1241,N_23386,N_24682);
xor UO_1242 (O_1242,N_24022,N_21337);
nand UO_1243 (O_1243,N_20508,N_20979);
nor UO_1244 (O_1244,N_22251,N_19006);
or UO_1245 (O_1245,N_21725,N_24593);
xor UO_1246 (O_1246,N_24492,N_20041);
nand UO_1247 (O_1247,N_20136,N_22994);
nand UO_1248 (O_1248,N_20319,N_23018);
or UO_1249 (O_1249,N_24069,N_20760);
nor UO_1250 (O_1250,N_22943,N_24852);
or UO_1251 (O_1251,N_19834,N_19425);
and UO_1252 (O_1252,N_21542,N_20394);
nand UO_1253 (O_1253,N_23968,N_21061);
xor UO_1254 (O_1254,N_19405,N_19233);
and UO_1255 (O_1255,N_18947,N_19476);
nor UO_1256 (O_1256,N_21967,N_19482);
xnor UO_1257 (O_1257,N_23554,N_20475);
and UO_1258 (O_1258,N_18861,N_24419);
nand UO_1259 (O_1259,N_23208,N_23665);
xnor UO_1260 (O_1260,N_24863,N_22211);
nand UO_1261 (O_1261,N_24267,N_24042);
xor UO_1262 (O_1262,N_19918,N_24639);
nand UO_1263 (O_1263,N_21043,N_23580);
and UO_1264 (O_1264,N_23801,N_22945);
nand UO_1265 (O_1265,N_18906,N_24992);
or UO_1266 (O_1266,N_24962,N_22527);
nand UO_1267 (O_1267,N_22857,N_19959);
and UO_1268 (O_1268,N_19609,N_21450);
and UO_1269 (O_1269,N_20558,N_22425);
or UO_1270 (O_1270,N_22536,N_22663);
xnor UO_1271 (O_1271,N_23757,N_22856);
and UO_1272 (O_1272,N_22236,N_23168);
nand UO_1273 (O_1273,N_23412,N_24501);
nand UO_1274 (O_1274,N_24136,N_22011);
or UO_1275 (O_1275,N_19649,N_21290);
nand UO_1276 (O_1276,N_23536,N_20334);
and UO_1277 (O_1277,N_24764,N_19479);
nor UO_1278 (O_1278,N_20739,N_20434);
or UO_1279 (O_1279,N_22057,N_21934);
nor UO_1280 (O_1280,N_21097,N_24816);
nor UO_1281 (O_1281,N_19541,N_23352);
and UO_1282 (O_1282,N_20314,N_20694);
nor UO_1283 (O_1283,N_23992,N_22122);
or UO_1284 (O_1284,N_18778,N_24540);
nand UO_1285 (O_1285,N_24891,N_19639);
and UO_1286 (O_1286,N_22429,N_23804);
nand UO_1287 (O_1287,N_19470,N_22768);
nor UO_1288 (O_1288,N_22588,N_20811);
and UO_1289 (O_1289,N_23716,N_21580);
nor UO_1290 (O_1290,N_24820,N_23659);
nor UO_1291 (O_1291,N_21896,N_24411);
nor UO_1292 (O_1292,N_22806,N_24422);
or UO_1293 (O_1293,N_20922,N_23074);
xnor UO_1294 (O_1294,N_24530,N_18752);
or UO_1295 (O_1295,N_22718,N_20651);
nor UO_1296 (O_1296,N_20358,N_24825);
nor UO_1297 (O_1297,N_22457,N_23433);
nor UO_1298 (O_1298,N_24655,N_22840);
xnor UO_1299 (O_1299,N_22179,N_20858);
and UO_1300 (O_1300,N_22767,N_20080);
xnor UO_1301 (O_1301,N_23170,N_23779);
nor UO_1302 (O_1302,N_18950,N_24497);
and UO_1303 (O_1303,N_21891,N_19705);
and UO_1304 (O_1304,N_19049,N_19071);
nor UO_1305 (O_1305,N_24018,N_21639);
nand UO_1306 (O_1306,N_22273,N_19145);
xnor UO_1307 (O_1307,N_21439,N_23788);
xnor UO_1308 (O_1308,N_20560,N_21085);
xnor UO_1309 (O_1309,N_21320,N_22354);
or UO_1310 (O_1310,N_19245,N_23318);
nand UO_1311 (O_1311,N_19854,N_19610);
or UO_1312 (O_1312,N_22104,N_21499);
nor UO_1313 (O_1313,N_19099,N_22063);
or UO_1314 (O_1314,N_23298,N_21815);
and UO_1315 (O_1315,N_18839,N_23184);
xnor UO_1316 (O_1316,N_22123,N_22723);
xor UO_1317 (O_1317,N_23637,N_24854);
nor UO_1318 (O_1318,N_24939,N_21259);
or UO_1319 (O_1319,N_20906,N_22955);
nor UO_1320 (O_1320,N_22041,N_22537);
nor UO_1321 (O_1321,N_22015,N_22341);
nor UO_1322 (O_1322,N_23141,N_22069);
nor UO_1323 (O_1323,N_22620,N_22628);
nor UO_1324 (O_1324,N_18994,N_21510);
and UO_1325 (O_1325,N_24273,N_22990);
nor UO_1326 (O_1326,N_19893,N_22075);
or UO_1327 (O_1327,N_19724,N_19883);
nor UO_1328 (O_1328,N_23263,N_20702);
xnor UO_1329 (O_1329,N_23773,N_24784);
nor UO_1330 (O_1330,N_21285,N_21951);
nand UO_1331 (O_1331,N_22894,N_23226);
nand UO_1332 (O_1332,N_22118,N_21869);
and UO_1333 (O_1333,N_24009,N_19735);
xnor UO_1334 (O_1334,N_21483,N_20186);
nand UO_1335 (O_1335,N_24807,N_24350);
xnor UO_1336 (O_1336,N_19456,N_22667);
and UO_1337 (O_1337,N_21454,N_24848);
nand UO_1338 (O_1338,N_24773,N_21713);
and UO_1339 (O_1339,N_21424,N_24506);
xnor UO_1340 (O_1340,N_20004,N_19776);
nand UO_1341 (O_1341,N_22308,N_19070);
nor UO_1342 (O_1342,N_20662,N_19927);
or UO_1343 (O_1343,N_23692,N_18834);
or UO_1344 (O_1344,N_22662,N_21897);
nand UO_1345 (O_1345,N_19634,N_21783);
and UO_1346 (O_1346,N_18929,N_21705);
and UO_1347 (O_1347,N_20767,N_23363);
nand UO_1348 (O_1348,N_22157,N_23494);
nand UO_1349 (O_1349,N_20350,N_22707);
xor UO_1350 (O_1350,N_21597,N_24172);
nor UO_1351 (O_1351,N_21345,N_22785);
nand UO_1352 (O_1352,N_20311,N_20025);
nand UO_1353 (O_1353,N_23192,N_23201);
nand UO_1354 (O_1354,N_24610,N_19034);
or UO_1355 (O_1355,N_24109,N_24116);
xnor UO_1356 (O_1356,N_19163,N_24262);
nor UO_1357 (O_1357,N_19333,N_20862);
nand UO_1358 (O_1358,N_20681,N_24790);
xor UO_1359 (O_1359,N_20420,N_22052);
nand UO_1360 (O_1360,N_23556,N_24876);
xnor UO_1361 (O_1361,N_19115,N_19994);
xnor UO_1362 (O_1362,N_22370,N_19339);
or UO_1363 (O_1363,N_21991,N_22221);
nor UO_1364 (O_1364,N_20365,N_19377);
nor UO_1365 (O_1365,N_21083,N_23476);
or UO_1366 (O_1366,N_24133,N_21065);
nand UO_1367 (O_1367,N_23325,N_21883);
nand UO_1368 (O_1368,N_21072,N_24296);
or UO_1369 (O_1369,N_19748,N_21111);
xor UO_1370 (O_1370,N_20949,N_22871);
and UO_1371 (O_1371,N_20904,N_22447);
xor UO_1372 (O_1372,N_21848,N_20198);
nor UO_1373 (O_1373,N_19257,N_20277);
nor UO_1374 (O_1374,N_20527,N_22017);
xnor UO_1375 (O_1375,N_21661,N_23511);
or UO_1376 (O_1376,N_24728,N_21018);
or UO_1377 (O_1377,N_24329,N_20450);
nand UO_1378 (O_1378,N_20549,N_21710);
xnor UO_1379 (O_1379,N_21852,N_18820);
or UO_1380 (O_1380,N_20821,N_21789);
xnor UO_1381 (O_1381,N_19500,N_24319);
or UO_1382 (O_1382,N_22272,N_24289);
xor UO_1383 (O_1383,N_22732,N_20304);
and UO_1384 (O_1384,N_22149,N_24302);
or UO_1385 (O_1385,N_20487,N_22438);
xor UO_1386 (O_1386,N_22938,N_19540);
nand UO_1387 (O_1387,N_19108,N_22556);
and UO_1388 (O_1388,N_23402,N_24837);
nor UO_1389 (O_1389,N_24468,N_21503);
and UO_1390 (O_1390,N_22812,N_19521);
xor UO_1391 (O_1391,N_20118,N_22084);
nand UO_1392 (O_1392,N_22933,N_21225);
nor UO_1393 (O_1393,N_22095,N_18758);
nor UO_1394 (O_1394,N_22680,N_21776);
nand UO_1395 (O_1395,N_24750,N_23076);
nor UO_1396 (O_1396,N_20095,N_23590);
nor UO_1397 (O_1397,N_21640,N_24446);
or UO_1398 (O_1398,N_19295,N_20429);
or UO_1399 (O_1399,N_23539,N_24851);
nor UO_1400 (O_1400,N_22749,N_19063);
or UO_1401 (O_1401,N_23116,N_24275);
nand UO_1402 (O_1402,N_23906,N_20998);
xnor UO_1403 (O_1403,N_24872,N_24543);
nor UO_1404 (O_1404,N_23075,N_23811);
xor UO_1405 (O_1405,N_21910,N_19427);
nand UO_1406 (O_1406,N_24294,N_19109);
nand UO_1407 (O_1407,N_24834,N_21046);
nor UO_1408 (O_1408,N_24952,N_21589);
xnor UO_1409 (O_1409,N_22033,N_21316);
nand UO_1410 (O_1410,N_19791,N_21845);
nor UO_1411 (O_1411,N_19996,N_22258);
nand UO_1412 (O_1412,N_21419,N_21262);
nor UO_1413 (O_1413,N_22875,N_19331);
nor UO_1414 (O_1414,N_20915,N_23642);
xnor UO_1415 (O_1415,N_20071,N_22100);
or UO_1416 (O_1416,N_22326,N_21000);
xor UO_1417 (O_1417,N_19408,N_18914);
or UO_1418 (O_1418,N_22245,N_24438);
xor UO_1419 (O_1419,N_22515,N_20403);
and UO_1420 (O_1420,N_22831,N_24114);
and UO_1421 (O_1421,N_23939,N_19693);
and UO_1422 (O_1422,N_22671,N_23312);
nand UO_1423 (O_1423,N_24624,N_21299);
xnor UO_1424 (O_1424,N_22484,N_19293);
nor UO_1425 (O_1425,N_24703,N_20903);
or UO_1426 (O_1426,N_19155,N_23490);
and UO_1427 (O_1427,N_22223,N_24710);
or UO_1428 (O_1428,N_22297,N_23829);
xor UO_1429 (O_1429,N_23956,N_23115);
and UO_1430 (O_1430,N_19948,N_21734);
or UO_1431 (O_1431,N_23745,N_23054);
or UO_1432 (O_1432,N_21242,N_20143);
nand UO_1433 (O_1433,N_24709,N_24587);
nand UO_1434 (O_1434,N_20867,N_21612);
or UO_1435 (O_1435,N_23373,N_21988);
and UO_1436 (O_1436,N_21900,N_23855);
nand UO_1437 (O_1437,N_21990,N_24247);
xor UO_1438 (O_1438,N_22554,N_22029);
or UO_1439 (O_1439,N_23671,N_21177);
nand UO_1440 (O_1440,N_20907,N_24324);
nor UO_1441 (O_1441,N_21239,N_21315);
and UO_1442 (O_1442,N_22775,N_19909);
and UO_1443 (O_1443,N_18959,N_21430);
nand UO_1444 (O_1444,N_23843,N_23153);
or UO_1445 (O_1445,N_21413,N_20703);
nand UO_1446 (O_1446,N_19326,N_24187);
or UO_1447 (O_1447,N_19384,N_22303);
nand UO_1448 (O_1448,N_22180,N_23015);
nor UO_1449 (O_1449,N_21671,N_19887);
xnor UO_1450 (O_1450,N_21922,N_22932);
nor UO_1451 (O_1451,N_22254,N_24255);
xor UO_1452 (O_1452,N_23035,N_20317);
nor UO_1453 (O_1453,N_20972,N_22607);
or UO_1454 (O_1454,N_24105,N_20625);
xor UO_1455 (O_1455,N_23910,N_21855);
nand UO_1456 (O_1456,N_19375,N_22269);
xnor UO_1457 (O_1457,N_24977,N_21162);
or UO_1458 (O_1458,N_19158,N_19056);
nor UO_1459 (O_1459,N_21462,N_21067);
nor UO_1460 (O_1460,N_19065,N_22412);
xor UO_1461 (O_1461,N_23013,N_24856);
xnor UO_1462 (O_1462,N_20241,N_22631);
nor UO_1463 (O_1463,N_24586,N_20688);
nor UO_1464 (O_1464,N_21936,N_22241);
and UO_1465 (O_1465,N_23485,N_24364);
nor UO_1466 (O_1466,N_20313,N_23924);
xnor UO_1467 (O_1467,N_24332,N_19391);
nor UO_1468 (O_1468,N_19302,N_23238);
and UO_1469 (O_1469,N_21492,N_20373);
xnor UO_1470 (O_1470,N_24693,N_18963);
nor UO_1471 (O_1471,N_19508,N_23002);
xor UO_1472 (O_1472,N_23058,N_23227);
and UO_1473 (O_1473,N_23569,N_20271);
nand UO_1474 (O_1474,N_22668,N_24295);
xnor UO_1475 (O_1475,N_19133,N_24250);
and UO_1476 (O_1476,N_19704,N_19096);
xor UO_1477 (O_1477,N_21611,N_19089);
or UO_1478 (O_1478,N_20840,N_20865);
nor UO_1479 (O_1479,N_19116,N_24253);
and UO_1480 (O_1480,N_20121,N_21694);
nor UO_1481 (O_1481,N_21344,N_19960);
xnor UO_1482 (O_1482,N_22023,N_22751);
xnor UO_1483 (O_1483,N_21853,N_20627);
xnor UO_1484 (O_1484,N_18984,N_23951);
or UO_1485 (O_1485,N_24179,N_24751);
nand UO_1486 (O_1486,N_21135,N_23281);
or UO_1487 (O_1487,N_22530,N_22608);
nand UO_1488 (O_1488,N_21292,N_19726);
and UO_1489 (O_1489,N_19813,N_21420);
nand UO_1490 (O_1490,N_18837,N_22524);
nand UO_1491 (O_1491,N_21992,N_20256);
or UO_1492 (O_1492,N_23881,N_21081);
nor UO_1493 (O_1493,N_22832,N_24041);
and UO_1494 (O_1494,N_24402,N_19597);
and UO_1495 (O_1495,N_22396,N_23033);
xnor UO_1496 (O_1496,N_21291,N_22818);
nand UO_1497 (O_1497,N_21079,N_21180);
xnor UO_1498 (O_1498,N_22584,N_19274);
or UO_1499 (O_1499,N_24321,N_22430);
nor UO_1500 (O_1500,N_23502,N_22478);
or UO_1501 (O_1501,N_20802,N_23963);
xor UO_1502 (O_1502,N_18845,N_19736);
and UO_1503 (O_1503,N_20312,N_24645);
and UO_1504 (O_1504,N_19304,N_23974);
and UO_1505 (O_1505,N_23666,N_21942);
xor UO_1506 (O_1506,N_18996,N_23911);
or UO_1507 (O_1507,N_20800,N_20911);
xor UO_1508 (O_1508,N_22682,N_22864);
or UO_1509 (O_1509,N_20799,N_21188);
xor UO_1510 (O_1510,N_22202,N_23461);
xor UO_1511 (O_1511,N_22352,N_22565);
or UO_1512 (O_1512,N_19984,N_23751);
nor UO_1513 (O_1513,N_22166,N_23454);
or UO_1514 (O_1514,N_22643,N_23629);
nor UO_1515 (O_1515,N_23500,N_21248);
nand UO_1516 (O_1516,N_24801,N_18776);
xnor UO_1517 (O_1517,N_21654,N_23256);
and UO_1518 (O_1518,N_21300,N_23398);
and UO_1519 (O_1519,N_23739,N_24897);
or UO_1520 (O_1520,N_21956,N_19193);
nand UO_1521 (O_1521,N_19999,N_20196);
nor UO_1522 (O_1522,N_20771,N_20093);
and UO_1523 (O_1523,N_22395,N_21565);
and UO_1524 (O_1524,N_23273,N_19712);
and UO_1525 (O_1525,N_21584,N_19962);
or UO_1526 (O_1526,N_24830,N_24566);
nor UO_1527 (O_1527,N_22470,N_23313);
or UO_1528 (O_1528,N_23728,N_22424);
xor UO_1529 (O_1529,N_24020,N_23770);
xnor UO_1530 (O_1530,N_21227,N_20138);
and UO_1531 (O_1531,N_19916,N_21319);
xnor UO_1532 (O_1532,N_21403,N_22918);
or UO_1533 (O_1533,N_19817,N_23314);
nand UO_1534 (O_1534,N_22575,N_21608);
xor UO_1535 (O_1535,N_24227,N_19797);
xor UO_1536 (O_1536,N_21773,N_21178);
nor UO_1537 (O_1537,N_20586,N_19979);
nand UO_1538 (O_1538,N_22072,N_20005);
nand UO_1539 (O_1539,N_23026,N_21443);
xor UO_1540 (O_1540,N_24972,N_23439);
and UO_1541 (O_1541,N_21915,N_19182);
and UO_1542 (O_1542,N_23540,N_23624);
or UO_1543 (O_1543,N_24771,N_21053);
or UO_1544 (O_1544,N_18803,N_24073);
nand UO_1545 (O_1545,N_23912,N_23332);
xor UO_1546 (O_1546,N_21818,N_19210);
and UO_1547 (O_1547,N_20023,N_24093);
and UO_1548 (O_1548,N_21870,N_23976);
or UO_1549 (O_1549,N_20199,N_24674);
nand UO_1550 (O_1550,N_19040,N_21431);
nand UO_1551 (O_1551,N_22031,N_20786);
xor UO_1552 (O_1552,N_18931,N_23291);
nand UO_1553 (O_1553,N_19372,N_24070);
and UO_1554 (O_1554,N_23841,N_21930);
nand UO_1555 (O_1555,N_23359,N_19237);
or UO_1556 (O_1556,N_19858,N_19239);
nand UO_1557 (O_1557,N_19226,N_24781);
nand UO_1558 (O_1558,N_19179,N_24447);
nand UO_1559 (O_1559,N_24129,N_21858);
and UO_1560 (O_1560,N_22816,N_24195);
xnor UO_1561 (O_1561,N_21877,N_20251);
nor UO_1562 (O_1562,N_19215,N_19991);
nor UO_1563 (O_1563,N_24539,N_19605);
nor UO_1564 (O_1564,N_20619,N_20448);
or UO_1565 (O_1565,N_22167,N_20864);
and UO_1566 (O_1566,N_22796,N_19031);
and UO_1567 (O_1567,N_24459,N_23616);
or UO_1568 (O_1568,N_23694,N_23840);
xor UO_1569 (O_1569,N_20073,N_21396);
nor UO_1570 (O_1570,N_20284,N_21780);
nor UO_1571 (O_1571,N_24888,N_19062);
or UO_1572 (O_1572,N_22685,N_20616);
xnor UO_1573 (O_1573,N_24832,N_22486);
nand UO_1574 (O_1574,N_24113,N_22393);
nor UO_1575 (O_1575,N_22329,N_21437);
xnor UO_1576 (O_1576,N_20103,N_23121);
nand UO_1577 (O_1577,N_22766,N_20064);
and UO_1578 (O_1578,N_19250,N_20128);
nor UO_1579 (O_1579,N_22134,N_19160);
nand UO_1580 (O_1580,N_22183,N_20281);
xnor UO_1581 (O_1581,N_22184,N_19297);
and UO_1582 (O_1582,N_22780,N_19527);
nor UO_1583 (O_1583,N_19354,N_23970);
nor UO_1584 (O_1584,N_21743,N_23120);
nor UO_1585 (O_1585,N_24865,N_24428);
xnor UO_1586 (O_1586,N_19851,N_20804);
and UO_1587 (O_1587,N_23340,N_19965);
and UO_1588 (O_1588,N_23812,N_18757);
or UO_1589 (O_1589,N_24376,N_18910);
and UO_1590 (O_1590,N_20632,N_24753);
nor UO_1591 (O_1591,N_21545,N_22040);
nand UO_1592 (O_1592,N_19298,N_20374);
nand UO_1593 (O_1593,N_22585,N_24796);
nor UO_1594 (O_1594,N_22798,N_22372);
nand UO_1595 (O_1595,N_23376,N_22493);
nand UO_1596 (O_1596,N_18924,N_19092);
xnor UO_1597 (O_1597,N_20656,N_23842);
or UO_1598 (O_1598,N_23234,N_23353);
xor UO_1599 (O_1599,N_24130,N_22842);
nor UO_1600 (O_1600,N_21995,N_20231);
or UO_1601 (O_1601,N_22992,N_22740);
nor UO_1602 (O_1602,N_21663,N_21241);
nand UO_1603 (O_1603,N_18793,N_19490);
or UO_1604 (O_1604,N_22580,N_18856);
nor UO_1605 (O_1605,N_21903,N_20644);
or UO_1606 (O_1606,N_23775,N_21257);
nor UO_1607 (O_1607,N_21863,N_22710);
and UO_1608 (O_1608,N_20072,N_23137);
or UO_1609 (O_1609,N_20039,N_19396);
nor UO_1610 (O_1610,N_23600,N_20253);
nand UO_1611 (O_1611,N_23890,N_23598);
or UO_1612 (O_1612,N_24197,N_23094);
and UO_1613 (O_1613,N_23421,N_19534);
or UO_1614 (O_1614,N_19757,N_22712);
and UO_1615 (O_1615,N_24415,N_21791);
or UO_1616 (O_1616,N_22633,N_20158);
nand UO_1617 (O_1617,N_21573,N_19783);
nand UO_1618 (O_1618,N_23632,N_22635);
nand UO_1619 (O_1619,N_19689,N_24342);
nor UO_1620 (O_1620,N_23096,N_22138);
nand UO_1621 (O_1621,N_19424,N_23451);
nand UO_1622 (O_1622,N_19719,N_23704);
nand UO_1623 (O_1623,N_20571,N_19498);
nor UO_1624 (O_1624,N_21254,N_24276);
xnor UO_1625 (O_1625,N_19709,N_22496);
nand UO_1626 (O_1626,N_19679,N_23711);
xnor UO_1627 (O_1627,N_22590,N_20962);
nand UO_1628 (O_1628,N_22071,N_19057);
or UO_1629 (O_1629,N_23157,N_24335);
and UO_1630 (O_1630,N_20955,N_18940);
and UO_1631 (O_1631,N_23183,N_19167);
xnor UO_1632 (O_1632,N_24039,N_23032);
and UO_1633 (O_1633,N_21306,N_18956);
nand UO_1634 (O_1634,N_22826,N_20507);
nor UO_1635 (O_1635,N_21745,N_19202);
and UO_1636 (O_1636,N_18934,N_23501);
and UO_1637 (O_1637,N_24940,N_24284);
nor UO_1638 (O_1638,N_22028,N_23794);
nand UO_1639 (O_1639,N_21487,N_21377);
or UO_1640 (O_1640,N_24663,N_19526);
xor UO_1641 (O_1641,N_20934,N_19980);
nor UO_1642 (O_1642,N_20445,N_20097);
nand UO_1643 (O_1643,N_21525,N_23735);
nand UO_1644 (O_1644,N_21012,N_24199);
nor UO_1645 (O_1645,N_20564,N_23876);
and UO_1646 (O_1646,N_20187,N_20596);
xnor UO_1647 (O_1647,N_20535,N_20824);
xnor UO_1648 (O_1648,N_23729,N_22417);
or UO_1649 (O_1649,N_22642,N_19827);
and UO_1650 (O_1650,N_21850,N_22357);
nand UO_1651 (O_1651,N_20435,N_23955);
xor UO_1652 (O_1652,N_23420,N_23134);
xor UO_1653 (O_1653,N_23292,N_18955);
nor UO_1654 (O_1654,N_19439,N_23962);
nand UO_1655 (O_1655,N_23434,N_23211);
xnor UO_1656 (O_1656,N_21201,N_24845);
nand UO_1657 (O_1657,N_20769,N_18938);
and UO_1658 (O_1658,N_24569,N_24749);
nor UO_1659 (O_1659,N_21471,N_21328);
and UO_1660 (O_1660,N_22036,N_22315);
or UO_1661 (O_1661,N_22390,N_21449);
nor UO_1662 (O_1662,N_23079,N_20871);
nor UO_1663 (O_1663,N_20088,N_24357);
nor UO_1664 (O_1664,N_23052,N_23311);
xor UO_1665 (O_1665,N_19464,N_20157);
nand UO_1666 (O_1666,N_23255,N_24556);
and UO_1667 (O_1667,N_22843,N_20386);
xor UO_1668 (O_1668,N_23952,N_21442);
and UO_1669 (O_1669,N_24912,N_21528);
xor UO_1670 (O_1670,N_20320,N_20970);
nand UO_1671 (O_1671,N_19039,N_20661);
or UO_1672 (O_1672,N_21635,N_22190);
and UO_1673 (O_1673,N_18753,N_18884);
or UO_1674 (O_1674,N_23080,N_21445);
or UO_1675 (O_1675,N_22985,N_18864);
and UO_1676 (O_1676,N_20282,N_21157);
and UO_1677 (O_1677,N_21609,N_21029);
nand UO_1678 (O_1678,N_23466,N_22105);
nor UO_1679 (O_1679,N_19767,N_20548);
nand UO_1680 (O_1680,N_20298,N_22909);
nand UO_1681 (O_1681,N_20660,N_24705);
or UO_1682 (O_1682,N_20028,N_20714);
xnor UO_1683 (O_1683,N_19583,N_19612);
or UO_1684 (O_1684,N_23844,N_23662);
nor UO_1685 (O_1685,N_21688,N_23477);
nor UO_1686 (O_1686,N_19652,N_23925);
nand UO_1687 (O_1687,N_24833,N_21324);
and UO_1688 (O_1688,N_21229,N_23675);
nand UO_1689 (O_1689,N_23185,N_20954);
nand UO_1690 (O_1690,N_20778,N_24955);
nand UO_1691 (O_1691,N_22121,N_22623);
xnor UO_1692 (O_1692,N_19598,N_20197);
xnor UO_1693 (O_1693,N_23555,N_24152);
or UO_1694 (O_1694,N_23922,N_24104);
and UO_1695 (O_1695,N_24340,N_23069);
or UO_1696 (O_1696,N_23593,N_24443);
nor UO_1697 (O_1697,N_19128,N_24240);
xor UO_1698 (O_1698,N_20675,N_24483);
xnor UO_1699 (O_1699,N_20179,N_22947);
xor UO_1700 (O_1700,N_19700,N_19881);
and UO_1701 (O_1701,N_19181,N_19539);
and UO_1702 (O_1702,N_19168,N_19656);
nor UO_1703 (O_1703,N_21763,N_24512);
and UO_1704 (O_1704,N_19125,N_19785);
nor UO_1705 (O_1705,N_22367,N_19685);
or UO_1706 (O_1706,N_21467,N_21576);
xor UO_1707 (O_1707,N_22928,N_18855);
xnor UO_1708 (O_1708,N_22042,N_18920);
xnor UO_1709 (O_1709,N_21786,N_22039);
and UO_1710 (O_1710,N_24272,N_20664);
or UO_1711 (O_1711,N_22934,N_23321);
nand UO_1712 (O_1712,N_22214,N_24234);
and UO_1713 (O_1713,N_19325,N_20410);
nand UO_1714 (O_1714,N_21145,N_22082);
xnor UO_1715 (O_1715,N_20577,N_22278);
or UO_1716 (O_1716,N_22834,N_22999);
nand UO_1717 (O_1717,N_24973,N_19054);
nand UO_1718 (O_1718,N_19205,N_22482);
xnor UO_1719 (O_1719,N_20684,N_23668);
and UO_1720 (O_1720,N_18868,N_24725);
and UO_1721 (O_1721,N_20630,N_19899);
nor UO_1722 (O_1722,N_24677,N_23150);
and UO_1723 (O_1723,N_22379,N_22225);
nand UO_1724 (O_1724,N_22265,N_19283);
and UO_1725 (O_1725,N_24054,N_24898);
nor UO_1726 (O_1726,N_20828,N_21940);
or UO_1727 (O_1727,N_24333,N_21862);
and UO_1728 (O_1728,N_23878,N_21757);
nand UO_1729 (O_1729,N_22735,N_24994);
or UO_1730 (O_1730,N_20592,N_23504);
xor UO_1731 (O_1731,N_22427,N_23101);
nand UO_1732 (O_1732,N_24414,N_22384);
nor UO_1733 (O_1733,N_19816,N_21270);
nand UO_1734 (O_1734,N_19954,N_20330);
nand UO_1735 (O_1735,N_24683,N_21214);
nand UO_1736 (O_1736,N_22440,N_19815);
or UO_1737 (O_1737,N_19170,N_24208);
nor UO_1738 (O_1738,N_21488,N_21700);
and UO_1739 (O_1739,N_24904,N_21417);
and UO_1740 (O_1740,N_21676,N_20961);
and UO_1741 (O_1741,N_22705,N_22262);
xnor UO_1742 (O_1742,N_22952,N_20200);
or UO_1743 (O_1743,N_23301,N_22733);
or UO_1744 (O_1744,N_24839,N_24058);
nor UO_1745 (O_1745,N_22453,N_20066);
and UO_1746 (O_1746,N_20740,N_19013);
nand UO_1747 (O_1747,N_19078,N_24061);
nor UO_1748 (O_1748,N_20345,N_21684);
nor UO_1749 (O_1749,N_22233,N_24517);
nor UO_1750 (O_1750,N_23894,N_21074);
nand UO_1751 (O_1751,N_23527,N_19287);
xor UO_1752 (O_1752,N_24236,N_19467);
or UO_1753 (O_1753,N_22389,N_19864);
nor UO_1754 (O_1754,N_24209,N_24778);
nand UO_1755 (O_1755,N_22307,N_20370);
or UO_1756 (O_1756,N_24334,N_19699);
xor UO_1757 (O_1757,N_22441,N_18976);
nand UO_1758 (O_1758,N_22020,N_23700);
nor UO_1759 (O_1759,N_23169,N_22255);
and UO_1760 (O_1760,N_19669,N_23994);
or UO_1761 (O_1761,N_24647,N_23215);
xnor UO_1762 (O_1762,N_21655,N_18879);
and UO_1763 (O_1763,N_22500,N_19141);
nand UO_1764 (O_1764,N_24180,N_19600);
nand UO_1765 (O_1765,N_20887,N_18936);
nand UO_1766 (O_1766,N_21354,N_23813);
nand UO_1767 (O_1767,N_22800,N_24351);
nor UO_1768 (O_1768,N_23333,N_24375);
nor UO_1769 (O_1769,N_22921,N_24762);
nor UO_1770 (O_1770,N_21047,N_19863);
and UO_1771 (O_1771,N_19602,N_19745);
nor UO_1772 (O_1772,N_21976,N_19805);
nand UO_1773 (O_1773,N_24600,N_24390);
or UO_1774 (O_1774,N_21948,N_21650);
nand UO_1775 (O_1775,N_24878,N_23450);
xor UO_1776 (O_1776,N_20399,N_22363);
xnor UO_1777 (O_1777,N_21532,N_20178);
or UO_1778 (O_1778,N_22034,N_20980);
nor UO_1779 (O_1779,N_20380,N_22728);
nor UO_1780 (O_1780,N_20581,N_23232);
nor UO_1781 (O_1781,N_24303,N_20065);
xnor UO_1782 (O_1782,N_23888,N_21371);
xor UO_1783 (O_1783,N_19080,N_20941);
nor UO_1784 (O_1784,N_24480,N_22647);
and UO_1785 (O_1785,N_21338,N_21184);
and UO_1786 (O_1786,N_23437,N_19177);
nand UO_1787 (O_1787,N_22009,N_24031);
and UO_1788 (O_1788,N_24754,N_18958);
nor UO_1789 (O_1789,N_20229,N_20533);
or UO_1790 (O_1790,N_20726,N_21638);
nor UO_1791 (O_1791,N_21150,N_21632);
and UO_1792 (O_1792,N_21050,N_21360);
nor UO_1793 (O_1793,N_24451,N_20725);
or UO_1794 (O_1794,N_24381,N_20122);
nor UO_1795 (O_1795,N_21756,N_18894);
or UO_1796 (O_1796,N_19001,N_21016);
nand UO_1797 (O_1797,N_21066,N_24395);
and UO_1798 (O_1798,N_18944,N_22361);
and UO_1799 (O_1799,N_23471,N_24996);
and UO_1800 (O_1800,N_24008,N_21985);
nand UO_1801 (O_1801,N_24978,N_19683);
and UO_1802 (O_1802,N_22841,N_23180);
nor UO_1803 (O_1803,N_19543,N_18781);
nand UO_1804 (O_1804,N_21293,N_20854);
xnor UO_1805 (O_1805,N_21731,N_24045);
nand UO_1806 (O_1806,N_21010,N_24442);
xor UO_1807 (O_1807,N_18977,N_21384);
or UO_1808 (O_1808,N_19303,N_22244);
xor UO_1809 (O_1809,N_21265,N_23720);
and UO_1810 (O_1810,N_21820,N_22170);
or UO_1811 (O_1811,N_23699,N_20745);
or UO_1812 (O_1812,N_22946,N_20792);
xor UO_1813 (O_1813,N_20622,N_22940);
xnor UO_1814 (O_1814,N_23508,N_18798);
and UO_1815 (O_1815,N_20716,N_24087);
xnor UO_1816 (O_1816,N_20615,N_24649);
nor UO_1817 (O_1817,N_24046,N_24853);
nand UO_1818 (O_1818,N_20400,N_21404);
xor UO_1819 (O_1819,N_19319,N_20860);
nor UO_1820 (O_1820,N_24841,N_19087);
xor UO_1821 (O_1821,N_18888,N_23320);
or UO_1822 (O_1822,N_20166,N_20561);
or UO_1823 (O_1823,N_23814,N_20276);
nand UO_1824 (O_1824,N_22353,N_20984);
xnor UO_1825 (O_1825,N_21790,N_24063);
and UO_1826 (O_1826,N_19877,N_23380);
or UO_1827 (O_1827,N_23931,N_23807);
and UO_1828 (O_1828,N_23919,N_22025);
nor UO_1829 (O_1829,N_19882,N_20306);
or UO_1830 (O_1830,N_23235,N_24358);
and UO_1831 (O_1831,N_24397,N_21868);
or UO_1832 (O_1832,N_21758,N_21682);
xor UO_1833 (O_1833,N_22825,N_19262);
nand UO_1834 (O_1834,N_20107,N_22270);
nor UO_1835 (O_1835,N_21920,N_20279);
nand UO_1836 (O_1836,N_23176,N_19974);
xnor UO_1837 (O_1837,N_24680,N_22388);
or UO_1838 (O_1838,N_19575,N_24953);
or UO_1839 (O_1839,N_22334,N_22589);
xnor UO_1840 (O_1840,N_19985,N_24736);
xor UO_1841 (O_1841,N_19166,N_20488);
or UO_1842 (O_1842,N_20996,N_23008);
nor UO_1843 (O_1843,N_23993,N_21271);
nand UO_1844 (O_1844,N_20946,N_20249);
nand UO_1845 (O_1845,N_24588,N_20826);
nand UO_1846 (O_1846,N_22006,N_21407);
and UO_1847 (O_1847,N_20363,N_20977);
nand UO_1848 (O_1848,N_24338,N_22456);
and UO_1849 (O_1849,N_20505,N_22874);
nand UO_1850 (O_1850,N_23837,N_20184);
or UO_1851 (O_1851,N_24140,N_23769);
or UO_1852 (O_1852,N_21837,N_22109);
xor UO_1853 (O_1853,N_18971,N_22906);
nor UO_1854 (O_1854,N_20757,N_19829);
or UO_1855 (O_1855,N_22621,N_21825);
or UO_1856 (O_1856,N_22074,N_23763);
nand UO_1857 (O_1857,N_20557,N_23530);
xor UO_1858 (O_1858,N_20442,N_24003);
or UO_1859 (O_1859,N_19058,N_21152);
nand UO_1860 (O_1860,N_19073,N_23174);
nor UO_1861 (O_1861,N_23059,N_19518);
nand UO_1862 (O_1862,N_23132,N_19992);
or UO_1863 (O_1863,N_19395,N_22048);
nand UO_1864 (O_1864,N_22653,N_22333);
and UO_1865 (O_1865,N_20917,N_21911);
nand UO_1866 (O_1866,N_23088,N_23519);
or UO_1867 (O_1867,N_21749,N_24503);
and UO_1868 (O_1868,N_24646,N_23784);
or UO_1869 (O_1869,N_23415,N_19252);
nor UO_1870 (O_1870,N_24220,N_20624);
nor UO_1871 (O_1871,N_20950,N_22626);
nand UO_1872 (O_1872,N_19389,N_22107);
xnor UO_1873 (O_1873,N_21954,N_20194);
nor UO_1874 (O_1874,N_23882,N_21495);
or UO_1875 (O_1875,N_22506,N_21329);
nand UO_1876 (O_1876,N_24826,N_23044);
or UO_1877 (O_1877,N_23061,N_20696);
nor UO_1878 (O_1878,N_23267,N_22923);
nand UO_1879 (O_1879,N_24673,N_23204);
or UO_1880 (O_1880,N_23246,N_19647);
nor UO_1881 (O_1881,N_21017,N_20459);
nand UO_1882 (O_1882,N_20787,N_20172);
nand UO_1883 (O_1883,N_23362,N_23868);
or UO_1884 (O_1884,N_19871,N_20807);
xor UO_1885 (O_1885,N_24330,N_22397);
xor UO_1886 (O_1886,N_24465,N_20000);
xor UO_1887 (O_1887,N_23656,N_22636);
nor UO_1888 (O_1888,N_24453,N_22459);
nand UO_1889 (O_1889,N_24076,N_22814);
nor UO_1890 (O_1890,N_20406,N_19730);
and UO_1891 (O_1891,N_20905,N_21198);
xnor UO_1892 (O_1892,N_21808,N_21469);
and UO_1893 (O_1893,N_19942,N_20502);
or UO_1894 (O_1894,N_24444,N_23541);
nand UO_1895 (O_1895,N_24921,N_24100);
nor UO_1896 (O_1896,N_22828,N_22915);
or UO_1897 (O_1897,N_19646,N_19247);
xnor UO_1898 (O_1898,N_20566,N_23827);
nand UO_1899 (O_1899,N_22364,N_20695);
nand UO_1900 (O_1900,N_20255,N_23173);
nand UO_1901 (O_1901,N_20500,N_19904);
nor UO_1902 (O_1902,N_18882,N_21131);
and UO_1903 (O_1903,N_24597,N_22335);
or UO_1904 (O_1904,N_20153,N_22344);
and UO_1905 (O_1905,N_23253,N_20944);
xnor UO_1906 (O_1906,N_21054,N_20418);
and UO_1907 (O_1907,N_22819,N_22517);
or UO_1908 (O_1908,N_20732,N_24942);
nand UO_1909 (O_1909,N_23495,N_21585);
or UO_1910 (O_1910,N_20245,N_24219);
or UO_1911 (O_1911,N_21030,N_19130);
nor UO_1912 (O_1912,N_23219,N_19261);
nor UO_1913 (O_1913,N_22713,N_22126);
nor UO_1914 (O_1914,N_20140,N_18905);
nor UO_1915 (O_1915,N_23286,N_24021);
xor UO_1916 (O_1916,N_19208,N_21719);
nand UO_1917 (O_1917,N_22708,N_19081);
nor UO_1918 (O_1918,N_19631,N_24990);
nor UO_1919 (O_1919,N_21823,N_20628);
and UO_1920 (O_1920,N_23175,N_20706);
or UO_1921 (O_1921,N_21944,N_20623);
nand UO_1922 (O_1922,N_24326,N_19008);
and UO_1923 (O_1923,N_22737,N_24900);
nand UO_1924 (O_1924,N_23507,N_20654);
and UO_1925 (O_1925,N_20798,N_20036);
or UO_1926 (O_1926,N_19189,N_22461);
and UO_1927 (O_1927,N_19192,N_18966);
nor UO_1928 (O_1928,N_23427,N_20235);
or UO_1929 (O_1929,N_22743,N_24644);
and UO_1930 (O_1930,N_23733,N_23657);
xor UO_1931 (O_1931,N_23221,N_20938);
xor UO_1932 (O_1932,N_21143,N_20378);
or UO_1933 (O_1933,N_21255,N_21564);
and UO_1934 (O_1934,N_24301,N_20598);
nor UO_1935 (O_1935,N_23288,N_24575);
nand UO_1936 (O_1936,N_22217,N_22391);
or UO_1937 (O_1937,N_21521,N_21243);
nor UO_1938 (O_1938,N_19848,N_19691);
or UO_1939 (O_1939,N_20774,N_20976);
nand UO_1940 (O_1940,N_23083,N_24734);
xnor UO_1941 (O_1941,N_24615,N_24676);
nand UO_1942 (O_1942,N_18771,N_19413);
nand UO_1943 (O_1943,N_22997,N_18867);
and UO_1944 (O_1944,N_19874,N_20337);
nand UO_1945 (O_1945,N_21194,N_24097);
nand UO_1946 (O_1946,N_21950,N_23649);
nor UO_1947 (O_1947,N_23480,N_23210);
xnor UO_1948 (O_1948,N_24721,N_19026);
nand UO_1949 (O_1949,N_20226,N_22615);
nor UO_1950 (O_1950,N_22571,N_18995);
and UO_1951 (O_1951,N_19447,N_22093);
nand UO_1952 (O_1952,N_24216,N_19675);
or UO_1953 (O_1953,N_20859,N_22907);
xnor UO_1954 (O_1954,N_21578,N_24211);
xnor UO_1955 (O_1955,N_20190,N_24059);
and UO_1956 (O_1956,N_19387,N_19272);
and UO_1957 (O_1957,N_21305,N_23717);
nor UO_1958 (O_1958,N_21836,N_19833);
nor UO_1959 (O_1959,N_20102,N_21130);
xor UO_1960 (O_1960,N_21916,N_21197);
and UO_1961 (O_1961,N_18863,N_20461);
and UO_1962 (O_1962,N_23513,N_22283);
and UO_1963 (O_1963,N_23606,N_20935);
nand UO_1964 (O_1964,N_24298,N_21297);
nand UO_1965 (O_1965,N_19284,N_18789);
xor UO_1966 (O_1966,N_19790,N_19024);
nand UO_1967 (O_1967,N_23691,N_20108);
and UO_1968 (O_1968,N_23663,N_19216);
nand UO_1969 (O_1969,N_20665,N_21906);
nand UO_1970 (O_1970,N_22759,N_21398);
nor UO_1971 (O_1971,N_24002,N_23343);
xor UO_1972 (O_1972,N_19094,N_18862);
and UO_1973 (O_1973,N_24367,N_22403);
nand UO_1974 (O_1974,N_19623,N_24374);
nor UO_1975 (O_1975,N_19571,N_24343);
and UO_1976 (O_1976,N_22373,N_20555);
nand UO_1977 (O_1977,N_19853,N_22629);
nor UO_1978 (O_1978,N_20991,N_20838);
and UO_1979 (O_1979,N_19067,N_20176);
and UO_1980 (O_1980,N_23742,N_20803);
and UO_1981 (O_1981,N_22331,N_22133);
and UO_1982 (O_1982,N_21912,N_19939);
xor UO_1983 (O_1983,N_18790,N_23200);
nor UO_1984 (O_1984,N_22502,N_24015);
nor UO_1985 (O_1985,N_19802,N_24618);
or UO_1986 (O_1986,N_22267,N_19242);
or UO_1987 (O_1987,N_19946,N_23159);
or UO_1988 (O_1988,N_18887,N_24251);
nand UO_1989 (O_1989,N_23441,N_24235);
and UO_1990 (O_1990,N_22410,N_24768);
nand UO_1991 (O_1991,N_24873,N_23045);
nor UO_1992 (O_1992,N_21089,N_24541);
or UO_1993 (O_1993,N_18818,N_20884);
nand UO_1994 (O_1994,N_24096,N_21019);
xor UO_1995 (O_1995,N_24926,N_24633);
or UO_1996 (O_1996,N_19593,N_21457);
and UO_1997 (O_1997,N_22304,N_23472);
xnor UO_1998 (O_1998,N_21309,N_24259);
and UO_1999 (O_1999,N_22786,N_23370);
or UO_2000 (O_2000,N_23067,N_24274);
xor UO_2001 (O_2001,N_24034,N_24192);
nor UO_2002 (O_2002,N_23534,N_23990);
nand UO_2003 (O_2003,N_20729,N_18835);
nand UO_2004 (O_2004,N_22998,N_22742);
nor UO_2005 (O_2005,N_24886,N_22688);
and UO_2006 (O_2006,N_19227,N_19332);
or UO_2007 (O_2007,N_21993,N_22158);
and UO_2008 (O_2008,N_20013,N_20721);
or UO_2009 (O_2009,N_21075,N_21125);
nand UO_2010 (O_2010,N_23428,N_18841);
xnor UO_2011 (O_2011,N_20149,N_22349);
or UO_2012 (O_2012,N_19867,N_24707);
xor UO_2013 (O_2013,N_21491,N_19418);
nor UO_2014 (O_2014,N_22618,N_20873);
nor UO_2015 (O_2015,N_24161,N_23635);
xor UO_2016 (O_2016,N_23296,N_20538);
xnor UO_2017 (O_2017,N_20513,N_24879);
nor UO_2018 (O_2018,N_20485,N_19430);
xnor UO_2019 (O_2019,N_22993,N_23634);
and UO_2020 (O_2020,N_20501,N_24858);
nand UO_2021 (O_2021,N_23839,N_24692);
nand UO_2022 (O_2022,N_23374,N_24440);
nor UO_2023 (O_2023,N_21548,N_24337);
nor UO_2024 (O_2024,N_20120,N_22696);
or UO_2025 (O_2025,N_18807,N_23250);
nand UO_2026 (O_2026,N_18949,N_21781);
xor UO_2027 (O_2027,N_20283,N_20170);
nor UO_2028 (O_2028,N_19457,N_23478);
nand UO_2029 (O_2029,N_20570,N_24559);
xnor UO_2030 (O_2030,N_22820,N_22351);
xnor UO_2031 (O_2031,N_24090,N_22398);
nor UO_2032 (O_2032,N_20162,N_19076);
and UO_2033 (O_2033,N_21839,N_19578);
and UO_2034 (O_2034,N_21006,N_23130);
xnor UO_2035 (O_2035,N_18942,N_21899);
and UO_2036 (O_2036,N_24723,N_24625);
nand UO_2037 (O_2037,N_18822,N_21102);
nor UO_2038 (O_2038,N_19821,N_21496);
or UO_2039 (O_2039,N_19486,N_21234);
nor UO_2040 (O_2040,N_24491,N_20712);
xor UO_2041 (O_2041,N_24477,N_23162);
xnor UO_2042 (O_2042,N_20059,N_23610);
and UO_2043 (O_2043,N_19672,N_24706);
nand UO_2044 (O_2044,N_24547,N_21681);
nand UO_2045 (O_2045,N_20866,N_20822);
nand UO_2046 (O_2046,N_21838,N_19542);
nor UO_2047 (O_2047,N_24399,N_19005);
nand UO_2048 (O_2048,N_19043,N_19379);
and UO_2049 (O_2049,N_21511,N_19020);
nor UO_2050 (O_2050,N_22893,N_22822);
xor UO_2051 (O_2051,N_19696,N_18999);
xor UO_2052 (O_2052,N_21427,N_19507);
nand UO_2053 (O_2053,N_24918,N_21785);
and UO_2054 (O_2054,N_23453,N_24407);
and UO_2055 (O_2055,N_22603,N_19964);
xnor UO_2056 (O_2056,N_18777,N_22092);
nor UO_2057 (O_2057,N_22552,N_24596);
nor UO_2058 (O_2058,N_24650,N_19638);
nor UO_2059 (O_2059,N_23791,N_20699);
nand UO_2060 (O_2060,N_23078,N_19136);
and UO_2061 (O_2061,N_20303,N_19107);
nor UO_2062 (O_2062,N_21357,N_22650);
nor UO_2063 (O_2063,N_22151,N_22851);
nand UO_2064 (O_2064,N_20735,N_19209);
nand UO_2065 (O_2065,N_22600,N_22788);
and UO_2066 (O_2066,N_21819,N_21717);
nor UO_2067 (O_2067,N_19512,N_24315);
nor UO_2068 (O_2068,N_22944,N_23317);
or UO_2069 (O_2069,N_23516,N_19154);
and UO_2070 (O_2070,N_21346,N_21103);
nand UO_2071 (O_2071,N_24454,N_21569);
nor UO_2072 (O_2072,N_24049,N_24325);
nor UO_2073 (O_2073,N_24408,N_19140);
nor UO_2074 (O_2074,N_24245,N_22734);
or UO_2075 (O_2075,N_24157,N_19924);
or UO_2076 (O_2076,N_21847,N_20529);
and UO_2077 (O_2077,N_23271,N_24120);
nand UO_2078 (O_2078,N_20493,N_21094);
nand UO_2079 (O_2079,N_23469,N_20544);
or UO_2080 (O_2080,N_24604,N_21390);
or UO_2081 (O_2081,N_21039,N_23252);
and UO_2082 (O_2082,N_20174,N_23835);
xnor UO_2083 (O_2083,N_18832,N_23528);
nor UO_2084 (O_2084,N_20964,N_19004);
or UO_2085 (O_2085,N_22162,N_21266);
and UO_2086 (O_2086,N_22542,N_19198);
xor UO_2087 (O_2087,N_22622,N_19799);
nand UO_2088 (O_2088,N_20263,N_24431);
nor UO_2089 (O_2089,N_21236,N_20447);
nand UO_2090 (O_2090,N_22927,N_21409);
nor UO_2091 (O_2091,N_20937,N_24690);
and UO_2092 (O_2092,N_20297,N_20146);
nor UO_2093 (O_2093,N_19510,N_20011);
nor UO_2094 (O_2094,N_23824,N_22234);
nor UO_2095 (O_2095,N_22325,N_19695);
nand UO_2096 (O_2096,N_24529,N_20747);
xor UO_2097 (O_2097,N_19869,N_24722);
nor UO_2098 (O_2098,N_22886,N_18847);
nand UO_2099 (O_2099,N_23892,N_21493);
and UO_2100 (O_2100,N_22887,N_23988);
or UO_2101 (O_2101,N_19808,N_23680);
nor UO_2102 (O_2102,N_20542,N_22972);
nand UO_2103 (O_2103,N_22434,N_24687);
xnor UO_2104 (O_2104,N_21714,N_24666);
nand UO_2105 (O_2105,N_22844,N_23679);
or UO_2106 (O_2106,N_20135,N_20469);
nor UO_2107 (O_2107,N_18907,N_23780);
xnor UO_2108 (O_2108,N_22698,N_22266);
nor UO_2109 (O_2109,N_20973,N_19481);
or UO_2110 (O_2110,N_21223,N_22231);
and UO_2111 (O_2111,N_20147,N_21109);
and UO_2112 (O_2112,N_24067,N_24471);
and UO_2113 (O_2113,N_20391,N_20559);
nand UO_2114 (O_2114,N_23938,N_22845);
xor UO_2115 (O_2115,N_19079,N_19644);
or UO_2116 (O_2116,N_21898,N_23012);
nand UO_2117 (O_2117,N_21670,N_20568);
and UO_2118 (O_2118,N_23392,N_24466);
nor UO_2119 (O_2119,N_21369,N_23986);
nor UO_2120 (O_2120,N_19308,N_21174);
or UO_2121 (O_2121,N_23512,N_21754);
xor UO_2122 (O_2122,N_24382,N_19868);
nand UO_2123 (O_2123,N_23166,N_22641);
xor UO_2124 (O_2124,N_19627,N_18997);
or UO_2125 (O_2125,N_18979,N_19911);
and UO_2126 (O_2126,N_20663,N_18930);
and UO_2127 (O_2127,N_21386,N_20929);
and UO_2128 (O_2128,N_21154,N_19875);
nor UO_2129 (O_2129,N_22119,N_20546);
or UO_2130 (O_2130,N_20908,N_23302);
xor UO_2131 (O_2131,N_18824,N_23636);
nor UO_2132 (O_2132,N_22630,N_24609);
nor UO_2133 (O_2133,N_19857,N_22644);
nand UO_2134 (O_2134,N_20594,N_19966);
or UO_2135 (O_2135,N_22513,N_19186);
nor UO_2136 (O_2136,N_22910,N_21722);
or UO_2137 (O_2137,N_19266,N_23996);
or UO_2138 (O_2138,N_18880,N_21193);
nor UO_2139 (O_2139,N_24359,N_20360);
xnor UO_2140 (O_2140,N_20110,N_20466);
or UO_2141 (O_2141,N_22914,N_23261);
or UO_2142 (O_2142,N_24500,N_21202);
or UO_2143 (O_2143,N_23605,N_20969);
nand UO_2144 (O_2144,N_19276,N_18801);
nor UO_2145 (O_2145,N_20405,N_19131);
and UO_2146 (O_2146,N_19789,N_22891);
xnor UO_2147 (O_2147,N_19129,N_22392);
nor UO_2148 (O_2148,N_24078,N_23202);
or UO_2149 (O_2149,N_20228,N_19765);
or UO_2150 (O_2150,N_20470,N_21997);
and UO_2151 (O_2151,N_22954,N_22448);
nand UO_2152 (O_2152,N_23336,N_20650);
nor UO_2153 (O_2153,N_20430,N_20697);
nor UO_2154 (O_2154,N_21062,N_24346);
nand UO_2155 (O_2155,N_20455,N_21210);
or UO_2156 (O_2156,N_22973,N_24439);
nor UO_2157 (O_2157,N_24237,N_22569);
nor UO_2158 (O_2158,N_21590,N_21423);
nor UO_2159 (O_2159,N_24880,N_23019);
or UO_2160 (O_2160,N_20620,N_21740);
nand UO_2161 (O_2161,N_22694,N_21388);
nor UO_2162 (O_2162,N_23048,N_24118);
xnor UO_2163 (O_2163,N_24306,N_23979);
nor UO_2164 (O_2164,N_20177,N_23959);
and UO_2165 (O_2165,N_20343,N_21843);
nor UO_2166 (O_2166,N_22656,N_24504);
xnor UO_2167 (O_2167,N_23859,N_23832);
nor UO_2168 (O_2168,N_22445,N_19194);
nor UO_2169 (O_2169,N_23620,N_21932);
or UO_2170 (O_2170,N_22345,N_19018);
or UO_2171 (O_2171,N_22560,N_22302);
nand UO_2172 (O_2172,N_19830,N_20056);
nand UO_2173 (O_2173,N_19640,N_18760);
or UO_2174 (O_2174,N_19390,N_22729);
xnor UO_2175 (O_2175,N_21099,N_23515);
nand UO_2176 (O_2176,N_21933,N_21232);
nor UO_2177 (O_2177,N_23575,N_21958);
or UO_2178 (O_2178,N_24982,N_23364);
nand UO_2179 (O_2179,N_23406,N_20239);
xor UO_2180 (O_2180,N_20727,N_24914);
xor UO_2181 (O_2181,N_22002,N_21826);
nand UO_2182 (O_2182,N_22406,N_18893);
nand UO_2183 (O_2183,N_18935,N_19291);
nor UO_2184 (O_2184,N_24190,N_22606);
nor UO_2185 (O_2185,N_21308,N_21258);
and UO_2186 (O_2186,N_22086,N_21484);
nor UO_2187 (O_2187,N_19232,N_21373);
xor UO_2188 (O_2188,N_19806,N_20894);
xnor UO_2189 (O_2189,N_24371,N_18810);
or UO_2190 (O_2190,N_21529,N_21587);
xor UO_2191 (O_2191,N_23443,N_23522);
nand UO_2192 (O_2192,N_23572,N_18808);
xnor UO_2193 (O_2193,N_23209,N_24735);
nand UO_2194 (O_2194,N_24810,N_20751);
or UO_2195 (O_2195,N_23361,N_23264);
and UO_2196 (O_2196,N_19083,N_18812);
nand UO_2197 (O_2197,N_19915,N_24744);
and UO_2198 (O_2198,N_19187,N_19235);
nand UO_2199 (O_2199,N_22294,N_20789);
nor UO_2200 (O_2200,N_23518,N_18828);
nor UO_2201 (O_2201,N_21165,N_22186);
nand UO_2202 (O_2202,N_24579,N_23042);
xor UO_2203 (O_2203,N_19769,N_22498);
nor UO_2204 (O_2204,N_20413,N_19892);
nand UO_2205 (O_2205,N_21474,N_22473);
nor UO_2206 (O_2206,N_22212,N_20511);
and UO_2207 (O_2207,N_18981,N_22206);
or UO_2208 (O_2208,N_22432,N_24470);
xnor UO_2209 (O_2209,N_22338,N_20207);
xor UO_2210 (O_2210,N_21860,N_24793);
nand UO_2211 (O_2211,N_19558,N_22690);
and UO_2212 (O_2212,N_20272,N_21553);
xnor UO_2213 (O_2213,N_23852,N_24228);
nor UO_2214 (O_2214,N_21359,N_23100);
and UO_2215 (O_2215,N_21975,N_19278);
or UO_2216 (O_2216,N_21372,N_24163);
and UO_2217 (O_2217,N_23687,N_24936);
nand UO_2218 (O_2218,N_23834,N_19010);
or UO_2219 (O_2219,N_22147,N_20683);
or UO_2220 (O_2220,N_19787,N_19599);
or UO_2221 (O_2221,N_23752,N_21631);
xnor UO_2222 (O_2222,N_24686,N_19990);
nand UO_2223 (O_2223,N_20562,N_20629);
and UO_2224 (O_2224,N_20183,N_23875);
nor UO_2225 (O_2225,N_24756,N_21224);
and UO_2226 (O_2226,N_20210,N_20322);
nor UO_2227 (O_2227,N_20670,N_21119);
or UO_2228 (O_2228,N_19742,N_22896);
xor UO_2229 (O_2229,N_20206,N_22394);
or UO_2230 (O_2230,N_22286,N_23570);
nor UO_2231 (O_2231,N_23546,N_21349);
or UO_2232 (O_2232,N_22651,N_21480);
nor UO_2233 (O_2233,N_23995,N_19241);
nor UO_2234 (O_2234,N_24043,N_19244);
and UO_2235 (O_2235,N_18902,N_19619);
xnor UO_2236 (O_2236,N_22802,N_22483);
or UO_2237 (O_2237,N_20388,N_22652);
or UO_2238 (O_2238,N_21960,N_21572);
or UO_2239 (O_2239,N_24798,N_18848);
nand UO_2240 (O_2240,N_20336,N_24162);
and UO_2241 (O_2241,N_20070,N_19914);
or UO_2242 (O_2242,N_23548,N_21465);
nor UO_2243 (O_2243,N_20713,N_24396);
xor UO_2244 (O_2244,N_20440,N_19444);
nor UO_2245 (O_2245,N_21559,N_20788);
or UO_2246 (O_2246,N_24207,N_23218);
and UO_2247 (O_2247,N_19347,N_20291);
nand UO_2248 (O_2248,N_23693,N_24217);
nor UO_2249 (O_2249,N_23191,N_22830);
or UO_2250 (O_2250,N_20640,N_19299);
nand UO_2251 (O_2251,N_23759,N_19273);
xnor UO_2252 (O_2252,N_23983,N_21881);
xnor UO_2253 (O_2253,N_21946,N_20756);
or UO_2254 (O_2254,N_22497,N_21879);
and UO_2255 (O_2255,N_20520,N_21013);
and UO_2256 (O_2256,N_22878,N_24304);
nor UO_2257 (O_2257,N_22811,N_19440);
or UO_2258 (O_2258,N_24032,N_18886);
nand UO_2259 (O_2259,N_23404,N_20637);
or UO_2260 (O_2260,N_22611,N_20523);
nor UO_2261 (O_2261,N_19341,N_18817);
nor UO_2262 (O_2262,N_22050,N_23594);
and UO_2263 (O_2263,N_19572,N_19466);
or UO_2264 (O_2264,N_24066,N_22639);
nor UO_2265 (O_2265,N_19934,N_19788);
and UO_2266 (O_2266,N_21261,N_23499);
nor UO_2267 (O_2267,N_19703,N_22277);
nor UO_2268 (O_2268,N_22499,N_23277);
xor UO_2269 (O_2269,N_21506,N_20913);
nand UO_2270 (O_2270,N_23899,N_24905);
and UO_2271 (O_2271,N_20175,N_19448);
xnor UO_2272 (O_2272,N_22684,N_23358);
and UO_2273 (O_2273,N_21001,N_23484);
and UO_2274 (O_2274,N_22285,N_19750);
xor UO_2275 (O_2275,N_20273,N_19035);
and UO_2276 (O_2276,N_20541,N_21286);
xnor UO_2277 (O_2277,N_20326,N_19012);
nor UO_2278 (O_2278,N_22462,N_23709);
or UO_2279 (O_2279,N_23566,N_23596);
nand UO_2280 (O_2280,N_23324,N_19832);
or UO_2281 (O_2281,N_21475,N_21536);
nand UO_2282 (O_2282,N_23497,N_23027);
nor UO_2283 (O_2283,N_19029,N_22835);
nand UO_2284 (O_2284,N_20015,N_22762);
and UO_2285 (O_2285,N_23479,N_22247);
nand UO_2286 (O_2286,N_20678,N_24013);
or UO_2287 (O_2287,N_20428,N_23369);
nand UO_2288 (O_2288,N_24523,N_23641);
nor UO_2289 (O_2289,N_24392,N_20874);
nand UO_2290 (O_2290,N_24791,N_21925);
nand UO_2291 (O_2291,N_22480,N_22634);
nand UO_2292 (O_2292,N_23239,N_20471);
and UO_2293 (O_2293,N_18878,N_23765);
nor UO_2294 (O_2294,N_24993,N_24787);
nor UO_2295 (O_2295,N_20154,N_19538);
and UO_2296 (O_2296,N_24766,N_24909);
nand UO_2297 (O_2297,N_21080,N_21744);
xnor UO_2298 (O_2298,N_22773,N_20193);
nor UO_2299 (O_2299,N_20655,N_24527);
nor UO_2300 (O_2300,N_22139,N_22779);
and UO_2301 (O_2301,N_22987,N_24804);
xor UO_2302 (O_2302,N_19472,N_19837);
or UO_2303 (O_2303,N_19741,N_18911);
and UO_2304 (O_2304,N_23652,N_23685);
and UO_2305 (O_2305,N_21383,N_20268);
or UO_2306 (O_2306,N_21570,N_19935);
and UO_2307 (O_2307,N_23831,N_24927);
nor UO_2308 (O_2308,N_23135,N_19363);
or UO_2309 (O_2309,N_21771,N_22346);
nor UO_2310 (O_2310,N_21800,N_22342);
nor UO_2311 (O_2311,N_22627,N_20201);
and UO_2312 (O_2312,N_21601,N_24581);
and UO_2313 (O_2313,N_20682,N_22018);
xor UO_2314 (O_2314,N_23609,N_20815);
xor UO_2315 (O_2315,N_23943,N_21418);
nand UO_2316 (O_2316,N_18901,N_23771);
and UO_2317 (O_2317,N_21208,N_19907);
and UO_2318 (O_2318,N_21273,N_24449);
xor UO_2319 (O_2319,N_20956,N_20849);
or UO_2320 (O_2320,N_21750,N_22324);
and UO_2321 (O_2321,N_23503,N_23199);
xor UO_2322 (O_2322,N_23631,N_19488);
nor UO_2323 (O_2323,N_21762,N_19311);
nor UO_2324 (O_2324,N_20744,N_24285);
xnor UO_2325 (O_2325,N_20458,N_22624);
or UO_2326 (O_2326,N_21865,N_23550);
nand UO_2327 (O_2327,N_19429,N_18792);
nor UO_2328 (O_2328,N_24929,N_21659);
xor UO_2329 (O_2329,N_20246,N_22970);
xor UO_2330 (O_2330,N_19548,N_21614);
or UO_2331 (O_2331,N_21627,N_21668);
xnor UO_2332 (O_2332,N_19292,N_23167);
nand UO_2333 (O_2333,N_23966,N_19688);
or UO_2334 (O_2334,N_23133,N_22144);
and UO_2335 (O_2335,N_20331,N_24525);
or UO_2336 (O_2336,N_20926,N_23473);
and UO_2337 (O_2337,N_21649,N_21325);
and UO_2338 (O_2338,N_19905,N_18918);
xnor UO_2339 (O_2339,N_23847,N_22317);
nand UO_2340 (O_2340,N_23896,N_21086);
nor UO_2341 (O_2341,N_20126,N_20928);
xnor UO_2342 (O_2342,N_19203,N_22905);
xor UO_2343 (O_2343,N_20909,N_20754);
nand UO_2344 (O_2344,N_22795,N_24971);
xor UO_2345 (O_2345,N_23070,N_24743);
and UO_2346 (O_2346,N_24156,N_23884);
xor UO_2347 (O_2347,N_23869,N_23113);
or UO_2348 (O_2348,N_21133,N_20053);
or UO_2349 (O_2349,N_23674,N_19415);
nand UO_2350 (O_2350,N_20286,N_20424);
or UO_2351 (O_2351,N_19438,N_24019);
and UO_2352 (O_2352,N_21961,N_24526);
or UO_2353 (O_2353,N_24355,N_22070);
or UO_2354 (O_2354,N_19713,N_19113);
nand UO_2355 (O_2355,N_23786,N_21703);
and UO_2356 (O_2356,N_22460,N_22436);
xor UO_2357 (O_2357,N_20633,N_19552);
nand UO_2358 (O_2358,N_22846,N_20919);
nor UO_2359 (O_2359,N_19775,N_24568);
and UO_2360 (O_2360,N_24083,N_19175);
nor UO_2361 (O_2361,N_21144,N_24695);
nor UO_2362 (O_2362,N_19818,N_23220);
and UO_2363 (O_2363,N_21056,N_21666);
xor UO_2364 (O_2364,N_22557,N_24051);
nand UO_2365 (O_2365,N_21893,N_18904);
nor UO_2366 (O_2366,N_21277,N_24613);
or UO_2367 (O_2367,N_21106,N_23081);
xnor UO_2368 (O_2368,N_21953,N_19038);
xnor UO_2369 (O_2369,N_22883,N_20982);
or UO_2370 (O_2370,N_22948,N_21155);
or UO_2371 (O_2371,N_20608,N_22274);
nor UO_2372 (O_2372,N_24085,N_20278);
xor UO_2373 (O_2373,N_24154,N_21871);
nand UO_2374 (O_2374,N_21615,N_20308);
nand UO_2375 (O_2375,N_24200,N_21272);
and UO_2376 (O_2376,N_20202,N_21237);
xor UO_2377 (O_2377,N_21561,N_18922);
nor UO_2378 (O_2378,N_21979,N_23713);
and UO_2379 (O_2379,N_19340,N_21501);
nor UO_2380 (O_2380,N_21246,N_20855);
nor UO_2381 (O_2381,N_21267,N_18964);
or UO_2382 (O_2382,N_21512,N_20939);
or UO_2383 (O_2383,N_24406,N_20621);
nor UO_2384 (O_2384,N_18898,N_19615);
nor UO_2385 (O_2385,N_18954,N_23205);
nor UO_2386 (O_2386,N_19585,N_21784);
and UO_2387 (O_2387,N_20783,N_24482);
and UO_2388 (O_2388,N_18941,N_24775);
nor UO_2389 (O_2389,N_22481,N_21864);
nand UO_2390 (O_2390,N_23351,N_22981);
nor UO_2391 (O_2391,N_21466,N_24123);
nand UO_2392 (O_2392,N_20219,N_24844);
xor UO_2393 (O_2393,N_19753,N_20671);
or UO_2394 (O_2394,N_20764,N_22337);
nor UO_2395 (O_2395,N_24591,N_21974);
xnor UO_2396 (O_2396,N_22275,N_20853);
and UO_2397 (O_2397,N_19290,N_20274);
nand UO_2398 (O_2398,N_24906,N_22340);
nor UO_2399 (O_2399,N_20090,N_21832);
nor UO_2400 (O_2400,N_22238,N_21538);
and UO_2401 (O_2401,N_24238,N_20089);
nor UO_2402 (O_2402,N_22348,N_20212);
and UO_2403 (O_2403,N_20900,N_24727);
or UO_2404 (O_2404,N_22366,N_21175);
xor UO_2405 (O_2405,N_24617,N_20020);
and UO_2406 (O_2406,N_22756,N_22476);
nand UO_2407 (O_2407,N_20763,N_20463);
nand UO_2408 (O_2408,N_21463,N_21982);
or UO_2409 (O_2409,N_24336,N_22765);
and UO_2410 (O_2410,N_24474,N_24110);
or UO_2411 (O_2411,N_20323,N_23367);
and UO_2412 (O_2412,N_22026,N_23537);
nand UO_2413 (O_2413,N_21987,N_19676);
and UO_2414 (O_2414,N_22089,N_22054);
nand UO_2415 (O_2415,N_21610,N_23316);
xor UO_2416 (O_2416,N_20437,N_22619);
and UO_2417 (O_2417,N_21678,N_19903);
xor UO_2418 (O_2418,N_23583,N_21939);
and UO_2419 (O_2419,N_21636,N_23935);
and UO_2420 (O_2420,N_20812,N_21643);
nand UO_2421 (O_2421,N_20891,N_24177);
and UO_2422 (O_2422,N_24204,N_22722);
and UO_2423 (O_2423,N_22715,N_23514);
or UO_2424 (O_2424,N_24840,N_20173);
or UO_2425 (O_2425,N_21341,N_23984);
nor UO_2426 (O_2426,N_19747,N_18875);
xnor UO_2427 (O_2427,N_21284,N_22996);
nand UO_2428 (O_2428,N_21355,N_24871);
and UO_2429 (O_2429,N_21882,N_19680);
xnor UO_2430 (O_2430,N_20236,N_19781);
or UO_2431 (O_2431,N_21282,N_22296);
or UO_2432 (O_2432,N_24776,N_23385);
or UO_2433 (O_2433,N_22085,N_23104);
xnor UO_2434 (O_2434,N_21031,N_19036);
or UO_2435 (O_2435,N_22055,N_22113);
or UO_2436 (O_2436,N_24759,N_20825);
and UO_2437 (O_2437,N_18968,N_21517);
nand UO_2438 (O_2438,N_22753,N_21658);
nand UO_2439 (O_2439,N_21112,N_20392);
nand UO_2440 (O_2440,N_23857,N_23568);
and UO_2441 (O_2441,N_19357,N_22681);
nand UO_2442 (O_2442,N_23510,N_24954);
or UO_2443 (O_2443,N_18900,N_21909);
and UO_2444 (O_2444,N_22450,N_20758);
or UO_2445 (O_2445,N_24910,N_24384);
and UO_2446 (O_2446,N_24429,N_19582);
xnor UO_2447 (O_2447,N_24970,N_18923);
nor UO_2448 (O_2448,N_24117,N_20536);
xnor UO_2449 (O_2449,N_22027,N_24522);
or UO_2450 (O_2450,N_22935,N_20579);
or UO_2451 (O_2451,N_20451,N_20209);
nor UO_2452 (O_2452,N_19987,N_21381);
or UO_2453 (O_2453,N_24448,N_20898);
and UO_2454 (O_2454,N_19873,N_19513);
nor UO_2455 (O_2455,N_24366,N_20701);
and UO_2456 (O_2456,N_22529,N_21653);
nor UO_2457 (O_2457,N_23388,N_19240);
or UO_2458 (O_2458,N_21831,N_21233);
or UO_2459 (O_2459,N_19397,N_23920);
nor UO_2460 (O_2460,N_23357,N_20752);
nand UO_2461 (O_2461,N_19433,N_19620);
nand UO_2462 (O_2462,N_23143,N_21712);
xor UO_2463 (O_2463,N_22387,N_23937);
nand UO_2464 (O_2464,N_18932,N_18773);
xnor UO_2465 (O_2465,N_22686,N_24554);
xor UO_2466 (O_2466,N_20920,N_22328);
and UO_2467 (O_2467,N_24241,N_18919);
nand UO_2468 (O_2468,N_20948,N_18854);
xor UO_2469 (O_2469,N_24027,N_21228);
nand UO_2470 (O_2470,N_21204,N_19007);
nand UO_2471 (O_2471,N_22386,N_24101);
xnor UO_2472 (O_2472,N_21191,N_22787);
or UO_2473 (O_2473,N_18916,N_22879);
or UO_2474 (O_2474,N_24528,N_24573);
and UO_2475 (O_2475,N_24986,N_23034);
nand UO_2476 (O_2476,N_20446,N_22165);
nor UO_2477 (O_2477,N_23223,N_22305);
nand UO_2478 (O_2478,N_21113,N_23833);
or UO_2479 (O_2479,N_21446,N_19684);
xnor UO_2480 (O_2480,N_20603,N_18786);
nor UO_2481 (O_2481,N_24515,N_24981);
nand UO_2482 (O_2482,N_20930,N_19463);
xnor UO_2483 (O_2483,N_18759,N_23946);
nand UO_2484 (O_2484,N_21751,N_23818);
nand UO_2485 (O_2485,N_22888,N_21892);
nand UO_2486 (O_2486,N_20514,N_23452);
or UO_2487 (O_2487,N_23964,N_20480);
and UO_2488 (O_2488,N_23913,N_19212);
or UO_2489 (O_2489,N_21742,N_24737);
nand UO_2490 (O_2490,N_21444,N_22672);
nor UO_2491 (O_2491,N_22689,N_22763);
and UO_2492 (O_2492,N_19147,N_18890);
nand UO_2493 (O_2493,N_22528,N_22807);
xnor UO_2494 (O_2494,N_22941,N_21101);
or UO_2495 (O_2495,N_19739,N_22776);
and UO_2496 (O_2496,N_20181,N_24892);
or UO_2497 (O_2497,N_21183,N_21240);
or UO_2498 (O_2498,N_19859,N_23748);
and UO_2499 (O_2499,N_24320,N_23401);
and UO_2500 (O_2500,N_24246,N_24030);
nor UO_2501 (O_2501,N_22239,N_18852);
and UO_2502 (O_2502,N_24979,N_19563);
nand UO_2503 (O_2503,N_18912,N_24288);
and UO_2504 (O_2504,N_19673,N_23889);
nand UO_2505 (O_2505,N_20383,N_22059);
nor UO_2506 (O_2506,N_24947,N_23071);
or UO_2507 (O_2507,N_24752,N_23549);
nand UO_2508 (O_2508,N_22492,N_23483);
nand UO_2509 (O_2509,N_19289,N_20673);
and UO_2510 (O_2510,N_21314,N_21775);
or UO_2511 (O_2511,N_22306,N_24040);
and UO_2512 (O_2512,N_20225,N_23886);
xnor UO_2513 (O_2513,N_20032,N_21333);
or UO_2514 (O_2514,N_24558,N_24222);
and UO_2515 (O_2515,N_18998,N_20465);
and UO_2516 (O_2516,N_23608,N_19051);
nor UO_2517 (O_2517,N_23776,N_22850);
nor UO_2518 (O_2518,N_19878,N_22645);
nor UO_2519 (O_2519,N_19327,N_23822);
or UO_2520 (O_2520,N_23247,N_20636);
xnor UO_2521 (O_2521,N_24349,N_21351);
or UO_2522 (O_2522,N_24499,N_24924);
nand UO_2523 (O_2523,N_23730,N_21118);
or UO_2524 (O_2524,N_24488,N_20780);
nor UO_2525 (O_2525,N_21665,N_23272);
xor UO_2526 (O_2526,N_21108,N_20857);
or UO_2527 (O_2527,N_19420,N_23701);
or UO_2528 (O_2528,N_23278,N_21907);
xnor UO_2529 (O_2529,N_19400,N_24231);
nand UO_2530 (O_2530,N_22692,N_22452);
nand UO_2531 (O_2531,N_21088,N_23658);
xnor UO_2532 (O_2532,N_19468,N_21537);
nor UO_2533 (O_2533,N_20646,N_20476);
xnor UO_2534 (O_2534,N_19569,N_23682);
nand UO_2535 (O_2535,N_24149,N_19933);
or UO_2536 (O_2536,N_21379,N_19211);
nand UO_2537 (O_2537,N_18816,N_19556);
xor UO_2538 (O_2538,N_22019,N_20524);
or UO_2539 (O_2539,N_21904,N_24792);
and UO_2540 (O_2540,N_21926,N_22037);
nand UO_2541 (O_2541,N_19978,N_23544);
xnor UO_2542 (O_2542,N_22411,N_22983);
xnor UO_2543 (O_2543,N_18788,N_20427);
xor UO_2544 (O_2544,N_24432,N_21817);
and UO_2545 (O_2545,N_22116,N_19888);
and UO_2546 (O_2546,N_24592,N_20574);
xor UO_2547 (O_2547,N_22193,N_21880);
nand UO_2548 (O_2548,N_21036,N_20161);
xnor UO_2549 (O_2549,N_22789,N_23447);
or UO_2550 (O_2550,N_23224,N_20782);
xnor UO_2551 (O_2551,N_21680,N_19144);
and UO_2552 (O_2552,N_24719,N_22368);
nand UO_2553 (O_2553,N_19373,N_21955);
and UO_2554 (O_2554,N_21391,N_24292);
and UO_2555 (O_2555,N_19917,N_24091);
or UO_2556 (O_2556,N_21092,N_23798);
and UO_2557 (O_2557,N_22360,N_20734);
nand UO_2558 (O_2558,N_24641,N_19260);
xnor UO_2559 (O_2559,N_23655,N_21599);
or UO_2560 (O_2560,N_20305,N_19015);
or UO_2561 (O_2561,N_19975,N_23602);
nand UO_2562 (O_2562,N_19551,N_21486);
nor UO_2563 (O_2563,N_19217,N_19342);
and UO_2564 (O_2564,N_22605,N_21196);
or UO_2565 (O_2565,N_23155,N_24472);
or UO_2566 (O_2566,N_21556,N_22974);
or UO_2567 (O_2567,N_19185,N_19648);
xnor UO_2568 (O_2568,N_20686,N_19075);
and UO_2569 (O_2569,N_22724,N_22771);
and UO_2570 (O_2570,N_21641,N_21802);
nor UO_2571 (O_2571,N_24946,N_22813);
nor UO_2572 (O_2572,N_24757,N_20288);
and UO_2573 (O_2573,N_21310,N_24985);
or UO_2574 (O_2574,N_23873,N_24679);
or UO_2575 (O_2575,N_20367,N_19126);
nand UO_2576 (O_2576,N_23732,N_20556);
or UO_2577 (O_2577,N_24874,N_22873);
or UO_2578 (O_2578,N_22805,N_23517);
nand UO_2579 (O_2579,N_18915,N_20718);
or UO_2580 (O_2580,N_24661,N_24881);
and UO_2581 (O_2581,N_22152,N_22885);
and UO_2582 (O_2582,N_19493,N_22219);
nand UO_2583 (O_2583,N_22838,N_19474);
nand UO_2584 (O_2584,N_23893,N_23003);
xnor UO_2585 (O_2585,N_22197,N_20341);
nand UO_2586 (O_2586,N_19124,N_20460);
nor UO_2587 (O_2587,N_21861,N_21287);
or UO_2588 (O_2588,N_21363,N_22014);
or UO_2589 (O_2589,N_22744,N_20055);
nor UO_2590 (O_2590,N_24988,N_21581);
nand UO_2591 (O_2591,N_22808,N_20610);
xor UO_2592 (O_2592,N_22979,N_23142);
nand UO_2593 (O_2593,N_24175,N_21213);
xor UO_2594 (O_2594,N_20398,N_20653);
and UO_2595 (O_2595,N_24369,N_19386);
or UO_2596 (O_2596,N_22490,N_19774);
and UO_2597 (O_2597,N_20994,N_19590);
nor UO_2598 (O_2598,N_21051,N_22196);
xor UO_2599 (O_2599,N_21365,N_23557);
or UO_2600 (O_2600,N_22327,N_24870);
xnor UO_2601 (O_2601,N_24779,N_19989);
and UO_2602 (O_2602,N_23009,N_18791);
nor UO_2603 (O_2603,N_23710,N_24712);
nand UO_2604 (O_2604,N_23097,N_24598);
xnor UO_2605 (O_2605,N_22665,N_22930);
nor UO_2606 (O_2606,N_24323,N_21726);
xnor UO_2607 (O_2607,N_24014,N_20366);
and UO_2608 (O_2608,N_20252,N_19060);
or UO_2609 (O_2609,N_20076,N_23365);
nor UO_2610 (O_2610,N_21664,N_21035);
nor UO_2611 (O_2611,N_21949,N_22268);
xnor UO_2612 (O_2612,N_24147,N_24555);
nor UO_2613 (O_2613,N_24126,N_24075);
xor UO_2614 (O_2614,N_23961,N_21140);
nand UO_2615 (O_2615,N_20096,N_23683);
or UO_2616 (O_2616,N_19164,N_24356);
and UO_2617 (O_2617,N_20952,N_19589);
or UO_2618 (O_2618,N_22849,N_21226);
nor UO_2619 (O_2619,N_22163,N_19515);
and UO_2620 (O_2620,N_23930,N_19454);
nor UO_2621 (O_2621,N_21727,N_18764);
nor UO_2622 (O_2622,N_20569,N_22124);
and UO_2623 (O_2623,N_23409,N_20237);
nand UO_2624 (O_2624,N_24875,N_22466);
xor UO_2625 (O_2625,N_21336,N_19947);
nand UO_2626 (O_2626,N_22477,N_21604);
nor UO_2627 (O_2627,N_19529,N_24370);
or UO_2628 (O_2628,N_18945,N_20547);
nand UO_2629 (O_2629,N_24387,N_21813);
and UO_2630 (O_2630,N_23681,N_23260);
or UO_2631 (O_2631,N_21217,N_19710);
nand UO_2632 (O_2632,N_21964,N_23339);
nor UO_2633 (O_2633,N_22558,N_21603);
xor UO_2634 (O_2634,N_23144,N_19238);
xor UO_2635 (O_2635,N_18838,N_23440);
and UO_2636 (O_2636,N_20674,N_20897);
or UO_2637 (O_2637,N_20499,N_21146);
and UO_2638 (O_2638,N_19069,N_22137);
xor UO_2639 (O_2639,N_22577,N_19740);
nand UO_2640 (O_2640,N_21311,N_23592);
nor UO_2641 (O_2641,N_19663,N_22892);
nand UO_2642 (O_2642,N_24048,N_24299);
xor UO_2643 (O_2643,N_23474,N_24580);
and UO_2644 (O_2644,N_20809,N_24901);
xor UO_2645 (O_2645,N_23390,N_18967);
nand UO_2646 (O_2646,N_19624,N_24842);
and UO_2647 (O_2647,N_20260,N_22112);
nor UO_2648 (O_2648,N_22062,N_24165);
xor UO_2649 (O_2649,N_19811,N_23772);
nor UO_2650 (O_2650,N_23777,N_18827);
or UO_2651 (O_2651,N_21887,N_23274);
nand UO_2652 (O_2652,N_20914,N_23387);
and UO_2653 (O_2653,N_22102,N_20753);
nor UO_2654 (O_2654,N_21307,N_24688);
xor UO_2655 (O_2655,N_23980,N_22757);
nand UO_2656 (O_2656,N_20988,N_18937);
nand UO_2657 (O_2657,N_22371,N_18858);
nor UO_2658 (O_2658,N_19222,N_18913);
or UO_2659 (O_2659,N_20517,N_22423);
and UO_2660 (O_2660,N_22669,N_22160);
nand UO_2661 (O_2661,N_21812,N_20046);
or UO_2662 (O_2662,N_21841,N_23828);
nand UO_2663 (O_2663,N_24260,N_22136);
or UO_2664 (O_2664,N_24360,N_20099);
xnor UO_2665 (O_2665,N_22988,N_23934);
nor UO_2666 (O_2666,N_21348,N_23127);
xor UO_2667 (O_2667,N_20119,N_22827);
nand UO_2668 (O_2668,N_19584,N_22761);
nand UO_2669 (O_2669,N_24181,N_21977);
nor UO_2670 (O_2670,N_22422,N_21647);
xor UO_2671 (O_2671,N_19751,N_22612);
xor UO_2672 (O_2672,N_19784,N_20896);
or UO_2673 (O_2673,N_19533,N_23050);
xor UO_2674 (O_2674,N_23128,N_20293);
nor UO_2675 (O_2675,N_24372,N_21406);
xor UO_2676 (O_2676,N_22754,N_19801);
nand UO_2677 (O_2677,N_21674,N_22984);
nand UO_2678 (O_2678,N_24567,N_20899);
xor UO_2679 (O_2679,N_24843,N_21402);
xnor UO_2680 (O_2680,N_24028,N_19111);
and UO_2681 (O_2681,N_24201,N_19201);
nand UO_2682 (O_2682,N_23582,N_20079);
nand UO_2683 (O_2683,N_19449,N_21691);
xnor UO_2684 (O_2684,N_23322,N_22823);
xnor UO_2685 (O_2685,N_21321,N_20433);
and UO_2686 (O_2686,N_23240,N_24595);
and UO_2687 (O_2687,N_19625,N_19847);
and UO_2688 (O_2688,N_20933,N_23793);
xor UO_2689 (O_2689,N_21264,N_23487);
nand UO_2690 (O_2690,N_22311,N_18836);
nor UO_2691 (O_2691,N_22659,N_24689);
xor UO_2692 (O_2692,N_22926,N_19458);
xnor UO_2693 (O_2693,N_19645,N_24859);
and UO_2694 (O_2694,N_20163,N_21026);
xnor UO_2695 (O_2695,N_22870,N_24590);
xor UO_2696 (O_2696,N_21606,N_22474);
nor UO_2697 (O_2697,N_19671,N_18872);
nor UO_2698 (O_2698,N_22881,N_20743);
nand UO_2699 (O_2699,N_23865,N_22003);
nor UO_2700 (O_2700,N_20242,N_21171);
or UO_2701 (O_2701,N_19044,N_24601);
or UO_2702 (O_2702,N_23989,N_23057);
nor UO_2703 (O_2703,N_20389,N_22801);
nand UO_2704 (O_2704,N_18842,N_20981);
xnor UO_2705 (O_2705,N_22494,N_23062);
and UO_2706 (O_2706,N_21456,N_24958);
nor UO_2707 (O_2707,N_22675,N_24684);
xor UO_2708 (O_2708,N_19728,N_24945);
nand UO_2709 (O_2709,N_19503,N_20050);
or UO_2710 (O_2710,N_22957,N_23744);
nand UO_2711 (O_2711,N_22257,N_22919);
xnor UO_2712 (O_2712,N_23707,N_20612);
nor UO_2713 (O_2713,N_24760,N_24081);
and UO_2714 (O_2714,N_24254,N_23024);
or UO_2715 (O_2715,N_22794,N_19642);
and UO_2716 (O_2716,N_23958,N_24473);
and UO_2717 (O_2717,N_19702,N_19729);
xnor UO_2718 (O_2718,N_19809,N_24846);
or UO_2719 (O_2719,N_23486,N_21927);
nor UO_2720 (O_2720,N_23160,N_22451);
or UO_2721 (O_2721,N_21943,N_21513);
xor UO_2722 (O_2722,N_20652,N_18761);
or UO_2723 (O_2723,N_19350,N_21071);
or UO_2724 (O_2724,N_21582,N_20599);
nand UO_2725 (O_2725,N_23630,N_19369);
nor UO_2726 (O_2726,N_23046,N_24316);
nand UO_2727 (O_2727,N_21405,N_22586);
xor UO_2728 (O_2728,N_23207,N_24903);
nor UO_2729 (O_2729,N_24612,N_20473);
or UO_2730 (O_2730,N_20959,N_21432);
or UO_2731 (O_2731,N_24037,N_23470);
xor UO_2732 (O_2732,N_22632,N_19944);
xnor UO_2733 (O_2733,N_20796,N_19306);
or UO_2734 (O_2734,N_24557,N_23883);
nand UO_2735 (O_2735,N_24068,N_23464);
nor UO_2736 (O_2736,N_22965,N_21730);
or UO_2737 (O_2737,N_24611,N_20018);
or UO_2738 (O_2738,N_20407,N_19230);
or UO_2739 (O_2739,N_21913,N_24805);
or UO_2740 (O_2740,N_23117,N_23948);
xor UO_2741 (O_2741,N_23489,N_22058);
or UO_2742 (O_2742,N_24822,N_24717);
and UO_2743 (O_2743,N_21042,N_19009);
nor UO_2744 (O_2744,N_22769,N_19495);
nand UO_2745 (O_2745,N_19178,N_21060);
or UO_2746 (O_2746,N_18784,N_23400);
and UO_2747 (O_2747,N_23755,N_20989);
or UO_2748 (O_2748,N_19422,N_19651);
nand UO_2749 (O_2749,N_21857,N_22237);
xor UO_2750 (O_2750,N_21115,N_21535);
or UO_2751 (O_2751,N_20453,N_23987);
nor UO_2752 (O_2752,N_23299,N_22777);
or UO_2753 (O_2753,N_19328,N_20040);
or UO_2754 (O_2754,N_21002,N_24106);
xnor UO_2755 (O_2755,N_23276,N_24809);
nor UO_2756 (O_2756,N_20185,N_23587);
or UO_2757 (O_2757,N_20881,N_20863);
xor UO_2758 (O_2758,N_24077,N_23010);
xor UO_2759 (O_2759,N_19754,N_22443);
xnor UO_2760 (O_2760,N_19943,N_23098);
or UO_2761 (O_2761,N_20257,N_24024);
and UO_2762 (O_2762,N_21138,N_24248);
and UO_2763 (O_2763,N_24479,N_21648);
and UO_2764 (O_2764,N_22216,N_23853);
or UO_2765 (O_2765,N_19957,N_22098);
xor UO_2766 (O_2766,N_20339,N_22227);
or UO_2767 (O_2767,N_19758,N_20017);
xor UO_2768 (O_2768,N_23714,N_22853);
xnor UO_2769 (O_2769,N_20218,N_20452);
or UO_2770 (O_2770,N_19708,N_19399);
nor UO_2771 (O_2771,N_21769,N_20112);
nand UO_2772 (O_2772,N_22176,N_21729);
or UO_2773 (O_2773,N_20422,N_22293);
nor UO_2774 (O_2774,N_22464,N_22772);
or UO_2775 (O_2775,N_18821,N_24824);
and UO_2776 (O_2776,N_21453,N_24244);
xor UO_2777 (O_2777,N_24016,N_22350);
or UO_2778 (O_2778,N_23158,N_19127);
xor UO_2779 (O_2779,N_21846,N_22531);
nor UO_2780 (O_2780,N_22322,N_20142);
and UO_2781 (O_2781,N_23672,N_21093);
and UO_2782 (O_2782,N_20890,N_19382);
nand UO_2783 (O_2783,N_18896,N_18975);
xor UO_2784 (O_2784,N_18767,N_21127);
xnor UO_2785 (O_2785,N_19550,N_22566);
nand UO_2786 (O_2786,N_24984,N_21340);
xnor UO_2787 (O_2787,N_18957,N_24398);
xnor UO_2788 (O_2788,N_21624,N_24155);
xor UO_2789 (O_2789,N_19091,N_22646);
and UO_2790 (O_2790,N_24056,N_20720);
xor UO_2791 (O_2791,N_21479,N_19557);
or UO_2792 (O_2792,N_24215,N_19121);
or UO_2793 (O_2793,N_22561,N_23023);
nand UO_2794 (O_2794,N_20728,N_24849);
and UO_2795 (O_2795,N_20572,N_21938);
nor UO_2796 (O_2796,N_22449,N_23524);
xnor UO_2797 (O_2797,N_24902,N_20576);
xnor UO_2798 (O_2798,N_19407,N_21685);
nand UO_2799 (O_2799,N_19635,N_23864);
nor UO_2800 (O_2800,N_19473,N_23505);
nor UO_2801 (O_2801,N_21167,N_21507);
nor UO_2802 (O_2802,N_21312,N_24800);
xor UO_2803 (O_2803,N_21343,N_23360);
nand UO_2804 (O_2804,N_21724,N_24697);
or UO_2805 (O_2805,N_19970,N_22377);
nand UO_2806 (O_2806,N_19756,N_21014);
and UO_2807 (O_2807,N_19352,N_22181);
or UO_2808 (O_2808,N_23424,N_19559);
xor UO_2809 (O_2809,N_19068,N_20797);
nand UO_2810 (O_2810,N_18928,N_24531);
and UO_2811 (O_2811,N_20259,N_21889);
nor UO_2812 (O_2812,N_19843,N_19723);
and UO_2813 (O_2813,N_23107,N_22073);
xnor UO_2814 (O_2814,N_19879,N_23573);
or UO_2815 (O_2815,N_21482,N_19716);
and UO_2816 (O_2816,N_21429,N_20921);
and UO_2817 (O_2817,N_21023,N_21833);
xor UO_2818 (O_2818,N_19469,N_22858);
xnor UO_2819 (O_2819,N_21049,N_23738);
xnor UO_2820 (O_2820,N_19973,N_23354);
nor UO_2821 (O_2821,N_21617,N_19176);
nor UO_2822 (O_2822,N_24884,N_19870);
nand UO_2823 (O_2823,N_21249,N_21076);
nand UO_2824 (O_2824,N_23998,N_20106);
xnor UO_2825 (O_2825,N_21438,N_19321);
xnor UO_2826 (O_2826,N_20001,N_20634);
xnor UO_2827 (O_2827,N_24920,N_23492);
or UO_2828 (O_2828,N_23041,N_18843);
nor UO_2829 (O_2829,N_21380,N_21984);
nand UO_2830 (O_2830,N_19214,N_19920);
xnor UO_2831 (O_2831,N_23754,N_21551);
and UO_2832 (O_2832,N_21669,N_24731);
or UO_2833 (O_2833,N_19666,N_19749);
xnor UO_2834 (O_2834,N_19353,N_19891);
nor UO_2835 (O_2835,N_18885,N_24519);
xnor UO_2836 (O_2836,N_21368,N_22609);
nor UO_2837 (O_2837,N_19053,N_24476);
and UO_2838 (O_2838,N_24761,N_20482);
and UO_2839 (O_2839,N_19275,N_24441);
xor UO_2840 (O_2840,N_22066,N_21289);
or UO_2841 (O_2841,N_22140,N_22784);
xor UO_2842 (O_2842,N_21394,N_24544);
and UO_2843 (O_2843,N_24354,N_20847);
or UO_2844 (O_2844,N_19953,N_23916);
nand UO_2845 (O_2845,N_19577,N_19370);
nor UO_2846 (O_2846,N_22154,N_18978);
xor UO_2847 (O_2847,N_21375,N_20749);
nand UO_2848 (O_2848,N_19000,N_24997);
nor UO_2849 (O_2849,N_23349,N_21508);
xnor UO_2850 (O_2850,N_22535,N_19323);
and UO_2851 (O_2851,N_22658,N_19461);
or UO_2852 (O_2852,N_19199,N_19931);
xnor UO_2853 (O_2853,N_19770,N_18993);
or UO_2854 (O_2854,N_22489,N_19555);
and UO_2855 (O_2855,N_21207,N_20902);
nor UO_2856 (O_2856,N_19643,N_22859);
nor UO_2857 (O_2857,N_22714,N_20519);
or UO_2858 (O_2858,N_19183,N_22076);
nor UO_2859 (O_2859,N_23049,N_23399);
and UO_2860 (O_2860,N_24934,N_24608);
xor UO_2861 (O_2861,N_22141,N_23190);
nand UO_2862 (O_2862,N_22770,N_23021);
and UO_2863 (O_2863,N_23251,N_21322);
and UO_2864 (O_2864,N_21924,N_21673);
nor UO_2865 (O_2865,N_24582,N_24662);
nor UO_2866 (O_2866,N_24659,N_21736);
or UO_2867 (O_2867,N_20883,N_24496);
xor UO_2868 (O_2868,N_21374,N_20497);
nand UO_2869 (O_2869,N_24258,N_21520);
nand UO_2870 (O_2870,N_20262,N_18826);
nor UO_2871 (O_2871,N_19849,N_20248);
nand UO_2872 (O_2872,N_23588,N_21505);
xor UO_2873 (O_2873,N_22614,N_23007);
xor UO_2874 (O_2874,N_19459,N_20316);
xnor UO_2875 (O_2875,N_21642,N_18825);
xor UO_2876 (O_2876,N_23403,N_18970);
xnor UO_2877 (O_2877,N_20965,N_20993);
nand UO_2878 (O_2878,N_20347,N_23014);
and UO_2879 (O_2879,N_23371,N_19348);
or UO_2880 (O_2880,N_21411,N_22911);
xor UO_2881 (O_2881,N_20588,N_20419);
nand UO_2882 (O_2882,N_21408,N_23877);
nor UO_2883 (O_2883,N_20687,N_21220);
xnor UO_2884 (O_2884,N_19120,N_20940);
nand UO_2885 (O_2885,N_21875,N_19862);
nand UO_2886 (O_2886,N_21005,N_22895);
nand UO_2887 (O_2887,N_21593,N_22625);
nor UO_2888 (O_2888,N_24060,N_22172);
nand UO_2889 (O_2889,N_24125,N_20289);
nand UO_2890 (O_2890,N_21672,N_22030);
and UO_2891 (O_2891,N_22655,N_24134);
nor UO_2892 (O_2892,N_23417,N_22598);
and UO_2893 (O_2893,N_21856,N_23908);
nor UO_2894 (O_2894,N_21854,N_22420);
xor UO_2895 (O_2895,N_23327,N_20123);
nor UO_2896 (O_2896,N_24733,N_21908);
or UO_2897 (O_2897,N_22064,N_19906);
and UO_2898 (O_2898,N_21793,N_23244);
or UO_2899 (O_2899,N_22249,N_22208);
nor UO_2900 (O_2900,N_21571,N_23782);
and UO_2901 (O_2901,N_21764,N_22284);
xnor UO_2902 (O_2902,N_20384,N_22755);
nand UO_2903 (O_2903,N_22758,N_19738);
nor UO_2904 (O_2904,N_20478,N_21472);
nand UO_2905 (O_2905,N_23904,N_19852);
and UO_2906 (O_2906,N_24044,N_24445);
nand UO_2907 (O_2907,N_21447,N_24882);
xor UO_2908 (O_2908,N_19603,N_22872);
xor UO_2909 (O_2909,N_19995,N_22967);
and UO_2910 (O_2910,N_21998,N_21935);
nor UO_2911 (O_2911,N_18853,N_24188);
nand UO_2912 (O_2912,N_20155,N_21149);
nand UO_2913 (O_2913,N_24614,N_24694);
nand UO_2914 (O_2914,N_24868,N_19714);
and UO_2915 (O_2915,N_22289,N_23090);
and UO_2916 (O_2916,N_23722,N_21247);
xor UO_2917 (O_2917,N_24998,N_18796);
xor UO_2918 (O_2918,N_21279,N_20402);
nand UO_2919 (O_2919,N_19506,N_24535);
nor UO_2920 (O_2920,N_21829,N_22220);
nand UO_2921 (O_2921,N_19746,N_23285);
or UO_2922 (O_2922,N_20342,N_20690);
or UO_2923 (O_2923,N_20310,N_23248);
nor UO_2924 (O_2924,N_23257,N_23140);
nor UO_2925 (O_2925,N_22792,N_22602);
nor UO_2926 (O_2926,N_24400,N_21816);
nand UO_2927 (O_2927,N_23254,N_19544);
or UO_2928 (O_2928,N_20614,N_22683);
or UO_2929 (O_2929,N_24631,N_21124);
xor UO_2930 (O_2930,N_18969,N_23001);
xnor UO_2931 (O_2931,N_21502,N_22810);
or UO_2932 (O_2932,N_19172,N_21966);
xor UO_2933 (O_2933,N_19658,N_18951);
and UO_2934 (O_2934,N_19324,N_22545);
xnor UO_2935 (O_2935,N_23498,N_20224);
or UO_2936 (O_2936,N_23172,N_21069);
nand UO_2937 (O_2937,N_20710,N_19711);
and UO_2938 (O_2938,N_22413,N_22115);
xor UO_2939 (O_2939,N_19661,N_23848);
or UO_2940 (O_2940,N_21592,N_21283);
xor UO_2941 (O_2941,N_22182,N_20325);
xnor UO_2942 (O_2942,N_24256,N_22150);
nor UO_2943 (O_2943,N_23747,N_19455);
or UO_2944 (O_2944,N_23727,N_20332);
or UO_2945 (O_2945,N_21008,N_20111);
or UO_2946 (O_2946,N_21748,N_21192);
nand UO_2947 (O_2947,N_20794,N_20167);
nor UO_2948 (O_2948,N_24817,N_23795);
xnor UO_2949 (O_2949,N_21123,N_21095);
and UO_2950 (O_2950,N_18860,N_23397);
nand UO_2951 (O_2951,N_23463,N_22563);
nand UO_2952 (O_2952,N_24108,N_21708);
nand UO_2953 (O_2953,N_24510,N_23836);
xor UO_2954 (O_2954,N_20772,N_22405);
xnor UO_2955 (O_2955,N_21473,N_24950);
or UO_2956 (O_2956,N_22409,N_20831);
or UO_2957 (O_2957,N_23446,N_20868);
xnor UO_2958 (O_2958,N_19002,N_21872);
nor UO_2959 (O_2959,N_22385,N_19686);
xor UO_2960 (O_2960,N_23626,N_23300);
xnor UO_2961 (O_2961,N_24883,N_24361);
or UO_2962 (O_2962,N_23491,N_23817);
and UO_2963 (O_2963,N_21034,N_24347);
nor UO_2964 (O_2964,N_20269,N_23923);
nand UO_2965 (O_2965,N_21562,N_24546);
xnor UO_2966 (O_2966,N_23563,N_23756);
nand UO_2967 (O_2967,N_23060,N_19100);
or UO_2968 (O_2968,N_22963,N_18980);
or UO_2969 (O_2969,N_22485,N_23262);
xor UO_2970 (O_2970,N_20575,N_20597);
and UO_2971 (O_2971,N_24127,N_20061);
xor UO_2972 (O_2972,N_20724,N_20680);
or UO_2973 (O_2973,N_23419,N_21362);
xnor UO_2974 (O_2974,N_23197,N_22007);
or UO_2975 (O_2975,N_22514,N_21723);
and UO_2976 (O_2976,N_20672,N_20057);
or UO_2977 (O_2977,N_20875,N_23467);
nand UO_2978 (O_2978,N_24001,N_18780);
nand UO_2979 (O_2979,N_22706,N_23559);
nand UO_2980 (O_2980,N_19378,N_24224);
and UO_2981 (O_2981,N_19061,N_19165);
nor UO_2982 (O_2982,N_22525,N_22592);
and UO_2983 (O_2983,N_21117,N_18804);
nor UO_2984 (O_2984,N_20230,N_20516);
and UO_2985 (O_2985,N_23909,N_21534);
nand UO_2986 (O_2986,N_21972,N_24339);
xnor UO_2987 (O_2987,N_21385,N_22596);
and UO_2988 (O_2988,N_23778,N_23171);
nor UO_2989 (O_2989,N_24632,N_19269);
nand UO_2990 (O_2990,N_24730,N_24205);
nor UO_2991 (O_2991,N_23161,N_23303);
xor UO_2992 (O_2992,N_19737,N_23785);
or UO_2993 (O_2993,N_23731,N_22581);
nand UO_2994 (O_2994,N_22719,N_19138);
nand UO_2995 (O_2995,N_23092,N_21451);
and UO_2996 (O_2996,N_24456,N_19860);
nand UO_2997 (O_2997,N_22177,N_19090);
nor UO_2998 (O_2998,N_18895,N_19733);
or UO_2999 (O_2999,N_19826,N_18782);
endmodule