module basic_500_3000_500_3_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_230,In_448);
nor U1 (N_1,In_342,In_189);
nor U2 (N_2,In_216,In_449);
and U3 (N_3,In_178,In_274);
nand U4 (N_4,In_144,In_392);
nand U5 (N_5,In_226,In_368);
and U6 (N_6,In_222,In_255);
nor U7 (N_7,In_286,In_263);
or U8 (N_8,In_159,In_271);
and U9 (N_9,In_420,In_139);
nor U10 (N_10,In_456,In_79);
or U11 (N_11,In_333,In_127);
or U12 (N_12,In_113,In_181);
nor U13 (N_13,In_206,In_151);
nand U14 (N_14,In_135,In_57);
nor U15 (N_15,In_229,In_409);
nand U16 (N_16,In_472,In_1);
nor U17 (N_17,In_356,In_129);
xnor U18 (N_18,In_395,In_498);
nor U19 (N_19,In_171,In_126);
nor U20 (N_20,In_68,In_265);
nand U21 (N_21,In_100,In_132);
or U22 (N_22,In_259,In_154);
nand U23 (N_23,In_417,In_370);
nor U24 (N_24,In_367,In_310);
or U25 (N_25,In_204,In_58);
and U26 (N_26,In_147,In_175);
nor U27 (N_27,In_190,In_492);
nand U28 (N_28,In_210,In_77);
or U29 (N_29,In_351,In_65);
or U30 (N_30,In_237,In_13);
or U31 (N_31,In_321,In_287);
and U32 (N_32,In_142,In_212);
nand U33 (N_33,In_258,In_386);
or U34 (N_34,In_439,In_359);
nand U35 (N_35,In_340,In_404);
and U36 (N_36,In_385,In_400);
nand U37 (N_37,In_88,In_481);
and U38 (N_38,In_408,In_249);
nand U39 (N_39,In_174,In_415);
and U40 (N_40,In_338,In_288);
or U41 (N_41,In_84,In_413);
or U42 (N_42,In_443,In_354);
nor U43 (N_43,In_8,In_183);
and U44 (N_44,In_170,In_350);
nand U45 (N_45,In_164,In_453);
nand U46 (N_46,In_149,In_12);
and U47 (N_47,In_3,In_124);
or U48 (N_48,In_290,In_32);
or U49 (N_49,In_223,In_327);
and U50 (N_50,In_238,In_125);
or U51 (N_51,In_433,In_285);
and U52 (N_52,In_99,In_411);
and U53 (N_53,In_316,In_198);
and U54 (N_54,In_442,In_387);
nand U55 (N_55,In_60,In_199);
or U56 (N_56,In_202,In_36);
or U57 (N_57,In_114,In_377);
nor U58 (N_58,In_203,In_362);
nor U59 (N_59,In_233,In_355);
or U60 (N_60,In_197,In_182);
nand U61 (N_61,In_388,In_282);
or U62 (N_62,In_251,In_179);
and U63 (N_63,In_87,In_85);
and U64 (N_64,In_266,In_252);
or U65 (N_65,In_76,In_301);
nor U66 (N_66,In_475,In_29);
and U67 (N_67,In_109,In_107);
nand U68 (N_68,In_261,In_314);
nor U69 (N_69,In_80,In_412);
nor U70 (N_70,In_457,In_378);
or U71 (N_71,In_236,In_103);
or U72 (N_72,In_372,In_161);
nor U73 (N_73,In_346,In_294);
nor U74 (N_74,In_19,In_48);
or U75 (N_75,In_451,In_247);
nor U76 (N_76,In_146,In_353);
and U77 (N_77,In_92,In_307);
or U78 (N_78,In_279,In_38);
and U79 (N_79,In_192,In_334);
or U80 (N_80,In_315,In_53);
nor U81 (N_81,In_27,In_205);
nor U82 (N_82,In_318,In_496);
or U83 (N_83,In_72,In_134);
nand U84 (N_84,In_471,In_269);
or U85 (N_85,In_138,In_276);
nor U86 (N_86,In_193,In_476);
or U87 (N_87,In_89,In_396);
and U88 (N_88,In_384,In_16);
nand U89 (N_89,In_158,In_165);
and U90 (N_90,In_101,In_156);
xnor U91 (N_91,In_153,In_130);
and U92 (N_92,In_264,In_423);
or U93 (N_93,In_106,In_26);
xnor U94 (N_94,In_41,In_234);
nand U95 (N_95,In_64,In_437);
and U96 (N_96,In_464,In_73);
or U97 (N_97,In_267,In_460);
nor U98 (N_98,In_455,In_257);
and U99 (N_99,In_21,In_260);
nand U100 (N_100,In_54,In_10);
or U101 (N_101,In_432,In_141);
nor U102 (N_102,In_108,In_360);
or U103 (N_103,In_292,In_487);
or U104 (N_104,In_461,In_50);
nor U105 (N_105,In_270,In_467);
or U106 (N_106,In_499,In_78);
and U107 (N_107,In_365,In_444);
or U108 (N_108,In_284,In_302);
or U109 (N_109,In_322,In_70);
nand U110 (N_110,In_379,In_200);
and U111 (N_111,In_136,In_300);
nor U112 (N_112,In_97,In_324);
and U113 (N_113,In_470,In_225);
or U114 (N_114,In_42,In_0);
and U115 (N_115,In_427,In_30);
and U116 (N_116,In_228,In_157);
and U117 (N_117,In_66,In_424);
or U118 (N_118,In_37,In_128);
nand U119 (N_119,In_440,In_383);
and U120 (N_120,In_401,In_195);
nand U121 (N_121,In_74,In_480);
or U122 (N_122,In_341,In_435);
and U123 (N_123,In_18,In_332);
or U124 (N_124,In_463,In_393);
nand U125 (N_125,In_361,In_120);
nor U126 (N_126,In_94,In_441);
or U127 (N_127,In_148,In_6);
nor U128 (N_128,In_357,In_336);
nor U129 (N_129,In_343,In_407);
or U130 (N_130,In_352,In_465);
nor U131 (N_131,In_140,In_214);
or U132 (N_132,In_173,In_311);
and U133 (N_133,In_201,In_207);
nor U134 (N_134,In_335,In_227);
nand U135 (N_135,In_312,In_116);
or U136 (N_136,In_122,In_44);
nand U137 (N_137,In_339,In_331);
or U138 (N_138,In_250,In_187);
nor U139 (N_139,In_105,In_391);
or U140 (N_140,In_25,In_218);
nor U141 (N_141,In_4,In_172);
or U142 (N_142,In_102,In_244);
and U143 (N_143,In_418,In_278);
nand U144 (N_144,In_414,In_93);
nor U145 (N_145,In_347,In_83);
nor U146 (N_146,In_320,In_313);
nand U147 (N_147,In_363,In_397);
nor U148 (N_148,In_430,In_348);
nand U149 (N_149,In_188,In_262);
and U150 (N_150,In_23,In_243);
nor U151 (N_151,In_382,In_434);
nor U152 (N_152,In_61,In_458);
nor U153 (N_153,In_35,In_31);
and U154 (N_154,In_117,In_308);
and U155 (N_155,In_45,In_220);
and U156 (N_156,In_82,In_494);
and U157 (N_157,In_69,In_268);
nand U158 (N_158,In_169,In_277);
or U159 (N_159,In_390,In_364);
or U160 (N_160,In_254,In_275);
nor U161 (N_161,In_303,In_474);
xnor U162 (N_162,In_438,In_358);
or U163 (N_163,In_296,In_241);
nor U164 (N_164,In_34,In_52);
and U165 (N_165,In_162,In_495);
or U166 (N_166,In_429,In_297);
xnor U167 (N_167,In_110,In_422);
and U168 (N_168,In_111,In_221);
or U169 (N_169,In_399,In_131);
nor U170 (N_170,In_329,In_493);
and U171 (N_171,In_224,In_49);
nor U172 (N_172,In_155,In_98);
nor U173 (N_173,In_91,In_215);
xor U174 (N_174,In_323,In_22);
nand U175 (N_175,In_375,In_373);
nand U176 (N_176,In_213,In_96);
or U177 (N_177,In_497,In_402);
or U178 (N_178,In_484,In_46);
nand U179 (N_179,In_403,In_39);
nor U180 (N_180,In_328,In_466);
nor U181 (N_181,In_217,In_369);
and U182 (N_182,In_15,In_298);
nor U183 (N_183,In_33,In_143);
nand U184 (N_184,In_299,In_47);
or U185 (N_185,In_479,In_191);
or U186 (N_186,In_425,In_235);
xnor U187 (N_187,In_75,In_289);
nand U188 (N_188,In_330,In_426);
and U189 (N_189,In_194,In_394);
or U190 (N_190,In_389,In_245);
nand U191 (N_191,In_371,In_152);
or U192 (N_192,In_63,In_410);
or U193 (N_193,In_483,In_337);
nor U194 (N_194,In_304,In_431);
nor U195 (N_195,In_118,In_185);
or U196 (N_196,In_24,In_305);
or U197 (N_197,In_231,In_344);
and U198 (N_198,In_436,In_283);
and U199 (N_199,In_326,In_115);
nor U200 (N_200,In_454,In_376);
nand U201 (N_201,In_291,In_280);
and U202 (N_202,In_56,In_349);
nor U203 (N_203,In_133,In_67);
or U204 (N_204,In_309,In_180);
or U205 (N_205,In_112,In_186);
or U206 (N_206,In_273,In_490);
and U207 (N_207,In_81,In_184);
nand U208 (N_208,In_428,In_240);
and U209 (N_209,In_406,In_398);
nand U210 (N_210,In_405,In_28);
and U211 (N_211,In_445,In_137);
or U212 (N_212,In_421,In_2);
nor U213 (N_213,In_374,In_485);
or U214 (N_214,In_121,In_459);
nand U215 (N_215,In_208,In_447);
and U216 (N_216,In_71,In_366);
and U217 (N_217,In_17,In_256);
and U218 (N_218,In_468,In_123);
or U219 (N_219,In_55,In_176);
or U220 (N_220,In_248,In_160);
nor U221 (N_221,In_486,In_95);
or U222 (N_222,In_5,In_163);
nor U223 (N_223,In_167,In_242);
nor U224 (N_224,In_209,In_86);
or U225 (N_225,In_325,In_491);
nand U226 (N_226,In_469,In_295);
xnor U227 (N_227,In_319,In_104);
or U228 (N_228,In_477,In_446);
nor U229 (N_229,In_253,In_317);
nor U230 (N_230,In_272,In_20);
and U231 (N_231,In_478,In_7);
and U232 (N_232,In_43,In_246);
and U233 (N_233,In_40,In_381);
nand U234 (N_234,In_473,In_419);
or U235 (N_235,In_416,In_119);
xor U236 (N_236,In_11,In_62);
nand U237 (N_237,In_14,In_168);
nor U238 (N_238,In_452,In_211);
and U239 (N_239,In_281,In_219);
or U240 (N_240,In_196,In_306);
nand U241 (N_241,In_51,In_232);
or U242 (N_242,In_145,In_293);
nor U243 (N_243,In_345,In_9);
nand U244 (N_244,In_488,In_59);
or U245 (N_245,In_380,In_177);
nand U246 (N_246,In_150,In_450);
or U247 (N_247,In_90,In_166);
and U248 (N_248,In_462,In_489);
nor U249 (N_249,In_239,In_482);
and U250 (N_250,In_61,In_225);
or U251 (N_251,In_297,In_193);
nor U252 (N_252,In_178,In_83);
and U253 (N_253,In_209,In_494);
nor U254 (N_254,In_136,In_31);
and U255 (N_255,In_477,In_49);
nand U256 (N_256,In_279,In_169);
xnor U257 (N_257,In_39,In_37);
xnor U258 (N_258,In_118,In_253);
and U259 (N_259,In_415,In_469);
nor U260 (N_260,In_364,In_418);
nor U261 (N_261,In_344,In_208);
xor U262 (N_262,In_494,In_248);
and U263 (N_263,In_100,In_330);
nand U264 (N_264,In_248,In_203);
nor U265 (N_265,In_205,In_389);
or U266 (N_266,In_224,In_174);
and U267 (N_267,In_218,In_394);
and U268 (N_268,In_17,In_444);
xnor U269 (N_269,In_416,In_166);
nand U270 (N_270,In_167,In_106);
and U271 (N_271,In_365,In_109);
nand U272 (N_272,In_342,In_0);
xnor U273 (N_273,In_434,In_21);
nor U274 (N_274,In_416,In_436);
nor U275 (N_275,In_146,In_174);
and U276 (N_276,In_154,In_231);
nand U277 (N_277,In_418,In_227);
nand U278 (N_278,In_87,In_382);
nor U279 (N_279,In_165,In_382);
nor U280 (N_280,In_474,In_136);
and U281 (N_281,In_50,In_69);
nor U282 (N_282,In_285,In_203);
or U283 (N_283,In_377,In_345);
nand U284 (N_284,In_312,In_45);
nand U285 (N_285,In_142,In_108);
nor U286 (N_286,In_256,In_268);
or U287 (N_287,In_372,In_38);
nor U288 (N_288,In_199,In_229);
or U289 (N_289,In_90,In_148);
nand U290 (N_290,In_98,In_472);
or U291 (N_291,In_174,In_408);
or U292 (N_292,In_82,In_171);
nor U293 (N_293,In_9,In_84);
nand U294 (N_294,In_268,In_94);
or U295 (N_295,In_338,In_141);
nor U296 (N_296,In_336,In_349);
and U297 (N_297,In_79,In_385);
and U298 (N_298,In_463,In_406);
nand U299 (N_299,In_204,In_76);
or U300 (N_300,In_225,In_10);
and U301 (N_301,In_33,In_122);
nor U302 (N_302,In_324,In_479);
nor U303 (N_303,In_86,In_236);
and U304 (N_304,In_15,In_237);
and U305 (N_305,In_365,In_231);
or U306 (N_306,In_494,In_238);
or U307 (N_307,In_144,In_457);
nor U308 (N_308,In_374,In_474);
nor U309 (N_309,In_256,In_459);
or U310 (N_310,In_282,In_232);
nand U311 (N_311,In_63,In_145);
and U312 (N_312,In_111,In_186);
and U313 (N_313,In_407,In_261);
or U314 (N_314,In_227,In_442);
and U315 (N_315,In_412,In_99);
or U316 (N_316,In_73,In_465);
and U317 (N_317,In_279,In_358);
nand U318 (N_318,In_379,In_98);
or U319 (N_319,In_192,In_78);
nor U320 (N_320,In_470,In_173);
and U321 (N_321,In_196,In_135);
or U322 (N_322,In_10,In_491);
nor U323 (N_323,In_88,In_184);
nor U324 (N_324,In_141,In_372);
and U325 (N_325,In_385,In_430);
nand U326 (N_326,In_195,In_49);
or U327 (N_327,In_5,In_460);
and U328 (N_328,In_406,In_286);
nand U329 (N_329,In_255,In_75);
nor U330 (N_330,In_180,In_429);
and U331 (N_331,In_335,In_189);
nand U332 (N_332,In_226,In_144);
nand U333 (N_333,In_31,In_250);
nor U334 (N_334,In_270,In_305);
or U335 (N_335,In_81,In_121);
or U336 (N_336,In_132,In_43);
and U337 (N_337,In_432,In_215);
nor U338 (N_338,In_373,In_129);
and U339 (N_339,In_390,In_429);
or U340 (N_340,In_184,In_272);
or U341 (N_341,In_19,In_474);
or U342 (N_342,In_198,In_209);
nor U343 (N_343,In_181,In_115);
or U344 (N_344,In_281,In_438);
nor U345 (N_345,In_215,In_97);
nand U346 (N_346,In_251,In_5);
or U347 (N_347,In_120,In_261);
nor U348 (N_348,In_153,In_226);
nand U349 (N_349,In_360,In_261);
nor U350 (N_350,In_81,In_77);
nand U351 (N_351,In_404,In_219);
nor U352 (N_352,In_321,In_408);
and U353 (N_353,In_317,In_301);
nand U354 (N_354,In_272,In_89);
nand U355 (N_355,In_309,In_99);
nor U356 (N_356,In_108,In_279);
or U357 (N_357,In_235,In_302);
nor U358 (N_358,In_275,In_244);
and U359 (N_359,In_300,In_465);
nor U360 (N_360,In_244,In_160);
or U361 (N_361,In_326,In_318);
and U362 (N_362,In_496,In_227);
nor U363 (N_363,In_58,In_18);
nand U364 (N_364,In_37,In_395);
nor U365 (N_365,In_158,In_5);
or U366 (N_366,In_47,In_240);
nand U367 (N_367,In_489,In_121);
and U368 (N_368,In_498,In_486);
nand U369 (N_369,In_322,In_400);
nand U370 (N_370,In_202,In_13);
nand U371 (N_371,In_31,In_137);
nor U372 (N_372,In_453,In_25);
nor U373 (N_373,In_400,In_237);
nor U374 (N_374,In_123,In_17);
nor U375 (N_375,In_139,In_494);
nor U376 (N_376,In_241,In_127);
and U377 (N_377,In_275,In_460);
nor U378 (N_378,In_461,In_55);
nand U379 (N_379,In_358,In_11);
nor U380 (N_380,In_83,In_419);
nand U381 (N_381,In_325,In_382);
nand U382 (N_382,In_4,In_295);
nand U383 (N_383,In_483,In_341);
nor U384 (N_384,In_414,In_151);
and U385 (N_385,In_188,In_169);
nand U386 (N_386,In_388,In_188);
or U387 (N_387,In_400,In_379);
nand U388 (N_388,In_139,In_172);
or U389 (N_389,In_161,In_328);
nor U390 (N_390,In_48,In_431);
and U391 (N_391,In_68,In_45);
nor U392 (N_392,In_375,In_16);
nand U393 (N_393,In_153,In_193);
and U394 (N_394,In_369,In_28);
or U395 (N_395,In_190,In_119);
nor U396 (N_396,In_478,In_2);
xor U397 (N_397,In_52,In_346);
xor U398 (N_398,In_359,In_367);
xnor U399 (N_399,In_156,In_260);
and U400 (N_400,In_366,In_218);
or U401 (N_401,In_80,In_334);
nor U402 (N_402,In_238,In_150);
or U403 (N_403,In_473,In_49);
or U404 (N_404,In_421,In_235);
nand U405 (N_405,In_420,In_2);
nor U406 (N_406,In_142,In_238);
nor U407 (N_407,In_63,In_87);
xnor U408 (N_408,In_248,In_108);
or U409 (N_409,In_70,In_378);
and U410 (N_410,In_288,In_296);
nor U411 (N_411,In_168,In_194);
nor U412 (N_412,In_69,In_11);
and U413 (N_413,In_458,In_487);
and U414 (N_414,In_408,In_340);
nor U415 (N_415,In_379,In_55);
nor U416 (N_416,In_258,In_131);
nand U417 (N_417,In_329,In_481);
nand U418 (N_418,In_399,In_437);
and U419 (N_419,In_256,In_249);
or U420 (N_420,In_155,In_340);
nand U421 (N_421,In_316,In_4);
or U422 (N_422,In_446,In_24);
or U423 (N_423,In_182,In_60);
nand U424 (N_424,In_487,In_193);
nor U425 (N_425,In_489,In_328);
nand U426 (N_426,In_320,In_85);
nand U427 (N_427,In_415,In_472);
nor U428 (N_428,In_187,In_124);
xnor U429 (N_429,In_22,In_180);
and U430 (N_430,In_261,In_6);
nand U431 (N_431,In_293,In_138);
nand U432 (N_432,In_386,In_180);
or U433 (N_433,In_52,In_220);
or U434 (N_434,In_218,In_348);
and U435 (N_435,In_120,In_271);
and U436 (N_436,In_325,In_479);
nor U437 (N_437,In_152,In_343);
or U438 (N_438,In_59,In_84);
nand U439 (N_439,In_35,In_476);
and U440 (N_440,In_369,In_240);
nand U441 (N_441,In_209,In_232);
or U442 (N_442,In_379,In_230);
or U443 (N_443,In_148,In_55);
nor U444 (N_444,In_121,In_460);
and U445 (N_445,In_393,In_385);
and U446 (N_446,In_89,In_283);
or U447 (N_447,In_194,In_278);
and U448 (N_448,In_124,In_47);
nor U449 (N_449,In_167,In_16);
and U450 (N_450,In_176,In_82);
or U451 (N_451,In_384,In_354);
nor U452 (N_452,In_74,In_44);
nand U453 (N_453,In_345,In_465);
nand U454 (N_454,In_162,In_461);
nor U455 (N_455,In_161,In_111);
nor U456 (N_456,In_10,In_418);
and U457 (N_457,In_384,In_9);
or U458 (N_458,In_42,In_210);
nor U459 (N_459,In_234,In_8);
or U460 (N_460,In_16,In_242);
or U461 (N_461,In_191,In_142);
nand U462 (N_462,In_4,In_471);
or U463 (N_463,In_144,In_89);
nor U464 (N_464,In_406,In_411);
nand U465 (N_465,In_437,In_398);
and U466 (N_466,In_340,In_259);
nor U467 (N_467,In_376,In_229);
nor U468 (N_468,In_460,In_291);
or U469 (N_469,In_218,In_135);
nor U470 (N_470,In_58,In_380);
and U471 (N_471,In_283,In_200);
nor U472 (N_472,In_177,In_406);
and U473 (N_473,In_453,In_156);
and U474 (N_474,In_89,In_331);
nor U475 (N_475,In_252,In_478);
nor U476 (N_476,In_395,In_120);
and U477 (N_477,In_25,In_243);
or U478 (N_478,In_405,In_187);
or U479 (N_479,In_361,In_464);
and U480 (N_480,In_196,In_223);
or U481 (N_481,In_403,In_13);
or U482 (N_482,In_56,In_439);
or U483 (N_483,In_252,In_153);
nor U484 (N_484,In_163,In_101);
and U485 (N_485,In_98,In_313);
or U486 (N_486,In_327,In_382);
and U487 (N_487,In_441,In_150);
nor U488 (N_488,In_262,In_251);
nor U489 (N_489,In_358,In_380);
nand U490 (N_490,In_128,In_499);
nor U491 (N_491,In_238,In_489);
nor U492 (N_492,In_72,In_481);
nand U493 (N_493,In_278,In_120);
and U494 (N_494,In_250,In_72);
and U495 (N_495,In_146,In_132);
or U496 (N_496,In_153,In_173);
or U497 (N_497,In_74,In_275);
nor U498 (N_498,In_475,In_113);
or U499 (N_499,In_13,In_464);
and U500 (N_500,In_171,In_231);
nand U501 (N_501,In_489,In_57);
nor U502 (N_502,In_494,In_205);
and U503 (N_503,In_365,In_65);
or U504 (N_504,In_272,In_352);
and U505 (N_505,In_48,In_323);
nor U506 (N_506,In_341,In_92);
or U507 (N_507,In_48,In_207);
nor U508 (N_508,In_24,In_451);
or U509 (N_509,In_220,In_300);
or U510 (N_510,In_350,In_307);
nor U511 (N_511,In_264,In_289);
nor U512 (N_512,In_377,In_335);
and U513 (N_513,In_24,In_167);
nand U514 (N_514,In_18,In_73);
nor U515 (N_515,In_19,In_277);
and U516 (N_516,In_468,In_252);
and U517 (N_517,In_59,In_216);
nor U518 (N_518,In_443,In_227);
or U519 (N_519,In_8,In_49);
and U520 (N_520,In_28,In_404);
and U521 (N_521,In_355,In_457);
nor U522 (N_522,In_374,In_8);
nor U523 (N_523,In_153,In_124);
or U524 (N_524,In_365,In_433);
nor U525 (N_525,In_101,In_165);
nand U526 (N_526,In_282,In_305);
xnor U527 (N_527,In_105,In_122);
and U528 (N_528,In_493,In_488);
nor U529 (N_529,In_441,In_235);
and U530 (N_530,In_316,In_278);
or U531 (N_531,In_181,In_355);
and U532 (N_532,In_248,In_376);
nor U533 (N_533,In_188,In_303);
and U534 (N_534,In_375,In_103);
xnor U535 (N_535,In_268,In_179);
nand U536 (N_536,In_226,In_379);
nand U537 (N_537,In_133,In_173);
or U538 (N_538,In_199,In_391);
or U539 (N_539,In_327,In_95);
nor U540 (N_540,In_360,In_231);
nand U541 (N_541,In_497,In_18);
nor U542 (N_542,In_8,In_350);
and U543 (N_543,In_114,In_212);
nand U544 (N_544,In_313,In_83);
nor U545 (N_545,In_197,In_177);
nand U546 (N_546,In_104,In_293);
and U547 (N_547,In_205,In_203);
nand U548 (N_548,In_64,In_19);
nor U549 (N_549,In_65,In_320);
or U550 (N_550,In_363,In_69);
nand U551 (N_551,In_84,In_448);
nor U552 (N_552,In_71,In_419);
and U553 (N_553,In_299,In_337);
nor U554 (N_554,In_162,In_452);
nand U555 (N_555,In_352,In_122);
or U556 (N_556,In_370,In_166);
xnor U557 (N_557,In_486,In_53);
or U558 (N_558,In_330,In_204);
or U559 (N_559,In_103,In_249);
or U560 (N_560,In_410,In_384);
and U561 (N_561,In_332,In_230);
and U562 (N_562,In_308,In_426);
and U563 (N_563,In_337,In_329);
or U564 (N_564,In_33,In_382);
and U565 (N_565,In_407,In_285);
and U566 (N_566,In_31,In_441);
nor U567 (N_567,In_203,In_86);
or U568 (N_568,In_417,In_435);
and U569 (N_569,In_83,In_269);
nor U570 (N_570,In_287,In_253);
and U571 (N_571,In_442,In_83);
and U572 (N_572,In_253,In_264);
or U573 (N_573,In_140,In_294);
and U574 (N_574,In_53,In_253);
and U575 (N_575,In_175,In_223);
nand U576 (N_576,In_301,In_120);
or U577 (N_577,In_408,In_24);
or U578 (N_578,In_9,In_399);
or U579 (N_579,In_226,In_446);
and U580 (N_580,In_10,In_50);
and U581 (N_581,In_324,In_491);
xnor U582 (N_582,In_454,In_406);
or U583 (N_583,In_439,In_255);
and U584 (N_584,In_488,In_236);
or U585 (N_585,In_471,In_66);
nor U586 (N_586,In_312,In_32);
and U587 (N_587,In_142,In_182);
and U588 (N_588,In_251,In_6);
nor U589 (N_589,In_376,In_340);
and U590 (N_590,In_324,In_430);
and U591 (N_591,In_38,In_433);
nor U592 (N_592,In_121,In_40);
and U593 (N_593,In_294,In_302);
nor U594 (N_594,In_64,In_195);
xor U595 (N_595,In_481,In_237);
nand U596 (N_596,In_230,In_98);
nand U597 (N_597,In_36,In_358);
or U598 (N_598,In_102,In_417);
or U599 (N_599,In_167,In_399);
nand U600 (N_600,In_176,In_110);
nor U601 (N_601,In_194,In_255);
or U602 (N_602,In_281,In_167);
nand U603 (N_603,In_469,In_50);
and U604 (N_604,In_138,In_420);
nor U605 (N_605,In_204,In_153);
or U606 (N_606,In_469,In_47);
nor U607 (N_607,In_69,In_416);
and U608 (N_608,In_159,In_412);
nand U609 (N_609,In_38,In_286);
nor U610 (N_610,In_132,In_9);
nor U611 (N_611,In_257,In_253);
nor U612 (N_612,In_290,In_310);
and U613 (N_613,In_418,In_346);
nand U614 (N_614,In_88,In_82);
nand U615 (N_615,In_139,In_232);
nand U616 (N_616,In_37,In_143);
and U617 (N_617,In_488,In_185);
nor U618 (N_618,In_365,In_135);
or U619 (N_619,In_253,In_148);
nand U620 (N_620,In_363,In_74);
nor U621 (N_621,In_200,In_169);
nor U622 (N_622,In_254,In_465);
and U623 (N_623,In_337,In_346);
and U624 (N_624,In_405,In_151);
nor U625 (N_625,In_490,In_177);
or U626 (N_626,In_11,In_308);
and U627 (N_627,In_402,In_278);
nor U628 (N_628,In_94,In_68);
or U629 (N_629,In_486,In_32);
nor U630 (N_630,In_33,In_232);
or U631 (N_631,In_241,In_485);
nand U632 (N_632,In_336,In_57);
and U633 (N_633,In_460,In_426);
or U634 (N_634,In_160,In_279);
or U635 (N_635,In_249,In_499);
or U636 (N_636,In_127,In_55);
and U637 (N_637,In_121,In_380);
nor U638 (N_638,In_174,In_130);
and U639 (N_639,In_107,In_408);
or U640 (N_640,In_289,In_277);
xnor U641 (N_641,In_192,In_418);
nand U642 (N_642,In_298,In_457);
xor U643 (N_643,In_328,In_492);
or U644 (N_644,In_261,In_190);
or U645 (N_645,In_497,In_354);
nand U646 (N_646,In_407,In_232);
nand U647 (N_647,In_31,In_245);
and U648 (N_648,In_19,In_223);
nor U649 (N_649,In_28,In_206);
nor U650 (N_650,In_324,In_147);
nand U651 (N_651,In_345,In_460);
xor U652 (N_652,In_148,In_189);
or U653 (N_653,In_90,In_176);
or U654 (N_654,In_373,In_290);
nand U655 (N_655,In_151,In_400);
nand U656 (N_656,In_210,In_341);
and U657 (N_657,In_25,In_434);
and U658 (N_658,In_292,In_167);
or U659 (N_659,In_290,In_114);
nor U660 (N_660,In_51,In_341);
or U661 (N_661,In_379,In_3);
or U662 (N_662,In_471,In_382);
and U663 (N_663,In_195,In_148);
nand U664 (N_664,In_299,In_484);
and U665 (N_665,In_216,In_475);
nor U666 (N_666,In_198,In_68);
nand U667 (N_667,In_470,In_303);
and U668 (N_668,In_382,In_6);
nor U669 (N_669,In_212,In_338);
and U670 (N_670,In_406,In_287);
nand U671 (N_671,In_34,In_54);
or U672 (N_672,In_68,In_71);
and U673 (N_673,In_117,In_436);
or U674 (N_674,In_245,In_157);
nor U675 (N_675,In_429,In_287);
nor U676 (N_676,In_403,In_20);
nor U677 (N_677,In_322,In_404);
or U678 (N_678,In_270,In_481);
nor U679 (N_679,In_448,In_261);
nor U680 (N_680,In_447,In_445);
nand U681 (N_681,In_485,In_31);
nor U682 (N_682,In_369,In_153);
nand U683 (N_683,In_476,In_444);
or U684 (N_684,In_493,In_135);
nand U685 (N_685,In_225,In_437);
and U686 (N_686,In_478,In_318);
nand U687 (N_687,In_248,In_197);
nor U688 (N_688,In_247,In_408);
xnor U689 (N_689,In_469,In_319);
or U690 (N_690,In_497,In_85);
or U691 (N_691,In_22,In_441);
xor U692 (N_692,In_24,In_339);
and U693 (N_693,In_283,In_9);
or U694 (N_694,In_487,In_212);
or U695 (N_695,In_263,In_252);
or U696 (N_696,In_280,In_32);
and U697 (N_697,In_52,In_374);
nor U698 (N_698,In_311,In_170);
nand U699 (N_699,In_212,In_446);
nand U700 (N_700,In_414,In_281);
nor U701 (N_701,In_32,In_64);
nor U702 (N_702,In_289,In_324);
and U703 (N_703,In_321,In_101);
and U704 (N_704,In_185,In_434);
nand U705 (N_705,In_486,In_275);
and U706 (N_706,In_8,In_130);
and U707 (N_707,In_286,In_306);
and U708 (N_708,In_333,In_148);
or U709 (N_709,In_70,In_277);
nor U710 (N_710,In_193,In_295);
and U711 (N_711,In_296,In_353);
and U712 (N_712,In_332,In_408);
nor U713 (N_713,In_208,In_180);
or U714 (N_714,In_178,In_330);
nand U715 (N_715,In_22,In_414);
nand U716 (N_716,In_309,In_304);
and U717 (N_717,In_218,In_385);
xor U718 (N_718,In_224,In_349);
nor U719 (N_719,In_274,In_438);
nand U720 (N_720,In_56,In_321);
nor U721 (N_721,In_278,In_323);
nor U722 (N_722,In_65,In_396);
and U723 (N_723,In_31,In_229);
or U724 (N_724,In_310,In_241);
nand U725 (N_725,In_97,In_355);
nand U726 (N_726,In_369,In_185);
and U727 (N_727,In_279,In_105);
and U728 (N_728,In_10,In_261);
and U729 (N_729,In_348,In_115);
nor U730 (N_730,In_153,In_387);
and U731 (N_731,In_53,In_217);
or U732 (N_732,In_339,In_444);
xor U733 (N_733,In_239,In_144);
nor U734 (N_734,In_137,In_53);
or U735 (N_735,In_30,In_94);
nor U736 (N_736,In_201,In_429);
nand U737 (N_737,In_344,In_203);
nand U738 (N_738,In_77,In_265);
nand U739 (N_739,In_99,In_440);
or U740 (N_740,In_410,In_465);
and U741 (N_741,In_357,In_377);
xnor U742 (N_742,In_365,In_376);
nand U743 (N_743,In_378,In_32);
nand U744 (N_744,In_224,In_499);
or U745 (N_745,In_183,In_174);
nor U746 (N_746,In_286,In_256);
or U747 (N_747,In_179,In_117);
or U748 (N_748,In_316,In_5);
nand U749 (N_749,In_286,In_184);
or U750 (N_750,In_242,In_107);
nor U751 (N_751,In_114,In_224);
nor U752 (N_752,In_154,In_234);
and U753 (N_753,In_263,In_340);
nand U754 (N_754,In_342,In_48);
and U755 (N_755,In_362,In_281);
or U756 (N_756,In_454,In_495);
nor U757 (N_757,In_212,In_130);
and U758 (N_758,In_120,In_451);
or U759 (N_759,In_331,In_211);
nor U760 (N_760,In_494,In_383);
and U761 (N_761,In_92,In_115);
or U762 (N_762,In_19,In_283);
nor U763 (N_763,In_3,In_329);
nand U764 (N_764,In_289,In_311);
nor U765 (N_765,In_404,In_146);
nor U766 (N_766,In_23,In_333);
nor U767 (N_767,In_161,In_225);
nor U768 (N_768,In_351,In_170);
nor U769 (N_769,In_319,In_396);
and U770 (N_770,In_411,In_497);
nand U771 (N_771,In_473,In_126);
nand U772 (N_772,In_109,In_28);
nand U773 (N_773,In_228,In_32);
xor U774 (N_774,In_264,In_213);
and U775 (N_775,In_0,In_454);
or U776 (N_776,In_394,In_375);
and U777 (N_777,In_61,In_232);
nor U778 (N_778,In_292,In_335);
or U779 (N_779,In_16,In_131);
nor U780 (N_780,In_32,In_388);
nand U781 (N_781,In_331,In_277);
or U782 (N_782,In_117,In_454);
or U783 (N_783,In_335,In_7);
nor U784 (N_784,In_277,In_3);
xor U785 (N_785,In_380,In_394);
or U786 (N_786,In_78,In_95);
or U787 (N_787,In_130,In_185);
xnor U788 (N_788,In_171,In_256);
or U789 (N_789,In_73,In_157);
or U790 (N_790,In_286,In_200);
nand U791 (N_791,In_60,In_150);
and U792 (N_792,In_27,In_346);
nor U793 (N_793,In_395,In_490);
xnor U794 (N_794,In_486,In_31);
nand U795 (N_795,In_281,In_328);
nor U796 (N_796,In_459,In_259);
or U797 (N_797,In_196,In_333);
or U798 (N_798,In_181,In_346);
nand U799 (N_799,In_394,In_214);
and U800 (N_800,In_443,In_112);
nand U801 (N_801,In_71,In_73);
nand U802 (N_802,In_147,In_408);
or U803 (N_803,In_451,In_418);
and U804 (N_804,In_392,In_485);
nor U805 (N_805,In_363,In_317);
or U806 (N_806,In_100,In_287);
nor U807 (N_807,In_442,In_152);
or U808 (N_808,In_71,In_470);
nand U809 (N_809,In_335,In_374);
nor U810 (N_810,In_252,In_186);
and U811 (N_811,In_93,In_366);
xnor U812 (N_812,In_179,In_473);
or U813 (N_813,In_98,In_87);
and U814 (N_814,In_107,In_328);
nand U815 (N_815,In_320,In_372);
or U816 (N_816,In_151,In_29);
nor U817 (N_817,In_329,In_207);
or U818 (N_818,In_122,In_447);
nor U819 (N_819,In_197,In_120);
or U820 (N_820,In_343,In_131);
and U821 (N_821,In_302,In_444);
nor U822 (N_822,In_138,In_27);
nor U823 (N_823,In_238,In_35);
nor U824 (N_824,In_272,In_491);
and U825 (N_825,In_481,In_10);
and U826 (N_826,In_458,In_228);
nand U827 (N_827,In_184,In_35);
nand U828 (N_828,In_32,In_95);
and U829 (N_829,In_112,In_243);
nand U830 (N_830,In_151,In_418);
nand U831 (N_831,In_155,In_338);
nor U832 (N_832,In_184,In_478);
nor U833 (N_833,In_160,In_476);
or U834 (N_834,In_102,In_320);
or U835 (N_835,In_255,In_262);
nand U836 (N_836,In_369,In_363);
and U837 (N_837,In_260,In_30);
nor U838 (N_838,In_449,In_58);
xor U839 (N_839,In_396,In_337);
nor U840 (N_840,In_0,In_22);
and U841 (N_841,In_7,In_193);
nor U842 (N_842,In_361,In_307);
nand U843 (N_843,In_63,In_339);
and U844 (N_844,In_408,In_421);
nor U845 (N_845,In_177,In_193);
nand U846 (N_846,In_371,In_402);
nor U847 (N_847,In_39,In_488);
nor U848 (N_848,In_160,In_425);
or U849 (N_849,In_302,In_296);
or U850 (N_850,In_249,In_218);
nand U851 (N_851,In_1,In_175);
nand U852 (N_852,In_322,In_137);
nor U853 (N_853,In_170,In_73);
nor U854 (N_854,In_315,In_267);
or U855 (N_855,In_342,In_105);
nor U856 (N_856,In_298,In_56);
nand U857 (N_857,In_440,In_141);
or U858 (N_858,In_496,In_494);
nand U859 (N_859,In_93,In_484);
or U860 (N_860,In_459,In_41);
nand U861 (N_861,In_224,In_330);
or U862 (N_862,In_74,In_303);
nor U863 (N_863,In_147,In_153);
and U864 (N_864,In_114,In_102);
and U865 (N_865,In_453,In_23);
or U866 (N_866,In_201,In_147);
nand U867 (N_867,In_41,In_212);
nor U868 (N_868,In_397,In_374);
and U869 (N_869,In_362,In_174);
or U870 (N_870,In_241,In_462);
nor U871 (N_871,In_85,In_464);
nand U872 (N_872,In_211,In_150);
or U873 (N_873,In_99,In_110);
nand U874 (N_874,In_439,In_187);
and U875 (N_875,In_338,In_230);
and U876 (N_876,In_40,In_471);
nand U877 (N_877,In_337,In_258);
and U878 (N_878,In_479,In_268);
nand U879 (N_879,In_106,In_227);
or U880 (N_880,In_353,In_198);
nor U881 (N_881,In_250,In_491);
or U882 (N_882,In_309,In_292);
or U883 (N_883,In_167,In_154);
nand U884 (N_884,In_161,In_425);
nand U885 (N_885,In_217,In_164);
and U886 (N_886,In_351,In_133);
or U887 (N_887,In_173,In_185);
nand U888 (N_888,In_415,In_414);
nor U889 (N_889,In_475,In_273);
nor U890 (N_890,In_297,In_198);
nand U891 (N_891,In_211,In_433);
nand U892 (N_892,In_40,In_360);
nor U893 (N_893,In_484,In_292);
nor U894 (N_894,In_317,In_479);
nand U895 (N_895,In_72,In_123);
nand U896 (N_896,In_10,In_371);
nor U897 (N_897,In_26,In_122);
nor U898 (N_898,In_468,In_421);
nand U899 (N_899,In_75,In_437);
nand U900 (N_900,In_21,In_68);
nor U901 (N_901,In_416,In_6);
nand U902 (N_902,In_96,In_50);
and U903 (N_903,In_67,In_91);
and U904 (N_904,In_499,In_404);
or U905 (N_905,In_221,In_63);
nor U906 (N_906,In_167,In_178);
or U907 (N_907,In_277,In_446);
nand U908 (N_908,In_441,In_213);
and U909 (N_909,In_371,In_83);
nand U910 (N_910,In_134,In_405);
and U911 (N_911,In_289,In_321);
nand U912 (N_912,In_239,In_378);
nor U913 (N_913,In_378,In_414);
and U914 (N_914,In_258,In_297);
nand U915 (N_915,In_241,In_153);
and U916 (N_916,In_2,In_359);
nor U917 (N_917,In_38,In_453);
and U918 (N_918,In_76,In_38);
or U919 (N_919,In_8,In_9);
and U920 (N_920,In_109,In_148);
nand U921 (N_921,In_209,In_412);
or U922 (N_922,In_467,In_14);
or U923 (N_923,In_185,In_94);
nor U924 (N_924,In_380,In_31);
and U925 (N_925,In_372,In_450);
nor U926 (N_926,In_60,In_294);
nand U927 (N_927,In_137,In_420);
nor U928 (N_928,In_373,In_51);
or U929 (N_929,In_290,In_223);
and U930 (N_930,In_380,In_161);
nand U931 (N_931,In_250,In_235);
nor U932 (N_932,In_161,In_260);
and U933 (N_933,In_439,In_153);
nor U934 (N_934,In_217,In_102);
and U935 (N_935,In_361,In_447);
nor U936 (N_936,In_115,In_241);
nor U937 (N_937,In_189,In_104);
and U938 (N_938,In_123,In_303);
or U939 (N_939,In_486,In_89);
and U940 (N_940,In_177,In_176);
nor U941 (N_941,In_65,In_69);
or U942 (N_942,In_392,In_255);
and U943 (N_943,In_202,In_83);
and U944 (N_944,In_46,In_443);
nand U945 (N_945,In_289,In_4);
or U946 (N_946,In_290,In_192);
nand U947 (N_947,In_26,In_351);
and U948 (N_948,In_321,In_136);
nand U949 (N_949,In_385,In_198);
nor U950 (N_950,In_390,In_313);
nor U951 (N_951,In_132,In_136);
and U952 (N_952,In_86,In_285);
or U953 (N_953,In_425,In_132);
and U954 (N_954,In_161,In_327);
nand U955 (N_955,In_178,In_387);
nand U956 (N_956,In_260,In_216);
nand U957 (N_957,In_10,In_307);
and U958 (N_958,In_408,In_150);
or U959 (N_959,In_360,In_383);
nand U960 (N_960,In_369,In_7);
or U961 (N_961,In_493,In_132);
and U962 (N_962,In_330,In_171);
nor U963 (N_963,In_490,In_462);
nand U964 (N_964,In_109,In_293);
nor U965 (N_965,In_135,In_81);
or U966 (N_966,In_243,In_279);
nand U967 (N_967,In_110,In_16);
xor U968 (N_968,In_73,In_242);
or U969 (N_969,In_186,In_204);
and U970 (N_970,In_298,In_132);
nor U971 (N_971,In_61,In_408);
and U972 (N_972,In_391,In_157);
or U973 (N_973,In_491,In_43);
nand U974 (N_974,In_284,In_334);
nor U975 (N_975,In_269,In_183);
nor U976 (N_976,In_217,In_435);
or U977 (N_977,In_152,In_341);
xor U978 (N_978,In_64,In_265);
or U979 (N_979,In_183,In_251);
xnor U980 (N_980,In_102,In_198);
and U981 (N_981,In_247,In_360);
or U982 (N_982,In_232,In_470);
nor U983 (N_983,In_123,In_99);
or U984 (N_984,In_246,In_314);
nand U985 (N_985,In_431,In_254);
nand U986 (N_986,In_328,In_204);
and U987 (N_987,In_56,In_292);
nand U988 (N_988,In_262,In_470);
nand U989 (N_989,In_400,In_219);
and U990 (N_990,In_370,In_430);
and U991 (N_991,In_477,In_476);
nor U992 (N_992,In_425,In_252);
nand U993 (N_993,In_455,In_388);
or U994 (N_994,In_8,In_59);
nand U995 (N_995,In_489,In_484);
or U996 (N_996,In_20,In_370);
or U997 (N_997,In_445,In_218);
or U998 (N_998,In_287,In_390);
nor U999 (N_999,In_248,In_4);
nand U1000 (N_1000,N_696,N_290);
nor U1001 (N_1001,N_993,N_951);
and U1002 (N_1002,N_816,N_37);
nor U1003 (N_1003,N_843,N_33);
nand U1004 (N_1004,N_525,N_40);
xnor U1005 (N_1005,N_3,N_540);
and U1006 (N_1006,N_679,N_336);
or U1007 (N_1007,N_957,N_315);
nand U1008 (N_1008,N_443,N_975);
or U1009 (N_1009,N_304,N_57);
nand U1010 (N_1010,N_420,N_846);
nor U1011 (N_1011,N_994,N_481);
nand U1012 (N_1012,N_681,N_647);
nand U1013 (N_1013,N_902,N_952);
xnor U1014 (N_1014,N_464,N_573);
or U1015 (N_1015,N_882,N_175);
or U1016 (N_1016,N_365,N_193);
nor U1017 (N_1017,N_91,N_161);
or U1018 (N_1018,N_276,N_463);
nor U1019 (N_1019,N_163,N_865);
and U1020 (N_1020,N_36,N_185);
and U1021 (N_1021,N_270,N_432);
and U1022 (N_1022,N_666,N_367);
nor U1023 (N_1023,N_318,N_296);
or U1024 (N_1024,N_947,N_845);
and U1025 (N_1025,N_724,N_285);
nand U1026 (N_1026,N_55,N_76);
nand U1027 (N_1027,N_383,N_140);
nand U1028 (N_1028,N_486,N_418);
xor U1029 (N_1029,N_65,N_563);
nor U1030 (N_1030,N_179,N_965);
nand U1031 (N_1031,N_349,N_38);
or U1032 (N_1032,N_901,N_8);
or U1033 (N_1033,N_580,N_321);
or U1034 (N_1034,N_803,N_457);
nor U1035 (N_1035,N_919,N_243);
xnor U1036 (N_1036,N_415,N_654);
nor U1037 (N_1037,N_257,N_222);
and U1038 (N_1038,N_303,N_670);
and U1039 (N_1039,N_271,N_949);
and U1040 (N_1040,N_896,N_472);
and U1041 (N_1041,N_95,N_967);
nand U1042 (N_1042,N_279,N_305);
and U1043 (N_1043,N_103,N_268);
or U1044 (N_1044,N_160,N_519);
nand U1045 (N_1045,N_876,N_748);
nand U1046 (N_1046,N_483,N_593);
and U1047 (N_1047,N_796,N_559);
nor U1048 (N_1048,N_466,N_578);
and U1049 (N_1049,N_314,N_135);
or U1050 (N_1050,N_604,N_996);
nand U1051 (N_1051,N_810,N_391);
and U1052 (N_1052,N_785,N_821);
and U1053 (N_1053,N_599,N_379);
and U1054 (N_1054,N_62,N_797);
nand U1055 (N_1055,N_572,N_564);
and U1056 (N_1056,N_515,N_799);
and U1057 (N_1057,N_783,N_671);
nand U1058 (N_1058,N_212,N_216);
nor U1059 (N_1059,N_207,N_12);
and U1060 (N_1060,N_849,N_120);
nand U1061 (N_1061,N_206,N_399);
and U1062 (N_1062,N_266,N_406);
or U1063 (N_1063,N_200,N_489);
and U1064 (N_1064,N_149,N_125);
nand U1065 (N_1065,N_422,N_780);
or U1066 (N_1066,N_236,N_98);
nand U1067 (N_1067,N_292,N_310);
nor U1068 (N_1068,N_475,N_982);
nor U1069 (N_1069,N_348,N_706);
nand U1070 (N_1070,N_337,N_112);
or U1071 (N_1071,N_789,N_790);
nand U1072 (N_1072,N_289,N_755);
nand U1073 (N_1073,N_771,N_259);
or U1074 (N_1074,N_128,N_491);
nor U1075 (N_1075,N_754,N_827);
nand U1076 (N_1076,N_743,N_832);
nor U1077 (N_1077,N_150,N_746);
nor U1078 (N_1078,N_499,N_211);
or U1079 (N_1079,N_824,N_508);
or U1080 (N_1080,N_946,N_675);
nor U1081 (N_1081,N_447,N_482);
nor U1082 (N_1082,N_809,N_232);
and U1083 (N_1083,N_116,N_351);
and U1084 (N_1084,N_1,N_977);
or U1085 (N_1085,N_465,N_644);
and U1086 (N_1086,N_403,N_145);
nor U1087 (N_1087,N_496,N_888);
or U1088 (N_1088,N_721,N_807);
nor U1089 (N_1089,N_998,N_115);
and U1090 (N_1090,N_963,N_651);
nand U1091 (N_1091,N_494,N_238);
and U1092 (N_1092,N_411,N_386);
nand U1093 (N_1093,N_948,N_543);
and U1094 (N_1094,N_246,N_56);
nor U1095 (N_1095,N_283,N_219);
nand U1096 (N_1096,N_772,N_583);
or U1097 (N_1097,N_278,N_579);
or U1098 (N_1098,N_134,N_920);
nor U1099 (N_1099,N_421,N_388);
nor U1100 (N_1100,N_68,N_931);
nand U1101 (N_1101,N_610,N_417);
or U1102 (N_1102,N_495,N_766);
nand U1103 (N_1103,N_669,N_7);
nand U1104 (N_1104,N_22,N_374);
or U1105 (N_1105,N_132,N_717);
nand U1106 (N_1106,N_362,N_42);
nor U1107 (N_1107,N_822,N_467);
and U1108 (N_1108,N_284,N_446);
nand U1109 (N_1109,N_445,N_894);
nand U1110 (N_1110,N_369,N_184);
nor U1111 (N_1111,N_646,N_554);
and U1112 (N_1112,N_682,N_879);
and U1113 (N_1113,N_926,N_237);
and U1114 (N_1114,N_356,N_209);
or U1115 (N_1115,N_917,N_177);
nand U1116 (N_1116,N_829,N_455);
nor U1117 (N_1117,N_102,N_652);
nand U1118 (N_1118,N_277,N_758);
and U1119 (N_1119,N_565,N_195);
and U1120 (N_1120,N_923,N_908);
nand U1121 (N_1121,N_172,N_428);
or U1122 (N_1122,N_251,N_661);
and U1123 (N_1123,N_286,N_871);
or U1124 (N_1124,N_781,N_956);
and U1125 (N_1125,N_518,N_954);
or U1126 (N_1126,N_479,N_619);
nand U1127 (N_1127,N_714,N_205);
or U1128 (N_1128,N_630,N_970);
or U1129 (N_1129,N_761,N_964);
nand U1130 (N_1130,N_312,N_69);
nand U1131 (N_1131,N_59,N_794);
or U1132 (N_1132,N_587,N_995);
and U1133 (N_1133,N_897,N_676);
or U1134 (N_1134,N_823,N_503);
nand U1135 (N_1135,N_181,N_439);
nor U1136 (N_1136,N_744,N_690);
and U1137 (N_1137,N_123,N_106);
nand U1138 (N_1138,N_659,N_942);
or U1139 (N_1139,N_155,N_941);
or U1140 (N_1140,N_224,N_441);
or U1141 (N_1141,N_886,N_101);
nand U1142 (N_1142,N_689,N_168);
xor U1143 (N_1143,N_493,N_512);
and U1144 (N_1144,N_297,N_906);
nor U1145 (N_1145,N_333,N_74);
nand U1146 (N_1146,N_334,N_19);
or U1147 (N_1147,N_176,N_932);
xnor U1148 (N_1148,N_364,N_358);
nor U1149 (N_1149,N_633,N_698);
xnor U1150 (N_1150,N_950,N_427);
or U1151 (N_1151,N_857,N_387);
or U1152 (N_1152,N_215,N_380);
or U1153 (N_1153,N_301,N_838);
or U1154 (N_1154,N_786,N_294);
nand U1155 (N_1155,N_450,N_987);
nor U1156 (N_1156,N_9,N_30);
nor U1157 (N_1157,N_914,N_751);
and U1158 (N_1158,N_288,N_608);
nor U1159 (N_1159,N_171,N_89);
and U1160 (N_1160,N_117,N_371);
and U1161 (N_1161,N_250,N_384);
nor U1162 (N_1162,N_597,N_672);
or U1163 (N_1163,N_342,N_320);
or U1164 (N_1164,N_108,N_504);
and U1165 (N_1165,N_739,N_858);
or U1166 (N_1166,N_426,N_598);
or U1167 (N_1167,N_298,N_861);
xnor U1168 (N_1168,N_221,N_770);
xor U1169 (N_1169,N_187,N_104);
or U1170 (N_1170,N_353,N_183);
and U1171 (N_1171,N_873,N_900);
nor U1172 (N_1172,N_694,N_93);
xnor U1173 (N_1173,N_622,N_174);
nor U1174 (N_1174,N_958,N_21);
and U1175 (N_1175,N_940,N_892);
and U1176 (N_1176,N_24,N_462);
nand U1177 (N_1177,N_898,N_801);
or U1178 (N_1178,N_686,N_359);
nand U1179 (N_1179,N_524,N_50);
nand U1180 (N_1180,N_156,N_264);
nand U1181 (N_1181,N_992,N_667);
or U1182 (N_1182,N_685,N_971);
nor U1183 (N_1183,N_620,N_204);
and U1184 (N_1184,N_726,N_444);
nand U1185 (N_1185,N_955,N_84);
nor U1186 (N_1186,N_96,N_627);
or U1187 (N_1187,N_368,N_167);
nor U1188 (N_1188,N_144,N_930);
nand U1189 (N_1189,N_71,N_614);
and U1190 (N_1190,N_642,N_571);
nand U1191 (N_1191,N_976,N_759);
or U1192 (N_1192,N_64,N_859);
or U1193 (N_1193,N_557,N_601);
or U1194 (N_1194,N_710,N_602);
or U1195 (N_1195,N_146,N_805);
nand U1196 (N_1196,N_373,N_352);
nor U1197 (N_1197,N_695,N_773);
or U1198 (N_1198,N_402,N_198);
and U1199 (N_1199,N_634,N_332);
nor U1200 (N_1200,N_966,N_86);
nor U1201 (N_1201,N_566,N_850);
nor U1202 (N_1202,N_953,N_727);
nor U1203 (N_1203,N_984,N_138);
or U1204 (N_1204,N_874,N_66);
nand U1205 (N_1205,N_218,N_723);
nand U1206 (N_1206,N_887,N_247);
and U1207 (N_1207,N_319,N_32);
nor U1208 (N_1208,N_983,N_506);
xor U1209 (N_1209,N_560,N_784);
and U1210 (N_1210,N_707,N_507);
or U1211 (N_1211,N_99,N_749);
nor U1212 (N_1212,N_110,N_728);
nor U1213 (N_1213,N_511,N_860);
and U1214 (N_1214,N_733,N_961);
or U1215 (N_1215,N_502,N_862);
nor U1216 (N_1216,N_490,N_330);
and U1217 (N_1217,N_613,N_664);
nor U1218 (N_1218,N_164,N_648);
nor U1219 (N_1219,N_615,N_818);
nand U1220 (N_1220,N_631,N_347);
or U1221 (N_1221,N_63,N_891);
nand U1222 (N_1222,N_210,N_480);
or U1223 (N_1223,N_67,N_35);
or U1224 (N_1224,N_692,N_223);
or U1225 (N_1225,N_229,N_324);
nor U1226 (N_1226,N_28,N_338);
or U1227 (N_1227,N_122,N_2);
and U1228 (N_1228,N_189,N_233);
nor U1229 (N_1229,N_485,N_878);
or U1230 (N_1230,N_737,N_814);
nand U1231 (N_1231,N_550,N_354);
or U1232 (N_1232,N_159,N_881);
nor U1233 (N_1233,N_684,N_335);
nor U1234 (N_1234,N_513,N_972);
and U1235 (N_1235,N_699,N_662);
nand U1236 (N_1236,N_768,N_867);
and U1237 (N_1237,N_655,N_641);
or U1238 (N_1238,N_49,N_582);
and U1239 (N_1239,N_239,N_214);
nor U1240 (N_1240,N_812,N_774);
or U1241 (N_1241,N_302,N_968);
and U1242 (N_1242,N_173,N_649);
nand U1243 (N_1243,N_416,N_741);
nor U1244 (N_1244,N_468,N_637);
or U1245 (N_1245,N_327,N_742);
nor U1246 (N_1246,N_703,N_309);
nand U1247 (N_1247,N_653,N_510);
or U1248 (N_1248,N_273,N_716);
and U1249 (N_1249,N_747,N_488);
and U1250 (N_1250,N_640,N_830);
nand U1251 (N_1251,N_718,N_474);
nor U1252 (N_1252,N_985,N_708);
nand U1253 (N_1253,N_817,N_568);
nor U1254 (N_1254,N_575,N_322);
and U1255 (N_1255,N_558,N_555);
or U1256 (N_1256,N_46,N_562);
or U1257 (N_1257,N_680,N_272);
nand U1258 (N_1258,N_750,N_178);
and U1259 (N_1259,N_851,N_197);
nor U1260 (N_1260,N_663,N_521);
nor U1261 (N_1261,N_240,N_889);
or U1262 (N_1262,N_847,N_346);
and U1263 (N_1263,N_139,N_325);
nor U1264 (N_1264,N_413,N_643);
or U1265 (N_1265,N_267,N_552);
nand U1266 (N_1266,N_492,N_788);
nand U1267 (N_1267,N_539,N_170);
or U1268 (N_1268,N_248,N_884);
nand U1269 (N_1269,N_143,N_944);
nand U1270 (N_1270,N_147,N_561);
or U1271 (N_1271,N_438,N_722);
and U1272 (N_1272,N_517,N_712);
or U1273 (N_1273,N_188,N_393);
and U1274 (N_1274,N_460,N_25);
nand U1275 (N_1275,N_603,N_905);
nand U1276 (N_1276,N_855,N_574);
and U1277 (N_1277,N_196,N_409);
nor U1278 (N_1278,N_734,N_126);
nand U1279 (N_1279,N_839,N_311);
or U1280 (N_1280,N_429,N_18);
or U1281 (N_1281,N_280,N_77);
nor U1282 (N_1282,N_629,N_945);
nand U1283 (N_1283,N_757,N_624);
or U1284 (N_1284,N_545,N_704);
nand U1285 (N_1285,N_804,N_343);
or U1286 (N_1286,N_674,N_530);
or U1287 (N_1287,N_43,N_534);
xnor U1288 (N_1288,N_300,N_235);
nand U1289 (N_1289,N_78,N_591);
nand U1290 (N_1290,N_153,N_922);
nor U1291 (N_1291,N_526,N_589);
nand U1292 (N_1292,N_841,N_124);
nor U1293 (N_1293,N_505,N_787);
nor U1294 (N_1294,N_192,N_85);
and U1295 (N_1295,N_870,N_0);
or U1296 (N_1296,N_535,N_618);
or U1297 (N_1297,N_638,N_244);
or U1298 (N_1298,N_114,N_933);
nor U1299 (N_1299,N_339,N_133);
xnor U1300 (N_1300,N_433,N_806);
or U1301 (N_1301,N_570,N_828);
and U1302 (N_1302,N_606,N_825);
and U1303 (N_1303,N_736,N_454);
or U1304 (N_1304,N_678,N_350);
nor U1305 (N_1305,N_72,N_732);
or U1306 (N_1306,N_281,N_997);
nand U1307 (N_1307,N_20,N_390);
or U1308 (N_1308,N_740,N_793);
or U1309 (N_1309,N_645,N_844);
or U1310 (N_1310,N_92,N_255);
and U1311 (N_1311,N_725,N_201);
nand U1312 (N_1312,N_478,N_58);
nand U1313 (N_1313,N_656,N_476);
and U1314 (N_1314,N_498,N_668);
and U1315 (N_1315,N_893,N_735);
nor U1316 (N_1316,N_231,N_912);
and U1317 (N_1317,N_107,N_811);
nor U1318 (N_1318,N_414,N_595);
and U1319 (N_1319,N_317,N_226);
nand U1320 (N_1320,N_73,N_826);
nand U1321 (N_1321,N_911,N_693);
and U1322 (N_1322,N_375,N_854);
or U1323 (N_1323,N_962,N_131);
nor U1324 (N_1324,N_306,N_556);
nand U1325 (N_1325,N_600,N_431);
and U1326 (N_1326,N_628,N_394);
nand U1327 (N_1327,N_842,N_111);
and U1328 (N_1328,N_477,N_592);
nor U1329 (N_1329,N_451,N_180);
nand U1330 (N_1330,N_875,N_756);
nand U1331 (N_1331,N_398,N_657);
and U1332 (N_1332,N_316,N_75);
and U1333 (N_1333,N_121,N_899);
nand U1334 (N_1334,N_528,N_609);
nand U1335 (N_1335,N_396,N_54);
nor U1336 (N_1336,N_590,N_500);
and U1337 (N_1337,N_199,N_711);
and U1338 (N_1338,N_228,N_400);
nor U1339 (N_1339,N_127,N_864);
or U1340 (N_1340,N_925,N_863);
and U1341 (N_1341,N_872,N_437);
and U1342 (N_1342,N_937,N_407);
nand U1343 (N_1343,N_777,N_397);
or U1344 (N_1344,N_837,N_658);
nand U1345 (N_1345,N_833,N_249);
nor U1346 (N_1346,N_459,N_263);
nor U1347 (N_1347,N_10,N_328);
nor U1348 (N_1348,N_381,N_713);
nand U1349 (N_1349,N_419,N_536);
or U1350 (N_1350,N_287,N_83);
and U1351 (N_1351,N_6,N_5);
nand U1352 (N_1352,N_434,N_795);
or U1353 (N_1353,N_973,N_436);
or U1354 (N_1354,N_27,N_252);
or U1355 (N_1355,N_382,N_635);
nand U1356 (N_1356,N_581,N_90);
and U1357 (N_1357,N_376,N_709);
or U1358 (N_1358,N_903,N_541);
or U1359 (N_1359,N_938,N_779);
and U1360 (N_1360,N_960,N_151);
xor U1361 (N_1361,N_410,N_136);
nor U1362 (N_1362,N_453,N_691);
and U1363 (N_1363,N_137,N_52);
nor U1364 (N_1364,N_617,N_883);
nor U1365 (N_1365,N_927,N_547);
or U1366 (N_1366,N_924,N_274);
or U1367 (N_1367,N_719,N_313);
and U1368 (N_1368,N_293,N_514);
or U1369 (N_1369,N_13,N_760);
or U1370 (N_1370,N_425,N_389);
nor U1371 (N_1371,N_202,N_834);
nand U1372 (N_1372,N_868,N_763);
or U1373 (N_1373,N_105,N_939);
nand U1374 (N_1374,N_542,N_29);
nand U1375 (N_1375,N_109,N_820);
nand U1376 (N_1376,N_625,N_934);
nor U1377 (N_1377,N_836,N_41);
nand U1378 (N_1378,N_687,N_999);
and U1379 (N_1379,N_522,N_730);
nor U1380 (N_1380,N_895,N_191);
nor U1381 (N_1381,N_607,N_372);
nor U1382 (N_1382,N_527,N_80);
and U1383 (N_1383,N_782,N_848);
nor U1384 (N_1384,N_612,N_745);
or U1385 (N_1385,N_769,N_190);
nor U1386 (N_1386,N_586,N_762);
nor U1387 (N_1387,N_130,N_165);
and U1388 (N_1388,N_449,N_45);
and U1389 (N_1389,N_509,N_404);
nand U1390 (N_1390,N_119,N_916);
nor U1391 (N_1391,N_169,N_986);
nand U1392 (N_1392,N_60,N_611);
or U1393 (N_1393,N_340,N_989);
nand U1394 (N_1394,N_148,N_907);
nand U1395 (N_1395,N_869,N_537);
or U1396 (N_1396,N_182,N_501);
or U1397 (N_1397,N_523,N_326);
and U1398 (N_1398,N_87,N_307);
or U1399 (N_1399,N_254,N_53);
or U1400 (N_1400,N_918,N_31);
and U1401 (N_1401,N_791,N_520);
or U1402 (N_1402,N_452,N_129);
nand U1403 (N_1403,N_935,N_51);
nand U1404 (N_1404,N_70,N_401);
and U1405 (N_1405,N_194,N_385);
and U1406 (N_1406,N_775,N_715);
nand U1407 (N_1407,N_341,N_261);
nor U1408 (N_1408,N_461,N_357);
or U1409 (N_1409,N_632,N_915);
nand U1410 (N_1410,N_234,N_697);
nor U1411 (N_1411,N_227,N_835);
xnor U1412 (N_1412,N_23,N_701);
or U1413 (N_1413,N_928,N_516);
nand U1414 (N_1414,N_113,N_988);
or U1415 (N_1415,N_909,N_308);
and U1416 (N_1416,N_14,N_208);
and U1417 (N_1417,N_688,N_88);
nand U1418 (N_1418,N_538,N_913);
or U1419 (N_1419,N_776,N_26);
nor U1420 (N_1420,N_546,N_242);
xor U1421 (N_1421,N_548,N_800);
and U1422 (N_1422,N_269,N_936);
nor U1423 (N_1423,N_331,N_577);
nor U1424 (N_1424,N_81,N_152);
and U1425 (N_1425,N_360,N_819);
nor U1426 (N_1426,N_533,N_626);
and U1427 (N_1427,N_753,N_904);
nand U1428 (N_1428,N_677,N_412);
nand U1429 (N_1429,N_47,N_299);
or U1430 (N_1430,N_370,N_448);
and U1431 (N_1431,N_974,N_980);
and U1432 (N_1432,N_623,N_700);
and U1433 (N_1433,N_345,N_162);
nor U1434 (N_1434,N_544,N_553);
and U1435 (N_1435,N_831,N_978);
and U1436 (N_1436,N_943,N_484);
nor U1437 (N_1437,N_392,N_576);
and U1438 (N_1438,N_531,N_329);
and U1439 (N_1439,N_487,N_621);
and U1440 (N_1440,N_840,N_665);
or U1441 (N_1441,N_94,N_702);
nand U1442 (N_1442,N_705,N_100);
xor U1443 (N_1443,N_979,N_245);
and U1444 (N_1444,N_778,N_921);
nand U1445 (N_1445,N_991,N_585);
or U1446 (N_1446,N_253,N_256);
nor U1447 (N_1447,N_225,N_473);
nand U1448 (N_1448,N_752,N_154);
and U1449 (N_1449,N_802,N_241);
nor U1450 (N_1450,N_767,N_423);
or U1451 (N_1451,N_260,N_720);
nor U1452 (N_1452,N_584,N_880);
and U1453 (N_1453,N_258,N_910);
nor U1454 (N_1454,N_532,N_471);
nor U1455 (N_1455,N_458,N_798);
and U1456 (N_1456,N_48,N_440);
or U1457 (N_1457,N_82,N_792);
or U1458 (N_1458,N_4,N_141);
nand U1459 (N_1459,N_230,N_435);
nand U1460 (N_1460,N_549,N_217);
or U1461 (N_1461,N_275,N_344);
nor U1462 (N_1462,N_683,N_497);
nand U1463 (N_1463,N_929,N_291);
nand U1464 (N_1464,N_660,N_366);
and U1465 (N_1465,N_395,N_97);
nand U1466 (N_1466,N_15,N_469);
and U1467 (N_1467,N_157,N_378);
or U1468 (N_1468,N_456,N_605);
or U1469 (N_1469,N_588,N_118);
or U1470 (N_1470,N_596,N_430);
or U1471 (N_1471,N_856,N_639);
and U1472 (N_1472,N_220,N_355);
or U1473 (N_1473,N_265,N_405);
and U1474 (N_1474,N_990,N_203);
or U1475 (N_1475,N_866,N_569);
nor U1476 (N_1476,N_11,N_16);
nand U1477 (N_1477,N_981,N_729);
nand U1478 (N_1478,N_17,N_853);
nor U1479 (N_1479,N_408,N_79);
or U1480 (N_1480,N_650,N_361);
nand U1481 (N_1481,N_363,N_567);
nand U1482 (N_1482,N_673,N_885);
or U1483 (N_1483,N_442,N_282);
nor U1484 (N_1484,N_61,N_959);
nor U1485 (N_1485,N_262,N_890);
nor U1486 (N_1486,N_852,N_594);
nand U1487 (N_1487,N_969,N_34);
or U1488 (N_1488,N_470,N_44);
nor U1489 (N_1489,N_815,N_39);
nor U1490 (N_1490,N_142,N_323);
or U1491 (N_1491,N_166,N_636);
xor U1492 (N_1492,N_529,N_551);
nand U1493 (N_1493,N_764,N_813);
nor U1494 (N_1494,N_877,N_738);
nand U1495 (N_1495,N_731,N_295);
and U1496 (N_1496,N_186,N_158);
nand U1497 (N_1497,N_213,N_808);
xnor U1498 (N_1498,N_424,N_616);
or U1499 (N_1499,N_377,N_765);
and U1500 (N_1500,N_911,N_711);
or U1501 (N_1501,N_892,N_827);
nor U1502 (N_1502,N_83,N_166);
nand U1503 (N_1503,N_280,N_349);
xor U1504 (N_1504,N_839,N_17);
and U1505 (N_1505,N_485,N_21);
nor U1506 (N_1506,N_620,N_724);
and U1507 (N_1507,N_96,N_175);
nor U1508 (N_1508,N_97,N_467);
nor U1509 (N_1509,N_402,N_401);
nand U1510 (N_1510,N_846,N_714);
or U1511 (N_1511,N_303,N_494);
xnor U1512 (N_1512,N_580,N_257);
nor U1513 (N_1513,N_133,N_181);
nand U1514 (N_1514,N_287,N_331);
or U1515 (N_1515,N_661,N_954);
and U1516 (N_1516,N_345,N_988);
nor U1517 (N_1517,N_360,N_880);
or U1518 (N_1518,N_296,N_845);
and U1519 (N_1519,N_402,N_930);
nand U1520 (N_1520,N_577,N_138);
nand U1521 (N_1521,N_64,N_761);
and U1522 (N_1522,N_815,N_271);
or U1523 (N_1523,N_30,N_513);
and U1524 (N_1524,N_950,N_158);
or U1525 (N_1525,N_138,N_285);
nor U1526 (N_1526,N_390,N_89);
or U1527 (N_1527,N_752,N_821);
nand U1528 (N_1528,N_492,N_901);
or U1529 (N_1529,N_690,N_510);
or U1530 (N_1530,N_986,N_655);
and U1531 (N_1531,N_615,N_191);
nor U1532 (N_1532,N_864,N_784);
and U1533 (N_1533,N_767,N_561);
or U1534 (N_1534,N_452,N_300);
nor U1535 (N_1535,N_195,N_883);
nand U1536 (N_1536,N_633,N_848);
and U1537 (N_1537,N_935,N_385);
or U1538 (N_1538,N_63,N_302);
nand U1539 (N_1539,N_703,N_124);
nand U1540 (N_1540,N_143,N_449);
or U1541 (N_1541,N_938,N_962);
or U1542 (N_1542,N_51,N_212);
or U1543 (N_1543,N_401,N_994);
nand U1544 (N_1544,N_368,N_762);
and U1545 (N_1545,N_530,N_451);
nor U1546 (N_1546,N_769,N_690);
or U1547 (N_1547,N_700,N_615);
nor U1548 (N_1548,N_299,N_686);
or U1549 (N_1549,N_443,N_648);
nand U1550 (N_1550,N_406,N_285);
or U1551 (N_1551,N_600,N_565);
nor U1552 (N_1552,N_480,N_950);
nand U1553 (N_1553,N_866,N_49);
or U1554 (N_1554,N_640,N_229);
and U1555 (N_1555,N_402,N_139);
nand U1556 (N_1556,N_118,N_459);
nor U1557 (N_1557,N_708,N_480);
nor U1558 (N_1558,N_25,N_564);
or U1559 (N_1559,N_529,N_526);
nor U1560 (N_1560,N_590,N_304);
or U1561 (N_1561,N_850,N_825);
nor U1562 (N_1562,N_670,N_749);
and U1563 (N_1563,N_178,N_713);
nand U1564 (N_1564,N_53,N_421);
nor U1565 (N_1565,N_761,N_367);
nand U1566 (N_1566,N_580,N_885);
nand U1567 (N_1567,N_444,N_871);
nand U1568 (N_1568,N_156,N_203);
nor U1569 (N_1569,N_856,N_663);
nor U1570 (N_1570,N_829,N_949);
nor U1571 (N_1571,N_480,N_353);
or U1572 (N_1572,N_516,N_868);
or U1573 (N_1573,N_752,N_502);
nor U1574 (N_1574,N_354,N_503);
nand U1575 (N_1575,N_941,N_121);
nor U1576 (N_1576,N_426,N_147);
nand U1577 (N_1577,N_989,N_21);
nor U1578 (N_1578,N_967,N_352);
and U1579 (N_1579,N_963,N_217);
nand U1580 (N_1580,N_751,N_901);
or U1581 (N_1581,N_214,N_402);
nor U1582 (N_1582,N_94,N_592);
nor U1583 (N_1583,N_243,N_135);
nor U1584 (N_1584,N_348,N_237);
nor U1585 (N_1585,N_366,N_913);
or U1586 (N_1586,N_548,N_603);
nor U1587 (N_1587,N_852,N_118);
nand U1588 (N_1588,N_294,N_926);
or U1589 (N_1589,N_440,N_403);
nand U1590 (N_1590,N_562,N_424);
nand U1591 (N_1591,N_523,N_330);
nand U1592 (N_1592,N_926,N_464);
nand U1593 (N_1593,N_104,N_556);
or U1594 (N_1594,N_118,N_259);
nor U1595 (N_1595,N_642,N_736);
nor U1596 (N_1596,N_360,N_233);
and U1597 (N_1597,N_727,N_340);
nor U1598 (N_1598,N_504,N_313);
nand U1599 (N_1599,N_930,N_621);
or U1600 (N_1600,N_414,N_120);
nand U1601 (N_1601,N_540,N_116);
or U1602 (N_1602,N_76,N_111);
and U1603 (N_1603,N_506,N_413);
or U1604 (N_1604,N_407,N_434);
nand U1605 (N_1605,N_353,N_71);
nor U1606 (N_1606,N_801,N_735);
nor U1607 (N_1607,N_315,N_468);
or U1608 (N_1608,N_898,N_272);
or U1609 (N_1609,N_248,N_476);
nor U1610 (N_1610,N_268,N_372);
and U1611 (N_1611,N_263,N_525);
nand U1612 (N_1612,N_936,N_864);
nand U1613 (N_1613,N_881,N_639);
or U1614 (N_1614,N_476,N_737);
nor U1615 (N_1615,N_325,N_559);
nor U1616 (N_1616,N_270,N_634);
nor U1617 (N_1617,N_16,N_473);
or U1618 (N_1618,N_931,N_43);
and U1619 (N_1619,N_19,N_851);
nor U1620 (N_1620,N_602,N_433);
or U1621 (N_1621,N_281,N_277);
and U1622 (N_1622,N_144,N_304);
nor U1623 (N_1623,N_261,N_579);
nor U1624 (N_1624,N_498,N_388);
or U1625 (N_1625,N_511,N_871);
or U1626 (N_1626,N_832,N_184);
xor U1627 (N_1627,N_251,N_221);
nand U1628 (N_1628,N_371,N_466);
and U1629 (N_1629,N_420,N_526);
nand U1630 (N_1630,N_662,N_372);
nand U1631 (N_1631,N_416,N_751);
nor U1632 (N_1632,N_111,N_538);
or U1633 (N_1633,N_472,N_73);
or U1634 (N_1634,N_722,N_884);
or U1635 (N_1635,N_955,N_294);
or U1636 (N_1636,N_563,N_125);
or U1637 (N_1637,N_69,N_100);
nor U1638 (N_1638,N_664,N_238);
nor U1639 (N_1639,N_555,N_331);
nor U1640 (N_1640,N_114,N_388);
and U1641 (N_1641,N_712,N_899);
or U1642 (N_1642,N_810,N_812);
nand U1643 (N_1643,N_526,N_103);
nand U1644 (N_1644,N_18,N_851);
and U1645 (N_1645,N_153,N_63);
nor U1646 (N_1646,N_306,N_265);
and U1647 (N_1647,N_347,N_187);
nand U1648 (N_1648,N_112,N_764);
nand U1649 (N_1649,N_142,N_527);
nand U1650 (N_1650,N_230,N_322);
and U1651 (N_1651,N_535,N_582);
nor U1652 (N_1652,N_183,N_905);
and U1653 (N_1653,N_711,N_190);
or U1654 (N_1654,N_42,N_299);
or U1655 (N_1655,N_897,N_307);
xnor U1656 (N_1656,N_67,N_621);
nand U1657 (N_1657,N_264,N_963);
nand U1658 (N_1658,N_469,N_413);
nand U1659 (N_1659,N_169,N_829);
nor U1660 (N_1660,N_815,N_407);
and U1661 (N_1661,N_475,N_173);
nor U1662 (N_1662,N_341,N_959);
nand U1663 (N_1663,N_875,N_45);
nand U1664 (N_1664,N_510,N_570);
or U1665 (N_1665,N_988,N_14);
or U1666 (N_1666,N_264,N_108);
xnor U1667 (N_1667,N_611,N_328);
or U1668 (N_1668,N_118,N_650);
and U1669 (N_1669,N_61,N_655);
and U1670 (N_1670,N_527,N_6);
nor U1671 (N_1671,N_959,N_387);
and U1672 (N_1672,N_360,N_854);
or U1673 (N_1673,N_926,N_541);
and U1674 (N_1674,N_442,N_150);
nor U1675 (N_1675,N_430,N_194);
and U1676 (N_1676,N_5,N_143);
or U1677 (N_1677,N_148,N_412);
or U1678 (N_1678,N_422,N_345);
nor U1679 (N_1679,N_59,N_169);
or U1680 (N_1680,N_11,N_471);
or U1681 (N_1681,N_691,N_247);
nand U1682 (N_1682,N_504,N_941);
and U1683 (N_1683,N_150,N_795);
and U1684 (N_1684,N_733,N_216);
or U1685 (N_1685,N_506,N_459);
or U1686 (N_1686,N_554,N_706);
nor U1687 (N_1687,N_956,N_355);
and U1688 (N_1688,N_852,N_718);
and U1689 (N_1689,N_256,N_830);
or U1690 (N_1690,N_836,N_481);
nand U1691 (N_1691,N_378,N_455);
nand U1692 (N_1692,N_963,N_670);
or U1693 (N_1693,N_263,N_95);
and U1694 (N_1694,N_720,N_671);
and U1695 (N_1695,N_33,N_250);
nor U1696 (N_1696,N_896,N_912);
and U1697 (N_1697,N_63,N_448);
or U1698 (N_1698,N_8,N_542);
nor U1699 (N_1699,N_931,N_810);
and U1700 (N_1700,N_858,N_335);
nor U1701 (N_1701,N_56,N_315);
and U1702 (N_1702,N_505,N_542);
or U1703 (N_1703,N_634,N_485);
nor U1704 (N_1704,N_27,N_655);
nor U1705 (N_1705,N_948,N_472);
nor U1706 (N_1706,N_225,N_769);
or U1707 (N_1707,N_392,N_545);
and U1708 (N_1708,N_804,N_954);
and U1709 (N_1709,N_806,N_285);
nand U1710 (N_1710,N_406,N_543);
or U1711 (N_1711,N_170,N_373);
nor U1712 (N_1712,N_775,N_860);
nand U1713 (N_1713,N_91,N_472);
nand U1714 (N_1714,N_678,N_494);
or U1715 (N_1715,N_473,N_319);
nor U1716 (N_1716,N_959,N_328);
or U1717 (N_1717,N_536,N_947);
nor U1718 (N_1718,N_175,N_590);
and U1719 (N_1719,N_134,N_656);
nor U1720 (N_1720,N_686,N_713);
nand U1721 (N_1721,N_889,N_856);
nand U1722 (N_1722,N_341,N_37);
nand U1723 (N_1723,N_188,N_213);
or U1724 (N_1724,N_517,N_913);
nor U1725 (N_1725,N_712,N_923);
or U1726 (N_1726,N_165,N_789);
and U1727 (N_1727,N_254,N_896);
nand U1728 (N_1728,N_341,N_597);
nand U1729 (N_1729,N_741,N_318);
nand U1730 (N_1730,N_739,N_108);
nor U1731 (N_1731,N_764,N_403);
and U1732 (N_1732,N_803,N_910);
nor U1733 (N_1733,N_251,N_732);
or U1734 (N_1734,N_45,N_760);
and U1735 (N_1735,N_397,N_781);
xor U1736 (N_1736,N_951,N_65);
or U1737 (N_1737,N_162,N_914);
nand U1738 (N_1738,N_686,N_402);
and U1739 (N_1739,N_571,N_608);
and U1740 (N_1740,N_894,N_223);
nor U1741 (N_1741,N_496,N_452);
nor U1742 (N_1742,N_498,N_422);
nor U1743 (N_1743,N_297,N_325);
nand U1744 (N_1744,N_611,N_541);
nand U1745 (N_1745,N_801,N_448);
xor U1746 (N_1746,N_26,N_904);
nor U1747 (N_1747,N_843,N_306);
nor U1748 (N_1748,N_588,N_138);
or U1749 (N_1749,N_248,N_60);
nand U1750 (N_1750,N_60,N_471);
nand U1751 (N_1751,N_227,N_93);
or U1752 (N_1752,N_523,N_700);
and U1753 (N_1753,N_677,N_142);
nor U1754 (N_1754,N_804,N_576);
nor U1755 (N_1755,N_150,N_258);
nand U1756 (N_1756,N_612,N_225);
nor U1757 (N_1757,N_849,N_571);
nor U1758 (N_1758,N_332,N_229);
nand U1759 (N_1759,N_517,N_728);
and U1760 (N_1760,N_923,N_413);
nor U1761 (N_1761,N_96,N_49);
or U1762 (N_1762,N_548,N_263);
and U1763 (N_1763,N_798,N_217);
nor U1764 (N_1764,N_994,N_729);
nor U1765 (N_1765,N_178,N_136);
xor U1766 (N_1766,N_304,N_176);
nor U1767 (N_1767,N_613,N_941);
or U1768 (N_1768,N_971,N_628);
nand U1769 (N_1769,N_79,N_560);
or U1770 (N_1770,N_269,N_253);
nand U1771 (N_1771,N_121,N_250);
nor U1772 (N_1772,N_415,N_756);
nand U1773 (N_1773,N_6,N_526);
and U1774 (N_1774,N_360,N_403);
and U1775 (N_1775,N_334,N_973);
or U1776 (N_1776,N_481,N_704);
or U1777 (N_1777,N_867,N_275);
and U1778 (N_1778,N_845,N_196);
nand U1779 (N_1779,N_570,N_61);
or U1780 (N_1780,N_255,N_867);
nor U1781 (N_1781,N_674,N_187);
or U1782 (N_1782,N_284,N_778);
xnor U1783 (N_1783,N_317,N_203);
and U1784 (N_1784,N_89,N_125);
nor U1785 (N_1785,N_143,N_667);
or U1786 (N_1786,N_802,N_254);
nor U1787 (N_1787,N_78,N_756);
nand U1788 (N_1788,N_587,N_985);
nand U1789 (N_1789,N_850,N_154);
or U1790 (N_1790,N_297,N_395);
and U1791 (N_1791,N_647,N_669);
nand U1792 (N_1792,N_392,N_750);
nand U1793 (N_1793,N_936,N_158);
nand U1794 (N_1794,N_345,N_536);
nand U1795 (N_1795,N_40,N_138);
xnor U1796 (N_1796,N_180,N_89);
or U1797 (N_1797,N_21,N_853);
or U1798 (N_1798,N_514,N_882);
nand U1799 (N_1799,N_15,N_22);
or U1800 (N_1800,N_205,N_207);
nor U1801 (N_1801,N_167,N_54);
nor U1802 (N_1802,N_694,N_119);
nor U1803 (N_1803,N_536,N_858);
or U1804 (N_1804,N_681,N_109);
nor U1805 (N_1805,N_738,N_490);
or U1806 (N_1806,N_795,N_765);
nor U1807 (N_1807,N_550,N_477);
xor U1808 (N_1808,N_538,N_685);
and U1809 (N_1809,N_787,N_250);
nor U1810 (N_1810,N_796,N_168);
nor U1811 (N_1811,N_990,N_842);
nand U1812 (N_1812,N_969,N_698);
or U1813 (N_1813,N_91,N_805);
nand U1814 (N_1814,N_209,N_552);
or U1815 (N_1815,N_130,N_461);
or U1816 (N_1816,N_376,N_364);
and U1817 (N_1817,N_222,N_505);
and U1818 (N_1818,N_35,N_854);
or U1819 (N_1819,N_940,N_143);
nand U1820 (N_1820,N_130,N_439);
nor U1821 (N_1821,N_132,N_494);
or U1822 (N_1822,N_968,N_573);
or U1823 (N_1823,N_547,N_47);
and U1824 (N_1824,N_675,N_318);
nor U1825 (N_1825,N_938,N_292);
nor U1826 (N_1826,N_189,N_711);
xor U1827 (N_1827,N_625,N_936);
nor U1828 (N_1828,N_59,N_901);
nor U1829 (N_1829,N_497,N_114);
or U1830 (N_1830,N_105,N_733);
and U1831 (N_1831,N_907,N_568);
nand U1832 (N_1832,N_984,N_422);
nand U1833 (N_1833,N_780,N_284);
nor U1834 (N_1834,N_963,N_989);
and U1835 (N_1835,N_680,N_82);
or U1836 (N_1836,N_783,N_742);
nor U1837 (N_1837,N_427,N_520);
nand U1838 (N_1838,N_821,N_936);
and U1839 (N_1839,N_30,N_149);
nand U1840 (N_1840,N_771,N_444);
and U1841 (N_1841,N_458,N_107);
and U1842 (N_1842,N_912,N_947);
and U1843 (N_1843,N_835,N_950);
nand U1844 (N_1844,N_520,N_392);
and U1845 (N_1845,N_262,N_817);
and U1846 (N_1846,N_977,N_308);
nand U1847 (N_1847,N_379,N_796);
and U1848 (N_1848,N_440,N_803);
and U1849 (N_1849,N_994,N_687);
nor U1850 (N_1850,N_973,N_484);
nand U1851 (N_1851,N_875,N_689);
and U1852 (N_1852,N_985,N_677);
nand U1853 (N_1853,N_176,N_655);
nor U1854 (N_1854,N_868,N_845);
or U1855 (N_1855,N_210,N_729);
nor U1856 (N_1856,N_75,N_680);
and U1857 (N_1857,N_50,N_544);
and U1858 (N_1858,N_915,N_385);
and U1859 (N_1859,N_144,N_132);
or U1860 (N_1860,N_89,N_79);
or U1861 (N_1861,N_251,N_708);
nor U1862 (N_1862,N_780,N_86);
nand U1863 (N_1863,N_389,N_416);
nor U1864 (N_1864,N_737,N_291);
or U1865 (N_1865,N_254,N_591);
and U1866 (N_1866,N_821,N_759);
or U1867 (N_1867,N_702,N_584);
nand U1868 (N_1868,N_513,N_23);
nand U1869 (N_1869,N_523,N_755);
nand U1870 (N_1870,N_141,N_424);
and U1871 (N_1871,N_231,N_801);
nor U1872 (N_1872,N_467,N_543);
nand U1873 (N_1873,N_251,N_152);
nor U1874 (N_1874,N_726,N_376);
or U1875 (N_1875,N_127,N_582);
or U1876 (N_1876,N_469,N_945);
nor U1877 (N_1877,N_801,N_238);
and U1878 (N_1878,N_716,N_538);
and U1879 (N_1879,N_124,N_705);
nand U1880 (N_1880,N_907,N_304);
and U1881 (N_1881,N_292,N_421);
nor U1882 (N_1882,N_191,N_516);
nor U1883 (N_1883,N_804,N_778);
nor U1884 (N_1884,N_941,N_41);
or U1885 (N_1885,N_941,N_823);
nand U1886 (N_1886,N_918,N_892);
and U1887 (N_1887,N_664,N_881);
or U1888 (N_1888,N_107,N_725);
nand U1889 (N_1889,N_742,N_250);
xor U1890 (N_1890,N_709,N_28);
nor U1891 (N_1891,N_534,N_168);
or U1892 (N_1892,N_650,N_928);
and U1893 (N_1893,N_290,N_76);
and U1894 (N_1894,N_381,N_841);
or U1895 (N_1895,N_763,N_747);
and U1896 (N_1896,N_720,N_972);
and U1897 (N_1897,N_386,N_899);
or U1898 (N_1898,N_329,N_1);
and U1899 (N_1899,N_945,N_626);
and U1900 (N_1900,N_410,N_285);
nor U1901 (N_1901,N_978,N_554);
nand U1902 (N_1902,N_200,N_599);
nand U1903 (N_1903,N_315,N_981);
and U1904 (N_1904,N_202,N_29);
nor U1905 (N_1905,N_177,N_443);
and U1906 (N_1906,N_621,N_280);
or U1907 (N_1907,N_870,N_701);
or U1908 (N_1908,N_907,N_629);
or U1909 (N_1909,N_892,N_920);
nand U1910 (N_1910,N_976,N_130);
and U1911 (N_1911,N_940,N_637);
and U1912 (N_1912,N_614,N_815);
nor U1913 (N_1913,N_494,N_574);
nand U1914 (N_1914,N_733,N_583);
nand U1915 (N_1915,N_643,N_865);
nor U1916 (N_1916,N_855,N_109);
or U1917 (N_1917,N_975,N_19);
and U1918 (N_1918,N_632,N_124);
xor U1919 (N_1919,N_955,N_492);
nand U1920 (N_1920,N_65,N_889);
nor U1921 (N_1921,N_877,N_198);
and U1922 (N_1922,N_676,N_268);
nand U1923 (N_1923,N_782,N_45);
or U1924 (N_1924,N_888,N_269);
or U1925 (N_1925,N_620,N_745);
or U1926 (N_1926,N_892,N_598);
or U1927 (N_1927,N_227,N_641);
nor U1928 (N_1928,N_41,N_360);
or U1929 (N_1929,N_960,N_170);
or U1930 (N_1930,N_150,N_645);
and U1931 (N_1931,N_220,N_772);
and U1932 (N_1932,N_551,N_539);
nor U1933 (N_1933,N_602,N_65);
and U1934 (N_1934,N_500,N_795);
nand U1935 (N_1935,N_677,N_981);
nand U1936 (N_1936,N_117,N_939);
nand U1937 (N_1937,N_545,N_22);
nand U1938 (N_1938,N_385,N_963);
or U1939 (N_1939,N_159,N_751);
nor U1940 (N_1940,N_228,N_628);
and U1941 (N_1941,N_699,N_961);
nand U1942 (N_1942,N_488,N_782);
or U1943 (N_1943,N_915,N_857);
or U1944 (N_1944,N_287,N_829);
or U1945 (N_1945,N_318,N_128);
and U1946 (N_1946,N_414,N_639);
xnor U1947 (N_1947,N_156,N_954);
nand U1948 (N_1948,N_380,N_137);
or U1949 (N_1949,N_795,N_61);
and U1950 (N_1950,N_951,N_11);
nand U1951 (N_1951,N_538,N_546);
nor U1952 (N_1952,N_724,N_342);
nor U1953 (N_1953,N_298,N_639);
or U1954 (N_1954,N_691,N_781);
or U1955 (N_1955,N_659,N_461);
nor U1956 (N_1956,N_297,N_65);
and U1957 (N_1957,N_77,N_510);
or U1958 (N_1958,N_519,N_631);
nor U1959 (N_1959,N_877,N_977);
nand U1960 (N_1960,N_768,N_253);
or U1961 (N_1961,N_562,N_39);
or U1962 (N_1962,N_718,N_631);
nand U1963 (N_1963,N_143,N_862);
nand U1964 (N_1964,N_41,N_548);
and U1965 (N_1965,N_940,N_278);
or U1966 (N_1966,N_797,N_73);
nand U1967 (N_1967,N_228,N_752);
nand U1968 (N_1968,N_235,N_223);
nand U1969 (N_1969,N_837,N_327);
nor U1970 (N_1970,N_937,N_221);
nor U1971 (N_1971,N_563,N_901);
and U1972 (N_1972,N_83,N_343);
nand U1973 (N_1973,N_779,N_802);
or U1974 (N_1974,N_635,N_782);
nand U1975 (N_1975,N_113,N_136);
nand U1976 (N_1976,N_774,N_862);
or U1977 (N_1977,N_944,N_772);
or U1978 (N_1978,N_528,N_575);
and U1979 (N_1979,N_998,N_523);
nor U1980 (N_1980,N_754,N_673);
nand U1981 (N_1981,N_611,N_313);
nand U1982 (N_1982,N_18,N_289);
nand U1983 (N_1983,N_817,N_467);
or U1984 (N_1984,N_81,N_50);
or U1985 (N_1985,N_442,N_925);
and U1986 (N_1986,N_150,N_696);
nand U1987 (N_1987,N_703,N_134);
and U1988 (N_1988,N_834,N_15);
nor U1989 (N_1989,N_890,N_350);
nand U1990 (N_1990,N_571,N_407);
and U1991 (N_1991,N_354,N_606);
or U1992 (N_1992,N_87,N_929);
nand U1993 (N_1993,N_768,N_851);
nor U1994 (N_1994,N_115,N_988);
nand U1995 (N_1995,N_833,N_591);
nor U1996 (N_1996,N_483,N_32);
and U1997 (N_1997,N_698,N_60);
nand U1998 (N_1998,N_933,N_439);
and U1999 (N_1999,N_612,N_420);
nor U2000 (N_2000,N_1604,N_1470);
nor U2001 (N_2001,N_1519,N_1273);
nor U2002 (N_2002,N_1988,N_1298);
nand U2003 (N_2003,N_1414,N_1576);
or U2004 (N_2004,N_1429,N_1067);
nand U2005 (N_2005,N_1627,N_1566);
or U2006 (N_2006,N_1233,N_1420);
nand U2007 (N_2007,N_1662,N_1919);
and U2008 (N_2008,N_1467,N_1186);
or U2009 (N_2009,N_1318,N_1504);
nor U2010 (N_2010,N_1471,N_1001);
and U2011 (N_2011,N_1833,N_1144);
or U2012 (N_2012,N_1054,N_1909);
and U2013 (N_2013,N_1128,N_1527);
or U2014 (N_2014,N_1291,N_1741);
nor U2015 (N_2015,N_1478,N_1285);
and U2016 (N_2016,N_1661,N_1161);
or U2017 (N_2017,N_1375,N_1350);
or U2018 (N_2018,N_1212,N_1850);
nand U2019 (N_2019,N_1931,N_1480);
or U2020 (N_2020,N_1776,N_1404);
or U2021 (N_2021,N_1500,N_1312);
and U2022 (N_2022,N_1171,N_1968);
nand U2023 (N_2023,N_1792,N_1704);
nand U2024 (N_2024,N_1226,N_1538);
or U2025 (N_2025,N_1256,N_1544);
nor U2026 (N_2026,N_1996,N_1723);
and U2027 (N_2027,N_1717,N_1410);
and U2028 (N_2028,N_1698,N_1006);
nand U2029 (N_2029,N_1643,N_1346);
nor U2030 (N_2030,N_1829,N_1022);
or U2031 (N_2031,N_1738,N_1481);
nand U2032 (N_2032,N_1063,N_1516);
nor U2033 (N_2033,N_1613,N_1959);
nor U2034 (N_2034,N_1526,N_1210);
nand U2035 (N_2035,N_1622,N_1250);
or U2036 (N_2036,N_1170,N_1834);
nand U2037 (N_2037,N_1916,N_1589);
nand U2038 (N_2038,N_1729,N_1407);
or U2039 (N_2039,N_1579,N_1882);
nand U2040 (N_2040,N_1458,N_1353);
nor U2041 (N_2041,N_1240,N_1672);
and U2042 (N_2042,N_1191,N_1711);
and U2043 (N_2043,N_1534,N_1096);
and U2044 (N_2044,N_1880,N_1267);
nor U2045 (N_2045,N_1227,N_1413);
nand U2046 (N_2046,N_1202,N_1980);
and U2047 (N_2047,N_1888,N_1749);
nand U2048 (N_2048,N_1449,N_1397);
nor U2049 (N_2049,N_1941,N_1724);
nor U2050 (N_2050,N_1015,N_1178);
and U2051 (N_2051,N_1571,N_1190);
or U2052 (N_2052,N_1563,N_1127);
nand U2053 (N_2053,N_1716,N_1751);
or U2054 (N_2054,N_1945,N_1646);
nand U2055 (N_2055,N_1088,N_1371);
nand U2056 (N_2056,N_1879,N_1506);
and U2057 (N_2057,N_1477,N_1638);
and U2058 (N_2058,N_1623,N_1344);
and U2059 (N_2059,N_1352,N_1854);
or U2060 (N_2060,N_1886,N_1020);
and U2061 (N_2061,N_1985,N_1466);
nand U2062 (N_2062,N_1666,N_1875);
nor U2063 (N_2063,N_1992,N_1361);
xor U2064 (N_2064,N_1671,N_1997);
nor U2065 (N_2065,N_1869,N_1765);
or U2066 (N_2066,N_1330,N_1338);
nand U2067 (N_2067,N_1373,N_1194);
nand U2068 (N_2068,N_1857,N_1129);
nand U2069 (N_2069,N_1933,N_1101);
xnor U2070 (N_2070,N_1138,N_1117);
or U2071 (N_2071,N_1952,N_1114);
nor U2072 (N_2072,N_1475,N_1680);
nor U2073 (N_2073,N_1356,N_1209);
nand U2074 (N_2074,N_1616,N_1349);
nor U2075 (N_2075,N_1657,N_1351);
nand U2076 (N_2076,N_1795,N_1339);
and U2077 (N_2077,N_1777,N_1440);
and U2078 (N_2078,N_1963,N_1447);
or U2079 (N_2079,N_1621,N_1663);
and U2080 (N_2080,N_1051,N_1214);
and U2081 (N_2081,N_1340,N_1756);
or U2082 (N_2082,N_1183,N_1456);
and U2083 (N_2083,N_1310,N_1848);
or U2084 (N_2084,N_1759,N_1454);
nand U2085 (N_2085,N_1327,N_1642);
or U2086 (N_2086,N_1625,N_1337);
nor U2087 (N_2087,N_1774,N_1826);
or U2088 (N_2088,N_1247,N_1173);
or U2089 (N_2089,N_1799,N_1253);
or U2090 (N_2090,N_1292,N_1842);
xor U2091 (N_2091,N_1103,N_1064);
nand U2092 (N_2092,N_1261,N_1592);
and U2093 (N_2093,N_1084,N_1168);
and U2094 (N_2094,N_1803,N_1892);
nand U2095 (N_2095,N_1607,N_1690);
nand U2096 (N_2096,N_1860,N_1374);
or U2097 (N_2097,N_1787,N_1090);
nand U2098 (N_2098,N_1043,N_1815);
and U2099 (N_2099,N_1201,N_1231);
nand U2100 (N_2100,N_1999,N_1583);
or U2101 (N_2101,N_1841,N_1881);
and U2102 (N_2102,N_1007,N_1619);
or U2103 (N_2103,N_1132,N_1602);
nand U2104 (N_2104,N_1739,N_1900);
xor U2105 (N_2105,N_1555,N_1794);
nand U2106 (N_2106,N_1781,N_1174);
nand U2107 (N_2107,N_1782,N_1328);
nor U2108 (N_2108,N_1029,N_1198);
or U2109 (N_2109,N_1089,N_1958);
or U2110 (N_2110,N_1610,N_1034);
nand U2111 (N_2111,N_1159,N_1038);
or U2112 (N_2112,N_1217,N_1725);
nor U2113 (N_2113,N_1530,N_1542);
and U2114 (N_2114,N_1259,N_1493);
nand U2115 (N_2115,N_1216,N_1193);
nor U2116 (N_2116,N_1649,N_1917);
or U2117 (N_2117,N_1389,N_1620);
nand U2118 (N_2118,N_1164,N_1744);
nand U2119 (N_2119,N_1736,N_1584);
and U2120 (N_2120,N_1961,N_1957);
or U2121 (N_2121,N_1052,N_1167);
nor U2122 (N_2122,N_1942,N_1760);
or U2123 (N_2123,N_1733,N_1807);
nor U2124 (N_2124,N_1861,N_1699);
nand U2125 (N_2125,N_1363,N_1130);
nand U2126 (N_2126,N_1232,N_1686);
and U2127 (N_2127,N_1747,N_1087);
or U2128 (N_2128,N_1396,N_1681);
nor U2129 (N_2129,N_1510,N_1796);
or U2130 (N_2130,N_1425,N_1545);
and U2131 (N_2131,N_1966,N_1742);
nand U2132 (N_2132,N_1061,N_1573);
nor U2133 (N_2133,N_1936,N_1111);
nand U2134 (N_2134,N_1487,N_1234);
nor U2135 (N_2135,N_1362,N_1484);
nor U2136 (N_2136,N_1368,N_1609);
nor U2137 (N_2137,N_1712,N_1639);
and U2138 (N_2138,N_1115,N_1982);
or U2139 (N_2139,N_1734,N_1012);
or U2140 (N_2140,N_1406,N_1827);
and U2141 (N_2141,N_1182,N_1463);
nor U2142 (N_2142,N_1731,N_1549);
or U2143 (N_2143,N_1011,N_1417);
nor U2144 (N_2144,N_1947,N_1370);
or U2145 (N_2145,N_1077,N_1165);
or U2146 (N_2146,N_1612,N_1753);
and U2147 (N_2147,N_1636,N_1002);
or U2148 (N_2148,N_1846,N_1319);
or U2149 (N_2149,N_1770,N_1539);
or U2150 (N_2150,N_1066,N_1994);
xor U2151 (N_2151,N_1778,N_1257);
or U2152 (N_2152,N_1313,N_1907);
nor U2153 (N_2153,N_1930,N_1412);
or U2154 (N_2154,N_1387,N_1058);
nor U2155 (N_2155,N_1239,N_1172);
nand U2156 (N_2156,N_1145,N_1940);
nand U2157 (N_2157,N_1856,N_1032);
or U2158 (N_2158,N_1868,N_1904);
and U2159 (N_2159,N_1503,N_1154);
and U2160 (N_2160,N_1139,N_1902);
or U2161 (N_2161,N_1564,N_1019);
nand U2162 (N_2162,N_1594,N_1677);
nand U2163 (N_2163,N_1099,N_1901);
and U2164 (N_2164,N_1093,N_1042);
nand U2165 (N_2165,N_1659,N_1687);
nor U2166 (N_2166,N_1301,N_1847);
and U2167 (N_2167,N_1763,N_1109);
or U2168 (N_2168,N_1498,N_1431);
or U2169 (N_2169,N_1142,N_1939);
and U2170 (N_2170,N_1702,N_1785);
and U2171 (N_2171,N_1320,N_1102);
nor U2172 (N_2172,N_1433,N_1331);
xnor U2173 (N_2173,N_1085,N_1804);
and U2174 (N_2174,N_1160,N_1325);
nand U2175 (N_2175,N_1153,N_1295);
and U2176 (N_2176,N_1461,N_1508);
or U2177 (N_2177,N_1673,N_1068);
or U2178 (N_2178,N_1211,N_1030);
or U2179 (N_2179,N_1131,N_1887);
nor U2180 (N_2180,N_1280,N_1260);
nand U2181 (N_2181,N_1568,N_1188);
nor U2182 (N_2182,N_1853,N_1514);
nand U2183 (N_2183,N_1578,N_1443);
and U2184 (N_2184,N_1469,N_1494);
or U2185 (N_2185,N_1163,N_1380);
and U2186 (N_2186,N_1924,N_1522);
nor U2187 (N_2187,N_1143,N_1392);
nor U2188 (N_2188,N_1755,N_1059);
and U2189 (N_2189,N_1665,N_1617);
and U2190 (N_2190,N_1121,N_1599);
nor U2191 (N_2191,N_1511,N_1452);
and U2192 (N_2192,N_1284,N_1246);
and U2193 (N_2193,N_1288,N_1849);
nand U2194 (N_2194,N_1376,N_1898);
and U2195 (N_2195,N_1048,N_1937);
nand U2196 (N_2196,N_1053,N_1683);
or U2197 (N_2197,N_1297,N_1046);
nor U2198 (N_2198,N_1772,N_1335);
nor U2199 (N_2199,N_1409,N_1306);
nand U2200 (N_2200,N_1446,N_1473);
and U2201 (N_2201,N_1014,N_1618);
or U2202 (N_2202,N_1520,N_1243);
nor U2203 (N_2203,N_1460,N_1601);
or U2204 (N_2204,N_1228,N_1737);
nor U2205 (N_2205,N_1040,N_1377);
or U2206 (N_2206,N_1070,N_1788);
and U2207 (N_2207,N_1444,N_1844);
nand U2208 (N_2208,N_1722,N_1141);
or U2209 (N_2209,N_1039,N_1714);
or U2210 (N_2210,N_1836,N_1864);
and U2211 (N_2211,N_1445,N_1329);
or U2212 (N_2212,N_1707,N_1010);
and U2213 (N_2213,N_1912,N_1586);
or U2214 (N_2214,N_1653,N_1728);
nand U2215 (N_2215,N_1667,N_1858);
nor U2216 (N_2216,N_1437,N_1220);
or U2217 (N_2217,N_1092,N_1264);
nor U2218 (N_2218,N_1422,N_1177);
or U2219 (N_2219,N_1700,N_1378);
nor U2220 (N_2220,N_1175,N_1013);
nand U2221 (N_2221,N_1105,N_1497);
and U2222 (N_2222,N_1802,N_1633);
or U2223 (N_2223,N_1730,N_1235);
nor U2224 (N_2224,N_1496,N_1541);
nand U2225 (N_2225,N_1743,N_1266);
and U2226 (N_2226,N_1254,N_1658);
or U2227 (N_2227,N_1786,N_1838);
xor U2228 (N_2228,N_1839,N_1840);
or U2229 (N_2229,N_1276,N_1364);
and U2230 (N_2230,N_1614,N_1877);
nor U2231 (N_2231,N_1465,N_1567);
nand U2232 (N_2232,N_1675,N_1157);
nor U2233 (N_2233,N_1322,N_1720);
or U2234 (N_2234,N_1082,N_1630);
nor U2235 (N_2235,N_1453,N_1867);
nor U2236 (N_2236,N_1537,N_1421);
or U2237 (N_2237,N_1348,N_1134);
and U2238 (N_2238,N_1265,N_1221);
nand U2239 (N_2239,N_1748,N_1071);
xnor U2240 (N_2240,N_1812,N_1791);
nand U2241 (N_2241,N_1780,N_1935);
nor U2242 (N_2242,N_1072,N_1296);
or U2243 (N_2243,N_1889,N_1208);
and U2244 (N_2244,N_1060,N_1492);
and U2245 (N_2245,N_1382,N_1823);
or U2246 (N_2246,N_1403,N_1789);
and U2247 (N_2247,N_1495,N_1577);
nand U2248 (N_2248,N_1028,N_1097);
nor U2249 (N_2249,N_1166,N_1689);
and U2250 (N_2250,N_1811,N_1464);
or U2251 (N_2251,N_1977,N_1628);
nor U2252 (N_2252,N_1830,N_1271);
nor U2253 (N_2253,N_1908,N_1552);
and U2254 (N_2254,N_1224,N_1278);
nand U2255 (N_2255,N_1423,N_1424);
nor U2256 (N_2256,N_1418,N_1925);
nand U2257 (N_2257,N_1018,N_1485);
nand U2258 (N_2258,N_1411,N_1715);
or U2259 (N_2259,N_1241,N_1113);
nor U2260 (N_2260,N_1771,N_1706);
nand U2261 (N_2261,N_1336,N_1648);
and U2262 (N_2262,N_1557,N_1929);
nor U2263 (N_2263,N_1651,N_1334);
or U2264 (N_2264,N_1691,N_1049);
or U2265 (N_2265,N_1441,N_1047);
nand U2266 (N_2266,N_1797,N_1927);
or U2267 (N_2267,N_1218,N_1822);
and U2268 (N_2268,N_1179,N_1915);
and U2269 (N_2269,N_1953,N_1585);
or U2270 (N_2270,N_1593,N_1535);
or U2271 (N_2271,N_1197,N_1180);
nor U2272 (N_2272,N_1415,N_1251);
or U2273 (N_2273,N_1595,N_1033);
and U2274 (N_2274,N_1512,N_1355);
nor U2275 (N_2275,N_1554,N_1360);
and U2276 (N_2276,N_1975,N_1314);
nand U2277 (N_2277,N_1004,N_1125);
nor U2278 (N_2278,N_1727,N_1600);
and U2279 (N_2279,N_1200,N_1920);
xnor U2280 (N_2280,N_1533,N_1199);
nor U2281 (N_2281,N_1969,N_1385);
nor U2282 (N_2282,N_1970,N_1307);
and U2283 (N_2283,N_1562,N_1597);
xor U2284 (N_2284,N_1079,N_1106);
nor U2285 (N_2285,N_1050,N_1281);
nand U2286 (N_2286,N_1548,N_1357);
or U2287 (N_2287,N_1365,N_1502);
nand U2288 (N_2288,N_1821,N_1393);
or U2289 (N_2289,N_1146,N_1289);
nand U2290 (N_2290,N_1685,N_1081);
or U2291 (N_2291,N_1779,N_1523);
and U2292 (N_2292,N_1998,N_1615);
nor U2293 (N_2293,N_1855,N_1991);
and U2294 (N_2294,N_1921,N_1442);
nor U2295 (N_2295,N_1835,N_1342);
and U2296 (N_2296,N_1000,N_1903);
nand U2297 (N_2297,N_1222,N_1637);
and U2298 (N_2298,N_1108,N_1701);
nor U2299 (N_2299,N_1474,N_1390);
nor U2300 (N_2300,N_1718,N_1906);
nand U2301 (N_2301,N_1509,N_1062);
nor U2302 (N_2302,N_1394,N_1640);
and U2303 (N_2303,N_1709,N_1080);
and U2304 (N_2304,N_1870,N_1323);
or U2305 (N_2305,N_1379,N_1434);
and U2306 (N_2306,N_1100,N_1343);
or U2307 (N_2307,N_1635,N_1315);
nor U2308 (N_2308,N_1317,N_1993);
and U2309 (N_2309,N_1225,N_1491);
nor U2310 (N_2310,N_1674,N_1551);
nand U2311 (N_2311,N_1974,N_1845);
nand U2312 (N_2312,N_1479,N_1899);
nand U2313 (N_2313,N_1345,N_1499);
or U2314 (N_2314,N_1556,N_1692);
or U2315 (N_2315,N_1017,N_1824);
or U2316 (N_2316,N_1565,N_1024);
nand U2317 (N_2317,N_1679,N_1457);
nand U2318 (N_2318,N_1603,N_1989);
or U2319 (N_2319,N_1775,N_1124);
nand U2320 (N_2320,N_1207,N_1978);
nand U2321 (N_2321,N_1489,N_1402);
and U2322 (N_2322,N_1761,N_1204);
nor U2323 (N_2323,N_1482,N_1416);
and U2324 (N_2324,N_1381,N_1044);
and U2325 (N_2325,N_1946,N_1932);
nor U2326 (N_2326,N_1950,N_1876);
xnor U2327 (N_2327,N_1255,N_1262);
or U2328 (N_2328,N_1719,N_1438);
nand U2329 (N_2329,N_1740,N_1045);
nor U2330 (N_2330,N_1488,N_1003);
or U2331 (N_2331,N_1388,N_1147);
nor U2332 (N_2332,N_1938,N_1203);
and U2333 (N_2333,N_1258,N_1341);
nor U2334 (N_2334,N_1123,N_1911);
nand U2335 (N_2335,N_1587,N_1238);
nand U2336 (N_2336,N_1268,N_1091);
or U2337 (N_2337,N_1140,N_1764);
or U2338 (N_2338,N_1660,N_1367);
nor U2339 (N_2339,N_1055,N_1518);
nand U2340 (N_2340,N_1229,N_1971);
nor U2341 (N_2341,N_1694,N_1831);
nand U2342 (N_2342,N_1647,N_1195);
or U2343 (N_2343,N_1558,N_1559);
xor U2344 (N_2344,N_1943,N_1400);
nand U2345 (N_2345,N_1427,N_1580);
and U2346 (N_2346,N_1158,N_1507);
nor U2347 (N_2347,N_1990,N_1611);
and U2348 (N_2348,N_1309,N_1501);
nor U2349 (N_2349,N_1196,N_1036);
and U2350 (N_2350,N_1213,N_1189);
nor U2351 (N_2351,N_1570,N_1629);
or U2352 (N_2352,N_1668,N_1819);
or U2353 (N_2353,N_1676,N_1472);
xnor U2354 (N_2354,N_1960,N_1076);
nand U2355 (N_2355,N_1656,N_1107);
nor U2356 (N_2356,N_1192,N_1752);
nand U2357 (N_2357,N_1283,N_1517);
and U2358 (N_2358,N_1769,N_1244);
nor U2359 (N_2359,N_1332,N_1074);
and U2360 (N_2360,N_1670,N_1126);
and U2361 (N_2361,N_1242,N_1543);
nor U2362 (N_2362,N_1928,N_1735);
and U2363 (N_2363,N_1754,N_1035);
or U2364 (N_2364,N_1949,N_1399);
or U2365 (N_2365,N_1531,N_1169);
or U2366 (N_2366,N_1326,N_1245);
nor U2367 (N_2367,N_1896,N_1184);
nand U2368 (N_2368,N_1574,N_1037);
nand U2369 (N_2369,N_1913,N_1118);
and U2370 (N_2370,N_1923,N_1793);
and U2371 (N_2371,N_1187,N_1528);
and U2372 (N_2372,N_1150,N_1626);
or U2373 (N_2373,N_1300,N_1333);
and U2374 (N_2374,N_1641,N_1550);
nor U2375 (N_2375,N_1133,N_1324);
nand U2376 (N_2376,N_1944,N_1995);
or U2377 (N_2377,N_1608,N_1311);
or U2378 (N_2378,N_1693,N_1710);
and U2379 (N_2379,N_1448,N_1591);
nand U2380 (N_2380,N_1155,N_1893);
or U2381 (N_2381,N_1708,N_1773);
or U2382 (N_2382,N_1758,N_1569);
nor U2383 (N_2383,N_1287,N_1490);
nand U2384 (N_2384,N_1814,N_1095);
and U2385 (N_2385,N_1269,N_1302);
nor U2386 (N_2386,N_1005,N_1372);
or U2387 (N_2387,N_1885,N_1401);
and U2388 (N_2388,N_1808,N_1818);
or U2389 (N_2389,N_1806,N_1408);
and U2390 (N_2390,N_1816,N_1391);
or U2391 (N_2391,N_1272,N_1695);
or U2392 (N_2392,N_1525,N_1964);
nand U2393 (N_2393,N_1486,N_1606);
nor U2394 (N_2394,N_1075,N_1865);
nand U2395 (N_2395,N_1984,N_1895);
xor U2396 (N_2396,N_1148,N_1468);
and U2397 (N_2397,N_1065,N_1483);
or U2398 (N_2398,N_1801,N_1540);
and U2399 (N_2399,N_1149,N_1572);
or U2400 (N_2400,N_1398,N_1800);
and U2401 (N_2401,N_1757,N_1832);
nand U2402 (N_2402,N_1874,N_1137);
nor U2403 (N_2403,N_1206,N_1450);
or U2404 (N_2404,N_1891,N_1986);
nor U2405 (N_2405,N_1532,N_1768);
or U2406 (N_2406,N_1745,N_1237);
nand U2407 (N_2407,N_1275,N_1021);
or U2408 (N_2408,N_1972,N_1926);
or U2409 (N_2409,N_1784,N_1878);
and U2410 (N_2410,N_1798,N_1951);
nor U2411 (N_2411,N_1426,N_1366);
and U2412 (N_2412,N_1098,N_1575);
or U2413 (N_2413,N_1016,N_1476);
nor U2414 (N_2414,N_1031,N_1027);
and U2415 (N_2415,N_1354,N_1817);
and U2416 (N_2416,N_1783,N_1897);
nor U2417 (N_2417,N_1185,N_1176);
nand U2418 (N_2418,N_1270,N_1455);
nor U2419 (N_2419,N_1654,N_1215);
nand U2420 (N_2420,N_1851,N_1152);
nor U2421 (N_2421,N_1073,N_1588);
nor U2422 (N_2422,N_1884,N_1436);
or U2423 (N_2423,N_1116,N_1598);
or U2424 (N_2424,N_1590,N_1041);
nor U2425 (N_2425,N_1967,N_1922);
or U2426 (N_2426,N_1650,N_1435);
or U2427 (N_2427,N_1866,N_1282);
nand U2428 (N_2428,N_1316,N_1384);
and U2429 (N_2429,N_1705,N_1299);
nor U2430 (N_2430,N_1162,N_1009);
nor U2431 (N_2431,N_1383,N_1008);
xor U2432 (N_2432,N_1369,N_1086);
or U2433 (N_2433,N_1713,N_1252);
or U2434 (N_2434,N_1120,N_1910);
nor U2435 (N_2435,N_1219,N_1805);
or U2436 (N_2436,N_1873,N_1462);
or U2437 (N_2437,N_1119,N_1918);
nor U2438 (N_2438,N_1954,N_1973);
nand U2439 (N_2439,N_1956,N_1451);
nand U2440 (N_2440,N_1632,N_1057);
nor U2441 (N_2441,N_1230,N_1820);
nand U2442 (N_2442,N_1684,N_1962);
nand U2443 (N_2443,N_1843,N_1948);
nand U2444 (N_2444,N_1652,N_1277);
nand U2445 (N_2445,N_1122,N_1529);
and U2446 (N_2446,N_1582,N_1026);
or U2447 (N_2447,N_1894,N_1883);
nand U2448 (N_2448,N_1809,N_1156);
and U2449 (N_2449,N_1682,N_1766);
nor U2450 (N_2450,N_1056,N_1645);
nor U2451 (N_2451,N_1669,N_1581);
or U2452 (N_2452,N_1069,N_1631);
or U2453 (N_2453,N_1181,N_1872);
nand U2454 (N_2454,N_1110,N_1746);
and U2455 (N_2455,N_1104,N_1767);
or U2456 (N_2456,N_1294,N_1762);
or U2457 (N_2457,N_1810,N_1305);
nand U2458 (N_2458,N_1987,N_1430);
nand U2459 (N_2459,N_1358,N_1905);
and U2460 (N_2460,N_1934,N_1308);
and U2461 (N_2461,N_1513,N_1852);
nand U2462 (N_2462,N_1863,N_1274);
nor U2463 (N_2463,N_1428,N_1521);
nand U2464 (N_2464,N_1303,N_1979);
nor U2465 (N_2465,N_1025,N_1678);
nor U2466 (N_2466,N_1135,N_1236);
and U2467 (N_2467,N_1432,N_1515);
nand U2468 (N_2468,N_1596,N_1983);
and U2469 (N_2469,N_1750,N_1248);
or U2470 (N_2470,N_1605,N_1688);
nand U2471 (N_2471,N_1263,N_1136);
nand U2472 (N_2472,N_1023,N_1293);
and U2473 (N_2473,N_1459,N_1151);
nand U2474 (N_2474,N_1560,N_1837);
and U2475 (N_2475,N_1634,N_1359);
and U2476 (N_2476,N_1703,N_1546);
and U2477 (N_2477,N_1955,N_1547);
or U2478 (N_2478,N_1419,N_1790);
and U2479 (N_2479,N_1078,N_1726);
nor U2480 (N_2480,N_1524,N_1505);
and U2481 (N_2481,N_1553,N_1981);
or U2482 (N_2482,N_1536,N_1914);
or U2483 (N_2483,N_1205,N_1813);
nand U2484 (N_2484,N_1439,N_1825);
nor U2485 (N_2485,N_1094,N_1732);
nor U2486 (N_2486,N_1304,N_1395);
or U2487 (N_2487,N_1286,N_1347);
or U2488 (N_2488,N_1696,N_1624);
or U2489 (N_2489,N_1112,N_1644);
xor U2490 (N_2490,N_1890,N_1279);
and U2491 (N_2491,N_1859,N_1386);
and U2492 (N_2492,N_1862,N_1697);
or U2493 (N_2493,N_1828,N_1290);
and U2494 (N_2494,N_1083,N_1664);
nor U2495 (N_2495,N_1321,N_1249);
or U2496 (N_2496,N_1965,N_1405);
and U2497 (N_2497,N_1655,N_1223);
or U2498 (N_2498,N_1976,N_1721);
nand U2499 (N_2499,N_1871,N_1561);
xnor U2500 (N_2500,N_1469,N_1545);
nand U2501 (N_2501,N_1124,N_1039);
nand U2502 (N_2502,N_1411,N_1435);
and U2503 (N_2503,N_1818,N_1830);
or U2504 (N_2504,N_1369,N_1030);
nand U2505 (N_2505,N_1106,N_1800);
or U2506 (N_2506,N_1139,N_1521);
or U2507 (N_2507,N_1271,N_1519);
nor U2508 (N_2508,N_1700,N_1832);
and U2509 (N_2509,N_1685,N_1541);
nand U2510 (N_2510,N_1334,N_1071);
nor U2511 (N_2511,N_1024,N_1374);
xor U2512 (N_2512,N_1818,N_1184);
nand U2513 (N_2513,N_1128,N_1285);
nor U2514 (N_2514,N_1555,N_1509);
nor U2515 (N_2515,N_1636,N_1792);
nand U2516 (N_2516,N_1875,N_1848);
nand U2517 (N_2517,N_1936,N_1535);
nand U2518 (N_2518,N_1447,N_1513);
and U2519 (N_2519,N_1377,N_1133);
nand U2520 (N_2520,N_1456,N_1347);
nor U2521 (N_2521,N_1933,N_1223);
nand U2522 (N_2522,N_1156,N_1889);
nand U2523 (N_2523,N_1774,N_1515);
and U2524 (N_2524,N_1694,N_1789);
nand U2525 (N_2525,N_1857,N_1475);
nand U2526 (N_2526,N_1782,N_1826);
nand U2527 (N_2527,N_1181,N_1807);
and U2528 (N_2528,N_1724,N_1524);
or U2529 (N_2529,N_1731,N_1946);
and U2530 (N_2530,N_1977,N_1258);
and U2531 (N_2531,N_1083,N_1209);
nor U2532 (N_2532,N_1310,N_1372);
nand U2533 (N_2533,N_1564,N_1514);
nor U2534 (N_2534,N_1962,N_1222);
and U2535 (N_2535,N_1024,N_1989);
and U2536 (N_2536,N_1957,N_1228);
and U2537 (N_2537,N_1265,N_1193);
nand U2538 (N_2538,N_1580,N_1166);
nor U2539 (N_2539,N_1792,N_1966);
and U2540 (N_2540,N_1348,N_1701);
and U2541 (N_2541,N_1234,N_1673);
and U2542 (N_2542,N_1460,N_1790);
and U2543 (N_2543,N_1154,N_1183);
or U2544 (N_2544,N_1880,N_1661);
nand U2545 (N_2545,N_1911,N_1690);
and U2546 (N_2546,N_1002,N_1345);
or U2547 (N_2547,N_1475,N_1452);
or U2548 (N_2548,N_1174,N_1749);
and U2549 (N_2549,N_1913,N_1053);
nor U2550 (N_2550,N_1186,N_1471);
nand U2551 (N_2551,N_1888,N_1364);
and U2552 (N_2552,N_1419,N_1058);
or U2553 (N_2553,N_1786,N_1530);
nor U2554 (N_2554,N_1557,N_1305);
nand U2555 (N_2555,N_1969,N_1622);
or U2556 (N_2556,N_1979,N_1040);
nand U2557 (N_2557,N_1097,N_1224);
and U2558 (N_2558,N_1330,N_1188);
nor U2559 (N_2559,N_1880,N_1374);
nand U2560 (N_2560,N_1630,N_1195);
nand U2561 (N_2561,N_1491,N_1379);
nor U2562 (N_2562,N_1360,N_1000);
nand U2563 (N_2563,N_1016,N_1093);
or U2564 (N_2564,N_1978,N_1278);
nor U2565 (N_2565,N_1973,N_1452);
nor U2566 (N_2566,N_1411,N_1421);
and U2567 (N_2567,N_1312,N_1675);
xor U2568 (N_2568,N_1477,N_1194);
and U2569 (N_2569,N_1875,N_1311);
or U2570 (N_2570,N_1028,N_1832);
nand U2571 (N_2571,N_1828,N_1297);
nand U2572 (N_2572,N_1642,N_1237);
nand U2573 (N_2573,N_1499,N_1644);
or U2574 (N_2574,N_1082,N_1016);
or U2575 (N_2575,N_1509,N_1830);
nor U2576 (N_2576,N_1873,N_1869);
and U2577 (N_2577,N_1710,N_1651);
or U2578 (N_2578,N_1150,N_1853);
nor U2579 (N_2579,N_1435,N_1469);
or U2580 (N_2580,N_1864,N_1238);
or U2581 (N_2581,N_1918,N_1811);
and U2582 (N_2582,N_1117,N_1837);
and U2583 (N_2583,N_1365,N_1294);
nor U2584 (N_2584,N_1891,N_1487);
nor U2585 (N_2585,N_1094,N_1735);
and U2586 (N_2586,N_1691,N_1560);
or U2587 (N_2587,N_1730,N_1221);
and U2588 (N_2588,N_1159,N_1380);
nand U2589 (N_2589,N_1213,N_1415);
nand U2590 (N_2590,N_1094,N_1541);
and U2591 (N_2591,N_1358,N_1192);
nand U2592 (N_2592,N_1098,N_1322);
and U2593 (N_2593,N_1580,N_1562);
and U2594 (N_2594,N_1529,N_1519);
or U2595 (N_2595,N_1064,N_1662);
nand U2596 (N_2596,N_1744,N_1873);
nand U2597 (N_2597,N_1456,N_1896);
and U2598 (N_2598,N_1010,N_1588);
nand U2599 (N_2599,N_1502,N_1246);
or U2600 (N_2600,N_1365,N_1650);
or U2601 (N_2601,N_1542,N_1218);
nand U2602 (N_2602,N_1333,N_1088);
nor U2603 (N_2603,N_1268,N_1283);
nor U2604 (N_2604,N_1235,N_1334);
and U2605 (N_2605,N_1249,N_1337);
and U2606 (N_2606,N_1121,N_1975);
and U2607 (N_2607,N_1304,N_1047);
nor U2608 (N_2608,N_1419,N_1247);
nand U2609 (N_2609,N_1050,N_1314);
nor U2610 (N_2610,N_1777,N_1092);
nand U2611 (N_2611,N_1993,N_1254);
or U2612 (N_2612,N_1104,N_1317);
nor U2613 (N_2613,N_1835,N_1164);
nor U2614 (N_2614,N_1380,N_1892);
and U2615 (N_2615,N_1023,N_1961);
and U2616 (N_2616,N_1883,N_1566);
nand U2617 (N_2617,N_1711,N_1247);
nand U2618 (N_2618,N_1371,N_1611);
nand U2619 (N_2619,N_1768,N_1799);
nand U2620 (N_2620,N_1063,N_1344);
and U2621 (N_2621,N_1441,N_1145);
nand U2622 (N_2622,N_1348,N_1660);
and U2623 (N_2623,N_1624,N_1003);
or U2624 (N_2624,N_1954,N_1723);
or U2625 (N_2625,N_1254,N_1002);
or U2626 (N_2626,N_1019,N_1588);
nand U2627 (N_2627,N_1093,N_1850);
or U2628 (N_2628,N_1133,N_1454);
nor U2629 (N_2629,N_1981,N_1805);
nor U2630 (N_2630,N_1203,N_1629);
nand U2631 (N_2631,N_1331,N_1588);
and U2632 (N_2632,N_1723,N_1093);
or U2633 (N_2633,N_1888,N_1335);
nand U2634 (N_2634,N_1444,N_1180);
and U2635 (N_2635,N_1989,N_1828);
nor U2636 (N_2636,N_1460,N_1215);
or U2637 (N_2637,N_1009,N_1750);
nand U2638 (N_2638,N_1205,N_1195);
and U2639 (N_2639,N_1508,N_1644);
nand U2640 (N_2640,N_1045,N_1568);
nand U2641 (N_2641,N_1584,N_1520);
or U2642 (N_2642,N_1265,N_1800);
and U2643 (N_2643,N_1053,N_1556);
and U2644 (N_2644,N_1600,N_1075);
and U2645 (N_2645,N_1657,N_1256);
nor U2646 (N_2646,N_1535,N_1108);
nor U2647 (N_2647,N_1699,N_1480);
and U2648 (N_2648,N_1933,N_1259);
and U2649 (N_2649,N_1761,N_1048);
nand U2650 (N_2650,N_1244,N_1968);
nand U2651 (N_2651,N_1811,N_1758);
or U2652 (N_2652,N_1579,N_1235);
nand U2653 (N_2653,N_1790,N_1365);
and U2654 (N_2654,N_1003,N_1530);
nand U2655 (N_2655,N_1907,N_1800);
and U2656 (N_2656,N_1110,N_1371);
or U2657 (N_2657,N_1197,N_1477);
and U2658 (N_2658,N_1391,N_1420);
nor U2659 (N_2659,N_1325,N_1383);
or U2660 (N_2660,N_1426,N_1393);
nor U2661 (N_2661,N_1442,N_1932);
nand U2662 (N_2662,N_1972,N_1643);
or U2663 (N_2663,N_1256,N_1622);
and U2664 (N_2664,N_1154,N_1025);
nand U2665 (N_2665,N_1044,N_1288);
nor U2666 (N_2666,N_1922,N_1536);
xnor U2667 (N_2667,N_1310,N_1193);
xnor U2668 (N_2668,N_1694,N_1885);
nor U2669 (N_2669,N_1103,N_1476);
nand U2670 (N_2670,N_1537,N_1911);
or U2671 (N_2671,N_1013,N_1910);
or U2672 (N_2672,N_1988,N_1931);
and U2673 (N_2673,N_1717,N_1172);
or U2674 (N_2674,N_1961,N_1579);
xnor U2675 (N_2675,N_1928,N_1505);
nor U2676 (N_2676,N_1827,N_1556);
nand U2677 (N_2677,N_1450,N_1011);
nor U2678 (N_2678,N_1311,N_1418);
nor U2679 (N_2679,N_1291,N_1830);
nor U2680 (N_2680,N_1313,N_1895);
or U2681 (N_2681,N_1633,N_1932);
and U2682 (N_2682,N_1720,N_1552);
nand U2683 (N_2683,N_1636,N_1774);
nand U2684 (N_2684,N_1014,N_1927);
nor U2685 (N_2685,N_1111,N_1703);
nand U2686 (N_2686,N_1373,N_1954);
or U2687 (N_2687,N_1715,N_1103);
or U2688 (N_2688,N_1010,N_1995);
nor U2689 (N_2689,N_1958,N_1420);
and U2690 (N_2690,N_1122,N_1985);
and U2691 (N_2691,N_1184,N_1137);
xnor U2692 (N_2692,N_1451,N_1744);
and U2693 (N_2693,N_1598,N_1368);
nand U2694 (N_2694,N_1235,N_1007);
nor U2695 (N_2695,N_1914,N_1237);
xnor U2696 (N_2696,N_1788,N_1413);
nand U2697 (N_2697,N_1843,N_1471);
or U2698 (N_2698,N_1165,N_1521);
nand U2699 (N_2699,N_1210,N_1022);
nor U2700 (N_2700,N_1127,N_1872);
and U2701 (N_2701,N_1141,N_1486);
nand U2702 (N_2702,N_1688,N_1076);
nor U2703 (N_2703,N_1278,N_1492);
nand U2704 (N_2704,N_1910,N_1344);
and U2705 (N_2705,N_1262,N_1377);
nor U2706 (N_2706,N_1425,N_1050);
or U2707 (N_2707,N_1379,N_1699);
nand U2708 (N_2708,N_1052,N_1951);
and U2709 (N_2709,N_1405,N_1857);
and U2710 (N_2710,N_1241,N_1600);
nand U2711 (N_2711,N_1376,N_1360);
nand U2712 (N_2712,N_1314,N_1160);
or U2713 (N_2713,N_1349,N_1910);
and U2714 (N_2714,N_1714,N_1236);
nand U2715 (N_2715,N_1634,N_1031);
nand U2716 (N_2716,N_1556,N_1498);
nand U2717 (N_2717,N_1970,N_1700);
or U2718 (N_2718,N_1688,N_1458);
or U2719 (N_2719,N_1395,N_1976);
and U2720 (N_2720,N_1939,N_1235);
nor U2721 (N_2721,N_1919,N_1226);
nor U2722 (N_2722,N_1089,N_1375);
and U2723 (N_2723,N_1681,N_1704);
nor U2724 (N_2724,N_1378,N_1356);
nand U2725 (N_2725,N_1482,N_1418);
nor U2726 (N_2726,N_1732,N_1244);
nand U2727 (N_2727,N_1294,N_1800);
nand U2728 (N_2728,N_1268,N_1967);
or U2729 (N_2729,N_1180,N_1227);
or U2730 (N_2730,N_1528,N_1052);
nand U2731 (N_2731,N_1128,N_1524);
and U2732 (N_2732,N_1450,N_1281);
and U2733 (N_2733,N_1455,N_1755);
or U2734 (N_2734,N_1951,N_1391);
or U2735 (N_2735,N_1027,N_1864);
nand U2736 (N_2736,N_1498,N_1974);
nor U2737 (N_2737,N_1388,N_1472);
nand U2738 (N_2738,N_1662,N_1623);
and U2739 (N_2739,N_1331,N_1050);
nand U2740 (N_2740,N_1418,N_1123);
or U2741 (N_2741,N_1768,N_1133);
nand U2742 (N_2742,N_1912,N_1498);
nand U2743 (N_2743,N_1591,N_1982);
nand U2744 (N_2744,N_1196,N_1544);
and U2745 (N_2745,N_1337,N_1259);
xor U2746 (N_2746,N_1034,N_1261);
nand U2747 (N_2747,N_1367,N_1242);
nand U2748 (N_2748,N_1662,N_1025);
or U2749 (N_2749,N_1717,N_1295);
nor U2750 (N_2750,N_1490,N_1899);
nor U2751 (N_2751,N_1157,N_1582);
nor U2752 (N_2752,N_1511,N_1639);
and U2753 (N_2753,N_1768,N_1106);
nand U2754 (N_2754,N_1397,N_1872);
and U2755 (N_2755,N_1262,N_1846);
and U2756 (N_2756,N_1870,N_1393);
nor U2757 (N_2757,N_1436,N_1671);
nand U2758 (N_2758,N_1687,N_1297);
nand U2759 (N_2759,N_1599,N_1968);
nor U2760 (N_2760,N_1878,N_1802);
and U2761 (N_2761,N_1321,N_1832);
nand U2762 (N_2762,N_1135,N_1228);
or U2763 (N_2763,N_1126,N_1287);
and U2764 (N_2764,N_1855,N_1395);
and U2765 (N_2765,N_1153,N_1414);
nor U2766 (N_2766,N_1635,N_1781);
nand U2767 (N_2767,N_1567,N_1538);
and U2768 (N_2768,N_1649,N_1852);
nor U2769 (N_2769,N_1978,N_1941);
nor U2770 (N_2770,N_1719,N_1585);
nor U2771 (N_2771,N_1183,N_1869);
or U2772 (N_2772,N_1664,N_1291);
nand U2773 (N_2773,N_1516,N_1365);
nor U2774 (N_2774,N_1575,N_1553);
and U2775 (N_2775,N_1094,N_1639);
and U2776 (N_2776,N_1021,N_1922);
and U2777 (N_2777,N_1118,N_1937);
xor U2778 (N_2778,N_1272,N_1095);
nand U2779 (N_2779,N_1036,N_1481);
nand U2780 (N_2780,N_1763,N_1289);
xnor U2781 (N_2781,N_1973,N_1057);
nand U2782 (N_2782,N_1667,N_1595);
nor U2783 (N_2783,N_1368,N_1995);
nor U2784 (N_2784,N_1566,N_1730);
nand U2785 (N_2785,N_1447,N_1604);
xor U2786 (N_2786,N_1406,N_1133);
nand U2787 (N_2787,N_1104,N_1582);
or U2788 (N_2788,N_1733,N_1406);
nand U2789 (N_2789,N_1160,N_1940);
and U2790 (N_2790,N_1262,N_1369);
or U2791 (N_2791,N_1743,N_1644);
nor U2792 (N_2792,N_1687,N_1880);
nand U2793 (N_2793,N_1346,N_1730);
and U2794 (N_2794,N_1811,N_1180);
nor U2795 (N_2795,N_1208,N_1132);
nand U2796 (N_2796,N_1037,N_1775);
nand U2797 (N_2797,N_1674,N_1985);
or U2798 (N_2798,N_1310,N_1988);
nand U2799 (N_2799,N_1781,N_1356);
and U2800 (N_2800,N_1000,N_1539);
nand U2801 (N_2801,N_1847,N_1084);
and U2802 (N_2802,N_1426,N_1510);
nor U2803 (N_2803,N_1854,N_1987);
nand U2804 (N_2804,N_1653,N_1554);
or U2805 (N_2805,N_1014,N_1356);
or U2806 (N_2806,N_1045,N_1205);
or U2807 (N_2807,N_1320,N_1134);
and U2808 (N_2808,N_1630,N_1475);
nand U2809 (N_2809,N_1543,N_1188);
nor U2810 (N_2810,N_1433,N_1666);
nand U2811 (N_2811,N_1233,N_1285);
and U2812 (N_2812,N_1863,N_1700);
nand U2813 (N_2813,N_1288,N_1626);
nor U2814 (N_2814,N_1956,N_1121);
nor U2815 (N_2815,N_1754,N_1157);
nor U2816 (N_2816,N_1752,N_1415);
nor U2817 (N_2817,N_1409,N_1402);
nand U2818 (N_2818,N_1214,N_1203);
or U2819 (N_2819,N_1780,N_1900);
or U2820 (N_2820,N_1080,N_1214);
and U2821 (N_2821,N_1405,N_1006);
and U2822 (N_2822,N_1699,N_1417);
or U2823 (N_2823,N_1167,N_1995);
or U2824 (N_2824,N_1987,N_1418);
or U2825 (N_2825,N_1950,N_1873);
nand U2826 (N_2826,N_1256,N_1244);
nand U2827 (N_2827,N_1627,N_1349);
and U2828 (N_2828,N_1409,N_1913);
and U2829 (N_2829,N_1619,N_1906);
nor U2830 (N_2830,N_1463,N_1718);
or U2831 (N_2831,N_1310,N_1300);
and U2832 (N_2832,N_1223,N_1416);
nand U2833 (N_2833,N_1603,N_1467);
nand U2834 (N_2834,N_1609,N_1435);
nand U2835 (N_2835,N_1288,N_1587);
nand U2836 (N_2836,N_1780,N_1564);
nand U2837 (N_2837,N_1491,N_1435);
and U2838 (N_2838,N_1551,N_1914);
nand U2839 (N_2839,N_1860,N_1008);
nor U2840 (N_2840,N_1903,N_1993);
nor U2841 (N_2841,N_1712,N_1375);
nand U2842 (N_2842,N_1437,N_1280);
nor U2843 (N_2843,N_1233,N_1193);
nor U2844 (N_2844,N_1772,N_1548);
nor U2845 (N_2845,N_1071,N_1929);
nor U2846 (N_2846,N_1753,N_1412);
nor U2847 (N_2847,N_1645,N_1703);
and U2848 (N_2848,N_1282,N_1673);
and U2849 (N_2849,N_1168,N_1955);
nor U2850 (N_2850,N_1460,N_1787);
xnor U2851 (N_2851,N_1439,N_1208);
nor U2852 (N_2852,N_1188,N_1118);
nor U2853 (N_2853,N_1605,N_1672);
nor U2854 (N_2854,N_1755,N_1127);
nor U2855 (N_2855,N_1099,N_1921);
and U2856 (N_2856,N_1369,N_1818);
nand U2857 (N_2857,N_1784,N_1714);
or U2858 (N_2858,N_1376,N_1729);
nor U2859 (N_2859,N_1050,N_1705);
and U2860 (N_2860,N_1271,N_1337);
nor U2861 (N_2861,N_1091,N_1260);
nor U2862 (N_2862,N_1581,N_1193);
or U2863 (N_2863,N_1427,N_1108);
nand U2864 (N_2864,N_1739,N_1100);
nand U2865 (N_2865,N_1841,N_1746);
nand U2866 (N_2866,N_1927,N_1786);
and U2867 (N_2867,N_1971,N_1696);
nand U2868 (N_2868,N_1739,N_1791);
and U2869 (N_2869,N_1584,N_1114);
xor U2870 (N_2870,N_1494,N_1708);
or U2871 (N_2871,N_1155,N_1138);
or U2872 (N_2872,N_1014,N_1277);
nand U2873 (N_2873,N_1783,N_1055);
and U2874 (N_2874,N_1776,N_1294);
nor U2875 (N_2875,N_1220,N_1199);
nor U2876 (N_2876,N_1135,N_1775);
nand U2877 (N_2877,N_1269,N_1635);
and U2878 (N_2878,N_1885,N_1367);
or U2879 (N_2879,N_1374,N_1021);
nand U2880 (N_2880,N_1540,N_1473);
or U2881 (N_2881,N_1564,N_1095);
and U2882 (N_2882,N_1358,N_1950);
and U2883 (N_2883,N_1614,N_1508);
nor U2884 (N_2884,N_1664,N_1441);
nand U2885 (N_2885,N_1533,N_1241);
or U2886 (N_2886,N_1910,N_1207);
nand U2887 (N_2887,N_1336,N_1122);
nor U2888 (N_2888,N_1803,N_1408);
and U2889 (N_2889,N_1090,N_1566);
and U2890 (N_2890,N_1719,N_1161);
nand U2891 (N_2891,N_1515,N_1909);
nand U2892 (N_2892,N_1849,N_1630);
nor U2893 (N_2893,N_1063,N_1956);
nand U2894 (N_2894,N_1664,N_1818);
or U2895 (N_2895,N_1424,N_1110);
xnor U2896 (N_2896,N_1235,N_1324);
or U2897 (N_2897,N_1609,N_1814);
or U2898 (N_2898,N_1269,N_1479);
nand U2899 (N_2899,N_1063,N_1272);
nor U2900 (N_2900,N_1149,N_1930);
or U2901 (N_2901,N_1823,N_1734);
or U2902 (N_2902,N_1351,N_1452);
and U2903 (N_2903,N_1865,N_1383);
nor U2904 (N_2904,N_1773,N_1368);
nand U2905 (N_2905,N_1024,N_1043);
xnor U2906 (N_2906,N_1615,N_1564);
nor U2907 (N_2907,N_1547,N_1379);
or U2908 (N_2908,N_1220,N_1914);
nor U2909 (N_2909,N_1507,N_1610);
and U2910 (N_2910,N_1034,N_1970);
nor U2911 (N_2911,N_1528,N_1206);
nand U2912 (N_2912,N_1540,N_1300);
nor U2913 (N_2913,N_1252,N_1545);
and U2914 (N_2914,N_1250,N_1707);
nor U2915 (N_2915,N_1440,N_1688);
and U2916 (N_2916,N_1047,N_1921);
and U2917 (N_2917,N_1902,N_1966);
and U2918 (N_2918,N_1491,N_1068);
nor U2919 (N_2919,N_1858,N_1958);
nand U2920 (N_2920,N_1463,N_1100);
nor U2921 (N_2921,N_1026,N_1216);
nor U2922 (N_2922,N_1081,N_1712);
nor U2923 (N_2923,N_1053,N_1458);
nand U2924 (N_2924,N_1787,N_1374);
and U2925 (N_2925,N_1626,N_1532);
nor U2926 (N_2926,N_1760,N_1764);
or U2927 (N_2927,N_1755,N_1463);
or U2928 (N_2928,N_1318,N_1911);
nand U2929 (N_2929,N_1440,N_1222);
nor U2930 (N_2930,N_1438,N_1721);
nand U2931 (N_2931,N_1694,N_1075);
or U2932 (N_2932,N_1954,N_1778);
nor U2933 (N_2933,N_1900,N_1145);
and U2934 (N_2934,N_1646,N_1248);
nor U2935 (N_2935,N_1786,N_1453);
or U2936 (N_2936,N_1080,N_1026);
or U2937 (N_2937,N_1138,N_1963);
and U2938 (N_2938,N_1641,N_1989);
or U2939 (N_2939,N_1367,N_1898);
nand U2940 (N_2940,N_1784,N_1299);
nand U2941 (N_2941,N_1512,N_1423);
and U2942 (N_2942,N_1612,N_1679);
nor U2943 (N_2943,N_1738,N_1166);
and U2944 (N_2944,N_1122,N_1468);
or U2945 (N_2945,N_1394,N_1491);
nor U2946 (N_2946,N_1724,N_1641);
and U2947 (N_2947,N_1258,N_1835);
nand U2948 (N_2948,N_1688,N_1851);
and U2949 (N_2949,N_1027,N_1628);
nand U2950 (N_2950,N_1863,N_1172);
or U2951 (N_2951,N_1820,N_1005);
nand U2952 (N_2952,N_1112,N_1818);
nor U2953 (N_2953,N_1508,N_1991);
or U2954 (N_2954,N_1564,N_1903);
and U2955 (N_2955,N_1159,N_1244);
nor U2956 (N_2956,N_1092,N_1399);
nand U2957 (N_2957,N_1868,N_1582);
and U2958 (N_2958,N_1305,N_1115);
nor U2959 (N_2959,N_1905,N_1509);
or U2960 (N_2960,N_1712,N_1889);
or U2961 (N_2961,N_1588,N_1318);
nor U2962 (N_2962,N_1450,N_1981);
nand U2963 (N_2963,N_1000,N_1408);
nand U2964 (N_2964,N_1090,N_1623);
nand U2965 (N_2965,N_1641,N_1877);
nor U2966 (N_2966,N_1495,N_1607);
nor U2967 (N_2967,N_1481,N_1576);
nand U2968 (N_2968,N_1384,N_1464);
nand U2969 (N_2969,N_1243,N_1827);
or U2970 (N_2970,N_1712,N_1193);
nand U2971 (N_2971,N_1264,N_1429);
nand U2972 (N_2972,N_1713,N_1927);
or U2973 (N_2973,N_1407,N_1107);
and U2974 (N_2974,N_1771,N_1015);
nand U2975 (N_2975,N_1531,N_1458);
nand U2976 (N_2976,N_1019,N_1561);
nor U2977 (N_2977,N_1665,N_1315);
nand U2978 (N_2978,N_1373,N_1587);
or U2979 (N_2979,N_1940,N_1847);
or U2980 (N_2980,N_1792,N_1317);
and U2981 (N_2981,N_1148,N_1442);
or U2982 (N_2982,N_1683,N_1554);
nor U2983 (N_2983,N_1423,N_1477);
and U2984 (N_2984,N_1498,N_1820);
or U2985 (N_2985,N_1705,N_1089);
nor U2986 (N_2986,N_1097,N_1914);
and U2987 (N_2987,N_1646,N_1331);
nand U2988 (N_2988,N_1000,N_1568);
nor U2989 (N_2989,N_1352,N_1083);
nand U2990 (N_2990,N_1823,N_1095);
nor U2991 (N_2991,N_1737,N_1053);
and U2992 (N_2992,N_1884,N_1175);
and U2993 (N_2993,N_1503,N_1413);
nand U2994 (N_2994,N_1232,N_1058);
nand U2995 (N_2995,N_1992,N_1568);
and U2996 (N_2996,N_1307,N_1063);
and U2997 (N_2997,N_1691,N_1887);
nand U2998 (N_2998,N_1755,N_1217);
nor U2999 (N_2999,N_1719,N_1631);
or UO_0 (O_0,N_2706,N_2889);
nor UO_1 (O_1,N_2430,N_2489);
nand UO_2 (O_2,N_2109,N_2285);
nand UO_3 (O_3,N_2659,N_2257);
and UO_4 (O_4,N_2241,N_2104);
and UO_5 (O_5,N_2772,N_2808);
and UO_6 (O_6,N_2433,N_2360);
nor UO_7 (O_7,N_2686,N_2338);
nor UO_8 (O_8,N_2969,N_2531);
nor UO_9 (O_9,N_2163,N_2983);
or UO_10 (O_10,N_2751,N_2054);
or UO_11 (O_11,N_2881,N_2414);
nand UO_12 (O_12,N_2766,N_2890);
nand UO_13 (O_13,N_2865,N_2830);
or UO_14 (O_14,N_2463,N_2700);
or UO_15 (O_15,N_2006,N_2643);
and UO_16 (O_16,N_2947,N_2987);
nor UO_17 (O_17,N_2316,N_2334);
nand UO_18 (O_18,N_2753,N_2549);
or UO_19 (O_19,N_2796,N_2500);
nand UO_20 (O_20,N_2041,N_2133);
nor UO_21 (O_21,N_2237,N_2178);
and UO_22 (O_22,N_2923,N_2413);
and UO_23 (O_23,N_2607,N_2261);
nor UO_24 (O_24,N_2359,N_2303);
nand UO_25 (O_25,N_2907,N_2708);
or UO_26 (O_26,N_2017,N_2797);
nor UO_27 (O_27,N_2053,N_2139);
xor UO_28 (O_28,N_2974,N_2354);
nor UO_29 (O_29,N_2355,N_2282);
and UO_30 (O_30,N_2441,N_2327);
and UO_31 (O_31,N_2204,N_2729);
or UO_32 (O_32,N_2863,N_2943);
or UO_33 (O_33,N_2228,N_2364);
xor UO_34 (O_34,N_2552,N_2744);
and UO_35 (O_35,N_2002,N_2994);
and UO_36 (O_36,N_2010,N_2530);
or UO_37 (O_37,N_2693,N_2353);
nand UO_38 (O_38,N_2995,N_2631);
nand UO_39 (O_39,N_2418,N_2810);
or UO_40 (O_40,N_2313,N_2019);
or UO_41 (O_41,N_2891,N_2249);
nor UO_42 (O_42,N_2428,N_2646);
nand UO_43 (O_43,N_2118,N_2378);
and UO_44 (O_44,N_2423,N_2080);
and UO_45 (O_45,N_2542,N_2505);
xor UO_46 (O_46,N_2874,N_2315);
or UO_47 (O_47,N_2314,N_2293);
nand UO_48 (O_48,N_2290,N_2370);
and UO_49 (O_49,N_2346,N_2246);
or UO_50 (O_50,N_2813,N_2880);
nor UO_51 (O_51,N_2373,N_2410);
nor UO_52 (O_52,N_2269,N_2778);
or UO_53 (O_53,N_2783,N_2658);
and UO_54 (O_54,N_2154,N_2539);
and UO_55 (O_55,N_2755,N_2136);
nand UO_56 (O_56,N_2915,N_2067);
nand UO_57 (O_57,N_2786,N_2690);
or UO_58 (O_58,N_2264,N_2048);
or UO_59 (O_59,N_2837,N_2034);
and UO_60 (O_60,N_2792,N_2305);
and UO_61 (O_61,N_2065,N_2595);
nand UO_62 (O_62,N_2193,N_2773);
nand UO_63 (O_63,N_2718,N_2450);
nor UO_64 (O_64,N_2510,N_2546);
nand UO_65 (O_65,N_2286,N_2826);
nor UO_66 (O_66,N_2005,N_2960);
and UO_67 (O_67,N_2040,N_2461);
and UO_68 (O_68,N_2710,N_2900);
and UO_69 (O_69,N_2168,N_2750);
nand UO_70 (O_70,N_2554,N_2165);
xnor UO_71 (O_71,N_2077,N_2196);
and UO_72 (O_72,N_2412,N_2634);
or UO_73 (O_73,N_2657,N_2222);
nand UO_74 (O_74,N_2024,N_2834);
nor UO_75 (O_75,N_2166,N_2388);
nand UO_76 (O_76,N_2978,N_2691);
nor UO_77 (O_77,N_2422,N_2798);
and UO_78 (O_78,N_2059,N_2190);
or UO_79 (O_79,N_2117,N_2565);
and UO_80 (O_80,N_2471,N_2704);
and UO_81 (O_81,N_2112,N_2090);
and UO_82 (O_82,N_2209,N_2609);
nor UO_83 (O_83,N_2114,N_2135);
nor UO_84 (O_84,N_2072,N_2426);
and UO_85 (O_85,N_2008,N_2288);
nand UO_86 (O_86,N_2919,N_2374);
or UO_87 (O_87,N_2663,N_2490);
nand UO_88 (O_88,N_2352,N_2765);
and UO_89 (O_89,N_2192,N_2211);
nor UO_90 (O_90,N_2523,N_2601);
nor UO_91 (O_91,N_2736,N_2582);
or UO_92 (O_92,N_2152,N_2042);
or UO_93 (O_93,N_2392,N_2970);
and UO_94 (O_94,N_2851,N_2205);
nand UO_95 (O_95,N_2624,N_2864);
nor UO_96 (O_96,N_2217,N_2534);
or UO_97 (O_97,N_2730,N_2733);
nor UO_98 (O_98,N_2876,N_2636);
or UO_99 (O_99,N_2940,N_2926);
and UO_100 (O_100,N_2666,N_2479);
or UO_101 (O_101,N_2091,N_2411);
or UO_102 (O_102,N_2897,N_2513);
nand UO_103 (O_103,N_2835,N_2220);
nand UO_104 (O_104,N_2898,N_2400);
and UO_105 (O_105,N_2920,N_2594);
nand UO_106 (O_106,N_2394,N_2930);
nand UO_107 (O_107,N_2300,N_2218);
and UO_108 (O_108,N_2195,N_2665);
or UO_109 (O_109,N_2329,N_2291);
or UO_110 (O_110,N_2320,N_2506);
nand UO_111 (O_111,N_2137,N_2103);
nand UO_112 (O_112,N_2215,N_2832);
nor UO_113 (O_113,N_2340,N_2802);
nor UO_114 (O_114,N_2862,N_2186);
nor UO_115 (O_115,N_2021,N_2870);
and UO_116 (O_116,N_2586,N_2683);
xnor UO_117 (O_117,N_2086,N_2424);
nor UO_118 (O_118,N_2000,N_2941);
or UO_119 (O_119,N_2973,N_2279);
nor UO_120 (O_120,N_2157,N_2158);
and UO_121 (O_121,N_2541,N_2653);
and UO_122 (O_122,N_2466,N_2520);
or UO_123 (O_123,N_2570,N_2715);
and UO_124 (O_124,N_2177,N_2633);
nand UO_125 (O_125,N_2677,N_2032);
nor UO_126 (O_126,N_2240,N_2629);
and UO_127 (O_127,N_2023,N_2082);
xnor UO_128 (O_128,N_2784,N_2815);
nand UO_129 (O_129,N_2442,N_2982);
nand UO_130 (O_130,N_2793,N_2669);
nand UO_131 (O_131,N_2265,N_2321);
or UO_132 (O_132,N_2516,N_2200);
nand UO_133 (O_133,N_2632,N_2939);
and UO_134 (O_134,N_2111,N_2169);
and UO_135 (O_135,N_2901,N_2097);
and UO_136 (O_136,N_2641,N_2130);
xnor UO_137 (O_137,N_2980,N_2122);
nor UO_138 (O_138,N_2229,N_2758);
and UO_139 (O_139,N_2203,N_2971);
and UO_140 (O_140,N_2230,N_2509);
and UO_141 (O_141,N_2532,N_2167);
or UO_142 (O_142,N_2391,N_2854);
or UO_143 (O_143,N_2698,N_2421);
and UO_144 (O_144,N_2039,N_2035);
nor UO_145 (O_145,N_2608,N_2262);
or UO_146 (O_146,N_2727,N_2613);
nor UO_147 (O_147,N_2376,N_2129);
nor UO_148 (O_148,N_2963,N_2892);
and UO_149 (O_149,N_2210,N_2676);
and UO_150 (O_150,N_2244,N_2670);
or UO_151 (O_151,N_2799,N_2990);
xnor UO_152 (O_152,N_2253,N_2991);
and UO_153 (O_153,N_2326,N_2110);
nand UO_154 (O_154,N_2831,N_2085);
and UO_155 (O_155,N_2825,N_2526);
nand UO_156 (O_156,N_2711,N_2660);
nor UO_157 (O_157,N_2180,N_2402);
nand UO_158 (O_158,N_2263,N_2393);
or UO_159 (O_159,N_2976,N_2487);
or UO_160 (O_160,N_2524,N_2324);
and UO_161 (O_161,N_2046,N_2173);
nor UO_162 (O_162,N_2183,N_2187);
xnor UO_163 (O_163,N_2143,N_2922);
and UO_164 (O_164,N_2233,N_2975);
nor UO_165 (O_165,N_2682,N_2829);
nor UO_166 (O_166,N_2914,N_2493);
nand UO_167 (O_167,N_2954,N_2107);
and UO_168 (O_168,N_2564,N_2061);
nor UO_169 (O_169,N_2757,N_2274);
nand UO_170 (O_170,N_2344,N_2071);
or UO_171 (O_171,N_2273,N_2981);
or UO_172 (O_172,N_2537,N_2869);
and UO_173 (O_173,N_2580,N_2406);
nor UO_174 (O_174,N_2299,N_2330);
or UO_175 (O_175,N_2989,N_2654);
or UO_176 (O_176,N_2087,N_2895);
nor UO_177 (O_177,N_2258,N_2208);
or UO_178 (O_178,N_2968,N_2126);
xor UO_179 (O_179,N_2064,N_2482);
or UO_180 (O_180,N_2348,N_2125);
and UO_181 (O_181,N_2127,N_2124);
nand UO_182 (O_182,N_2875,N_2221);
and UO_183 (O_183,N_2885,N_2088);
nor UO_184 (O_184,N_2335,N_2800);
xor UO_185 (O_185,N_2456,N_2816);
and UO_186 (O_186,N_2967,N_2671);
nor UO_187 (O_187,N_2673,N_2953);
and UO_188 (O_188,N_2142,N_2894);
and UO_189 (O_189,N_2382,N_2602);
and UO_190 (O_190,N_2791,N_2444);
nor UO_191 (O_191,N_2419,N_2502);
and UO_192 (O_192,N_2469,N_2503);
and UO_193 (O_193,N_2095,N_2839);
nor UO_194 (O_194,N_2649,N_2100);
nand UO_195 (O_195,N_2302,N_2425);
and UO_196 (O_196,N_2473,N_2459);
and UO_197 (O_197,N_2533,N_2153);
and UO_198 (O_198,N_2047,N_2492);
nand UO_199 (O_199,N_2866,N_2507);
and UO_200 (O_200,N_2223,N_2840);
nor UO_201 (O_201,N_2824,N_2957);
nor UO_202 (O_202,N_2771,N_2339);
and UO_203 (O_203,N_2144,N_2958);
nand UO_204 (O_204,N_2518,N_2345);
nand UO_205 (O_205,N_2369,N_2709);
xor UO_206 (O_206,N_2172,N_2235);
nand UO_207 (O_207,N_2569,N_2746);
or UO_208 (O_208,N_2779,N_2248);
or UO_209 (O_209,N_2543,N_2079);
and UO_210 (O_210,N_2514,N_2899);
or UO_211 (O_211,N_2031,N_2319);
and UO_212 (O_212,N_2821,N_2908);
nor UO_213 (O_213,N_2956,N_2702);
nor UO_214 (O_214,N_2341,N_2576);
or UO_215 (O_215,N_2009,N_2647);
xnor UO_216 (O_216,N_2164,N_2435);
nand UO_217 (O_217,N_2707,N_2574);
nand UO_218 (O_218,N_2882,N_2656);
and UO_219 (O_219,N_2266,N_2236);
and UO_220 (O_220,N_2460,N_2050);
nor UO_221 (O_221,N_2777,N_2439);
and UO_222 (O_222,N_2724,N_2936);
nand UO_223 (O_223,N_2925,N_2921);
nor UO_224 (O_224,N_2276,N_2906);
nor UO_225 (O_225,N_2701,N_2007);
nor UO_226 (O_226,N_2872,N_2572);
nand UO_227 (O_227,N_2384,N_2726);
or UO_228 (O_228,N_2383,N_2026);
or UO_229 (O_229,N_2368,N_2199);
or UO_230 (O_230,N_2593,N_2226);
nand UO_231 (O_231,N_2295,N_2232);
nand UO_232 (O_232,N_2612,N_2497);
nand UO_233 (O_233,N_2281,N_2182);
or UO_234 (O_234,N_2561,N_2664);
and UO_235 (O_235,N_2011,N_2655);
nor UO_236 (O_236,N_2437,N_2015);
nand UO_237 (O_237,N_2092,N_2756);
or UO_238 (O_238,N_2025,N_2672);
and UO_239 (O_239,N_2687,N_2774);
or UO_240 (O_240,N_2488,N_2213);
or UO_241 (O_241,N_2651,N_2775);
or UO_242 (O_242,N_2650,N_2202);
nor UO_243 (O_243,N_2860,N_2508);
and UO_244 (O_244,N_2078,N_2845);
nor UO_245 (O_245,N_2357,N_2855);
nand UO_246 (O_246,N_2737,N_2247);
nor UO_247 (O_247,N_2294,N_2847);
nand UO_248 (O_248,N_2310,N_2038);
nand UO_249 (O_249,N_2674,N_2148);
or UO_250 (O_250,N_2045,N_2578);
nor UO_251 (O_251,N_2113,N_2259);
or UO_252 (O_252,N_2787,N_2499);
or UO_253 (O_253,N_2734,N_2801);
or UO_254 (O_254,N_2563,N_2417);
nand UO_255 (O_255,N_2557,N_2462);
and UO_256 (O_256,N_2058,N_2332);
nand UO_257 (O_257,N_2909,N_2688);
nor UO_258 (O_258,N_2404,N_2022);
nor UO_259 (O_259,N_2197,N_2961);
nor UO_260 (O_260,N_2395,N_2804);
nand UO_261 (O_261,N_2764,N_2309);
nor UO_262 (O_262,N_2361,N_2794);
or UO_263 (O_263,N_2093,N_2243);
nor UO_264 (O_264,N_2703,N_2938);
and UO_265 (O_265,N_2191,N_2741);
nor UO_266 (O_266,N_2198,N_2696);
nor UO_267 (O_267,N_2379,N_2848);
nand UO_268 (O_268,N_2887,N_2828);
and UO_269 (O_269,N_2188,N_2933);
nor UO_270 (O_270,N_2619,N_2977);
and UO_271 (O_271,N_2820,N_2171);
and UO_272 (O_272,N_2063,N_2141);
and UO_273 (O_273,N_2668,N_2996);
and UO_274 (O_274,N_2752,N_2161);
or UO_275 (O_275,N_2283,N_2453);
and UO_276 (O_276,N_2581,N_2844);
nand UO_277 (O_277,N_2474,N_2252);
nor UO_278 (O_278,N_2589,N_2336);
or UO_279 (O_279,N_2720,N_2458);
and UO_280 (O_280,N_2074,N_2596);
nor UO_281 (O_281,N_2689,N_2556);
nor UO_282 (O_282,N_2056,N_2878);
xnor UO_283 (O_283,N_2342,N_2445);
and UO_284 (O_284,N_2494,N_2776);
or UO_285 (O_285,N_2728,N_2485);
and UO_286 (O_286,N_2277,N_2108);
nor UO_287 (O_287,N_2396,N_2918);
and UO_288 (O_288,N_2287,N_2789);
or UO_289 (O_289,N_2681,N_2372);
or UO_290 (O_290,N_2811,N_2833);
or UO_291 (O_291,N_2317,N_2356);
nand UO_292 (O_292,N_2224,N_2160);
or UO_293 (O_293,N_2179,N_2731);
or UO_294 (O_294,N_2451,N_2610);
nand UO_295 (O_295,N_2822,N_2511);
and UO_296 (O_296,N_2478,N_2725);
nor UO_297 (O_297,N_2603,N_2910);
nand UO_298 (O_298,N_2408,N_2297);
nand UO_299 (O_299,N_2571,N_2529);
and UO_300 (O_300,N_2251,N_2446);
nor UO_301 (O_301,N_2020,N_2517);
nand UO_302 (O_302,N_2623,N_2853);
and UO_303 (O_303,N_2739,N_2250);
and UO_304 (O_304,N_2156,N_2814);
nor UO_305 (O_305,N_2486,N_2904);
xnor UO_306 (O_306,N_2748,N_2037);
and UO_307 (O_307,N_2611,N_2194);
or UO_308 (O_308,N_2390,N_2377);
or UO_309 (O_309,N_2984,N_2852);
or UO_310 (O_310,N_2325,N_2694);
or UO_311 (O_311,N_2680,N_2652);
nor UO_312 (O_312,N_2823,N_2427);
nand UO_313 (O_313,N_2732,N_2785);
nor UO_314 (O_314,N_2292,N_2405);
nand UO_315 (O_315,N_2836,N_2931);
and UO_316 (O_316,N_2367,N_2858);
nor UO_317 (O_317,N_2640,N_2070);
and UO_318 (O_318,N_2268,N_2762);
and UO_319 (O_319,N_2401,N_2884);
nand UO_320 (O_320,N_2522,N_2949);
nor UO_321 (O_321,N_2298,N_2591);
and UO_322 (O_322,N_2028,N_2362);
nor UO_323 (O_323,N_2573,N_2296);
and UO_324 (O_324,N_2598,N_2176);
nand UO_325 (O_325,N_2366,N_2448);
nor UO_326 (O_326,N_2057,N_2945);
nor UO_327 (O_327,N_2639,N_2052);
and UO_328 (O_328,N_2398,N_2301);
nor UO_329 (O_329,N_2504,N_2599);
nor UO_330 (O_330,N_2780,N_2212);
nand UO_331 (O_331,N_2712,N_2644);
nor UO_332 (O_332,N_2770,N_2371);
nand UO_333 (O_333,N_2115,N_2272);
or UO_334 (O_334,N_2579,N_2407);
xor UO_335 (O_335,N_2722,N_2231);
and UO_336 (O_336,N_2684,N_2484);
and UO_337 (O_337,N_2495,N_2083);
xor UO_338 (O_338,N_2558,N_2912);
nor UO_339 (O_339,N_2457,N_2151);
or UO_340 (O_340,N_2438,N_2588);
and UO_341 (O_341,N_2012,N_2567);
and UO_342 (O_342,N_2060,N_2879);
or UO_343 (O_343,N_2645,N_2841);
and UO_344 (O_344,N_2454,N_2201);
nor UO_345 (O_345,N_2162,N_2049);
and UO_346 (O_346,N_2622,N_2545);
nor UO_347 (O_347,N_2027,N_2763);
and UO_348 (O_348,N_2600,N_2289);
or UO_349 (O_349,N_2769,N_2999);
or UO_350 (O_350,N_2951,N_2304);
and UO_351 (O_351,N_2242,N_2911);
or UO_352 (O_352,N_2467,N_2358);
nor UO_353 (O_353,N_2409,N_2306);
and UO_354 (O_354,N_2311,N_2014);
nor UO_355 (O_355,N_2886,N_2099);
nor UO_356 (O_356,N_2544,N_2089);
nor UO_357 (O_357,N_2630,N_2470);
nor UO_358 (O_358,N_2284,N_2761);
or UO_359 (O_359,N_2323,N_2527);
and UO_360 (O_360,N_2849,N_2979);
nor UO_361 (O_361,N_2033,N_2365);
and UO_362 (O_362,N_2343,N_2175);
and UO_363 (O_363,N_2893,N_2084);
nor UO_364 (O_364,N_2159,N_2924);
nand UO_365 (O_365,N_2846,N_2480);
or UO_366 (O_366,N_2604,N_2819);
or UO_367 (O_367,N_2431,N_2525);
or UO_368 (O_368,N_2416,N_2935);
nor UO_369 (O_369,N_2397,N_2128);
nor UO_370 (O_370,N_2934,N_2184);
nor UO_371 (O_371,N_2386,N_2868);
and UO_372 (O_372,N_2551,N_2932);
or UO_373 (O_373,N_2081,N_2443);
nor UO_374 (O_374,N_2719,N_2678);
and UO_375 (O_375,N_2464,N_2695);
or UO_376 (O_376,N_2616,N_2942);
and UO_377 (O_377,N_2562,N_2806);
nand UO_378 (O_378,N_2986,N_2449);
and UO_379 (O_379,N_2455,N_2308);
or UO_380 (O_380,N_2016,N_2350);
nand UO_381 (O_381,N_2481,N_2859);
nor UO_382 (O_382,N_2705,N_2548);
or UO_383 (O_383,N_2817,N_2838);
or UO_384 (O_384,N_2206,N_2667);
and UO_385 (O_385,N_2723,N_2399);
nand UO_386 (O_386,N_2992,N_2121);
nand UO_387 (O_387,N_2754,N_2132);
or UO_388 (O_388,N_2946,N_2432);
nand UO_389 (O_389,N_2123,N_2120);
or UO_390 (O_390,N_2842,N_2337);
nand UO_391 (O_391,N_2717,N_2692);
and UO_392 (O_392,N_2101,N_2434);
nor UO_393 (O_393,N_2312,N_2515);
or UO_394 (O_394,N_2997,N_2181);
nor UO_395 (O_395,N_2818,N_2928);
nor UO_396 (O_396,N_2966,N_2238);
nor UO_397 (O_397,N_2747,N_2150);
nand UO_398 (O_398,N_2149,N_2387);
nor UO_399 (O_399,N_2721,N_2003);
and UO_400 (O_400,N_2096,N_2597);
or UO_401 (O_401,N_2716,N_2584);
nand UO_402 (O_402,N_2227,N_2498);
or UO_403 (O_403,N_2883,N_2575);
nor UO_404 (O_404,N_2621,N_2962);
or UO_405 (O_405,N_2795,N_2170);
nor UO_406 (O_406,N_2475,N_2512);
and UO_407 (O_407,N_2955,N_2585);
nand UO_408 (O_408,N_2917,N_2536);
or UO_409 (O_409,N_2055,N_2521);
and UO_410 (O_410,N_2929,N_2625);
and UO_411 (O_411,N_2685,N_2952);
nor UO_412 (O_412,N_2528,N_2349);
or UO_413 (O_413,N_2568,N_2256);
and UO_414 (O_414,N_2333,N_2743);
nand UO_415 (O_415,N_2965,N_2559);
nor UO_416 (O_416,N_2465,N_2590);
nand UO_417 (O_417,N_2742,N_2260);
or UO_418 (O_418,N_2381,N_2044);
or UO_419 (O_419,N_2102,N_2270);
and UO_420 (O_420,N_2066,N_2856);
and UO_421 (O_421,N_2927,N_2675);
and UO_422 (O_422,N_2146,N_2073);
nor UO_423 (O_423,N_2147,N_2781);
or UO_424 (O_424,N_2385,N_2767);
nor UO_425 (O_425,N_2043,N_2626);
or UO_426 (O_426,N_2760,N_2843);
nor UO_427 (O_427,N_2903,N_2699);
or UO_428 (O_428,N_2638,N_2004);
nand UO_429 (O_429,N_2661,N_2809);
or UO_430 (O_430,N_2902,N_2577);
nand UO_431 (O_431,N_2587,N_2807);
or UO_432 (O_432,N_2592,N_2267);
and UO_433 (O_433,N_2745,N_2318);
nor UO_434 (O_434,N_2105,N_2403);
or UO_435 (O_435,N_2948,N_2322);
nand UO_436 (O_436,N_2620,N_2540);
or UO_437 (O_437,N_2913,N_2476);
or UO_438 (O_438,N_2075,N_2447);
nand UO_439 (O_439,N_2662,N_2440);
nor UO_440 (O_440,N_2420,N_2916);
nor UO_441 (O_441,N_2959,N_2328);
nor UO_442 (O_442,N_2873,N_2138);
and UO_443 (O_443,N_2850,N_2351);
or UO_444 (O_444,N_2553,N_2628);
and UO_445 (O_445,N_2768,N_2749);
and UO_446 (O_446,N_2477,N_2275);
nand UO_447 (O_447,N_2905,N_2415);
or UO_448 (O_448,N_2782,N_2759);
nor UO_449 (O_449,N_2331,N_2896);
or UO_450 (O_450,N_2271,N_2857);
nand UO_451 (O_451,N_2174,N_2614);
nand UO_452 (O_452,N_2119,N_2069);
nor UO_453 (O_453,N_2713,N_2094);
nor UO_454 (O_454,N_2606,N_2635);
nor UO_455 (O_455,N_2134,N_2496);
or UO_456 (O_456,N_2452,N_2867);
nor UO_457 (O_457,N_2347,N_2062);
nor UO_458 (O_458,N_2566,N_2013);
nor UO_459 (O_459,N_2714,N_2219);
nor UO_460 (O_460,N_2803,N_2648);
and UO_461 (O_461,N_2030,N_2245);
and UO_462 (O_462,N_2735,N_2145);
xnor UO_463 (O_463,N_2029,N_2216);
nor UO_464 (O_464,N_2788,N_2988);
nand UO_465 (O_465,N_2001,N_2155);
nor UO_466 (O_466,N_2225,N_2550);
and UO_467 (O_467,N_2018,N_2740);
and UO_468 (O_468,N_2937,N_2888);
or UO_469 (O_469,N_2051,N_2036);
or UO_470 (O_470,N_2993,N_2116);
and UO_471 (O_471,N_2790,N_2627);
nand UO_472 (O_472,N_2185,N_2429);
and UO_473 (O_473,N_2189,N_2483);
nand UO_474 (O_474,N_2207,N_2501);
or UO_475 (O_475,N_2615,N_2106);
xnor UO_476 (O_476,N_2555,N_2234);
nor UO_477 (O_477,N_2972,N_2068);
nor UO_478 (O_478,N_2519,N_2535);
nand UO_479 (O_479,N_2950,N_2697);
nor UO_480 (O_480,N_2076,N_2827);
and UO_481 (O_481,N_2255,N_2944);
or UO_482 (O_482,N_2547,N_2642);
and UO_483 (O_483,N_2239,N_2436);
nand UO_484 (O_484,N_2363,N_2738);
or UO_485 (O_485,N_2998,N_2812);
nor UO_486 (O_486,N_2861,N_2618);
nand UO_487 (O_487,N_2254,N_2583);
nor UO_488 (O_488,N_2214,N_2468);
nand UO_489 (O_489,N_2375,N_2637);
nor UO_490 (O_490,N_2140,N_2605);
and UO_491 (O_491,N_2538,N_2871);
and UO_492 (O_492,N_2280,N_2617);
nor UO_493 (O_493,N_2389,N_2964);
and UO_494 (O_494,N_2131,N_2278);
nand UO_495 (O_495,N_2472,N_2805);
nor UO_496 (O_496,N_2985,N_2491);
or UO_497 (O_497,N_2380,N_2877);
nor UO_498 (O_498,N_2679,N_2307);
nand UO_499 (O_499,N_2560,N_2098);
endmodule