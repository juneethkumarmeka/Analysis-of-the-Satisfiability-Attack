module basic_1500_15000_2000_30_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_702,In_365);
and U1 (N_1,In_675,In_420);
nor U2 (N_2,In_524,In_1461);
or U3 (N_3,In_509,In_358);
xor U4 (N_4,In_691,In_476);
xor U5 (N_5,In_1373,In_856);
and U6 (N_6,In_1386,In_129);
nor U7 (N_7,In_1284,In_176);
xor U8 (N_8,In_1465,In_1403);
xnor U9 (N_9,In_999,In_439);
nand U10 (N_10,In_525,In_1329);
nand U11 (N_11,In_268,In_271);
nand U12 (N_12,In_514,In_297);
and U13 (N_13,In_1027,In_411);
or U14 (N_14,In_1209,In_535);
nand U15 (N_15,In_577,In_89);
and U16 (N_16,In_1424,In_869);
nand U17 (N_17,In_1071,In_910);
or U18 (N_18,In_208,In_1167);
nand U19 (N_19,In_11,In_804);
xnor U20 (N_20,In_903,In_854);
or U21 (N_21,In_904,In_79);
and U22 (N_22,In_1306,In_622);
and U23 (N_23,In_426,In_292);
or U24 (N_24,In_403,In_1002);
or U25 (N_25,In_1164,In_651);
or U26 (N_26,In_395,In_897);
nand U27 (N_27,In_1222,In_1402);
and U28 (N_28,In_669,In_785);
xor U29 (N_29,In_289,In_1178);
nand U30 (N_30,In_128,In_1250);
nand U31 (N_31,In_922,In_328);
nand U32 (N_32,In_492,In_1150);
nor U33 (N_33,In_991,In_1234);
and U34 (N_34,In_797,In_1253);
nand U35 (N_35,In_687,In_1367);
and U36 (N_36,In_580,In_19);
nand U37 (N_37,In_318,In_1314);
and U38 (N_38,In_1259,In_1126);
xnor U39 (N_39,In_477,In_1088);
nand U40 (N_40,In_878,In_728);
nor U41 (N_41,In_723,In_106);
nor U42 (N_42,In_644,In_1076);
or U43 (N_43,In_346,In_712);
nor U44 (N_44,In_987,In_132);
or U45 (N_45,In_327,In_383);
and U46 (N_46,In_589,In_469);
or U47 (N_47,In_1409,In_655);
xor U48 (N_48,In_2,In_893);
or U49 (N_49,In_938,In_585);
and U50 (N_50,In_473,In_966);
nor U51 (N_51,In_1175,In_1362);
nand U52 (N_52,In_446,In_1184);
xnor U53 (N_53,In_1288,In_902);
or U54 (N_54,In_1374,In_234);
and U55 (N_55,In_1158,In_164);
or U56 (N_56,In_506,In_547);
nor U57 (N_57,In_342,In_1022);
xor U58 (N_58,In_43,In_716);
xor U59 (N_59,In_435,In_778);
or U60 (N_60,In_1108,In_882);
nor U61 (N_61,In_617,In_1012);
nand U62 (N_62,In_1417,In_110);
and U63 (N_63,In_1313,In_627);
and U64 (N_64,In_175,In_13);
and U65 (N_65,In_430,In_850);
nor U66 (N_66,In_1225,In_1220);
nor U67 (N_67,In_737,In_188);
xor U68 (N_68,In_1142,In_360);
and U69 (N_69,In_361,In_9);
and U70 (N_70,In_1464,In_863);
nor U71 (N_71,In_1303,In_1331);
nor U72 (N_72,In_1173,In_422);
xor U73 (N_73,In_145,In_1411);
or U74 (N_74,In_300,In_183);
and U75 (N_75,In_185,In_159);
nor U76 (N_76,In_150,In_369);
nor U77 (N_77,In_925,In_994);
nor U78 (N_78,In_692,In_194);
xnor U79 (N_79,In_248,In_551);
nand U80 (N_80,In_940,In_1065);
nor U81 (N_81,In_400,In_853);
nand U82 (N_82,In_1112,In_1199);
or U83 (N_83,In_359,In_1160);
and U84 (N_84,In_276,In_5);
xnor U85 (N_85,In_385,In_877);
or U86 (N_86,In_490,In_1015);
nand U87 (N_87,In_575,In_1145);
and U88 (N_88,In_275,In_1491);
nand U89 (N_89,In_881,In_1185);
xor U90 (N_90,In_199,In_845);
xor U91 (N_91,In_1020,In_6);
nand U92 (N_92,In_1172,In_1266);
or U93 (N_93,In_206,In_337);
nand U94 (N_94,In_99,In_1192);
nand U95 (N_95,In_1385,In_1177);
or U96 (N_96,In_610,In_769);
and U97 (N_97,In_565,In_70);
and U98 (N_98,In_345,In_1169);
nor U99 (N_99,In_495,In_1423);
or U100 (N_100,In_824,In_351);
xnor U101 (N_101,In_1005,In_173);
nand U102 (N_102,In_834,In_710);
or U103 (N_103,In_419,In_738);
and U104 (N_104,In_852,In_1292);
and U105 (N_105,In_1382,In_388);
or U106 (N_106,In_281,In_660);
nor U107 (N_107,In_623,In_724);
xnor U108 (N_108,In_918,In_67);
nor U109 (N_109,In_170,In_875);
xor U110 (N_110,In_643,In_133);
xnor U111 (N_111,In_1335,In_1033);
and U112 (N_112,In_1154,In_636);
nand U113 (N_113,In_195,In_1193);
nor U114 (N_114,In_1486,In_848);
nand U115 (N_115,In_876,In_1183);
and U116 (N_116,In_215,In_870);
nand U117 (N_117,In_1325,In_463);
nor U118 (N_118,In_325,In_513);
nand U119 (N_119,In_408,In_611);
xnor U120 (N_120,In_1407,In_407);
xor U121 (N_121,In_731,In_331);
nor U122 (N_122,In_387,In_1077);
and U123 (N_123,In_1047,In_304);
and U124 (N_124,In_1000,In_1346);
or U125 (N_125,In_1134,In_621);
xnor U126 (N_126,In_896,In_1141);
nand U127 (N_127,In_568,In_349);
xor U128 (N_128,In_149,In_890);
nor U129 (N_129,In_76,In_354);
nor U130 (N_130,In_1358,In_375);
nand U131 (N_131,In_1434,In_736);
xnor U132 (N_132,In_593,In_650);
nor U133 (N_133,In_972,In_1125);
and U134 (N_134,In_775,In_1073);
nand U135 (N_135,In_1179,In_1355);
nand U136 (N_136,In_1099,In_969);
nor U137 (N_137,In_1147,In_811);
and U138 (N_138,In_25,In_204);
nand U139 (N_139,In_243,In_656);
and U140 (N_140,In_851,In_131);
xnor U141 (N_141,In_900,In_55);
nor U142 (N_142,In_745,In_373);
xnor U143 (N_143,In_190,In_47);
and U144 (N_144,In_1070,In_947);
and U145 (N_145,In_698,In_1489);
and U146 (N_146,In_550,In_1243);
and U147 (N_147,In_117,In_1280);
and U148 (N_148,In_1097,In_51);
xnor U149 (N_149,In_978,In_1232);
xor U150 (N_150,In_1143,In_571);
or U151 (N_151,In_899,In_272);
nand U152 (N_152,In_865,In_293);
xor U153 (N_153,In_1466,In_105);
nand U154 (N_154,In_1347,In_450);
nand U155 (N_155,In_1004,In_631);
nor U156 (N_156,In_127,In_620);
and U157 (N_157,In_122,In_549);
nor U158 (N_158,In_366,In_711);
or U159 (N_159,In_211,In_787);
nor U160 (N_160,In_233,In_86);
nor U161 (N_161,In_116,In_998);
xnor U162 (N_162,In_1315,In_412);
and U163 (N_163,In_258,In_1274);
nor U164 (N_164,In_813,In_1136);
nand U165 (N_165,In_59,In_444);
nand U166 (N_166,In_356,In_1378);
nand U167 (N_167,In_29,In_1404);
or U168 (N_168,In_1282,In_1273);
nor U169 (N_169,In_42,In_1194);
nor U170 (N_170,In_1345,In_988);
nor U171 (N_171,In_36,In_1202);
nand U172 (N_172,In_1216,In_1157);
xnor U173 (N_173,In_227,In_434);
nor U174 (N_174,In_497,In_112);
or U175 (N_175,In_914,In_61);
nand U176 (N_176,In_929,In_511);
nand U177 (N_177,In_313,In_1302);
nand U178 (N_178,In_1035,In_52);
and U179 (N_179,In_168,In_1080);
xor U180 (N_180,In_534,In_570);
or U181 (N_181,In_88,In_1363);
or U182 (N_182,In_406,In_1151);
or U183 (N_183,In_413,In_826);
nor U184 (N_184,In_717,In_371);
and U185 (N_185,In_1051,In_859);
xnor U186 (N_186,In_372,In_729);
or U187 (N_187,In_1389,In_1170);
or U188 (N_188,In_1487,In_567);
and U189 (N_189,In_146,In_100);
or U190 (N_190,In_755,In_703);
nand U191 (N_191,In_1361,In_1233);
xnor U192 (N_192,In_1354,In_144);
nand U193 (N_193,In_809,In_20);
nor U194 (N_194,In_895,In_504);
nor U195 (N_195,In_1296,In_1416);
xnor U196 (N_196,In_517,In_15);
xnor U197 (N_197,In_1421,In_392);
nand U198 (N_198,In_353,In_637);
and U199 (N_199,In_1484,In_202);
nor U200 (N_200,In_143,In_1082);
nor U201 (N_201,In_1351,In_855);
nand U202 (N_202,In_493,In_75);
or U203 (N_203,In_1456,In_254);
and U204 (N_204,In_503,In_44);
nor U205 (N_205,In_1032,In_1387);
nand U206 (N_206,In_125,In_518);
xor U207 (N_207,In_217,In_1072);
nand U208 (N_208,In_618,In_427);
or U209 (N_209,In_1068,In_860);
nand U210 (N_210,In_561,In_955);
nand U211 (N_211,In_66,In_1330);
nor U212 (N_212,In_1471,In_652);
nor U213 (N_213,In_1377,In_1341);
and U214 (N_214,In_1352,In_1226);
nand U215 (N_215,In_46,In_256);
and U216 (N_216,In_884,In_58);
or U217 (N_217,In_908,In_1079);
xor U218 (N_218,In_629,In_382);
nor U219 (N_219,In_722,In_468);
xor U220 (N_220,In_746,In_1120);
nand U221 (N_221,In_1210,In_792);
nor U222 (N_222,In_148,In_1375);
nor U223 (N_223,In_1426,In_1398);
or U224 (N_224,In_213,In_704);
or U225 (N_225,In_399,In_84);
xor U226 (N_226,In_1161,In_798);
nor U227 (N_227,In_71,In_253);
or U228 (N_228,In_730,In_1086);
nor U229 (N_229,In_1023,In_1252);
xor U230 (N_230,In_1492,In_726);
xor U231 (N_231,In_971,In_121);
nor U232 (N_232,In_1153,In_218);
or U233 (N_233,In_1460,In_1241);
and U234 (N_234,In_180,In_941);
nor U235 (N_235,In_1050,In_1269);
or U236 (N_236,In_838,In_321);
nand U237 (N_237,In_814,In_1052);
and U238 (N_238,In_1412,In_1045);
or U239 (N_239,In_1420,In_1208);
xor U240 (N_240,In_662,In_817);
nor U241 (N_241,In_498,In_739);
and U242 (N_242,In_437,In_364);
or U243 (N_243,In_39,In_537);
xor U244 (N_244,In_33,In_1096);
nor U245 (N_245,In_799,In_628);
and U246 (N_246,In_1093,In_1287);
nand U247 (N_247,In_808,In_1422);
or U248 (N_248,In_1436,In_1452);
nand U249 (N_249,In_1413,In_416);
and U250 (N_250,In_515,In_63);
or U251 (N_251,In_224,In_975);
or U252 (N_252,In_680,In_684);
and U253 (N_253,In_749,In_483);
nand U254 (N_254,In_31,In_1174);
xor U255 (N_255,In_1053,In_1083);
or U256 (N_256,In_1181,In_600);
and U257 (N_257,In_807,In_294);
or U258 (N_258,In_480,In_1206);
nand U259 (N_259,In_37,In_1203);
nor U260 (N_260,In_171,In_574);
nor U261 (N_261,In_1334,In_1479);
or U262 (N_262,In_683,In_948);
and U263 (N_263,In_725,In_1454);
and U264 (N_264,In_376,In_788);
xor U265 (N_265,In_378,In_441);
nor U266 (N_266,In_1496,In_138);
nand U267 (N_267,In_10,In_805);
xor U268 (N_268,In_560,In_1327);
and U269 (N_269,In_827,In_639);
and U270 (N_270,In_1455,In_1293);
nand U271 (N_271,In_414,In_136);
and U272 (N_272,In_1283,In_649);
and U273 (N_273,In_1211,In_1443);
and U274 (N_274,In_1391,In_734);
nand U275 (N_275,In_793,In_714);
or U276 (N_276,In_250,In_1488);
xor U277 (N_277,In_699,In_640);
xor U278 (N_278,In_415,In_1030);
nand U279 (N_279,In_1006,In_1074);
and U280 (N_280,In_990,In_1118);
and U281 (N_281,In_576,In_1343);
and U282 (N_282,In_1029,In_840);
nand U283 (N_283,In_829,In_1063);
and U284 (N_284,In_1294,In_220);
and U285 (N_285,In_830,In_1264);
xor U286 (N_286,In_1415,In_678);
nand U287 (N_287,In_1396,In_163);
nor U288 (N_288,In_1224,In_1307);
and U289 (N_289,In_151,In_977);
and U290 (N_290,In_1021,In_315);
xor U291 (N_291,In_73,In_285);
nand U292 (N_292,In_1171,In_979);
xnor U293 (N_293,In_1453,In_613);
nor U294 (N_294,In_847,In_1103);
xor U295 (N_295,In_27,In_210);
or U296 (N_296,In_521,In_16);
nand U297 (N_297,In_754,In_527);
and U298 (N_298,In_1247,In_1235);
or U299 (N_299,In_1430,In_682);
nand U300 (N_300,In_960,In_107);
nor U301 (N_301,In_1446,In_1291);
and U302 (N_302,In_284,In_229);
and U303 (N_303,In_1110,In_1044);
and U304 (N_304,In_40,In_68);
nand U305 (N_305,In_1326,In_0);
nor U306 (N_306,In_1311,In_486);
and U307 (N_307,In_23,In_866);
or U308 (N_308,In_1350,In_1165);
nor U309 (N_309,In_954,In_894);
xor U310 (N_310,In_1001,In_1301);
nand U311 (N_311,In_671,In_310);
nor U312 (N_312,In_1480,In_330);
and U313 (N_313,In_996,In_843);
and U314 (N_314,In_225,In_53);
and U315 (N_315,In_587,In_1248);
nor U316 (N_316,In_543,In_608);
xnor U317 (N_317,In_1467,In_1495);
or U318 (N_318,In_241,In_1449);
xnor U319 (N_319,In_861,In_612);
and U320 (N_320,In_1107,In_937);
xor U321 (N_321,In_7,In_431);
and U322 (N_322,In_926,In_781);
nor U323 (N_323,In_257,In_264);
xor U324 (N_324,In_1379,In_796);
nor U325 (N_325,In_238,In_689);
or U326 (N_326,In_1207,In_1246);
nand U327 (N_327,In_114,In_1217);
and U328 (N_328,In_460,In_1318);
or U329 (N_329,In_1256,In_1039);
xnor U330 (N_330,In_1135,In_1289);
nor U331 (N_331,In_445,In_456);
nor U332 (N_332,In_768,In_1061);
and U333 (N_333,In_928,In_1100);
nand U334 (N_334,In_209,In_464);
xor U335 (N_335,In_1388,In_1268);
and U336 (N_336,In_633,In_26);
nand U337 (N_337,In_436,In_306);
or U338 (N_338,In_449,In_892);
xor U339 (N_339,In_654,In_952);
xor U340 (N_340,In_1046,In_54);
nor U341 (N_341,In_763,In_986);
xnor U342 (N_342,In_590,In_983);
xnor U343 (N_343,In_1010,In_1237);
and U344 (N_344,In_791,In_958);
xnor U345 (N_345,In_849,In_302);
xnor U346 (N_346,In_1419,In_77);
and U347 (N_347,In_1114,In_1137);
and U348 (N_348,In_816,In_533);
and U349 (N_349,In_1109,In_1316);
or U350 (N_350,In_102,In_638);
nand U351 (N_351,In_279,In_765);
nor U352 (N_352,In_1163,In_582);
or U353 (N_353,In_1401,In_605);
nand U354 (N_354,In_667,In_423);
nor U355 (N_355,In_228,In_288);
nor U356 (N_356,In_1337,In_949);
and U357 (N_357,In_507,In_973);
nand U358 (N_358,In_389,In_523);
nor U359 (N_359,In_566,In_1482);
xnor U360 (N_360,In_742,In_786);
nor U361 (N_361,In_822,In_214);
nand U362 (N_362,In_1490,In_461);
or U363 (N_363,In_803,In_1081);
or U364 (N_364,In_1236,In_21);
nand U365 (N_365,In_440,In_812);
nand U366 (N_366,In_1320,In_544);
or U367 (N_367,In_80,In_601);
and U368 (N_368,In_1267,In_65);
and U369 (N_369,In_597,In_453);
nor U370 (N_370,In_1336,In_231);
xnor U371 (N_371,In_794,In_1129);
or U372 (N_372,In_564,In_1095);
or U373 (N_373,In_1117,In_599);
nand U374 (N_374,In_632,In_665);
and U375 (N_375,In_324,In_1049);
xnor U376 (N_376,In_1297,In_705);
nand U377 (N_377,In_178,In_273);
nand U378 (N_378,In_1272,In_1383);
or U379 (N_379,In_197,In_679);
nor U380 (N_380,In_317,In_1007);
nor U381 (N_381,In_959,In_1189);
nor U382 (N_382,In_706,In_278);
nor U383 (N_383,In_614,In_438);
or U384 (N_384,In_1356,In_1498);
or U385 (N_385,In_1428,In_531);
or U386 (N_386,In_24,In_56);
or U387 (N_387,In_748,In_1087);
nand U388 (N_388,In_1384,In_287);
and U389 (N_389,In_62,In_91);
nand U390 (N_390,In_1370,In_980);
and U391 (N_391,In_993,In_1285);
nor U392 (N_392,In_901,In_226);
nor U393 (N_393,In_883,In_642);
xor U394 (N_394,In_124,In_1312);
and U395 (N_395,In_340,In_141);
xor U396 (N_396,In_312,In_484);
nor U397 (N_397,In_90,In_465);
or U398 (N_398,In_69,In_707);
and U399 (N_399,In_964,In_177);
nor U400 (N_400,In_1458,In_474);
xor U401 (N_401,In_1457,In_907);
nor U402 (N_402,In_442,In_556);
and U403 (N_403,In_18,In_761);
nor U404 (N_404,In_835,In_1438);
xor U405 (N_405,In_1043,In_405);
and U406 (N_406,In_995,In_686);
and U407 (N_407,In_283,In_1380);
nor U408 (N_408,In_800,In_1376);
nor U409 (N_409,In_8,In_1214);
xor U410 (N_410,In_887,In_267);
nand U411 (N_411,In_424,In_833);
nand U412 (N_412,In_591,In_237);
xnor U413 (N_413,In_1368,In_539);
nor U414 (N_414,In_1215,In_1102);
or U415 (N_415,In_397,In_740);
or U416 (N_416,In_626,In_1089);
and U417 (N_417,In_223,In_1092);
or U418 (N_418,In_625,In_489);
nor U419 (N_419,In_1405,In_1008);
nor U420 (N_420,In_810,In_1324);
nor U421 (N_421,In_1190,In_48);
nand U422 (N_422,In_1290,In_886);
nor U423 (N_423,In_203,In_596);
and U424 (N_424,In_367,In_108);
nand U425 (N_425,In_488,In_917);
nor U426 (N_426,In_137,In_391);
xor U427 (N_427,In_562,In_1481);
nand U428 (N_428,In_305,In_134);
xor U429 (N_429,In_83,In_485);
nand U430 (N_430,In_192,In_1186);
and U431 (N_431,In_823,In_913);
xor U432 (N_432,In_1144,In_584);
or U433 (N_433,In_572,In_247);
nor U434 (N_434,In_338,In_927);
xnor U435 (N_435,In_261,In_1011);
nor U436 (N_436,In_1156,In_355);
nor U437 (N_437,In_1451,In_997);
or U438 (N_438,In_1255,In_1414);
xor U439 (N_439,In_1124,In_147);
nand U440 (N_440,In_1369,In_579);
and U441 (N_441,In_298,In_789);
xor U442 (N_442,In_759,In_491);
nand U443 (N_443,In_1182,In_1275);
xnor U444 (N_444,In_653,In_207);
xnor U445 (N_445,In_943,In_316);
nand U446 (N_446,In_1249,In_1231);
xnor U447 (N_447,In_1149,In_911);
and U448 (N_448,In_295,In_98);
or U449 (N_449,In_735,In_1475);
nor U450 (N_450,In_118,In_774);
nor U451 (N_451,In_1372,In_1399);
xnor U452 (N_452,In_715,In_874);
or U453 (N_453,In_751,In_1119);
nand U454 (N_454,In_119,In_974);
and U455 (N_455,In_4,In_1198);
xor U456 (N_456,In_274,In_1310);
xor U457 (N_457,In_957,In_1254);
or U458 (N_458,In_992,In_1353);
nor U459 (N_459,In_846,In_433);
or U460 (N_460,In_158,In_255);
or U461 (N_461,In_1016,In_38);
xnor U462 (N_462,In_681,In_50);
and U463 (N_463,In_663,In_1064);
nor U464 (N_464,In_221,In_1339);
nand U465 (N_465,In_909,In_244);
or U466 (N_466,In_239,In_719);
nor U467 (N_467,In_296,In_140);
or U468 (N_468,In_619,In_1060);
nor U469 (N_469,In_624,In_165);
xor U470 (N_470,In_142,In_1101);
nand U471 (N_471,In_1371,In_970);
xnor U472 (N_472,In_953,In_752);
and U473 (N_473,In_1003,In_915);
and U474 (N_474,In_1317,In_520);
or U475 (N_475,In_1094,In_985);
nor U476 (N_476,In_1393,In_45);
or U477 (N_477,In_443,In_428);
nor U478 (N_478,In_377,In_1227);
nand U479 (N_479,In_1017,In_916);
nor U480 (N_480,In_384,In_1058);
nor U481 (N_481,In_693,In_187);
xnor U482 (N_482,In_1239,In_1219);
or U483 (N_483,In_832,In_1483);
nand U484 (N_484,In_828,In_1328);
and U485 (N_485,In_783,In_676);
nor U486 (N_486,In_429,In_658);
nor U487 (N_487,In_806,In_396);
xor U488 (N_488,In_1340,In_1104);
nand U489 (N_489,In_1308,In_459);
and U490 (N_490,In_697,In_981);
or U491 (N_491,In_472,In_139);
or U492 (N_492,In_1359,In_1036);
and U493 (N_493,In_516,In_266);
and U494 (N_494,In_1286,In_688);
xnor U495 (N_495,In_1084,In_868);
xor U496 (N_496,In_242,In_1195);
nor U497 (N_497,In_604,In_81);
xnor U498 (N_498,In_402,In_198);
and U499 (N_499,In_155,In_205);
nor U500 (N_500,N_400,In_169);
or U501 (N_501,In_1240,In_819);
xor U502 (N_502,N_487,N_118);
xor U503 (N_503,N_254,N_458);
nor U504 (N_504,In_961,In_418);
xor U505 (N_505,In_1470,N_170);
and U506 (N_506,N_143,N_359);
and U507 (N_507,In_1091,N_307);
nor U508 (N_508,N_353,N_75);
nand U509 (N_509,N_134,In_475);
xnor U510 (N_510,In_762,N_102);
or U511 (N_511,In_1121,N_59);
nand U512 (N_512,In_363,N_288);
xor U513 (N_513,In_594,N_408);
or U514 (N_514,In_1342,In_93);
nor U515 (N_515,In_270,N_220);
nand U516 (N_516,In_573,N_135);
xor U517 (N_517,In_347,In_528);
nor U518 (N_518,In_1201,In_401);
nor U519 (N_519,N_96,N_127);
nor U520 (N_520,N_491,In_326);
or U521 (N_521,N_426,N_464);
nor U522 (N_522,In_499,In_1477);
or U523 (N_523,N_200,In_989);
or U524 (N_524,N_105,In_744);
nor U525 (N_525,N_66,In_303);
nor U526 (N_526,N_15,In_481);
and U527 (N_527,In_417,In_380);
or U528 (N_528,In_530,In_196);
nor U529 (N_529,N_334,In_932);
and U530 (N_530,In_1078,In_501);
and U531 (N_531,In_747,In_269);
nor U532 (N_532,In_12,In_1066);
and U533 (N_533,N_492,In_670);
or U534 (N_534,In_542,In_545);
nand U535 (N_535,N_76,N_296);
or U536 (N_536,In_1271,N_14);
nor U537 (N_537,N_237,In_641);
or U538 (N_538,In_837,N_452);
nand U539 (N_539,In_1166,In_1055);
or U540 (N_540,N_277,N_498);
nand U541 (N_541,N_215,N_56);
and U542 (N_542,In_592,In_944);
nand U543 (N_543,In_1418,In_448);
nor U544 (N_544,N_247,N_19);
nor U545 (N_545,N_301,N_283);
nand U546 (N_546,N_138,N_490);
nor U547 (N_547,In_1067,In_646);
and U548 (N_548,N_425,In_286);
xnor U549 (N_549,N_146,N_238);
or U550 (N_550,N_499,N_295);
or U551 (N_551,N_291,N_279);
xnor U552 (N_552,N_412,In_339);
nor U553 (N_553,N_258,N_304);
and U554 (N_554,N_465,N_354);
and U555 (N_555,In_1013,In_344);
and U556 (N_556,N_202,N_483);
or U557 (N_557,N_12,In_1196);
nand U558 (N_558,In_1360,N_114);
or U559 (N_559,In_35,In_708);
and U560 (N_560,In_404,In_889);
xnor U561 (N_561,N_191,In_323);
or U562 (N_562,N_207,N_375);
nor U563 (N_563,In_1260,In_1218);
nand U564 (N_564,In_802,N_453);
or U565 (N_565,N_350,N_415);
or U566 (N_566,N_183,In_496);
nor U567 (N_567,N_182,In_529);
xnor U568 (N_568,In_569,N_24);
or U569 (N_569,In_532,N_124);
or U570 (N_570,N_228,In_1349);
nor U571 (N_571,N_16,N_206);
nor U572 (N_572,In_332,In_49);
nor U573 (N_573,N_461,N_449);
and U574 (N_574,In_767,N_298);
nand U575 (N_575,In_771,N_351);
nor U576 (N_576,In_1123,N_136);
xor U577 (N_577,N_367,In_152);
and U578 (N_578,N_115,N_317);
nor U579 (N_579,In_1494,In_880);
xor U580 (N_580,N_339,In_713);
or U581 (N_581,N_193,N_406);
or U582 (N_582,In_290,In_635);
xor U583 (N_583,In_603,N_72);
nand U584 (N_584,N_28,In_968);
nand U585 (N_585,N_213,In_82);
nand U586 (N_586,N_368,In_334);
and U587 (N_587,N_119,In_588);
nor U588 (N_588,N_180,In_216);
nor U589 (N_589,In_1300,In_17);
nand U590 (N_590,In_1159,In_200);
nand U591 (N_591,N_171,N_274);
and U592 (N_592,In_458,In_240);
and U593 (N_593,N_436,N_417);
or U594 (N_594,N_432,N_323);
nand U595 (N_595,N_306,N_83);
nor U596 (N_596,In_1298,In_779);
xnor U597 (N_597,In_750,In_130);
nand U598 (N_598,In_457,In_554);
or U599 (N_599,N_451,In_172);
or U600 (N_600,In_92,N_244);
nand U601 (N_601,In_1244,N_35);
and U602 (N_602,N_418,In_1447);
or U603 (N_603,N_107,In_1348);
and U604 (N_604,In_1,N_370);
xor U605 (N_605,In_1155,In_425);
nand U606 (N_606,In_844,In_984);
or U607 (N_607,N_260,In_607);
nand U608 (N_608,N_489,N_2);
and U609 (N_609,In_1057,In_1392);
and U610 (N_610,In_1439,N_360);
and U611 (N_611,In_1221,In_906);
xnor U612 (N_612,N_89,N_176);
or U613 (N_613,In_606,N_294);
xnor U614 (N_614,In_784,N_148);
xor U615 (N_615,In_30,N_303);
xnor U616 (N_616,In_1168,In_236);
or U617 (N_617,N_91,In_410);
and U618 (N_618,N_239,In_1034);
or U619 (N_619,In_951,In_666);
nand U620 (N_620,In_78,In_1026);
and U621 (N_621,N_497,N_164);
and U622 (N_622,N_71,In_432);
xor U623 (N_623,N_356,In_482);
nor U624 (N_624,In_942,In_362);
xor U625 (N_625,N_431,In_756);
nor U626 (N_626,In_609,In_873);
xnor U627 (N_627,In_478,In_1429);
nor U628 (N_628,N_427,N_233);
nor U629 (N_629,In_1322,In_1162);
nand U630 (N_630,N_256,In_578);
and U631 (N_631,In_976,In_1146);
xnor U632 (N_632,N_199,In_753);
and U633 (N_633,N_478,N_371);
and U634 (N_634,N_44,N_476);
nand U635 (N_635,In_1180,N_217);
and U636 (N_636,N_302,In_1111);
and U637 (N_637,N_190,N_411);
nand U638 (N_638,N_99,N_30);
xnor U639 (N_639,In_885,In_154);
and U640 (N_640,In_598,In_28);
nand U641 (N_641,N_34,In_1040);
or U642 (N_642,N_420,In_508);
and U643 (N_643,N_313,N_225);
nand U644 (N_644,In_1140,In_1344);
nor U645 (N_645,In_777,N_398);
nor U646 (N_646,In_709,In_581);
nand U647 (N_647,N_227,N_284);
nor U648 (N_648,In_764,In_1056);
and U649 (N_649,In_1019,N_343);
nand U650 (N_650,N_29,In_1400);
xnor U651 (N_651,In_668,N_162);
nand U652 (N_652,In_352,In_946);
nor U653 (N_653,In_648,In_162);
nor U654 (N_654,N_116,In_1469);
xor U655 (N_655,In_3,N_401);
and U656 (N_656,N_23,N_457);
nand U657 (N_657,N_63,In_546);
and U658 (N_658,In_60,N_468);
xor U659 (N_659,N_242,In_879);
nand U660 (N_660,N_333,N_329);
nand U661 (N_661,N_315,N_93);
nor U662 (N_662,In_370,In_602);
and U663 (N_663,In_780,N_396);
or U664 (N_664,In_277,N_322);
nand U665 (N_665,N_479,In_1200);
nor U666 (N_666,N_152,N_149);
and U667 (N_667,N_173,In_1213);
nor U668 (N_668,In_394,In_212);
nand U669 (N_669,In_872,In_1261);
and U670 (N_670,In_1463,In_72);
nand U671 (N_671,N_108,In_191);
nand U672 (N_672,N_42,N_495);
nand U673 (N_673,N_330,In_1018);
nor U674 (N_674,In_695,N_161);
nand U675 (N_675,In_1238,N_210);
nand U676 (N_676,N_160,N_234);
xor U677 (N_677,In_487,In_522);
and U678 (N_678,N_224,In_96);
nor U679 (N_679,In_891,In_1075);
and U680 (N_680,N_297,N_221);
xor U681 (N_681,N_157,In_282);
nand U682 (N_682,In_1277,N_265);
or U683 (N_683,In_1042,N_25);
and U684 (N_684,N_20,N_209);
and U685 (N_685,N_399,N_447);
and U686 (N_686,N_130,N_455);
and U687 (N_687,In_1395,In_1176);
or U688 (N_688,N_179,In_109);
and U689 (N_689,In_181,In_1132);
or U690 (N_690,In_1437,N_230);
nor U691 (N_691,In_757,N_106);
xor U692 (N_692,In_1191,In_1257);
nor U693 (N_693,N_235,In_825);
and U694 (N_694,N_214,In_502);
nor U695 (N_695,In_1427,In_479);
or U696 (N_696,In_1037,N_270);
nand U697 (N_697,N_169,N_163);
nand U698 (N_698,In_1299,N_397);
nand U699 (N_699,N_268,N_141);
nor U700 (N_700,In_343,In_1188);
or U701 (N_701,In_97,N_204);
nor U702 (N_702,In_758,N_462);
nand U703 (N_703,N_208,N_459);
xor U704 (N_704,In_368,In_1251);
xor U705 (N_705,N_300,In_1048);
nand U706 (N_706,N_477,N_249);
and U707 (N_707,N_413,In_694);
or U708 (N_708,In_320,In_661);
xnor U709 (N_709,N_448,N_36);
or U710 (N_710,In_923,N_95);
nand U711 (N_711,In_1445,N_186);
or U712 (N_712,N_10,N_101);
or U713 (N_713,In_454,In_184);
nor U714 (N_714,In_14,In_1139);
nand U715 (N_715,In_1054,N_113);
nor U716 (N_716,N_430,N_154);
and U717 (N_717,In_409,N_262);
xor U718 (N_718,In_557,N_203);
xor U719 (N_719,In_1265,In_309);
or U720 (N_720,In_1262,N_494);
nor U721 (N_721,N_111,N_50);
nand U722 (N_722,In_1212,N_345);
and U723 (N_723,In_905,In_659);
or U724 (N_724,N_441,N_17);
or U725 (N_725,N_31,N_391);
xor U726 (N_726,In_1304,N_43);
and U727 (N_727,In_1090,N_81);
or U728 (N_728,N_328,N_97);
nand U729 (N_729,N_13,N_358);
xor U730 (N_730,In_235,In_950);
nor U731 (N_731,In_1365,In_930);
and U732 (N_732,N_85,N_65);
nand U733 (N_733,N_198,In_512);
nand U734 (N_734,In_864,N_424);
xor U735 (N_735,N_364,N_67);
nor U736 (N_736,N_305,In_262);
nand U737 (N_737,In_1009,N_439);
xnor U738 (N_738,In_540,N_442);
or U739 (N_739,N_48,In_1038);
nand U740 (N_740,In_1106,In_308);
xnor U741 (N_741,N_485,N_327);
xor U742 (N_742,N_421,In_157);
nor U743 (N_743,In_350,In_1440);
and U744 (N_744,In_935,N_311);
or U745 (N_745,In_1131,In_393);
nand U746 (N_746,In_732,In_1450);
and U747 (N_747,N_137,In_1127);
xnor U748 (N_748,N_445,N_471);
nor U749 (N_749,N_147,In_842);
nor U750 (N_750,N_54,In_967);
nand U751 (N_751,N_484,In_1408);
nand U752 (N_752,N_21,In_120);
nor U753 (N_753,In_1130,N_145);
and U754 (N_754,N_61,In_280);
and U755 (N_755,N_4,In_1223);
or U756 (N_756,In_167,In_645);
xor U757 (N_757,N_201,In_963);
nor U758 (N_758,In_519,In_1410);
or U759 (N_759,N_325,N_379);
xnor U760 (N_760,N_251,In_790);
nand U761 (N_761,In_664,In_690);
nor U762 (N_762,In_945,In_696);
xor U763 (N_763,In_795,In_772);
and U764 (N_764,In_727,N_77);
nor U765 (N_765,N_128,N_338);
nor U766 (N_766,N_87,N_45);
nor U767 (N_767,N_150,N_444);
and U768 (N_768,In_956,N_267);
xor U769 (N_769,In_57,In_1441);
or U770 (N_770,In_526,N_32);
xor U771 (N_771,In_87,In_505);
and U772 (N_772,N_433,N_275);
and U773 (N_773,In_398,In_815);
nor U774 (N_774,In_563,N_434);
nor U775 (N_775,N_126,In_1497);
xor U776 (N_776,In_1459,In_818);
or U777 (N_777,N_429,In_329);
or U778 (N_778,In_1270,N_355);
xnor U779 (N_779,In_455,N_222);
and U780 (N_780,In_115,In_1406);
xnor U781 (N_781,In_1323,In_553);
xnor U782 (N_782,N_409,N_51);
and U783 (N_783,In_201,N_6);
nor U784 (N_784,N_131,In_101);
xor U785 (N_785,N_419,N_142);
and U786 (N_786,N_156,N_374);
and U787 (N_787,N_273,In_857);
nand U788 (N_788,In_103,In_1476);
nand U789 (N_789,In_1138,N_46);
nor U790 (N_790,N_414,N_80);
and U791 (N_791,N_469,In_160);
or U792 (N_792,In_672,In_1397);
nand U793 (N_793,N_5,In_558);
xor U794 (N_794,N_272,In_307);
or U795 (N_795,In_1321,N_276);
nor U796 (N_796,In_831,N_37);
or U797 (N_797,In_898,N_39);
nor U798 (N_798,N_122,In_219);
xnor U799 (N_799,In_471,In_921);
or U800 (N_800,In_1105,N_92);
nor U801 (N_801,N_292,N_446);
nand U802 (N_802,In_1228,N_88);
xor U803 (N_803,N_9,In_1113);
xnor U804 (N_804,N_403,In_1279);
nand U805 (N_805,N_178,N_181);
or U806 (N_806,In_452,N_211);
xor U807 (N_807,In_1128,N_416);
or U808 (N_808,N_454,In_1187);
xnor U809 (N_809,N_310,In_1278);
or U810 (N_810,N_280,In_867);
xnor U811 (N_811,N_389,In_1364);
nand U812 (N_812,N_123,N_312);
xnor U813 (N_813,N_383,N_187);
nand U814 (N_814,N_98,In_770);
xnor U815 (N_815,In_595,In_559);
xor U816 (N_816,In_1116,In_1041);
and U817 (N_817,N_361,N_68);
nor U818 (N_818,In_246,In_322);
or U819 (N_819,N_331,N_365);
nand U820 (N_820,N_188,N_486);
and U821 (N_821,In_841,N_259);
xor U822 (N_822,N_287,In_1338);
nor U823 (N_823,N_269,In_1152);
xor U824 (N_824,N_404,N_49);
and U825 (N_825,N_70,In_741);
or U826 (N_826,N_440,N_53);
nor U827 (N_827,N_229,N_335);
and U828 (N_828,In_912,In_1473);
nand U829 (N_829,N_481,In_379);
xor U830 (N_830,N_373,N_405);
nor U831 (N_831,In_1478,In_263);
or U832 (N_832,In_1357,In_462);
nor U833 (N_833,In_936,In_161);
or U834 (N_834,N_27,N_382);
and U835 (N_835,N_264,In_1242);
or U836 (N_836,N_112,In_701);
and U837 (N_837,N_324,In_1493);
and U838 (N_838,N_52,N_363);
or U839 (N_839,N_344,N_393);
xor U840 (N_840,In_674,N_316);
xor U841 (N_841,In_74,In_390);
or U842 (N_842,In_466,In_743);
and U843 (N_843,In_1366,In_630);
xnor U844 (N_844,In_336,In_1031);
nand U845 (N_845,In_189,In_616);
and U846 (N_846,In_773,N_40);
xnor U847 (N_847,N_437,N_473);
nand U848 (N_848,N_381,In_348);
nor U849 (N_849,N_320,N_384);
nor U850 (N_850,N_226,In_179);
nand U851 (N_851,N_336,N_347);
xnor U852 (N_852,In_249,N_94);
and U853 (N_853,In_291,In_776);
nand U854 (N_854,In_1433,In_470);
nor U855 (N_855,N_271,N_319);
nand U856 (N_856,In_1197,N_8);
nand U857 (N_857,N_410,N_496);
and U858 (N_858,In_1444,N_460);
and U859 (N_859,In_583,In_319);
or U860 (N_860,N_321,In_839);
xor U861 (N_861,N_69,N_349);
nor U862 (N_862,In_41,N_62);
nand U863 (N_863,In_720,In_1381);
xor U864 (N_864,In_153,N_480);
nand U865 (N_865,N_282,In_451);
nor U866 (N_866,N_192,In_500);
or U867 (N_867,N_165,In_919);
xnor U868 (N_868,In_447,N_174);
nor U869 (N_869,In_1148,In_924);
nand U870 (N_870,N_392,In_801);
or U871 (N_871,N_443,N_26);
or U872 (N_872,In_1085,In_314);
xor U873 (N_873,In_1122,In_386);
nand U874 (N_874,In_1435,In_333);
nor U875 (N_875,N_195,In_1062);
or U876 (N_876,N_475,N_248);
nor U877 (N_877,N_352,In_1425);
nor U878 (N_878,In_615,N_423);
xnor U879 (N_879,In_335,N_231);
or U880 (N_880,In_821,In_1390);
xnor U881 (N_881,N_388,In_94);
nor U882 (N_882,N_140,In_555);
nor U883 (N_883,N_407,In_113);
nor U884 (N_884,N_309,In_156);
nand U885 (N_885,In_934,N_332);
and U886 (N_886,In_421,N_395);
nor U887 (N_887,N_185,N_177);
xor U888 (N_888,N_348,In_182);
or U889 (N_889,In_1115,N_155);
xnor U890 (N_890,In_341,N_467);
nor U891 (N_891,N_120,N_218);
nor U892 (N_892,N_263,N_278);
or U893 (N_893,N_73,N_194);
and U894 (N_894,In_836,In_1432);
nor U895 (N_895,N_385,In_32);
and U896 (N_896,In_920,In_700);
xnor U897 (N_897,N_33,N_246);
nand U898 (N_898,In_962,In_858);
and U899 (N_899,N_470,N_103);
xor U900 (N_900,N_47,In_1468);
xor U901 (N_901,In_862,N_281);
xnor U902 (N_902,In_1448,In_381);
nand U903 (N_903,In_251,N_257);
or U904 (N_904,In_166,In_982);
nand U905 (N_905,In_1442,In_252);
nor U906 (N_906,In_673,N_144);
nand U907 (N_907,In_174,N_175);
and U908 (N_908,N_241,N_121);
nand U909 (N_909,N_232,N_380);
and U910 (N_910,N_18,N_450);
xnor U911 (N_911,N_318,In_685);
and U912 (N_912,N_377,N_466);
xnor U913 (N_913,In_95,N_11);
nor U914 (N_914,N_285,N_255);
nor U915 (N_915,In_1230,N_261);
and U916 (N_916,N_196,In_22);
and U917 (N_917,N_159,In_1474);
nor U918 (N_918,In_299,N_57);
or U919 (N_919,N_125,In_1332);
and U920 (N_920,In_1472,In_104);
or U921 (N_921,In_135,N_493);
nand U922 (N_922,N_402,N_286);
nand U923 (N_923,N_197,In_232);
xnor U924 (N_924,N_435,N_341);
nand U925 (N_925,N_100,N_438);
or U926 (N_926,In_647,N_266);
or U927 (N_927,N_153,In_1333);
xor U928 (N_928,In_357,N_172);
or U929 (N_929,In_1025,In_721);
xor U930 (N_930,N_133,In_1245);
xnor U931 (N_931,In_245,N_166);
or U932 (N_932,In_766,N_212);
xnor U933 (N_933,N_236,N_205);
nand U934 (N_934,In_939,In_186);
or U935 (N_935,N_378,N_151);
or U936 (N_936,N_372,N_79);
or U937 (N_937,In_1394,N_290);
and U938 (N_938,N_387,In_552);
nand U939 (N_939,In_510,In_1258);
nand U940 (N_940,N_129,N_41);
nor U941 (N_941,In_1499,In_260);
or U942 (N_942,In_1024,In_1069);
or U943 (N_943,N_1,N_110);
nor U944 (N_944,In_193,In_34);
or U945 (N_945,N_22,In_311);
or U946 (N_946,In_634,N_472);
nand U947 (N_947,N_340,N_369);
or U948 (N_948,In_230,In_1014);
nand U949 (N_949,N_456,In_677);
xnor U950 (N_950,In_718,N_184);
and U951 (N_951,In_126,In_374);
xnor U952 (N_952,In_933,In_1319);
nor U953 (N_953,N_482,N_84);
or U954 (N_954,In_1305,In_265);
xor U955 (N_955,N_289,N_223);
and U956 (N_956,N_314,In_1133);
nand U957 (N_957,N_104,In_494);
or U958 (N_958,In_1462,N_366);
nor U959 (N_959,N_463,In_733);
xnor U960 (N_960,N_253,In_541);
nand U961 (N_961,N_386,N_428);
nor U962 (N_962,In_1485,N_167);
and U963 (N_963,In_1276,In_1295);
xor U964 (N_964,N_58,In_301);
and U965 (N_965,N_337,N_240);
or U966 (N_966,N_74,N_376);
nor U967 (N_967,N_250,In_85);
nand U968 (N_968,N_243,In_760);
and U969 (N_969,N_422,N_326);
or U970 (N_970,In_657,N_299);
nand U971 (N_971,N_390,N_189);
and U972 (N_972,In_538,In_1229);
xor U973 (N_973,In_111,N_139);
nor U974 (N_974,N_158,N_64);
and U975 (N_975,In_888,In_259);
xnor U976 (N_976,In_536,In_1205);
nand U977 (N_977,In_1263,In_1098);
or U978 (N_978,N_117,In_548);
nor U979 (N_979,In_1309,N_219);
and U980 (N_980,In_467,N_346);
xor U981 (N_981,In_64,In_820);
or U982 (N_982,N_55,N_78);
nand U983 (N_983,In_1431,N_90);
nand U984 (N_984,N_0,N_86);
nor U985 (N_985,N_3,In_1204);
nand U986 (N_986,N_245,N_109);
nor U987 (N_987,In_965,N_7);
xor U988 (N_988,N_293,N_342);
and U989 (N_989,N_308,In_871);
and U990 (N_990,In_586,N_394);
nor U991 (N_991,N_82,N_474);
and U992 (N_992,In_1059,In_782);
nor U993 (N_993,N_488,N_132);
and U994 (N_994,N_38,N_362);
and U995 (N_995,N_60,In_931);
or U996 (N_996,In_222,N_216);
and U997 (N_997,N_252,In_123);
xor U998 (N_998,N_357,N_168);
xor U999 (N_999,In_1281,In_1028);
or U1000 (N_1000,N_913,N_939);
and U1001 (N_1001,N_567,N_729);
or U1002 (N_1002,N_536,N_970);
and U1003 (N_1003,N_807,N_901);
nand U1004 (N_1004,N_915,N_507);
xnor U1005 (N_1005,N_920,N_515);
or U1006 (N_1006,N_821,N_767);
nor U1007 (N_1007,N_831,N_693);
and U1008 (N_1008,N_513,N_545);
or U1009 (N_1009,N_849,N_846);
nor U1010 (N_1010,N_618,N_699);
nand U1011 (N_1011,N_940,N_591);
or U1012 (N_1012,N_617,N_832);
nand U1013 (N_1013,N_654,N_739);
nor U1014 (N_1014,N_630,N_575);
nand U1015 (N_1015,N_525,N_780);
or U1016 (N_1016,N_876,N_741);
and U1017 (N_1017,N_889,N_855);
nor U1018 (N_1018,N_822,N_932);
nor U1019 (N_1019,N_823,N_927);
nand U1020 (N_1020,N_647,N_596);
and U1021 (N_1021,N_713,N_895);
xnor U1022 (N_1022,N_590,N_706);
and U1023 (N_1023,N_884,N_563);
nand U1024 (N_1024,N_830,N_973);
nor U1025 (N_1025,N_806,N_829);
nand U1026 (N_1026,N_828,N_540);
or U1027 (N_1027,N_526,N_725);
nor U1028 (N_1028,N_658,N_599);
or U1029 (N_1029,N_752,N_714);
xor U1030 (N_1030,N_888,N_809);
and U1031 (N_1031,N_632,N_665);
nand U1032 (N_1032,N_577,N_985);
or U1033 (N_1033,N_698,N_730);
and U1034 (N_1034,N_711,N_580);
nand U1035 (N_1035,N_709,N_892);
xor U1036 (N_1036,N_673,N_523);
xor U1037 (N_1037,N_687,N_695);
xnor U1038 (N_1038,N_535,N_847);
xor U1039 (N_1039,N_502,N_933);
and U1040 (N_1040,N_505,N_508);
xnor U1041 (N_1041,N_878,N_848);
xnor U1042 (N_1042,N_655,N_863);
and U1043 (N_1043,N_597,N_980);
or U1044 (N_1044,N_799,N_668);
or U1045 (N_1045,N_923,N_842);
nand U1046 (N_1046,N_872,N_975);
or U1047 (N_1047,N_773,N_991);
nor U1048 (N_1048,N_858,N_735);
and U1049 (N_1049,N_688,N_760);
nor U1050 (N_1050,N_528,N_541);
and U1051 (N_1051,N_899,N_659);
or U1052 (N_1052,N_601,N_820);
and U1053 (N_1053,N_734,N_917);
nor U1054 (N_1054,N_790,N_782);
xnor U1055 (N_1055,N_983,N_835);
xor U1056 (N_1056,N_969,N_750);
or U1057 (N_1057,N_690,N_845);
xor U1058 (N_1058,N_839,N_979);
xnor U1059 (N_1059,N_623,N_615);
nor U1060 (N_1060,N_958,N_930);
nor U1061 (N_1061,N_624,N_784);
or U1062 (N_1062,N_906,N_569);
or U1063 (N_1063,N_724,N_747);
or U1064 (N_1064,N_988,N_501);
xnor U1065 (N_1065,N_961,N_742);
xor U1066 (N_1066,N_804,N_873);
nand U1067 (N_1067,N_953,N_573);
nor U1068 (N_1068,N_946,N_818);
nand U1069 (N_1069,N_914,N_753);
nand U1070 (N_1070,N_891,N_907);
nor U1071 (N_1071,N_707,N_902);
nor U1072 (N_1072,N_783,N_534);
and U1073 (N_1073,N_910,N_531);
nor U1074 (N_1074,N_594,N_749);
or U1075 (N_1075,N_826,N_954);
or U1076 (N_1076,N_613,N_656);
or U1077 (N_1077,N_748,N_585);
nor U1078 (N_1078,N_982,N_755);
nor U1079 (N_1079,N_827,N_527);
and U1080 (N_1080,N_797,N_789);
xnor U1081 (N_1081,N_674,N_637);
nand U1082 (N_1082,N_894,N_696);
nand U1083 (N_1083,N_675,N_893);
nor U1084 (N_1084,N_628,N_791);
and U1085 (N_1085,N_678,N_887);
or U1086 (N_1086,N_683,N_705);
nand U1087 (N_1087,N_704,N_861);
and U1088 (N_1088,N_517,N_712);
and U1089 (N_1089,N_986,N_571);
or U1090 (N_1090,N_824,N_918);
xor U1091 (N_1091,N_518,N_838);
nand U1092 (N_1092,N_745,N_777);
nand U1093 (N_1093,N_833,N_864);
or U1094 (N_1094,N_609,N_542);
xnor U1095 (N_1095,N_560,N_813);
and U1096 (N_1096,N_589,N_511);
or U1097 (N_1097,N_661,N_795);
and U1098 (N_1098,N_948,N_756);
xor U1099 (N_1099,N_786,N_717);
or U1100 (N_1100,N_552,N_625);
and U1101 (N_1101,N_633,N_787);
nand U1102 (N_1102,N_976,N_532);
or U1103 (N_1103,N_544,N_740);
or U1104 (N_1104,N_556,N_619);
or U1105 (N_1105,N_869,N_880);
nor U1106 (N_1106,N_916,N_667);
or U1107 (N_1107,N_595,N_557);
nor U1108 (N_1108,N_775,N_865);
nand U1109 (N_1109,N_691,N_928);
nand U1110 (N_1110,N_792,N_905);
nand U1111 (N_1111,N_997,N_978);
and U1112 (N_1112,N_931,N_757);
nor U1113 (N_1113,N_904,N_924);
nor U1114 (N_1114,N_934,N_620);
nor U1115 (N_1115,N_751,N_680);
nand U1116 (N_1116,N_952,N_937);
nor U1117 (N_1117,N_945,N_641);
nand U1118 (N_1118,N_605,N_614);
nor U1119 (N_1119,N_771,N_957);
nand U1120 (N_1120,N_972,N_685);
xor U1121 (N_1121,N_631,N_785);
nor U1122 (N_1122,N_852,N_660);
xnor U1123 (N_1123,N_684,N_758);
nor U1124 (N_1124,N_722,N_581);
nand U1125 (N_1125,N_836,N_759);
and U1126 (N_1126,N_627,N_938);
or U1127 (N_1127,N_859,N_692);
nor U1128 (N_1128,N_516,N_801);
xor U1129 (N_1129,N_761,N_744);
and U1130 (N_1130,N_561,N_862);
or U1131 (N_1131,N_732,N_837);
xor U1132 (N_1132,N_943,N_768);
and U1133 (N_1133,N_682,N_681);
and U1134 (N_1134,N_956,N_593);
xor U1135 (N_1135,N_676,N_564);
nand U1136 (N_1136,N_964,N_817);
nor U1137 (N_1137,N_908,N_548);
nand U1138 (N_1138,N_506,N_524);
xnor U1139 (N_1139,N_576,N_586);
nand U1140 (N_1140,N_960,N_935);
and U1141 (N_1141,N_968,N_951);
nor U1142 (N_1142,N_689,N_606);
nor U1143 (N_1143,N_922,N_881);
xor U1144 (N_1144,N_950,N_570);
and U1145 (N_1145,N_521,N_883);
nand U1146 (N_1146,N_999,N_736);
nor U1147 (N_1147,N_640,N_959);
or U1148 (N_1148,N_981,N_592);
nor U1149 (N_1149,N_866,N_860);
and U1150 (N_1150,N_720,N_737);
xor U1151 (N_1151,N_582,N_875);
xor U1152 (N_1152,N_886,N_686);
nand U1153 (N_1153,N_811,N_700);
nand U1154 (N_1154,N_921,N_778);
nor U1155 (N_1155,N_776,N_697);
nor U1156 (N_1156,N_514,N_583);
nor U1157 (N_1157,N_549,N_764);
nor U1158 (N_1158,N_509,N_947);
xor U1159 (N_1159,N_805,N_984);
nor U1160 (N_1160,N_537,N_612);
nand U1161 (N_1161,N_559,N_844);
nor U1162 (N_1162,N_798,N_634);
and U1163 (N_1163,N_635,N_942);
xnor U1164 (N_1164,N_611,N_772);
nor U1165 (N_1165,N_879,N_510);
nand U1166 (N_1166,N_616,N_834);
or U1167 (N_1167,N_648,N_754);
xnor U1168 (N_1168,N_912,N_642);
nand U1169 (N_1169,N_738,N_679);
xor U1170 (N_1170,N_971,N_562);
or U1171 (N_1171,N_529,N_566);
or U1172 (N_1172,N_520,N_638);
xnor U1173 (N_1173,N_963,N_565);
xor U1174 (N_1174,N_998,N_603);
xnor U1175 (N_1175,N_766,N_578);
or U1176 (N_1176,N_825,N_649);
xor U1177 (N_1177,N_547,N_987);
nand U1178 (N_1178,N_769,N_555);
or U1179 (N_1179,N_671,N_670);
or U1180 (N_1180,N_909,N_977);
or U1181 (N_1181,N_543,N_610);
and U1182 (N_1182,N_803,N_644);
nor U1183 (N_1183,N_993,N_650);
or U1184 (N_1184,N_992,N_721);
nand U1185 (N_1185,N_819,N_900);
nand U1186 (N_1186,N_702,N_746);
xor U1187 (N_1187,N_701,N_574);
nor U1188 (N_1188,N_810,N_604);
and U1189 (N_1189,N_962,N_600);
or U1190 (N_1190,N_967,N_636);
xor U1191 (N_1191,N_926,N_897);
xnor U1192 (N_1192,N_584,N_890);
xnor U1193 (N_1193,N_854,N_955);
nor U1194 (N_1194,N_794,N_710);
nor U1195 (N_1195,N_602,N_588);
nand U1196 (N_1196,N_718,N_598);
or U1197 (N_1197,N_533,N_622);
or U1198 (N_1198,N_896,N_770);
or U1199 (N_1199,N_512,N_911);
and U1200 (N_1200,N_572,N_587);
xor U1201 (N_1201,N_877,N_885);
xnor U1202 (N_1202,N_919,N_949);
and U1203 (N_1203,N_857,N_608);
or U1204 (N_1204,N_965,N_551);
xnor U1205 (N_1205,N_653,N_974);
nor U1206 (N_1206,N_733,N_723);
or U1207 (N_1207,N_874,N_867);
or U1208 (N_1208,N_996,N_743);
or U1209 (N_1209,N_731,N_814);
or U1210 (N_1210,N_853,N_639);
xor U1211 (N_1211,N_558,N_672);
nor U1212 (N_1212,N_788,N_850);
xor U1213 (N_1213,N_652,N_936);
and U1214 (N_1214,N_925,N_870);
nand U1215 (N_1215,N_941,N_694);
nor U1216 (N_1216,N_793,N_666);
nand U1217 (N_1217,N_530,N_779);
nor U1218 (N_1218,N_815,N_621);
and U1219 (N_1219,N_703,N_802);
and U1220 (N_1220,N_868,N_763);
and U1221 (N_1221,N_990,N_553);
and U1222 (N_1222,N_646,N_663);
xor U1223 (N_1223,N_774,N_995);
and U1224 (N_1224,N_843,N_664);
nor U1225 (N_1225,N_841,N_840);
nand U1226 (N_1226,N_626,N_762);
or U1227 (N_1227,N_882,N_503);
or U1228 (N_1228,N_662,N_851);
nor U1229 (N_1229,N_856,N_812);
nor U1230 (N_1230,N_765,N_989);
and U1231 (N_1231,N_579,N_898);
nand U1232 (N_1232,N_554,N_546);
nand U1233 (N_1233,N_726,N_645);
and U1234 (N_1234,N_716,N_568);
nand U1235 (N_1235,N_728,N_504);
nand U1236 (N_1236,N_781,N_994);
or U1237 (N_1237,N_651,N_929);
xor U1238 (N_1238,N_796,N_607);
and U1239 (N_1239,N_800,N_727);
and U1240 (N_1240,N_871,N_522);
nand U1241 (N_1241,N_669,N_816);
or U1242 (N_1242,N_657,N_708);
nor U1243 (N_1243,N_966,N_677);
nand U1244 (N_1244,N_643,N_944);
nor U1245 (N_1245,N_719,N_539);
nor U1246 (N_1246,N_715,N_538);
xor U1247 (N_1247,N_550,N_808);
and U1248 (N_1248,N_629,N_500);
or U1249 (N_1249,N_519,N_903);
or U1250 (N_1250,N_791,N_933);
xor U1251 (N_1251,N_791,N_960);
and U1252 (N_1252,N_858,N_925);
or U1253 (N_1253,N_520,N_675);
xor U1254 (N_1254,N_528,N_753);
and U1255 (N_1255,N_718,N_757);
and U1256 (N_1256,N_804,N_532);
nand U1257 (N_1257,N_763,N_811);
nand U1258 (N_1258,N_931,N_753);
and U1259 (N_1259,N_873,N_862);
nand U1260 (N_1260,N_831,N_976);
xor U1261 (N_1261,N_547,N_575);
xnor U1262 (N_1262,N_864,N_872);
and U1263 (N_1263,N_674,N_630);
nor U1264 (N_1264,N_858,N_891);
nor U1265 (N_1265,N_705,N_928);
and U1266 (N_1266,N_932,N_713);
nor U1267 (N_1267,N_879,N_581);
nor U1268 (N_1268,N_918,N_910);
or U1269 (N_1269,N_854,N_623);
nor U1270 (N_1270,N_836,N_598);
or U1271 (N_1271,N_837,N_733);
nand U1272 (N_1272,N_722,N_697);
or U1273 (N_1273,N_931,N_988);
nand U1274 (N_1274,N_949,N_540);
nand U1275 (N_1275,N_970,N_919);
xor U1276 (N_1276,N_609,N_616);
nand U1277 (N_1277,N_969,N_725);
nor U1278 (N_1278,N_628,N_876);
nand U1279 (N_1279,N_935,N_669);
and U1280 (N_1280,N_705,N_628);
or U1281 (N_1281,N_887,N_940);
nand U1282 (N_1282,N_964,N_926);
or U1283 (N_1283,N_785,N_538);
and U1284 (N_1284,N_526,N_642);
nand U1285 (N_1285,N_569,N_910);
or U1286 (N_1286,N_740,N_612);
and U1287 (N_1287,N_759,N_940);
and U1288 (N_1288,N_791,N_765);
and U1289 (N_1289,N_848,N_994);
xor U1290 (N_1290,N_618,N_716);
xor U1291 (N_1291,N_943,N_937);
and U1292 (N_1292,N_924,N_876);
nor U1293 (N_1293,N_898,N_725);
nor U1294 (N_1294,N_520,N_858);
or U1295 (N_1295,N_562,N_526);
nand U1296 (N_1296,N_874,N_737);
nor U1297 (N_1297,N_913,N_827);
xnor U1298 (N_1298,N_606,N_893);
nand U1299 (N_1299,N_585,N_814);
nand U1300 (N_1300,N_866,N_624);
or U1301 (N_1301,N_804,N_669);
xnor U1302 (N_1302,N_636,N_618);
and U1303 (N_1303,N_896,N_521);
xnor U1304 (N_1304,N_805,N_547);
or U1305 (N_1305,N_768,N_608);
nand U1306 (N_1306,N_643,N_684);
or U1307 (N_1307,N_542,N_691);
or U1308 (N_1308,N_732,N_568);
xor U1309 (N_1309,N_621,N_613);
or U1310 (N_1310,N_532,N_980);
or U1311 (N_1311,N_530,N_797);
nand U1312 (N_1312,N_785,N_557);
nand U1313 (N_1313,N_774,N_659);
xnor U1314 (N_1314,N_844,N_841);
nor U1315 (N_1315,N_683,N_764);
nand U1316 (N_1316,N_845,N_904);
nand U1317 (N_1317,N_686,N_843);
and U1318 (N_1318,N_774,N_618);
or U1319 (N_1319,N_874,N_632);
or U1320 (N_1320,N_569,N_613);
nor U1321 (N_1321,N_701,N_661);
or U1322 (N_1322,N_745,N_554);
nor U1323 (N_1323,N_889,N_785);
or U1324 (N_1324,N_640,N_594);
xnor U1325 (N_1325,N_821,N_503);
xor U1326 (N_1326,N_660,N_642);
xnor U1327 (N_1327,N_858,N_510);
nand U1328 (N_1328,N_826,N_753);
or U1329 (N_1329,N_913,N_944);
nor U1330 (N_1330,N_543,N_860);
nor U1331 (N_1331,N_983,N_523);
nand U1332 (N_1332,N_909,N_693);
nand U1333 (N_1333,N_953,N_744);
xor U1334 (N_1334,N_929,N_562);
xnor U1335 (N_1335,N_616,N_826);
xnor U1336 (N_1336,N_947,N_886);
nand U1337 (N_1337,N_768,N_985);
xnor U1338 (N_1338,N_831,N_630);
or U1339 (N_1339,N_652,N_682);
xor U1340 (N_1340,N_853,N_858);
and U1341 (N_1341,N_706,N_518);
and U1342 (N_1342,N_742,N_981);
nand U1343 (N_1343,N_883,N_650);
nor U1344 (N_1344,N_714,N_548);
nor U1345 (N_1345,N_823,N_587);
nor U1346 (N_1346,N_830,N_997);
xnor U1347 (N_1347,N_837,N_873);
nor U1348 (N_1348,N_823,N_907);
xnor U1349 (N_1349,N_676,N_822);
nand U1350 (N_1350,N_705,N_732);
xnor U1351 (N_1351,N_810,N_875);
nand U1352 (N_1352,N_890,N_751);
xnor U1353 (N_1353,N_547,N_589);
xor U1354 (N_1354,N_512,N_783);
nand U1355 (N_1355,N_827,N_557);
and U1356 (N_1356,N_810,N_727);
nand U1357 (N_1357,N_693,N_882);
and U1358 (N_1358,N_813,N_804);
nand U1359 (N_1359,N_917,N_712);
xnor U1360 (N_1360,N_591,N_602);
nor U1361 (N_1361,N_899,N_535);
and U1362 (N_1362,N_532,N_720);
nand U1363 (N_1363,N_889,N_762);
xor U1364 (N_1364,N_950,N_548);
nand U1365 (N_1365,N_921,N_869);
nor U1366 (N_1366,N_955,N_932);
nor U1367 (N_1367,N_882,N_802);
nand U1368 (N_1368,N_555,N_601);
nand U1369 (N_1369,N_566,N_910);
or U1370 (N_1370,N_606,N_649);
or U1371 (N_1371,N_571,N_756);
nor U1372 (N_1372,N_586,N_572);
nand U1373 (N_1373,N_856,N_666);
and U1374 (N_1374,N_953,N_831);
xor U1375 (N_1375,N_642,N_734);
xnor U1376 (N_1376,N_831,N_517);
xnor U1377 (N_1377,N_525,N_901);
nand U1378 (N_1378,N_708,N_739);
and U1379 (N_1379,N_972,N_843);
and U1380 (N_1380,N_996,N_862);
or U1381 (N_1381,N_607,N_542);
nand U1382 (N_1382,N_883,N_931);
nand U1383 (N_1383,N_518,N_912);
or U1384 (N_1384,N_995,N_689);
xor U1385 (N_1385,N_578,N_908);
nor U1386 (N_1386,N_951,N_841);
nor U1387 (N_1387,N_816,N_654);
nand U1388 (N_1388,N_931,N_843);
or U1389 (N_1389,N_795,N_617);
xor U1390 (N_1390,N_581,N_612);
or U1391 (N_1391,N_581,N_930);
or U1392 (N_1392,N_771,N_860);
nand U1393 (N_1393,N_646,N_630);
and U1394 (N_1394,N_906,N_962);
or U1395 (N_1395,N_697,N_886);
nor U1396 (N_1396,N_681,N_615);
or U1397 (N_1397,N_639,N_936);
and U1398 (N_1398,N_984,N_962);
nor U1399 (N_1399,N_745,N_988);
xnor U1400 (N_1400,N_796,N_941);
nand U1401 (N_1401,N_804,N_620);
nor U1402 (N_1402,N_564,N_500);
nor U1403 (N_1403,N_667,N_898);
and U1404 (N_1404,N_631,N_787);
nand U1405 (N_1405,N_848,N_802);
nor U1406 (N_1406,N_534,N_573);
and U1407 (N_1407,N_856,N_982);
or U1408 (N_1408,N_894,N_501);
xnor U1409 (N_1409,N_789,N_541);
nand U1410 (N_1410,N_977,N_792);
or U1411 (N_1411,N_936,N_649);
xnor U1412 (N_1412,N_600,N_550);
xor U1413 (N_1413,N_549,N_706);
nand U1414 (N_1414,N_687,N_811);
xnor U1415 (N_1415,N_699,N_823);
or U1416 (N_1416,N_524,N_922);
and U1417 (N_1417,N_573,N_588);
or U1418 (N_1418,N_725,N_674);
or U1419 (N_1419,N_585,N_731);
nor U1420 (N_1420,N_511,N_654);
nand U1421 (N_1421,N_563,N_875);
or U1422 (N_1422,N_529,N_833);
nor U1423 (N_1423,N_931,N_824);
and U1424 (N_1424,N_768,N_570);
and U1425 (N_1425,N_841,N_779);
nand U1426 (N_1426,N_535,N_560);
and U1427 (N_1427,N_797,N_608);
nor U1428 (N_1428,N_780,N_734);
or U1429 (N_1429,N_617,N_841);
or U1430 (N_1430,N_582,N_539);
or U1431 (N_1431,N_945,N_684);
xor U1432 (N_1432,N_813,N_807);
and U1433 (N_1433,N_865,N_631);
or U1434 (N_1434,N_846,N_991);
and U1435 (N_1435,N_693,N_850);
nor U1436 (N_1436,N_909,N_808);
nor U1437 (N_1437,N_704,N_651);
or U1438 (N_1438,N_610,N_655);
nand U1439 (N_1439,N_953,N_595);
or U1440 (N_1440,N_999,N_552);
or U1441 (N_1441,N_782,N_661);
and U1442 (N_1442,N_557,N_696);
and U1443 (N_1443,N_828,N_982);
or U1444 (N_1444,N_534,N_943);
and U1445 (N_1445,N_805,N_618);
or U1446 (N_1446,N_791,N_922);
nand U1447 (N_1447,N_640,N_692);
nor U1448 (N_1448,N_770,N_510);
nand U1449 (N_1449,N_647,N_939);
nor U1450 (N_1450,N_506,N_754);
nand U1451 (N_1451,N_627,N_646);
or U1452 (N_1452,N_926,N_857);
or U1453 (N_1453,N_690,N_978);
nand U1454 (N_1454,N_868,N_563);
xnor U1455 (N_1455,N_605,N_673);
and U1456 (N_1456,N_611,N_672);
or U1457 (N_1457,N_974,N_937);
xor U1458 (N_1458,N_866,N_776);
nor U1459 (N_1459,N_693,N_607);
nand U1460 (N_1460,N_904,N_720);
or U1461 (N_1461,N_945,N_667);
nand U1462 (N_1462,N_940,N_637);
nand U1463 (N_1463,N_981,N_992);
xnor U1464 (N_1464,N_546,N_988);
and U1465 (N_1465,N_617,N_973);
and U1466 (N_1466,N_697,N_729);
xor U1467 (N_1467,N_866,N_669);
xnor U1468 (N_1468,N_724,N_765);
or U1469 (N_1469,N_797,N_516);
xnor U1470 (N_1470,N_519,N_565);
xnor U1471 (N_1471,N_559,N_936);
nor U1472 (N_1472,N_522,N_786);
and U1473 (N_1473,N_644,N_816);
nor U1474 (N_1474,N_616,N_656);
nor U1475 (N_1475,N_946,N_958);
and U1476 (N_1476,N_540,N_820);
or U1477 (N_1477,N_744,N_872);
nand U1478 (N_1478,N_912,N_631);
nand U1479 (N_1479,N_523,N_889);
or U1480 (N_1480,N_556,N_654);
or U1481 (N_1481,N_791,N_700);
and U1482 (N_1482,N_825,N_815);
xor U1483 (N_1483,N_757,N_540);
and U1484 (N_1484,N_623,N_837);
nand U1485 (N_1485,N_581,N_706);
xor U1486 (N_1486,N_543,N_838);
nor U1487 (N_1487,N_895,N_703);
nand U1488 (N_1488,N_508,N_593);
and U1489 (N_1489,N_745,N_532);
or U1490 (N_1490,N_772,N_676);
nand U1491 (N_1491,N_521,N_734);
and U1492 (N_1492,N_901,N_812);
and U1493 (N_1493,N_774,N_519);
xnor U1494 (N_1494,N_746,N_926);
xnor U1495 (N_1495,N_888,N_816);
nand U1496 (N_1496,N_957,N_803);
nor U1497 (N_1497,N_975,N_547);
xnor U1498 (N_1498,N_803,N_535);
nor U1499 (N_1499,N_597,N_719);
xor U1500 (N_1500,N_1277,N_1464);
xor U1501 (N_1501,N_1062,N_1362);
and U1502 (N_1502,N_1018,N_1027);
nor U1503 (N_1503,N_1003,N_1143);
xnor U1504 (N_1504,N_1070,N_1310);
or U1505 (N_1505,N_1250,N_1407);
xnor U1506 (N_1506,N_1151,N_1110);
xor U1507 (N_1507,N_1431,N_1067);
xnor U1508 (N_1508,N_1488,N_1425);
nor U1509 (N_1509,N_1296,N_1429);
nor U1510 (N_1510,N_1242,N_1440);
xnor U1511 (N_1511,N_1372,N_1186);
nor U1512 (N_1512,N_1273,N_1320);
nand U1513 (N_1513,N_1017,N_1040);
or U1514 (N_1514,N_1265,N_1384);
and U1515 (N_1515,N_1031,N_1115);
nand U1516 (N_1516,N_1157,N_1267);
or U1517 (N_1517,N_1393,N_1126);
nand U1518 (N_1518,N_1466,N_1252);
nor U1519 (N_1519,N_1283,N_1288);
nand U1520 (N_1520,N_1079,N_1301);
xnor U1521 (N_1521,N_1063,N_1140);
nand U1522 (N_1522,N_1076,N_1181);
xor U1523 (N_1523,N_1292,N_1453);
nand U1524 (N_1524,N_1212,N_1246);
and U1525 (N_1525,N_1467,N_1385);
or U1526 (N_1526,N_1161,N_1328);
or U1527 (N_1527,N_1218,N_1111);
or U1528 (N_1528,N_1166,N_1034);
nand U1529 (N_1529,N_1257,N_1086);
xnor U1530 (N_1530,N_1089,N_1160);
nand U1531 (N_1531,N_1112,N_1432);
and U1532 (N_1532,N_1411,N_1336);
xnor U1533 (N_1533,N_1182,N_1338);
nand U1534 (N_1534,N_1285,N_1239);
xor U1535 (N_1535,N_1479,N_1287);
nor U1536 (N_1536,N_1356,N_1061);
xor U1537 (N_1537,N_1321,N_1081);
and U1538 (N_1538,N_1282,N_1192);
or U1539 (N_1539,N_1006,N_1108);
or U1540 (N_1540,N_1322,N_1378);
or U1541 (N_1541,N_1225,N_1430);
nor U1542 (N_1542,N_1189,N_1305);
nand U1543 (N_1543,N_1323,N_1256);
nand U1544 (N_1544,N_1368,N_1307);
nand U1545 (N_1545,N_1461,N_1355);
or U1546 (N_1546,N_1105,N_1138);
xnor U1547 (N_1547,N_1381,N_1291);
and U1548 (N_1548,N_1096,N_1264);
nand U1549 (N_1549,N_1318,N_1304);
xor U1550 (N_1550,N_1153,N_1162);
and U1551 (N_1551,N_1276,N_1102);
nor U1552 (N_1552,N_1200,N_1369);
nor U1553 (N_1553,N_1156,N_1021);
or U1554 (N_1554,N_1493,N_1434);
and U1555 (N_1555,N_1492,N_1275);
nor U1556 (N_1556,N_1311,N_1042);
nor U1557 (N_1557,N_1465,N_1316);
nor U1558 (N_1558,N_1187,N_1147);
nand U1559 (N_1559,N_1423,N_1215);
xnor U1560 (N_1560,N_1382,N_1405);
nand U1561 (N_1561,N_1216,N_1077);
or U1562 (N_1562,N_1404,N_1289);
and U1563 (N_1563,N_1145,N_1367);
xor U1564 (N_1564,N_1064,N_1202);
or U1565 (N_1565,N_1116,N_1066);
nor U1566 (N_1566,N_1420,N_1243);
and U1567 (N_1567,N_1317,N_1154);
or U1568 (N_1568,N_1005,N_1445);
nor U1569 (N_1569,N_1001,N_1053);
nor U1570 (N_1570,N_1210,N_1137);
or U1571 (N_1571,N_1051,N_1418);
or U1572 (N_1572,N_1417,N_1071);
nand U1573 (N_1573,N_1459,N_1130);
or U1574 (N_1574,N_1201,N_1188);
or U1575 (N_1575,N_1233,N_1036);
or U1576 (N_1576,N_1203,N_1221);
xnor U1577 (N_1577,N_1446,N_1023);
nor U1578 (N_1578,N_1073,N_1358);
xnor U1579 (N_1579,N_1414,N_1455);
nand U1580 (N_1580,N_1360,N_1072);
nand U1581 (N_1581,N_1350,N_1007);
and U1582 (N_1582,N_1090,N_1469);
nor U1583 (N_1583,N_1314,N_1004);
nor U1584 (N_1584,N_1100,N_1397);
and U1585 (N_1585,N_1364,N_1206);
or U1586 (N_1586,N_1424,N_1261);
and U1587 (N_1587,N_1389,N_1359);
and U1588 (N_1588,N_1391,N_1045);
and U1589 (N_1589,N_1290,N_1148);
xor U1590 (N_1590,N_1088,N_1176);
and U1591 (N_1591,N_1470,N_1142);
or U1592 (N_1592,N_1232,N_1178);
nand U1593 (N_1593,N_1085,N_1433);
and U1594 (N_1594,N_1244,N_1306);
nor U1595 (N_1595,N_1268,N_1131);
nor U1596 (N_1596,N_1030,N_1222);
nor U1597 (N_1597,N_1032,N_1150);
and U1598 (N_1598,N_1238,N_1341);
nand U1599 (N_1599,N_1240,N_1348);
and U1600 (N_1600,N_1164,N_1410);
xor U1601 (N_1601,N_1269,N_1334);
xnor U1602 (N_1602,N_1106,N_1319);
and U1603 (N_1603,N_1297,N_1002);
nor U1604 (N_1604,N_1228,N_1388);
xor U1605 (N_1605,N_1448,N_1068);
and U1606 (N_1606,N_1235,N_1226);
or U1607 (N_1607,N_1037,N_1443);
or U1608 (N_1608,N_1295,N_1398);
nand U1609 (N_1609,N_1191,N_1428);
xor U1610 (N_1610,N_1449,N_1353);
xnor U1611 (N_1611,N_1375,N_1029);
nor U1612 (N_1612,N_1020,N_1444);
nand U1613 (N_1613,N_1139,N_1167);
nor U1614 (N_1614,N_1195,N_1000);
or U1615 (N_1615,N_1087,N_1286);
or U1616 (N_1616,N_1011,N_1041);
or U1617 (N_1617,N_1128,N_1422);
xor U1618 (N_1618,N_1097,N_1019);
nand U1619 (N_1619,N_1025,N_1190);
nor U1620 (N_1620,N_1333,N_1121);
nand U1621 (N_1621,N_1141,N_1183);
and U1622 (N_1622,N_1075,N_1409);
and U1623 (N_1623,N_1386,N_1284);
or U1624 (N_1624,N_1241,N_1223);
nor U1625 (N_1625,N_1207,N_1024);
nand U1626 (N_1626,N_1117,N_1456);
nand U1627 (N_1627,N_1331,N_1408);
or U1628 (N_1628,N_1308,N_1315);
nand U1629 (N_1629,N_1054,N_1229);
and U1630 (N_1630,N_1083,N_1069);
xnor U1631 (N_1631,N_1109,N_1294);
and U1632 (N_1632,N_1494,N_1281);
and U1633 (N_1633,N_1196,N_1047);
or U1634 (N_1634,N_1374,N_1342);
and U1635 (N_1635,N_1033,N_1026);
and U1636 (N_1636,N_1132,N_1199);
or U1637 (N_1637,N_1171,N_1124);
and U1638 (N_1638,N_1149,N_1234);
nand U1639 (N_1639,N_1413,N_1330);
xor U1640 (N_1640,N_1078,N_1458);
nor U1641 (N_1641,N_1114,N_1415);
nand U1642 (N_1642,N_1123,N_1379);
or U1643 (N_1643,N_1231,N_1399);
xor U1644 (N_1644,N_1266,N_1390);
and U1645 (N_1645,N_1122,N_1103);
nand U1646 (N_1646,N_1274,N_1476);
nor U1647 (N_1647,N_1058,N_1474);
nor U1648 (N_1648,N_1173,N_1401);
nand U1649 (N_1649,N_1133,N_1043);
nor U1650 (N_1650,N_1230,N_1349);
and U1651 (N_1651,N_1208,N_1329);
and U1652 (N_1652,N_1074,N_1158);
and U1653 (N_1653,N_1416,N_1412);
nor U1654 (N_1654,N_1254,N_1022);
nand U1655 (N_1655,N_1155,N_1302);
and U1656 (N_1656,N_1351,N_1473);
nor U1657 (N_1657,N_1457,N_1056);
or U1658 (N_1658,N_1480,N_1094);
nor U1659 (N_1659,N_1028,N_1263);
nor U1660 (N_1660,N_1344,N_1193);
and U1661 (N_1661,N_1332,N_1435);
nand U1662 (N_1662,N_1272,N_1335);
nor U1663 (N_1663,N_1395,N_1146);
and U1664 (N_1664,N_1217,N_1471);
nand U1665 (N_1665,N_1454,N_1259);
xor U1666 (N_1666,N_1481,N_1120);
xor U1667 (N_1667,N_1213,N_1484);
xor U1668 (N_1668,N_1441,N_1144);
and U1669 (N_1669,N_1490,N_1383);
or U1670 (N_1670,N_1371,N_1487);
nor U1671 (N_1671,N_1013,N_1377);
xnor U1672 (N_1672,N_1361,N_1278);
xor U1673 (N_1673,N_1326,N_1271);
and U1674 (N_1674,N_1038,N_1236);
nor U1675 (N_1675,N_1249,N_1224);
xnor U1676 (N_1676,N_1172,N_1245);
nand U1677 (N_1677,N_1468,N_1169);
and U1678 (N_1678,N_1387,N_1175);
nand U1679 (N_1679,N_1402,N_1299);
and U1680 (N_1680,N_1174,N_1127);
nor U1681 (N_1681,N_1039,N_1357);
nand U1682 (N_1682,N_1309,N_1486);
or U1683 (N_1683,N_1303,N_1060);
nand U1684 (N_1684,N_1477,N_1209);
and U1685 (N_1685,N_1101,N_1119);
xor U1686 (N_1686,N_1248,N_1496);
nor U1687 (N_1687,N_1392,N_1099);
and U1688 (N_1688,N_1159,N_1373);
nand U1689 (N_1689,N_1170,N_1394);
nand U1690 (N_1690,N_1179,N_1452);
and U1691 (N_1691,N_1253,N_1055);
nand U1692 (N_1692,N_1442,N_1214);
and U1693 (N_1693,N_1312,N_1168);
xnor U1694 (N_1694,N_1472,N_1046);
or U1695 (N_1695,N_1135,N_1107);
nand U1696 (N_1696,N_1498,N_1439);
or U1697 (N_1697,N_1325,N_1211);
xnor U1698 (N_1698,N_1491,N_1050);
or U1699 (N_1699,N_1363,N_1009);
or U1700 (N_1700,N_1340,N_1347);
nand U1701 (N_1701,N_1258,N_1300);
xor U1702 (N_1702,N_1419,N_1237);
xor U1703 (N_1703,N_1082,N_1365);
xnor U1704 (N_1704,N_1447,N_1396);
nor U1705 (N_1705,N_1016,N_1092);
nand U1706 (N_1706,N_1354,N_1197);
xnor U1707 (N_1707,N_1483,N_1205);
xor U1708 (N_1708,N_1093,N_1380);
xor U1709 (N_1709,N_1184,N_1489);
or U1710 (N_1710,N_1052,N_1339);
and U1711 (N_1711,N_1298,N_1293);
and U1712 (N_1712,N_1014,N_1015);
nor U1713 (N_1713,N_1482,N_1426);
nor U1714 (N_1714,N_1185,N_1163);
nand U1715 (N_1715,N_1366,N_1012);
or U1716 (N_1716,N_1352,N_1194);
xnor U1717 (N_1717,N_1048,N_1497);
nor U1718 (N_1718,N_1118,N_1437);
xnor U1719 (N_1719,N_1057,N_1421);
or U1720 (N_1720,N_1251,N_1113);
xnor U1721 (N_1721,N_1403,N_1136);
nand U1722 (N_1722,N_1080,N_1499);
and U1723 (N_1723,N_1125,N_1345);
nand U1724 (N_1724,N_1427,N_1152);
xor U1725 (N_1725,N_1084,N_1436);
or U1726 (N_1726,N_1337,N_1262);
xnor U1727 (N_1727,N_1279,N_1327);
nand U1728 (N_1728,N_1462,N_1280);
and U1729 (N_1729,N_1495,N_1400);
nor U1730 (N_1730,N_1451,N_1460);
or U1731 (N_1731,N_1247,N_1227);
nor U1732 (N_1732,N_1091,N_1478);
or U1733 (N_1733,N_1165,N_1270);
or U1734 (N_1734,N_1219,N_1065);
nor U1735 (N_1735,N_1049,N_1044);
or U1736 (N_1736,N_1346,N_1485);
nor U1737 (N_1737,N_1475,N_1059);
xor U1738 (N_1738,N_1260,N_1343);
and U1739 (N_1739,N_1129,N_1095);
xnor U1740 (N_1740,N_1134,N_1010);
nor U1741 (N_1741,N_1104,N_1180);
nand U1742 (N_1742,N_1204,N_1324);
xor U1743 (N_1743,N_1376,N_1406);
nand U1744 (N_1744,N_1198,N_1008);
nand U1745 (N_1745,N_1255,N_1438);
xnor U1746 (N_1746,N_1463,N_1220);
nand U1747 (N_1747,N_1450,N_1313);
and U1748 (N_1748,N_1177,N_1370);
or U1749 (N_1749,N_1098,N_1035);
nor U1750 (N_1750,N_1324,N_1121);
nor U1751 (N_1751,N_1336,N_1222);
and U1752 (N_1752,N_1362,N_1181);
xor U1753 (N_1753,N_1429,N_1242);
nand U1754 (N_1754,N_1469,N_1101);
and U1755 (N_1755,N_1074,N_1391);
nand U1756 (N_1756,N_1325,N_1064);
nand U1757 (N_1757,N_1420,N_1328);
nand U1758 (N_1758,N_1193,N_1327);
and U1759 (N_1759,N_1061,N_1339);
xor U1760 (N_1760,N_1048,N_1181);
xnor U1761 (N_1761,N_1249,N_1170);
and U1762 (N_1762,N_1136,N_1438);
nand U1763 (N_1763,N_1245,N_1461);
nand U1764 (N_1764,N_1259,N_1152);
xnor U1765 (N_1765,N_1121,N_1453);
nand U1766 (N_1766,N_1437,N_1482);
nand U1767 (N_1767,N_1143,N_1451);
or U1768 (N_1768,N_1409,N_1303);
or U1769 (N_1769,N_1388,N_1007);
nor U1770 (N_1770,N_1141,N_1146);
or U1771 (N_1771,N_1015,N_1372);
xor U1772 (N_1772,N_1062,N_1363);
nand U1773 (N_1773,N_1347,N_1189);
nand U1774 (N_1774,N_1177,N_1487);
nor U1775 (N_1775,N_1184,N_1209);
xor U1776 (N_1776,N_1032,N_1197);
or U1777 (N_1777,N_1304,N_1238);
or U1778 (N_1778,N_1266,N_1115);
nor U1779 (N_1779,N_1167,N_1208);
nor U1780 (N_1780,N_1441,N_1246);
and U1781 (N_1781,N_1368,N_1084);
and U1782 (N_1782,N_1179,N_1462);
or U1783 (N_1783,N_1144,N_1387);
or U1784 (N_1784,N_1336,N_1042);
nor U1785 (N_1785,N_1202,N_1177);
xnor U1786 (N_1786,N_1297,N_1384);
and U1787 (N_1787,N_1459,N_1478);
nand U1788 (N_1788,N_1262,N_1324);
xor U1789 (N_1789,N_1142,N_1219);
nor U1790 (N_1790,N_1070,N_1449);
xor U1791 (N_1791,N_1426,N_1195);
nor U1792 (N_1792,N_1165,N_1356);
nor U1793 (N_1793,N_1310,N_1231);
xnor U1794 (N_1794,N_1371,N_1460);
nand U1795 (N_1795,N_1114,N_1175);
nor U1796 (N_1796,N_1226,N_1085);
and U1797 (N_1797,N_1063,N_1468);
and U1798 (N_1798,N_1466,N_1206);
or U1799 (N_1799,N_1104,N_1394);
xnor U1800 (N_1800,N_1009,N_1372);
or U1801 (N_1801,N_1215,N_1004);
nor U1802 (N_1802,N_1034,N_1457);
nor U1803 (N_1803,N_1437,N_1196);
or U1804 (N_1804,N_1096,N_1417);
xnor U1805 (N_1805,N_1407,N_1495);
nor U1806 (N_1806,N_1045,N_1281);
xnor U1807 (N_1807,N_1031,N_1060);
or U1808 (N_1808,N_1142,N_1459);
nor U1809 (N_1809,N_1054,N_1495);
and U1810 (N_1810,N_1313,N_1081);
or U1811 (N_1811,N_1449,N_1294);
xnor U1812 (N_1812,N_1071,N_1014);
xor U1813 (N_1813,N_1233,N_1140);
nand U1814 (N_1814,N_1155,N_1484);
xor U1815 (N_1815,N_1033,N_1084);
xor U1816 (N_1816,N_1009,N_1331);
nand U1817 (N_1817,N_1363,N_1454);
nand U1818 (N_1818,N_1190,N_1330);
nand U1819 (N_1819,N_1317,N_1435);
and U1820 (N_1820,N_1143,N_1080);
nand U1821 (N_1821,N_1243,N_1466);
nand U1822 (N_1822,N_1135,N_1196);
nor U1823 (N_1823,N_1473,N_1340);
xor U1824 (N_1824,N_1024,N_1052);
nor U1825 (N_1825,N_1290,N_1208);
nand U1826 (N_1826,N_1099,N_1066);
or U1827 (N_1827,N_1047,N_1358);
nor U1828 (N_1828,N_1099,N_1032);
and U1829 (N_1829,N_1092,N_1169);
or U1830 (N_1830,N_1467,N_1430);
nand U1831 (N_1831,N_1491,N_1361);
and U1832 (N_1832,N_1043,N_1165);
xnor U1833 (N_1833,N_1145,N_1496);
nor U1834 (N_1834,N_1023,N_1077);
nand U1835 (N_1835,N_1448,N_1026);
and U1836 (N_1836,N_1454,N_1312);
or U1837 (N_1837,N_1260,N_1415);
and U1838 (N_1838,N_1346,N_1407);
xor U1839 (N_1839,N_1022,N_1027);
and U1840 (N_1840,N_1343,N_1419);
nand U1841 (N_1841,N_1022,N_1196);
nor U1842 (N_1842,N_1441,N_1182);
nand U1843 (N_1843,N_1167,N_1196);
and U1844 (N_1844,N_1252,N_1357);
and U1845 (N_1845,N_1178,N_1153);
nand U1846 (N_1846,N_1208,N_1097);
nand U1847 (N_1847,N_1079,N_1227);
and U1848 (N_1848,N_1490,N_1373);
nand U1849 (N_1849,N_1486,N_1189);
nor U1850 (N_1850,N_1272,N_1394);
nor U1851 (N_1851,N_1093,N_1112);
nor U1852 (N_1852,N_1392,N_1150);
or U1853 (N_1853,N_1346,N_1273);
nor U1854 (N_1854,N_1226,N_1275);
and U1855 (N_1855,N_1039,N_1199);
and U1856 (N_1856,N_1003,N_1245);
and U1857 (N_1857,N_1402,N_1138);
nand U1858 (N_1858,N_1225,N_1008);
or U1859 (N_1859,N_1113,N_1436);
xnor U1860 (N_1860,N_1100,N_1385);
and U1861 (N_1861,N_1174,N_1258);
and U1862 (N_1862,N_1216,N_1199);
xor U1863 (N_1863,N_1154,N_1186);
or U1864 (N_1864,N_1230,N_1238);
nor U1865 (N_1865,N_1422,N_1147);
nand U1866 (N_1866,N_1300,N_1482);
nor U1867 (N_1867,N_1012,N_1104);
xnor U1868 (N_1868,N_1100,N_1414);
and U1869 (N_1869,N_1274,N_1287);
xor U1870 (N_1870,N_1336,N_1001);
and U1871 (N_1871,N_1384,N_1068);
nor U1872 (N_1872,N_1065,N_1416);
xor U1873 (N_1873,N_1497,N_1411);
nand U1874 (N_1874,N_1412,N_1417);
and U1875 (N_1875,N_1319,N_1167);
nor U1876 (N_1876,N_1251,N_1104);
or U1877 (N_1877,N_1084,N_1024);
xor U1878 (N_1878,N_1366,N_1356);
or U1879 (N_1879,N_1027,N_1158);
nor U1880 (N_1880,N_1104,N_1492);
or U1881 (N_1881,N_1493,N_1115);
and U1882 (N_1882,N_1176,N_1321);
xnor U1883 (N_1883,N_1396,N_1091);
xor U1884 (N_1884,N_1069,N_1255);
xnor U1885 (N_1885,N_1407,N_1107);
and U1886 (N_1886,N_1125,N_1301);
nand U1887 (N_1887,N_1471,N_1177);
nor U1888 (N_1888,N_1474,N_1138);
or U1889 (N_1889,N_1314,N_1137);
nor U1890 (N_1890,N_1126,N_1213);
or U1891 (N_1891,N_1458,N_1312);
nor U1892 (N_1892,N_1207,N_1450);
nor U1893 (N_1893,N_1125,N_1269);
or U1894 (N_1894,N_1039,N_1027);
or U1895 (N_1895,N_1378,N_1279);
nor U1896 (N_1896,N_1132,N_1151);
nor U1897 (N_1897,N_1418,N_1096);
and U1898 (N_1898,N_1189,N_1391);
or U1899 (N_1899,N_1346,N_1434);
xnor U1900 (N_1900,N_1392,N_1024);
xnor U1901 (N_1901,N_1458,N_1347);
nand U1902 (N_1902,N_1022,N_1217);
or U1903 (N_1903,N_1443,N_1263);
nor U1904 (N_1904,N_1356,N_1100);
nand U1905 (N_1905,N_1080,N_1396);
or U1906 (N_1906,N_1390,N_1290);
and U1907 (N_1907,N_1377,N_1473);
or U1908 (N_1908,N_1439,N_1447);
nor U1909 (N_1909,N_1125,N_1425);
xor U1910 (N_1910,N_1435,N_1446);
or U1911 (N_1911,N_1002,N_1050);
xor U1912 (N_1912,N_1028,N_1200);
xnor U1913 (N_1913,N_1059,N_1378);
xor U1914 (N_1914,N_1357,N_1316);
or U1915 (N_1915,N_1344,N_1028);
nand U1916 (N_1916,N_1300,N_1344);
or U1917 (N_1917,N_1465,N_1139);
nand U1918 (N_1918,N_1018,N_1396);
nor U1919 (N_1919,N_1390,N_1301);
xor U1920 (N_1920,N_1258,N_1371);
nand U1921 (N_1921,N_1438,N_1230);
nand U1922 (N_1922,N_1100,N_1417);
nand U1923 (N_1923,N_1319,N_1345);
and U1924 (N_1924,N_1039,N_1362);
nand U1925 (N_1925,N_1445,N_1052);
and U1926 (N_1926,N_1074,N_1472);
xnor U1927 (N_1927,N_1253,N_1453);
nand U1928 (N_1928,N_1299,N_1427);
nor U1929 (N_1929,N_1215,N_1201);
nand U1930 (N_1930,N_1406,N_1227);
or U1931 (N_1931,N_1358,N_1417);
and U1932 (N_1932,N_1484,N_1367);
nand U1933 (N_1933,N_1283,N_1372);
or U1934 (N_1934,N_1363,N_1056);
or U1935 (N_1935,N_1073,N_1128);
and U1936 (N_1936,N_1059,N_1096);
nand U1937 (N_1937,N_1012,N_1146);
nand U1938 (N_1938,N_1145,N_1102);
xnor U1939 (N_1939,N_1016,N_1103);
nor U1940 (N_1940,N_1237,N_1154);
nor U1941 (N_1941,N_1174,N_1224);
or U1942 (N_1942,N_1010,N_1031);
or U1943 (N_1943,N_1469,N_1223);
nor U1944 (N_1944,N_1417,N_1360);
nand U1945 (N_1945,N_1395,N_1266);
or U1946 (N_1946,N_1151,N_1369);
xnor U1947 (N_1947,N_1048,N_1323);
nand U1948 (N_1948,N_1024,N_1290);
nand U1949 (N_1949,N_1371,N_1417);
nor U1950 (N_1950,N_1343,N_1108);
nor U1951 (N_1951,N_1477,N_1311);
nand U1952 (N_1952,N_1115,N_1481);
xnor U1953 (N_1953,N_1373,N_1163);
nand U1954 (N_1954,N_1344,N_1127);
xnor U1955 (N_1955,N_1317,N_1300);
and U1956 (N_1956,N_1257,N_1337);
xor U1957 (N_1957,N_1175,N_1290);
nor U1958 (N_1958,N_1114,N_1405);
and U1959 (N_1959,N_1340,N_1272);
or U1960 (N_1960,N_1405,N_1066);
and U1961 (N_1961,N_1085,N_1027);
or U1962 (N_1962,N_1218,N_1246);
or U1963 (N_1963,N_1116,N_1158);
nor U1964 (N_1964,N_1113,N_1450);
or U1965 (N_1965,N_1431,N_1179);
and U1966 (N_1966,N_1345,N_1257);
and U1967 (N_1967,N_1234,N_1335);
xnor U1968 (N_1968,N_1241,N_1378);
nand U1969 (N_1969,N_1192,N_1157);
and U1970 (N_1970,N_1413,N_1364);
xnor U1971 (N_1971,N_1393,N_1191);
xor U1972 (N_1972,N_1172,N_1300);
or U1973 (N_1973,N_1456,N_1419);
nand U1974 (N_1974,N_1203,N_1106);
xor U1975 (N_1975,N_1352,N_1482);
xnor U1976 (N_1976,N_1486,N_1094);
xor U1977 (N_1977,N_1477,N_1247);
and U1978 (N_1978,N_1069,N_1165);
or U1979 (N_1979,N_1042,N_1256);
nor U1980 (N_1980,N_1041,N_1117);
or U1981 (N_1981,N_1002,N_1340);
nand U1982 (N_1982,N_1021,N_1143);
nand U1983 (N_1983,N_1399,N_1308);
nand U1984 (N_1984,N_1354,N_1037);
nand U1985 (N_1985,N_1409,N_1129);
xor U1986 (N_1986,N_1168,N_1293);
xnor U1987 (N_1987,N_1041,N_1105);
xnor U1988 (N_1988,N_1155,N_1462);
nor U1989 (N_1989,N_1422,N_1086);
nand U1990 (N_1990,N_1379,N_1137);
nor U1991 (N_1991,N_1270,N_1111);
and U1992 (N_1992,N_1170,N_1183);
nand U1993 (N_1993,N_1117,N_1096);
or U1994 (N_1994,N_1490,N_1311);
xor U1995 (N_1995,N_1083,N_1420);
xnor U1996 (N_1996,N_1352,N_1432);
xor U1997 (N_1997,N_1120,N_1192);
xor U1998 (N_1998,N_1375,N_1282);
or U1999 (N_1999,N_1395,N_1260);
xnor U2000 (N_2000,N_1899,N_1877);
nor U2001 (N_2001,N_1663,N_1523);
nand U2002 (N_2002,N_1551,N_1774);
or U2003 (N_2003,N_1506,N_1697);
or U2004 (N_2004,N_1565,N_1511);
and U2005 (N_2005,N_1768,N_1696);
and U2006 (N_2006,N_1924,N_1786);
xnor U2007 (N_2007,N_1821,N_1519);
nor U2008 (N_2008,N_1871,N_1676);
and U2009 (N_2009,N_1829,N_1524);
nand U2010 (N_2010,N_1571,N_1955);
nand U2011 (N_2011,N_1935,N_1732);
nand U2012 (N_2012,N_1549,N_1628);
xor U2013 (N_2013,N_1531,N_1545);
and U2014 (N_2014,N_1611,N_1974);
nand U2015 (N_2015,N_1804,N_1714);
xnor U2016 (N_2016,N_1527,N_1603);
nor U2017 (N_2017,N_1558,N_1639);
nor U2018 (N_2018,N_1529,N_1843);
or U2019 (N_2019,N_1929,N_1751);
xnor U2020 (N_2020,N_1823,N_1706);
and U2021 (N_2021,N_1852,N_1967);
and U2022 (N_2022,N_1678,N_1770);
nor U2023 (N_2023,N_1728,N_1956);
and U2024 (N_2024,N_1841,N_1637);
nor U2025 (N_2025,N_1691,N_1937);
xor U2026 (N_2026,N_1972,N_1857);
and U2027 (N_2027,N_1689,N_1906);
nor U2028 (N_2028,N_1748,N_1606);
nor U2029 (N_2029,N_1550,N_1954);
nand U2030 (N_2030,N_1862,N_1579);
nand U2031 (N_2031,N_1573,N_1503);
nand U2032 (N_2032,N_1743,N_1810);
nor U2033 (N_2033,N_1828,N_1636);
and U2034 (N_2034,N_1787,N_1845);
xor U2035 (N_2035,N_1807,N_1630);
xnor U2036 (N_2036,N_1576,N_1615);
nand U2037 (N_2037,N_1819,N_1960);
xor U2038 (N_2038,N_1713,N_1502);
and U2039 (N_2039,N_1923,N_1522);
xor U2040 (N_2040,N_1901,N_1759);
and U2041 (N_2041,N_1656,N_1802);
and U2042 (N_2042,N_1648,N_1936);
nor U2043 (N_2043,N_1569,N_1831);
xnor U2044 (N_2044,N_1913,N_1780);
xor U2045 (N_2045,N_1538,N_1561);
nor U2046 (N_2046,N_1870,N_1632);
nor U2047 (N_2047,N_1698,N_1994);
or U2048 (N_2048,N_1948,N_1757);
and U2049 (N_2049,N_1659,N_1957);
or U2050 (N_2050,N_1812,N_1905);
or U2051 (N_2051,N_1629,N_1747);
or U2052 (N_2052,N_1730,N_1863);
nor U2053 (N_2053,N_1613,N_1975);
nand U2054 (N_2054,N_1799,N_1682);
nand U2055 (N_2055,N_1512,N_1825);
xnor U2056 (N_2056,N_1866,N_1992);
nor U2057 (N_2057,N_1540,N_1851);
or U2058 (N_2058,N_1530,N_1782);
nor U2059 (N_2059,N_1702,N_1800);
nor U2060 (N_2060,N_1820,N_1650);
or U2061 (N_2061,N_1541,N_1814);
and U2062 (N_2062,N_1575,N_1869);
xnor U2063 (N_2063,N_1720,N_1601);
nor U2064 (N_2064,N_1670,N_1796);
or U2065 (N_2065,N_1805,N_1900);
or U2066 (N_2066,N_1641,N_1791);
nor U2067 (N_2067,N_1908,N_1574);
nand U2068 (N_2068,N_1947,N_1764);
xnor U2069 (N_2069,N_1915,N_1944);
xor U2070 (N_2070,N_1710,N_1931);
nand U2071 (N_2071,N_1535,N_1942);
xnor U2072 (N_2072,N_1912,N_1625);
nand U2073 (N_2073,N_1976,N_1952);
nand U2074 (N_2074,N_1722,N_1649);
and U2075 (N_2075,N_1539,N_1508);
and U2076 (N_2076,N_1513,N_1958);
or U2077 (N_2077,N_1723,N_1874);
or U2078 (N_2078,N_1635,N_1612);
nor U2079 (N_2079,N_1907,N_1623);
nor U2080 (N_2080,N_1662,N_1679);
or U2081 (N_2081,N_1646,N_1701);
xnor U2082 (N_2082,N_1904,N_1660);
xor U2083 (N_2083,N_1963,N_1744);
nor U2084 (N_2084,N_1991,N_1693);
and U2085 (N_2085,N_1520,N_1617);
nand U2086 (N_2086,N_1951,N_1703);
nand U2087 (N_2087,N_1563,N_1627);
nand U2088 (N_2088,N_1634,N_1669);
nor U2089 (N_2089,N_1980,N_1715);
and U2090 (N_2090,N_1822,N_1528);
xnor U2091 (N_2091,N_1890,N_1811);
nand U2092 (N_2092,N_1547,N_1622);
xor U2093 (N_2093,N_1762,N_1880);
nand U2094 (N_2094,N_1784,N_1927);
and U2095 (N_2095,N_1969,N_1752);
xor U2096 (N_2096,N_1582,N_1883);
or U2097 (N_2097,N_1794,N_1911);
or U2098 (N_2098,N_1775,N_1917);
xnor U2099 (N_2099,N_1626,N_1729);
nor U2100 (N_2100,N_1847,N_1655);
nor U2101 (N_2101,N_1588,N_1769);
nor U2102 (N_2102,N_1586,N_1504);
and U2103 (N_2103,N_1643,N_1647);
nor U2104 (N_2104,N_1688,N_1946);
xor U2105 (N_2105,N_1716,N_1602);
or U2106 (N_2106,N_1749,N_1882);
xnor U2107 (N_2107,N_1705,N_1711);
nor U2108 (N_2108,N_1961,N_1846);
nor U2109 (N_2109,N_1718,N_1884);
or U2110 (N_2110,N_1939,N_1661);
nand U2111 (N_2111,N_1526,N_1704);
xnor U2112 (N_2112,N_1887,N_1808);
or U2113 (N_2113,N_1839,N_1872);
nand U2114 (N_2114,N_1668,N_1973);
nor U2115 (N_2115,N_1577,N_1681);
nor U2116 (N_2116,N_1949,N_1971);
nand U2117 (N_2117,N_1848,N_1785);
and U2118 (N_2118,N_1950,N_1754);
nor U2119 (N_2119,N_1885,N_1867);
xnor U2120 (N_2120,N_1733,N_1806);
xor U2121 (N_2121,N_1532,N_1817);
or U2122 (N_2122,N_1608,N_1621);
or U2123 (N_2123,N_1683,N_1832);
xnor U2124 (N_2124,N_1798,N_1809);
nor U2125 (N_2125,N_1797,N_1999);
nor U2126 (N_2126,N_1510,N_1584);
and U2127 (N_2127,N_1836,N_1654);
xnor U2128 (N_2128,N_1858,N_1793);
and U2129 (N_2129,N_1690,N_1583);
nand U2130 (N_2130,N_1645,N_1995);
nand U2131 (N_2131,N_1566,N_1940);
xnor U2132 (N_2132,N_1578,N_1624);
and U2133 (N_2133,N_1966,N_1544);
nand U2134 (N_2134,N_1835,N_1983);
nand U2135 (N_2135,N_1868,N_1607);
xor U2136 (N_2136,N_1855,N_1505);
nor U2137 (N_2137,N_1988,N_1902);
xnor U2138 (N_2138,N_1555,N_1777);
and U2139 (N_2139,N_1968,N_1631);
and U2140 (N_2140,N_1542,N_1554);
and U2141 (N_2141,N_1614,N_1761);
nor U2142 (N_2142,N_1861,N_1543);
or U2143 (N_2143,N_1776,N_1596);
xor U2144 (N_2144,N_1687,N_1840);
and U2145 (N_2145,N_1739,N_1604);
xnor U2146 (N_2146,N_1965,N_1515);
or U2147 (N_2147,N_1772,N_1842);
nand U2148 (N_2148,N_1894,N_1984);
nor U2149 (N_2149,N_1849,N_1589);
or U2150 (N_2150,N_1640,N_1767);
and U2151 (N_2151,N_1572,N_1964);
or U2152 (N_2152,N_1897,N_1712);
xnor U2153 (N_2153,N_1516,N_1719);
or U2154 (N_2154,N_1620,N_1567);
and U2155 (N_2155,N_1844,N_1667);
or U2156 (N_2156,N_1920,N_1664);
or U2157 (N_2157,N_1593,N_1826);
or U2158 (N_2158,N_1982,N_1735);
and U2159 (N_2159,N_1738,N_1537);
or U2160 (N_2160,N_1933,N_1909);
xor U2161 (N_2161,N_1673,N_1953);
xor U2162 (N_2162,N_1765,N_1993);
or U2163 (N_2163,N_1590,N_1921);
or U2164 (N_2164,N_1987,N_1671);
or U2165 (N_2165,N_1830,N_1592);
nor U2166 (N_2166,N_1680,N_1824);
and U2167 (N_2167,N_1600,N_1658);
nor U2168 (N_2168,N_1896,N_1653);
and U2169 (N_2169,N_1779,N_1928);
or U2170 (N_2170,N_1657,N_1865);
nor U2171 (N_2171,N_1795,N_1644);
nor U2172 (N_2172,N_1708,N_1979);
nand U2173 (N_2173,N_1756,N_1591);
xor U2174 (N_2174,N_1943,N_1781);
and U2175 (N_2175,N_1707,N_1803);
xor U2176 (N_2176,N_1815,N_1986);
xor U2177 (N_2177,N_1652,N_1609);
nand U2178 (N_2178,N_1737,N_1699);
and U2179 (N_2179,N_1580,N_1721);
nor U2180 (N_2180,N_1709,N_1546);
nor U2181 (N_2181,N_1587,N_1694);
xnor U2182 (N_2182,N_1916,N_1695);
nor U2183 (N_2183,N_1557,N_1918);
or U2184 (N_2184,N_1568,N_1534);
nand U2185 (N_2185,N_1581,N_1521);
and U2186 (N_2186,N_1789,N_1878);
and U2187 (N_2187,N_1881,N_1903);
or U2188 (N_2188,N_1941,N_1560);
xnor U2189 (N_2189,N_1758,N_1585);
xnor U2190 (N_2190,N_1919,N_1666);
xnor U2191 (N_2191,N_1850,N_1597);
or U2192 (N_2192,N_1753,N_1598);
and U2193 (N_2193,N_1684,N_1638);
or U2194 (N_2194,N_1605,N_1856);
xor U2195 (N_2195,N_1700,N_1938);
and U2196 (N_2196,N_1834,N_1788);
xnor U2197 (N_2197,N_1562,N_1692);
and U2198 (N_2198,N_1559,N_1792);
xnor U2199 (N_2199,N_1893,N_1518);
or U2200 (N_2200,N_1734,N_1517);
nor U2201 (N_2201,N_1766,N_1548);
and U2202 (N_2202,N_1594,N_1536);
nor U2203 (N_2203,N_1818,N_1886);
nor U2204 (N_2204,N_1990,N_1790);
nand U2205 (N_2205,N_1783,N_1760);
or U2206 (N_2206,N_1686,N_1501);
nand U2207 (N_2207,N_1827,N_1771);
or U2208 (N_2208,N_1962,N_1926);
or U2209 (N_2209,N_1595,N_1533);
xnor U2210 (N_2210,N_1552,N_1860);
nor U2211 (N_2211,N_1778,N_1674);
nor U2212 (N_2212,N_1616,N_1977);
and U2213 (N_2213,N_1833,N_1736);
nand U2214 (N_2214,N_1997,N_1816);
nor U2215 (N_2215,N_1932,N_1981);
nand U2216 (N_2216,N_1672,N_1888);
nor U2217 (N_2217,N_1556,N_1685);
or U2218 (N_2218,N_1970,N_1898);
or U2219 (N_2219,N_1876,N_1773);
and U2220 (N_2220,N_1910,N_1813);
and U2221 (N_2221,N_1922,N_1746);
nand U2222 (N_2222,N_1665,N_1989);
nor U2223 (N_2223,N_1564,N_1740);
or U2224 (N_2224,N_1837,N_1642);
nor U2225 (N_2225,N_1978,N_1500);
nor U2226 (N_2226,N_1755,N_1717);
nand U2227 (N_2227,N_1725,N_1879);
and U2228 (N_2228,N_1891,N_1873);
nor U2229 (N_2229,N_1763,N_1934);
nor U2230 (N_2230,N_1619,N_1914);
or U2231 (N_2231,N_1864,N_1745);
nand U2232 (N_2232,N_1742,N_1727);
nor U2233 (N_2233,N_1618,N_1859);
xor U2234 (N_2234,N_1930,N_1854);
nor U2235 (N_2235,N_1750,N_1677);
xnor U2236 (N_2236,N_1875,N_1525);
or U2237 (N_2237,N_1925,N_1895);
nor U2238 (N_2238,N_1675,N_1945);
nand U2239 (N_2239,N_1801,N_1892);
and U2240 (N_2240,N_1853,N_1726);
nor U2241 (N_2241,N_1509,N_1998);
nor U2242 (N_2242,N_1553,N_1889);
or U2243 (N_2243,N_1570,N_1724);
nor U2244 (N_2244,N_1514,N_1507);
and U2245 (N_2245,N_1633,N_1651);
nand U2246 (N_2246,N_1741,N_1838);
xor U2247 (N_2247,N_1985,N_1599);
nand U2248 (N_2248,N_1731,N_1996);
and U2249 (N_2249,N_1610,N_1959);
nor U2250 (N_2250,N_1981,N_1575);
or U2251 (N_2251,N_1789,N_1504);
or U2252 (N_2252,N_1913,N_1906);
xor U2253 (N_2253,N_1599,N_1663);
nand U2254 (N_2254,N_1703,N_1666);
nor U2255 (N_2255,N_1538,N_1638);
or U2256 (N_2256,N_1823,N_1767);
and U2257 (N_2257,N_1997,N_1697);
or U2258 (N_2258,N_1681,N_1758);
and U2259 (N_2259,N_1820,N_1800);
nand U2260 (N_2260,N_1941,N_1764);
xor U2261 (N_2261,N_1563,N_1788);
and U2262 (N_2262,N_1735,N_1903);
xor U2263 (N_2263,N_1586,N_1607);
or U2264 (N_2264,N_1539,N_1623);
xnor U2265 (N_2265,N_1919,N_1870);
nand U2266 (N_2266,N_1985,N_1929);
and U2267 (N_2267,N_1762,N_1970);
nand U2268 (N_2268,N_1873,N_1559);
and U2269 (N_2269,N_1548,N_1837);
xor U2270 (N_2270,N_1992,N_1942);
xor U2271 (N_2271,N_1761,N_1815);
or U2272 (N_2272,N_1649,N_1975);
and U2273 (N_2273,N_1521,N_1906);
or U2274 (N_2274,N_1964,N_1780);
nor U2275 (N_2275,N_1762,N_1655);
xnor U2276 (N_2276,N_1507,N_1622);
or U2277 (N_2277,N_1958,N_1826);
nand U2278 (N_2278,N_1975,N_1631);
nand U2279 (N_2279,N_1966,N_1754);
nand U2280 (N_2280,N_1642,N_1552);
or U2281 (N_2281,N_1692,N_1955);
or U2282 (N_2282,N_1903,N_1714);
xor U2283 (N_2283,N_1857,N_1763);
xnor U2284 (N_2284,N_1707,N_1534);
nor U2285 (N_2285,N_1833,N_1933);
or U2286 (N_2286,N_1740,N_1744);
or U2287 (N_2287,N_1605,N_1602);
and U2288 (N_2288,N_1684,N_1544);
nor U2289 (N_2289,N_1972,N_1549);
xor U2290 (N_2290,N_1782,N_1635);
or U2291 (N_2291,N_1734,N_1818);
nand U2292 (N_2292,N_1739,N_1583);
nor U2293 (N_2293,N_1855,N_1799);
nand U2294 (N_2294,N_1875,N_1943);
xor U2295 (N_2295,N_1562,N_1733);
xor U2296 (N_2296,N_1548,N_1598);
and U2297 (N_2297,N_1679,N_1894);
xnor U2298 (N_2298,N_1642,N_1503);
and U2299 (N_2299,N_1747,N_1799);
nand U2300 (N_2300,N_1714,N_1523);
nand U2301 (N_2301,N_1969,N_1771);
nand U2302 (N_2302,N_1807,N_1913);
or U2303 (N_2303,N_1549,N_1873);
nand U2304 (N_2304,N_1659,N_1960);
nor U2305 (N_2305,N_1711,N_1875);
nand U2306 (N_2306,N_1637,N_1885);
and U2307 (N_2307,N_1720,N_1646);
xor U2308 (N_2308,N_1664,N_1990);
nand U2309 (N_2309,N_1779,N_1880);
nand U2310 (N_2310,N_1894,N_1738);
and U2311 (N_2311,N_1714,N_1855);
nor U2312 (N_2312,N_1930,N_1945);
xnor U2313 (N_2313,N_1958,N_1976);
nand U2314 (N_2314,N_1617,N_1708);
nand U2315 (N_2315,N_1514,N_1970);
or U2316 (N_2316,N_1852,N_1543);
or U2317 (N_2317,N_1723,N_1676);
nor U2318 (N_2318,N_1625,N_1558);
xnor U2319 (N_2319,N_1817,N_1848);
nor U2320 (N_2320,N_1991,N_1529);
or U2321 (N_2321,N_1890,N_1883);
nand U2322 (N_2322,N_1577,N_1997);
nand U2323 (N_2323,N_1609,N_1619);
xor U2324 (N_2324,N_1614,N_1999);
xnor U2325 (N_2325,N_1580,N_1503);
nand U2326 (N_2326,N_1761,N_1683);
nor U2327 (N_2327,N_1563,N_1637);
and U2328 (N_2328,N_1541,N_1938);
or U2329 (N_2329,N_1665,N_1513);
or U2330 (N_2330,N_1706,N_1789);
nor U2331 (N_2331,N_1608,N_1638);
xnor U2332 (N_2332,N_1771,N_1534);
xnor U2333 (N_2333,N_1762,N_1605);
xnor U2334 (N_2334,N_1735,N_1984);
or U2335 (N_2335,N_1911,N_1945);
or U2336 (N_2336,N_1997,N_1803);
and U2337 (N_2337,N_1901,N_1951);
or U2338 (N_2338,N_1933,N_1616);
nand U2339 (N_2339,N_1630,N_1639);
or U2340 (N_2340,N_1529,N_1976);
nand U2341 (N_2341,N_1503,N_1707);
xor U2342 (N_2342,N_1878,N_1975);
nor U2343 (N_2343,N_1771,N_1736);
xnor U2344 (N_2344,N_1824,N_1559);
xnor U2345 (N_2345,N_1543,N_1525);
xor U2346 (N_2346,N_1769,N_1654);
or U2347 (N_2347,N_1528,N_1740);
nor U2348 (N_2348,N_1873,N_1646);
xor U2349 (N_2349,N_1970,N_1609);
xor U2350 (N_2350,N_1857,N_1684);
nor U2351 (N_2351,N_1770,N_1504);
xnor U2352 (N_2352,N_1664,N_1851);
nor U2353 (N_2353,N_1537,N_1784);
and U2354 (N_2354,N_1761,N_1992);
nand U2355 (N_2355,N_1920,N_1810);
nor U2356 (N_2356,N_1508,N_1702);
and U2357 (N_2357,N_1769,N_1722);
nand U2358 (N_2358,N_1780,N_1868);
nand U2359 (N_2359,N_1896,N_1944);
nand U2360 (N_2360,N_1938,N_1638);
nand U2361 (N_2361,N_1929,N_1731);
nor U2362 (N_2362,N_1718,N_1775);
and U2363 (N_2363,N_1593,N_1644);
nor U2364 (N_2364,N_1652,N_1616);
nor U2365 (N_2365,N_1850,N_1946);
xnor U2366 (N_2366,N_1756,N_1512);
nor U2367 (N_2367,N_1937,N_1524);
xnor U2368 (N_2368,N_1501,N_1733);
nor U2369 (N_2369,N_1563,N_1975);
and U2370 (N_2370,N_1516,N_1579);
or U2371 (N_2371,N_1845,N_1738);
nand U2372 (N_2372,N_1736,N_1582);
or U2373 (N_2373,N_1555,N_1631);
xor U2374 (N_2374,N_1666,N_1630);
xor U2375 (N_2375,N_1545,N_1606);
and U2376 (N_2376,N_1681,N_1633);
nand U2377 (N_2377,N_1856,N_1715);
or U2378 (N_2378,N_1996,N_1854);
or U2379 (N_2379,N_1719,N_1885);
nand U2380 (N_2380,N_1744,N_1915);
and U2381 (N_2381,N_1556,N_1974);
nor U2382 (N_2382,N_1948,N_1533);
or U2383 (N_2383,N_1888,N_1705);
and U2384 (N_2384,N_1581,N_1968);
and U2385 (N_2385,N_1725,N_1689);
or U2386 (N_2386,N_1902,N_1958);
or U2387 (N_2387,N_1740,N_1713);
and U2388 (N_2388,N_1692,N_1738);
nand U2389 (N_2389,N_1870,N_1845);
nand U2390 (N_2390,N_1964,N_1981);
and U2391 (N_2391,N_1680,N_1840);
or U2392 (N_2392,N_1555,N_1637);
nor U2393 (N_2393,N_1995,N_1712);
nor U2394 (N_2394,N_1991,N_1981);
nor U2395 (N_2395,N_1948,N_1596);
and U2396 (N_2396,N_1553,N_1609);
nor U2397 (N_2397,N_1710,N_1810);
nand U2398 (N_2398,N_1830,N_1540);
and U2399 (N_2399,N_1747,N_1505);
nand U2400 (N_2400,N_1933,N_1969);
nor U2401 (N_2401,N_1600,N_1897);
nor U2402 (N_2402,N_1748,N_1885);
xnor U2403 (N_2403,N_1510,N_1519);
and U2404 (N_2404,N_1759,N_1740);
or U2405 (N_2405,N_1729,N_1978);
and U2406 (N_2406,N_1863,N_1921);
nor U2407 (N_2407,N_1881,N_1615);
nand U2408 (N_2408,N_1860,N_1846);
and U2409 (N_2409,N_1540,N_1785);
or U2410 (N_2410,N_1576,N_1554);
nor U2411 (N_2411,N_1708,N_1666);
and U2412 (N_2412,N_1639,N_1930);
xnor U2413 (N_2413,N_1694,N_1757);
nand U2414 (N_2414,N_1574,N_1501);
nor U2415 (N_2415,N_1733,N_1675);
nand U2416 (N_2416,N_1822,N_1924);
or U2417 (N_2417,N_1573,N_1956);
or U2418 (N_2418,N_1814,N_1619);
nor U2419 (N_2419,N_1667,N_1989);
nand U2420 (N_2420,N_1533,N_1659);
nand U2421 (N_2421,N_1673,N_1961);
nor U2422 (N_2422,N_1503,N_1636);
or U2423 (N_2423,N_1562,N_1756);
nor U2424 (N_2424,N_1733,N_1784);
and U2425 (N_2425,N_1674,N_1833);
nand U2426 (N_2426,N_1557,N_1897);
and U2427 (N_2427,N_1812,N_1959);
and U2428 (N_2428,N_1555,N_1886);
and U2429 (N_2429,N_1992,N_1581);
or U2430 (N_2430,N_1808,N_1600);
or U2431 (N_2431,N_1608,N_1520);
nand U2432 (N_2432,N_1807,N_1646);
xor U2433 (N_2433,N_1672,N_1938);
or U2434 (N_2434,N_1927,N_1747);
xor U2435 (N_2435,N_1844,N_1738);
xnor U2436 (N_2436,N_1684,N_1998);
and U2437 (N_2437,N_1737,N_1778);
nor U2438 (N_2438,N_1887,N_1735);
xor U2439 (N_2439,N_1999,N_1924);
xor U2440 (N_2440,N_1946,N_1657);
nand U2441 (N_2441,N_1784,N_1813);
nand U2442 (N_2442,N_1733,N_1974);
xnor U2443 (N_2443,N_1546,N_1783);
nor U2444 (N_2444,N_1598,N_1794);
and U2445 (N_2445,N_1589,N_1809);
or U2446 (N_2446,N_1760,N_1587);
nor U2447 (N_2447,N_1820,N_1547);
or U2448 (N_2448,N_1773,N_1704);
xor U2449 (N_2449,N_1895,N_1719);
nor U2450 (N_2450,N_1876,N_1915);
nor U2451 (N_2451,N_1608,N_1800);
and U2452 (N_2452,N_1710,N_1532);
xor U2453 (N_2453,N_1902,N_1510);
nand U2454 (N_2454,N_1747,N_1568);
nor U2455 (N_2455,N_1641,N_1690);
nor U2456 (N_2456,N_1965,N_1871);
xor U2457 (N_2457,N_1680,N_1799);
or U2458 (N_2458,N_1968,N_1930);
nor U2459 (N_2459,N_1591,N_1835);
nand U2460 (N_2460,N_1825,N_1763);
xnor U2461 (N_2461,N_1546,N_1743);
xnor U2462 (N_2462,N_1697,N_1910);
xnor U2463 (N_2463,N_1750,N_1715);
and U2464 (N_2464,N_1566,N_1912);
nand U2465 (N_2465,N_1999,N_1708);
xnor U2466 (N_2466,N_1572,N_1929);
and U2467 (N_2467,N_1998,N_1544);
and U2468 (N_2468,N_1524,N_1538);
and U2469 (N_2469,N_1798,N_1574);
and U2470 (N_2470,N_1847,N_1631);
nand U2471 (N_2471,N_1527,N_1931);
xnor U2472 (N_2472,N_1687,N_1809);
and U2473 (N_2473,N_1996,N_1511);
and U2474 (N_2474,N_1770,N_1945);
nand U2475 (N_2475,N_1972,N_1934);
and U2476 (N_2476,N_1993,N_1597);
nor U2477 (N_2477,N_1872,N_1860);
nand U2478 (N_2478,N_1681,N_1938);
and U2479 (N_2479,N_1863,N_1650);
nand U2480 (N_2480,N_1617,N_1715);
and U2481 (N_2481,N_1842,N_1649);
xor U2482 (N_2482,N_1530,N_1660);
nor U2483 (N_2483,N_1877,N_1648);
xnor U2484 (N_2484,N_1509,N_1992);
or U2485 (N_2485,N_1809,N_1591);
or U2486 (N_2486,N_1860,N_1819);
nor U2487 (N_2487,N_1724,N_1978);
nor U2488 (N_2488,N_1968,N_1607);
nand U2489 (N_2489,N_1779,N_1600);
and U2490 (N_2490,N_1893,N_1842);
xnor U2491 (N_2491,N_1849,N_1921);
or U2492 (N_2492,N_1660,N_1928);
nor U2493 (N_2493,N_1747,N_1680);
nor U2494 (N_2494,N_1546,N_1708);
nand U2495 (N_2495,N_1720,N_1548);
xnor U2496 (N_2496,N_1670,N_1845);
xnor U2497 (N_2497,N_1673,N_1908);
xnor U2498 (N_2498,N_1760,N_1740);
nand U2499 (N_2499,N_1683,N_1835);
xor U2500 (N_2500,N_2091,N_2296);
and U2501 (N_2501,N_2099,N_2057);
nor U2502 (N_2502,N_2050,N_2216);
nand U2503 (N_2503,N_2171,N_2055);
xnor U2504 (N_2504,N_2108,N_2426);
or U2505 (N_2505,N_2373,N_2226);
and U2506 (N_2506,N_2053,N_2397);
nor U2507 (N_2507,N_2051,N_2147);
nor U2508 (N_2508,N_2123,N_2459);
xor U2509 (N_2509,N_2469,N_2046);
xnor U2510 (N_2510,N_2014,N_2101);
and U2511 (N_2511,N_2346,N_2180);
xor U2512 (N_2512,N_2305,N_2234);
xor U2513 (N_2513,N_2339,N_2256);
nor U2514 (N_2514,N_2075,N_2432);
or U2515 (N_2515,N_2009,N_2270);
and U2516 (N_2516,N_2220,N_2472);
and U2517 (N_2517,N_2263,N_2487);
xor U2518 (N_2518,N_2241,N_2463);
nor U2519 (N_2519,N_2295,N_2258);
or U2520 (N_2520,N_2284,N_2303);
or U2521 (N_2521,N_2213,N_2079);
nor U2522 (N_2522,N_2315,N_2273);
and U2523 (N_2523,N_2011,N_2097);
nor U2524 (N_2524,N_2290,N_2034);
nand U2525 (N_2525,N_2347,N_2370);
xnor U2526 (N_2526,N_2000,N_2435);
nor U2527 (N_2527,N_2385,N_2194);
nand U2528 (N_2528,N_2423,N_2403);
or U2529 (N_2529,N_2132,N_2280);
or U2530 (N_2530,N_2161,N_2054);
nor U2531 (N_2531,N_2490,N_2390);
xor U2532 (N_2532,N_2479,N_2340);
and U2533 (N_2533,N_2449,N_2279);
nor U2534 (N_2534,N_2417,N_2369);
or U2535 (N_2535,N_2088,N_2229);
xor U2536 (N_2536,N_2165,N_2387);
nand U2537 (N_2537,N_2059,N_2382);
and U2538 (N_2538,N_2041,N_2440);
or U2539 (N_2539,N_2355,N_2453);
or U2540 (N_2540,N_2249,N_2411);
or U2541 (N_2541,N_2089,N_2248);
nand U2542 (N_2542,N_2441,N_2211);
nand U2543 (N_2543,N_2391,N_2413);
xor U2544 (N_2544,N_2062,N_2306);
or U2545 (N_2545,N_2086,N_2364);
xor U2546 (N_2546,N_2465,N_2321);
and U2547 (N_2547,N_2473,N_2230);
xor U2548 (N_2548,N_2257,N_2228);
nor U2549 (N_2549,N_2483,N_2087);
or U2550 (N_2550,N_2071,N_2264);
xnor U2551 (N_2551,N_2478,N_2033);
nor U2552 (N_2552,N_2204,N_2004);
xor U2553 (N_2553,N_2095,N_2322);
or U2554 (N_2554,N_2304,N_2218);
nor U2555 (N_2555,N_2197,N_2145);
nand U2556 (N_2556,N_2060,N_2177);
nor U2557 (N_2557,N_2259,N_2386);
nand U2558 (N_2558,N_2358,N_2098);
nand U2559 (N_2559,N_2252,N_2024);
and U2560 (N_2560,N_2193,N_2327);
or U2561 (N_2561,N_2038,N_2462);
nand U2562 (N_2562,N_2470,N_2117);
and U2563 (N_2563,N_2126,N_2400);
nand U2564 (N_2564,N_2082,N_2238);
nor U2565 (N_2565,N_2410,N_2100);
or U2566 (N_2566,N_2113,N_2496);
xnor U2567 (N_2567,N_2210,N_2481);
xnor U2568 (N_2568,N_2162,N_2081);
or U2569 (N_2569,N_2439,N_2337);
or U2570 (N_2570,N_2170,N_2294);
nand U2571 (N_2571,N_2227,N_2124);
and U2572 (N_2572,N_2302,N_2148);
and U2573 (N_2573,N_2277,N_2104);
nand U2574 (N_2574,N_2319,N_2452);
nor U2575 (N_2575,N_2458,N_2128);
nand U2576 (N_2576,N_2408,N_2242);
and U2577 (N_2577,N_2331,N_2077);
xor U2578 (N_2578,N_2299,N_2292);
xor U2579 (N_2579,N_2395,N_2007);
xor U2580 (N_2580,N_2336,N_2010);
xor U2581 (N_2581,N_2187,N_2027);
nand U2582 (N_2582,N_2414,N_2291);
nor U2583 (N_2583,N_2419,N_2129);
or U2584 (N_2584,N_2489,N_2484);
or U2585 (N_2585,N_2298,N_2085);
or U2586 (N_2586,N_2164,N_2118);
or U2587 (N_2587,N_2399,N_2184);
and U2588 (N_2588,N_2112,N_2495);
or U2589 (N_2589,N_2130,N_2047);
xnor U2590 (N_2590,N_2313,N_2188);
nor U2591 (N_2591,N_2486,N_2061);
nand U2592 (N_2592,N_2428,N_2335);
and U2593 (N_2593,N_2325,N_2246);
or U2594 (N_2594,N_2389,N_2032);
xor U2595 (N_2595,N_2182,N_2398);
or U2596 (N_2596,N_2353,N_2328);
xnor U2597 (N_2597,N_2392,N_2239);
and U2598 (N_2598,N_2151,N_2172);
and U2599 (N_2599,N_2157,N_2377);
nor U2600 (N_2600,N_2155,N_2365);
and U2601 (N_2601,N_2424,N_2283);
or U2602 (N_2602,N_2267,N_2438);
nor U2603 (N_2603,N_2429,N_2437);
or U2604 (N_2604,N_2378,N_2198);
and U2605 (N_2605,N_2203,N_2471);
nand U2606 (N_2606,N_2348,N_2135);
xnor U2607 (N_2607,N_2492,N_2013);
xor U2608 (N_2608,N_2497,N_2351);
nor U2609 (N_2609,N_2311,N_2425);
and U2610 (N_2610,N_2368,N_2448);
xor U2611 (N_2611,N_2214,N_2396);
xor U2612 (N_2612,N_2276,N_2111);
nor U2613 (N_2613,N_2317,N_2116);
nand U2614 (N_2614,N_2215,N_2225);
or U2615 (N_2615,N_2043,N_2427);
nand U2616 (N_2616,N_2195,N_2064);
nor U2617 (N_2617,N_2431,N_2454);
or U2618 (N_2618,N_2375,N_2201);
nand U2619 (N_2619,N_2312,N_2205);
xnor U2620 (N_2620,N_2360,N_2045);
nand U2621 (N_2621,N_2329,N_2156);
nor U2622 (N_2622,N_2153,N_2036);
nor U2623 (N_2623,N_2342,N_2106);
xnor U2624 (N_2624,N_2464,N_2192);
xor U2625 (N_2625,N_2323,N_2207);
or U2626 (N_2626,N_2443,N_2015);
nor U2627 (N_2627,N_2002,N_2048);
xnor U2628 (N_2628,N_2115,N_2405);
xor U2629 (N_2629,N_2480,N_2093);
xnor U2630 (N_2630,N_2208,N_2003);
nor U2631 (N_2631,N_2488,N_2404);
xnor U2632 (N_2632,N_2200,N_2016);
nor U2633 (N_2633,N_2407,N_2185);
nand U2634 (N_2634,N_2149,N_2297);
and U2635 (N_2635,N_2065,N_2401);
or U2636 (N_2636,N_2455,N_2447);
and U2637 (N_2637,N_2056,N_2212);
nor U2638 (N_2638,N_2160,N_2028);
nand U2639 (N_2639,N_2006,N_2159);
nor U2640 (N_2640,N_2309,N_2072);
xnor U2641 (N_2641,N_2076,N_2467);
nand U2642 (N_2642,N_2272,N_2493);
nor U2643 (N_2643,N_2314,N_2120);
xnor U2644 (N_2644,N_2236,N_2107);
xor U2645 (N_2645,N_2243,N_2476);
nor U2646 (N_2646,N_2363,N_2466);
and U2647 (N_2647,N_2144,N_2436);
and U2648 (N_2648,N_2183,N_2025);
xor U2649 (N_2649,N_2357,N_2012);
or U2650 (N_2650,N_2231,N_2078);
or U2651 (N_2651,N_2285,N_2301);
nand U2652 (N_2652,N_2334,N_2268);
and U2653 (N_2653,N_2444,N_2475);
xnor U2654 (N_2654,N_2154,N_2163);
nand U2655 (N_2655,N_2372,N_2219);
or U2656 (N_2656,N_2402,N_2199);
nand U2657 (N_2657,N_2103,N_2450);
or U2658 (N_2658,N_2482,N_2167);
and U2659 (N_2659,N_2412,N_2260);
nand U2660 (N_2660,N_2232,N_2173);
nor U2661 (N_2661,N_2451,N_2430);
xor U2662 (N_2662,N_2359,N_2371);
xor U2663 (N_2663,N_2066,N_2023);
nand U2664 (N_2664,N_2031,N_2383);
nor U2665 (N_2665,N_2109,N_2131);
nand U2666 (N_2666,N_2376,N_2247);
xor U2667 (N_2667,N_2029,N_2019);
nor U2668 (N_2668,N_2421,N_2384);
nor U2669 (N_2669,N_2265,N_2068);
nor U2670 (N_2670,N_2141,N_2017);
or U2671 (N_2671,N_2189,N_2158);
and U2672 (N_2672,N_2244,N_2084);
and U2673 (N_2673,N_2393,N_2001);
and U2674 (N_2674,N_2253,N_2310);
or U2675 (N_2675,N_2381,N_2461);
xor U2676 (N_2676,N_2394,N_2022);
nor U2677 (N_2677,N_2042,N_2251);
nor U2678 (N_2678,N_2380,N_2350);
xnor U2679 (N_2679,N_2491,N_2224);
xnor U2680 (N_2680,N_2138,N_2121);
nand U2681 (N_2681,N_2422,N_2318);
or U2682 (N_2682,N_2221,N_2166);
nand U2683 (N_2683,N_2030,N_2102);
nand U2684 (N_2684,N_2049,N_2237);
nand U2685 (N_2685,N_2275,N_2456);
xor U2686 (N_2686,N_2361,N_2110);
nand U2687 (N_2687,N_2070,N_2067);
or U2688 (N_2688,N_2320,N_2286);
and U2689 (N_2689,N_2352,N_2498);
xnor U2690 (N_2690,N_2343,N_2287);
nor U2691 (N_2691,N_2345,N_2191);
xor U2692 (N_2692,N_2152,N_2460);
nand U2693 (N_2693,N_2209,N_2005);
xnor U2694 (N_2694,N_2338,N_2434);
nand U2695 (N_2695,N_2196,N_2125);
nor U2696 (N_2696,N_2494,N_2416);
nor U2697 (N_2697,N_2142,N_2037);
and U2698 (N_2698,N_2474,N_2039);
and U2699 (N_2699,N_2094,N_2250);
nor U2700 (N_2700,N_2245,N_2262);
or U2701 (N_2701,N_2308,N_2271);
nand U2702 (N_2702,N_2418,N_2119);
and U2703 (N_2703,N_2114,N_2134);
or U2704 (N_2704,N_2136,N_2040);
xor U2705 (N_2705,N_2074,N_2235);
and U2706 (N_2706,N_2388,N_2058);
nor U2707 (N_2707,N_2445,N_2362);
or U2708 (N_2708,N_2176,N_2333);
and U2709 (N_2709,N_2477,N_2442);
xnor U2710 (N_2710,N_2332,N_2137);
xor U2711 (N_2711,N_2330,N_2433);
xnor U2712 (N_2712,N_2181,N_2190);
nand U2713 (N_2713,N_2052,N_2139);
and U2714 (N_2714,N_2300,N_2288);
nand U2715 (N_2715,N_2096,N_2293);
nand U2716 (N_2716,N_2069,N_2354);
or U2717 (N_2717,N_2026,N_2008);
nand U2718 (N_2718,N_2083,N_2090);
xor U2719 (N_2719,N_2341,N_2063);
nand U2720 (N_2720,N_2240,N_2092);
xor U2721 (N_2721,N_2222,N_2140);
xor U2722 (N_2722,N_2326,N_2186);
and U2723 (N_2723,N_2217,N_2420);
nor U2724 (N_2724,N_2020,N_2168);
nor U2725 (N_2725,N_2374,N_2178);
and U2726 (N_2726,N_2274,N_2344);
xnor U2727 (N_2727,N_2366,N_2266);
xnor U2728 (N_2728,N_2018,N_2406);
nand U2729 (N_2729,N_2261,N_2133);
nor U2730 (N_2730,N_2324,N_2021);
xnor U2731 (N_2731,N_2179,N_2356);
xor U2732 (N_2732,N_2409,N_2206);
xor U2733 (N_2733,N_2143,N_2499);
nor U2734 (N_2734,N_2073,N_2278);
xnor U2735 (N_2735,N_2146,N_2367);
nor U2736 (N_2736,N_2127,N_2468);
xor U2737 (N_2737,N_2269,N_2415);
nor U2738 (N_2738,N_2379,N_2457);
or U2739 (N_2739,N_2349,N_2175);
xor U2740 (N_2740,N_2255,N_2150);
and U2741 (N_2741,N_2174,N_2316);
nand U2742 (N_2742,N_2169,N_2080);
nand U2743 (N_2743,N_2044,N_2223);
nor U2744 (N_2744,N_2202,N_2485);
xnor U2745 (N_2745,N_2282,N_2446);
nand U2746 (N_2746,N_2307,N_2281);
nand U2747 (N_2747,N_2035,N_2289);
nand U2748 (N_2748,N_2122,N_2254);
nor U2749 (N_2749,N_2233,N_2105);
or U2750 (N_2750,N_2283,N_2066);
nor U2751 (N_2751,N_2118,N_2385);
nor U2752 (N_2752,N_2235,N_2183);
or U2753 (N_2753,N_2456,N_2382);
xnor U2754 (N_2754,N_2216,N_2157);
xnor U2755 (N_2755,N_2433,N_2274);
or U2756 (N_2756,N_2303,N_2125);
xnor U2757 (N_2757,N_2155,N_2213);
nand U2758 (N_2758,N_2278,N_2248);
nor U2759 (N_2759,N_2093,N_2412);
xnor U2760 (N_2760,N_2405,N_2315);
or U2761 (N_2761,N_2343,N_2293);
or U2762 (N_2762,N_2017,N_2380);
or U2763 (N_2763,N_2334,N_2477);
nor U2764 (N_2764,N_2456,N_2175);
xor U2765 (N_2765,N_2144,N_2210);
xnor U2766 (N_2766,N_2108,N_2179);
xnor U2767 (N_2767,N_2279,N_2322);
nor U2768 (N_2768,N_2481,N_2114);
nor U2769 (N_2769,N_2398,N_2233);
nand U2770 (N_2770,N_2140,N_2274);
or U2771 (N_2771,N_2311,N_2286);
nand U2772 (N_2772,N_2021,N_2042);
xnor U2773 (N_2773,N_2096,N_2267);
or U2774 (N_2774,N_2028,N_2427);
nand U2775 (N_2775,N_2326,N_2429);
nor U2776 (N_2776,N_2310,N_2149);
and U2777 (N_2777,N_2358,N_2486);
nor U2778 (N_2778,N_2170,N_2061);
xnor U2779 (N_2779,N_2437,N_2385);
nor U2780 (N_2780,N_2034,N_2404);
and U2781 (N_2781,N_2167,N_2389);
and U2782 (N_2782,N_2435,N_2089);
or U2783 (N_2783,N_2291,N_2429);
nor U2784 (N_2784,N_2092,N_2099);
nor U2785 (N_2785,N_2149,N_2262);
and U2786 (N_2786,N_2207,N_2132);
or U2787 (N_2787,N_2494,N_2411);
nand U2788 (N_2788,N_2200,N_2017);
or U2789 (N_2789,N_2450,N_2388);
nor U2790 (N_2790,N_2427,N_2384);
xor U2791 (N_2791,N_2285,N_2372);
or U2792 (N_2792,N_2068,N_2319);
nor U2793 (N_2793,N_2465,N_2337);
nor U2794 (N_2794,N_2410,N_2248);
and U2795 (N_2795,N_2103,N_2264);
nor U2796 (N_2796,N_2327,N_2225);
nand U2797 (N_2797,N_2054,N_2135);
and U2798 (N_2798,N_2462,N_2308);
nand U2799 (N_2799,N_2250,N_2137);
nand U2800 (N_2800,N_2096,N_2440);
nand U2801 (N_2801,N_2185,N_2400);
and U2802 (N_2802,N_2258,N_2067);
nor U2803 (N_2803,N_2261,N_2126);
nor U2804 (N_2804,N_2242,N_2114);
nand U2805 (N_2805,N_2079,N_2123);
nand U2806 (N_2806,N_2481,N_2107);
nor U2807 (N_2807,N_2387,N_2246);
nor U2808 (N_2808,N_2001,N_2491);
and U2809 (N_2809,N_2469,N_2077);
or U2810 (N_2810,N_2154,N_2247);
nand U2811 (N_2811,N_2289,N_2224);
or U2812 (N_2812,N_2066,N_2429);
and U2813 (N_2813,N_2360,N_2186);
xnor U2814 (N_2814,N_2356,N_2374);
or U2815 (N_2815,N_2316,N_2295);
xnor U2816 (N_2816,N_2014,N_2389);
xnor U2817 (N_2817,N_2419,N_2491);
nor U2818 (N_2818,N_2338,N_2222);
and U2819 (N_2819,N_2067,N_2205);
or U2820 (N_2820,N_2293,N_2024);
xor U2821 (N_2821,N_2248,N_2116);
nand U2822 (N_2822,N_2473,N_2175);
or U2823 (N_2823,N_2477,N_2232);
and U2824 (N_2824,N_2127,N_2383);
xor U2825 (N_2825,N_2337,N_2043);
xnor U2826 (N_2826,N_2212,N_2301);
and U2827 (N_2827,N_2319,N_2386);
and U2828 (N_2828,N_2470,N_2184);
xnor U2829 (N_2829,N_2463,N_2069);
nor U2830 (N_2830,N_2230,N_2170);
nor U2831 (N_2831,N_2457,N_2450);
nor U2832 (N_2832,N_2498,N_2075);
nand U2833 (N_2833,N_2079,N_2149);
nand U2834 (N_2834,N_2492,N_2220);
xor U2835 (N_2835,N_2355,N_2255);
and U2836 (N_2836,N_2220,N_2306);
nand U2837 (N_2837,N_2402,N_2461);
nand U2838 (N_2838,N_2329,N_2361);
and U2839 (N_2839,N_2271,N_2052);
and U2840 (N_2840,N_2323,N_2171);
nand U2841 (N_2841,N_2086,N_2336);
or U2842 (N_2842,N_2301,N_2062);
nand U2843 (N_2843,N_2435,N_2377);
and U2844 (N_2844,N_2263,N_2215);
xor U2845 (N_2845,N_2319,N_2342);
and U2846 (N_2846,N_2494,N_2076);
or U2847 (N_2847,N_2122,N_2233);
nor U2848 (N_2848,N_2060,N_2446);
xnor U2849 (N_2849,N_2350,N_2412);
nand U2850 (N_2850,N_2330,N_2412);
nor U2851 (N_2851,N_2338,N_2417);
nand U2852 (N_2852,N_2039,N_2192);
nor U2853 (N_2853,N_2012,N_2024);
nor U2854 (N_2854,N_2360,N_2334);
or U2855 (N_2855,N_2026,N_2432);
nor U2856 (N_2856,N_2016,N_2479);
and U2857 (N_2857,N_2452,N_2314);
xnor U2858 (N_2858,N_2146,N_2426);
or U2859 (N_2859,N_2484,N_2032);
nand U2860 (N_2860,N_2472,N_2348);
xor U2861 (N_2861,N_2198,N_2329);
nor U2862 (N_2862,N_2035,N_2371);
nor U2863 (N_2863,N_2182,N_2051);
and U2864 (N_2864,N_2239,N_2435);
or U2865 (N_2865,N_2179,N_2358);
and U2866 (N_2866,N_2389,N_2058);
nand U2867 (N_2867,N_2089,N_2013);
nand U2868 (N_2868,N_2099,N_2334);
nor U2869 (N_2869,N_2049,N_2184);
or U2870 (N_2870,N_2411,N_2389);
nand U2871 (N_2871,N_2135,N_2396);
and U2872 (N_2872,N_2226,N_2140);
or U2873 (N_2873,N_2388,N_2069);
nand U2874 (N_2874,N_2268,N_2353);
or U2875 (N_2875,N_2423,N_2127);
nand U2876 (N_2876,N_2165,N_2310);
nor U2877 (N_2877,N_2396,N_2334);
nand U2878 (N_2878,N_2319,N_2113);
xor U2879 (N_2879,N_2458,N_2066);
nor U2880 (N_2880,N_2108,N_2243);
nand U2881 (N_2881,N_2345,N_2103);
nand U2882 (N_2882,N_2197,N_2479);
and U2883 (N_2883,N_2070,N_2421);
and U2884 (N_2884,N_2345,N_2173);
nor U2885 (N_2885,N_2335,N_2458);
or U2886 (N_2886,N_2039,N_2178);
or U2887 (N_2887,N_2399,N_2459);
nand U2888 (N_2888,N_2316,N_2313);
xor U2889 (N_2889,N_2044,N_2227);
or U2890 (N_2890,N_2177,N_2479);
nor U2891 (N_2891,N_2155,N_2075);
and U2892 (N_2892,N_2053,N_2238);
xnor U2893 (N_2893,N_2459,N_2386);
xor U2894 (N_2894,N_2419,N_2189);
xor U2895 (N_2895,N_2414,N_2028);
nor U2896 (N_2896,N_2303,N_2450);
xnor U2897 (N_2897,N_2228,N_2283);
nor U2898 (N_2898,N_2026,N_2130);
and U2899 (N_2899,N_2146,N_2263);
nor U2900 (N_2900,N_2005,N_2301);
nand U2901 (N_2901,N_2492,N_2352);
nor U2902 (N_2902,N_2219,N_2381);
and U2903 (N_2903,N_2019,N_2142);
nor U2904 (N_2904,N_2471,N_2321);
nor U2905 (N_2905,N_2263,N_2470);
nor U2906 (N_2906,N_2226,N_2344);
xnor U2907 (N_2907,N_2237,N_2181);
and U2908 (N_2908,N_2459,N_2367);
or U2909 (N_2909,N_2215,N_2184);
and U2910 (N_2910,N_2078,N_2323);
and U2911 (N_2911,N_2217,N_2045);
nor U2912 (N_2912,N_2144,N_2165);
xnor U2913 (N_2913,N_2233,N_2474);
nor U2914 (N_2914,N_2050,N_2063);
or U2915 (N_2915,N_2034,N_2183);
nand U2916 (N_2916,N_2241,N_2123);
and U2917 (N_2917,N_2105,N_2023);
nand U2918 (N_2918,N_2362,N_2316);
and U2919 (N_2919,N_2325,N_2186);
nand U2920 (N_2920,N_2270,N_2360);
xnor U2921 (N_2921,N_2196,N_2188);
and U2922 (N_2922,N_2008,N_2151);
or U2923 (N_2923,N_2304,N_2308);
and U2924 (N_2924,N_2350,N_2455);
xor U2925 (N_2925,N_2271,N_2253);
or U2926 (N_2926,N_2026,N_2218);
or U2927 (N_2927,N_2174,N_2220);
nand U2928 (N_2928,N_2060,N_2144);
xnor U2929 (N_2929,N_2305,N_2122);
and U2930 (N_2930,N_2284,N_2280);
nor U2931 (N_2931,N_2421,N_2148);
nor U2932 (N_2932,N_2098,N_2229);
nor U2933 (N_2933,N_2295,N_2417);
nor U2934 (N_2934,N_2055,N_2473);
or U2935 (N_2935,N_2092,N_2292);
nand U2936 (N_2936,N_2439,N_2177);
nand U2937 (N_2937,N_2348,N_2496);
nor U2938 (N_2938,N_2023,N_2309);
nor U2939 (N_2939,N_2224,N_2364);
xor U2940 (N_2940,N_2045,N_2258);
nor U2941 (N_2941,N_2368,N_2013);
and U2942 (N_2942,N_2017,N_2245);
and U2943 (N_2943,N_2488,N_2346);
nand U2944 (N_2944,N_2073,N_2107);
or U2945 (N_2945,N_2006,N_2177);
xnor U2946 (N_2946,N_2279,N_2492);
and U2947 (N_2947,N_2421,N_2052);
nor U2948 (N_2948,N_2474,N_2271);
nand U2949 (N_2949,N_2294,N_2196);
or U2950 (N_2950,N_2309,N_2490);
or U2951 (N_2951,N_2139,N_2022);
xnor U2952 (N_2952,N_2058,N_2274);
xnor U2953 (N_2953,N_2038,N_2384);
nand U2954 (N_2954,N_2020,N_2017);
or U2955 (N_2955,N_2058,N_2320);
xor U2956 (N_2956,N_2364,N_2488);
and U2957 (N_2957,N_2231,N_2286);
or U2958 (N_2958,N_2211,N_2141);
or U2959 (N_2959,N_2176,N_2369);
nor U2960 (N_2960,N_2190,N_2255);
xor U2961 (N_2961,N_2145,N_2417);
xor U2962 (N_2962,N_2171,N_2363);
nor U2963 (N_2963,N_2400,N_2267);
xnor U2964 (N_2964,N_2045,N_2146);
and U2965 (N_2965,N_2258,N_2288);
or U2966 (N_2966,N_2203,N_2007);
nand U2967 (N_2967,N_2438,N_2204);
nor U2968 (N_2968,N_2173,N_2168);
nor U2969 (N_2969,N_2140,N_2026);
nand U2970 (N_2970,N_2384,N_2255);
nand U2971 (N_2971,N_2105,N_2261);
or U2972 (N_2972,N_2486,N_2215);
and U2973 (N_2973,N_2378,N_2264);
xor U2974 (N_2974,N_2294,N_2334);
xnor U2975 (N_2975,N_2331,N_2248);
and U2976 (N_2976,N_2139,N_2468);
nor U2977 (N_2977,N_2469,N_2348);
nand U2978 (N_2978,N_2440,N_2100);
nor U2979 (N_2979,N_2166,N_2052);
or U2980 (N_2980,N_2103,N_2406);
xnor U2981 (N_2981,N_2234,N_2471);
nor U2982 (N_2982,N_2192,N_2125);
nor U2983 (N_2983,N_2322,N_2498);
nor U2984 (N_2984,N_2299,N_2206);
nor U2985 (N_2985,N_2408,N_2004);
and U2986 (N_2986,N_2050,N_2406);
xor U2987 (N_2987,N_2032,N_2357);
xor U2988 (N_2988,N_2014,N_2254);
xnor U2989 (N_2989,N_2311,N_2012);
or U2990 (N_2990,N_2139,N_2136);
nand U2991 (N_2991,N_2112,N_2357);
nand U2992 (N_2992,N_2359,N_2162);
and U2993 (N_2993,N_2428,N_2078);
nand U2994 (N_2994,N_2305,N_2430);
xor U2995 (N_2995,N_2065,N_2453);
nand U2996 (N_2996,N_2360,N_2399);
nand U2997 (N_2997,N_2061,N_2146);
and U2998 (N_2998,N_2155,N_2042);
and U2999 (N_2999,N_2195,N_2048);
nor U3000 (N_3000,N_2669,N_2635);
or U3001 (N_3001,N_2756,N_2911);
and U3002 (N_3002,N_2801,N_2976);
or U3003 (N_3003,N_2685,N_2691);
xnor U3004 (N_3004,N_2968,N_2858);
xnor U3005 (N_3005,N_2663,N_2649);
nand U3006 (N_3006,N_2792,N_2793);
xnor U3007 (N_3007,N_2738,N_2974);
nand U3008 (N_3008,N_2782,N_2903);
and U3009 (N_3009,N_2621,N_2596);
or U3010 (N_3010,N_2712,N_2764);
or U3011 (N_3011,N_2655,N_2749);
xnor U3012 (N_3012,N_2671,N_2996);
nor U3013 (N_3013,N_2560,N_2571);
xnor U3014 (N_3014,N_2570,N_2926);
and U3015 (N_3015,N_2753,N_2931);
xnor U3016 (N_3016,N_2653,N_2638);
and U3017 (N_3017,N_2529,N_2746);
or U3018 (N_3018,N_2766,N_2802);
nand U3019 (N_3019,N_2803,N_2696);
nand U3020 (N_3020,N_2535,N_2847);
xnor U3021 (N_3021,N_2886,N_2841);
nand U3022 (N_3022,N_2779,N_2948);
or U3023 (N_3023,N_2845,N_2634);
nor U3024 (N_3024,N_2999,N_2618);
and U3025 (N_3025,N_2904,N_2693);
nand U3026 (N_3026,N_2787,N_2918);
and U3027 (N_3027,N_2657,N_2942);
or U3028 (N_3028,N_2966,N_2615);
nand U3029 (N_3029,N_2688,N_2599);
and U3030 (N_3030,N_2923,N_2833);
nand U3031 (N_3031,N_2572,N_2717);
nand U3032 (N_3032,N_2537,N_2625);
xor U3033 (N_3033,N_2523,N_2761);
nor U3034 (N_3034,N_2794,N_2737);
or U3035 (N_3035,N_2729,N_2991);
nand U3036 (N_3036,N_2935,N_2664);
or U3037 (N_3037,N_2993,N_2639);
nand U3038 (N_3038,N_2505,N_2513);
nand U3039 (N_3039,N_2889,N_2973);
nor U3040 (N_3040,N_2878,N_2521);
nand U3041 (N_3041,N_2775,N_2979);
nand U3042 (N_3042,N_2702,N_2617);
xor U3043 (N_3043,N_2825,N_2706);
nor U3044 (N_3044,N_2733,N_2573);
nor U3045 (N_3045,N_2703,N_2917);
xor U3046 (N_3046,N_2589,N_2791);
or U3047 (N_3047,N_2862,N_2575);
and U3048 (N_3048,N_2546,N_2928);
and U3049 (N_3049,N_2827,N_2568);
and U3050 (N_3050,N_2656,N_2666);
nor U3051 (N_3051,N_2719,N_2882);
and U3052 (N_3052,N_2716,N_2588);
nor U3053 (N_3053,N_2540,N_2632);
or U3054 (N_3054,N_2912,N_2800);
nor U3055 (N_3055,N_2820,N_2661);
or U3056 (N_3056,N_2541,N_2796);
xor U3057 (N_3057,N_2644,N_2929);
or U3058 (N_3058,N_2808,N_2557);
nor U3059 (N_3059,N_2839,N_2699);
xnor U3060 (N_3060,N_2501,N_2643);
xor U3061 (N_3061,N_2832,N_2772);
nor U3062 (N_3062,N_2780,N_2823);
nand U3063 (N_3063,N_2778,N_2872);
nor U3064 (N_3064,N_2844,N_2956);
or U3065 (N_3065,N_2939,N_2885);
nor U3066 (N_3066,N_2641,N_2861);
and U3067 (N_3067,N_2893,N_2654);
or U3068 (N_3068,N_2743,N_2810);
nor U3069 (N_3069,N_2500,N_2970);
nand U3070 (N_3070,N_2927,N_2777);
nor U3071 (N_3071,N_2842,N_2910);
xnor U3072 (N_3072,N_2936,N_2946);
and U3073 (N_3073,N_2809,N_2564);
or U3074 (N_3074,N_2819,N_2765);
xnor U3075 (N_3075,N_2605,N_2818);
and U3076 (N_3076,N_2548,N_2616);
nor U3077 (N_3077,N_2709,N_2652);
xor U3078 (N_3078,N_2902,N_2516);
nand U3079 (N_3079,N_2914,N_2595);
or U3080 (N_3080,N_2678,N_2840);
or U3081 (N_3081,N_2742,N_2785);
and U3082 (N_3082,N_2507,N_2817);
xor U3083 (N_3083,N_2843,N_2553);
xnor U3084 (N_3084,N_2567,N_2525);
xor U3085 (N_3085,N_2806,N_2745);
xnor U3086 (N_3086,N_2887,N_2905);
or U3087 (N_3087,N_2650,N_2807);
nand U3088 (N_3088,N_2680,N_2795);
or U3089 (N_3089,N_2579,N_2682);
nor U3090 (N_3090,N_2648,N_2837);
xnor U3091 (N_3091,N_2799,N_2606);
nand U3092 (N_3092,N_2754,N_2526);
nor U3093 (N_3093,N_2614,N_2998);
xnor U3094 (N_3094,N_2628,N_2934);
xor U3095 (N_3095,N_2955,N_2597);
or U3096 (N_3096,N_2985,N_2708);
xor U3097 (N_3097,N_2972,N_2763);
or U3098 (N_3098,N_2707,N_2877);
xnor U3099 (N_3099,N_2860,N_2975);
and U3100 (N_3100,N_2555,N_2725);
or U3101 (N_3101,N_2978,N_2988);
nor U3102 (N_3102,N_2890,N_2602);
or U3103 (N_3103,N_2875,N_2762);
and U3104 (N_3104,N_2610,N_2950);
and U3105 (N_3105,N_2609,N_2740);
and U3106 (N_3106,N_2874,N_2947);
xor U3107 (N_3107,N_2536,N_2888);
nand U3108 (N_3108,N_2969,N_2668);
nor U3109 (N_3109,N_2915,N_2550);
and U3110 (N_3110,N_2994,N_2879);
xnor U3111 (N_3111,N_2816,N_2594);
xor U3112 (N_3112,N_2622,N_2880);
nand U3113 (N_3113,N_2590,N_2951);
or U3114 (N_3114,N_2720,N_2629);
and U3115 (N_3115,N_2750,N_2549);
nor U3116 (N_3116,N_2620,N_2534);
or U3117 (N_3117,N_2721,N_2527);
nor U3118 (N_3118,N_2736,N_2562);
and U3119 (N_3119,N_2522,N_2925);
xnor U3120 (N_3120,N_2989,N_2876);
nor U3121 (N_3121,N_2665,N_2962);
or U3122 (N_3122,N_2831,N_2611);
xor U3123 (N_3123,N_2630,N_2854);
nand U3124 (N_3124,N_2683,N_2604);
nand U3125 (N_3125,N_2857,N_2959);
xor U3126 (N_3126,N_2583,N_2667);
xnor U3127 (N_3127,N_2677,N_2675);
nand U3128 (N_3128,N_2834,N_2633);
nand U3129 (N_3129,N_2982,N_2533);
or U3130 (N_3130,N_2734,N_2958);
nand U3131 (N_3131,N_2612,N_2577);
xnor U3132 (N_3132,N_2853,N_2730);
or U3133 (N_3133,N_2714,N_2937);
nor U3134 (N_3134,N_2971,N_2711);
nand U3135 (N_3135,N_2545,N_2582);
nand U3136 (N_3136,N_2797,N_2770);
and U3137 (N_3137,N_2891,N_2952);
nand U3138 (N_3138,N_2695,N_2759);
nor U3139 (N_3139,N_2760,N_2578);
xnor U3140 (N_3140,N_2715,N_2941);
and U3141 (N_3141,N_2576,N_2676);
nor U3142 (N_3142,N_2580,N_2869);
nand U3143 (N_3143,N_2566,N_2517);
xor U3144 (N_3144,N_2528,N_2694);
nand U3145 (N_3145,N_2957,N_2506);
and U3146 (N_3146,N_2909,N_2789);
xnor U3147 (N_3147,N_2944,N_2776);
and U3148 (N_3148,N_2690,N_2768);
nand U3149 (N_3149,N_2859,N_2940);
xnor U3150 (N_3150,N_2987,N_2731);
xnor U3151 (N_3151,N_2518,N_2697);
nor U3152 (N_3152,N_2892,N_2601);
nor U3153 (N_3153,N_2773,N_2623);
and U3154 (N_3154,N_2977,N_2774);
xnor U3155 (N_3155,N_2524,N_2873);
nand U3156 (N_3156,N_2906,N_2689);
nand U3157 (N_3157,N_2613,N_2901);
xor U3158 (N_3158,N_2790,N_2757);
nor U3159 (N_3159,N_2556,N_2646);
nor U3160 (N_3160,N_2949,N_2726);
or U3161 (N_3161,N_2559,N_2681);
nor U3162 (N_3162,N_2896,N_2836);
xor U3163 (N_3163,N_2514,N_2698);
nor U3164 (N_3164,N_2916,N_2674);
and U3165 (N_3165,N_2986,N_2748);
or U3166 (N_3166,N_2598,N_2771);
nand U3167 (N_3167,N_2552,N_2569);
xor U3168 (N_3168,N_2728,N_2551);
xnor U3169 (N_3169,N_2532,N_2945);
or U3170 (N_3170,N_2504,N_2826);
or U3171 (N_3171,N_2531,N_2701);
and U3172 (N_3172,N_2747,N_2783);
nor U3173 (N_3173,N_2647,N_2997);
nor U3174 (N_3174,N_2960,N_2913);
and U3175 (N_3175,N_2883,N_2930);
xnor U3176 (N_3176,N_2866,N_2636);
and U3177 (N_3177,N_2990,N_2627);
and U3178 (N_3178,N_2884,N_2995);
or U3179 (N_3179,N_2642,N_2700);
or U3180 (N_3180,N_2838,N_2502);
nor U3181 (N_3181,N_2626,N_2741);
xnor U3182 (N_3182,N_2835,N_2932);
xnor U3183 (N_3183,N_2984,N_2755);
nand U3184 (N_3184,N_2822,N_2980);
and U3185 (N_3185,N_2724,N_2804);
nand U3186 (N_3186,N_2919,N_2871);
or U3187 (N_3187,N_2963,N_2581);
xnor U3188 (N_3188,N_2718,N_2558);
and U3189 (N_3189,N_2704,N_2593);
or U3190 (N_3190,N_2600,N_2895);
nand U3191 (N_3191,N_2670,N_2705);
and U3192 (N_3192,N_2865,N_2744);
nor U3193 (N_3193,N_2954,N_2786);
and U3194 (N_3194,N_2660,N_2563);
nand U3195 (N_3195,N_2864,N_2603);
or U3196 (N_3196,N_2992,N_2624);
and U3197 (N_3197,N_2586,N_2821);
or U3198 (N_3198,N_2672,N_2964);
xor U3199 (N_3199,N_2519,N_2710);
nor U3200 (N_3200,N_2897,N_2723);
nand U3201 (N_3201,N_2784,N_2686);
and U3202 (N_3202,N_2863,N_2850);
or U3203 (N_3203,N_2815,N_2651);
nor U3204 (N_3204,N_2544,N_2659);
xnor U3205 (N_3205,N_2554,N_2539);
or U3206 (N_3206,N_2965,N_2848);
xor U3207 (N_3207,N_2828,N_2658);
xnor U3208 (N_3208,N_2855,N_2673);
and U3209 (N_3209,N_2587,N_2509);
nand U3210 (N_3210,N_2981,N_2637);
nand U3211 (N_3211,N_2983,N_2868);
and U3212 (N_3212,N_2574,N_2781);
or U3213 (N_3213,N_2565,N_2846);
and U3214 (N_3214,N_2684,N_2758);
nor U3215 (N_3215,N_2530,N_2713);
nor U3216 (N_3216,N_2856,N_2592);
xnor U3217 (N_3217,N_2503,N_2515);
nand U3218 (N_3218,N_2584,N_2921);
nor U3219 (N_3219,N_2812,N_2908);
or U3220 (N_3220,N_2899,N_2508);
xor U3221 (N_3221,N_2619,N_2510);
or U3222 (N_3222,N_2631,N_2788);
nor U3223 (N_3223,N_2561,N_2953);
or U3224 (N_3224,N_2645,N_2798);
nor U3225 (N_3225,N_2640,N_2943);
or U3226 (N_3226,N_2900,N_2542);
xnor U3227 (N_3227,N_2811,N_2591);
nor U3228 (N_3228,N_2767,N_2920);
or U3229 (N_3229,N_2732,N_2722);
nor U3230 (N_3230,N_2543,N_2961);
xor U3231 (N_3231,N_2769,N_2829);
and U3232 (N_3232,N_2752,N_2692);
xor U3233 (N_3233,N_2512,N_2870);
nand U3234 (N_3234,N_2607,N_2830);
xor U3235 (N_3235,N_2662,N_2735);
xor U3236 (N_3236,N_2538,N_2881);
xnor U3237 (N_3237,N_2851,N_2585);
xor U3238 (N_3238,N_2907,N_2751);
nor U3239 (N_3239,N_2849,N_2813);
xor U3240 (N_3240,N_2814,N_2922);
nor U3241 (N_3241,N_2727,N_2894);
or U3242 (N_3242,N_2867,N_2933);
nor U3243 (N_3243,N_2511,N_2687);
nand U3244 (N_3244,N_2520,N_2608);
or U3245 (N_3245,N_2898,N_2924);
or U3246 (N_3246,N_2938,N_2547);
xnor U3247 (N_3247,N_2824,N_2967);
or U3248 (N_3248,N_2805,N_2852);
or U3249 (N_3249,N_2739,N_2679);
and U3250 (N_3250,N_2523,N_2674);
or U3251 (N_3251,N_2959,N_2604);
or U3252 (N_3252,N_2802,N_2894);
xnor U3253 (N_3253,N_2559,N_2656);
or U3254 (N_3254,N_2587,N_2802);
and U3255 (N_3255,N_2547,N_2731);
and U3256 (N_3256,N_2675,N_2993);
nand U3257 (N_3257,N_2724,N_2550);
or U3258 (N_3258,N_2779,N_2815);
xor U3259 (N_3259,N_2735,N_2612);
nor U3260 (N_3260,N_2760,N_2985);
and U3261 (N_3261,N_2569,N_2718);
nand U3262 (N_3262,N_2577,N_2932);
nand U3263 (N_3263,N_2822,N_2960);
or U3264 (N_3264,N_2834,N_2738);
nand U3265 (N_3265,N_2673,N_2634);
or U3266 (N_3266,N_2816,N_2744);
nor U3267 (N_3267,N_2630,N_2901);
xnor U3268 (N_3268,N_2674,N_2749);
xor U3269 (N_3269,N_2793,N_2789);
nand U3270 (N_3270,N_2634,N_2960);
and U3271 (N_3271,N_2570,N_2538);
xnor U3272 (N_3272,N_2763,N_2518);
xor U3273 (N_3273,N_2816,N_2693);
xnor U3274 (N_3274,N_2783,N_2728);
or U3275 (N_3275,N_2983,N_2703);
or U3276 (N_3276,N_2993,N_2876);
nor U3277 (N_3277,N_2979,N_2702);
and U3278 (N_3278,N_2965,N_2869);
xnor U3279 (N_3279,N_2996,N_2725);
and U3280 (N_3280,N_2597,N_2823);
nor U3281 (N_3281,N_2505,N_2760);
and U3282 (N_3282,N_2969,N_2564);
and U3283 (N_3283,N_2937,N_2729);
xor U3284 (N_3284,N_2532,N_2794);
xnor U3285 (N_3285,N_2711,N_2905);
xor U3286 (N_3286,N_2832,N_2766);
nand U3287 (N_3287,N_2575,N_2699);
xor U3288 (N_3288,N_2560,N_2831);
nand U3289 (N_3289,N_2643,N_2831);
nor U3290 (N_3290,N_2828,N_2832);
nand U3291 (N_3291,N_2720,N_2813);
xnor U3292 (N_3292,N_2707,N_2902);
nand U3293 (N_3293,N_2925,N_2821);
nor U3294 (N_3294,N_2530,N_2769);
nor U3295 (N_3295,N_2505,N_2619);
xor U3296 (N_3296,N_2754,N_2998);
and U3297 (N_3297,N_2692,N_2823);
or U3298 (N_3298,N_2992,N_2844);
or U3299 (N_3299,N_2792,N_2939);
nand U3300 (N_3300,N_2615,N_2595);
nand U3301 (N_3301,N_2745,N_2533);
nor U3302 (N_3302,N_2540,N_2690);
xor U3303 (N_3303,N_2540,N_2967);
and U3304 (N_3304,N_2548,N_2669);
nand U3305 (N_3305,N_2541,N_2550);
nor U3306 (N_3306,N_2998,N_2857);
or U3307 (N_3307,N_2962,N_2976);
xnor U3308 (N_3308,N_2601,N_2823);
nor U3309 (N_3309,N_2857,N_2593);
nor U3310 (N_3310,N_2984,N_2957);
nor U3311 (N_3311,N_2661,N_2925);
or U3312 (N_3312,N_2817,N_2676);
and U3313 (N_3313,N_2656,N_2794);
xnor U3314 (N_3314,N_2914,N_2651);
xnor U3315 (N_3315,N_2510,N_2940);
and U3316 (N_3316,N_2867,N_2548);
nand U3317 (N_3317,N_2736,N_2668);
nor U3318 (N_3318,N_2856,N_2766);
or U3319 (N_3319,N_2516,N_2644);
or U3320 (N_3320,N_2682,N_2822);
or U3321 (N_3321,N_2558,N_2578);
xnor U3322 (N_3322,N_2970,N_2788);
or U3323 (N_3323,N_2663,N_2944);
nand U3324 (N_3324,N_2554,N_2934);
nand U3325 (N_3325,N_2704,N_2818);
nand U3326 (N_3326,N_2751,N_2703);
nand U3327 (N_3327,N_2596,N_2986);
or U3328 (N_3328,N_2670,N_2543);
xnor U3329 (N_3329,N_2710,N_2520);
and U3330 (N_3330,N_2773,N_2736);
or U3331 (N_3331,N_2620,N_2548);
and U3332 (N_3332,N_2562,N_2907);
or U3333 (N_3333,N_2842,N_2602);
xnor U3334 (N_3334,N_2913,N_2596);
nor U3335 (N_3335,N_2840,N_2681);
nand U3336 (N_3336,N_2738,N_2814);
and U3337 (N_3337,N_2891,N_2608);
nor U3338 (N_3338,N_2540,N_2754);
nor U3339 (N_3339,N_2971,N_2554);
and U3340 (N_3340,N_2691,N_2962);
xor U3341 (N_3341,N_2814,N_2804);
nand U3342 (N_3342,N_2545,N_2874);
and U3343 (N_3343,N_2531,N_2698);
nand U3344 (N_3344,N_2957,N_2661);
and U3345 (N_3345,N_2541,N_2816);
nand U3346 (N_3346,N_2881,N_2895);
and U3347 (N_3347,N_2504,N_2536);
nor U3348 (N_3348,N_2756,N_2705);
xor U3349 (N_3349,N_2705,N_2523);
nor U3350 (N_3350,N_2613,N_2668);
or U3351 (N_3351,N_2658,N_2986);
or U3352 (N_3352,N_2892,N_2850);
or U3353 (N_3353,N_2659,N_2976);
nor U3354 (N_3354,N_2628,N_2747);
nand U3355 (N_3355,N_2897,N_2814);
xor U3356 (N_3356,N_2924,N_2862);
nor U3357 (N_3357,N_2570,N_2886);
xnor U3358 (N_3358,N_2908,N_2918);
xnor U3359 (N_3359,N_2889,N_2725);
and U3360 (N_3360,N_2647,N_2707);
xnor U3361 (N_3361,N_2993,N_2572);
and U3362 (N_3362,N_2941,N_2518);
or U3363 (N_3363,N_2963,N_2518);
xnor U3364 (N_3364,N_2741,N_2984);
and U3365 (N_3365,N_2926,N_2799);
xor U3366 (N_3366,N_2680,N_2744);
xnor U3367 (N_3367,N_2878,N_2874);
and U3368 (N_3368,N_2610,N_2508);
or U3369 (N_3369,N_2892,N_2657);
or U3370 (N_3370,N_2966,N_2569);
nor U3371 (N_3371,N_2548,N_2911);
xnor U3372 (N_3372,N_2726,N_2871);
nor U3373 (N_3373,N_2793,N_2638);
or U3374 (N_3374,N_2676,N_2895);
nand U3375 (N_3375,N_2539,N_2836);
xor U3376 (N_3376,N_2627,N_2706);
or U3377 (N_3377,N_2929,N_2526);
nand U3378 (N_3378,N_2680,N_2979);
or U3379 (N_3379,N_2819,N_2815);
xnor U3380 (N_3380,N_2696,N_2663);
nor U3381 (N_3381,N_2508,N_2557);
xor U3382 (N_3382,N_2902,N_2942);
nand U3383 (N_3383,N_2850,N_2925);
nor U3384 (N_3384,N_2883,N_2814);
nand U3385 (N_3385,N_2527,N_2612);
and U3386 (N_3386,N_2947,N_2571);
and U3387 (N_3387,N_2952,N_2633);
nand U3388 (N_3388,N_2677,N_2779);
xnor U3389 (N_3389,N_2624,N_2953);
nor U3390 (N_3390,N_2523,N_2738);
nor U3391 (N_3391,N_2683,N_2975);
and U3392 (N_3392,N_2969,N_2927);
and U3393 (N_3393,N_2721,N_2601);
nor U3394 (N_3394,N_2724,N_2813);
xor U3395 (N_3395,N_2981,N_2852);
or U3396 (N_3396,N_2965,N_2805);
or U3397 (N_3397,N_2955,N_2807);
or U3398 (N_3398,N_2948,N_2837);
or U3399 (N_3399,N_2693,N_2640);
or U3400 (N_3400,N_2633,N_2850);
xor U3401 (N_3401,N_2981,N_2873);
nor U3402 (N_3402,N_2706,N_2978);
or U3403 (N_3403,N_2632,N_2914);
or U3404 (N_3404,N_2777,N_2653);
or U3405 (N_3405,N_2899,N_2502);
and U3406 (N_3406,N_2511,N_2779);
or U3407 (N_3407,N_2812,N_2926);
nand U3408 (N_3408,N_2765,N_2577);
and U3409 (N_3409,N_2946,N_2567);
nor U3410 (N_3410,N_2570,N_2802);
or U3411 (N_3411,N_2994,N_2660);
and U3412 (N_3412,N_2934,N_2809);
and U3413 (N_3413,N_2562,N_2580);
nor U3414 (N_3414,N_2690,N_2947);
xor U3415 (N_3415,N_2891,N_2814);
and U3416 (N_3416,N_2947,N_2663);
and U3417 (N_3417,N_2899,N_2532);
xnor U3418 (N_3418,N_2866,N_2846);
xor U3419 (N_3419,N_2612,N_2530);
or U3420 (N_3420,N_2603,N_2767);
or U3421 (N_3421,N_2823,N_2934);
and U3422 (N_3422,N_2719,N_2607);
nand U3423 (N_3423,N_2713,N_2594);
nor U3424 (N_3424,N_2844,N_2812);
nor U3425 (N_3425,N_2625,N_2781);
or U3426 (N_3426,N_2508,N_2663);
and U3427 (N_3427,N_2668,N_2531);
nand U3428 (N_3428,N_2733,N_2542);
and U3429 (N_3429,N_2640,N_2592);
xnor U3430 (N_3430,N_2738,N_2969);
or U3431 (N_3431,N_2871,N_2929);
and U3432 (N_3432,N_2729,N_2530);
nor U3433 (N_3433,N_2653,N_2895);
or U3434 (N_3434,N_2517,N_2547);
nor U3435 (N_3435,N_2675,N_2663);
nand U3436 (N_3436,N_2515,N_2706);
and U3437 (N_3437,N_2768,N_2745);
or U3438 (N_3438,N_2903,N_2769);
and U3439 (N_3439,N_2662,N_2978);
nor U3440 (N_3440,N_2774,N_2904);
and U3441 (N_3441,N_2514,N_2595);
nand U3442 (N_3442,N_2992,N_2982);
nor U3443 (N_3443,N_2741,N_2551);
or U3444 (N_3444,N_2915,N_2921);
nand U3445 (N_3445,N_2895,N_2661);
nand U3446 (N_3446,N_2845,N_2835);
nor U3447 (N_3447,N_2859,N_2752);
and U3448 (N_3448,N_2538,N_2847);
or U3449 (N_3449,N_2630,N_2839);
and U3450 (N_3450,N_2660,N_2583);
nand U3451 (N_3451,N_2962,N_2600);
and U3452 (N_3452,N_2927,N_2984);
or U3453 (N_3453,N_2565,N_2945);
nor U3454 (N_3454,N_2920,N_2745);
and U3455 (N_3455,N_2662,N_2508);
xor U3456 (N_3456,N_2874,N_2865);
or U3457 (N_3457,N_2721,N_2963);
or U3458 (N_3458,N_2868,N_2582);
and U3459 (N_3459,N_2994,N_2792);
and U3460 (N_3460,N_2941,N_2806);
nand U3461 (N_3461,N_2616,N_2907);
xnor U3462 (N_3462,N_2919,N_2743);
nand U3463 (N_3463,N_2988,N_2942);
or U3464 (N_3464,N_2901,N_2745);
and U3465 (N_3465,N_2547,N_2647);
and U3466 (N_3466,N_2869,N_2964);
xor U3467 (N_3467,N_2951,N_2985);
xor U3468 (N_3468,N_2595,N_2998);
xor U3469 (N_3469,N_2841,N_2575);
and U3470 (N_3470,N_2767,N_2540);
nor U3471 (N_3471,N_2953,N_2545);
or U3472 (N_3472,N_2727,N_2696);
nor U3473 (N_3473,N_2628,N_2667);
or U3474 (N_3474,N_2921,N_2952);
or U3475 (N_3475,N_2577,N_2637);
nor U3476 (N_3476,N_2683,N_2994);
nand U3477 (N_3477,N_2994,N_2912);
and U3478 (N_3478,N_2520,N_2862);
xnor U3479 (N_3479,N_2683,N_2743);
and U3480 (N_3480,N_2709,N_2925);
nor U3481 (N_3481,N_2913,N_2565);
nand U3482 (N_3482,N_2546,N_2711);
nand U3483 (N_3483,N_2582,N_2899);
nand U3484 (N_3484,N_2632,N_2596);
or U3485 (N_3485,N_2825,N_2975);
xor U3486 (N_3486,N_2835,N_2588);
nor U3487 (N_3487,N_2858,N_2552);
and U3488 (N_3488,N_2730,N_2776);
nand U3489 (N_3489,N_2758,N_2932);
and U3490 (N_3490,N_2978,N_2860);
xnor U3491 (N_3491,N_2778,N_2545);
nor U3492 (N_3492,N_2895,N_2725);
and U3493 (N_3493,N_2897,N_2600);
xor U3494 (N_3494,N_2956,N_2630);
nand U3495 (N_3495,N_2813,N_2743);
nand U3496 (N_3496,N_2635,N_2888);
nand U3497 (N_3497,N_2536,N_2592);
nand U3498 (N_3498,N_2991,N_2530);
xnor U3499 (N_3499,N_2838,N_2672);
nand U3500 (N_3500,N_3386,N_3020);
nand U3501 (N_3501,N_3091,N_3115);
nand U3502 (N_3502,N_3157,N_3273);
and U3503 (N_3503,N_3352,N_3397);
nor U3504 (N_3504,N_3121,N_3443);
and U3505 (N_3505,N_3034,N_3106);
nand U3506 (N_3506,N_3040,N_3127);
or U3507 (N_3507,N_3399,N_3084);
xor U3508 (N_3508,N_3264,N_3388);
and U3509 (N_3509,N_3039,N_3174);
or U3510 (N_3510,N_3315,N_3165);
nor U3511 (N_3511,N_3151,N_3013);
or U3512 (N_3512,N_3043,N_3134);
xnor U3513 (N_3513,N_3160,N_3304);
nor U3514 (N_3514,N_3063,N_3338);
nand U3515 (N_3515,N_3221,N_3009);
xor U3516 (N_3516,N_3495,N_3163);
xnor U3517 (N_3517,N_3267,N_3000);
nand U3518 (N_3518,N_3290,N_3204);
nand U3519 (N_3519,N_3045,N_3396);
or U3520 (N_3520,N_3008,N_3177);
nor U3521 (N_3521,N_3414,N_3027);
nor U3522 (N_3522,N_3311,N_3012);
or U3523 (N_3523,N_3108,N_3317);
nand U3524 (N_3524,N_3448,N_3498);
and U3525 (N_3525,N_3103,N_3131);
xnor U3526 (N_3526,N_3047,N_3014);
nor U3527 (N_3527,N_3413,N_3240);
xor U3528 (N_3528,N_3085,N_3024);
or U3529 (N_3529,N_3345,N_3324);
or U3530 (N_3530,N_3441,N_3263);
and U3531 (N_3531,N_3143,N_3124);
and U3532 (N_3532,N_3220,N_3036);
or U3533 (N_3533,N_3493,N_3011);
nor U3534 (N_3534,N_3403,N_3444);
nor U3535 (N_3535,N_3382,N_3342);
nand U3536 (N_3536,N_3050,N_3455);
nor U3537 (N_3537,N_3445,N_3195);
and U3538 (N_3538,N_3051,N_3225);
xnor U3539 (N_3539,N_3364,N_3281);
nand U3540 (N_3540,N_3019,N_3420);
nor U3541 (N_3541,N_3351,N_3052);
and U3542 (N_3542,N_3276,N_3496);
nand U3543 (N_3543,N_3083,N_3330);
nand U3544 (N_3544,N_3437,N_3175);
or U3545 (N_3545,N_3298,N_3410);
xor U3546 (N_3546,N_3480,N_3499);
and U3547 (N_3547,N_3142,N_3172);
and U3548 (N_3548,N_3046,N_3042);
or U3549 (N_3549,N_3132,N_3468);
xnor U3550 (N_3550,N_3446,N_3004);
and U3551 (N_3551,N_3377,N_3023);
nand U3552 (N_3552,N_3442,N_3246);
xor U3553 (N_3553,N_3475,N_3400);
and U3554 (N_3554,N_3375,N_3378);
nor U3555 (N_3555,N_3275,N_3032);
nand U3556 (N_3556,N_3236,N_3238);
or U3557 (N_3557,N_3439,N_3357);
and U3558 (N_3558,N_3299,N_3206);
or U3559 (N_3559,N_3099,N_3379);
nor U3560 (N_3560,N_3073,N_3322);
xor U3561 (N_3561,N_3173,N_3458);
xnor U3562 (N_3562,N_3485,N_3309);
nor U3563 (N_3563,N_3079,N_3104);
xor U3564 (N_3564,N_3018,N_3430);
and U3565 (N_3565,N_3144,N_3270);
and U3566 (N_3566,N_3207,N_3295);
and U3567 (N_3567,N_3257,N_3249);
nor U3568 (N_3568,N_3006,N_3334);
and U3569 (N_3569,N_3097,N_3340);
nor U3570 (N_3570,N_3055,N_3321);
nor U3571 (N_3571,N_3093,N_3323);
nand U3572 (N_3572,N_3128,N_3069);
xor U3573 (N_3573,N_3201,N_3152);
and U3574 (N_3574,N_3194,N_3021);
or U3575 (N_3575,N_3117,N_3002);
nor U3576 (N_3576,N_3030,N_3261);
or U3577 (N_3577,N_3426,N_3456);
and U3578 (N_3578,N_3348,N_3251);
and U3579 (N_3579,N_3433,N_3466);
nor U3580 (N_3580,N_3478,N_3297);
and U3581 (N_3581,N_3428,N_3164);
and U3582 (N_3582,N_3429,N_3041);
xnor U3583 (N_3583,N_3343,N_3349);
or U3584 (N_3584,N_3112,N_3028);
xnor U3585 (N_3585,N_3044,N_3235);
or U3586 (N_3586,N_3368,N_3453);
or U3587 (N_3587,N_3440,N_3260);
or U3588 (N_3588,N_3048,N_3398);
and U3589 (N_3589,N_3471,N_3469);
xnor U3590 (N_3590,N_3365,N_3185);
nor U3591 (N_3591,N_3037,N_3149);
nor U3592 (N_3592,N_3353,N_3059);
nor U3593 (N_3593,N_3347,N_3331);
nand U3594 (N_3594,N_3064,N_3186);
nor U3595 (N_3595,N_3158,N_3150);
and U3596 (N_3596,N_3291,N_3215);
or U3597 (N_3597,N_3286,N_3213);
and U3598 (N_3598,N_3184,N_3129);
nand U3599 (N_3599,N_3393,N_3003);
xnor U3600 (N_3600,N_3136,N_3071);
and U3601 (N_3601,N_3082,N_3133);
xor U3602 (N_3602,N_3060,N_3373);
or U3603 (N_3603,N_3459,N_3216);
nand U3604 (N_3604,N_3384,N_3326);
nor U3605 (N_3605,N_3171,N_3359);
nand U3606 (N_3606,N_3226,N_3248);
nor U3607 (N_3607,N_3422,N_3355);
nand U3608 (N_3608,N_3395,N_3411);
and U3609 (N_3609,N_3409,N_3125);
xnor U3610 (N_3610,N_3107,N_3109);
xnor U3611 (N_3611,N_3056,N_3483);
or U3612 (N_3612,N_3457,N_3095);
xor U3613 (N_3613,N_3391,N_3031);
xor U3614 (N_3614,N_3102,N_3074);
nand U3615 (N_3615,N_3360,N_3168);
nand U3616 (N_3616,N_3310,N_3068);
or U3617 (N_3617,N_3203,N_3219);
nor U3618 (N_3618,N_3147,N_3176);
or U3619 (N_3619,N_3313,N_3341);
or U3620 (N_3620,N_3146,N_3241);
xor U3621 (N_3621,N_3209,N_3022);
and U3622 (N_3622,N_3244,N_3462);
xor U3623 (N_3623,N_3421,N_3490);
or U3624 (N_3624,N_3318,N_3332);
or U3625 (N_3625,N_3271,N_3202);
or U3626 (N_3626,N_3161,N_3029);
and U3627 (N_3627,N_3312,N_3416);
or U3628 (N_3628,N_3007,N_3372);
and U3629 (N_3629,N_3081,N_3450);
nand U3630 (N_3630,N_3156,N_3086);
nand U3631 (N_3631,N_3141,N_3371);
or U3632 (N_3632,N_3301,N_3350);
and U3633 (N_3633,N_3245,N_3138);
xor U3634 (N_3634,N_3366,N_3182);
or U3635 (N_3635,N_3401,N_3300);
or U3636 (N_3636,N_3474,N_3277);
xnor U3637 (N_3637,N_3449,N_3385);
or U3638 (N_3638,N_3199,N_3228);
nand U3639 (N_3639,N_3424,N_3288);
nor U3640 (N_3640,N_3354,N_3337);
xnor U3641 (N_3641,N_3053,N_3427);
nor U3642 (N_3642,N_3162,N_3239);
nand U3643 (N_3643,N_3061,N_3287);
and U3644 (N_3644,N_3408,N_3285);
xnor U3645 (N_3645,N_3392,N_3335);
and U3646 (N_3646,N_3434,N_3234);
xor U3647 (N_3647,N_3314,N_3284);
or U3648 (N_3648,N_3394,N_3080);
nor U3649 (N_3649,N_3049,N_3178);
nand U3650 (N_3650,N_3319,N_3497);
nor U3651 (N_3651,N_3405,N_3463);
xor U3652 (N_3652,N_3296,N_3118);
and U3653 (N_3653,N_3283,N_3200);
and U3654 (N_3654,N_3247,N_3122);
nor U3655 (N_3655,N_3001,N_3035);
or U3656 (N_3656,N_3193,N_3017);
and U3657 (N_3657,N_3197,N_3180);
nand U3658 (N_3658,N_3016,N_3460);
and U3659 (N_3659,N_3269,N_3482);
nand U3660 (N_3660,N_3033,N_3077);
or U3661 (N_3661,N_3205,N_3419);
and U3662 (N_3662,N_3302,N_3417);
or U3663 (N_3663,N_3087,N_3452);
nor U3664 (N_3664,N_3328,N_3005);
xnor U3665 (N_3665,N_3113,N_3116);
nor U3666 (N_3666,N_3015,N_3362);
or U3667 (N_3667,N_3230,N_3383);
and U3668 (N_3668,N_3252,N_3096);
or U3669 (N_3669,N_3438,N_3232);
and U3670 (N_3670,N_3038,N_3320);
xnor U3671 (N_3671,N_3293,N_3489);
xor U3672 (N_3672,N_3306,N_3370);
nor U3673 (N_3673,N_3189,N_3242);
nand U3674 (N_3674,N_3488,N_3307);
nand U3675 (N_3675,N_3222,N_3363);
xnor U3676 (N_3676,N_3358,N_3167);
and U3677 (N_3677,N_3303,N_3123);
or U3678 (N_3678,N_3447,N_3211);
and U3679 (N_3679,N_3436,N_3327);
or U3680 (N_3680,N_3254,N_3208);
xor U3681 (N_3681,N_3090,N_3407);
or U3682 (N_3682,N_3120,N_3272);
nand U3683 (N_3683,N_3105,N_3231);
xor U3684 (N_3684,N_3058,N_3253);
or U3685 (N_3685,N_3406,N_3089);
nand U3686 (N_3686,N_3196,N_3210);
nand U3687 (N_3687,N_3119,N_3153);
nor U3688 (N_3688,N_3227,N_3088);
and U3689 (N_3689,N_3470,N_3479);
and U3690 (N_3690,N_3250,N_3237);
xor U3691 (N_3691,N_3380,N_3130);
or U3692 (N_3692,N_3333,N_3265);
and U3693 (N_3693,N_3187,N_3212);
nor U3694 (N_3694,N_3078,N_3170);
or U3695 (N_3695,N_3188,N_3473);
xor U3696 (N_3696,N_3191,N_3140);
nand U3697 (N_3697,N_3491,N_3435);
or U3698 (N_3698,N_3404,N_3477);
xnor U3699 (N_3699,N_3329,N_3390);
nor U3700 (N_3700,N_3361,N_3316);
nor U3701 (N_3701,N_3486,N_3070);
nand U3702 (N_3702,N_3094,N_3101);
nand U3703 (N_3703,N_3278,N_3339);
nor U3704 (N_3704,N_3381,N_3075);
xnor U3705 (N_3705,N_3465,N_3256);
or U3706 (N_3706,N_3100,N_3266);
or U3707 (N_3707,N_3279,N_3259);
nor U3708 (N_3708,N_3192,N_3305);
xor U3709 (N_3709,N_3282,N_3217);
nor U3710 (N_3710,N_3092,N_3110);
or U3711 (N_3711,N_3476,N_3255);
or U3712 (N_3712,N_3423,N_3218);
nor U3713 (N_3713,N_3415,N_3389);
xor U3714 (N_3714,N_3487,N_3214);
xor U3715 (N_3715,N_3198,N_3154);
xor U3716 (N_3716,N_3135,N_3467);
nor U3717 (N_3717,N_3454,N_3472);
or U3718 (N_3718,N_3268,N_3484);
or U3719 (N_3719,N_3292,N_3367);
and U3720 (N_3720,N_3374,N_3233);
xnor U3721 (N_3721,N_3148,N_3065);
nand U3722 (N_3722,N_3464,N_3344);
and U3723 (N_3723,N_3169,N_3114);
and U3724 (N_3724,N_3224,N_3258);
nor U3725 (N_3725,N_3274,N_3183);
nand U3726 (N_3726,N_3067,N_3076);
xnor U3727 (N_3727,N_3126,N_3387);
or U3728 (N_3728,N_3159,N_3376);
xnor U3729 (N_3729,N_3026,N_3179);
xnor U3730 (N_3730,N_3451,N_3098);
nand U3731 (N_3731,N_3425,N_3432);
and U3732 (N_3732,N_3431,N_3072);
nor U3733 (N_3733,N_3294,N_3418);
nor U3734 (N_3734,N_3229,N_3280);
nor U3735 (N_3735,N_3137,N_3166);
nor U3736 (N_3736,N_3062,N_3402);
nor U3737 (N_3737,N_3369,N_3262);
xnor U3738 (N_3738,N_3190,N_3181);
or U3739 (N_3739,N_3155,N_3139);
and U3740 (N_3740,N_3308,N_3346);
nor U3741 (N_3741,N_3025,N_3461);
nand U3742 (N_3742,N_3356,N_3289);
and U3743 (N_3743,N_3336,N_3243);
and U3744 (N_3744,N_3325,N_3492);
nor U3745 (N_3745,N_3066,N_3054);
and U3746 (N_3746,N_3494,N_3412);
xor U3747 (N_3747,N_3223,N_3057);
nand U3748 (N_3748,N_3481,N_3145);
or U3749 (N_3749,N_3111,N_3010);
or U3750 (N_3750,N_3185,N_3122);
nor U3751 (N_3751,N_3436,N_3051);
nor U3752 (N_3752,N_3009,N_3373);
nand U3753 (N_3753,N_3117,N_3108);
and U3754 (N_3754,N_3353,N_3175);
and U3755 (N_3755,N_3028,N_3068);
and U3756 (N_3756,N_3070,N_3491);
or U3757 (N_3757,N_3232,N_3153);
xnor U3758 (N_3758,N_3370,N_3455);
and U3759 (N_3759,N_3142,N_3414);
nand U3760 (N_3760,N_3478,N_3463);
and U3761 (N_3761,N_3177,N_3055);
nand U3762 (N_3762,N_3132,N_3492);
nand U3763 (N_3763,N_3284,N_3145);
and U3764 (N_3764,N_3295,N_3435);
nand U3765 (N_3765,N_3181,N_3177);
and U3766 (N_3766,N_3220,N_3330);
nand U3767 (N_3767,N_3456,N_3100);
or U3768 (N_3768,N_3257,N_3297);
and U3769 (N_3769,N_3408,N_3044);
nand U3770 (N_3770,N_3146,N_3064);
nor U3771 (N_3771,N_3226,N_3467);
and U3772 (N_3772,N_3032,N_3168);
xnor U3773 (N_3773,N_3403,N_3204);
or U3774 (N_3774,N_3427,N_3092);
nor U3775 (N_3775,N_3111,N_3329);
nand U3776 (N_3776,N_3135,N_3074);
nor U3777 (N_3777,N_3489,N_3453);
nand U3778 (N_3778,N_3270,N_3012);
nor U3779 (N_3779,N_3227,N_3334);
and U3780 (N_3780,N_3162,N_3303);
and U3781 (N_3781,N_3298,N_3235);
or U3782 (N_3782,N_3032,N_3031);
nor U3783 (N_3783,N_3261,N_3224);
nor U3784 (N_3784,N_3393,N_3035);
and U3785 (N_3785,N_3213,N_3059);
and U3786 (N_3786,N_3441,N_3234);
xor U3787 (N_3787,N_3461,N_3093);
and U3788 (N_3788,N_3173,N_3089);
xnor U3789 (N_3789,N_3242,N_3151);
and U3790 (N_3790,N_3091,N_3183);
xnor U3791 (N_3791,N_3104,N_3346);
and U3792 (N_3792,N_3052,N_3324);
and U3793 (N_3793,N_3318,N_3099);
nand U3794 (N_3794,N_3362,N_3283);
and U3795 (N_3795,N_3177,N_3462);
and U3796 (N_3796,N_3047,N_3408);
and U3797 (N_3797,N_3055,N_3482);
or U3798 (N_3798,N_3449,N_3172);
xnor U3799 (N_3799,N_3335,N_3255);
nor U3800 (N_3800,N_3056,N_3256);
or U3801 (N_3801,N_3302,N_3422);
nand U3802 (N_3802,N_3131,N_3424);
and U3803 (N_3803,N_3200,N_3087);
nor U3804 (N_3804,N_3417,N_3005);
and U3805 (N_3805,N_3302,N_3442);
and U3806 (N_3806,N_3045,N_3325);
nand U3807 (N_3807,N_3480,N_3210);
nand U3808 (N_3808,N_3040,N_3083);
nand U3809 (N_3809,N_3102,N_3031);
and U3810 (N_3810,N_3245,N_3200);
xnor U3811 (N_3811,N_3343,N_3383);
and U3812 (N_3812,N_3340,N_3266);
xnor U3813 (N_3813,N_3436,N_3143);
nor U3814 (N_3814,N_3245,N_3484);
or U3815 (N_3815,N_3033,N_3412);
and U3816 (N_3816,N_3078,N_3168);
and U3817 (N_3817,N_3074,N_3172);
or U3818 (N_3818,N_3150,N_3119);
xnor U3819 (N_3819,N_3339,N_3319);
and U3820 (N_3820,N_3368,N_3007);
nand U3821 (N_3821,N_3417,N_3194);
nor U3822 (N_3822,N_3101,N_3297);
nand U3823 (N_3823,N_3330,N_3030);
xor U3824 (N_3824,N_3399,N_3132);
nor U3825 (N_3825,N_3074,N_3335);
nand U3826 (N_3826,N_3189,N_3070);
nand U3827 (N_3827,N_3048,N_3234);
and U3828 (N_3828,N_3497,N_3114);
xnor U3829 (N_3829,N_3386,N_3018);
nand U3830 (N_3830,N_3413,N_3280);
nand U3831 (N_3831,N_3224,N_3106);
xor U3832 (N_3832,N_3455,N_3066);
nand U3833 (N_3833,N_3202,N_3034);
nor U3834 (N_3834,N_3218,N_3048);
nor U3835 (N_3835,N_3327,N_3484);
nor U3836 (N_3836,N_3267,N_3374);
nand U3837 (N_3837,N_3005,N_3199);
or U3838 (N_3838,N_3182,N_3223);
nor U3839 (N_3839,N_3010,N_3114);
and U3840 (N_3840,N_3410,N_3367);
and U3841 (N_3841,N_3274,N_3270);
and U3842 (N_3842,N_3355,N_3302);
nor U3843 (N_3843,N_3182,N_3323);
nand U3844 (N_3844,N_3219,N_3393);
and U3845 (N_3845,N_3188,N_3250);
and U3846 (N_3846,N_3343,N_3157);
nor U3847 (N_3847,N_3163,N_3457);
nor U3848 (N_3848,N_3310,N_3185);
xor U3849 (N_3849,N_3274,N_3340);
nand U3850 (N_3850,N_3119,N_3074);
xnor U3851 (N_3851,N_3258,N_3384);
nor U3852 (N_3852,N_3290,N_3220);
or U3853 (N_3853,N_3127,N_3409);
and U3854 (N_3854,N_3406,N_3077);
nand U3855 (N_3855,N_3130,N_3493);
nand U3856 (N_3856,N_3203,N_3104);
nor U3857 (N_3857,N_3034,N_3069);
or U3858 (N_3858,N_3416,N_3372);
xor U3859 (N_3859,N_3224,N_3305);
xnor U3860 (N_3860,N_3364,N_3441);
or U3861 (N_3861,N_3062,N_3093);
or U3862 (N_3862,N_3413,N_3372);
xnor U3863 (N_3863,N_3067,N_3195);
or U3864 (N_3864,N_3002,N_3383);
nand U3865 (N_3865,N_3166,N_3321);
nor U3866 (N_3866,N_3128,N_3443);
nand U3867 (N_3867,N_3138,N_3229);
xor U3868 (N_3868,N_3281,N_3028);
and U3869 (N_3869,N_3100,N_3174);
or U3870 (N_3870,N_3193,N_3461);
or U3871 (N_3871,N_3112,N_3088);
or U3872 (N_3872,N_3442,N_3299);
or U3873 (N_3873,N_3250,N_3234);
nand U3874 (N_3874,N_3464,N_3267);
xor U3875 (N_3875,N_3139,N_3452);
or U3876 (N_3876,N_3490,N_3164);
and U3877 (N_3877,N_3121,N_3042);
xor U3878 (N_3878,N_3294,N_3163);
nand U3879 (N_3879,N_3123,N_3317);
xnor U3880 (N_3880,N_3154,N_3363);
nor U3881 (N_3881,N_3006,N_3245);
nor U3882 (N_3882,N_3213,N_3230);
nand U3883 (N_3883,N_3325,N_3073);
and U3884 (N_3884,N_3199,N_3478);
xnor U3885 (N_3885,N_3302,N_3188);
xor U3886 (N_3886,N_3208,N_3097);
or U3887 (N_3887,N_3105,N_3335);
or U3888 (N_3888,N_3295,N_3184);
xnor U3889 (N_3889,N_3111,N_3380);
nor U3890 (N_3890,N_3061,N_3484);
nor U3891 (N_3891,N_3117,N_3410);
nor U3892 (N_3892,N_3356,N_3480);
xnor U3893 (N_3893,N_3344,N_3373);
nand U3894 (N_3894,N_3052,N_3335);
xor U3895 (N_3895,N_3484,N_3321);
and U3896 (N_3896,N_3180,N_3221);
and U3897 (N_3897,N_3197,N_3218);
xnor U3898 (N_3898,N_3436,N_3126);
nand U3899 (N_3899,N_3435,N_3117);
or U3900 (N_3900,N_3303,N_3246);
and U3901 (N_3901,N_3391,N_3413);
xor U3902 (N_3902,N_3204,N_3474);
or U3903 (N_3903,N_3432,N_3079);
nor U3904 (N_3904,N_3250,N_3010);
nand U3905 (N_3905,N_3470,N_3322);
nand U3906 (N_3906,N_3152,N_3313);
nor U3907 (N_3907,N_3090,N_3110);
nand U3908 (N_3908,N_3444,N_3158);
and U3909 (N_3909,N_3487,N_3179);
nand U3910 (N_3910,N_3394,N_3181);
nor U3911 (N_3911,N_3028,N_3209);
or U3912 (N_3912,N_3267,N_3346);
nand U3913 (N_3913,N_3290,N_3062);
xor U3914 (N_3914,N_3171,N_3188);
or U3915 (N_3915,N_3490,N_3477);
nor U3916 (N_3916,N_3026,N_3209);
and U3917 (N_3917,N_3379,N_3448);
nand U3918 (N_3918,N_3241,N_3401);
or U3919 (N_3919,N_3282,N_3347);
or U3920 (N_3920,N_3197,N_3241);
or U3921 (N_3921,N_3324,N_3451);
nand U3922 (N_3922,N_3494,N_3330);
nor U3923 (N_3923,N_3113,N_3415);
nand U3924 (N_3924,N_3418,N_3027);
xor U3925 (N_3925,N_3045,N_3232);
nand U3926 (N_3926,N_3177,N_3102);
or U3927 (N_3927,N_3069,N_3213);
nand U3928 (N_3928,N_3315,N_3432);
and U3929 (N_3929,N_3256,N_3132);
nand U3930 (N_3930,N_3000,N_3396);
and U3931 (N_3931,N_3151,N_3276);
xor U3932 (N_3932,N_3229,N_3207);
and U3933 (N_3933,N_3170,N_3102);
nand U3934 (N_3934,N_3402,N_3209);
or U3935 (N_3935,N_3407,N_3123);
nand U3936 (N_3936,N_3217,N_3240);
or U3937 (N_3937,N_3417,N_3235);
nand U3938 (N_3938,N_3057,N_3022);
xnor U3939 (N_3939,N_3018,N_3396);
and U3940 (N_3940,N_3331,N_3339);
nand U3941 (N_3941,N_3000,N_3378);
nand U3942 (N_3942,N_3378,N_3069);
nand U3943 (N_3943,N_3417,N_3225);
and U3944 (N_3944,N_3091,N_3469);
xnor U3945 (N_3945,N_3313,N_3430);
and U3946 (N_3946,N_3022,N_3234);
nand U3947 (N_3947,N_3430,N_3311);
and U3948 (N_3948,N_3111,N_3317);
and U3949 (N_3949,N_3149,N_3054);
nand U3950 (N_3950,N_3288,N_3376);
nor U3951 (N_3951,N_3361,N_3058);
xor U3952 (N_3952,N_3005,N_3120);
and U3953 (N_3953,N_3136,N_3002);
and U3954 (N_3954,N_3020,N_3342);
xor U3955 (N_3955,N_3071,N_3302);
xnor U3956 (N_3956,N_3475,N_3045);
or U3957 (N_3957,N_3226,N_3018);
nor U3958 (N_3958,N_3002,N_3288);
xor U3959 (N_3959,N_3287,N_3277);
and U3960 (N_3960,N_3136,N_3249);
nor U3961 (N_3961,N_3078,N_3479);
nand U3962 (N_3962,N_3272,N_3186);
nand U3963 (N_3963,N_3082,N_3168);
nand U3964 (N_3964,N_3064,N_3174);
nor U3965 (N_3965,N_3120,N_3441);
nor U3966 (N_3966,N_3159,N_3216);
or U3967 (N_3967,N_3449,N_3261);
xnor U3968 (N_3968,N_3180,N_3341);
and U3969 (N_3969,N_3348,N_3357);
or U3970 (N_3970,N_3082,N_3342);
or U3971 (N_3971,N_3283,N_3285);
or U3972 (N_3972,N_3398,N_3362);
and U3973 (N_3973,N_3318,N_3320);
or U3974 (N_3974,N_3480,N_3440);
nor U3975 (N_3975,N_3464,N_3011);
xnor U3976 (N_3976,N_3115,N_3449);
nor U3977 (N_3977,N_3377,N_3087);
and U3978 (N_3978,N_3463,N_3110);
nand U3979 (N_3979,N_3168,N_3318);
nor U3980 (N_3980,N_3196,N_3076);
nand U3981 (N_3981,N_3492,N_3459);
xor U3982 (N_3982,N_3405,N_3381);
or U3983 (N_3983,N_3264,N_3038);
or U3984 (N_3984,N_3184,N_3089);
nand U3985 (N_3985,N_3407,N_3413);
or U3986 (N_3986,N_3285,N_3049);
nor U3987 (N_3987,N_3374,N_3222);
nor U3988 (N_3988,N_3012,N_3319);
nand U3989 (N_3989,N_3302,N_3124);
xnor U3990 (N_3990,N_3465,N_3088);
or U3991 (N_3991,N_3362,N_3188);
or U3992 (N_3992,N_3260,N_3046);
or U3993 (N_3993,N_3353,N_3193);
and U3994 (N_3994,N_3027,N_3029);
nand U3995 (N_3995,N_3137,N_3074);
and U3996 (N_3996,N_3132,N_3170);
xor U3997 (N_3997,N_3348,N_3315);
nor U3998 (N_3998,N_3119,N_3430);
nand U3999 (N_3999,N_3428,N_3224);
and U4000 (N_4000,N_3842,N_3507);
nor U4001 (N_4001,N_3591,N_3856);
or U4002 (N_4002,N_3623,N_3931);
and U4003 (N_4003,N_3892,N_3697);
xnor U4004 (N_4004,N_3846,N_3734);
xnor U4005 (N_4005,N_3740,N_3940);
nand U4006 (N_4006,N_3612,N_3925);
xnor U4007 (N_4007,N_3943,N_3702);
and U4008 (N_4008,N_3561,N_3773);
and U4009 (N_4009,N_3744,N_3748);
or U4010 (N_4010,N_3954,N_3634);
xor U4011 (N_4011,N_3909,N_3535);
or U4012 (N_4012,N_3795,N_3516);
xor U4013 (N_4013,N_3813,N_3621);
or U4014 (N_4014,N_3839,N_3581);
or U4015 (N_4015,N_3917,N_3709);
or U4016 (N_4016,N_3999,N_3769);
and U4017 (N_4017,N_3731,N_3645);
and U4018 (N_4018,N_3970,N_3550);
or U4019 (N_4019,N_3721,N_3760);
and U4020 (N_4020,N_3725,N_3743);
nor U4021 (N_4021,N_3669,N_3872);
nand U4022 (N_4022,N_3800,N_3880);
xor U4023 (N_4023,N_3753,N_3891);
or U4024 (N_4024,N_3761,N_3907);
or U4025 (N_4025,N_3622,N_3831);
nor U4026 (N_4026,N_3936,N_3592);
nand U4027 (N_4027,N_3508,N_3662);
nand U4028 (N_4028,N_3884,N_3541);
and U4029 (N_4029,N_3780,N_3918);
xor U4030 (N_4030,N_3652,N_3549);
and U4031 (N_4031,N_3853,N_3902);
and U4032 (N_4032,N_3914,N_3804);
nand U4033 (N_4033,N_3688,N_3611);
xor U4034 (N_4034,N_3677,N_3716);
xor U4035 (N_4035,N_3826,N_3701);
xor U4036 (N_4036,N_3745,N_3724);
and U4037 (N_4037,N_3971,N_3871);
or U4038 (N_4038,N_3758,N_3674);
or U4039 (N_4039,N_3757,N_3765);
nand U4040 (N_4040,N_3963,N_3738);
nor U4041 (N_4041,N_3947,N_3997);
or U4042 (N_4042,N_3858,N_3503);
and U4043 (N_4043,N_3563,N_3961);
nor U4044 (N_4044,N_3567,N_3712);
nor U4045 (N_4045,N_3916,N_3610);
or U4046 (N_4046,N_3949,N_3861);
nor U4047 (N_4047,N_3819,N_3518);
nor U4048 (N_4048,N_3684,N_3569);
nor U4049 (N_4049,N_3723,N_3983);
or U4050 (N_4050,N_3635,N_3864);
nand U4051 (N_4051,N_3938,N_3806);
or U4052 (N_4052,N_3865,N_3633);
or U4053 (N_4053,N_3525,N_3548);
and U4054 (N_4054,N_3551,N_3703);
nand U4055 (N_4055,N_3718,N_3829);
nor U4056 (N_4056,N_3968,N_3735);
xnor U4057 (N_4057,N_3578,N_3692);
or U4058 (N_4058,N_3512,N_3899);
or U4059 (N_4059,N_3841,N_3542);
or U4060 (N_4060,N_3646,N_3589);
nor U4061 (N_4061,N_3523,N_3910);
nand U4062 (N_4062,N_3977,N_3720);
xnor U4063 (N_4063,N_3547,N_3650);
xnor U4064 (N_4064,N_3536,N_3615);
or U4065 (N_4065,N_3774,N_3572);
or U4066 (N_4066,N_3998,N_3875);
nor U4067 (N_4067,N_3568,N_3805);
and U4068 (N_4068,N_3691,N_3653);
or U4069 (N_4069,N_3895,N_3845);
xnor U4070 (N_4070,N_3717,N_3576);
or U4071 (N_4071,N_3617,N_3575);
xor U4072 (N_4072,N_3848,N_3739);
nor U4073 (N_4073,N_3501,N_3649);
nor U4074 (N_4074,N_3700,N_3854);
xor U4075 (N_4075,N_3832,N_3852);
nand U4076 (N_4076,N_3647,N_3671);
xnor U4077 (N_4077,N_3840,N_3678);
nor U4078 (N_4078,N_3526,N_3657);
nor U4079 (N_4079,N_3799,N_3510);
nand U4080 (N_4080,N_3851,N_3834);
nand U4081 (N_4081,N_3811,N_3596);
nand U4082 (N_4082,N_3866,N_3557);
xnor U4083 (N_4083,N_3582,N_3989);
xor U4084 (N_4084,N_3835,N_3893);
xnor U4085 (N_4085,N_3524,N_3887);
and U4086 (N_4086,N_3752,N_3641);
nor U4087 (N_4087,N_3620,N_3978);
nor U4088 (N_4088,N_3859,N_3616);
and U4089 (N_4089,N_3944,N_3539);
nor U4090 (N_4090,N_3517,N_3624);
nand U4091 (N_4091,N_3640,N_3915);
xor U4092 (N_4092,N_3544,N_3959);
xnor U4093 (N_4093,N_3877,N_3511);
or U4094 (N_4094,N_3791,N_3528);
nor U4095 (N_4095,N_3930,N_3847);
and U4096 (N_4096,N_3602,N_3537);
and U4097 (N_4097,N_3670,N_3981);
and U4098 (N_4098,N_3996,N_3682);
nor U4099 (N_4099,N_3975,N_3661);
or U4100 (N_4100,N_3911,N_3798);
xnor U4101 (N_4101,N_3986,N_3823);
nand U4102 (N_4102,N_3625,N_3704);
and U4103 (N_4103,N_3991,N_3782);
nand U4104 (N_4104,N_3648,N_3985);
and U4105 (N_4105,N_3945,N_3843);
and U4106 (N_4106,N_3824,N_3802);
or U4107 (N_4107,N_3500,N_3626);
or U4108 (N_4108,N_3600,N_3552);
and U4109 (N_4109,N_3787,N_3747);
nand U4110 (N_4110,N_3594,N_3900);
and U4111 (N_4111,N_3792,N_3584);
nor U4112 (N_4112,N_3808,N_3957);
xor U4113 (N_4113,N_3814,N_3862);
nand U4114 (N_4114,N_3637,N_3913);
xnor U4115 (N_4115,N_3663,N_3643);
nand U4116 (N_4116,N_3767,N_3816);
nor U4117 (N_4117,N_3570,N_3696);
nor U4118 (N_4118,N_3828,N_3574);
or U4119 (N_4119,N_3873,N_3759);
nand U4120 (N_4120,N_3545,N_3679);
nand U4121 (N_4121,N_3689,N_3726);
nor U4122 (N_4122,N_3651,N_3939);
nor U4123 (N_4123,N_3556,N_3972);
or U4124 (N_4124,N_3868,N_3710);
and U4125 (N_4125,N_3857,N_3553);
and U4126 (N_4126,N_3897,N_3778);
nand U4127 (N_4127,N_3715,N_3932);
xor U4128 (N_4128,N_3667,N_3719);
nor U4129 (N_4129,N_3789,N_3825);
nor U4130 (N_4130,N_3874,N_3713);
or U4131 (N_4131,N_3794,N_3830);
or U4132 (N_4132,N_3888,N_3807);
nand U4133 (N_4133,N_3527,N_3905);
or U4134 (N_4134,N_3706,N_3566);
nor U4135 (N_4135,N_3777,N_3966);
and U4136 (N_4136,N_3514,N_3733);
xor U4137 (N_4137,N_3521,N_3796);
xor U4138 (N_4138,N_3681,N_3630);
and U4139 (N_4139,N_3921,N_3749);
nand U4140 (N_4140,N_3515,N_3776);
or U4141 (N_4141,N_3506,N_3604);
xor U4142 (N_4142,N_3558,N_3520);
xnor U4143 (N_4143,N_3901,N_3564);
nor U4144 (N_4144,N_3827,N_3870);
nand U4145 (N_4145,N_3995,N_3598);
nor U4146 (N_4146,N_3699,N_3912);
or U4147 (N_4147,N_3967,N_3770);
xnor U4148 (N_4148,N_3766,N_3636);
nand U4149 (N_4149,N_3577,N_3976);
nand U4150 (N_4150,N_3755,N_3919);
nor U4151 (N_4151,N_3560,N_3929);
nor U4152 (N_4152,N_3964,N_3855);
nand U4153 (N_4153,N_3772,N_3965);
nand U4154 (N_4154,N_3573,N_3729);
xnor U4155 (N_4155,N_3942,N_3629);
and U4156 (N_4156,N_3613,N_3683);
xor U4157 (N_4157,N_3742,N_3941);
or U4158 (N_4158,N_3779,N_3922);
or U4159 (N_4159,N_3962,N_3987);
and U4160 (N_4160,N_3705,N_3898);
or U4161 (N_4161,N_3601,N_3658);
or U4162 (N_4162,N_3644,N_3937);
xnor U4163 (N_4163,N_3529,N_3934);
nand U4164 (N_4164,N_3756,N_3737);
xnor U4165 (N_4165,N_3894,N_3815);
nor U4166 (N_4166,N_3730,N_3953);
or U4167 (N_4167,N_3672,N_3546);
nor U4168 (N_4168,N_3890,N_3538);
nor U4169 (N_4169,N_3982,N_3979);
and U4170 (N_4170,N_3533,N_3605);
xnor U4171 (N_4171,N_3579,N_3952);
and U4172 (N_4172,N_3746,N_3849);
xor U4173 (N_4173,N_3708,N_3750);
xor U4174 (N_4174,N_3631,N_3509);
nand U4175 (N_4175,N_3906,N_3519);
nand U4176 (N_4176,N_3974,N_3803);
xor U4177 (N_4177,N_3793,N_3896);
nand U4178 (N_4178,N_3562,N_3768);
nand U4179 (N_4179,N_3958,N_3948);
nor U4180 (N_4180,N_3505,N_3883);
nor U4181 (N_4181,N_3994,N_3876);
xnor U4182 (N_4182,N_3775,N_3754);
nor U4183 (N_4183,N_3588,N_3513);
nor U4184 (N_4184,N_3614,N_3590);
nand U4185 (N_4185,N_3736,N_3531);
nor U4186 (N_4186,N_3889,N_3608);
nor U4187 (N_4187,N_3722,N_3786);
or U4188 (N_4188,N_3973,N_3522);
or U4189 (N_4189,N_3820,N_3585);
xor U4190 (N_4190,N_3781,N_3543);
and U4191 (N_4191,N_3502,N_3686);
or U4192 (N_4192,N_3728,N_3607);
and U4193 (N_4193,N_3869,N_3822);
xnor U4194 (N_4194,N_3580,N_3583);
or U4195 (N_4195,N_3727,N_3660);
nand U4196 (N_4196,N_3924,N_3530);
and U4197 (N_4197,N_3771,N_3821);
or U4198 (N_4198,N_3812,N_3593);
and U4199 (N_4199,N_3627,N_3693);
nand U4200 (N_4200,N_3599,N_3664);
nand U4201 (N_4201,N_3659,N_3764);
nand U4202 (N_4202,N_3988,N_3908);
xnor U4203 (N_4203,N_3790,N_3801);
nand U4204 (N_4204,N_3694,N_3980);
xnor U4205 (N_4205,N_3993,N_3879);
xnor U4206 (N_4206,N_3656,N_3655);
and U4207 (N_4207,N_3928,N_3878);
nand U4208 (N_4208,N_3885,N_3707);
xnor U4209 (N_4209,N_3837,N_3867);
nor U4210 (N_4210,N_3833,N_3540);
nor U4211 (N_4211,N_3609,N_3555);
xor U4212 (N_4212,N_3850,N_3860);
and U4213 (N_4213,N_3904,N_3817);
nand U4214 (N_4214,N_3763,N_3628);
or U4215 (N_4215,N_3685,N_3886);
nor U4216 (N_4216,N_3984,N_3638);
and U4217 (N_4217,N_3810,N_3619);
or U4218 (N_4218,N_3990,N_3687);
xor U4219 (N_4219,N_3595,N_3534);
and U4220 (N_4220,N_3668,N_3504);
nor U4221 (N_4221,N_3741,N_3935);
nor U4222 (N_4222,N_3698,N_3955);
xnor U4223 (N_4223,N_3732,N_3666);
or U4224 (N_4224,N_3923,N_3788);
xnor U4225 (N_4225,N_3642,N_3920);
or U4226 (N_4226,N_3680,N_3951);
nor U4227 (N_4227,N_3571,N_3797);
and U4228 (N_4228,N_3654,N_3784);
nor U4229 (N_4229,N_3844,N_3587);
nand U4230 (N_4230,N_3946,N_3926);
xnor U4231 (N_4231,N_3751,N_3863);
and U4232 (N_4232,N_3818,N_3695);
xnor U4233 (N_4233,N_3606,N_3618);
xnor U4234 (N_4234,N_3992,N_3950);
xnor U4235 (N_4235,N_3881,N_3690);
xnor U4236 (N_4236,N_3838,N_3639);
or U4237 (N_4237,N_3565,N_3676);
or U4238 (N_4238,N_3632,N_3836);
xnor U4239 (N_4239,N_3809,N_3960);
xor U4240 (N_4240,N_3559,N_3675);
and U4241 (N_4241,N_3586,N_3762);
nor U4242 (N_4242,N_3933,N_3597);
or U4243 (N_4243,N_3673,N_3882);
xor U4244 (N_4244,N_3783,N_3603);
or U4245 (N_4245,N_3554,N_3956);
xor U4246 (N_4246,N_3903,N_3665);
or U4247 (N_4247,N_3532,N_3714);
or U4248 (N_4248,N_3969,N_3785);
or U4249 (N_4249,N_3711,N_3927);
xor U4250 (N_4250,N_3556,N_3912);
nand U4251 (N_4251,N_3603,N_3613);
or U4252 (N_4252,N_3613,N_3700);
and U4253 (N_4253,N_3641,N_3594);
nand U4254 (N_4254,N_3654,N_3574);
and U4255 (N_4255,N_3898,N_3727);
xor U4256 (N_4256,N_3954,N_3723);
nand U4257 (N_4257,N_3522,N_3584);
xnor U4258 (N_4258,N_3956,N_3769);
or U4259 (N_4259,N_3865,N_3879);
and U4260 (N_4260,N_3537,N_3558);
or U4261 (N_4261,N_3782,N_3662);
xor U4262 (N_4262,N_3685,N_3631);
and U4263 (N_4263,N_3545,N_3586);
and U4264 (N_4264,N_3639,N_3833);
xor U4265 (N_4265,N_3844,N_3758);
nor U4266 (N_4266,N_3750,N_3831);
nor U4267 (N_4267,N_3625,N_3626);
nand U4268 (N_4268,N_3801,N_3985);
nor U4269 (N_4269,N_3633,N_3976);
nand U4270 (N_4270,N_3520,N_3811);
and U4271 (N_4271,N_3552,N_3734);
nand U4272 (N_4272,N_3926,N_3834);
nor U4273 (N_4273,N_3562,N_3933);
xnor U4274 (N_4274,N_3861,N_3536);
and U4275 (N_4275,N_3865,N_3569);
nand U4276 (N_4276,N_3651,N_3735);
xor U4277 (N_4277,N_3704,N_3831);
or U4278 (N_4278,N_3739,N_3564);
or U4279 (N_4279,N_3788,N_3940);
and U4280 (N_4280,N_3583,N_3699);
and U4281 (N_4281,N_3850,N_3703);
xnor U4282 (N_4282,N_3830,N_3750);
xor U4283 (N_4283,N_3972,N_3872);
nor U4284 (N_4284,N_3955,N_3984);
or U4285 (N_4285,N_3922,N_3842);
xnor U4286 (N_4286,N_3976,N_3628);
nand U4287 (N_4287,N_3877,N_3723);
nand U4288 (N_4288,N_3990,N_3880);
and U4289 (N_4289,N_3770,N_3950);
or U4290 (N_4290,N_3708,N_3729);
and U4291 (N_4291,N_3867,N_3893);
xor U4292 (N_4292,N_3765,N_3865);
nor U4293 (N_4293,N_3730,N_3661);
or U4294 (N_4294,N_3618,N_3796);
or U4295 (N_4295,N_3888,N_3712);
or U4296 (N_4296,N_3818,N_3847);
and U4297 (N_4297,N_3845,N_3535);
xnor U4298 (N_4298,N_3562,N_3826);
and U4299 (N_4299,N_3594,N_3962);
nor U4300 (N_4300,N_3891,N_3572);
or U4301 (N_4301,N_3516,N_3782);
xor U4302 (N_4302,N_3691,N_3568);
xnor U4303 (N_4303,N_3657,N_3506);
nor U4304 (N_4304,N_3635,N_3670);
nor U4305 (N_4305,N_3935,N_3853);
nand U4306 (N_4306,N_3753,N_3502);
and U4307 (N_4307,N_3613,N_3848);
nor U4308 (N_4308,N_3551,N_3524);
xnor U4309 (N_4309,N_3817,N_3541);
and U4310 (N_4310,N_3897,N_3681);
or U4311 (N_4311,N_3714,N_3591);
and U4312 (N_4312,N_3935,N_3838);
nor U4313 (N_4313,N_3625,N_3617);
nor U4314 (N_4314,N_3713,N_3922);
and U4315 (N_4315,N_3931,N_3750);
xnor U4316 (N_4316,N_3704,N_3729);
xor U4317 (N_4317,N_3503,N_3799);
or U4318 (N_4318,N_3990,N_3968);
nand U4319 (N_4319,N_3987,N_3984);
nor U4320 (N_4320,N_3781,N_3596);
and U4321 (N_4321,N_3887,N_3529);
and U4322 (N_4322,N_3894,N_3813);
nor U4323 (N_4323,N_3772,N_3628);
nor U4324 (N_4324,N_3889,N_3881);
nor U4325 (N_4325,N_3845,N_3886);
and U4326 (N_4326,N_3997,N_3759);
nand U4327 (N_4327,N_3895,N_3836);
xnor U4328 (N_4328,N_3984,N_3814);
or U4329 (N_4329,N_3714,N_3869);
or U4330 (N_4330,N_3927,N_3743);
nor U4331 (N_4331,N_3973,N_3559);
nor U4332 (N_4332,N_3766,N_3923);
and U4333 (N_4333,N_3549,N_3858);
or U4334 (N_4334,N_3799,N_3552);
xnor U4335 (N_4335,N_3641,N_3895);
xor U4336 (N_4336,N_3726,N_3848);
nand U4337 (N_4337,N_3714,N_3877);
or U4338 (N_4338,N_3665,N_3989);
or U4339 (N_4339,N_3842,N_3912);
xnor U4340 (N_4340,N_3939,N_3678);
nor U4341 (N_4341,N_3692,N_3589);
nor U4342 (N_4342,N_3629,N_3720);
nor U4343 (N_4343,N_3717,N_3698);
xor U4344 (N_4344,N_3551,N_3787);
and U4345 (N_4345,N_3567,N_3835);
xor U4346 (N_4346,N_3864,N_3538);
or U4347 (N_4347,N_3920,N_3970);
and U4348 (N_4348,N_3855,N_3780);
nor U4349 (N_4349,N_3645,N_3624);
or U4350 (N_4350,N_3786,N_3596);
xnor U4351 (N_4351,N_3724,N_3742);
xnor U4352 (N_4352,N_3949,N_3996);
xnor U4353 (N_4353,N_3512,N_3549);
or U4354 (N_4354,N_3599,N_3551);
nor U4355 (N_4355,N_3724,N_3798);
and U4356 (N_4356,N_3952,N_3768);
nand U4357 (N_4357,N_3961,N_3886);
and U4358 (N_4358,N_3876,N_3789);
nor U4359 (N_4359,N_3525,N_3930);
nand U4360 (N_4360,N_3672,N_3777);
nand U4361 (N_4361,N_3934,N_3919);
or U4362 (N_4362,N_3607,N_3945);
xnor U4363 (N_4363,N_3782,N_3500);
or U4364 (N_4364,N_3702,N_3897);
nor U4365 (N_4365,N_3930,N_3976);
xnor U4366 (N_4366,N_3962,N_3569);
or U4367 (N_4367,N_3663,N_3789);
and U4368 (N_4368,N_3586,N_3582);
and U4369 (N_4369,N_3943,N_3978);
and U4370 (N_4370,N_3972,N_3756);
and U4371 (N_4371,N_3708,N_3678);
nor U4372 (N_4372,N_3975,N_3511);
or U4373 (N_4373,N_3614,N_3798);
and U4374 (N_4374,N_3984,N_3616);
nand U4375 (N_4375,N_3622,N_3904);
or U4376 (N_4376,N_3516,N_3934);
nand U4377 (N_4377,N_3970,N_3816);
nand U4378 (N_4378,N_3982,N_3884);
xor U4379 (N_4379,N_3748,N_3514);
nor U4380 (N_4380,N_3578,N_3570);
nand U4381 (N_4381,N_3955,N_3766);
or U4382 (N_4382,N_3576,N_3608);
nand U4383 (N_4383,N_3646,N_3592);
nor U4384 (N_4384,N_3715,N_3547);
or U4385 (N_4385,N_3674,N_3792);
and U4386 (N_4386,N_3823,N_3672);
nor U4387 (N_4387,N_3845,N_3640);
or U4388 (N_4388,N_3899,N_3745);
nand U4389 (N_4389,N_3914,N_3980);
and U4390 (N_4390,N_3779,N_3729);
xnor U4391 (N_4391,N_3754,N_3630);
nand U4392 (N_4392,N_3986,N_3579);
nor U4393 (N_4393,N_3812,N_3936);
xor U4394 (N_4394,N_3774,N_3786);
xor U4395 (N_4395,N_3766,N_3799);
nor U4396 (N_4396,N_3899,N_3814);
xor U4397 (N_4397,N_3586,N_3780);
and U4398 (N_4398,N_3776,N_3768);
or U4399 (N_4399,N_3716,N_3592);
or U4400 (N_4400,N_3830,N_3711);
nor U4401 (N_4401,N_3737,N_3894);
nand U4402 (N_4402,N_3541,N_3557);
xnor U4403 (N_4403,N_3985,N_3892);
nand U4404 (N_4404,N_3729,N_3740);
nor U4405 (N_4405,N_3951,N_3739);
xnor U4406 (N_4406,N_3912,N_3658);
xnor U4407 (N_4407,N_3523,N_3575);
or U4408 (N_4408,N_3691,N_3859);
nand U4409 (N_4409,N_3699,N_3740);
nand U4410 (N_4410,N_3572,N_3576);
or U4411 (N_4411,N_3797,N_3912);
and U4412 (N_4412,N_3638,N_3949);
or U4413 (N_4413,N_3728,N_3635);
nor U4414 (N_4414,N_3640,N_3812);
nor U4415 (N_4415,N_3534,N_3848);
nor U4416 (N_4416,N_3974,N_3771);
xnor U4417 (N_4417,N_3782,N_3505);
nand U4418 (N_4418,N_3854,N_3761);
nor U4419 (N_4419,N_3985,N_3821);
xnor U4420 (N_4420,N_3536,N_3553);
nor U4421 (N_4421,N_3655,N_3765);
or U4422 (N_4422,N_3945,N_3591);
nand U4423 (N_4423,N_3849,N_3577);
nor U4424 (N_4424,N_3979,N_3521);
nor U4425 (N_4425,N_3673,N_3502);
nor U4426 (N_4426,N_3925,N_3555);
xor U4427 (N_4427,N_3821,N_3950);
nand U4428 (N_4428,N_3736,N_3681);
or U4429 (N_4429,N_3575,N_3825);
nor U4430 (N_4430,N_3902,N_3956);
nor U4431 (N_4431,N_3622,N_3555);
or U4432 (N_4432,N_3771,N_3885);
or U4433 (N_4433,N_3743,N_3514);
nand U4434 (N_4434,N_3839,N_3730);
nand U4435 (N_4435,N_3775,N_3818);
nor U4436 (N_4436,N_3666,N_3779);
xnor U4437 (N_4437,N_3519,N_3646);
nand U4438 (N_4438,N_3984,N_3973);
nand U4439 (N_4439,N_3795,N_3599);
nand U4440 (N_4440,N_3988,N_3826);
or U4441 (N_4441,N_3524,N_3888);
or U4442 (N_4442,N_3509,N_3988);
nand U4443 (N_4443,N_3923,N_3729);
and U4444 (N_4444,N_3528,N_3723);
nand U4445 (N_4445,N_3576,N_3787);
and U4446 (N_4446,N_3644,N_3648);
nand U4447 (N_4447,N_3703,N_3802);
nand U4448 (N_4448,N_3584,N_3814);
nor U4449 (N_4449,N_3793,N_3762);
and U4450 (N_4450,N_3739,N_3694);
or U4451 (N_4451,N_3924,N_3988);
xnor U4452 (N_4452,N_3932,N_3839);
xnor U4453 (N_4453,N_3647,N_3786);
xnor U4454 (N_4454,N_3886,N_3655);
nand U4455 (N_4455,N_3999,N_3840);
nor U4456 (N_4456,N_3756,N_3827);
nand U4457 (N_4457,N_3725,N_3712);
nand U4458 (N_4458,N_3994,N_3575);
nor U4459 (N_4459,N_3695,N_3688);
nor U4460 (N_4460,N_3596,N_3517);
nor U4461 (N_4461,N_3993,N_3715);
nand U4462 (N_4462,N_3965,N_3854);
nor U4463 (N_4463,N_3976,N_3870);
xor U4464 (N_4464,N_3579,N_3545);
nor U4465 (N_4465,N_3979,N_3556);
nand U4466 (N_4466,N_3972,N_3759);
nor U4467 (N_4467,N_3964,N_3531);
nor U4468 (N_4468,N_3913,N_3853);
xnor U4469 (N_4469,N_3538,N_3561);
or U4470 (N_4470,N_3667,N_3931);
or U4471 (N_4471,N_3846,N_3583);
and U4472 (N_4472,N_3883,N_3639);
or U4473 (N_4473,N_3787,N_3658);
and U4474 (N_4474,N_3704,N_3808);
nand U4475 (N_4475,N_3868,N_3717);
nand U4476 (N_4476,N_3818,N_3885);
xor U4477 (N_4477,N_3572,N_3784);
xor U4478 (N_4478,N_3569,N_3585);
nand U4479 (N_4479,N_3724,N_3574);
nor U4480 (N_4480,N_3639,N_3579);
nor U4481 (N_4481,N_3975,N_3569);
nor U4482 (N_4482,N_3674,N_3978);
nand U4483 (N_4483,N_3507,N_3746);
xnor U4484 (N_4484,N_3641,N_3987);
nor U4485 (N_4485,N_3829,N_3747);
nand U4486 (N_4486,N_3723,N_3648);
or U4487 (N_4487,N_3572,N_3806);
nand U4488 (N_4488,N_3741,N_3991);
nand U4489 (N_4489,N_3538,N_3727);
or U4490 (N_4490,N_3693,N_3895);
and U4491 (N_4491,N_3585,N_3784);
or U4492 (N_4492,N_3536,N_3865);
or U4493 (N_4493,N_3650,N_3590);
xor U4494 (N_4494,N_3590,N_3743);
nand U4495 (N_4495,N_3629,N_3510);
xor U4496 (N_4496,N_3759,N_3875);
xor U4497 (N_4497,N_3841,N_3605);
nand U4498 (N_4498,N_3717,N_3947);
or U4499 (N_4499,N_3963,N_3732);
and U4500 (N_4500,N_4094,N_4376);
and U4501 (N_4501,N_4130,N_4194);
or U4502 (N_4502,N_4444,N_4188);
and U4503 (N_4503,N_4328,N_4020);
xor U4504 (N_4504,N_4026,N_4414);
nand U4505 (N_4505,N_4406,N_4469);
nand U4506 (N_4506,N_4449,N_4385);
xnor U4507 (N_4507,N_4104,N_4079);
and U4508 (N_4508,N_4357,N_4486);
or U4509 (N_4509,N_4343,N_4342);
and U4510 (N_4510,N_4189,N_4454);
xor U4511 (N_4511,N_4157,N_4370);
xor U4512 (N_4512,N_4495,N_4181);
nor U4513 (N_4513,N_4143,N_4291);
nand U4514 (N_4514,N_4288,N_4299);
xnor U4515 (N_4515,N_4358,N_4464);
and U4516 (N_4516,N_4309,N_4246);
and U4517 (N_4517,N_4037,N_4416);
xnor U4518 (N_4518,N_4007,N_4493);
xor U4519 (N_4519,N_4412,N_4073);
nand U4520 (N_4520,N_4253,N_4098);
and U4521 (N_4521,N_4310,N_4336);
or U4522 (N_4522,N_4201,N_4019);
nand U4523 (N_4523,N_4408,N_4302);
or U4524 (N_4524,N_4002,N_4361);
xnor U4525 (N_4525,N_4295,N_4044);
or U4526 (N_4526,N_4040,N_4333);
nand U4527 (N_4527,N_4141,N_4455);
and U4528 (N_4528,N_4056,N_4351);
and U4529 (N_4529,N_4274,N_4331);
or U4530 (N_4530,N_4321,N_4476);
nand U4531 (N_4531,N_4364,N_4083);
and U4532 (N_4532,N_4437,N_4198);
xor U4533 (N_4533,N_4232,N_4137);
and U4534 (N_4534,N_4100,N_4413);
xor U4535 (N_4535,N_4147,N_4230);
nand U4536 (N_4536,N_4126,N_4494);
and U4537 (N_4537,N_4275,N_4018);
nand U4538 (N_4538,N_4380,N_4293);
or U4539 (N_4539,N_4210,N_4039);
xor U4540 (N_4540,N_4125,N_4059);
nor U4541 (N_4541,N_4430,N_4278);
nor U4542 (N_4542,N_4303,N_4187);
nand U4543 (N_4543,N_4021,N_4186);
and U4544 (N_4544,N_4255,N_4436);
and U4545 (N_4545,N_4145,N_4304);
xnor U4546 (N_4546,N_4123,N_4459);
xor U4547 (N_4547,N_4170,N_4359);
or U4548 (N_4548,N_4382,N_4131);
and U4549 (N_4549,N_4387,N_4216);
xnor U4550 (N_4550,N_4377,N_4393);
or U4551 (N_4551,N_4245,N_4330);
or U4552 (N_4552,N_4256,N_4050);
or U4553 (N_4553,N_4227,N_4270);
xnor U4554 (N_4554,N_4177,N_4116);
xor U4555 (N_4555,N_4159,N_4033);
nor U4556 (N_4556,N_4133,N_4067);
or U4557 (N_4557,N_4338,N_4499);
nand U4558 (N_4558,N_4207,N_4425);
or U4559 (N_4559,N_4167,N_4128);
or U4560 (N_4560,N_4114,N_4028);
nor U4561 (N_4561,N_4289,N_4399);
nand U4562 (N_4562,N_4443,N_4068);
xnor U4563 (N_4563,N_4217,N_4337);
or U4564 (N_4564,N_4318,N_4221);
xnor U4565 (N_4565,N_4488,N_4390);
and U4566 (N_4566,N_4322,N_4185);
nor U4567 (N_4567,N_4355,N_4257);
or U4568 (N_4568,N_4203,N_4320);
or U4569 (N_4569,N_4316,N_4268);
nor U4570 (N_4570,N_4281,N_4347);
xnor U4571 (N_4571,N_4162,N_4243);
nand U4572 (N_4572,N_4410,N_4372);
or U4573 (N_4573,N_4024,N_4031);
nor U4574 (N_4574,N_4086,N_4001);
and U4575 (N_4575,N_4060,N_4233);
xnor U4576 (N_4576,N_4264,N_4466);
and U4577 (N_4577,N_4280,N_4415);
nand U4578 (N_4578,N_4419,N_4052);
xnor U4579 (N_4579,N_4456,N_4082);
nand U4580 (N_4580,N_4152,N_4417);
nand U4581 (N_4581,N_4345,N_4065);
nor U4582 (N_4582,N_4122,N_4169);
or U4583 (N_4583,N_4247,N_4332);
nand U4584 (N_4584,N_4467,N_4009);
and U4585 (N_4585,N_4451,N_4151);
xnor U4586 (N_4586,N_4176,N_4150);
nand U4587 (N_4587,N_4120,N_4239);
or U4588 (N_4588,N_4090,N_4054);
and U4589 (N_4589,N_4206,N_4272);
or U4590 (N_4590,N_4038,N_4202);
xor U4591 (N_4591,N_4434,N_4356);
or U4592 (N_4592,N_4235,N_4146);
xnor U4593 (N_4593,N_4231,N_4213);
nor U4594 (N_4594,N_4395,N_4173);
nor U4595 (N_4595,N_4244,N_4062);
and U4596 (N_4596,N_4134,N_4315);
or U4597 (N_4597,N_4006,N_4371);
nor U4598 (N_4598,N_4214,N_4398);
nor U4599 (N_4599,N_4487,N_4142);
xnor U4600 (N_4600,N_4226,N_4097);
or U4601 (N_4601,N_4025,N_4103);
or U4602 (N_4602,N_4180,N_4388);
and U4603 (N_4603,N_4077,N_4057);
nand U4604 (N_4604,N_4386,N_4259);
xnor U4605 (N_4605,N_4403,N_4421);
and U4606 (N_4606,N_4129,N_4252);
and U4607 (N_4607,N_4363,N_4212);
nand U4608 (N_4608,N_4285,N_4383);
nand U4609 (N_4609,N_4089,N_4477);
xor U4610 (N_4610,N_4265,N_4135);
xor U4611 (N_4611,N_4424,N_4179);
and U4612 (N_4612,N_4117,N_4250);
nor U4613 (N_4613,N_4350,N_4153);
xor U4614 (N_4614,N_4271,N_4155);
nor U4615 (N_4615,N_4400,N_4029);
nand U4616 (N_4616,N_4475,N_4254);
nor U4617 (N_4617,N_4158,N_4010);
and U4618 (N_4618,N_4096,N_4016);
nor U4619 (N_4619,N_4045,N_4088);
nand U4620 (N_4620,N_4498,N_4258);
or U4621 (N_4621,N_4301,N_4081);
and U4622 (N_4622,N_4017,N_4085);
nand U4623 (N_4623,N_4327,N_4148);
xor U4624 (N_4624,N_4237,N_4394);
or U4625 (N_4625,N_4109,N_4178);
nor U4626 (N_4626,N_4470,N_4489);
nor U4627 (N_4627,N_4220,N_4209);
nor U4628 (N_4628,N_4360,N_4218);
and U4629 (N_4629,N_4340,N_4182);
and U4630 (N_4630,N_4119,N_4353);
nor U4631 (N_4631,N_4113,N_4277);
nor U4632 (N_4632,N_4108,N_4004);
or U4633 (N_4633,N_4426,N_4325);
xor U4634 (N_4634,N_4305,N_4276);
nand U4635 (N_4635,N_4111,N_4463);
nor U4636 (N_4636,N_4205,N_4481);
and U4637 (N_4637,N_4034,N_4228);
and U4638 (N_4638,N_4234,N_4296);
or U4639 (N_4639,N_4236,N_4204);
xor U4640 (N_4640,N_4047,N_4166);
nand U4641 (N_4641,N_4368,N_4314);
xor U4642 (N_4642,N_4012,N_4366);
or U4643 (N_4643,N_4431,N_4269);
xnor U4644 (N_4644,N_4461,N_4225);
or U4645 (N_4645,N_4238,N_4294);
or U4646 (N_4646,N_4460,N_4433);
or U4647 (N_4647,N_4248,N_4101);
or U4648 (N_4648,N_4080,N_4049);
nor U4649 (N_4649,N_4110,N_4384);
and U4650 (N_4650,N_4472,N_4215);
nand U4651 (N_4651,N_4492,N_4087);
xnor U4652 (N_4652,N_4267,N_4192);
xor U4653 (N_4653,N_4445,N_4106);
and U4654 (N_4654,N_4200,N_4480);
nand U4655 (N_4655,N_4334,N_4211);
nand U4656 (N_4656,N_4478,N_4136);
and U4657 (N_4657,N_4423,N_4251);
nor U4658 (N_4658,N_4219,N_4118);
xor U4659 (N_4659,N_4196,N_4442);
xor U4660 (N_4660,N_4319,N_4076);
nand U4661 (N_4661,N_4160,N_4174);
or U4662 (N_4662,N_4446,N_4300);
xnor U4663 (N_4663,N_4341,N_4263);
nand U4664 (N_4664,N_4354,N_4324);
nor U4665 (N_4665,N_4462,N_4308);
and U4666 (N_4666,N_4048,N_4290);
and U4667 (N_4667,N_4015,N_4323);
nor U4668 (N_4668,N_4420,N_4063);
or U4669 (N_4669,N_4409,N_4144);
nand U4670 (N_4670,N_4471,N_4042);
and U4671 (N_4671,N_4240,N_4043);
xnor U4672 (N_4672,N_4055,N_4389);
or U4673 (N_4673,N_4317,N_4069);
nor U4674 (N_4674,N_4241,N_4139);
nor U4675 (N_4675,N_4362,N_4473);
or U4676 (N_4676,N_4161,N_4132);
nand U4677 (N_4677,N_4095,N_4208);
xnor U4678 (N_4678,N_4344,N_4326);
and U4679 (N_4679,N_4313,N_4224);
and U4680 (N_4680,N_4051,N_4485);
nor U4681 (N_4681,N_4156,N_4286);
or U4682 (N_4682,N_4053,N_4283);
xor U4683 (N_4683,N_4392,N_4093);
and U4684 (N_4684,N_4438,N_4441);
xor U4685 (N_4685,N_4260,N_4003);
nand U4686 (N_4686,N_4497,N_4479);
and U4687 (N_4687,N_4484,N_4458);
and U4688 (N_4688,N_4391,N_4011);
or U4689 (N_4689,N_4222,N_4023);
and U4690 (N_4690,N_4292,N_4175);
xor U4691 (N_4691,N_4138,N_4022);
or U4692 (N_4692,N_4405,N_4307);
nor U4693 (N_4693,N_4261,N_4066);
nand U4694 (N_4694,N_4284,N_4105);
nand U4695 (N_4695,N_4164,N_4418);
and U4696 (N_4696,N_4035,N_4349);
or U4697 (N_4697,N_4163,N_4474);
and U4698 (N_4698,N_4422,N_4242);
nor U4699 (N_4699,N_4374,N_4199);
nor U4700 (N_4700,N_4071,N_4014);
xor U4701 (N_4701,N_4282,N_4072);
nand U4702 (N_4702,N_4032,N_4452);
nand U4703 (N_4703,N_4262,N_4183);
xor U4704 (N_4704,N_4378,N_4190);
nand U4705 (N_4705,N_4329,N_4468);
xnor U4706 (N_4706,N_4396,N_4064);
xor U4707 (N_4707,N_4084,N_4375);
xnor U4708 (N_4708,N_4482,N_4154);
or U4709 (N_4709,N_4172,N_4453);
and U4710 (N_4710,N_4448,N_4102);
or U4711 (N_4711,N_4490,N_4223);
or U4712 (N_4712,N_4457,N_4000);
nand U4713 (N_4713,N_4407,N_4184);
nand U4714 (N_4714,N_4483,N_4197);
xor U4715 (N_4715,N_4027,N_4058);
nand U4716 (N_4716,N_4099,N_4311);
or U4717 (N_4717,N_4149,N_4107);
or U4718 (N_4718,N_4041,N_4348);
nor U4719 (N_4719,N_4381,N_4429);
and U4720 (N_4720,N_4191,N_4140);
nand U4721 (N_4721,N_4121,N_4440);
and U4722 (N_4722,N_4411,N_4008);
nor U4723 (N_4723,N_4402,N_4091);
and U4724 (N_4724,N_4078,N_4312);
nand U4725 (N_4725,N_4365,N_4491);
nand U4726 (N_4726,N_4297,N_4061);
and U4727 (N_4727,N_4112,N_4171);
nor U4728 (N_4728,N_4124,N_4379);
and U4729 (N_4729,N_4127,N_4306);
or U4730 (N_4730,N_4013,N_4287);
nand U4731 (N_4731,N_4404,N_4273);
xor U4732 (N_4732,N_4229,N_4373);
nor U4733 (N_4733,N_4266,N_4030);
and U4734 (N_4734,N_4352,N_4193);
and U4735 (N_4735,N_4036,N_4168);
or U4736 (N_4736,N_4439,N_4046);
or U4737 (N_4737,N_4496,N_4279);
nor U4738 (N_4738,N_4195,N_4249);
nand U4739 (N_4739,N_4465,N_4432);
xor U4740 (N_4740,N_4335,N_4450);
nor U4741 (N_4741,N_4005,N_4369);
nand U4742 (N_4742,N_4339,N_4447);
nor U4743 (N_4743,N_4070,N_4346);
or U4744 (N_4744,N_4165,N_4115);
or U4745 (N_4745,N_4401,N_4367);
nand U4746 (N_4746,N_4092,N_4075);
and U4747 (N_4747,N_4428,N_4435);
or U4748 (N_4748,N_4298,N_4397);
nor U4749 (N_4749,N_4074,N_4427);
nor U4750 (N_4750,N_4409,N_4427);
or U4751 (N_4751,N_4222,N_4197);
xnor U4752 (N_4752,N_4439,N_4208);
nand U4753 (N_4753,N_4470,N_4067);
and U4754 (N_4754,N_4020,N_4141);
nand U4755 (N_4755,N_4415,N_4353);
xor U4756 (N_4756,N_4481,N_4372);
xor U4757 (N_4757,N_4166,N_4025);
nand U4758 (N_4758,N_4295,N_4098);
xnor U4759 (N_4759,N_4141,N_4254);
and U4760 (N_4760,N_4188,N_4310);
nor U4761 (N_4761,N_4166,N_4359);
or U4762 (N_4762,N_4272,N_4315);
or U4763 (N_4763,N_4198,N_4341);
xnor U4764 (N_4764,N_4321,N_4226);
nand U4765 (N_4765,N_4303,N_4222);
and U4766 (N_4766,N_4254,N_4402);
or U4767 (N_4767,N_4399,N_4306);
and U4768 (N_4768,N_4225,N_4337);
or U4769 (N_4769,N_4214,N_4466);
and U4770 (N_4770,N_4232,N_4428);
or U4771 (N_4771,N_4074,N_4475);
xor U4772 (N_4772,N_4070,N_4407);
xor U4773 (N_4773,N_4154,N_4110);
xor U4774 (N_4774,N_4138,N_4312);
nor U4775 (N_4775,N_4072,N_4482);
nor U4776 (N_4776,N_4084,N_4082);
xnor U4777 (N_4777,N_4377,N_4358);
nor U4778 (N_4778,N_4497,N_4446);
or U4779 (N_4779,N_4244,N_4168);
nor U4780 (N_4780,N_4066,N_4047);
xor U4781 (N_4781,N_4265,N_4214);
nand U4782 (N_4782,N_4118,N_4027);
xnor U4783 (N_4783,N_4205,N_4001);
or U4784 (N_4784,N_4299,N_4173);
nand U4785 (N_4785,N_4424,N_4270);
or U4786 (N_4786,N_4296,N_4388);
and U4787 (N_4787,N_4187,N_4142);
or U4788 (N_4788,N_4183,N_4251);
and U4789 (N_4789,N_4281,N_4431);
and U4790 (N_4790,N_4339,N_4191);
nor U4791 (N_4791,N_4200,N_4397);
xnor U4792 (N_4792,N_4262,N_4146);
or U4793 (N_4793,N_4142,N_4242);
or U4794 (N_4794,N_4291,N_4230);
or U4795 (N_4795,N_4123,N_4068);
or U4796 (N_4796,N_4296,N_4206);
nand U4797 (N_4797,N_4407,N_4420);
xor U4798 (N_4798,N_4165,N_4269);
xnor U4799 (N_4799,N_4080,N_4414);
xor U4800 (N_4800,N_4103,N_4208);
nor U4801 (N_4801,N_4071,N_4174);
or U4802 (N_4802,N_4189,N_4178);
xnor U4803 (N_4803,N_4344,N_4345);
nand U4804 (N_4804,N_4128,N_4457);
xnor U4805 (N_4805,N_4325,N_4448);
and U4806 (N_4806,N_4246,N_4088);
and U4807 (N_4807,N_4292,N_4481);
or U4808 (N_4808,N_4346,N_4017);
nor U4809 (N_4809,N_4286,N_4138);
or U4810 (N_4810,N_4308,N_4058);
xnor U4811 (N_4811,N_4382,N_4433);
nand U4812 (N_4812,N_4125,N_4025);
and U4813 (N_4813,N_4390,N_4095);
nand U4814 (N_4814,N_4214,N_4193);
xnor U4815 (N_4815,N_4306,N_4329);
and U4816 (N_4816,N_4222,N_4233);
xor U4817 (N_4817,N_4461,N_4150);
nand U4818 (N_4818,N_4182,N_4249);
or U4819 (N_4819,N_4491,N_4156);
nand U4820 (N_4820,N_4168,N_4098);
and U4821 (N_4821,N_4315,N_4127);
xnor U4822 (N_4822,N_4026,N_4270);
xor U4823 (N_4823,N_4162,N_4290);
and U4824 (N_4824,N_4385,N_4492);
nand U4825 (N_4825,N_4370,N_4321);
xor U4826 (N_4826,N_4000,N_4224);
nor U4827 (N_4827,N_4017,N_4342);
nand U4828 (N_4828,N_4454,N_4299);
nand U4829 (N_4829,N_4427,N_4028);
nor U4830 (N_4830,N_4414,N_4180);
nor U4831 (N_4831,N_4344,N_4042);
nor U4832 (N_4832,N_4050,N_4332);
nand U4833 (N_4833,N_4124,N_4049);
or U4834 (N_4834,N_4124,N_4277);
xor U4835 (N_4835,N_4416,N_4257);
or U4836 (N_4836,N_4083,N_4343);
nand U4837 (N_4837,N_4285,N_4218);
xor U4838 (N_4838,N_4479,N_4174);
or U4839 (N_4839,N_4278,N_4416);
nor U4840 (N_4840,N_4322,N_4051);
and U4841 (N_4841,N_4374,N_4127);
xnor U4842 (N_4842,N_4054,N_4112);
xor U4843 (N_4843,N_4450,N_4307);
xor U4844 (N_4844,N_4146,N_4008);
nand U4845 (N_4845,N_4444,N_4471);
nor U4846 (N_4846,N_4234,N_4304);
nand U4847 (N_4847,N_4314,N_4006);
or U4848 (N_4848,N_4305,N_4141);
and U4849 (N_4849,N_4194,N_4442);
and U4850 (N_4850,N_4267,N_4080);
and U4851 (N_4851,N_4094,N_4330);
or U4852 (N_4852,N_4138,N_4049);
and U4853 (N_4853,N_4026,N_4115);
and U4854 (N_4854,N_4241,N_4167);
or U4855 (N_4855,N_4495,N_4436);
nor U4856 (N_4856,N_4199,N_4362);
nand U4857 (N_4857,N_4059,N_4378);
and U4858 (N_4858,N_4472,N_4240);
and U4859 (N_4859,N_4491,N_4486);
and U4860 (N_4860,N_4247,N_4400);
or U4861 (N_4861,N_4268,N_4151);
nor U4862 (N_4862,N_4249,N_4269);
nand U4863 (N_4863,N_4472,N_4456);
or U4864 (N_4864,N_4246,N_4085);
or U4865 (N_4865,N_4357,N_4052);
or U4866 (N_4866,N_4189,N_4138);
xnor U4867 (N_4867,N_4169,N_4125);
xnor U4868 (N_4868,N_4227,N_4256);
nor U4869 (N_4869,N_4438,N_4339);
xnor U4870 (N_4870,N_4054,N_4332);
xnor U4871 (N_4871,N_4281,N_4019);
nand U4872 (N_4872,N_4298,N_4455);
nor U4873 (N_4873,N_4189,N_4469);
xnor U4874 (N_4874,N_4419,N_4079);
and U4875 (N_4875,N_4019,N_4137);
and U4876 (N_4876,N_4127,N_4196);
and U4877 (N_4877,N_4263,N_4350);
or U4878 (N_4878,N_4365,N_4316);
and U4879 (N_4879,N_4343,N_4044);
nor U4880 (N_4880,N_4193,N_4316);
xor U4881 (N_4881,N_4441,N_4076);
xnor U4882 (N_4882,N_4418,N_4014);
or U4883 (N_4883,N_4197,N_4051);
or U4884 (N_4884,N_4028,N_4274);
xnor U4885 (N_4885,N_4353,N_4078);
and U4886 (N_4886,N_4245,N_4340);
xor U4887 (N_4887,N_4121,N_4436);
nor U4888 (N_4888,N_4239,N_4469);
nand U4889 (N_4889,N_4010,N_4200);
and U4890 (N_4890,N_4132,N_4001);
and U4891 (N_4891,N_4334,N_4354);
nor U4892 (N_4892,N_4171,N_4330);
or U4893 (N_4893,N_4278,N_4440);
and U4894 (N_4894,N_4422,N_4469);
or U4895 (N_4895,N_4274,N_4138);
nand U4896 (N_4896,N_4256,N_4159);
nor U4897 (N_4897,N_4402,N_4465);
or U4898 (N_4898,N_4305,N_4243);
or U4899 (N_4899,N_4136,N_4473);
nor U4900 (N_4900,N_4109,N_4171);
nand U4901 (N_4901,N_4270,N_4066);
nor U4902 (N_4902,N_4496,N_4315);
xnor U4903 (N_4903,N_4316,N_4217);
nor U4904 (N_4904,N_4302,N_4018);
nor U4905 (N_4905,N_4192,N_4206);
or U4906 (N_4906,N_4479,N_4424);
xor U4907 (N_4907,N_4333,N_4350);
xnor U4908 (N_4908,N_4322,N_4419);
and U4909 (N_4909,N_4099,N_4166);
or U4910 (N_4910,N_4464,N_4317);
and U4911 (N_4911,N_4210,N_4404);
and U4912 (N_4912,N_4154,N_4079);
or U4913 (N_4913,N_4439,N_4165);
and U4914 (N_4914,N_4209,N_4082);
and U4915 (N_4915,N_4131,N_4470);
and U4916 (N_4916,N_4128,N_4054);
nand U4917 (N_4917,N_4338,N_4053);
or U4918 (N_4918,N_4328,N_4161);
nor U4919 (N_4919,N_4228,N_4211);
xnor U4920 (N_4920,N_4232,N_4222);
or U4921 (N_4921,N_4378,N_4328);
and U4922 (N_4922,N_4024,N_4227);
xnor U4923 (N_4923,N_4438,N_4194);
xnor U4924 (N_4924,N_4210,N_4064);
nand U4925 (N_4925,N_4485,N_4095);
and U4926 (N_4926,N_4015,N_4120);
and U4927 (N_4927,N_4356,N_4141);
nand U4928 (N_4928,N_4352,N_4167);
nor U4929 (N_4929,N_4374,N_4073);
and U4930 (N_4930,N_4063,N_4048);
nand U4931 (N_4931,N_4306,N_4323);
xnor U4932 (N_4932,N_4296,N_4342);
or U4933 (N_4933,N_4487,N_4338);
or U4934 (N_4934,N_4157,N_4132);
nand U4935 (N_4935,N_4152,N_4281);
nor U4936 (N_4936,N_4306,N_4208);
nor U4937 (N_4937,N_4265,N_4024);
xnor U4938 (N_4938,N_4299,N_4120);
and U4939 (N_4939,N_4411,N_4233);
nor U4940 (N_4940,N_4422,N_4211);
nand U4941 (N_4941,N_4428,N_4417);
nand U4942 (N_4942,N_4337,N_4304);
nor U4943 (N_4943,N_4337,N_4011);
and U4944 (N_4944,N_4154,N_4005);
nand U4945 (N_4945,N_4343,N_4095);
and U4946 (N_4946,N_4443,N_4302);
or U4947 (N_4947,N_4036,N_4233);
xnor U4948 (N_4948,N_4224,N_4070);
and U4949 (N_4949,N_4217,N_4158);
nand U4950 (N_4950,N_4121,N_4388);
or U4951 (N_4951,N_4268,N_4219);
nand U4952 (N_4952,N_4488,N_4251);
nand U4953 (N_4953,N_4319,N_4052);
nand U4954 (N_4954,N_4494,N_4401);
and U4955 (N_4955,N_4319,N_4140);
and U4956 (N_4956,N_4072,N_4331);
nand U4957 (N_4957,N_4472,N_4155);
nand U4958 (N_4958,N_4429,N_4181);
nand U4959 (N_4959,N_4233,N_4059);
or U4960 (N_4960,N_4396,N_4359);
and U4961 (N_4961,N_4439,N_4108);
and U4962 (N_4962,N_4499,N_4334);
or U4963 (N_4963,N_4014,N_4057);
and U4964 (N_4964,N_4025,N_4054);
or U4965 (N_4965,N_4347,N_4126);
nand U4966 (N_4966,N_4275,N_4052);
and U4967 (N_4967,N_4362,N_4024);
or U4968 (N_4968,N_4400,N_4267);
and U4969 (N_4969,N_4210,N_4296);
nand U4970 (N_4970,N_4123,N_4477);
nand U4971 (N_4971,N_4033,N_4210);
xor U4972 (N_4972,N_4212,N_4195);
or U4973 (N_4973,N_4410,N_4228);
nor U4974 (N_4974,N_4196,N_4071);
xnor U4975 (N_4975,N_4111,N_4146);
or U4976 (N_4976,N_4137,N_4440);
xor U4977 (N_4977,N_4069,N_4241);
nor U4978 (N_4978,N_4130,N_4222);
nor U4979 (N_4979,N_4249,N_4132);
and U4980 (N_4980,N_4412,N_4063);
nand U4981 (N_4981,N_4154,N_4277);
nor U4982 (N_4982,N_4286,N_4115);
nand U4983 (N_4983,N_4011,N_4121);
and U4984 (N_4984,N_4425,N_4209);
and U4985 (N_4985,N_4402,N_4274);
or U4986 (N_4986,N_4377,N_4263);
and U4987 (N_4987,N_4076,N_4100);
nor U4988 (N_4988,N_4330,N_4029);
nor U4989 (N_4989,N_4103,N_4276);
xnor U4990 (N_4990,N_4216,N_4444);
nor U4991 (N_4991,N_4121,N_4228);
xor U4992 (N_4992,N_4199,N_4348);
and U4993 (N_4993,N_4292,N_4056);
xnor U4994 (N_4994,N_4020,N_4003);
nand U4995 (N_4995,N_4113,N_4494);
nor U4996 (N_4996,N_4174,N_4224);
nor U4997 (N_4997,N_4267,N_4128);
xnor U4998 (N_4998,N_4370,N_4330);
xor U4999 (N_4999,N_4043,N_4361);
xor U5000 (N_5000,N_4951,N_4872);
nor U5001 (N_5001,N_4577,N_4965);
and U5002 (N_5002,N_4734,N_4950);
nor U5003 (N_5003,N_4569,N_4974);
and U5004 (N_5004,N_4810,N_4645);
and U5005 (N_5005,N_4861,N_4985);
or U5006 (N_5006,N_4797,N_4586);
or U5007 (N_5007,N_4643,N_4910);
nand U5008 (N_5008,N_4824,N_4812);
or U5009 (N_5009,N_4502,N_4845);
nand U5010 (N_5010,N_4952,N_4763);
nor U5011 (N_5011,N_4724,N_4543);
or U5012 (N_5012,N_4539,N_4510);
nor U5013 (N_5013,N_4942,N_4585);
nand U5014 (N_5014,N_4630,N_4752);
or U5015 (N_5015,N_4640,N_4730);
xor U5016 (N_5016,N_4878,N_4729);
or U5017 (N_5017,N_4975,N_4669);
or U5018 (N_5018,N_4789,N_4750);
and U5019 (N_5019,N_4979,N_4682);
xnor U5020 (N_5020,N_4527,N_4781);
nor U5021 (N_5021,N_4744,N_4567);
nor U5022 (N_5022,N_4604,N_4970);
and U5023 (N_5023,N_4707,N_4743);
and U5024 (N_5024,N_4868,N_4546);
or U5025 (N_5025,N_4946,N_4801);
nor U5026 (N_5026,N_4830,N_4825);
or U5027 (N_5027,N_4580,N_4613);
nor U5028 (N_5028,N_4826,N_4841);
and U5029 (N_5029,N_4737,N_4873);
nand U5030 (N_5030,N_4968,N_4513);
xor U5031 (N_5031,N_4815,N_4637);
nand U5032 (N_5032,N_4892,N_4887);
and U5033 (N_5033,N_4578,N_4501);
xnor U5034 (N_5034,N_4504,N_4927);
xnor U5035 (N_5035,N_4668,N_4600);
nor U5036 (N_5036,N_4639,N_4655);
xor U5037 (N_5037,N_4791,N_4686);
nand U5038 (N_5038,N_4780,N_4820);
xnor U5039 (N_5039,N_4902,N_4623);
nor U5040 (N_5040,N_4944,N_4949);
nor U5041 (N_5041,N_4762,N_4545);
and U5042 (N_5042,N_4904,N_4866);
nand U5043 (N_5043,N_4525,N_4774);
xor U5044 (N_5044,N_4976,N_4990);
nor U5045 (N_5045,N_4778,N_4628);
or U5046 (N_5046,N_4561,N_4701);
or U5047 (N_5047,N_4782,N_4665);
nand U5048 (N_5048,N_4775,N_4823);
nor U5049 (N_5049,N_4739,N_4692);
or U5050 (N_5050,N_4695,N_4533);
nand U5051 (N_5051,N_4874,N_4662);
xor U5052 (N_5052,N_4690,N_4936);
nand U5053 (N_5053,N_4940,N_4619);
and U5054 (N_5054,N_4846,N_4961);
nor U5055 (N_5055,N_4583,N_4827);
nor U5056 (N_5056,N_4538,N_4659);
xnor U5057 (N_5057,N_4786,N_4515);
and U5058 (N_5058,N_4829,N_4999);
or U5059 (N_5059,N_4671,N_4957);
and U5060 (N_5060,N_4636,N_4631);
nand U5061 (N_5061,N_4960,N_4652);
xnor U5062 (N_5062,N_4728,N_4749);
xor U5063 (N_5063,N_4733,N_4981);
and U5064 (N_5064,N_4656,N_4687);
nor U5065 (N_5065,N_4528,N_4712);
nor U5066 (N_5066,N_4530,N_4983);
nor U5067 (N_5067,N_4660,N_4865);
or U5068 (N_5068,N_4608,N_4647);
xor U5069 (N_5069,N_4986,N_4929);
and U5070 (N_5070,N_4971,N_4978);
nand U5071 (N_5071,N_4556,N_4703);
nand U5072 (N_5072,N_4776,N_4727);
nand U5073 (N_5073,N_4931,N_4955);
nand U5074 (N_5074,N_4560,N_4715);
and U5075 (N_5075,N_4787,N_4761);
nor U5076 (N_5076,N_4848,N_4984);
or U5077 (N_5077,N_4766,N_4633);
xnor U5078 (N_5078,N_4610,N_4685);
nor U5079 (N_5079,N_4783,N_4875);
xnor U5080 (N_5080,N_4666,N_4993);
nand U5081 (N_5081,N_4622,N_4948);
and U5082 (N_5082,N_4909,N_4954);
or U5083 (N_5083,N_4847,N_4511);
or U5084 (N_5084,N_4512,N_4748);
xnor U5085 (N_5085,N_4570,N_4885);
or U5086 (N_5086,N_4911,N_4813);
xor U5087 (N_5087,N_4764,N_4849);
or U5088 (N_5088,N_4680,N_4906);
nor U5089 (N_5089,N_4822,N_4895);
or U5090 (N_5090,N_4877,N_4907);
xnor U5091 (N_5091,N_4844,N_4657);
nand U5092 (N_5092,N_4616,N_4725);
xnor U5093 (N_5093,N_4593,N_4551);
or U5094 (N_5094,N_4842,N_4881);
or U5095 (N_5095,N_4856,N_4880);
nand U5096 (N_5096,N_4935,N_4629);
or U5097 (N_5097,N_4833,N_4765);
xnor U5098 (N_5098,N_4508,N_4535);
nor U5099 (N_5099,N_4700,N_4788);
and U5100 (N_5100,N_4507,N_4928);
or U5101 (N_5101,N_4839,N_4943);
xor U5102 (N_5102,N_4869,N_4925);
nor U5103 (N_5103,N_4916,N_4811);
nor U5104 (N_5104,N_4814,N_4799);
nor U5105 (N_5105,N_4723,N_4751);
nand U5106 (N_5106,N_4550,N_4972);
and U5107 (N_5107,N_4900,N_4796);
xor U5108 (N_5108,N_4930,N_4576);
nand U5109 (N_5109,N_4708,N_4720);
nor U5110 (N_5110,N_4590,N_4884);
xnor U5111 (N_5111,N_4571,N_4635);
xnor U5112 (N_5112,N_4641,N_4926);
or U5113 (N_5113,N_4518,N_4790);
or U5114 (N_5114,N_4973,N_4638);
and U5115 (N_5115,N_4644,N_4558);
nor U5116 (N_5116,N_4651,N_4836);
and U5117 (N_5117,N_4903,N_4611);
or U5118 (N_5118,N_4905,N_4777);
or U5119 (N_5119,N_4620,N_4650);
nand U5120 (N_5120,N_4614,N_4958);
nand U5121 (N_5121,N_4532,N_4771);
or U5122 (N_5122,N_4595,N_4514);
and U5123 (N_5123,N_4599,N_4860);
xor U5124 (N_5124,N_4838,N_4859);
nor U5125 (N_5125,N_4863,N_4832);
and U5126 (N_5126,N_4834,N_4584);
xnor U5127 (N_5127,N_4773,N_4582);
nand U5128 (N_5128,N_4718,N_4606);
xor U5129 (N_5129,N_4615,N_4785);
and U5130 (N_5130,N_4889,N_4563);
nor U5131 (N_5131,N_4805,N_4540);
xnor U5132 (N_5132,N_4573,N_4794);
xnor U5133 (N_5133,N_4520,N_4850);
nor U5134 (N_5134,N_4987,N_4964);
xnor U5135 (N_5135,N_4915,N_4517);
nor U5136 (N_5136,N_4617,N_4598);
xnor U5137 (N_5137,N_4531,N_4602);
nand U5138 (N_5138,N_4624,N_4988);
and U5139 (N_5139,N_4721,N_4760);
or U5140 (N_5140,N_4663,N_4867);
or U5141 (N_5141,N_4919,N_4607);
xor U5142 (N_5142,N_4956,N_4591);
nand U5143 (N_5143,N_4819,N_4557);
or U5144 (N_5144,N_4753,N_4800);
or U5145 (N_5145,N_4713,N_4821);
xnor U5146 (N_5146,N_4547,N_4882);
nand U5147 (N_5147,N_4677,N_4802);
or U5148 (N_5148,N_4989,N_4816);
nor U5149 (N_5149,N_4862,N_4793);
or U5150 (N_5150,N_4947,N_4843);
or U5151 (N_5151,N_4917,N_4853);
or U5152 (N_5152,N_4828,N_4977);
and U5153 (N_5153,N_4770,N_4597);
and U5154 (N_5154,N_4756,N_4691);
or U5155 (N_5155,N_4953,N_4592);
and U5156 (N_5156,N_4553,N_4982);
xnor U5157 (N_5157,N_4676,N_4642);
nor U5158 (N_5158,N_4831,N_4697);
or U5159 (N_5159,N_4534,N_4698);
and U5160 (N_5160,N_4678,N_4807);
nand U5161 (N_5161,N_4709,N_4879);
and U5162 (N_5162,N_4704,N_4516);
and U5163 (N_5163,N_4564,N_4893);
xor U5164 (N_5164,N_4719,N_4920);
and U5165 (N_5165,N_4738,N_4670);
nand U5166 (N_5166,N_4673,N_4541);
or U5167 (N_5167,N_4587,N_4932);
and U5168 (N_5168,N_4688,N_4552);
nand U5169 (N_5169,N_4526,N_4890);
xor U5170 (N_5170,N_4684,N_4536);
nand U5171 (N_5171,N_4529,N_4769);
and U5172 (N_5172,N_4858,N_4699);
nand U5173 (N_5173,N_4808,N_4896);
nor U5174 (N_5174,N_4609,N_4997);
and U5175 (N_5175,N_4959,N_4933);
or U5176 (N_5176,N_4711,N_4740);
or U5177 (N_5177,N_4693,N_4901);
and U5178 (N_5178,N_4555,N_4938);
or U5179 (N_5179,N_4649,N_4918);
nand U5180 (N_5180,N_4548,N_4664);
xor U5181 (N_5181,N_4646,N_4559);
and U5182 (N_5182,N_4694,N_4710);
nor U5183 (N_5183,N_4897,N_4996);
and U5184 (N_5184,N_4626,N_4746);
xor U5185 (N_5185,N_4992,N_4922);
or U5186 (N_5186,N_4566,N_4779);
nand U5187 (N_5187,N_4741,N_4579);
nor U5188 (N_5188,N_4894,N_4505);
nand U5189 (N_5189,N_4939,N_4735);
nand U5190 (N_5190,N_4913,N_4519);
xor U5191 (N_5191,N_4549,N_4809);
xnor U5192 (N_5192,N_4625,N_4632);
and U5193 (N_5193,N_4562,N_4731);
or U5194 (N_5194,N_4605,N_4742);
or U5195 (N_5195,N_4876,N_4565);
nand U5196 (N_5196,N_4689,N_4509);
or U5197 (N_5197,N_4716,N_4601);
xor U5198 (N_5198,N_4589,N_4835);
or U5199 (N_5199,N_4672,N_4870);
nor U5200 (N_5200,N_4732,N_4806);
nor U5201 (N_5201,N_4772,N_4798);
or U5202 (N_5202,N_4726,N_4705);
nand U5203 (N_5203,N_4803,N_4755);
and U5204 (N_5204,N_4544,N_4702);
nand U5205 (N_5205,N_4898,N_4851);
nor U5206 (N_5206,N_4854,N_4588);
xor U5207 (N_5207,N_4855,N_4658);
nand U5208 (N_5208,N_4594,N_4969);
xnor U5209 (N_5209,N_4500,N_4554);
nand U5210 (N_5210,N_4714,N_4722);
or U5211 (N_5211,N_4627,N_4980);
xnor U5212 (N_5212,N_4795,N_4914);
nand U5213 (N_5213,N_4994,N_4888);
and U5214 (N_5214,N_4792,N_4574);
xnor U5215 (N_5215,N_4891,N_4768);
nor U5216 (N_5216,N_4675,N_4581);
and U5217 (N_5217,N_4864,N_4661);
nor U5218 (N_5218,N_4522,N_4524);
and U5219 (N_5219,N_4817,N_4654);
and U5220 (N_5220,N_4945,N_4674);
and U5221 (N_5221,N_4937,N_4679);
nand U5222 (N_5222,N_4991,N_4568);
xor U5223 (N_5223,N_4621,N_4857);
nand U5224 (N_5224,N_4912,N_4852);
nand U5225 (N_5225,N_4908,N_4804);
and U5226 (N_5226,N_4921,N_4941);
nor U5227 (N_5227,N_4717,N_4634);
xor U5228 (N_5228,N_4871,N_4648);
xnor U5229 (N_5229,N_4963,N_4506);
xnor U5230 (N_5230,N_4934,N_4537);
or U5231 (N_5231,N_4757,N_4995);
nor U5232 (N_5232,N_4840,N_4618);
nor U5233 (N_5233,N_4572,N_4523);
and U5234 (N_5234,N_4924,N_4962);
nor U5235 (N_5235,N_4837,N_4747);
xor U5236 (N_5236,N_4998,N_4603);
nor U5237 (N_5237,N_4503,N_4967);
xnor U5238 (N_5238,N_4696,N_4542);
or U5239 (N_5239,N_4759,N_4653);
nand U5240 (N_5240,N_4758,N_4612);
xnor U5241 (N_5241,N_4784,N_4923);
and U5242 (N_5242,N_4818,N_4899);
and U5243 (N_5243,N_4575,N_4683);
nor U5244 (N_5244,N_4754,N_4596);
xnor U5245 (N_5245,N_4681,N_4767);
or U5246 (N_5246,N_4745,N_4883);
nand U5247 (N_5247,N_4736,N_4667);
nor U5248 (N_5248,N_4706,N_4966);
and U5249 (N_5249,N_4886,N_4521);
nand U5250 (N_5250,N_4979,N_4912);
nor U5251 (N_5251,N_4753,N_4805);
nor U5252 (N_5252,N_4670,N_4746);
or U5253 (N_5253,N_4765,N_4627);
xor U5254 (N_5254,N_4967,N_4985);
nor U5255 (N_5255,N_4602,N_4557);
and U5256 (N_5256,N_4781,N_4973);
nand U5257 (N_5257,N_4917,N_4620);
xor U5258 (N_5258,N_4607,N_4907);
nand U5259 (N_5259,N_4590,N_4525);
or U5260 (N_5260,N_4660,N_4991);
and U5261 (N_5261,N_4963,N_4753);
and U5262 (N_5262,N_4960,N_4713);
xnor U5263 (N_5263,N_4657,N_4767);
nand U5264 (N_5264,N_4648,N_4960);
xor U5265 (N_5265,N_4579,N_4653);
or U5266 (N_5266,N_4935,N_4850);
nand U5267 (N_5267,N_4748,N_4583);
or U5268 (N_5268,N_4579,N_4511);
and U5269 (N_5269,N_4691,N_4954);
or U5270 (N_5270,N_4710,N_4576);
or U5271 (N_5271,N_4928,N_4584);
or U5272 (N_5272,N_4942,N_4850);
and U5273 (N_5273,N_4673,N_4645);
nand U5274 (N_5274,N_4737,N_4866);
and U5275 (N_5275,N_4606,N_4599);
nor U5276 (N_5276,N_4686,N_4526);
nand U5277 (N_5277,N_4918,N_4866);
or U5278 (N_5278,N_4673,N_4945);
or U5279 (N_5279,N_4904,N_4617);
nor U5280 (N_5280,N_4920,N_4998);
or U5281 (N_5281,N_4835,N_4709);
nor U5282 (N_5282,N_4840,N_4685);
xor U5283 (N_5283,N_4695,N_4551);
or U5284 (N_5284,N_4658,N_4806);
and U5285 (N_5285,N_4756,N_4962);
or U5286 (N_5286,N_4975,N_4606);
xor U5287 (N_5287,N_4631,N_4795);
nand U5288 (N_5288,N_4935,N_4895);
or U5289 (N_5289,N_4651,N_4811);
and U5290 (N_5290,N_4889,N_4785);
and U5291 (N_5291,N_4797,N_4701);
and U5292 (N_5292,N_4745,N_4531);
nand U5293 (N_5293,N_4716,N_4948);
xor U5294 (N_5294,N_4969,N_4530);
nand U5295 (N_5295,N_4618,N_4930);
xnor U5296 (N_5296,N_4691,N_4818);
nor U5297 (N_5297,N_4809,N_4858);
xnor U5298 (N_5298,N_4829,N_4632);
nand U5299 (N_5299,N_4655,N_4528);
or U5300 (N_5300,N_4778,N_4664);
nand U5301 (N_5301,N_4578,N_4635);
or U5302 (N_5302,N_4899,N_4807);
nand U5303 (N_5303,N_4658,N_4809);
and U5304 (N_5304,N_4953,N_4975);
nor U5305 (N_5305,N_4884,N_4651);
xor U5306 (N_5306,N_4781,N_4916);
xor U5307 (N_5307,N_4852,N_4988);
nor U5308 (N_5308,N_4690,N_4772);
xnor U5309 (N_5309,N_4871,N_4850);
nand U5310 (N_5310,N_4784,N_4741);
nand U5311 (N_5311,N_4958,N_4995);
xor U5312 (N_5312,N_4663,N_4901);
and U5313 (N_5313,N_4515,N_4987);
or U5314 (N_5314,N_4566,N_4805);
and U5315 (N_5315,N_4847,N_4708);
or U5316 (N_5316,N_4816,N_4535);
or U5317 (N_5317,N_4531,N_4934);
and U5318 (N_5318,N_4836,N_4775);
or U5319 (N_5319,N_4754,N_4727);
or U5320 (N_5320,N_4551,N_4507);
or U5321 (N_5321,N_4835,N_4711);
nor U5322 (N_5322,N_4986,N_4606);
nor U5323 (N_5323,N_4847,N_4610);
xor U5324 (N_5324,N_4807,N_4993);
and U5325 (N_5325,N_4755,N_4895);
xnor U5326 (N_5326,N_4774,N_4802);
and U5327 (N_5327,N_4970,N_4762);
xor U5328 (N_5328,N_4966,N_4530);
nor U5329 (N_5329,N_4811,N_4776);
nand U5330 (N_5330,N_4789,N_4957);
nor U5331 (N_5331,N_4986,N_4738);
or U5332 (N_5332,N_4830,N_4726);
nand U5333 (N_5333,N_4881,N_4539);
and U5334 (N_5334,N_4573,N_4525);
nor U5335 (N_5335,N_4782,N_4852);
xor U5336 (N_5336,N_4794,N_4645);
or U5337 (N_5337,N_4921,N_4893);
nor U5338 (N_5338,N_4940,N_4594);
or U5339 (N_5339,N_4874,N_4960);
or U5340 (N_5340,N_4943,N_4583);
nor U5341 (N_5341,N_4904,N_4812);
xnor U5342 (N_5342,N_4598,N_4651);
or U5343 (N_5343,N_4803,N_4615);
nand U5344 (N_5344,N_4897,N_4825);
nand U5345 (N_5345,N_4843,N_4698);
nand U5346 (N_5346,N_4625,N_4602);
or U5347 (N_5347,N_4545,N_4596);
xor U5348 (N_5348,N_4566,N_4735);
nand U5349 (N_5349,N_4889,N_4863);
xnor U5350 (N_5350,N_4656,N_4972);
or U5351 (N_5351,N_4549,N_4963);
or U5352 (N_5352,N_4689,N_4759);
or U5353 (N_5353,N_4978,N_4770);
or U5354 (N_5354,N_4602,N_4521);
nand U5355 (N_5355,N_4562,N_4994);
or U5356 (N_5356,N_4709,N_4595);
nor U5357 (N_5357,N_4911,N_4555);
xnor U5358 (N_5358,N_4725,N_4522);
xor U5359 (N_5359,N_4979,N_4569);
xnor U5360 (N_5360,N_4702,N_4845);
nor U5361 (N_5361,N_4599,N_4621);
nand U5362 (N_5362,N_4708,N_4550);
or U5363 (N_5363,N_4710,N_4737);
nor U5364 (N_5364,N_4669,N_4523);
or U5365 (N_5365,N_4527,N_4598);
and U5366 (N_5366,N_4992,N_4941);
xnor U5367 (N_5367,N_4904,N_4883);
xor U5368 (N_5368,N_4759,N_4956);
nand U5369 (N_5369,N_4957,N_4750);
nor U5370 (N_5370,N_4671,N_4803);
xor U5371 (N_5371,N_4917,N_4969);
and U5372 (N_5372,N_4755,N_4561);
nor U5373 (N_5373,N_4854,N_4540);
nor U5374 (N_5374,N_4965,N_4792);
and U5375 (N_5375,N_4748,N_4735);
nor U5376 (N_5376,N_4729,N_4803);
xor U5377 (N_5377,N_4550,N_4979);
xor U5378 (N_5378,N_4768,N_4562);
nor U5379 (N_5379,N_4771,N_4681);
or U5380 (N_5380,N_4864,N_4507);
xnor U5381 (N_5381,N_4564,N_4786);
and U5382 (N_5382,N_4793,N_4969);
nand U5383 (N_5383,N_4598,N_4735);
or U5384 (N_5384,N_4629,N_4950);
nor U5385 (N_5385,N_4929,N_4799);
nand U5386 (N_5386,N_4673,N_4973);
nor U5387 (N_5387,N_4980,N_4691);
xor U5388 (N_5388,N_4895,N_4715);
nor U5389 (N_5389,N_4746,N_4868);
nand U5390 (N_5390,N_4914,N_4652);
or U5391 (N_5391,N_4503,N_4607);
xor U5392 (N_5392,N_4913,N_4762);
nand U5393 (N_5393,N_4548,N_4914);
nor U5394 (N_5394,N_4516,N_4793);
or U5395 (N_5395,N_4994,N_4702);
xnor U5396 (N_5396,N_4988,N_4555);
and U5397 (N_5397,N_4675,N_4560);
or U5398 (N_5398,N_4573,N_4510);
or U5399 (N_5399,N_4643,N_4599);
nor U5400 (N_5400,N_4706,N_4522);
and U5401 (N_5401,N_4712,N_4757);
nor U5402 (N_5402,N_4633,N_4878);
or U5403 (N_5403,N_4557,N_4826);
nor U5404 (N_5404,N_4808,N_4814);
and U5405 (N_5405,N_4969,N_4551);
or U5406 (N_5406,N_4687,N_4566);
or U5407 (N_5407,N_4873,N_4874);
or U5408 (N_5408,N_4821,N_4886);
or U5409 (N_5409,N_4832,N_4958);
and U5410 (N_5410,N_4975,N_4963);
nand U5411 (N_5411,N_4898,N_4722);
and U5412 (N_5412,N_4526,N_4803);
nor U5413 (N_5413,N_4701,N_4934);
nand U5414 (N_5414,N_4709,N_4845);
nor U5415 (N_5415,N_4817,N_4613);
or U5416 (N_5416,N_4623,N_4877);
nor U5417 (N_5417,N_4965,N_4849);
nand U5418 (N_5418,N_4950,N_4500);
and U5419 (N_5419,N_4860,N_4628);
and U5420 (N_5420,N_4941,N_4614);
xnor U5421 (N_5421,N_4915,N_4872);
and U5422 (N_5422,N_4796,N_4540);
nand U5423 (N_5423,N_4763,N_4894);
xnor U5424 (N_5424,N_4805,N_4899);
or U5425 (N_5425,N_4535,N_4840);
nand U5426 (N_5426,N_4667,N_4908);
and U5427 (N_5427,N_4836,N_4510);
nor U5428 (N_5428,N_4896,N_4845);
or U5429 (N_5429,N_4758,N_4600);
nor U5430 (N_5430,N_4973,N_4969);
and U5431 (N_5431,N_4556,N_4665);
nand U5432 (N_5432,N_4519,N_4822);
xnor U5433 (N_5433,N_4556,N_4911);
nand U5434 (N_5434,N_4976,N_4834);
xor U5435 (N_5435,N_4696,N_4883);
xor U5436 (N_5436,N_4936,N_4802);
nor U5437 (N_5437,N_4509,N_4936);
nand U5438 (N_5438,N_4644,N_4831);
or U5439 (N_5439,N_4793,N_4980);
or U5440 (N_5440,N_4700,N_4800);
nand U5441 (N_5441,N_4648,N_4643);
nand U5442 (N_5442,N_4889,N_4620);
and U5443 (N_5443,N_4668,N_4700);
nand U5444 (N_5444,N_4725,N_4872);
xor U5445 (N_5445,N_4726,N_4596);
xnor U5446 (N_5446,N_4601,N_4898);
nand U5447 (N_5447,N_4711,N_4816);
xnor U5448 (N_5448,N_4563,N_4542);
nor U5449 (N_5449,N_4779,N_4589);
or U5450 (N_5450,N_4593,N_4818);
or U5451 (N_5451,N_4780,N_4781);
or U5452 (N_5452,N_4569,N_4924);
or U5453 (N_5453,N_4652,N_4814);
nor U5454 (N_5454,N_4822,N_4521);
or U5455 (N_5455,N_4815,N_4622);
nor U5456 (N_5456,N_4950,N_4907);
and U5457 (N_5457,N_4601,N_4982);
nand U5458 (N_5458,N_4671,N_4879);
xnor U5459 (N_5459,N_4956,N_4778);
nor U5460 (N_5460,N_4999,N_4509);
xor U5461 (N_5461,N_4917,N_4600);
nor U5462 (N_5462,N_4790,N_4757);
xor U5463 (N_5463,N_4604,N_4804);
xnor U5464 (N_5464,N_4738,N_4860);
or U5465 (N_5465,N_4523,N_4963);
nor U5466 (N_5466,N_4590,N_4576);
and U5467 (N_5467,N_4527,N_4984);
and U5468 (N_5468,N_4621,N_4606);
and U5469 (N_5469,N_4858,N_4535);
xor U5470 (N_5470,N_4837,N_4567);
and U5471 (N_5471,N_4927,N_4699);
and U5472 (N_5472,N_4870,N_4910);
or U5473 (N_5473,N_4608,N_4576);
xnor U5474 (N_5474,N_4563,N_4533);
nor U5475 (N_5475,N_4512,N_4796);
xor U5476 (N_5476,N_4513,N_4876);
nand U5477 (N_5477,N_4531,N_4925);
or U5478 (N_5478,N_4980,N_4955);
xor U5479 (N_5479,N_4848,N_4722);
and U5480 (N_5480,N_4694,N_4636);
xor U5481 (N_5481,N_4608,N_4788);
or U5482 (N_5482,N_4652,N_4730);
and U5483 (N_5483,N_4933,N_4633);
xor U5484 (N_5484,N_4526,N_4811);
or U5485 (N_5485,N_4665,N_4593);
nor U5486 (N_5486,N_4870,N_4777);
xnor U5487 (N_5487,N_4641,N_4626);
or U5488 (N_5488,N_4926,N_4646);
or U5489 (N_5489,N_4623,N_4990);
nor U5490 (N_5490,N_4530,N_4682);
or U5491 (N_5491,N_4877,N_4713);
xor U5492 (N_5492,N_4949,N_4557);
or U5493 (N_5493,N_4728,N_4783);
nor U5494 (N_5494,N_4795,N_4698);
or U5495 (N_5495,N_4566,N_4869);
or U5496 (N_5496,N_4898,N_4787);
nand U5497 (N_5497,N_4802,N_4772);
or U5498 (N_5498,N_4657,N_4600);
or U5499 (N_5499,N_4925,N_4722);
xor U5500 (N_5500,N_5202,N_5122);
nand U5501 (N_5501,N_5413,N_5142);
nor U5502 (N_5502,N_5146,N_5438);
nand U5503 (N_5503,N_5174,N_5027);
and U5504 (N_5504,N_5215,N_5435);
and U5505 (N_5505,N_5424,N_5051);
and U5506 (N_5506,N_5071,N_5101);
and U5507 (N_5507,N_5035,N_5442);
and U5508 (N_5508,N_5437,N_5136);
nand U5509 (N_5509,N_5068,N_5197);
nand U5510 (N_5510,N_5496,N_5168);
nor U5511 (N_5511,N_5310,N_5107);
or U5512 (N_5512,N_5212,N_5133);
nor U5513 (N_5513,N_5388,N_5391);
xor U5514 (N_5514,N_5216,N_5063);
xnor U5515 (N_5515,N_5186,N_5259);
or U5516 (N_5516,N_5052,N_5324);
nand U5517 (N_5517,N_5015,N_5184);
and U5518 (N_5518,N_5139,N_5147);
and U5519 (N_5519,N_5152,N_5018);
nand U5520 (N_5520,N_5114,N_5355);
or U5521 (N_5521,N_5225,N_5099);
and U5522 (N_5522,N_5489,N_5112);
xnor U5523 (N_5523,N_5464,N_5246);
nand U5524 (N_5524,N_5214,N_5237);
and U5525 (N_5525,N_5299,N_5012);
xnor U5526 (N_5526,N_5157,N_5276);
or U5527 (N_5527,N_5378,N_5493);
and U5528 (N_5528,N_5195,N_5439);
or U5529 (N_5529,N_5316,N_5069);
nand U5530 (N_5530,N_5188,N_5308);
or U5531 (N_5531,N_5321,N_5406);
nand U5532 (N_5532,N_5042,N_5028);
nand U5533 (N_5533,N_5491,N_5089);
xnor U5534 (N_5534,N_5066,N_5292);
nand U5535 (N_5535,N_5084,N_5425);
nand U5536 (N_5536,N_5078,N_5016);
xnor U5537 (N_5537,N_5342,N_5135);
and U5538 (N_5538,N_5247,N_5148);
nand U5539 (N_5539,N_5492,N_5466);
nor U5540 (N_5540,N_5106,N_5248);
nor U5541 (N_5541,N_5185,N_5109);
nand U5542 (N_5542,N_5469,N_5362);
nor U5543 (N_5543,N_5095,N_5178);
nor U5544 (N_5544,N_5386,N_5271);
or U5545 (N_5545,N_5451,N_5262);
nand U5546 (N_5546,N_5023,N_5475);
and U5547 (N_5547,N_5367,N_5119);
or U5548 (N_5548,N_5088,N_5403);
nor U5549 (N_5549,N_5428,N_5251);
nor U5550 (N_5550,N_5243,N_5490);
or U5551 (N_5551,N_5346,N_5004);
or U5552 (N_5552,N_5264,N_5085);
or U5553 (N_5553,N_5477,N_5410);
xnor U5554 (N_5554,N_5010,N_5213);
xor U5555 (N_5555,N_5481,N_5319);
nand U5556 (N_5556,N_5008,N_5003);
and U5557 (N_5557,N_5427,N_5463);
xor U5558 (N_5558,N_5181,N_5453);
nor U5559 (N_5559,N_5080,N_5059);
or U5560 (N_5560,N_5098,N_5209);
or U5561 (N_5561,N_5141,N_5331);
xor U5562 (N_5562,N_5056,N_5171);
and U5563 (N_5563,N_5205,N_5250);
xnor U5564 (N_5564,N_5121,N_5289);
or U5565 (N_5565,N_5423,N_5011);
or U5566 (N_5566,N_5211,N_5086);
or U5567 (N_5567,N_5039,N_5232);
xnor U5568 (N_5568,N_5431,N_5175);
nor U5569 (N_5569,N_5082,N_5231);
and U5570 (N_5570,N_5207,N_5030);
nor U5571 (N_5571,N_5471,N_5034);
nand U5572 (N_5572,N_5091,N_5255);
or U5573 (N_5573,N_5499,N_5001);
and U5574 (N_5574,N_5260,N_5294);
nor U5575 (N_5575,N_5100,N_5094);
nor U5576 (N_5576,N_5019,N_5317);
xnor U5577 (N_5577,N_5291,N_5339);
or U5578 (N_5578,N_5313,N_5375);
nor U5579 (N_5579,N_5074,N_5105);
xor U5580 (N_5580,N_5358,N_5282);
or U5581 (N_5581,N_5046,N_5456);
nand U5582 (N_5582,N_5345,N_5445);
and U5583 (N_5583,N_5194,N_5239);
or U5584 (N_5584,N_5470,N_5049);
xnor U5585 (N_5585,N_5256,N_5199);
xnor U5586 (N_5586,N_5108,N_5222);
nor U5587 (N_5587,N_5269,N_5061);
nor U5588 (N_5588,N_5189,N_5238);
xor U5589 (N_5589,N_5393,N_5261);
xnor U5590 (N_5590,N_5155,N_5401);
nor U5591 (N_5591,N_5050,N_5409);
and U5592 (N_5592,N_5006,N_5405);
xor U5593 (N_5593,N_5138,N_5177);
and U5594 (N_5594,N_5065,N_5455);
or U5595 (N_5595,N_5240,N_5287);
nand U5596 (N_5596,N_5352,N_5433);
xnor U5597 (N_5597,N_5309,N_5395);
or U5598 (N_5598,N_5040,N_5480);
xnor U5599 (N_5599,N_5230,N_5187);
and U5600 (N_5600,N_5371,N_5130);
xor U5601 (N_5601,N_5379,N_5415);
or U5602 (N_5602,N_5322,N_5220);
nand U5603 (N_5603,N_5191,N_5092);
or U5604 (N_5604,N_5295,N_5278);
xnor U5605 (N_5605,N_5458,N_5103);
nor U5606 (N_5606,N_5485,N_5498);
nor U5607 (N_5607,N_5134,N_5219);
and U5608 (N_5608,N_5389,N_5311);
and U5609 (N_5609,N_5359,N_5173);
nand U5610 (N_5610,N_5430,N_5486);
nand U5611 (N_5611,N_5497,N_5380);
nand U5612 (N_5612,N_5446,N_5224);
and U5613 (N_5613,N_5307,N_5340);
nor U5614 (N_5614,N_5396,N_5303);
nor U5615 (N_5615,N_5318,N_5125);
nand U5616 (N_5616,N_5229,N_5400);
xnor U5617 (N_5617,N_5422,N_5000);
nor U5618 (N_5618,N_5038,N_5128);
and U5619 (N_5619,N_5387,N_5280);
or U5620 (N_5620,N_5296,N_5479);
and U5621 (N_5621,N_5143,N_5131);
nor U5622 (N_5622,N_5353,N_5418);
xnor U5623 (N_5623,N_5073,N_5198);
xor U5624 (N_5624,N_5279,N_5245);
xnor U5625 (N_5625,N_5167,N_5045);
or U5626 (N_5626,N_5154,N_5144);
or U5627 (N_5627,N_5033,N_5054);
or U5628 (N_5628,N_5356,N_5335);
nand U5629 (N_5629,N_5221,N_5366);
or U5630 (N_5630,N_5459,N_5460);
nor U5631 (N_5631,N_5283,N_5301);
nand U5632 (N_5632,N_5123,N_5163);
xor U5633 (N_5633,N_5162,N_5374);
nor U5634 (N_5634,N_5223,N_5273);
nor U5635 (N_5635,N_5032,N_5372);
and U5636 (N_5636,N_5160,N_5441);
xor U5637 (N_5637,N_5129,N_5031);
and U5638 (N_5638,N_5025,N_5275);
nor U5639 (N_5639,N_5377,N_5349);
and U5640 (N_5640,N_5081,N_5290);
or U5641 (N_5641,N_5265,N_5302);
or U5642 (N_5642,N_5270,N_5013);
and U5643 (N_5643,N_5233,N_5093);
and U5644 (N_5644,N_5210,N_5404);
or U5645 (N_5645,N_5036,N_5382);
nand U5646 (N_5646,N_5159,N_5151);
and U5647 (N_5647,N_5426,N_5126);
xnor U5648 (N_5648,N_5192,N_5258);
and U5649 (N_5649,N_5369,N_5137);
nand U5650 (N_5650,N_5457,N_5333);
nand U5651 (N_5651,N_5320,N_5312);
or U5652 (N_5652,N_5343,N_5483);
or U5653 (N_5653,N_5495,N_5452);
and U5654 (N_5654,N_5043,N_5293);
nand U5655 (N_5655,N_5272,N_5286);
or U5656 (N_5656,N_5115,N_5473);
or U5657 (N_5657,N_5204,N_5454);
nor U5658 (N_5658,N_5242,N_5416);
nand U5659 (N_5659,N_5300,N_5053);
and U5660 (N_5660,N_5326,N_5392);
or U5661 (N_5661,N_5044,N_5196);
or U5662 (N_5662,N_5076,N_5145);
or U5663 (N_5663,N_5474,N_5306);
or U5664 (N_5664,N_5060,N_5234);
nor U5665 (N_5665,N_5357,N_5487);
xor U5666 (N_5666,N_5421,N_5407);
nor U5667 (N_5667,N_5390,N_5048);
or U5668 (N_5668,N_5218,N_5315);
nor U5669 (N_5669,N_5017,N_5118);
or U5670 (N_5670,N_5370,N_5166);
or U5671 (N_5671,N_5104,N_5450);
xnor U5672 (N_5672,N_5236,N_5228);
nor U5673 (N_5673,N_5079,N_5170);
xor U5674 (N_5674,N_5005,N_5399);
or U5675 (N_5675,N_5444,N_5090);
nand U5676 (N_5676,N_5348,N_5361);
xnor U5677 (N_5677,N_5336,N_5014);
and U5678 (N_5678,N_5029,N_5385);
or U5679 (N_5679,N_5344,N_5411);
nand U5680 (N_5680,N_5206,N_5398);
nand U5681 (N_5681,N_5096,N_5200);
and U5682 (N_5682,N_5448,N_5288);
nand U5683 (N_5683,N_5443,N_5334);
nor U5684 (N_5684,N_5183,N_5179);
nand U5685 (N_5685,N_5140,N_5332);
and U5686 (N_5686,N_5111,N_5408);
nand U5687 (N_5687,N_5075,N_5341);
and U5688 (N_5688,N_5476,N_5329);
nor U5689 (N_5689,N_5007,N_5417);
and U5690 (N_5690,N_5298,N_5465);
or U5691 (N_5691,N_5077,N_5284);
xor U5692 (N_5692,N_5057,N_5203);
nor U5693 (N_5693,N_5462,N_5067);
or U5694 (N_5694,N_5235,N_5447);
or U5695 (N_5695,N_5420,N_5190);
xnor U5696 (N_5696,N_5024,N_5397);
nor U5697 (N_5697,N_5156,N_5472);
xnor U5698 (N_5698,N_5110,N_5161);
and U5699 (N_5699,N_5394,N_5150);
xnor U5700 (N_5700,N_5347,N_5325);
nor U5701 (N_5701,N_5263,N_5266);
nand U5702 (N_5702,N_5201,N_5097);
nor U5703 (N_5703,N_5120,N_5376);
nand U5704 (N_5704,N_5062,N_5281);
xnor U5705 (N_5705,N_5297,N_5305);
or U5706 (N_5706,N_5365,N_5338);
or U5707 (N_5707,N_5072,N_5373);
or U5708 (N_5708,N_5182,N_5037);
nand U5709 (N_5709,N_5440,N_5165);
xnor U5710 (N_5710,N_5381,N_5124);
xnor U5711 (N_5711,N_5327,N_5337);
nor U5712 (N_5712,N_5368,N_5217);
xor U5713 (N_5713,N_5083,N_5070);
xnor U5714 (N_5714,N_5468,N_5064);
and U5715 (N_5715,N_5172,N_5252);
or U5716 (N_5716,N_5314,N_5277);
nor U5717 (N_5717,N_5304,N_5022);
nand U5718 (N_5718,N_5208,N_5364);
nand U5719 (N_5719,N_5226,N_5384);
xnor U5720 (N_5720,N_5412,N_5047);
xnor U5721 (N_5721,N_5149,N_5116);
nand U5722 (N_5722,N_5020,N_5021);
nand U5723 (N_5723,N_5132,N_5002);
xnor U5724 (N_5724,N_5274,N_5488);
nand U5725 (N_5725,N_5127,N_5169);
xnor U5726 (N_5726,N_5419,N_5102);
nor U5727 (N_5727,N_5176,N_5434);
nor U5728 (N_5728,N_5323,N_5041);
nor U5729 (N_5729,N_5354,N_5402);
xor U5730 (N_5730,N_5268,N_5193);
nor U5731 (N_5731,N_5249,N_5153);
and U5732 (N_5732,N_5383,N_5227);
or U5733 (N_5733,N_5026,N_5241);
xnor U5734 (N_5734,N_5180,N_5436);
xor U5735 (N_5735,N_5267,N_5254);
nand U5736 (N_5736,N_5478,N_5461);
or U5737 (N_5737,N_5449,N_5285);
nand U5738 (N_5738,N_5113,N_5328);
nor U5739 (N_5739,N_5432,N_5482);
and U5740 (N_5740,N_5158,N_5484);
nand U5741 (N_5741,N_5350,N_5117);
nor U5742 (N_5742,N_5429,N_5244);
or U5743 (N_5743,N_5414,N_5055);
nand U5744 (N_5744,N_5087,N_5494);
nor U5745 (N_5745,N_5363,N_5360);
and U5746 (N_5746,N_5351,N_5253);
nor U5747 (N_5747,N_5058,N_5467);
nor U5748 (N_5748,N_5330,N_5009);
or U5749 (N_5749,N_5257,N_5164);
or U5750 (N_5750,N_5155,N_5282);
nor U5751 (N_5751,N_5492,N_5067);
xnor U5752 (N_5752,N_5249,N_5387);
and U5753 (N_5753,N_5151,N_5430);
and U5754 (N_5754,N_5069,N_5387);
nor U5755 (N_5755,N_5297,N_5264);
xnor U5756 (N_5756,N_5445,N_5105);
or U5757 (N_5757,N_5103,N_5373);
nand U5758 (N_5758,N_5041,N_5463);
and U5759 (N_5759,N_5080,N_5314);
or U5760 (N_5760,N_5218,N_5307);
xor U5761 (N_5761,N_5246,N_5244);
nand U5762 (N_5762,N_5121,N_5476);
nor U5763 (N_5763,N_5466,N_5288);
or U5764 (N_5764,N_5120,N_5231);
and U5765 (N_5765,N_5059,N_5240);
nand U5766 (N_5766,N_5082,N_5242);
xnor U5767 (N_5767,N_5447,N_5469);
nor U5768 (N_5768,N_5029,N_5405);
xor U5769 (N_5769,N_5248,N_5021);
nor U5770 (N_5770,N_5007,N_5400);
nand U5771 (N_5771,N_5004,N_5382);
xnor U5772 (N_5772,N_5003,N_5187);
nor U5773 (N_5773,N_5237,N_5314);
nor U5774 (N_5774,N_5183,N_5291);
xnor U5775 (N_5775,N_5138,N_5031);
nand U5776 (N_5776,N_5129,N_5385);
and U5777 (N_5777,N_5065,N_5004);
and U5778 (N_5778,N_5164,N_5278);
nand U5779 (N_5779,N_5128,N_5423);
or U5780 (N_5780,N_5066,N_5486);
nor U5781 (N_5781,N_5406,N_5472);
nand U5782 (N_5782,N_5050,N_5336);
xnor U5783 (N_5783,N_5015,N_5141);
or U5784 (N_5784,N_5332,N_5326);
nand U5785 (N_5785,N_5030,N_5397);
or U5786 (N_5786,N_5001,N_5154);
and U5787 (N_5787,N_5181,N_5252);
nand U5788 (N_5788,N_5432,N_5290);
nor U5789 (N_5789,N_5010,N_5282);
nand U5790 (N_5790,N_5473,N_5161);
nor U5791 (N_5791,N_5190,N_5178);
and U5792 (N_5792,N_5498,N_5444);
xnor U5793 (N_5793,N_5442,N_5309);
or U5794 (N_5794,N_5142,N_5078);
or U5795 (N_5795,N_5340,N_5150);
xnor U5796 (N_5796,N_5003,N_5055);
and U5797 (N_5797,N_5366,N_5016);
and U5798 (N_5798,N_5020,N_5093);
and U5799 (N_5799,N_5028,N_5131);
xor U5800 (N_5800,N_5425,N_5343);
or U5801 (N_5801,N_5117,N_5305);
xnor U5802 (N_5802,N_5356,N_5460);
nor U5803 (N_5803,N_5104,N_5381);
and U5804 (N_5804,N_5362,N_5129);
and U5805 (N_5805,N_5214,N_5384);
nor U5806 (N_5806,N_5417,N_5356);
and U5807 (N_5807,N_5084,N_5349);
and U5808 (N_5808,N_5271,N_5335);
nand U5809 (N_5809,N_5407,N_5313);
or U5810 (N_5810,N_5208,N_5247);
nand U5811 (N_5811,N_5337,N_5319);
or U5812 (N_5812,N_5399,N_5351);
nor U5813 (N_5813,N_5305,N_5419);
or U5814 (N_5814,N_5320,N_5103);
nand U5815 (N_5815,N_5124,N_5207);
or U5816 (N_5816,N_5072,N_5055);
xor U5817 (N_5817,N_5439,N_5277);
or U5818 (N_5818,N_5213,N_5107);
and U5819 (N_5819,N_5038,N_5408);
or U5820 (N_5820,N_5483,N_5361);
or U5821 (N_5821,N_5341,N_5358);
nor U5822 (N_5822,N_5047,N_5192);
and U5823 (N_5823,N_5472,N_5094);
nand U5824 (N_5824,N_5021,N_5454);
nor U5825 (N_5825,N_5446,N_5218);
nand U5826 (N_5826,N_5364,N_5167);
and U5827 (N_5827,N_5020,N_5293);
nor U5828 (N_5828,N_5329,N_5207);
nand U5829 (N_5829,N_5286,N_5085);
and U5830 (N_5830,N_5198,N_5159);
nand U5831 (N_5831,N_5105,N_5288);
and U5832 (N_5832,N_5186,N_5335);
xor U5833 (N_5833,N_5434,N_5283);
or U5834 (N_5834,N_5047,N_5304);
nand U5835 (N_5835,N_5473,N_5356);
and U5836 (N_5836,N_5314,N_5177);
or U5837 (N_5837,N_5162,N_5210);
and U5838 (N_5838,N_5479,N_5006);
nand U5839 (N_5839,N_5424,N_5198);
and U5840 (N_5840,N_5053,N_5337);
nor U5841 (N_5841,N_5425,N_5046);
nand U5842 (N_5842,N_5412,N_5438);
xnor U5843 (N_5843,N_5460,N_5020);
nand U5844 (N_5844,N_5179,N_5134);
nor U5845 (N_5845,N_5169,N_5008);
or U5846 (N_5846,N_5182,N_5243);
nand U5847 (N_5847,N_5234,N_5332);
and U5848 (N_5848,N_5084,N_5181);
nor U5849 (N_5849,N_5064,N_5183);
nand U5850 (N_5850,N_5014,N_5040);
nand U5851 (N_5851,N_5064,N_5192);
and U5852 (N_5852,N_5489,N_5016);
and U5853 (N_5853,N_5009,N_5433);
or U5854 (N_5854,N_5284,N_5231);
nand U5855 (N_5855,N_5045,N_5189);
xor U5856 (N_5856,N_5087,N_5355);
xnor U5857 (N_5857,N_5213,N_5293);
nor U5858 (N_5858,N_5032,N_5055);
nand U5859 (N_5859,N_5202,N_5074);
or U5860 (N_5860,N_5220,N_5238);
nand U5861 (N_5861,N_5201,N_5092);
nand U5862 (N_5862,N_5272,N_5462);
nor U5863 (N_5863,N_5476,N_5342);
or U5864 (N_5864,N_5356,N_5279);
and U5865 (N_5865,N_5137,N_5032);
nor U5866 (N_5866,N_5323,N_5121);
xor U5867 (N_5867,N_5144,N_5421);
or U5868 (N_5868,N_5127,N_5036);
nor U5869 (N_5869,N_5357,N_5378);
xor U5870 (N_5870,N_5237,N_5149);
xor U5871 (N_5871,N_5403,N_5266);
xor U5872 (N_5872,N_5137,N_5264);
xnor U5873 (N_5873,N_5057,N_5202);
and U5874 (N_5874,N_5282,N_5225);
xnor U5875 (N_5875,N_5427,N_5260);
or U5876 (N_5876,N_5301,N_5242);
and U5877 (N_5877,N_5130,N_5178);
nor U5878 (N_5878,N_5493,N_5376);
nand U5879 (N_5879,N_5023,N_5198);
and U5880 (N_5880,N_5080,N_5452);
nor U5881 (N_5881,N_5003,N_5311);
nand U5882 (N_5882,N_5172,N_5391);
nor U5883 (N_5883,N_5094,N_5351);
and U5884 (N_5884,N_5355,N_5276);
and U5885 (N_5885,N_5044,N_5346);
and U5886 (N_5886,N_5314,N_5488);
nand U5887 (N_5887,N_5313,N_5076);
and U5888 (N_5888,N_5087,N_5129);
nor U5889 (N_5889,N_5461,N_5120);
xor U5890 (N_5890,N_5499,N_5435);
and U5891 (N_5891,N_5348,N_5117);
nor U5892 (N_5892,N_5180,N_5421);
nand U5893 (N_5893,N_5419,N_5126);
or U5894 (N_5894,N_5112,N_5029);
or U5895 (N_5895,N_5055,N_5383);
nand U5896 (N_5896,N_5098,N_5155);
nand U5897 (N_5897,N_5128,N_5324);
and U5898 (N_5898,N_5300,N_5261);
or U5899 (N_5899,N_5361,N_5093);
nand U5900 (N_5900,N_5342,N_5258);
nor U5901 (N_5901,N_5033,N_5433);
nor U5902 (N_5902,N_5361,N_5353);
and U5903 (N_5903,N_5008,N_5357);
or U5904 (N_5904,N_5215,N_5471);
nor U5905 (N_5905,N_5327,N_5321);
nor U5906 (N_5906,N_5278,N_5137);
nand U5907 (N_5907,N_5374,N_5018);
xnor U5908 (N_5908,N_5432,N_5153);
xor U5909 (N_5909,N_5439,N_5051);
nand U5910 (N_5910,N_5135,N_5195);
and U5911 (N_5911,N_5012,N_5006);
nor U5912 (N_5912,N_5352,N_5475);
xor U5913 (N_5913,N_5315,N_5423);
xor U5914 (N_5914,N_5148,N_5299);
nand U5915 (N_5915,N_5225,N_5168);
nand U5916 (N_5916,N_5257,N_5326);
or U5917 (N_5917,N_5360,N_5454);
nand U5918 (N_5918,N_5370,N_5210);
or U5919 (N_5919,N_5319,N_5493);
xor U5920 (N_5920,N_5487,N_5235);
or U5921 (N_5921,N_5069,N_5483);
xnor U5922 (N_5922,N_5298,N_5253);
or U5923 (N_5923,N_5289,N_5128);
and U5924 (N_5924,N_5073,N_5255);
xor U5925 (N_5925,N_5042,N_5430);
or U5926 (N_5926,N_5382,N_5281);
or U5927 (N_5927,N_5207,N_5402);
nor U5928 (N_5928,N_5240,N_5185);
xnor U5929 (N_5929,N_5031,N_5319);
nor U5930 (N_5930,N_5373,N_5208);
or U5931 (N_5931,N_5361,N_5451);
or U5932 (N_5932,N_5188,N_5167);
or U5933 (N_5933,N_5123,N_5213);
or U5934 (N_5934,N_5193,N_5065);
xnor U5935 (N_5935,N_5220,N_5036);
or U5936 (N_5936,N_5134,N_5036);
and U5937 (N_5937,N_5135,N_5283);
xnor U5938 (N_5938,N_5180,N_5353);
or U5939 (N_5939,N_5386,N_5034);
or U5940 (N_5940,N_5174,N_5357);
and U5941 (N_5941,N_5153,N_5461);
nor U5942 (N_5942,N_5141,N_5137);
nor U5943 (N_5943,N_5172,N_5259);
nor U5944 (N_5944,N_5327,N_5465);
and U5945 (N_5945,N_5299,N_5265);
nor U5946 (N_5946,N_5479,N_5358);
or U5947 (N_5947,N_5139,N_5226);
nand U5948 (N_5948,N_5433,N_5167);
xnor U5949 (N_5949,N_5256,N_5070);
nor U5950 (N_5950,N_5104,N_5051);
xor U5951 (N_5951,N_5257,N_5440);
and U5952 (N_5952,N_5087,N_5266);
xor U5953 (N_5953,N_5357,N_5468);
xor U5954 (N_5954,N_5132,N_5206);
and U5955 (N_5955,N_5325,N_5315);
xnor U5956 (N_5956,N_5441,N_5009);
nor U5957 (N_5957,N_5307,N_5388);
nand U5958 (N_5958,N_5363,N_5042);
nand U5959 (N_5959,N_5093,N_5310);
nand U5960 (N_5960,N_5486,N_5299);
nor U5961 (N_5961,N_5310,N_5343);
and U5962 (N_5962,N_5068,N_5029);
xor U5963 (N_5963,N_5300,N_5363);
nand U5964 (N_5964,N_5373,N_5014);
nor U5965 (N_5965,N_5308,N_5256);
and U5966 (N_5966,N_5280,N_5017);
xnor U5967 (N_5967,N_5322,N_5364);
or U5968 (N_5968,N_5014,N_5131);
nor U5969 (N_5969,N_5016,N_5218);
nand U5970 (N_5970,N_5410,N_5065);
nand U5971 (N_5971,N_5234,N_5003);
or U5972 (N_5972,N_5378,N_5115);
xor U5973 (N_5973,N_5488,N_5378);
and U5974 (N_5974,N_5194,N_5023);
nand U5975 (N_5975,N_5255,N_5307);
nand U5976 (N_5976,N_5165,N_5429);
xnor U5977 (N_5977,N_5365,N_5280);
or U5978 (N_5978,N_5185,N_5289);
xnor U5979 (N_5979,N_5071,N_5450);
and U5980 (N_5980,N_5271,N_5344);
nand U5981 (N_5981,N_5197,N_5124);
nor U5982 (N_5982,N_5142,N_5140);
or U5983 (N_5983,N_5028,N_5232);
and U5984 (N_5984,N_5191,N_5282);
or U5985 (N_5985,N_5431,N_5196);
or U5986 (N_5986,N_5467,N_5165);
and U5987 (N_5987,N_5301,N_5016);
nor U5988 (N_5988,N_5205,N_5067);
nor U5989 (N_5989,N_5233,N_5314);
nand U5990 (N_5990,N_5321,N_5485);
and U5991 (N_5991,N_5169,N_5376);
nor U5992 (N_5992,N_5376,N_5206);
or U5993 (N_5993,N_5298,N_5204);
nand U5994 (N_5994,N_5006,N_5202);
nor U5995 (N_5995,N_5118,N_5225);
nor U5996 (N_5996,N_5214,N_5247);
xor U5997 (N_5997,N_5148,N_5220);
xnor U5998 (N_5998,N_5111,N_5383);
xnor U5999 (N_5999,N_5171,N_5448);
or U6000 (N_6000,N_5878,N_5630);
or U6001 (N_6001,N_5660,N_5749);
nand U6002 (N_6002,N_5599,N_5898);
nand U6003 (N_6003,N_5983,N_5782);
xor U6004 (N_6004,N_5729,N_5925);
or U6005 (N_6005,N_5927,N_5674);
xnor U6006 (N_6006,N_5512,N_5566);
nor U6007 (N_6007,N_5681,N_5994);
nor U6008 (N_6008,N_5569,N_5648);
xnor U6009 (N_6009,N_5704,N_5777);
xnor U6010 (N_6010,N_5572,N_5944);
nand U6011 (N_6011,N_5941,N_5862);
nand U6012 (N_6012,N_5707,N_5523);
nand U6013 (N_6013,N_5762,N_5905);
xnor U6014 (N_6014,N_5766,N_5594);
xor U6015 (N_6015,N_5595,N_5918);
nand U6016 (N_6016,N_5664,N_5814);
nand U6017 (N_6017,N_5682,N_5781);
or U6018 (N_6018,N_5529,N_5570);
xnor U6019 (N_6019,N_5635,N_5637);
nand U6020 (N_6020,N_5615,N_5913);
or U6021 (N_6021,N_5693,N_5860);
nor U6022 (N_6022,N_5536,N_5698);
and U6023 (N_6023,N_5550,N_5665);
nand U6024 (N_6024,N_5702,N_5916);
and U6025 (N_6025,N_5980,N_5919);
nor U6026 (N_6026,N_5624,N_5596);
xnor U6027 (N_6027,N_5593,N_5619);
and U6028 (N_6028,N_5845,N_5666);
xor U6029 (N_6029,N_5722,N_5575);
nor U6030 (N_6030,N_5700,N_5694);
xor U6031 (N_6031,N_5792,N_5757);
or U6032 (N_6032,N_5793,N_5894);
nor U6033 (N_6033,N_5640,N_5772);
and U6034 (N_6034,N_5826,N_5836);
nor U6035 (N_6035,N_5568,N_5577);
and U6036 (N_6036,N_5923,N_5554);
or U6037 (N_6037,N_5954,N_5824);
or U6038 (N_6038,N_5745,N_5855);
nor U6039 (N_6039,N_5991,N_5653);
xnor U6040 (N_6040,N_5758,N_5510);
and U6041 (N_6041,N_5920,N_5747);
xor U6042 (N_6042,N_5587,N_5671);
nand U6043 (N_6043,N_5579,N_5505);
xor U6044 (N_6044,N_5713,N_5932);
or U6045 (N_6045,N_5709,N_5879);
xor U6046 (N_6046,N_5813,N_5869);
nor U6047 (N_6047,N_5724,N_5688);
and U6048 (N_6048,N_5807,N_5975);
nor U6049 (N_6049,N_5833,N_5816);
xor U6050 (N_6050,N_5904,N_5746);
or U6051 (N_6051,N_5794,N_5958);
xnor U6052 (N_6052,N_5875,N_5931);
or U6053 (N_6053,N_5996,N_5884);
nor U6054 (N_6054,N_5810,N_5645);
or U6055 (N_6055,N_5684,N_5871);
or U6056 (N_6056,N_5502,N_5669);
nor U6057 (N_6057,N_5597,N_5525);
nor U6058 (N_6058,N_5830,N_5543);
xor U6059 (N_6059,N_5851,N_5728);
nor U6060 (N_6060,N_5842,N_5797);
xnor U6061 (N_6061,N_5679,N_5784);
nand U6062 (N_6062,N_5955,N_5541);
nand U6063 (N_6063,N_5610,N_5647);
nand U6064 (N_6064,N_5725,N_5573);
nand U6065 (N_6065,N_5985,N_5775);
xnor U6066 (N_6066,N_5734,N_5513);
nor U6067 (N_6067,N_5580,N_5960);
nand U6068 (N_6068,N_5945,N_5854);
xor U6069 (N_6069,N_5697,N_5534);
or U6070 (N_6070,N_5742,N_5730);
nand U6071 (N_6071,N_5533,N_5625);
nand U6072 (N_6072,N_5902,N_5685);
or U6073 (N_6073,N_5765,N_5504);
or U6074 (N_6074,N_5532,N_5803);
and U6075 (N_6075,N_5926,N_5809);
or U6076 (N_6076,N_5943,N_5780);
nand U6077 (N_6077,N_5893,N_5507);
xor U6078 (N_6078,N_5535,N_5603);
xnor U6079 (N_6079,N_5522,N_5719);
nand U6080 (N_6080,N_5652,N_5999);
nand U6081 (N_6081,N_5744,N_5825);
xnor U6082 (N_6082,N_5969,N_5618);
or U6083 (N_6083,N_5733,N_5576);
xnor U6084 (N_6084,N_5870,N_5859);
and U6085 (N_6085,N_5872,N_5956);
nor U6086 (N_6086,N_5658,N_5708);
xor U6087 (N_6087,N_5891,N_5874);
and U6088 (N_6088,N_5751,N_5548);
nor U6089 (N_6089,N_5578,N_5839);
nand U6090 (N_6090,N_5668,N_5558);
or U6091 (N_6091,N_5977,N_5804);
and U6092 (N_6092,N_5817,N_5514);
or U6093 (N_6093,N_5584,N_5656);
and U6094 (N_6094,N_5952,N_5583);
nor U6095 (N_6095,N_5538,N_5873);
nand U6096 (N_6096,N_5582,N_5695);
nor U6097 (N_6097,N_5808,N_5990);
nor U6098 (N_6098,N_5767,N_5776);
xor U6099 (N_6099,N_5831,N_5965);
xor U6100 (N_6100,N_5963,N_5720);
or U6101 (N_6101,N_5951,N_5606);
xor U6102 (N_6102,N_5737,N_5740);
or U6103 (N_6103,N_5616,N_5849);
and U6104 (N_6104,N_5520,N_5636);
and U6105 (N_6105,N_5946,N_5544);
nand U6106 (N_6106,N_5562,N_5663);
and U6107 (N_6107,N_5822,N_5799);
nor U6108 (N_6108,N_5667,N_5889);
xor U6109 (N_6109,N_5787,N_5815);
and U6110 (N_6110,N_5993,N_5614);
nand U6111 (N_6111,N_5989,N_5861);
nor U6112 (N_6112,N_5723,N_5511);
and U6113 (N_6113,N_5731,N_5646);
or U6114 (N_6114,N_5752,N_5771);
nor U6115 (N_6115,N_5892,N_5936);
nand U6116 (N_6116,N_5911,N_5612);
xor U6117 (N_6117,N_5828,N_5877);
nor U6118 (N_6118,N_5706,N_5853);
or U6119 (N_6119,N_5718,N_5800);
or U6120 (N_6120,N_5680,N_5967);
and U6121 (N_6121,N_5586,N_5978);
xnor U6122 (N_6122,N_5930,N_5526);
or U6123 (N_6123,N_5605,N_5938);
nor U6124 (N_6124,N_5712,N_5690);
nor U6125 (N_6125,N_5929,N_5542);
or U6126 (N_6126,N_5633,N_5796);
and U6127 (N_6127,N_5754,N_5617);
nor U6128 (N_6128,N_5769,N_5726);
xor U6129 (N_6129,N_5988,N_5632);
or U6130 (N_6130,N_5995,N_5838);
and U6131 (N_6131,N_5972,N_5974);
and U6132 (N_6132,N_5687,N_5959);
or U6133 (N_6133,N_5506,N_5966);
nand U6134 (N_6134,N_5834,N_5798);
xnor U6135 (N_6135,N_5638,N_5961);
or U6136 (N_6136,N_5973,N_5976);
and U6137 (N_6137,N_5546,N_5883);
and U6138 (N_6138,N_5736,N_5998);
nand U6139 (N_6139,N_5727,N_5968);
and U6140 (N_6140,N_5867,N_5866);
nand U6141 (N_6141,N_5773,N_5590);
nor U6142 (N_6142,N_5717,N_5739);
nand U6143 (N_6143,N_5649,N_5806);
nand U6144 (N_6144,N_5818,N_5805);
and U6145 (N_6145,N_5756,N_5785);
and U6146 (N_6146,N_5589,N_5759);
nand U6147 (N_6147,N_5992,N_5827);
xnor U6148 (N_6148,N_5984,N_5521);
and U6149 (N_6149,N_5858,N_5601);
nand U6150 (N_6150,N_5711,N_5527);
and U6151 (N_6151,N_5840,N_5627);
xor U6152 (N_6152,N_5942,N_5921);
nand U6153 (N_6153,N_5997,N_5686);
and U6154 (N_6154,N_5609,N_5516);
and U6155 (N_6155,N_5906,N_5598);
nor U6156 (N_6156,N_5829,N_5783);
nor U6157 (N_6157,N_5537,N_5934);
nor U6158 (N_6158,N_5567,N_5500);
nor U6159 (N_6159,N_5721,N_5837);
and U6160 (N_6160,N_5672,N_5949);
or U6161 (N_6161,N_5651,N_5947);
and U6162 (N_6162,N_5650,N_5670);
or U6163 (N_6163,N_5508,N_5795);
xnor U6164 (N_6164,N_5689,N_5865);
and U6165 (N_6165,N_5705,N_5540);
or U6166 (N_6166,N_5683,N_5556);
or U6167 (N_6167,N_5691,N_5547);
nor U6168 (N_6168,N_5900,N_5899);
or U6169 (N_6169,N_5701,N_5774);
xor U6170 (N_6170,N_5628,N_5802);
nand U6171 (N_6171,N_5852,N_5778);
xor U6172 (N_6172,N_5957,N_5574);
nand U6173 (N_6173,N_5761,N_5909);
or U6174 (N_6174,N_5864,N_5937);
and U6175 (N_6175,N_5788,N_5820);
xor U6176 (N_6176,N_5553,N_5885);
nor U6177 (N_6177,N_5501,N_5987);
nor U6178 (N_6178,N_5823,N_5981);
and U6179 (N_6179,N_5848,N_5979);
or U6180 (N_6180,N_5644,N_5716);
nand U6181 (N_6181,N_5524,N_5760);
or U6182 (N_6182,N_5912,N_5886);
nor U6183 (N_6183,N_5821,N_5801);
nor U6184 (N_6184,N_5897,N_5654);
or U6185 (N_6185,N_5673,N_5748);
nand U6186 (N_6186,N_5623,N_5655);
or U6187 (N_6187,N_5528,N_5950);
or U6188 (N_6188,N_5779,N_5518);
xor U6189 (N_6189,N_5642,N_5503);
xnor U6190 (N_6190,N_5560,N_5970);
nor U6191 (N_6191,N_5948,N_5868);
or U6192 (N_6192,N_5764,N_5850);
nand U6193 (N_6193,N_5592,N_5812);
and U6194 (N_6194,N_5847,N_5678);
xnor U6195 (N_6195,N_5895,N_5675);
xnor U6196 (N_6196,N_5602,N_5888);
xnor U6197 (N_6197,N_5515,N_5551);
nand U6198 (N_6198,N_5564,N_5585);
xnor U6199 (N_6199,N_5832,N_5621);
and U6200 (N_6200,N_5715,N_5661);
xnor U6201 (N_6201,N_5622,N_5843);
and U6202 (N_6202,N_5545,N_5928);
xnor U6203 (N_6203,N_5896,N_5581);
nand U6204 (N_6204,N_5743,N_5629);
or U6205 (N_6205,N_5791,N_5881);
or U6206 (N_6206,N_5657,N_5917);
xnor U6207 (N_6207,N_5908,N_5924);
nor U6208 (N_6208,N_5882,N_5753);
xnor U6209 (N_6209,N_5819,N_5571);
or U6210 (N_6210,N_5509,N_5933);
xor U6211 (N_6211,N_5953,N_5735);
or U6212 (N_6212,N_5922,N_5789);
nand U6213 (N_6213,N_5643,N_5863);
and U6214 (N_6214,N_5876,N_5530);
or U6215 (N_6215,N_5557,N_5841);
and U6216 (N_6216,N_5659,N_5631);
nor U6217 (N_6217,N_5790,N_5857);
nor U6218 (N_6218,N_5738,N_5964);
nand U6219 (N_6219,N_5750,N_5914);
nand U6220 (N_6220,N_5692,N_5768);
and U6221 (N_6221,N_5588,N_5835);
xor U6222 (N_6222,N_5626,N_5641);
and U6223 (N_6223,N_5517,N_5531);
xnor U6224 (N_6224,N_5608,N_5786);
nor U6225 (N_6225,N_5549,N_5676);
and U6226 (N_6226,N_5600,N_5741);
nor U6227 (N_6227,N_5846,N_5770);
xor U6228 (N_6228,N_5971,N_5519);
xor U6229 (N_6229,N_5607,N_5714);
xor U6230 (N_6230,N_5613,N_5710);
nand U6231 (N_6231,N_5639,N_5880);
and U6232 (N_6232,N_5962,N_5699);
and U6233 (N_6233,N_5986,N_5634);
nor U6234 (N_6234,N_5552,N_5939);
nand U6235 (N_6235,N_5662,N_5591);
and U6236 (N_6236,N_5935,N_5604);
and U6237 (N_6237,N_5696,N_5620);
nand U6238 (N_6238,N_5907,N_5563);
nand U6239 (N_6239,N_5677,N_5561);
xnor U6240 (N_6240,N_5755,N_5555);
xor U6241 (N_6241,N_5844,N_5611);
and U6242 (N_6242,N_5703,N_5901);
nor U6243 (N_6243,N_5915,N_5856);
or U6244 (N_6244,N_5903,N_5559);
or U6245 (N_6245,N_5763,N_5887);
nor U6246 (N_6246,N_5982,N_5565);
nand U6247 (N_6247,N_5539,N_5940);
or U6248 (N_6248,N_5732,N_5910);
xor U6249 (N_6249,N_5811,N_5890);
and U6250 (N_6250,N_5811,N_5546);
and U6251 (N_6251,N_5852,N_5555);
and U6252 (N_6252,N_5712,N_5634);
nor U6253 (N_6253,N_5782,N_5845);
or U6254 (N_6254,N_5780,N_5555);
xor U6255 (N_6255,N_5747,N_5895);
or U6256 (N_6256,N_5610,N_5816);
or U6257 (N_6257,N_5984,N_5651);
nor U6258 (N_6258,N_5777,N_5862);
nand U6259 (N_6259,N_5783,N_5636);
nand U6260 (N_6260,N_5912,N_5877);
and U6261 (N_6261,N_5888,N_5926);
xnor U6262 (N_6262,N_5555,N_5729);
or U6263 (N_6263,N_5841,N_5885);
nor U6264 (N_6264,N_5969,N_5756);
nor U6265 (N_6265,N_5669,N_5545);
nand U6266 (N_6266,N_5603,N_5640);
xor U6267 (N_6267,N_5570,N_5859);
nand U6268 (N_6268,N_5639,N_5537);
or U6269 (N_6269,N_5946,N_5529);
or U6270 (N_6270,N_5528,N_5620);
nor U6271 (N_6271,N_5913,N_5977);
nand U6272 (N_6272,N_5543,N_5892);
nor U6273 (N_6273,N_5933,N_5827);
and U6274 (N_6274,N_5634,N_5635);
and U6275 (N_6275,N_5994,N_5690);
nor U6276 (N_6276,N_5673,N_5521);
xor U6277 (N_6277,N_5840,N_5537);
or U6278 (N_6278,N_5602,N_5564);
and U6279 (N_6279,N_5562,N_5507);
or U6280 (N_6280,N_5631,N_5912);
or U6281 (N_6281,N_5535,N_5617);
nor U6282 (N_6282,N_5733,N_5800);
nor U6283 (N_6283,N_5789,N_5687);
nand U6284 (N_6284,N_5587,N_5845);
nand U6285 (N_6285,N_5644,N_5746);
nor U6286 (N_6286,N_5690,N_5630);
nor U6287 (N_6287,N_5586,N_5670);
or U6288 (N_6288,N_5738,N_5657);
nor U6289 (N_6289,N_5965,N_5671);
nor U6290 (N_6290,N_5941,N_5569);
nor U6291 (N_6291,N_5514,N_5853);
or U6292 (N_6292,N_5796,N_5819);
nor U6293 (N_6293,N_5575,N_5789);
or U6294 (N_6294,N_5841,N_5867);
and U6295 (N_6295,N_5787,N_5734);
and U6296 (N_6296,N_5973,N_5518);
or U6297 (N_6297,N_5686,N_5523);
or U6298 (N_6298,N_5877,N_5973);
or U6299 (N_6299,N_5503,N_5613);
or U6300 (N_6300,N_5577,N_5667);
xnor U6301 (N_6301,N_5732,N_5944);
nor U6302 (N_6302,N_5607,N_5588);
and U6303 (N_6303,N_5887,N_5549);
xnor U6304 (N_6304,N_5967,N_5781);
or U6305 (N_6305,N_5733,N_5774);
or U6306 (N_6306,N_5699,N_5536);
or U6307 (N_6307,N_5698,N_5576);
or U6308 (N_6308,N_5902,N_5545);
nor U6309 (N_6309,N_5876,N_5721);
nor U6310 (N_6310,N_5731,N_5909);
nor U6311 (N_6311,N_5690,N_5804);
and U6312 (N_6312,N_5559,N_5887);
or U6313 (N_6313,N_5919,N_5815);
or U6314 (N_6314,N_5904,N_5603);
or U6315 (N_6315,N_5991,N_5624);
nand U6316 (N_6316,N_5943,N_5612);
nor U6317 (N_6317,N_5813,N_5981);
or U6318 (N_6318,N_5842,N_5912);
nand U6319 (N_6319,N_5540,N_5818);
and U6320 (N_6320,N_5584,N_5934);
or U6321 (N_6321,N_5636,N_5671);
xor U6322 (N_6322,N_5760,N_5840);
or U6323 (N_6323,N_5786,N_5518);
and U6324 (N_6324,N_5759,N_5900);
nor U6325 (N_6325,N_5921,N_5859);
or U6326 (N_6326,N_5979,N_5650);
xor U6327 (N_6327,N_5537,N_5776);
nor U6328 (N_6328,N_5973,N_5913);
or U6329 (N_6329,N_5745,N_5853);
xor U6330 (N_6330,N_5540,N_5688);
and U6331 (N_6331,N_5991,N_5819);
nor U6332 (N_6332,N_5684,N_5810);
and U6333 (N_6333,N_5663,N_5968);
nand U6334 (N_6334,N_5786,N_5769);
nor U6335 (N_6335,N_5631,N_5543);
nor U6336 (N_6336,N_5615,N_5618);
or U6337 (N_6337,N_5784,N_5678);
nor U6338 (N_6338,N_5899,N_5684);
nand U6339 (N_6339,N_5627,N_5807);
and U6340 (N_6340,N_5892,N_5807);
xor U6341 (N_6341,N_5864,N_5535);
and U6342 (N_6342,N_5966,N_5501);
and U6343 (N_6343,N_5760,N_5832);
nor U6344 (N_6344,N_5803,N_5767);
nand U6345 (N_6345,N_5570,N_5975);
xnor U6346 (N_6346,N_5772,N_5646);
or U6347 (N_6347,N_5938,N_5752);
nor U6348 (N_6348,N_5792,N_5923);
and U6349 (N_6349,N_5892,N_5809);
nand U6350 (N_6350,N_5877,N_5524);
and U6351 (N_6351,N_5568,N_5700);
and U6352 (N_6352,N_5806,N_5878);
nand U6353 (N_6353,N_5631,N_5953);
or U6354 (N_6354,N_5962,N_5534);
nand U6355 (N_6355,N_5635,N_5864);
xnor U6356 (N_6356,N_5643,N_5860);
xor U6357 (N_6357,N_5592,N_5597);
nor U6358 (N_6358,N_5613,N_5608);
nand U6359 (N_6359,N_5942,N_5757);
nand U6360 (N_6360,N_5670,N_5575);
or U6361 (N_6361,N_5734,N_5815);
xnor U6362 (N_6362,N_5627,N_5693);
nand U6363 (N_6363,N_5557,N_5537);
or U6364 (N_6364,N_5593,N_5790);
or U6365 (N_6365,N_5600,N_5555);
nand U6366 (N_6366,N_5532,N_5995);
nor U6367 (N_6367,N_5523,N_5856);
nand U6368 (N_6368,N_5872,N_5750);
nand U6369 (N_6369,N_5634,N_5821);
nand U6370 (N_6370,N_5742,N_5940);
or U6371 (N_6371,N_5766,N_5695);
and U6372 (N_6372,N_5689,N_5805);
and U6373 (N_6373,N_5770,N_5992);
or U6374 (N_6374,N_5678,N_5892);
nor U6375 (N_6375,N_5714,N_5519);
nor U6376 (N_6376,N_5533,N_5549);
nand U6377 (N_6377,N_5644,N_5601);
nand U6378 (N_6378,N_5785,N_5861);
nand U6379 (N_6379,N_5992,N_5882);
or U6380 (N_6380,N_5977,N_5643);
nand U6381 (N_6381,N_5936,N_5732);
and U6382 (N_6382,N_5942,N_5870);
or U6383 (N_6383,N_5920,N_5918);
nand U6384 (N_6384,N_5795,N_5761);
nand U6385 (N_6385,N_5579,N_5930);
nand U6386 (N_6386,N_5827,N_5988);
and U6387 (N_6387,N_5626,N_5660);
xor U6388 (N_6388,N_5772,N_5727);
or U6389 (N_6389,N_5607,N_5999);
nand U6390 (N_6390,N_5516,N_5700);
nor U6391 (N_6391,N_5835,N_5727);
xnor U6392 (N_6392,N_5667,N_5747);
or U6393 (N_6393,N_5728,N_5898);
nor U6394 (N_6394,N_5560,N_5558);
nand U6395 (N_6395,N_5877,N_5695);
or U6396 (N_6396,N_5616,N_5776);
xnor U6397 (N_6397,N_5705,N_5707);
nand U6398 (N_6398,N_5667,N_5758);
xor U6399 (N_6399,N_5943,N_5879);
or U6400 (N_6400,N_5767,N_5682);
nor U6401 (N_6401,N_5598,N_5812);
and U6402 (N_6402,N_5818,N_5732);
or U6403 (N_6403,N_5859,N_5917);
or U6404 (N_6404,N_5763,N_5639);
nor U6405 (N_6405,N_5839,N_5525);
and U6406 (N_6406,N_5739,N_5977);
or U6407 (N_6407,N_5915,N_5604);
or U6408 (N_6408,N_5931,N_5800);
and U6409 (N_6409,N_5633,N_5745);
or U6410 (N_6410,N_5557,N_5514);
and U6411 (N_6411,N_5662,N_5924);
or U6412 (N_6412,N_5980,N_5744);
xor U6413 (N_6413,N_5579,N_5706);
nor U6414 (N_6414,N_5876,N_5781);
or U6415 (N_6415,N_5560,N_5952);
xor U6416 (N_6416,N_5849,N_5547);
xor U6417 (N_6417,N_5512,N_5923);
or U6418 (N_6418,N_5580,N_5594);
or U6419 (N_6419,N_5815,N_5657);
xnor U6420 (N_6420,N_5703,N_5671);
xnor U6421 (N_6421,N_5927,N_5614);
nor U6422 (N_6422,N_5793,N_5935);
and U6423 (N_6423,N_5885,N_5578);
nand U6424 (N_6424,N_5531,N_5777);
xnor U6425 (N_6425,N_5543,N_5719);
and U6426 (N_6426,N_5842,N_5731);
and U6427 (N_6427,N_5932,N_5923);
and U6428 (N_6428,N_5925,N_5709);
xnor U6429 (N_6429,N_5639,N_5571);
or U6430 (N_6430,N_5585,N_5974);
and U6431 (N_6431,N_5832,N_5636);
xnor U6432 (N_6432,N_5775,N_5641);
or U6433 (N_6433,N_5826,N_5560);
and U6434 (N_6434,N_5791,N_5932);
and U6435 (N_6435,N_5776,N_5565);
xor U6436 (N_6436,N_5670,N_5592);
nand U6437 (N_6437,N_5512,N_5724);
nand U6438 (N_6438,N_5962,N_5649);
nand U6439 (N_6439,N_5527,N_5977);
nor U6440 (N_6440,N_5680,N_5768);
and U6441 (N_6441,N_5599,N_5825);
nor U6442 (N_6442,N_5746,N_5801);
nor U6443 (N_6443,N_5985,N_5625);
nor U6444 (N_6444,N_5505,N_5907);
nand U6445 (N_6445,N_5526,N_5819);
xnor U6446 (N_6446,N_5552,N_5678);
and U6447 (N_6447,N_5547,N_5860);
or U6448 (N_6448,N_5530,N_5687);
nand U6449 (N_6449,N_5898,N_5642);
or U6450 (N_6450,N_5650,N_5857);
nand U6451 (N_6451,N_5848,N_5618);
and U6452 (N_6452,N_5550,N_5918);
nor U6453 (N_6453,N_5927,N_5627);
or U6454 (N_6454,N_5748,N_5703);
nand U6455 (N_6455,N_5810,N_5637);
nand U6456 (N_6456,N_5894,N_5954);
xor U6457 (N_6457,N_5787,N_5821);
xor U6458 (N_6458,N_5609,N_5886);
or U6459 (N_6459,N_5502,N_5864);
nand U6460 (N_6460,N_5671,N_5990);
nand U6461 (N_6461,N_5977,N_5659);
nand U6462 (N_6462,N_5790,N_5708);
or U6463 (N_6463,N_5603,N_5994);
nand U6464 (N_6464,N_5938,N_5948);
or U6465 (N_6465,N_5603,N_5833);
xnor U6466 (N_6466,N_5657,N_5610);
or U6467 (N_6467,N_5985,N_5536);
nor U6468 (N_6468,N_5828,N_5751);
xnor U6469 (N_6469,N_5574,N_5646);
and U6470 (N_6470,N_5607,N_5587);
and U6471 (N_6471,N_5802,N_5539);
or U6472 (N_6472,N_5664,N_5635);
and U6473 (N_6473,N_5644,N_5565);
and U6474 (N_6474,N_5705,N_5500);
or U6475 (N_6475,N_5604,N_5612);
or U6476 (N_6476,N_5708,N_5817);
and U6477 (N_6477,N_5566,N_5706);
nand U6478 (N_6478,N_5960,N_5642);
nor U6479 (N_6479,N_5839,N_5994);
nor U6480 (N_6480,N_5676,N_5594);
nand U6481 (N_6481,N_5720,N_5945);
or U6482 (N_6482,N_5570,N_5639);
or U6483 (N_6483,N_5767,N_5585);
or U6484 (N_6484,N_5944,N_5525);
or U6485 (N_6485,N_5593,N_5931);
xnor U6486 (N_6486,N_5935,N_5710);
nand U6487 (N_6487,N_5647,N_5655);
xor U6488 (N_6488,N_5966,N_5767);
or U6489 (N_6489,N_5902,N_5615);
nand U6490 (N_6490,N_5845,N_5880);
and U6491 (N_6491,N_5665,N_5892);
and U6492 (N_6492,N_5782,N_5650);
xor U6493 (N_6493,N_5584,N_5835);
nand U6494 (N_6494,N_5750,N_5505);
xor U6495 (N_6495,N_5978,N_5962);
nand U6496 (N_6496,N_5822,N_5656);
or U6497 (N_6497,N_5888,N_5741);
nand U6498 (N_6498,N_5646,N_5532);
xnor U6499 (N_6499,N_5516,N_5606);
nand U6500 (N_6500,N_6379,N_6078);
nand U6501 (N_6501,N_6465,N_6361);
nor U6502 (N_6502,N_6422,N_6087);
xor U6503 (N_6503,N_6265,N_6247);
nand U6504 (N_6504,N_6479,N_6016);
or U6505 (N_6505,N_6142,N_6056);
xnor U6506 (N_6506,N_6424,N_6272);
nor U6507 (N_6507,N_6374,N_6220);
nand U6508 (N_6508,N_6290,N_6381);
and U6509 (N_6509,N_6472,N_6298);
nand U6510 (N_6510,N_6029,N_6403);
xnor U6511 (N_6511,N_6080,N_6366);
and U6512 (N_6512,N_6450,N_6214);
nor U6513 (N_6513,N_6127,N_6475);
and U6514 (N_6514,N_6447,N_6279);
or U6515 (N_6515,N_6204,N_6227);
nor U6516 (N_6516,N_6481,N_6253);
and U6517 (N_6517,N_6449,N_6476);
and U6518 (N_6518,N_6362,N_6074);
nand U6519 (N_6519,N_6477,N_6024);
xor U6520 (N_6520,N_6002,N_6110);
and U6521 (N_6521,N_6445,N_6244);
xnor U6522 (N_6522,N_6027,N_6008);
or U6523 (N_6523,N_6275,N_6098);
xor U6524 (N_6524,N_6224,N_6116);
and U6525 (N_6525,N_6398,N_6178);
or U6526 (N_6526,N_6267,N_6208);
xor U6527 (N_6527,N_6269,N_6393);
and U6528 (N_6528,N_6073,N_6489);
and U6529 (N_6529,N_6287,N_6277);
and U6530 (N_6530,N_6294,N_6451);
xor U6531 (N_6531,N_6130,N_6286);
nand U6532 (N_6532,N_6363,N_6229);
nor U6533 (N_6533,N_6484,N_6312);
nor U6534 (N_6534,N_6210,N_6443);
xor U6535 (N_6535,N_6187,N_6421);
or U6536 (N_6536,N_6478,N_6232);
or U6537 (N_6537,N_6463,N_6076);
and U6538 (N_6538,N_6297,N_6365);
xnor U6539 (N_6539,N_6406,N_6175);
nor U6540 (N_6540,N_6164,N_6119);
and U6541 (N_6541,N_6207,N_6355);
xnor U6542 (N_6542,N_6216,N_6263);
or U6543 (N_6543,N_6123,N_6072);
or U6544 (N_6544,N_6011,N_6439);
xor U6545 (N_6545,N_6293,N_6097);
nor U6546 (N_6546,N_6154,N_6303);
nor U6547 (N_6547,N_6181,N_6332);
xnor U6548 (N_6548,N_6436,N_6360);
nor U6549 (N_6549,N_6033,N_6274);
nand U6550 (N_6550,N_6282,N_6161);
nor U6551 (N_6551,N_6452,N_6165);
and U6552 (N_6552,N_6377,N_6431);
and U6553 (N_6553,N_6050,N_6048);
nand U6554 (N_6554,N_6030,N_6409);
xor U6555 (N_6555,N_6068,N_6045);
xor U6556 (N_6556,N_6474,N_6041);
xnor U6557 (N_6557,N_6236,N_6213);
xnor U6558 (N_6558,N_6205,N_6042);
nand U6559 (N_6559,N_6032,N_6378);
and U6560 (N_6560,N_6411,N_6237);
or U6561 (N_6561,N_6020,N_6141);
xor U6562 (N_6562,N_6368,N_6299);
or U6563 (N_6563,N_6330,N_6083);
nor U6564 (N_6564,N_6261,N_6319);
nand U6565 (N_6565,N_6199,N_6099);
nand U6566 (N_6566,N_6367,N_6356);
or U6567 (N_6567,N_6334,N_6081);
nor U6568 (N_6568,N_6037,N_6348);
and U6569 (N_6569,N_6155,N_6483);
or U6570 (N_6570,N_6113,N_6462);
nand U6571 (N_6571,N_6103,N_6292);
and U6572 (N_6572,N_6322,N_6053);
nor U6573 (N_6573,N_6400,N_6309);
nand U6574 (N_6574,N_6318,N_6352);
and U6575 (N_6575,N_6316,N_6039);
nor U6576 (N_6576,N_6440,N_6225);
nand U6577 (N_6577,N_6469,N_6276);
xnor U6578 (N_6578,N_6211,N_6082);
nor U6579 (N_6579,N_6174,N_6306);
or U6580 (N_6580,N_6133,N_6243);
nand U6581 (N_6581,N_6414,N_6031);
nor U6582 (N_6582,N_6308,N_6285);
xor U6583 (N_6583,N_6284,N_6304);
xnor U6584 (N_6584,N_6240,N_6057);
nand U6585 (N_6585,N_6115,N_6486);
or U6586 (N_6586,N_6248,N_6004);
and U6587 (N_6587,N_6258,N_6091);
and U6588 (N_6588,N_6249,N_6109);
nand U6589 (N_6589,N_6129,N_6071);
or U6590 (N_6590,N_6467,N_6497);
and U6591 (N_6591,N_6254,N_6438);
nor U6592 (N_6592,N_6490,N_6149);
nand U6593 (N_6593,N_6327,N_6487);
and U6594 (N_6594,N_6172,N_6397);
xnor U6595 (N_6595,N_6245,N_6035);
or U6596 (N_6596,N_6280,N_6173);
xnor U6597 (N_6597,N_6320,N_6215);
or U6598 (N_6598,N_6460,N_6212);
or U6599 (N_6599,N_6353,N_6444);
nor U6600 (N_6600,N_6346,N_6455);
or U6601 (N_6601,N_6291,N_6435);
xor U6602 (N_6602,N_6264,N_6093);
nand U6603 (N_6603,N_6192,N_6184);
xnor U6604 (N_6604,N_6310,N_6364);
and U6605 (N_6605,N_6420,N_6022);
nor U6606 (N_6606,N_6335,N_6168);
nor U6607 (N_6607,N_6301,N_6122);
xnor U6608 (N_6608,N_6102,N_6454);
or U6609 (N_6609,N_6058,N_6195);
or U6610 (N_6610,N_6494,N_6009);
nand U6611 (N_6611,N_6038,N_6217);
and U6612 (N_6612,N_6437,N_6121);
nand U6613 (N_6613,N_6458,N_6186);
nand U6614 (N_6614,N_6166,N_6125);
nand U6615 (N_6615,N_6390,N_6021);
nor U6616 (N_6616,N_6104,N_6295);
xor U6617 (N_6617,N_6001,N_6108);
and U6618 (N_6618,N_6075,N_6158);
nand U6619 (N_6619,N_6111,N_6179);
nand U6620 (N_6620,N_6343,N_6090);
or U6621 (N_6621,N_6105,N_6006);
xnor U6622 (N_6622,N_6170,N_6466);
xor U6623 (N_6623,N_6473,N_6266);
or U6624 (N_6624,N_6413,N_6176);
or U6625 (N_6625,N_6140,N_6281);
or U6626 (N_6626,N_6014,N_6059);
xnor U6627 (N_6627,N_6350,N_6230);
xor U6628 (N_6628,N_6156,N_6325);
and U6629 (N_6629,N_6448,N_6496);
nor U6630 (N_6630,N_6391,N_6468);
and U6631 (N_6631,N_6339,N_6314);
nand U6632 (N_6632,N_6259,N_6470);
nand U6633 (N_6633,N_6415,N_6047);
or U6634 (N_6634,N_6197,N_6410);
and U6635 (N_6635,N_6376,N_6372);
and U6636 (N_6636,N_6333,N_6498);
nor U6637 (N_6637,N_6000,N_6499);
or U6638 (N_6638,N_6066,N_6340);
nor U6639 (N_6639,N_6412,N_6423);
nand U6640 (N_6640,N_6126,N_6321);
and U6641 (N_6641,N_6446,N_6416);
and U6642 (N_6642,N_6025,N_6338);
and U6643 (N_6643,N_6380,N_6384);
xor U6644 (N_6644,N_6271,N_6117);
nor U6645 (N_6645,N_6329,N_6369);
nand U6646 (N_6646,N_6182,N_6200);
nor U6647 (N_6647,N_6358,N_6088);
or U6648 (N_6648,N_6132,N_6302);
xor U6649 (N_6649,N_6150,N_6433);
or U6650 (N_6650,N_6069,N_6148);
nor U6651 (N_6651,N_6019,N_6387);
nor U6652 (N_6652,N_6417,N_6337);
nor U6653 (N_6653,N_6430,N_6112);
and U6654 (N_6654,N_6100,N_6300);
nor U6655 (N_6655,N_6062,N_6485);
or U6656 (N_6656,N_6235,N_6251);
or U6657 (N_6657,N_6015,N_6311);
xnor U6658 (N_6658,N_6060,N_6394);
nand U6659 (N_6659,N_6250,N_6101);
or U6660 (N_6660,N_6064,N_6492);
and U6661 (N_6661,N_6138,N_6392);
xor U6662 (N_6662,N_6396,N_6324);
xnor U6663 (N_6663,N_6370,N_6228);
nand U6664 (N_6664,N_6456,N_6052);
and U6665 (N_6665,N_6296,N_6453);
nor U6666 (N_6666,N_6395,N_6005);
xnor U6667 (N_6667,N_6180,N_6218);
xnor U6668 (N_6668,N_6043,N_6375);
and U6669 (N_6669,N_6077,N_6023);
nand U6670 (N_6670,N_6094,N_6386);
nor U6671 (N_6671,N_6070,N_6034);
or U6672 (N_6672,N_6151,N_6238);
nor U6673 (N_6673,N_6233,N_6190);
nand U6674 (N_6674,N_6252,N_6313);
nand U6675 (N_6675,N_6131,N_6345);
and U6676 (N_6676,N_6203,N_6188);
nor U6677 (N_6677,N_6134,N_6341);
and U6678 (N_6678,N_6418,N_6471);
nand U6679 (N_6679,N_6012,N_6089);
nand U6680 (N_6680,N_6044,N_6028);
nand U6681 (N_6681,N_6221,N_6429);
and U6682 (N_6682,N_6177,N_6139);
xor U6683 (N_6683,N_6336,N_6357);
nand U6684 (N_6684,N_6171,N_6241);
and U6685 (N_6685,N_6144,N_6488);
and U6686 (N_6686,N_6383,N_6326);
xor U6687 (N_6687,N_6007,N_6427);
xnor U6688 (N_6688,N_6079,N_6193);
xor U6689 (N_6689,N_6457,N_6136);
nor U6690 (N_6690,N_6096,N_6354);
xnor U6691 (N_6691,N_6226,N_6153);
or U6692 (N_6692,N_6242,N_6183);
xor U6693 (N_6693,N_6107,N_6389);
nor U6694 (N_6694,N_6349,N_6194);
and U6695 (N_6695,N_6273,N_6480);
xnor U6696 (N_6696,N_6323,N_6114);
and U6697 (N_6697,N_6347,N_6118);
nand U6698 (N_6698,N_6201,N_6189);
nand U6699 (N_6699,N_6160,N_6305);
xor U6700 (N_6700,N_6428,N_6441);
xor U6701 (N_6701,N_6373,N_6092);
nand U6702 (N_6702,N_6425,N_6185);
or U6703 (N_6703,N_6371,N_6426);
xnor U6704 (N_6704,N_6404,N_6464);
nor U6705 (N_6705,N_6268,N_6388);
nor U6706 (N_6706,N_6124,N_6106);
nand U6707 (N_6707,N_6482,N_6010);
xor U6708 (N_6708,N_6419,N_6159);
and U6709 (N_6709,N_6408,N_6491);
nand U6710 (N_6710,N_6169,N_6328);
xor U6711 (N_6711,N_6086,N_6036);
xor U6712 (N_6712,N_6442,N_6399);
nor U6713 (N_6713,N_6157,N_6026);
nand U6714 (N_6714,N_6401,N_6003);
xnor U6715 (N_6715,N_6065,N_6288);
and U6716 (N_6716,N_6342,N_6128);
nor U6717 (N_6717,N_6351,N_6493);
nor U6718 (N_6718,N_6051,N_6054);
or U6719 (N_6719,N_6206,N_6067);
or U6720 (N_6720,N_6063,N_6084);
or U6721 (N_6721,N_6163,N_6146);
nor U6722 (N_6722,N_6095,N_6120);
nor U6723 (N_6723,N_6198,N_6135);
nor U6724 (N_6724,N_6256,N_6018);
or U6725 (N_6725,N_6017,N_6143);
and U6726 (N_6726,N_6402,N_6331);
xor U6727 (N_6727,N_6385,N_6209);
and U6728 (N_6728,N_6495,N_6262);
nand U6729 (N_6729,N_6257,N_6145);
or U6730 (N_6730,N_6061,N_6152);
or U6731 (N_6731,N_6246,N_6270);
nor U6732 (N_6732,N_6307,N_6432);
and U6733 (N_6733,N_6255,N_6162);
nor U6734 (N_6734,N_6202,N_6239);
nor U6735 (N_6735,N_6167,N_6382);
or U6736 (N_6736,N_6137,N_6344);
nand U6737 (N_6737,N_6234,N_6461);
nand U6738 (N_6738,N_6085,N_6317);
nand U6739 (N_6739,N_6191,N_6283);
nand U6740 (N_6740,N_6219,N_6049);
nor U6741 (N_6741,N_6359,N_6315);
xor U6742 (N_6742,N_6459,N_6260);
xnor U6743 (N_6743,N_6013,N_6434);
and U6744 (N_6744,N_6046,N_6147);
xnor U6745 (N_6745,N_6231,N_6040);
or U6746 (N_6746,N_6222,N_6196);
or U6747 (N_6747,N_6278,N_6405);
and U6748 (N_6748,N_6055,N_6407);
and U6749 (N_6749,N_6289,N_6223);
nor U6750 (N_6750,N_6490,N_6276);
or U6751 (N_6751,N_6071,N_6476);
and U6752 (N_6752,N_6378,N_6180);
nor U6753 (N_6753,N_6471,N_6361);
nand U6754 (N_6754,N_6007,N_6313);
xnor U6755 (N_6755,N_6124,N_6099);
and U6756 (N_6756,N_6138,N_6266);
and U6757 (N_6757,N_6295,N_6428);
nand U6758 (N_6758,N_6311,N_6151);
or U6759 (N_6759,N_6359,N_6207);
or U6760 (N_6760,N_6361,N_6023);
nor U6761 (N_6761,N_6307,N_6380);
nor U6762 (N_6762,N_6156,N_6369);
and U6763 (N_6763,N_6453,N_6015);
xnor U6764 (N_6764,N_6208,N_6041);
and U6765 (N_6765,N_6399,N_6105);
nor U6766 (N_6766,N_6433,N_6107);
xor U6767 (N_6767,N_6135,N_6257);
nor U6768 (N_6768,N_6415,N_6222);
or U6769 (N_6769,N_6137,N_6301);
nor U6770 (N_6770,N_6352,N_6203);
and U6771 (N_6771,N_6132,N_6146);
and U6772 (N_6772,N_6437,N_6102);
nand U6773 (N_6773,N_6315,N_6392);
xor U6774 (N_6774,N_6056,N_6190);
nor U6775 (N_6775,N_6146,N_6456);
xnor U6776 (N_6776,N_6330,N_6137);
or U6777 (N_6777,N_6140,N_6313);
nand U6778 (N_6778,N_6002,N_6123);
nand U6779 (N_6779,N_6139,N_6468);
or U6780 (N_6780,N_6131,N_6202);
nand U6781 (N_6781,N_6477,N_6080);
or U6782 (N_6782,N_6112,N_6479);
xor U6783 (N_6783,N_6353,N_6010);
or U6784 (N_6784,N_6020,N_6302);
and U6785 (N_6785,N_6383,N_6054);
xnor U6786 (N_6786,N_6364,N_6311);
or U6787 (N_6787,N_6182,N_6082);
and U6788 (N_6788,N_6246,N_6394);
and U6789 (N_6789,N_6190,N_6037);
nand U6790 (N_6790,N_6252,N_6228);
nand U6791 (N_6791,N_6271,N_6324);
or U6792 (N_6792,N_6398,N_6066);
xnor U6793 (N_6793,N_6213,N_6074);
xnor U6794 (N_6794,N_6304,N_6372);
xor U6795 (N_6795,N_6497,N_6156);
and U6796 (N_6796,N_6069,N_6429);
or U6797 (N_6797,N_6107,N_6297);
or U6798 (N_6798,N_6259,N_6020);
nor U6799 (N_6799,N_6376,N_6082);
and U6800 (N_6800,N_6375,N_6054);
or U6801 (N_6801,N_6236,N_6298);
and U6802 (N_6802,N_6286,N_6157);
nand U6803 (N_6803,N_6374,N_6468);
and U6804 (N_6804,N_6494,N_6291);
xor U6805 (N_6805,N_6164,N_6266);
nand U6806 (N_6806,N_6293,N_6149);
nor U6807 (N_6807,N_6293,N_6228);
and U6808 (N_6808,N_6189,N_6006);
nor U6809 (N_6809,N_6379,N_6278);
nor U6810 (N_6810,N_6364,N_6191);
or U6811 (N_6811,N_6398,N_6457);
or U6812 (N_6812,N_6087,N_6213);
or U6813 (N_6813,N_6035,N_6039);
xor U6814 (N_6814,N_6318,N_6116);
nor U6815 (N_6815,N_6168,N_6155);
xor U6816 (N_6816,N_6062,N_6227);
xnor U6817 (N_6817,N_6128,N_6260);
nand U6818 (N_6818,N_6201,N_6407);
or U6819 (N_6819,N_6036,N_6004);
nor U6820 (N_6820,N_6368,N_6373);
xnor U6821 (N_6821,N_6457,N_6307);
or U6822 (N_6822,N_6049,N_6157);
xor U6823 (N_6823,N_6431,N_6135);
and U6824 (N_6824,N_6354,N_6338);
nand U6825 (N_6825,N_6108,N_6180);
and U6826 (N_6826,N_6464,N_6311);
xnor U6827 (N_6827,N_6211,N_6170);
xor U6828 (N_6828,N_6271,N_6367);
nand U6829 (N_6829,N_6309,N_6159);
xor U6830 (N_6830,N_6395,N_6382);
or U6831 (N_6831,N_6137,N_6480);
and U6832 (N_6832,N_6295,N_6024);
xnor U6833 (N_6833,N_6046,N_6159);
and U6834 (N_6834,N_6460,N_6191);
xor U6835 (N_6835,N_6448,N_6416);
nor U6836 (N_6836,N_6058,N_6094);
xor U6837 (N_6837,N_6279,N_6087);
nand U6838 (N_6838,N_6365,N_6192);
nor U6839 (N_6839,N_6098,N_6410);
and U6840 (N_6840,N_6195,N_6261);
or U6841 (N_6841,N_6184,N_6127);
xnor U6842 (N_6842,N_6060,N_6284);
nor U6843 (N_6843,N_6062,N_6114);
or U6844 (N_6844,N_6244,N_6472);
and U6845 (N_6845,N_6366,N_6496);
nand U6846 (N_6846,N_6313,N_6083);
nor U6847 (N_6847,N_6036,N_6226);
and U6848 (N_6848,N_6070,N_6279);
nor U6849 (N_6849,N_6110,N_6127);
and U6850 (N_6850,N_6100,N_6367);
and U6851 (N_6851,N_6495,N_6145);
or U6852 (N_6852,N_6422,N_6283);
or U6853 (N_6853,N_6210,N_6252);
or U6854 (N_6854,N_6298,N_6141);
nand U6855 (N_6855,N_6486,N_6244);
xor U6856 (N_6856,N_6018,N_6281);
nor U6857 (N_6857,N_6374,N_6044);
nand U6858 (N_6858,N_6365,N_6002);
nand U6859 (N_6859,N_6132,N_6303);
or U6860 (N_6860,N_6100,N_6093);
and U6861 (N_6861,N_6120,N_6264);
or U6862 (N_6862,N_6242,N_6085);
nand U6863 (N_6863,N_6399,N_6393);
xor U6864 (N_6864,N_6183,N_6140);
xnor U6865 (N_6865,N_6281,N_6309);
nor U6866 (N_6866,N_6082,N_6067);
nand U6867 (N_6867,N_6009,N_6190);
or U6868 (N_6868,N_6094,N_6295);
nor U6869 (N_6869,N_6069,N_6153);
nand U6870 (N_6870,N_6490,N_6476);
and U6871 (N_6871,N_6224,N_6422);
xnor U6872 (N_6872,N_6434,N_6485);
or U6873 (N_6873,N_6041,N_6062);
or U6874 (N_6874,N_6473,N_6414);
and U6875 (N_6875,N_6164,N_6246);
nand U6876 (N_6876,N_6372,N_6189);
nor U6877 (N_6877,N_6324,N_6220);
nand U6878 (N_6878,N_6435,N_6070);
nor U6879 (N_6879,N_6160,N_6269);
or U6880 (N_6880,N_6310,N_6122);
nor U6881 (N_6881,N_6227,N_6460);
xor U6882 (N_6882,N_6443,N_6208);
xnor U6883 (N_6883,N_6096,N_6278);
and U6884 (N_6884,N_6355,N_6120);
nand U6885 (N_6885,N_6249,N_6157);
and U6886 (N_6886,N_6104,N_6316);
and U6887 (N_6887,N_6078,N_6003);
nor U6888 (N_6888,N_6155,N_6360);
nand U6889 (N_6889,N_6206,N_6282);
or U6890 (N_6890,N_6417,N_6071);
and U6891 (N_6891,N_6005,N_6025);
nor U6892 (N_6892,N_6095,N_6241);
or U6893 (N_6893,N_6163,N_6330);
xor U6894 (N_6894,N_6193,N_6097);
and U6895 (N_6895,N_6143,N_6207);
and U6896 (N_6896,N_6409,N_6182);
xor U6897 (N_6897,N_6251,N_6231);
nand U6898 (N_6898,N_6090,N_6492);
nand U6899 (N_6899,N_6333,N_6347);
nor U6900 (N_6900,N_6249,N_6313);
nor U6901 (N_6901,N_6305,N_6193);
nand U6902 (N_6902,N_6156,N_6183);
nor U6903 (N_6903,N_6424,N_6076);
nor U6904 (N_6904,N_6457,N_6293);
and U6905 (N_6905,N_6105,N_6205);
nor U6906 (N_6906,N_6447,N_6222);
nor U6907 (N_6907,N_6341,N_6425);
nor U6908 (N_6908,N_6017,N_6467);
or U6909 (N_6909,N_6036,N_6414);
nand U6910 (N_6910,N_6263,N_6096);
nand U6911 (N_6911,N_6493,N_6162);
nor U6912 (N_6912,N_6059,N_6211);
xor U6913 (N_6913,N_6241,N_6164);
nor U6914 (N_6914,N_6483,N_6128);
xnor U6915 (N_6915,N_6045,N_6443);
and U6916 (N_6916,N_6067,N_6498);
nor U6917 (N_6917,N_6346,N_6088);
nand U6918 (N_6918,N_6180,N_6300);
xor U6919 (N_6919,N_6171,N_6085);
xnor U6920 (N_6920,N_6485,N_6035);
and U6921 (N_6921,N_6139,N_6251);
nand U6922 (N_6922,N_6435,N_6489);
and U6923 (N_6923,N_6059,N_6222);
and U6924 (N_6924,N_6063,N_6427);
and U6925 (N_6925,N_6309,N_6165);
nor U6926 (N_6926,N_6207,N_6441);
and U6927 (N_6927,N_6448,N_6145);
nor U6928 (N_6928,N_6121,N_6057);
and U6929 (N_6929,N_6247,N_6340);
nand U6930 (N_6930,N_6265,N_6156);
and U6931 (N_6931,N_6499,N_6186);
or U6932 (N_6932,N_6172,N_6231);
xnor U6933 (N_6933,N_6183,N_6419);
nor U6934 (N_6934,N_6416,N_6419);
nand U6935 (N_6935,N_6392,N_6130);
and U6936 (N_6936,N_6220,N_6227);
nand U6937 (N_6937,N_6005,N_6403);
or U6938 (N_6938,N_6286,N_6046);
xor U6939 (N_6939,N_6452,N_6473);
xor U6940 (N_6940,N_6173,N_6428);
nand U6941 (N_6941,N_6378,N_6043);
or U6942 (N_6942,N_6271,N_6001);
nor U6943 (N_6943,N_6234,N_6191);
xnor U6944 (N_6944,N_6242,N_6114);
or U6945 (N_6945,N_6203,N_6489);
xor U6946 (N_6946,N_6134,N_6160);
and U6947 (N_6947,N_6396,N_6117);
nor U6948 (N_6948,N_6198,N_6304);
nor U6949 (N_6949,N_6161,N_6053);
and U6950 (N_6950,N_6293,N_6172);
and U6951 (N_6951,N_6160,N_6466);
nand U6952 (N_6952,N_6257,N_6495);
and U6953 (N_6953,N_6200,N_6244);
nor U6954 (N_6954,N_6280,N_6463);
or U6955 (N_6955,N_6295,N_6320);
or U6956 (N_6956,N_6037,N_6018);
nor U6957 (N_6957,N_6006,N_6344);
or U6958 (N_6958,N_6281,N_6278);
xor U6959 (N_6959,N_6083,N_6414);
xnor U6960 (N_6960,N_6336,N_6401);
nand U6961 (N_6961,N_6371,N_6443);
xor U6962 (N_6962,N_6095,N_6463);
and U6963 (N_6963,N_6136,N_6113);
xnor U6964 (N_6964,N_6499,N_6308);
xnor U6965 (N_6965,N_6287,N_6022);
or U6966 (N_6966,N_6200,N_6483);
nand U6967 (N_6967,N_6050,N_6172);
nand U6968 (N_6968,N_6179,N_6158);
and U6969 (N_6969,N_6151,N_6477);
nand U6970 (N_6970,N_6216,N_6056);
or U6971 (N_6971,N_6148,N_6300);
nand U6972 (N_6972,N_6002,N_6178);
nor U6973 (N_6973,N_6252,N_6032);
xnor U6974 (N_6974,N_6137,N_6133);
or U6975 (N_6975,N_6305,N_6128);
xnor U6976 (N_6976,N_6008,N_6310);
nand U6977 (N_6977,N_6095,N_6268);
or U6978 (N_6978,N_6492,N_6216);
nor U6979 (N_6979,N_6003,N_6273);
and U6980 (N_6980,N_6279,N_6477);
xor U6981 (N_6981,N_6251,N_6344);
xnor U6982 (N_6982,N_6384,N_6030);
and U6983 (N_6983,N_6096,N_6470);
xnor U6984 (N_6984,N_6272,N_6303);
xor U6985 (N_6985,N_6141,N_6093);
xnor U6986 (N_6986,N_6118,N_6248);
nand U6987 (N_6987,N_6263,N_6302);
xor U6988 (N_6988,N_6015,N_6255);
or U6989 (N_6989,N_6000,N_6436);
nor U6990 (N_6990,N_6443,N_6160);
or U6991 (N_6991,N_6450,N_6050);
or U6992 (N_6992,N_6408,N_6136);
nor U6993 (N_6993,N_6113,N_6109);
and U6994 (N_6994,N_6268,N_6214);
or U6995 (N_6995,N_6035,N_6094);
nor U6996 (N_6996,N_6014,N_6020);
or U6997 (N_6997,N_6347,N_6368);
and U6998 (N_6998,N_6269,N_6364);
and U6999 (N_6999,N_6319,N_6313);
nand U7000 (N_7000,N_6873,N_6565);
nand U7001 (N_7001,N_6673,N_6876);
xnor U7002 (N_7002,N_6974,N_6536);
and U7003 (N_7003,N_6702,N_6560);
nor U7004 (N_7004,N_6802,N_6645);
nand U7005 (N_7005,N_6507,N_6526);
and U7006 (N_7006,N_6892,N_6927);
nor U7007 (N_7007,N_6527,N_6879);
nand U7008 (N_7008,N_6520,N_6674);
or U7009 (N_7009,N_6906,N_6680);
nor U7010 (N_7010,N_6602,N_6523);
and U7011 (N_7011,N_6577,N_6812);
xnor U7012 (N_7012,N_6706,N_6994);
nand U7013 (N_7013,N_6529,N_6938);
nor U7014 (N_7014,N_6593,N_6775);
xor U7015 (N_7015,N_6984,N_6584);
nand U7016 (N_7016,N_6754,N_6929);
nor U7017 (N_7017,N_6948,N_6514);
nor U7018 (N_7018,N_6612,N_6937);
nor U7019 (N_7019,N_6830,N_6962);
or U7020 (N_7020,N_6646,N_6557);
nor U7021 (N_7021,N_6890,N_6945);
and U7022 (N_7022,N_6715,N_6666);
and U7023 (N_7023,N_6925,N_6651);
nand U7024 (N_7024,N_6505,N_6548);
or U7025 (N_7025,N_6883,N_6722);
or U7026 (N_7026,N_6664,N_6820);
and U7027 (N_7027,N_6899,N_6778);
nor U7028 (N_7028,N_6961,N_6955);
xor U7029 (N_7029,N_6840,N_6877);
nand U7030 (N_7030,N_6744,N_6695);
nor U7031 (N_7031,N_6796,N_6518);
and U7032 (N_7032,N_6894,N_6941);
nand U7033 (N_7033,N_6575,N_6758);
xnor U7034 (N_7034,N_6530,N_6832);
xnor U7035 (N_7035,N_6632,N_6697);
and U7036 (N_7036,N_6630,N_6528);
nand U7037 (N_7037,N_6968,N_6886);
or U7038 (N_7038,N_6772,N_6782);
nand U7039 (N_7039,N_6777,N_6599);
nor U7040 (N_7040,N_6547,N_6689);
and U7041 (N_7041,N_6932,N_6639);
or U7042 (N_7042,N_6606,N_6851);
nand U7043 (N_7043,N_6717,N_6719);
xor U7044 (N_7044,N_6977,N_6848);
or U7045 (N_7045,N_6972,N_6787);
nand U7046 (N_7046,N_6956,N_6742);
nand U7047 (N_7047,N_6978,N_6862);
nand U7048 (N_7048,N_6784,N_6506);
and U7049 (N_7049,N_6764,N_6912);
nor U7050 (N_7050,N_6953,N_6756);
xnor U7051 (N_7051,N_6677,N_6916);
nor U7052 (N_7052,N_6844,N_6985);
or U7053 (N_7053,N_6939,N_6700);
and U7054 (N_7054,N_6740,N_6684);
nand U7055 (N_7055,N_6752,N_6556);
and U7056 (N_7056,N_6672,N_6736);
and U7057 (N_7057,N_6753,N_6853);
nand U7058 (N_7058,N_6838,N_6720);
and U7059 (N_7059,N_6751,N_6936);
xnor U7060 (N_7060,N_6662,N_6635);
nor U7061 (N_7061,N_6611,N_6931);
nor U7062 (N_7062,N_6683,N_6889);
nor U7063 (N_7063,N_6551,N_6538);
xor U7064 (N_7064,N_6767,N_6667);
xnor U7065 (N_7065,N_6696,N_6976);
xor U7066 (N_7066,N_6549,N_6841);
or U7067 (N_7067,N_6813,N_6852);
nand U7068 (N_7068,N_6582,N_6511);
or U7069 (N_7069,N_6607,N_6998);
or U7070 (N_7070,N_6516,N_6587);
and U7071 (N_7071,N_6738,N_6896);
nor U7072 (N_7072,N_6571,N_6641);
nand U7073 (N_7073,N_6746,N_6703);
xnor U7074 (N_7074,N_6681,N_6731);
nand U7075 (N_7075,N_6735,N_6712);
nand U7076 (N_7076,N_6979,N_6901);
xor U7077 (N_7077,N_6816,N_6687);
nand U7078 (N_7078,N_6629,N_6966);
nand U7079 (N_7079,N_6967,N_6934);
xnor U7080 (N_7080,N_6589,N_6855);
xor U7081 (N_7081,N_6888,N_6847);
xnor U7082 (N_7082,N_6915,N_6884);
and U7083 (N_7083,N_6874,N_6686);
or U7084 (N_7084,N_6709,N_6918);
and U7085 (N_7085,N_6519,N_6643);
nor U7086 (N_7086,N_6842,N_6950);
nor U7087 (N_7087,N_6621,N_6585);
nor U7088 (N_7088,N_6729,N_6613);
and U7089 (N_7089,N_6597,N_6710);
nand U7090 (N_7090,N_6903,N_6546);
xor U7091 (N_7091,N_6980,N_6574);
and U7092 (N_7092,N_6502,N_6581);
xnor U7093 (N_7093,N_6623,N_6598);
or U7094 (N_7094,N_6821,N_6963);
or U7095 (N_7095,N_6657,N_6943);
and U7096 (N_7096,N_6576,N_6570);
nor U7097 (N_7097,N_6940,N_6922);
and U7098 (N_7098,N_6871,N_6914);
and U7099 (N_7099,N_6792,N_6648);
nor U7100 (N_7100,N_6745,N_6615);
nor U7101 (N_7101,N_6776,N_6590);
or U7102 (N_7102,N_6803,N_6951);
or U7103 (N_7103,N_6552,N_6804);
and U7104 (N_7104,N_6724,N_6878);
nor U7105 (N_7105,N_6992,N_6504);
nand U7106 (N_7106,N_6875,N_6647);
xor U7107 (N_7107,N_6555,N_6983);
nand U7108 (N_7108,N_6671,N_6868);
or U7109 (N_7109,N_6670,N_6592);
xnor U7110 (N_7110,N_6627,N_6701);
or U7111 (N_7111,N_6898,N_6793);
xor U7112 (N_7112,N_6935,N_6869);
nand U7113 (N_7113,N_6824,N_6655);
and U7114 (N_7114,N_6870,N_6788);
or U7115 (N_7115,N_6762,N_6624);
nor U7116 (N_7116,N_6827,N_6653);
and U7117 (N_7117,N_6917,N_6880);
and U7118 (N_7118,N_6679,N_6781);
nand U7119 (N_7119,N_6760,N_6825);
or U7120 (N_7120,N_6763,N_6975);
xor U7121 (N_7121,N_6849,N_6521);
or U7122 (N_7122,N_6944,N_6801);
and U7123 (N_7123,N_6583,N_6734);
and U7124 (N_7124,N_6791,N_6866);
and U7125 (N_7125,N_6969,N_6900);
nor U7126 (N_7126,N_6790,N_6616);
or U7127 (N_7127,N_6532,N_6881);
nand U7128 (N_7128,N_6947,N_6522);
and U7129 (N_7129,N_6910,N_6996);
nor U7130 (N_7130,N_6640,N_6805);
nand U7131 (N_7131,N_6800,N_6794);
nand U7132 (N_7132,N_6911,N_6885);
and U7133 (N_7133,N_6887,N_6893);
xnor U7134 (N_7134,N_6661,N_6858);
xor U7135 (N_7135,N_6609,N_6748);
nor U7136 (N_7136,N_6924,N_6721);
xor U7137 (N_7137,N_6601,N_6688);
and U7138 (N_7138,N_6786,N_6524);
nand U7139 (N_7139,N_6535,N_6770);
or U7140 (N_7140,N_6861,N_6542);
or U7141 (N_7141,N_6743,N_6831);
or U7142 (N_7142,N_6988,N_6822);
nand U7143 (N_7143,N_6867,N_6652);
or U7144 (N_7144,N_6676,N_6559);
nor U7145 (N_7145,N_6923,N_6649);
xnor U7146 (N_7146,N_6780,N_6895);
or U7147 (N_7147,N_6995,N_6891);
and U7148 (N_7148,N_6755,N_6540);
or U7149 (N_7149,N_6628,N_6926);
or U7150 (N_7150,N_6897,N_6904);
or U7151 (N_7151,N_6865,N_6818);
xnor U7152 (N_7152,N_6919,N_6579);
and U7153 (N_7153,N_6508,N_6839);
nor U7154 (N_7154,N_6588,N_6964);
nor U7155 (N_7155,N_6779,N_6603);
nor U7156 (N_7156,N_6991,N_6586);
or U7157 (N_7157,N_6930,N_6659);
and U7158 (N_7158,N_6625,N_6563);
nand U7159 (N_7159,N_6795,N_6958);
or U7160 (N_7160,N_6739,N_6699);
nand U7161 (N_7161,N_6642,N_6704);
nor U7162 (N_7162,N_6741,N_6761);
nand U7163 (N_7163,N_6531,N_6626);
or U7164 (N_7164,N_6810,N_6726);
and U7165 (N_7165,N_6733,N_6614);
nor U7166 (N_7166,N_6675,N_6633);
or U7167 (N_7167,N_6631,N_6959);
and U7168 (N_7168,N_6872,N_6971);
or U7169 (N_7169,N_6845,N_6716);
and U7170 (N_7170,N_6909,N_6834);
nand U7171 (N_7171,N_6814,N_6771);
or U7172 (N_7172,N_6545,N_6863);
and U7173 (N_7173,N_6638,N_6989);
xnor U7174 (N_7174,N_6533,N_6510);
nor U7175 (N_7175,N_6564,N_6750);
and U7176 (N_7176,N_6694,N_6990);
nand U7177 (N_7177,N_6713,N_6622);
xor U7178 (N_7178,N_6833,N_6567);
xor U7179 (N_7179,N_6634,N_6512);
nand U7180 (N_7180,N_6554,N_6905);
nor U7181 (N_7181,N_6882,N_6658);
nand U7182 (N_7182,N_6856,N_6809);
nor U7183 (N_7183,N_6660,N_6811);
and U7184 (N_7184,N_6707,N_6501);
nor U7185 (N_7185,N_6591,N_6569);
and U7186 (N_7186,N_6543,N_6798);
xnor U7187 (N_7187,N_6580,N_6541);
or U7188 (N_7188,N_6749,N_6544);
xnor U7189 (N_7189,N_6783,N_6942);
and U7190 (N_7190,N_6690,N_6509);
nor U7191 (N_7191,N_6768,N_6513);
or U7192 (N_7192,N_6920,N_6558);
nand U7193 (N_7193,N_6807,N_6728);
nor U7194 (N_7194,N_6785,N_6952);
nor U7195 (N_7195,N_6596,N_6553);
nor U7196 (N_7196,N_6859,N_6600);
nor U7197 (N_7197,N_6561,N_6836);
or U7198 (N_7198,N_6823,N_6981);
and U7199 (N_7199,N_6973,N_6685);
nor U7200 (N_7200,N_6620,N_6997);
or U7201 (N_7201,N_6503,N_6757);
nand U7202 (N_7202,N_6765,N_6682);
nor U7203 (N_7203,N_6698,N_6797);
nor U7204 (N_7204,N_6982,N_6747);
nand U7205 (N_7205,N_6846,N_6921);
xor U7206 (N_7206,N_6789,N_6986);
xor U7207 (N_7207,N_6730,N_6668);
nor U7208 (N_7208,N_6714,N_6573);
and U7209 (N_7209,N_6525,N_6817);
or U7210 (N_7210,N_6578,N_6644);
or U7211 (N_7211,N_6737,N_6769);
or U7212 (N_7212,N_6678,N_6534);
nor U7213 (N_7213,N_6949,N_6605);
xnor U7214 (N_7214,N_6725,N_6957);
or U7215 (N_7215,N_6669,N_6993);
nor U7216 (N_7216,N_6808,N_6608);
or U7217 (N_7217,N_6727,N_6960);
xnor U7218 (N_7218,N_6568,N_6954);
and U7219 (N_7219,N_6732,N_6850);
xor U7220 (N_7220,N_6595,N_6718);
xor U7221 (N_7221,N_6773,N_6843);
or U7222 (N_7222,N_6946,N_6618);
and U7223 (N_7223,N_6774,N_6860);
and U7224 (N_7224,N_6650,N_6799);
nor U7225 (N_7225,N_6654,N_6636);
nor U7226 (N_7226,N_6766,N_6705);
and U7227 (N_7227,N_6908,N_6835);
nor U7228 (N_7228,N_6987,N_6902);
and U7229 (N_7229,N_6965,N_6663);
nand U7230 (N_7230,N_6515,N_6759);
or U7231 (N_7231,N_6610,N_6815);
nor U7232 (N_7232,N_6864,N_6691);
and U7233 (N_7233,N_6819,N_6933);
or U7234 (N_7234,N_6806,N_6913);
xnor U7235 (N_7235,N_6537,N_6828);
and U7236 (N_7236,N_6692,N_6999);
nor U7237 (N_7237,N_6837,N_6619);
and U7238 (N_7238,N_6826,N_6711);
xnor U7239 (N_7239,N_6566,N_6604);
xnor U7240 (N_7240,N_6500,N_6637);
nand U7241 (N_7241,N_6550,N_6928);
or U7242 (N_7242,N_6907,N_6708);
nand U7243 (N_7243,N_6617,N_6572);
xor U7244 (N_7244,N_6562,N_6665);
xnor U7245 (N_7245,N_6829,N_6594);
and U7246 (N_7246,N_6656,N_6854);
or U7247 (N_7247,N_6693,N_6723);
nand U7248 (N_7248,N_6517,N_6970);
nor U7249 (N_7249,N_6539,N_6857);
nor U7250 (N_7250,N_6670,N_6958);
nor U7251 (N_7251,N_6596,N_6749);
or U7252 (N_7252,N_6698,N_6770);
xor U7253 (N_7253,N_6525,N_6621);
nand U7254 (N_7254,N_6624,N_6746);
and U7255 (N_7255,N_6528,N_6612);
and U7256 (N_7256,N_6774,N_6743);
nand U7257 (N_7257,N_6628,N_6752);
and U7258 (N_7258,N_6713,N_6935);
xnor U7259 (N_7259,N_6531,N_6671);
nor U7260 (N_7260,N_6948,N_6672);
nor U7261 (N_7261,N_6620,N_6931);
nand U7262 (N_7262,N_6564,N_6908);
nand U7263 (N_7263,N_6589,N_6659);
nand U7264 (N_7264,N_6506,N_6668);
xor U7265 (N_7265,N_6899,N_6971);
nand U7266 (N_7266,N_6946,N_6662);
and U7267 (N_7267,N_6843,N_6660);
nor U7268 (N_7268,N_6702,N_6535);
and U7269 (N_7269,N_6654,N_6598);
nand U7270 (N_7270,N_6777,N_6713);
nor U7271 (N_7271,N_6814,N_6808);
xor U7272 (N_7272,N_6680,N_6951);
nand U7273 (N_7273,N_6740,N_6777);
nor U7274 (N_7274,N_6607,N_6619);
or U7275 (N_7275,N_6549,N_6877);
or U7276 (N_7276,N_6875,N_6951);
nor U7277 (N_7277,N_6770,N_6784);
xnor U7278 (N_7278,N_6627,N_6948);
or U7279 (N_7279,N_6738,N_6787);
xor U7280 (N_7280,N_6639,N_6621);
xnor U7281 (N_7281,N_6792,N_6856);
xor U7282 (N_7282,N_6836,N_6544);
and U7283 (N_7283,N_6819,N_6839);
nor U7284 (N_7284,N_6875,N_6510);
xnor U7285 (N_7285,N_6607,N_6601);
nor U7286 (N_7286,N_6979,N_6814);
xor U7287 (N_7287,N_6802,N_6641);
xor U7288 (N_7288,N_6660,N_6775);
nand U7289 (N_7289,N_6845,N_6898);
nor U7290 (N_7290,N_6661,N_6849);
xor U7291 (N_7291,N_6928,N_6722);
or U7292 (N_7292,N_6599,N_6768);
nand U7293 (N_7293,N_6596,N_6607);
nor U7294 (N_7294,N_6508,N_6588);
nor U7295 (N_7295,N_6729,N_6942);
nand U7296 (N_7296,N_6708,N_6733);
and U7297 (N_7297,N_6741,N_6722);
xor U7298 (N_7298,N_6783,N_6633);
or U7299 (N_7299,N_6961,N_6569);
xnor U7300 (N_7300,N_6938,N_6619);
and U7301 (N_7301,N_6884,N_6710);
and U7302 (N_7302,N_6992,N_6829);
xor U7303 (N_7303,N_6512,N_6530);
and U7304 (N_7304,N_6711,N_6976);
xor U7305 (N_7305,N_6614,N_6670);
nand U7306 (N_7306,N_6955,N_6971);
nand U7307 (N_7307,N_6625,N_6662);
or U7308 (N_7308,N_6547,N_6842);
and U7309 (N_7309,N_6637,N_6791);
nand U7310 (N_7310,N_6583,N_6960);
xnor U7311 (N_7311,N_6892,N_6878);
or U7312 (N_7312,N_6917,N_6876);
or U7313 (N_7313,N_6618,N_6769);
nand U7314 (N_7314,N_6957,N_6601);
nor U7315 (N_7315,N_6714,N_6547);
and U7316 (N_7316,N_6919,N_6877);
nor U7317 (N_7317,N_6570,N_6849);
xnor U7318 (N_7318,N_6801,N_6608);
and U7319 (N_7319,N_6583,N_6853);
nor U7320 (N_7320,N_6751,N_6815);
or U7321 (N_7321,N_6678,N_6721);
or U7322 (N_7322,N_6701,N_6575);
and U7323 (N_7323,N_6920,N_6918);
xor U7324 (N_7324,N_6946,N_6747);
and U7325 (N_7325,N_6781,N_6892);
nand U7326 (N_7326,N_6957,N_6781);
and U7327 (N_7327,N_6659,N_6729);
xnor U7328 (N_7328,N_6937,N_6751);
or U7329 (N_7329,N_6737,N_6690);
or U7330 (N_7330,N_6623,N_6676);
xor U7331 (N_7331,N_6828,N_6506);
nand U7332 (N_7332,N_6659,N_6513);
or U7333 (N_7333,N_6667,N_6848);
nand U7334 (N_7334,N_6985,N_6628);
nand U7335 (N_7335,N_6647,N_6587);
xnor U7336 (N_7336,N_6741,N_6980);
nor U7337 (N_7337,N_6648,N_6864);
nor U7338 (N_7338,N_6811,N_6940);
and U7339 (N_7339,N_6507,N_6983);
or U7340 (N_7340,N_6533,N_6761);
xnor U7341 (N_7341,N_6699,N_6629);
nand U7342 (N_7342,N_6931,N_6662);
xnor U7343 (N_7343,N_6731,N_6758);
nand U7344 (N_7344,N_6930,N_6687);
xnor U7345 (N_7345,N_6938,N_6859);
nand U7346 (N_7346,N_6644,N_6608);
nand U7347 (N_7347,N_6500,N_6906);
xnor U7348 (N_7348,N_6596,N_6921);
xnor U7349 (N_7349,N_6841,N_6716);
or U7350 (N_7350,N_6746,N_6676);
nor U7351 (N_7351,N_6620,N_6659);
xnor U7352 (N_7352,N_6886,N_6712);
or U7353 (N_7353,N_6865,N_6728);
and U7354 (N_7354,N_6773,N_6651);
xnor U7355 (N_7355,N_6748,N_6962);
or U7356 (N_7356,N_6708,N_6521);
nor U7357 (N_7357,N_6787,N_6587);
or U7358 (N_7358,N_6627,N_6513);
nor U7359 (N_7359,N_6788,N_6560);
and U7360 (N_7360,N_6657,N_6836);
xor U7361 (N_7361,N_6836,N_6923);
and U7362 (N_7362,N_6884,N_6797);
xor U7363 (N_7363,N_6770,N_6685);
and U7364 (N_7364,N_6875,N_6919);
or U7365 (N_7365,N_6536,N_6706);
or U7366 (N_7366,N_6561,N_6559);
nand U7367 (N_7367,N_6756,N_6712);
and U7368 (N_7368,N_6981,N_6784);
nor U7369 (N_7369,N_6609,N_6749);
nand U7370 (N_7370,N_6763,N_6890);
nor U7371 (N_7371,N_6912,N_6854);
nor U7372 (N_7372,N_6871,N_6595);
nor U7373 (N_7373,N_6513,N_6617);
nand U7374 (N_7374,N_6788,N_6707);
nand U7375 (N_7375,N_6924,N_6830);
or U7376 (N_7376,N_6503,N_6849);
nor U7377 (N_7377,N_6931,N_6618);
nand U7378 (N_7378,N_6772,N_6672);
nor U7379 (N_7379,N_6940,N_6818);
or U7380 (N_7380,N_6517,N_6679);
and U7381 (N_7381,N_6529,N_6894);
and U7382 (N_7382,N_6895,N_6734);
and U7383 (N_7383,N_6758,N_6680);
or U7384 (N_7384,N_6798,N_6810);
nand U7385 (N_7385,N_6576,N_6535);
nor U7386 (N_7386,N_6908,N_6561);
nor U7387 (N_7387,N_6780,N_6658);
nand U7388 (N_7388,N_6910,N_6877);
nor U7389 (N_7389,N_6660,N_6886);
nor U7390 (N_7390,N_6733,N_6660);
xnor U7391 (N_7391,N_6830,N_6874);
nor U7392 (N_7392,N_6655,N_6643);
or U7393 (N_7393,N_6710,N_6880);
or U7394 (N_7394,N_6626,N_6534);
nand U7395 (N_7395,N_6924,N_6828);
nand U7396 (N_7396,N_6578,N_6739);
xor U7397 (N_7397,N_6534,N_6828);
nor U7398 (N_7398,N_6519,N_6849);
xnor U7399 (N_7399,N_6854,N_6865);
and U7400 (N_7400,N_6561,N_6767);
xnor U7401 (N_7401,N_6792,N_6826);
nor U7402 (N_7402,N_6803,N_6932);
nand U7403 (N_7403,N_6989,N_6828);
nand U7404 (N_7404,N_6768,N_6719);
or U7405 (N_7405,N_6907,N_6825);
or U7406 (N_7406,N_6929,N_6926);
or U7407 (N_7407,N_6982,N_6921);
and U7408 (N_7408,N_6885,N_6993);
or U7409 (N_7409,N_6597,N_6976);
nand U7410 (N_7410,N_6601,N_6961);
nand U7411 (N_7411,N_6503,N_6536);
xnor U7412 (N_7412,N_6586,N_6530);
and U7413 (N_7413,N_6849,N_6985);
and U7414 (N_7414,N_6657,N_6894);
and U7415 (N_7415,N_6619,N_6760);
nand U7416 (N_7416,N_6516,N_6672);
and U7417 (N_7417,N_6535,N_6941);
nand U7418 (N_7418,N_6839,N_6718);
nor U7419 (N_7419,N_6573,N_6877);
or U7420 (N_7420,N_6710,N_6767);
xnor U7421 (N_7421,N_6988,N_6672);
or U7422 (N_7422,N_6802,N_6932);
or U7423 (N_7423,N_6846,N_6510);
nor U7424 (N_7424,N_6622,N_6815);
and U7425 (N_7425,N_6678,N_6538);
nand U7426 (N_7426,N_6849,N_6828);
nor U7427 (N_7427,N_6713,N_6726);
nor U7428 (N_7428,N_6556,N_6529);
and U7429 (N_7429,N_6791,N_6690);
or U7430 (N_7430,N_6945,N_6787);
and U7431 (N_7431,N_6933,N_6964);
xnor U7432 (N_7432,N_6671,N_6706);
nor U7433 (N_7433,N_6803,N_6677);
xor U7434 (N_7434,N_6519,N_6755);
or U7435 (N_7435,N_6811,N_6625);
and U7436 (N_7436,N_6911,N_6693);
or U7437 (N_7437,N_6500,N_6892);
or U7438 (N_7438,N_6977,N_6546);
or U7439 (N_7439,N_6548,N_6656);
and U7440 (N_7440,N_6679,N_6547);
or U7441 (N_7441,N_6923,N_6944);
and U7442 (N_7442,N_6999,N_6661);
nand U7443 (N_7443,N_6548,N_6919);
and U7444 (N_7444,N_6723,N_6596);
xnor U7445 (N_7445,N_6642,N_6606);
xor U7446 (N_7446,N_6878,N_6564);
nand U7447 (N_7447,N_6739,N_6796);
and U7448 (N_7448,N_6660,N_6556);
nand U7449 (N_7449,N_6863,N_6985);
or U7450 (N_7450,N_6779,N_6777);
or U7451 (N_7451,N_6550,N_6824);
and U7452 (N_7452,N_6796,N_6928);
xor U7453 (N_7453,N_6589,N_6766);
nor U7454 (N_7454,N_6864,N_6724);
and U7455 (N_7455,N_6604,N_6606);
nor U7456 (N_7456,N_6916,N_6761);
xor U7457 (N_7457,N_6902,N_6759);
and U7458 (N_7458,N_6895,N_6837);
xnor U7459 (N_7459,N_6690,N_6868);
xor U7460 (N_7460,N_6835,N_6870);
xor U7461 (N_7461,N_6929,N_6724);
and U7462 (N_7462,N_6630,N_6653);
xor U7463 (N_7463,N_6594,N_6658);
and U7464 (N_7464,N_6967,N_6850);
xnor U7465 (N_7465,N_6724,N_6676);
nand U7466 (N_7466,N_6789,N_6998);
and U7467 (N_7467,N_6650,N_6626);
and U7468 (N_7468,N_6682,N_6743);
or U7469 (N_7469,N_6918,N_6525);
nor U7470 (N_7470,N_6873,N_6542);
and U7471 (N_7471,N_6889,N_6839);
and U7472 (N_7472,N_6513,N_6975);
and U7473 (N_7473,N_6543,N_6995);
and U7474 (N_7474,N_6858,N_6682);
nand U7475 (N_7475,N_6740,N_6548);
nor U7476 (N_7476,N_6598,N_6642);
xnor U7477 (N_7477,N_6577,N_6533);
nor U7478 (N_7478,N_6588,N_6568);
or U7479 (N_7479,N_6979,N_6953);
nand U7480 (N_7480,N_6849,N_6668);
nor U7481 (N_7481,N_6801,N_6500);
or U7482 (N_7482,N_6992,N_6679);
or U7483 (N_7483,N_6581,N_6631);
nand U7484 (N_7484,N_6564,N_6865);
nor U7485 (N_7485,N_6770,N_6558);
and U7486 (N_7486,N_6854,N_6908);
or U7487 (N_7487,N_6886,N_6961);
nand U7488 (N_7488,N_6647,N_6511);
nor U7489 (N_7489,N_6519,N_6640);
and U7490 (N_7490,N_6981,N_6588);
nor U7491 (N_7491,N_6911,N_6692);
nand U7492 (N_7492,N_6812,N_6996);
or U7493 (N_7493,N_6880,N_6599);
nor U7494 (N_7494,N_6554,N_6547);
nor U7495 (N_7495,N_6602,N_6597);
nand U7496 (N_7496,N_6540,N_6589);
or U7497 (N_7497,N_6958,N_6842);
xnor U7498 (N_7498,N_6750,N_6519);
nand U7499 (N_7499,N_6611,N_6890);
xor U7500 (N_7500,N_7433,N_7006);
xor U7501 (N_7501,N_7298,N_7209);
and U7502 (N_7502,N_7243,N_7383);
and U7503 (N_7503,N_7220,N_7049);
xnor U7504 (N_7504,N_7344,N_7125);
nor U7505 (N_7505,N_7030,N_7240);
and U7506 (N_7506,N_7069,N_7406);
and U7507 (N_7507,N_7495,N_7258);
and U7508 (N_7508,N_7200,N_7428);
nand U7509 (N_7509,N_7287,N_7124);
and U7510 (N_7510,N_7087,N_7466);
nor U7511 (N_7511,N_7073,N_7392);
nor U7512 (N_7512,N_7063,N_7436);
nor U7513 (N_7513,N_7247,N_7452);
xnor U7514 (N_7514,N_7170,N_7234);
xnor U7515 (N_7515,N_7017,N_7145);
xor U7516 (N_7516,N_7133,N_7486);
or U7517 (N_7517,N_7116,N_7393);
nor U7518 (N_7518,N_7369,N_7283);
or U7519 (N_7519,N_7147,N_7329);
xnor U7520 (N_7520,N_7489,N_7016);
or U7521 (N_7521,N_7110,N_7041);
and U7522 (N_7522,N_7427,N_7152);
nor U7523 (N_7523,N_7107,N_7195);
nand U7524 (N_7524,N_7260,N_7176);
nand U7525 (N_7525,N_7191,N_7192);
or U7526 (N_7526,N_7231,N_7096);
or U7527 (N_7527,N_7174,N_7168);
nor U7528 (N_7528,N_7481,N_7440);
nand U7529 (N_7529,N_7375,N_7022);
and U7530 (N_7530,N_7336,N_7280);
and U7531 (N_7531,N_7018,N_7417);
nand U7532 (N_7532,N_7267,N_7345);
nand U7533 (N_7533,N_7294,N_7015);
nor U7534 (N_7534,N_7108,N_7216);
xnor U7535 (N_7535,N_7215,N_7488);
or U7536 (N_7536,N_7480,N_7071);
nor U7537 (N_7537,N_7162,N_7288);
or U7538 (N_7538,N_7461,N_7212);
nor U7539 (N_7539,N_7270,N_7410);
or U7540 (N_7540,N_7400,N_7444);
xor U7541 (N_7541,N_7164,N_7402);
xor U7542 (N_7542,N_7142,N_7084);
or U7543 (N_7543,N_7448,N_7307);
or U7544 (N_7544,N_7381,N_7050);
xor U7545 (N_7545,N_7246,N_7103);
and U7546 (N_7546,N_7225,N_7420);
and U7547 (N_7547,N_7470,N_7059);
xor U7548 (N_7548,N_7151,N_7169);
nor U7549 (N_7549,N_7377,N_7439);
nand U7550 (N_7550,N_7154,N_7370);
and U7551 (N_7551,N_7180,N_7324);
and U7552 (N_7552,N_7476,N_7187);
and U7553 (N_7553,N_7379,N_7237);
nor U7554 (N_7554,N_7399,N_7353);
xnor U7555 (N_7555,N_7356,N_7218);
and U7556 (N_7556,N_7214,N_7358);
nand U7557 (N_7557,N_7348,N_7323);
or U7558 (N_7558,N_7019,N_7135);
or U7559 (N_7559,N_7366,N_7424);
or U7560 (N_7560,N_7198,N_7227);
and U7561 (N_7561,N_7331,N_7000);
and U7562 (N_7562,N_7100,N_7499);
or U7563 (N_7563,N_7357,N_7408);
or U7564 (N_7564,N_7469,N_7349);
nor U7565 (N_7565,N_7091,N_7411);
or U7566 (N_7566,N_7241,N_7458);
nand U7567 (N_7567,N_7045,N_7001);
xnor U7568 (N_7568,N_7484,N_7075);
and U7569 (N_7569,N_7184,N_7447);
or U7570 (N_7570,N_7313,N_7360);
nor U7571 (N_7571,N_7141,N_7423);
and U7572 (N_7572,N_7095,N_7014);
xnor U7573 (N_7573,N_7304,N_7264);
xor U7574 (N_7574,N_7013,N_7396);
nor U7575 (N_7575,N_7414,N_7046);
xor U7576 (N_7576,N_7204,N_7009);
nand U7577 (N_7577,N_7099,N_7032);
xor U7578 (N_7578,N_7378,N_7438);
xnor U7579 (N_7579,N_7111,N_7020);
and U7580 (N_7580,N_7354,N_7351);
and U7581 (N_7581,N_7306,N_7315);
and U7582 (N_7582,N_7232,N_7121);
xnor U7583 (N_7583,N_7413,N_7337);
nor U7584 (N_7584,N_7387,N_7181);
nand U7585 (N_7585,N_7449,N_7493);
nor U7586 (N_7586,N_7285,N_7021);
nand U7587 (N_7587,N_7043,N_7418);
or U7588 (N_7588,N_7295,N_7165);
or U7589 (N_7589,N_7189,N_7425);
nand U7590 (N_7590,N_7202,N_7211);
nand U7591 (N_7591,N_7056,N_7185);
nand U7592 (N_7592,N_7465,N_7302);
nand U7593 (N_7593,N_7037,N_7085);
or U7594 (N_7594,N_7341,N_7002);
and U7595 (N_7595,N_7036,N_7093);
nand U7596 (N_7596,N_7109,N_7359);
nand U7597 (N_7597,N_7042,N_7311);
nor U7598 (N_7598,N_7308,N_7397);
nand U7599 (N_7599,N_7299,N_7060);
nand U7600 (N_7600,N_7117,N_7248);
or U7601 (N_7601,N_7319,N_7072);
nand U7602 (N_7602,N_7389,N_7317);
and U7603 (N_7603,N_7228,N_7415);
nor U7604 (N_7604,N_7419,N_7496);
and U7605 (N_7605,N_7441,N_7213);
nand U7606 (N_7606,N_7177,N_7094);
nor U7607 (N_7607,N_7450,N_7179);
or U7608 (N_7608,N_7482,N_7089);
and U7609 (N_7609,N_7472,N_7498);
or U7610 (N_7610,N_7146,N_7004);
xor U7611 (N_7611,N_7158,N_7340);
nand U7612 (N_7612,N_7123,N_7404);
or U7613 (N_7613,N_7274,N_7321);
or U7614 (N_7614,N_7455,N_7265);
nand U7615 (N_7615,N_7376,N_7318);
nand U7616 (N_7616,N_7055,N_7077);
or U7617 (N_7617,N_7062,N_7303);
or U7618 (N_7618,N_7497,N_7080);
or U7619 (N_7619,N_7430,N_7088);
nor U7620 (N_7620,N_7083,N_7028);
and U7621 (N_7621,N_7188,N_7309);
nor U7622 (N_7622,N_7473,N_7058);
or U7623 (N_7623,N_7183,N_7252);
or U7624 (N_7624,N_7244,N_7391);
and U7625 (N_7625,N_7273,N_7171);
and U7626 (N_7626,N_7401,N_7143);
and U7627 (N_7627,N_7190,N_7076);
nor U7628 (N_7628,N_7118,N_7445);
nand U7629 (N_7629,N_7325,N_7460);
nand U7630 (N_7630,N_7047,N_7459);
and U7631 (N_7631,N_7233,N_7160);
and U7632 (N_7632,N_7350,N_7372);
or U7633 (N_7633,N_7039,N_7464);
nor U7634 (N_7634,N_7422,N_7483);
or U7635 (N_7635,N_7194,N_7024);
xor U7636 (N_7636,N_7296,N_7398);
or U7637 (N_7637,N_7205,N_7355);
or U7638 (N_7638,N_7167,N_7451);
and U7639 (N_7639,N_7412,N_7173);
nor U7640 (N_7640,N_7082,N_7196);
nand U7641 (N_7641,N_7338,N_7035);
nand U7642 (N_7642,N_7012,N_7380);
nand U7643 (N_7643,N_7003,N_7395);
xnor U7644 (N_7644,N_7286,N_7104);
nand U7645 (N_7645,N_7025,N_7256);
nor U7646 (N_7646,N_7182,N_7262);
xor U7647 (N_7647,N_7407,N_7051);
or U7648 (N_7648,N_7301,N_7106);
and U7649 (N_7649,N_7334,N_7268);
and U7650 (N_7650,N_7253,N_7092);
xnor U7651 (N_7651,N_7312,N_7266);
xnor U7652 (N_7652,N_7224,N_7197);
and U7653 (N_7653,N_7305,N_7153);
nand U7654 (N_7654,N_7250,N_7186);
and U7655 (N_7655,N_7219,N_7172);
nor U7656 (N_7656,N_7081,N_7409);
xor U7657 (N_7657,N_7175,N_7065);
nand U7658 (N_7658,N_7367,N_7127);
nand U7659 (N_7659,N_7434,N_7097);
nand U7660 (N_7660,N_7139,N_7442);
and U7661 (N_7661,N_7166,N_7029);
xor U7662 (N_7662,N_7475,N_7140);
or U7663 (N_7663,N_7269,N_7238);
xor U7664 (N_7664,N_7326,N_7487);
nand U7665 (N_7665,N_7226,N_7038);
nor U7666 (N_7666,N_7272,N_7163);
xor U7667 (N_7667,N_7136,N_7291);
nand U7668 (N_7668,N_7388,N_7245);
and U7669 (N_7669,N_7208,N_7207);
and U7670 (N_7670,N_7462,N_7382);
nand U7671 (N_7671,N_7130,N_7115);
nand U7672 (N_7672,N_7333,N_7474);
or U7673 (N_7673,N_7132,N_7054);
or U7674 (N_7674,N_7282,N_7254);
or U7675 (N_7675,N_7101,N_7284);
nor U7676 (N_7676,N_7330,N_7279);
nand U7677 (N_7677,N_7027,N_7031);
nand U7678 (N_7678,N_7431,N_7206);
or U7679 (N_7679,N_7229,N_7098);
nand U7680 (N_7680,N_7048,N_7068);
or U7681 (N_7681,N_7339,N_7131);
or U7682 (N_7682,N_7119,N_7421);
or U7683 (N_7683,N_7390,N_7137);
nand U7684 (N_7684,N_7230,N_7102);
or U7685 (N_7685,N_7454,N_7492);
nor U7686 (N_7686,N_7271,N_7010);
or U7687 (N_7687,N_7007,N_7343);
nand U7688 (N_7688,N_7485,N_7149);
nor U7689 (N_7689,N_7426,N_7086);
and U7690 (N_7690,N_7249,N_7079);
and U7691 (N_7691,N_7067,N_7005);
and U7692 (N_7692,N_7314,N_7052);
nand U7693 (N_7693,N_7126,N_7134);
nand U7694 (N_7694,N_7394,N_7105);
nor U7695 (N_7695,N_7471,N_7144);
xnor U7696 (N_7696,N_7361,N_7332);
xnor U7697 (N_7697,N_7453,N_7263);
or U7698 (N_7698,N_7386,N_7429);
or U7699 (N_7699,N_7373,N_7368);
xnor U7700 (N_7700,N_7011,N_7328);
xor U7701 (N_7701,N_7148,N_7385);
and U7702 (N_7702,N_7457,N_7316);
nor U7703 (N_7703,N_7026,N_7278);
nor U7704 (N_7704,N_7159,N_7310);
and U7705 (N_7705,N_7289,N_7384);
xnor U7706 (N_7706,N_7074,N_7157);
and U7707 (N_7707,N_7405,N_7352);
nor U7708 (N_7708,N_7479,N_7199);
and U7709 (N_7709,N_7374,N_7090);
or U7710 (N_7710,N_7365,N_7128);
or U7711 (N_7711,N_7033,N_7178);
or U7712 (N_7712,N_7362,N_7057);
nand U7713 (N_7713,N_7477,N_7120);
nor U7714 (N_7714,N_7346,N_7297);
and U7715 (N_7715,N_7223,N_7203);
nand U7716 (N_7716,N_7320,N_7201);
or U7717 (N_7717,N_7078,N_7138);
or U7718 (N_7718,N_7255,N_7403);
nand U7719 (N_7719,N_7277,N_7478);
nor U7720 (N_7720,N_7463,N_7161);
xor U7721 (N_7721,N_7235,N_7034);
nor U7722 (N_7722,N_7112,N_7491);
and U7723 (N_7723,N_7150,N_7221);
xor U7724 (N_7724,N_7114,N_7040);
xor U7725 (N_7725,N_7281,N_7432);
xor U7726 (N_7726,N_7193,N_7217);
or U7727 (N_7727,N_7064,N_7456);
nand U7728 (N_7728,N_7276,N_7293);
and U7729 (N_7729,N_7044,N_7053);
or U7730 (N_7730,N_7061,N_7008);
and U7731 (N_7731,N_7300,N_7468);
nor U7732 (N_7732,N_7261,N_7210);
nand U7733 (N_7733,N_7239,N_7467);
or U7734 (N_7734,N_7259,N_7122);
or U7735 (N_7735,N_7364,N_7070);
nand U7736 (N_7736,N_7494,N_7416);
and U7737 (N_7737,N_7342,N_7066);
nand U7738 (N_7738,N_7129,N_7371);
and U7739 (N_7739,N_7322,N_7236);
or U7740 (N_7740,N_7335,N_7446);
or U7741 (N_7741,N_7327,N_7257);
nor U7742 (N_7742,N_7437,N_7251);
or U7743 (N_7743,N_7156,N_7242);
nor U7744 (N_7744,N_7222,N_7290);
nor U7745 (N_7745,N_7113,N_7023);
xnor U7746 (N_7746,N_7155,N_7347);
nor U7747 (N_7747,N_7443,N_7363);
and U7748 (N_7748,N_7490,N_7292);
and U7749 (N_7749,N_7435,N_7275);
or U7750 (N_7750,N_7143,N_7445);
nand U7751 (N_7751,N_7472,N_7254);
or U7752 (N_7752,N_7409,N_7176);
or U7753 (N_7753,N_7080,N_7039);
nor U7754 (N_7754,N_7234,N_7422);
nor U7755 (N_7755,N_7173,N_7358);
xnor U7756 (N_7756,N_7455,N_7219);
nor U7757 (N_7757,N_7487,N_7312);
and U7758 (N_7758,N_7433,N_7067);
nand U7759 (N_7759,N_7304,N_7388);
xor U7760 (N_7760,N_7367,N_7350);
and U7761 (N_7761,N_7278,N_7172);
or U7762 (N_7762,N_7047,N_7413);
nand U7763 (N_7763,N_7067,N_7297);
xnor U7764 (N_7764,N_7156,N_7085);
or U7765 (N_7765,N_7232,N_7448);
or U7766 (N_7766,N_7367,N_7218);
xnor U7767 (N_7767,N_7051,N_7164);
or U7768 (N_7768,N_7107,N_7209);
nand U7769 (N_7769,N_7240,N_7119);
xor U7770 (N_7770,N_7274,N_7256);
xnor U7771 (N_7771,N_7250,N_7351);
nand U7772 (N_7772,N_7046,N_7495);
and U7773 (N_7773,N_7474,N_7133);
nor U7774 (N_7774,N_7318,N_7167);
xor U7775 (N_7775,N_7484,N_7205);
or U7776 (N_7776,N_7235,N_7167);
or U7777 (N_7777,N_7260,N_7131);
xnor U7778 (N_7778,N_7008,N_7126);
or U7779 (N_7779,N_7263,N_7305);
or U7780 (N_7780,N_7267,N_7107);
nor U7781 (N_7781,N_7009,N_7422);
nor U7782 (N_7782,N_7498,N_7054);
xnor U7783 (N_7783,N_7286,N_7435);
nand U7784 (N_7784,N_7301,N_7340);
nor U7785 (N_7785,N_7145,N_7369);
or U7786 (N_7786,N_7457,N_7247);
nor U7787 (N_7787,N_7470,N_7370);
nor U7788 (N_7788,N_7378,N_7009);
and U7789 (N_7789,N_7164,N_7421);
and U7790 (N_7790,N_7315,N_7435);
nor U7791 (N_7791,N_7333,N_7465);
or U7792 (N_7792,N_7034,N_7133);
nor U7793 (N_7793,N_7390,N_7066);
nand U7794 (N_7794,N_7262,N_7066);
or U7795 (N_7795,N_7202,N_7027);
nand U7796 (N_7796,N_7488,N_7217);
or U7797 (N_7797,N_7011,N_7068);
or U7798 (N_7798,N_7382,N_7262);
and U7799 (N_7799,N_7108,N_7177);
nand U7800 (N_7800,N_7477,N_7003);
and U7801 (N_7801,N_7104,N_7486);
nand U7802 (N_7802,N_7133,N_7416);
and U7803 (N_7803,N_7152,N_7360);
nor U7804 (N_7804,N_7377,N_7042);
nor U7805 (N_7805,N_7274,N_7114);
and U7806 (N_7806,N_7149,N_7026);
xor U7807 (N_7807,N_7427,N_7173);
xor U7808 (N_7808,N_7062,N_7256);
xnor U7809 (N_7809,N_7097,N_7453);
or U7810 (N_7810,N_7129,N_7488);
and U7811 (N_7811,N_7011,N_7444);
and U7812 (N_7812,N_7352,N_7013);
nand U7813 (N_7813,N_7477,N_7065);
and U7814 (N_7814,N_7310,N_7442);
or U7815 (N_7815,N_7341,N_7263);
xnor U7816 (N_7816,N_7029,N_7188);
and U7817 (N_7817,N_7377,N_7167);
nor U7818 (N_7818,N_7055,N_7084);
or U7819 (N_7819,N_7094,N_7034);
xnor U7820 (N_7820,N_7185,N_7374);
and U7821 (N_7821,N_7450,N_7044);
and U7822 (N_7822,N_7321,N_7326);
nor U7823 (N_7823,N_7247,N_7001);
nand U7824 (N_7824,N_7295,N_7152);
xor U7825 (N_7825,N_7419,N_7377);
nand U7826 (N_7826,N_7242,N_7132);
and U7827 (N_7827,N_7371,N_7162);
or U7828 (N_7828,N_7235,N_7482);
nor U7829 (N_7829,N_7482,N_7210);
and U7830 (N_7830,N_7395,N_7176);
nand U7831 (N_7831,N_7365,N_7429);
and U7832 (N_7832,N_7072,N_7430);
and U7833 (N_7833,N_7051,N_7389);
nand U7834 (N_7834,N_7405,N_7481);
nor U7835 (N_7835,N_7306,N_7362);
xor U7836 (N_7836,N_7433,N_7264);
and U7837 (N_7837,N_7339,N_7332);
nor U7838 (N_7838,N_7440,N_7405);
nor U7839 (N_7839,N_7449,N_7201);
or U7840 (N_7840,N_7146,N_7131);
nor U7841 (N_7841,N_7024,N_7076);
nand U7842 (N_7842,N_7401,N_7135);
xor U7843 (N_7843,N_7114,N_7392);
nand U7844 (N_7844,N_7059,N_7188);
and U7845 (N_7845,N_7396,N_7070);
and U7846 (N_7846,N_7345,N_7201);
nand U7847 (N_7847,N_7433,N_7200);
and U7848 (N_7848,N_7393,N_7323);
or U7849 (N_7849,N_7311,N_7227);
nand U7850 (N_7850,N_7438,N_7236);
or U7851 (N_7851,N_7223,N_7222);
and U7852 (N_7852,N_7450,N_7444);
xnor U7853 (N_7853,N_7114,N_7353);
or U7854 (N_7854,N_7175,N_7461);
xnor U7855 (N_7855,N_7156,N_7213);
nor U7856 (N_7856,N_7336,N_7436);
nor U7857 (N_7857,N_7364,N_7441);
nor U7858 (N_7858,N_7191,N_7264);
nor U7859 (N_7859,N_7465,N_7382);
and U7860 (N_7860,N_7146,N_7180);
and U7861 (N_7861,N_7061,N_7257);
xor U7862 (N_7862,N_7032,N_7001);
nand U7863 (N_7863,N_7415,N_7456);
nor U7864 (N_7864,N_7317,N_7471);
nor U7865 (N_7865,N_7270,N_7082);
or U7866 (N_7866,N_7199,N_7029);
or U7867 (N_7867,N_7121,N_7117);
nand U7868 (N_7868,N_7152,N_7084);
xor U7869 (N_7869,N_7172,N_7122);
or U7870 (N_7870,N_7475,N_7261);
xnor U7871 (N_7871,N_7388,N_7167);
and U7872 (N_7872,N_7180,N_7177);
and U7873 (N_7873,N_7032,N_7479);
nor U7874 (N_7874,N_7099,N_7154);
nand U7875 (N_7875,N_7249,N_7125);
and U7876 (N_7876,N_7247,N_7238);
nand U7877 (N_7877,N_7134,N_7240);
or U7878 (N_7878,N_7341,N_7056);
nand U7879 (N_7879,N_7478,N_7261);
nand U7880 (N_7880,N_7437,N_7014);
xnor U7881 (N_7881,N_7095,N_7083);
or U7882 (N_7882,N_7198,N_7431);
and U7883 (N_7883,N_7363,N_7453);
nor U7884 (N_7884,N_7282,N_7416);
nor U7885 (N_7885,N_7428,N_7481);
or U7886 (N_7886,N_7475,N_7217);
and U7887 (N_7887,N_7445,N_7479);
or U7888 (N_7888,N_7051,N_7453);
and U7889 (N_7889,N_7110,N_7379);
xnor U7890 (N_7890,N_7475,N_7081);
xnor U7891 (N_7891,N_7113,N_7394);
xor U7892 (N_7892,N_7311,N_7202);
xnor U7893 (N_7893,N_7275,N_7048);
and U7894 (N_7894,N_7276,N_7349);
and U7895 (N_7895,N_7056,N_7451);
nand U7896 (N_7896,N_7274,N_7039);
and U7897 (N_7897,N_7375,N_7251);
nor U7898 (N_7898,N_7364,N_7428);
and U7899 (N_7899,N_7136,N_7253);
and U7900 (N_7900,N_7263,N_7016);
nor U7901 (N_7901,N_7355,N_7235);
or U7902 (N_7902,N_7385,N_7153);
and U7903 (N_7903,N_7280,N_7106);
nor U7904 (N_7904,N_7279,N_7164);
xor U7905 (N_7905,N_7360,N_7107);
nand U7906 (N_7906,N_7217,N_7167);
and U7907 (N_7907,N_7043,N_7321);
and U7908 (N_7908,N_7019,N_7129);
or U7909 (N_7909,N_7069,N_7465);
nor U7910 (N_7910,N_7039,N_7277);
xnor U7911 (N_7911,N_7126,N_7268);
and U7912 (N_7912,N_7281,N_7385);
xnor U7913 (N_7913,N_7051,N_7264);
and U7914 (N_7914,N_7427,N_7185);
or U7915 (N_7915,N_7484,N_7083);
nand U7916 (N_7916,N_7315,N_7324);
or U7917 (N_7917,N_7217,N_7470);
xnor U7918 (N_7918,N_7421,N_7494);
or U7919 (N_7919,N_7058,N_7086);
or U7920 (N_7920,N_7032,N_7179);
nand U7921 (N_7921,N_7118,N_7483);
and U7922 (N_7922,N_7385,N_7127);
xnor U7923 (N_7923,N_7492,N_7451);
and U7924 (N_7924,N_7129,N_7411);
and U7925 (N_7925,N_7435,N_7100);
nand U7926 (N_7926,N_7293,N_7399);
and U7927 (N_7927,N_7317,N_7324);
nand U7928 (N_7928,N_7017,N_7104);
or U7929 (N_7929,N_7064,N_7329);
nand U7930 (N_7930,N_7342,N_7029);
or U7931 (N_7931,N_7115,N_7126);
or U7932 (N_7932,N_7462,N_7203);
nand U7933 (N_7933,N_7238,N_7121);
xnor U7934 (N_7934,N_7327,N_7275);
nand U7935 (N_7935,N_7455,N_7185);
nor U7936 (N_7936,N_7399,N_7078);
xor U7937 (N_7937,N_7448,N_7057);
nand U7938 (N_7938,N_7343,N_7164);
or U7939 (N_7939,N_7094,N_7159);
and U7940 (N_7940,N_7031,N_7133);
xnor U7941 (N_7941,N_7091,N_7447);
and U7942 (N_7942,N_7132,N_7076);
nor U7943 (N_7943,N_7417,N_7160);
and U7944 (N_7944,N_7020,N_7323);
or U7945 (N_7945,N_7131,N_7465);
nor U7946 (N_7946,N_7209,N_7181);
nand U7947 (N_7947,N_7393,N_7268);
nor U7948 (N_7948,N_7197,N_7249);
nand U7949 (N_7949,N_7295,N_7147);
nand U7950 (N_7950,N_7119,N_7408);
or U7951 (N_7951,N_7368,N_7179);
or U7952 (N_7952,N_7182,N_7406);
nand U7953 (N_7953,N_7205,N_7361);
xor U7954 (N_7954,N_7302,N_7206);
nand U7955 (N_7955,N_7398,N_7285);
nor U7956 (N_7956,N_7439,N_7029);
or U7957 (N_7957,N_7170,N_7492);
xnor U7958 (N_7958,N_7304,N_7119);
xnor U7959 (N_7959,N_7134,N_7330);
nor U7960 (N_7960,N_7452,N_7362);
or U7961 (N_7961,N_7161,N_7346);
nand U7962 (N_7962,N_7246,N_7199);
or U7963 (N_7963,N_7065,N_7291);
nor U7964 (N_7964,N_7234,N_7374);
nand U7965 (N_7965,N_7058,N_7135);
xor U7966 (N_7966,N_7162,N_7390);
nor U7967 (N_7967,N_7009,N_7235);
or U7968 (N_7968,N_7177,N_7319);
nor U7969 (N_7969,N_7220,N_7118);
nand U7970 (N_7970,N_7240,N_7300);
or U7971 (N_7971,N_7381,N_7079);
and U7972 (N_7972,N_7190,N_7288);
and U7973 (N_7973,N_7421,N_7162);
xor U7974 (N_7974,N_7013,N_7343);
nand U7975 (N_7975,N_7103,N_7387);
or U7976 (N_7976,N_7138,N_7266);
or U7977 (N_7977,N_7455,N_7477);
xnor U7978 (N_7978,N_7124,N_7435);
and U7979 (N_7979,N_7420,N_7448);
xor U7980 (N_7980,N_7429,N_7497);
nor U7981 (N_7981,N_7330,N_7206);
and U7982 (N_7982,N_7166,N_7066);
or U7983 (N_7983,N_7488,N_7164);
and U7984 (N_7984,N_7291,N_7472);
or U7985 (N_7985,N_7086,N_7456);
or U7986 (N_7986,N_7493,N_7307);
and U7987 (N_7987,N_7491,N_7362);
or U7988 (N_7988,N_7219,N_7352);
and U7989 (N_7989,N_7262,N_7268);
xor U7990 (N_7990,N_7408,N_7064);
and U7991 (N_7991,N_7437,N_7284);
xnor U7992 (N_7992,N_7012,N_7090);
or U7993 (N_7993,N_7452,N_7116);
xnor U7994 (N_7994,N_7202,N_7251);
and U7995 (N_7995,N_7224,N_7302);
and U7996 (N_7996,N_7170,N_7194);
xnor U7997 (N_7997,N_7134,N_7002);
nor U7998 (N_7998,N_7367,N_7426);
nor U7999 (N_7999,N_7057,N_7381);
nand U8000 (N_8000,N_7729,N_7685);
or U8001 (N_8001,N_7642,N_7573);
nor U8002 (N_8002,N_7779,N_7548);
nand U8003 (N_8003,N_7993,N_7668);
nand U8004 (N_8004,N_7813,N_7751);
nor U8005 (N_8005,N_7737,N_7741);
xnor U8006 (N_8006,N_7513,N_7827);
nand U8007 (N_8007,N_7522,N_7671);
nand U8008 (N_8008,N_7625,N_7539);
or U8009 (N_8009,N_7780,N_7787);
nand U8010 (N_8010,N_7790,N_7773);
or U8011 (N_8011,N_7555,N_7979);
nor U8012 (N_8012,N_7772,N_7783);
nor U8013 (N_8013,N_7726,N_7932);
and U8014 (N_8014,N_7564,N_7686);
xnor U8015 (N_8015,N_7621,N_7643);
and U8016 (N_8016,N_7805,N_7849);
nand U8017 (N_8017,N_7961,N_7927);
nand U8018 (N_8018,N_7609,N_7535);
nand U8019 (N_8019,N_7945,N_7518);
xor U8020 (N_8020,N_7524,N_7923);
xnor U8021 (N_8021,N_7906,N_7763);
or U8022 (N_8022,N_7968,N_7848);
and U8023 (N_8023,N_7701,N_7692);
and U8024 (N_8024,N_7965,N_7577);
nand U8025 (N_8025,N_7782,N_7630);
and U8026 (N_8026,N_7786,N_7820);
and U8027 (N_8027,N_7917,N_7620);
xnor U8028 (N_8028,N_7959,N_7706);
nand U8029 (N_8029,N_7595,N_7750);
or U8030 (N_8030,N_7559,N_7528);
or U8031 (N_8031,N_7985,N_7584);
nor U8032 (N_8032,N_7930,N_7908);
or U8033 (N_8033,N_7947,N_7624);
nand U8034 (N_8034,N_7694,N_7594);
or U8035 (N_8035,N_7900,N_7590);
nor U8036 (N_8036,N_7865,N_7626);
xnor U8037 (N_8037,N_7898,N_7834);
and U8038 (N_8038,N_7884,N_7822);
xnor U8039 (N_8039,N_7869,N_7596);
nor U8040 (N_8040,N_7514,N_7851);
nor U8041 (N_8041,N_7558,N_7759);
or U8042 (N_8042,N_7943,N_7975);
nor U8043 (N_8043,N_7736,N_7669);
or U8044 (N_8044,N_7617,N_7619);
or U8045 (N_8045,N_7637,N_7845);
nand U8046 (N_8046,N_7714,N_7536);
and U8047 (N_8047,N_7856,N_7921);
nor U8048 (N_8048,N_7659,N_7939);
nor U8049 (N_8049,N_7846,N_7891);
nor U8050 (N_8050,N_7651,N_7854);
nor U8051 (N_8051,N_7622,N_7838);
and U8052 (N_8052,N_7833,N_7720);
xnor U8053 (N_8053,N_7678,N_7852);
or U8054 (N_8054,N_7660,N_7814);
nand U8055 (N_8055,N_7537,N_7552);
nor U8056 (N_8056,N_7735,N_7871);
or U8057 (N_8057,N_7875,N_7591);
and U8058 (N_8058,N_7995,N_7699);
or U8059 (N_8059,N_7665,N_7661);
nor U8060 (N_8060,N_7918,N_7676);
nor U8061 (N_8061,N_7646,N_7738);
or U8062 (N_8062,N_7655,N_7821);
xor U8063 (N_8063,N_7769,N_7843);
nor U8064 (N_8064,N_7672,N_7935);
nor U8065 (N_8065,N_7842,N_7853);
nor U8066 (N_8066,N_7907,N_7929);
or U8067 (N_8067,N_7886,N_7996);
nor U8068 (N_8068,N_7964,N_7811);
or U8069 (N_8069,N_7766,N_7952);
nor U8070 (N_8070,N_7915,N_7713);
or U8071 (N_8071,N_7809,N_7687);
xnor U8072 (N_8072,N_7519,N_7926);
xnor U8073 (N_8073,N_7658,N_7673);
nand U8074 (N_8074,N_7893,N_7941);
nand U8075 (N_8075,N_7533,N_7580);
or U8076 (N_8076,N_7615,N_7544);
or U8077 (N_8077,N_7931,N_7565);
xnor U8078 (N_8078,N_7525,N_7791);
and U8079 (N_8079,N_7710,N_7994);
or U8080 (N_8080,N_7500,N_7832);
and U8081 (N_8081,N_7888,N_7798);
xor U8082 (N_8082,N_7958,N_7545);
nor U8083 (N_8083,N_7777,N_7508);
or U8084 (N_8084,N_7753,N_7864);
and U8085 (N_8085,N_7670,N_7635);
and U8086 (N_8086,N_7542,N_7745);
and U8087 (N_8087,N_7896,N_7803);
and U8088 (N_8088,N_7883,N_7835);
nor U8089 (N_8089,N_7828,N_7956);
nand U8090 (N_8090,N_7755,N_7632);
or U8091 (N_8091,N_7815,N_7982);
xor U8092 (N_8092,N_7902,N_7693);
and U8093 (N_8093,N_7722,N_7579);
xnor U8094 (N_8094,N_7607,N_7649);
nand U8095 (N_8095,N_7654,N_7861);
and U8096 (N_8096,N_7928,N_7733);
xnor U8097 (N_8097,N_7895,N_7645);
or U8098 (N_8098,N_7689,N_7758);
or U8099 (N_8099,N_7817,N_7797);
or U8100 (N_8100,N_7572,N_7633);
nand U8101 (N_8101,N_7618,N_7844);
and U8102 (N_8102,N_7516,N_7818);
or U8103 (N_8103,N_7899,N_7598);
xnor U8104 (N_8104,N_7695,N_7910);
nand U8105 (N_8105,N_7520,N_7796);
xor U8106 (N_8106,N_7631,N_7966);
xnor U8107 (N_8107,N_7775,N_7904);
and U8108 (N_8108,N_7581,N_7505);
xor U8109 (N_8109,N_7638,N_7734);
or U8110 (N_8110,N_7727,N_7606);
or U8111 (N_8111,N_7876,N_7717);
nor U8112 (N_8112,N_7934,N_7705);
or U8113 (N_8113,N_7568,N_7909);
nor U8114 (N_8114,N_7897,N_7534);
or U8115 (N_8115,N_7510,N_7718);
or U8116 (N_8116,N_7788,N_7744);
xor U8117 (N_8117,N_7860,N_7688);
or U8118 (N_8118,N_7719,N_7762);
or U8119 (N_8119,N_7754,N_7937);
and U8120 (N_8120,N_7569,N_7839);
nand U8121 (N_8121,N_7674,N_7873);
and U8122 (N_8122,N_7816,N_7882);
nand U8123 (N_8123,N_7628,N_7903);
nor U8124 (N_8124,N_7948,N_7690);
and U8125 (N_8125,N_7704,N_7697);
or U8126 (N_8126,N_7739,N_7795);
or U8127 (N_8127,N_7976,N_7949);
xor U8128 (N_8128,N_7515,N_7770);
nor U8129 (N_8129,N_7551,N_7605);
xnor U8130 (N_8130,N_7583,N_7707);
and U8131 (N_8131,N_7683,N_7560);
and U8132 (N_8132,N_7550,N_7972);
nor U8133 (N_8133,N_7831,N_7675);
and U8134 (N_8134,N_7878,N_7989);
nand U8135 (N_8135,N_7785,N_7957);
nand U8136 (N_8136,N_7504,N_7990);
and U8137 (N_8137,N_7664,N_7614);
and U8138 (N_8138,N_7503,N_7824);
nand U8139 (N_8139,N_7682,N_7644);
nand U8140 (N_8140,N_7760,N_7502);
nand U8141 (N_8141,N_7725,N_7530);
nor U8142 (N_8142,N_7810,N_7567);
nand U8143 (N_8143,N_7911,N_7752);
xnor U8144 (N_8144,N_7794,N_7799);
nor U8145 (N_8145,N_7702,N_7634);
xor U8146 (N_8146,N_7916,N_7978);
xor U8147 (N_8147,N_7586,N_7894);
nor U8148 (N_8148,N_7823,N_7987);
nand U8149 (N_8149,N_7872,N_7715);
xnor U8150 (N_8150,N_7999,N_7698);
or U8151 (N_8151,N_7602,N_7540);
nand U8152 (N_8152,N_7563,N_7747);
and U8153 (N_8153,N_7973,N_7593);
or U8154 (N_8154,N_7901,N_7703);
nor U8155 (N_8155,N_7837,N_7553);
nand U8156 (N_8156,N_7807,N_7647);
nor U8157 (N_8157,N_7667,N_7983);
nor U8158 (N_8158,N_7765,N_7512);
or U8159 (N_8159,N_7740,N_7601);
and U8160 (N_8160,N_7998,N_7812);
nor U8161 (N_8161,N_7962,N_7506);
nand U8162 (N_8162,N_7716,N_7731);
or U8163 (N_8163,N_7951,N_7639);
or U8164 (N_8164,N_7742,N_7604);
nand U8165 (N_8165,N_7857,N_7627);
and U8166 (N_8166,N_7723,N_7984);
nor U8167 (N_8167,N_7603,N_7963);
xnor U8168 (N_8168,N_7521,N_7771);
or U8169 (N_8169,N_7889,N_7677);
or U8170 (N_8170,N_7746,N_7585);
or U8171 (N_8171,N_7507,N_7804);
nor U8172 (N_8172,N_7885,N_7879);
nor U8173 (N_8173,N_7801,N_7890);
and U8174 (N_8174,N_7862,N_7840);
nand U8175 (N_8175,N_7571,N_7556);
nor U8176 (N_8176,N_7600,N_7608);
or U8177 (N_8177,N_7992,N_7546);
and U8178 (N_8178,N_7696,N_7543);
nand U8179 (N_8179,N_7562,N_7953);
xnor U8180 (N_8180,N_7588,N_7778);
nor U8181 (N_8181,N_7527,N_7781);
or U8182 (N_8182,N_7652,N_7582);
xnor U8183 (N_8183,N_7599,N_7868);
nand U8184 (N_8184,N_7561,N_7808);
nor U8185 (N_8185,N_7977,N_7566);
nor U8186 (N_8186,N_7597,N_7730);
and U8187 (N_8187,N_7924,N_7728);
or U8188 (N_8188,N_7776,N_7919);
and U8189 (N_8189,N_7905,N_7679);
nand U8190 (N_8190,N_7743,N_7611);
and U8191 (N_8191,N_7640,N_7836);
xnor U8192 (N_8192,N_7792,N_7800);
and U8193 (N_8193,N_7589,N_7870);
xor U8194 (N_8194,N_7933,N_7855);
and U8195 (N_8195,N_7756,N_7666);
nand U8196 (N_8196,N_7950,N_7648);
nand U8197 (N_8197,N_7819,N_7650);
nor U8198 (N_8198,N_7942,N_7767);
or U8199 (N_8199,N_7991,N_7557);
and U8200 (N_8200,N_7657,N_7538);
nand U8201 (N_8201,N_7867,N_7501);
nand U8202 (N_8202,N_7541,N_7663);
nor U8203 (N_8203,N_7691,N_7863);
nand U8204 (N_8204,N_7523,N_7880);
or U8205 (N_8205,N_7940,N_7859);
xnor U8206 (N_8206,N_7768,N_7592);
nand U8207 (N_8207,N_7980,N_7570);
or U8208 (N_8208,N_7576,N_7858);
and U8209 (N_8209,N_7892,N_7946);
or U8210 (N_8210,N_7925,N_7700);
or U8211 (N_8211,N_7613,N_7517);
and U8212 (N_8212,N_7578,N_7825);
nor U8213 (N_8213,N_7887,N_7641);
nand U8214 (N_8214,N_7711,N_7532);
and U8215 (N_8215,N_7877,N_7841);
nand U8216 (N_8216,N_7850,N_7681);
or U8217 (N_8217,N_7749,N_7761);
or U8218 (N_8218,N_7997,N_7574);
nor U8219 (N_8219,N_7971,N_7721);
xor U8220 (N_8220,N_7732,N_7912);
nand U8221 (N_8221,N_7547,N_7774);
nand U8222 (N_8222,N_7922,N_7830);
xnor U8223 (N_8223,N_7610,N_7847);
xor U8224 (N_8224,N_7748,N_7653);
or U8225 (N_8225,N_7724,N_7866);
nand U8226 (N_8226,N_7826,N_7526);
and U8227 (N_8227,N_7974,N_7684);
and U8228 (N_8228,N_7969,N_7988);
nand U8229 (N_8229,N_7967,N_7636);
or U8230 (N_8230,N_7549,N_7793);
and U8231 (N_8231,N_7806,N_7914);
and U8232 (N_8232,N_7575,N_7802);
nor U8233 (N_8233,N_7981,N_7612);
or U8234 (N_8234,N_7954,N_7960);
and U8235 (N_8235,N_7709,N_7920);
nand U8236 (N_8236,N_7936,N_7662);
nand U8237 (N_8237,N_7656,N_7757);
nor U8238 (N_8238,N_7680,N_7511);
or U8239 (N_8239,N_7986,N_7913);
and U8240 (N_8240,N_7784,N_7529);
or U8241 (N_8241,N_7881,N_7509);
and U8242 (N_8242,N_7616,N_7587);
xnor U8243 (N_8243,N_7764,N_7829);
and U8244 (N_8244,N_7712,N_7970);
and U8245 (N_8245,N_7944,N_7629);
or U8246 (N_8246,N_7708,N_7938);
and U8247 (N_8247,N_7955,N_7623);
nand U8248 (N_8248,N_7531,N_7554);
xor U8249 (N_8249,N_7789,N_7874);
or U8250 (N_8250,N_7975,N_7743);
and U8251 (N_8251,N_7905,N_7674);
xor U8252 (N_8252,N_7593,N_7930);
nand U8253 (N_8253,N_7692,N_7847);
nand U8254 (N_8254,N_7609,N_7644);
nor U8255 (N_8255,N_7992,N_7705);
and U8256 (N_8256,N_7855,N_7570);
nand U8257 (N_8257,N_7783,N_7615);
nor U8258 (N_8258,N_7666,N_7647);
xnor U8259 (N_8259,N_7530,N_7518);
nor U8260 (N_8260,N_7610,N_7613);
xnor U8261 (N_8261,N_7985,N_7973);
or U8262 (N_8262,N_7874,N_7703);
or U8263 (N_8263,N_7728,N_7992);
nand U8264 (N_8264,N_7887,N_7885);
nor U8265 (N_8265,N_7756,N_7587);
nor U8266 (N_8266,N_7754,N_7520);
xnor U8267 (N_8267,N_7820,N_7660);
nand U8268 (N_8268,N_7786,N_7523);
nor U8269 (N_8269,N_7806,N_7732);
nand U8270 (N_8270,N_7538,N_7680);
nor U8271 (N_8271,N_7520,N_7715);
nor U8272 (N_8272,N_7770,N_7709);
nor U8273 (N_8273,N_7601,N_7780);
nand U8274 (N_8274,N_7747,N_7649);
and U8275 (N_8275,N_7650,N_7946);
nand U8276 (N_8276,N_7906,N_7755);
xor U8277 (N_8277,N_7539,N_7615);
nand U8278 (N_8278,N_7679,N_7639);
nor U8279 (N_8279,N_7600,N_7591);
or U8280 (N_8280,N_7726,N_7905);
nor U8281 (N_8281,N_7618,N_7562);
xor U8282 (N_8282,N_7810,N_7818);
xor U8283 (N_8283,N_7604,N_7728);
nand U8284 (N_8284,N_7903,N_7827);
nand U8285 (N_8285,N_7831,N_7651);
xor U8286 (N_8286,N_7654,N_7573);
and U8287 (N_8287,N_7522,N_7983);
nand U8288 (N_8288,N_7689,N_7572);
or U8289 (N_8289,N_7880,N_7579);
nand U8290 (N_8290,N_7550,N_7714);
nand U8291 (N_8291,N_7960,N_7648);
xor U8292 (N_8292,N_7562,N_7558);
nand U8293 (N_8293,N_7715,N_7837);
nand U8294 (N_8294,N_7679,N_7574);
xor U8295 (N_8295,N_7765,N_7923);
nand U8296 (N_8296,N_7753,N_7866);
nor U8297 (N_8297,N_7790,N_7751);
or U8298 (N_8298,N_7813,N_7680);
nor U8299 (N_8299,N_7527,N_7782);
nor U8300 (N_8300,N_7849,N_7630);
xor U8301 (N_8301,N_7535,N_7896);
nand U8302 (N_8302,N_7947,N_7929);
nor U8303 (N_8303,N_7855,N_7991);
nand U8304 (N_8304,N_7676,N_7803);
or U8305 (N_8305,N_7995,N_7602);
nand U8306 (N_8306,N_7872,N_7511);
or U8307 (N_8307,N_7887,N_7523);
nand U8308 (N_8308,N_7624,N_7920);
nor U8309 (N_8309,N_7783,N_7560);
and U8310 (N_8310,N_7937,N_7989);
xnor U8311 (N_8311,N_7908,N_7562);
xor U8312 (N_8312,N_7902,N_7678);
or U8313 (N_8313,N_7702,N_7642);
nand U8314 (N_8314,N_7953,N_7827);
and U8315 (N_8315,N_7586,N_7875);
and U8316 (N_8316,N_7808,N_7677);
or U8317 (N_8317,N_7913,N_7740);
nand U8318 (N_8318,N_7798,N_7870);
xor U8319 (N_8319,N_7904,N_7893);
nand U8320 (N_8320,N_7771,N_7960);
or U8321 (N_8321,N_7596,N_7737);
nand U8322 (N_8322,N_7746,N_7849);
or U8323 (N_8323,N_7897,N_7629);
or U8324 (N_8324,N_7594,N_7816);
or U8325 (N_8325,N_7628,N_7525);
xor U8326 (N_8326,N_7869,N_7601);
or U8327 (N_8327,N_7870,N_7831);
and U8328 (N_8328,N_7544,N_7959);
xor U8329 (N_8329,N_7785,N_7674);
xor U8330 (N_8330,N_7722,N_7572);
and U8331 (N_8331,N_7543,N_7667);
or U8332 (N_8332,N_7952,N_7710);
nand U8333 (N_8333,N_7810,N_7994);
xnor U8334 (N_8334,N_7911,N_7631);
and U8335 (N_8335,N_7691,N_7813);
or U8336 (N_8336,N_7513,N_7570);
xor U8337 (N_8337,N_7808,N_7729);
xor U8338 (N_8338,N_7688,N_7702);
nor U8339 (N_8339,N_7773,N_7983);
or U8340 (N_8340,N_7608,N_7620);
or U8341 (N_8341,N_7558,N_7951);
xnor U8342 (N_8342,N_7566,N_7961);
or U8343 (N_8343,N_7847,N_7636);
or U8344 (N_8344,N_7943,N_7794);
or U8345 (N_8345,N_7763,N_7571);
nor U8346 (N_8346,N_7593,N_7817);
xnor U8347 (N_8347,N_7991,N_7976);
xnor U8348 (N_8348,N_7622,N_7840);
or U8349 (N_8349,N_7960,N_7761);
or U8350 (N_8350,N_7900,N_7748);
nor U8351 (N_8351,N_7823,N_7743);
xor U8352 (N_8352,N_7720,N_7845);
and U8353 (N_8353,N_7784,N_7775);
and U8354 (N_8354,N_7769,N_7627);
or U8355 (N_8355,N_7960,N_7825);
nor U8356 (N_8356,N_7675,N_7995);
or U8357 (N_8357,N_7589,N_7524);
or U8358 (N_8358,N_7529,N_7807);
nor U8359 (N_8359,N_7563,N_7798);
or U8360 (N_8360,N_7652,N_7684);
nor U8361 (N_8361,N_7977,N_7891);
xnor U8362 (N_8362,N_7822,N_7944);
nor U8363 (N_8363,N_7838,N_7631);
or U8364 (N_8364,N_7896,N_7801);
nand U8365 (N_8365,N_7705,N_7574);
or U8366 (N_8366,N_7590,N_7704);
and U8367 (N_8367,N_7521,N_7946);
xor U8368 (N_8368,N_7632,N_7560);
xor U8369 (N_8369,N_7984,N_7784);
or U8370 (N_8370,N_7559,N_7709);
xnor U8371 (N_8371,N_7573,N_7717);
xnor U8372 (N_8372,N_7533,N_7860);
nand U8373 (N_8373,N_7939,N_7923);
and U8374 (N_8374,N_7591,N_7617);
xnor U8375 (N_8375,N_7534,N_7978);
xor U8376 (N_8376,N_7981,N_7833);
nand U8377 (N_8377,N_7877,N_7972);
nand U8378 (N_8378,N_7556,N_7515);
or U8379 (N_8379,N_7686,N_7824);
nand U8380 (N_8380,N_7713,N_7793);
or U8381 (N_8381,N_7851,N_7948);
or U8382 (N_8382,N_7971,N_7535);
and U8383 (N_8383,N_7866,N_7674);
or U8384 (N_8384,N_7846,N_7939);
or U8385 (N_8385,N_7865,N_7719);
or U8386 (N_8386,N_7868,N_7626);
and U8387 (N_8387,N_7685,N_7988);
and U8388 (N_8388,N_7602,N_7631);
nor U8389 (N_8389,N_7631,N_7686);
xor U8390 (N_8390,N_7943,N_7605);
xor U8391 (N_8391,N_7956,N_7699);
nand U8392 (N_8392,N_7506,N_7566);
nor U8393 (N_8393,N_7942,N_7750);
or U8394 (N_8394,N_7778,N_7938);
nor U8395 (N_8395,N_7658,N_7501);
xnor U8396 (N_8396,N_7618,N_7569);
or U8397 (N_8397,N_7941,N_7756);
nand U8398 (N_8398,N_7830,N_7913);
and U8399 (N_8399,N_7704,N_7678);
and U8400 (N_8400,N_7582,N_7747);
xnor U8401 (N_8401,N_7744,N_7677);
nor U8402 (N_8402,N_7638,N_7964);
or U8403 (N_8403,N_7666,N_7734);
or U8404 (N_8404,N_7867,N_7774);
xnor U8405 (N_8405,N_7788,N_7872);
xnor U8406 (N_8406,N_7704,N_7587);
and U8407 (N_8407,N_7618,N_7944);
and U8408 (N_8408,N_7771,N_7989);
or U8409 (N_8409,N_7582,N_7526);
nor U8410 (N_8410,N_7511,N_7512);
xor U8411 (N_8411,N_7931,N_7742);
nand U8412 (N_8412,N_7980,N_7718);
nor U8413 (N_8413,N_7847,N_7743);
or U8414 (N_8414,N_7870,N_7890);
or U8415 (N_8415,N_7588,N_7734);
xor U8416 (N_8416,N_7590,N_7541);
nand U8417 (N_8417,N_7508,N_7948);
nor U8418 (N_8418,N_7617,N_7594);
xnor U8419 (N_8419,N_7561,N_7954);
xor U8420 (N_8420,N_7673,N_7825);
xor U8421 (N_8421,N_7886,N_7540);
nand U8422 (N_8422,N_7504,N_7914);
and U8423 (N_8423,N_7747,N_7862);
xnor U8424 (N_8424,N_7504,N_7733);
xnor U8425 (N_8425,N_7804,N_7934);
nand U8426 (N_8426,N_7650,N_7518);
and U8427 (N_8427,N_7841,N_7710);
and U8428 (N_8428,N_7565,N_7618);
and U8429 (N_8429,N_7693,N_7772);
and U8430 (N_8430,N_7719,N_7634);
nor U8431 (N_8431,N_7523,N_7552);
and U8432 (N_8432,N_7543,N_7685);
or U8433 (N_8433,N_7865,N_7876);
or U8434 (N_8434,N_7684,N_7834);
nor U8435 (N_8435,N_7740,N_7978);
and U8436 (N_8436,N_7636,N_7581);
nor U8437 (N_8437,N_7787,N_7707);
nor U8438 (N_8438,N_7941,N_7993);
or U8439 (N_8439,N_7612,N_7636);
xnor U8440 (N_8440,N_7983,N_7734);
nand U8441 (N_8441,N_7824,N_7506);
nor U8442 (N_8442,N_7875,N_7545);
xnor U8443 (N_8443,N_7879,N_7699);
and U8444 (N_8444,N_7569,N_7630);
nor U8445 (N_8445,N_7656,N_7613);
xor U8446 (N_8446,N_7898,N_7954);
and U8447 (N_8447,N_7502,N_7939);
and U8448 (N_8448,N_7527,N_7507);
xor U8449 (N_8449,N_7875,N_7890);
or U8450 (N_8450,N_7679,N_7968);
nand U8451 (N_8451,N_7836,N_7690);
nor U8452 (N_8452,N_7626,N_7821);
or U8453 (N_8453,N_7838,N_7618);
nor U8454 (N_8454,N_7969,N_7840);
xnor U8455 (N_8455,N_7673,N_7781);
nor U8456 (N_8456,N_7959,N_7704);
nor U8457 (N_8457,N_7948,N_7784);
nand U8458 (N_8458,N_7610,N_7575);
and U8459 (N_8459,N_7912,N_7510);
and U8460 (N_8460,N_7842,N_7738);
nand U8461 (N_8461,N_7905,N_7884);
or U8462 (N_8462,N_7545,N_7638);
xnor U8463 (N_8463,N_7957,N_7958);
nor U8464 (N_8464,N_7658,N_7703);
and U8465 (N_8465,N_7918,N_7892);
nor U8466 (N_8466,N_7744,N_7698);
xor U8467 (N_8467,N_7869,N_7576);
nand U8468 (N_8468,N_7520,N_7848);
nand U8469 (N_8469,N_7539,N_7861);
nor U8470 (N_8470,N_7722,N_7584);
nor U8471 (N_8471,N_7697,N_7647);
and U8472 (N_8472,N_7640,N_7838);
xnor U8473 (N_8473,N_7847,N_7821);
xor U8474 (N_8474,N_7884,N_7896);
nor U8475 (N_8475,N_7986,N_7571);
and U8476 (N_8476,N_7639,N_7654);
or U8477 (N_8477,N_7818,N_7521);
and U8478 (N_8478,N_7883,N_7812);
xor U8479 (N_8479,N_7985,N_7771);
nor U8480 (N_8480,N_7798,N_7847);
nand U8481 (N_8481,N_7603,N_7736);
nor U8482 (N_8482,N_7564,N_7605);
nand U8483 (N_8483,N_7914,N_7634);
or U8484 (N_8484,N_7891,N_7949);
nand U8485 (N_8485,N_7876,N_7835);
or U8486 (N_8486,N_7845,N_7572);
or U8487 (N_8487,N_7826,N_7667);
xnor U8488 (N_8488,N_7515,N_7917);
and U8489 (N_8489,N_7539,N_7521);
or U8490 (N_8490,N_7671,N_7681);
xnor U8491 (N_8491,N_7540,N_7527);
or U8492 (N_8492,N_7835,N_7755);
and U8493 (N_8493,N_7878,N_7595);
and U8494 (N_8494,N_7627,N_7916);
and U8495 (N_8495,N_7853,N_7851);
xnor U8496 (N_8496,N_7851,N_7996);
or U8497 (N_8497,N_7916,N_7554);
nor U8498 (N_8498,N_7755,N_7896);
nor U8499 (N_8499,N_7610,N_7889);
or U8500 (N_8500,N_8487,N_8414);
and U8501 (N_8501,N_8402,N_8083);
and U8502 (N_8502,N_8302,N_8086);
nand U8503 (N_8503,N_8091,N_8303);
or U8504 (N_8504,N_8132,N_8445);
xnor U8505 (N_8505,N_8113,N_8022);
nand U8506 (N_8506,N_8189,N_8215);
nand U8507 (N_8507,N_8028,N_8385);
and U8508 (N_8508,N_8155,N_8390);
nor U8509 (N_8509,N_8059,N_8260);
xor U8510 (N_8510,N_8158,N_8250);
nand U8511 (N_8511,N_8437,N_8239);
nand U8512 (N_8512,N_8478,N_8165);
nand U8513 (N_8513,N_8248,N_8288);
xnor U8514 (N_8514,N_8055,N_8245);
nor U8515 (N_8515,N_8072,N_8344);
and U8516 (N_8516,N_8384,N_8470);
nand U8517 (N_8517,N_8000,N_8401);
nand U8518 (N_8518,N_8221,N_8271);
or U8519 (N_8519,N_8289,N_8297);
nand U8520 (N_8520,N_8228,N_8004);
xor U8521 (N_8521,N_8448,N_8143);
xnor U8522 (N_8522,N_8298,N_8047);
nor U8523 (N_8523,N_8197,N_8495);
nand U8524 (N_8524,N_8074,N_8415);
nand U8525 (N_8525,N_8396,N_8227);
nor U8526 (N_8526,N_8099,N_8032);
xor U8527 (N_8527,N_8188,N_8326);
and U8528 (N_8528,N_8244,N_8089);
nand U8529 (N_8529,N_8411,N_8482);
nor U8530 (N_8530,N_8125,N_8264);
and U8531 (N_8531,N_8345,N_8167);
or U8532 (N_8532,N_8233,N_8397);
nand U8533 (N_8533,N_8035,N_8333);
or U8534 (N_8534,N_8217,N_8229);
xor U8535 (N_8535,N_8472,N_8037);
or U8536 (N_8536,N_8494,N_8433);
xor U8537 (N_8537,N_8013,N_8316);
and U8538 (N_8538,N_8340,N_8422);
nor U8539 (N_8539,N_8080,N_8408);
nand U8540 (N_8540,N_8262,N_8452);
nand U8541 (N_8541,N_8023,N_8182);
nor U8542 (N_8542,N_8446,N_8123);
and U8543 (N_8543,N_8281,N_8025);
and U8544 (N_8544,N_8336,N_8351);
nor U8545 (N_8545,N_8142,N_8034);
nand U8546 (N_8546,N_8153,N_8421);
nor U8547 (N_8547,N_8021,N_8195);
and U8548 (N_8548,N_8010,N_8413);
nand U8549 (N_8549,N_8135,N_8111);
or U8550 (N_8550,N_8443,N_8367);
nor U8551 (N_8551,N_8436,N_8139);
nor U8552 (N_8552,N_8290,N_8134);
and U8553 (N_8553,N_8185,N_8180);
nand U8554 (N_8554,N_8184,N_8343);
nand U8555 (N_8555,N_8369,N_8358);
xor U8556 (N_8556,N_8283,N_8451);
or U8557 (N_8557,N_8231,N_8306);
xor U8558 (N_8558,N_8323,N_8160);
or U8559 (N_8559,N_8027,N_8218);
nand U8560 (N_8560,N_8002,N_8320);
nor U8561 (N_8561,N_8166,N_8267);
xnor U8562 (N_8562,N_8026,N_8430);
nor U8563 (N_8563,N_8104,N_8040);
nand U8564 (N_8564,N_8109,N_8088);
or U8565 (N_8565,N_8243,N_8151);
nor U8566 (N_8566,N_8129,N_8148);
nor U8567 (N_8567,N_8386,N_8137);
or U8568 (N_8568,N_8416,N_8489);
xor U8569 (N_8569,N_8439,N_8405);
or U8570 (N_8570,N_8168,N_8014);
or U8571 (N_8571,N_8241,N_8286);
xnor U8572 (N_8572,N_8057,N_8033);
or U8573 (N_8573,N_8361,N_8442);
nand U8574 (N_8574,N_8273,N_8467);
and U8575 (N_8575,N_8092,N_8146);
xnor U8576 (N_8576,N_8419,N_8031);
and U8577 (N_8577,N_8349,N_8206);
nand U8578 (N_8578,N_8268,N_8363);
or U8579 (N_8579,N_8331,N_8308);
or U8580 (N_8580,N_8276,N_8012);
or U8581 (N_8581,N_8424,N_8496);
nand U8582 (N_8582,N_8486,N_8199);
xnor U8583 (N_8583,N_8310,N_8152);
xnor U8584 (N_8584,N_8140,N_8087);
xnor U8585 (N_8585,N_8178,N_8058);
and U8586 (N_8586,N_8275,N_8319);
nand U8587 (N_8587,N_8485,N_8157);
xor U8588 (N_8588,N_8019,N_8016);
nor U8589 (N_8589,N_8200,N_8079);
and U8590 (N_8590,N_8247,N_8252);
nor U8591 (N_8591,N_8391,N_8253);
or U8592 (N_8592,N_8371,N_8440);
nor U8593 (N_8593,N_8350,N_8382);
or U8594 (N_8594,N_8327,N_8145);
nand U8595 (N_8595,N_8270,N_8300);
nor U8596 (N_8596,N_8175,N_8434);
xnor U8597 (N_8597,N_8054,N_8214);
xor U8598 (N_8598,N_8417,N_8194);
and U8599 (N_8599,N_8108,N_8362);
xnor U8600 (N_8600,N_8220,N_8469);
nor U8601 (N_8601,N_8406,N_8041);
or U8602 (N_8602,N_8438,N_8435);
nand U8603 (N_8603,N_8115,N_8201);
or U8604 (N_8604,N_8211,N_8096);
or U8605 (N_8605,N_8387,N_8461);
or U8606 (N_8606,N_8093,N_8173);
and U8607 (N_8607,N_8258,N_8141);
nor U8608 (N_8608,N_8128,N_8193);
nor U8609 (N_8609,N_8466,N_8352);
nor U8610 (N_8610,N_8492,N_8068);
or U8611 (N_8611,N_8429,N_8063);
nor U8612 (N_8612,N_8324,N_8179);
nand U8613 (N_8613,N_8024,N_8356);
nor U8614 (N_8614,N_8118,N_8381);
nand U8615 (N_8615,N_8368,N_8069);
or U8616 (N_8616,N_8280,N_8263);
and U8617 (N_8617,N_8164,N_8081);
nand U8618 (N_8618,N_8348,N_8293);
nor U8619 (N_8619,N_8427,N_8048);
xor U8620 (N_8620,N_8307,N_8388);
and U8621 (N_8621,N_8045,N_8374);
xor U8622 (N_8622,N_8360,N_8066);
or U8623 (N_8623,N_8464,N_8292);
xnor U8624 (N_8624,N_8106,N_8432);
and U8625 (N_8625,N_8428,N_8236);
nor U8626 (N_8626,N_8459,N_8001);
nor U8627 (N_8627,N_8061,N_8299);
xnor U8628 (N_8628,N_8313,N_8304);
and U8629 (N_8629,N_8084,N_8062);
xnor U8630 (N_8630,N_8223,N_8107);
and U8631 (N_8631,N_8038,N_8412);
nor U8632 (N_8632,N_8491,N_8124);
xor U8633 (N_8633,N_8242,N_8208);
and U8634 (N_8634,N_8377,N_8196);
or U8635 (N_8635,N_8046,N_8156);
and U8636 (N_8636,N_8015,N_8207);
nor U8637 (N_8637,N_8269,N_8305);
or U8638 (N_8638,N_8373,N_8121);
and U8639 (N_8639,N_8076,N_8234);
and U8640 (N_8640,N_8176,N_8477);
xor U8641 (N_8641,N_8119,N_8383);
or U8642 (N_8642,N_8117,N_8257);
xor U8643 (N_8643,N_8481,N_8105);
nand U8644 (N_8644,N_8449,N_8409);
or U8645 (N_8645,N_8030,N_8431);
nand U8646 (N_8646,N_8222,N_8232);
xnor U8647 (N_8647,N_8177,N_8100);
or U8648 (N_8648,N_8169,N_8309);
nor U8649 (N_8649,N_8353,N_8296);
xor U8650 (N_8650,N_8237,N_8370);
nor U8651 (N_8651,N_8455,N_8127);
or U8652 (N_8652,N_8005,N_8407);
nor U8653 (N_8653,N_8454,N_8395);
xor U8654 (N_8654,N_8339,N_8204);
or U8655 (N_8655,N_8183,N_8056);
nor U8656 (N_8656,N_8103,N_8163);
or U8657 (N_8657,N_8488,N_8457);
xnor U8658 (N_8658,N_8050,N_8404);
nor U8659 (N_8659,N_8380,N_8065);
nand U8660 (N_8660,N_8301,N_8479);
xor U8661 (N_8661,N_8256,N_8161);
or U8662 (N_8662,N_8147,N_8219);
xor U8663 (N_8663,N_8043,N_8097);
nor U8664 (N_8664,N_8272,N_8473);
or U8665 (N_8665,N_8060,N_8044);
or U8666 (N_8666,N_8354,N_8052);
or U8667 (N_8667,N_8372,N_8235);
xnor U8668 (N_8668,N_8483,N_8498);
or U8669 (N_8669,N_8322,N_8202);
or U8670 (N_8670,N_8480,N_8493);
nor U8671 (N_8671,N_8205,N_8246);
nand U8672 (N_8672,N_8364,N_8213);
nand U8673 (N_8673,N_8447,N_8330);
nor U8674 (N_8674,N_8067,N_8410);
xnor U8675 (N_8675,N_8116,N_8418);
or U8676 (N_8676,N_8029,N_8328);
xnor U8677 (N_8677,N_8334,N_8441);
xor U8678 (N_8678,N_8475,N_8036);
or U8679 (N_8679,N_8006,N_8130);
or U8680 (N_8680,N_8332,N_8203);
nor U8681 (N_8681,N_8314,N_8317);
and U8682 (N_8682,N_8463,N_8138);
and U8683 (N_8683,N_8020,N_8376);
or U8684 (N_8684,N_8378,N_8359);
and U8685 (N_8685,N_8277,N_8077);
or U8686 (N_8686,N_8017,N_8249);
nor U8687 (N_8687,N_8484,N_8174);
nand U8688 (N_8688,N_8279,N_8321);
nand U8689 (N_8689,N_8133,N_8171);
nor U8690 (N_8690,N_8187,N_8122);
nand U8691 (N_8691,N_8366,N_8311);
and U8692 (N_8692,N_8450,N_8254);
xnor U8693 (N_8693,N_8460,N_8073);
or U8694 (N_8694,N_8325,N_8216);
and U8695 (N_8695,N_8192,N_8315);
and U8696 (N_8696,N_8008,N_8172);
nand U8697 (N_8697,N_8346,N_8042);
and U8698 (N_8698,N_8393,N_8265);
nor U8699 (N_8699,N_8468,N_8101);
or U8700 (N_8700,N_8394,N_8181);
nor U8701 (N_8701,N_8126,N_8347);
nor U8702 (N_8702,N_8085,N_8186);
nor U8703 (N_8703,N_8078,N_8259);
nor U8704 (N_8704,N_8170,N_8357);
nand U8705 (N_8705,N_8120,N_8154);
nor U8706 (N_8706,N_8114,N_8190);
nor U8707 (N_8707,N_8497,N_8337);
or U8708 (N_8708,N_8039,N_8426);
nor U8709 (N_8709,N_8284,N_8490);
nor U8710 (N_8710,N_8191,N_8110);
or U8711 (N_8711,N_8285,N_8458);
xnor U8712 (N_8712,N_8075,N_8212);
nand U8713 (N_8713,N_8420,N_8341);
nor U8714 (N_8714,N_8112,N_8082);
nand U8715 (N_8715,N_8403,N_8294);
nor U8716 (N_8716,N_8499,N_8365);
and U8717 (N_8717,N_8329,N_8266);
and U8718 (N_8718,N_8282,N_8102);
nor U8719 (N_8719,N_8098,N_8136);
or U8720 (N_8720,N_8342,N_8150);
xnor U8721 (N_8721,N_8226,N_8159);
and U8722 (N_8722,N_8251,N_8453);
xnor U8723 (N_8723,N_8274,N_8291);
and U8724 (N_8724,N_8425,N_8476);
and U8725 (N_8725,N_8240,N_8144);
or U8726 (N_8726,N_8198,N_8399);
nand U8727 (N_8727,N_8278,N_8295);
nand U8728 (N_8728,N_8011,N_8465);
and U8729 (N_8729,N_8287,N_8095);
xor U8730 (N_8730,N_8312,N_8462);
or U8731 (N_8731,N_8375,N_8009);
xor U8732 (N_8732,N_8051,N_8444);
and U8733 (N_8733,N_8355,N_8335);
and U8734 (N_8734,N_8094,N_8053);
and U8735 (N_8735,N_8400,N_8090);
xor U8736 (N_8736,N_8224,N_8003);
nand U8737 (N_8737,N_8070,N_8389);
and U8738 (N_8738,N_8162,N_8474);
nor U8739 (N_8739,N_8209,N_8338);
nand U8740 (N_8740,N_8423,N_8261);
and U8741 (N_8741,N_8225,N_8149);
xnor U8742 (N_8742,N_8318,N_8456);
nand U8743 (N_8743,N_8131,N_8018);
or U8744 (N_8744,N_8238,N_8379);
nor U8745 (N_8745,N_8471,N_8392);
nor U8746 (N_8746,N_8398,N_8007);
xnor U8747 (N_8747,N_8210,N_8049);
or U8748 (N_8748,N_8255,N_8071);
or U8749 (N_8749,N_8064,N_8230);
or U8750 (N_8750,N_8405,N_8253);
and U8751 (N_8751,N_8218,N_8019);
nand U8752 (N_8752,N_8069,N_8105);
nand U8753 (N_8753,N_8111,N_8171);
or U8754 (N_8754,N_8008,N_8183);
xor U8755 (N_8755,N_8130,N_8393);
nand U8756 (N_8756,N_8245,N_8472);
or U8757 (N_8757,N_8236,N_8283);
or U8758 (N_8758,N_8358,N_8312);
nor U8759 (N_8759,N_8361,N_8377);
nand U8760 (N_8760,N_8212,N_8432);
nand U8761 (N_8761,N_8464,N_8146);
and U8762 (N_8762,N_8381,N_8439);
xor U8763 (N_8763,N_8309,N_8388);
xor U8764 (N_8764,N_8135,N_8002);
nand U8765 (N_8765,N_8322,N_8111);
and U8766 (N_8766,N_8046,N_8257);
xnor U8767 (N_8767,N_8116,N_8024);
nand U8768 (N_8768,N_8164,N_8151);
or U8769 (N_8769,N_8446,N_8432);
or U8770 (N_8770,N_8254,N_8277);
nor U8771 (N_8771,N_8136,N_8075);
or U8772 (N_8772,N_8052,N_8398);
nor U8773 (N_8773,N_8478,N_8090);
nand U8774 (N_8774,N_8258,N_8315);
nand U8775 (N_8775,N_8368,N_8158);
xnor U8776 (N_8776,N_8131,N_8401);
xor U8777 (N_8777,N_8428,N_8037);
and U8778 (N_8778,N_8323,N_8296);
or U8779 (N_8779,N_8267,N_8365);
xor U8780 (N_8780,N_8358,N_8016);
xnor U8781 (N_8781,N_8020,N_8123);
and U8782 (N_8782,N_8366,N_8386);
and U8783 (N_8783,N_8169,N_8425);
nand U8784 (N_8784,N_8366,N_8290);
xor U8785 (N_8785,N_8011,N_8313);
xor U8786 (N_8786,N_8468,N_8195);
and U8787 (N_8787,N_8451,N_8245);
nor U8788 (N_8788,N_8136,N_8349);
xnor U8789 (N_8789,N_8461,N_8120);
or U8790 (N_8790,N_8273,N_8449);
xnor U8791 (N_8791,N_8151,N_8256);
nor U8792 (N_8792,N_8416,N_8258);
nor U8793 (N_8793,N_8158,N_8283);
xnor U8794 (N_8794,N_8217,N_8189);
nor U8795 (N_8795,N_8366,N_8310);
nand U8796 (N_8796,N_8181,N_8239);
or U8797 (N_8797,N_8397,N_8371);
nor U8798 (N_8798,N_8069,N_8440);
or U8799 (N_8799,N_8044,N_8018);
xnor U8800 (N_8800,N_8048,N_8035);
xor U8801 (N_8801,N_8498,N_8447);
or U8802 (N_8802,N_8044,N_8299);
nor U8803 (N_8803,N_8222,N_8475);
or U8804 (N_8804,N_8038,N_8161);
nand U8805 (N_8805,N_8461,N_8133);
nand U8806 (N_8806,N_8320,N_8005);
nor U8807 (N_8807,N_8205,N_8018);
nor U8808 (N_8808,N_8181,N_8416);
or U8809 (N_8809,N_8127,N_8401);
nor U8810 (N_8810,N_8224,N_8371);
xnor U8811 (N_8811,N_8464,N_8127);
nor U8812 (N_8812,N_8447,N_8452);
nor U8813 (N_8813,N_8381,N_8013);
and U8814 (N_8814,N_8158,N_8219);
nand U8815 (N_8815,N_8356,N_8206);
and U8816 (N_8816,N_8231,N_8132);
nor U8817 (N_8817,N_8423,N_8409);
xor U8818 (N_8818,N_8343,N_8125);
nor U8819 (N_8819,N_8278,N_8473);
nor U8820 (N_8820,N_8117,N_8439);
or U8821 (N_8821,N_8498,N_8213);
nor U8822 (N_8822,N_8218,N_8407);
xnor U8823 (N_8823,N_8287,N_8442);
and U8824 (N_8824,N_8349,N_8215);
nor U8825 (N_8825,N_8141,N_8467);
nor U8826 (N_8826,N_8457,N_8296);
and U8827 (N_8827,N_8275,N_8271);
xnor U8828 (N_8828,N_8320,N_8256);
nand U8829 (N_8829,N_8443,N_8139);
nor U8830 (N_8830,N_8430,N_8055);
nor U8831 (N_8831,N_8436,N_8112);
xor U8832 (N_8832,N_8482,N_8367);
or U8833 (N_8833,N_8214,N_8296);
nand U8834 (N_8834,N_8318,N_8396);
nor U8835 (N_8835,N_8158,N_8278);
nand U8836 (N_8836,N_8265,N_8296);
xor U8837 (N_8837,N_8187,N_8302);
and U8838 (N_8838,N_8153,N_8408);
nand U8839 (N_8839,N_8497,N_8480);
nand U8840 (N_8840,N_8048,N_8434);
xnor U8841 (N_8841,N_8174,N_8061);
xnor U8842 (N_8842,N_8364,N_8244);
and U8843 (N_8843,N_8325,N_8376);
nor U8844 (N_8844,N_8151,N_8159);
nor U8845 (N_8845,N_8234,N_8469);
and U8846 (N_8846,N_8429,N_8170);
xor U8847 (N_8847,N_8394,N_8446);
nor U8848 (N_8848,N_8122,N_8430);
nor U8849 (N_8849,N_8444,N_8213);
and U8850 (N_8850,N_8150,N_8113);
nor U8851 (N_8851,N_8285,N_8035);
nand U8852 (N_8852,N_8319,N_8231);
and U8853 (N_8853,N_8021,N_8392);
xnor U8854 (N_8854,N_8232,N_8420);
or U8855 (N_8855,N_8182,N_8218);
nor U8856 (N_8856,N_8171,N_8381);
or U8857 (N_8857,N_8439,N_8409);
or U8858 (N_8858,N_8301,N_8092);
or U8859 (N_8859,N_8367,N_8152);
and U8860 (N_8860,N_8206,N_8016);
and U8861 (N_8861,N_8013,N_8336);
nand U8862 (N_8862,N_8299,N_8078);
nor U8863 (N_8863,N_8440,N_8280);
nand U8864 (N_8864,N_8069,N_8435);
nand U8865 (N_8865,N_8389,N_8313);
nor U8866 (N_8866,N_8098,N_8195);
xor U8867 (N_8867,N_8467,N_8377);
nor U8868 (N_8868,N_8159,N_8413);
or U8869 (N_8869,N_8456,N_8187);
and U8870 (N_8870,N_8211,N_8369);
and U8871 (N_8871,N_8348,N_8063);
nor U8872 (N_8872,N_8061,N_8217);
xnor U8873 (N_8873,N_8226,N_8134);
xnor U8874 (N_8874,N_8220,N_8459);
nor U8875 (N_8875,N_8122,N_8327);
nor U8876 (N_8876,N_8088,N_8259);
nor U8877 (N_8877,N_8217,N_8162);
nand U8878 (N_8878,N_8003,N_8181);
and U8879 (N_8879,N_8472,N_8203);
and U8880 (N_8880,N_8164,N_8057);
nor U8881 (N_8881,N_8205,N_8307);
nor U8882 (N_8882,N_8143,N_8285);
nand U8883 (N_8883,N_8273,N_8109);
or U8884 (N_8884,N_8462,N_8426);
nor U8885 (N_8885,N_8061,N_8068);
xnor U8886 (N_8886,N_8462,N_8220);
nor U8887 (N_8887,N_8258,N_8471);
and U8888 (N_8888,N_8331,N_8435);
nand U8889 (N_8889,N_8361,N_8414);
and U8890 (N_8890,N_8363,N_8113);
and U8891 (N_8891,N_8352,N_8105);
and U8892 (N_8892,N_8141,N_8013);
or U8893 (N_8893,N_8377,N_8396);
and U8894 (N_8894,N_8055,N_8469);
nor U8895 (N_8895,N_8281,N_8331);
xor U8896 (N_8896,N_8093,N_8218);
nand U8897 (N_8897,N_8393,N_8357);
or U8898 (N_8898,N_8123,N_8420);
and U8899 (N_8899,N_8249,N_8496);
or U8900 (N_8900,N_8075,N_8323);
or U8901 (N_8901,N_8220,N_8104);
nand U8902 (N_8902,N_8283,N_8171);
or U8903 (N_8903,N_8271,N_8159);
and U8904 (N_8904,N_8352,N_8128);
and U8905 (N_8905,N_8451,N_8016);
and U8906 (N_8906,N_8021,N_8001);
or U8907 (N_8907,N_8198,N_8152);
nor U8908 (N_8908,N_8240,N_8314);
nand U8909 (N_8909,N_8238,N_8256);
and U8910 (N_8910,N_8428,N_8427);
nor U8911 (N_8911,N_8000,N_8166);
nand U8912 (N_8912,N_8234,N_8120);
and U8913 (N_8913,N_8431,N_8248);
xor U8914 (N_8914,N_8357,N_8440);
or U8915 (N_8915,N_8077,N_8310);
or U8916 (N_8916,N_8319,N_8389);
nand U8917 (N_8917,N_8046,N_8236);
xor U8918 (N_8918,N_8011,N_8411);
nand U8919 (N_8919,N_8066,N_8499);
nor U8920 (N_8920,N_8061,N_8355);
or U8921 (N_8921,N_8180,N_8458);
xor U8922 (N_8922,N_8418,N_8361);
xor U8923 (N_8923,N_8271,N_8134);
or U8924 (N_8924,N_8047,N_8244);
and U8925 (N_8925,N_8475,N_8185);
nand U8926 (N_8926,N_8193,N_8084);
nor U8927 (N_8927,N_8306,N_8152);
nor U8928 (N_8928,N_8090,N_8065);
and U8929 (N_8929,N_8330,N_8445);
and U8930 (N_8930,N_8474,N_8287);
xnor U8931 (N_8931,N_8003,N_8438);
and U8932 (N_8932,N_8280,N_8057);
xor U8933 (N_8933,N_8196,N_8001);
and U8934 (N_8934,N_8070,N_8207);
xor U8935 (N_8935,N_8265,N_8088);
xor U8936 (N_8936,N_8376,N_8472);
and U8937 (N_8937,N_8159,N_8175);
or U8938 (N_8938,N_8315,N_8424);
and U8939 (N_8939,N_8300,N_8236);
nand U8940 (N_8940,N_8058,N_8258);
nor U8941 (N_8941,N_8045,N_8057);
nor U8942 (N_8942,N_8410,N_8360);
nor U8943 (N_8943,N_8188,N_8467);
xor U8944 (N_8944,N_8377,N_8344);
nand U8945 (N_8945,N_8499,N_8487);
xnor U8946 (N_8946,N_8182,N_8149);
nor U8947 (N_8947,N_8264,N_8386);
xor U8948 (N_8948,N_8306,N_8390);
xor U8949 (N_8949,N_8241,N_8090);
and U8950 (N_8950,N_8335,N_8346);
and U8951 (N_8951,N_8061,N_8110);
and U8952 (N_8952,N_8417,N_8240);
xor U8953 (N_8953,N_8447,N_8410);
or U8954 (N_8954,N_8270,N_8206);
xnor U8955 (N_8955,N_8174,N_8157);
or U8956 (N_8956,N_8463,N_8391);
xor U8957 (N_8957,N_8426,N_8409);
nor U8958 (N_8958,N_8427,N_8307);
and U8959 (N_8959,N_8178,N_8121);
nand U8960 (N_8960,N_8090,N_8358);
nor U8961 (N_8961,N_8485,N_8371);
xnor U8962 (N_8962,N_8470,N_8227);
nor U8963 (N_8963,N_8248,N_8103);
or U8964 (N_8964,N_8436,N_8073);
nor U8965 (N_8965,N_8284,N_8313);
or U8966 (N_8966,N_8302,N_8251);
and U8967 (N_8967,N_8222,N_8089);
and U8968 (N_8968,N_8088,N_8171);
or U8969 (N_8969,N_8301,N_8009);
nor U8970 (N_8970,N_8436,N_8393);
or U8971 (N_8971,N_8474,N_8236);
nand U8972 (N_8972,N_8152,N_8173);
nand U8973 (N_8973,N_8302,N_8039);
or U8974 (N_8974,N_8432,N_8002);
nand U8975 (N_8975,N_8087,N_8441);
and U8976 (N_8976,N_8034,N_8398);
or U8977 (N_8977,N_8257,N_8144);
nor U8978 (N_8978,N_8361,N_8245);
nand U8979 (N_8979,N_8499,N_8332);
or U8980 (N_8980,N_8140,N_8463);
xnor U8981 (N_8981,N_8095,N_8239);
or U8982 (N_8982,N_8110,N_8308);
nand U8983 (N_8983,N_8437,N_8490);
nor U8984 (N_8984,N_8113,N_8013);
or U8985 (N_8985,N_8038,N_8003);
nor U8986 (N_8986,N_8002,N_8024);
or U8987 (N_8987,N_8495,N_8116);
and U8988 (N_8988,N_8014,N_8459);
nor U8989 (N_8989,N_8207,N_8151);
nor U8990 (N_8990,N_8338,N_8380);
and U8991 (N_8991,N_8021,N_8428);
or U8992 (N_8992,N_8469,N_8136);
nor U8993 (N_8993,N_8146,N_8396);
nor U8994 (N_8994,N_8267,N_8061);
and U8995 (N_8995,N_8265,N_8176);
nand U8996 (N_8996,N_8223,N_8344);
nor U8997 (N_8997,N_8448,N_8266);
and U8998 (N_8998,N_8386,N_8176);
or U8999 (N_8999,N_8041,N_8304);
xor U9000 (N_9000,N_8699,N_8558);
xnor U9001 (N_9001,N_8506,N_8955);
or U9002 (N_9002,N_8711,N_8574);
nor U9003 (N_9003,N_8872,N_8912);
xor U9004 (N_9004,N_8635,N_8556);
or U9005 (N_9005,N_8938,N_8777);
nand U9006 (N_9006,N_8819,N_8508);
and U9007 (N_9007,N_8946,N_8940);
xor U9008 (N_9008,N_8573,N_8809);
xor U9009 (N_9009,N_8862,N_8870);
nor U9010 (N_9010,N_8646,N_8701);
nor U9011 (N_9011,N_8666,N_8764);
nand U9012 (N_9012,N_8902,N_8947);
nor U9013 (N_9013,N_8697,N_8683);
xor U9014 (N_9014,N_8948,N_8869);
nand U9015 (N_9015,N_8537,N_8682);
nor U9016 (N_9016,N_8518,N_8904);
or U9017 (N_9017,N_8734,N_8964);
nand U9018 (N_9018,N_8926,N_8694);
nor U9019 (N_9019,N_8905,N_8765);
or U9020 (N_9020,N_8957,N_8769);
xnor U9021 (N_9021,N_8873,N_8929);
nand U9022 (N_9022,N_8811,N_8989);
and U9023 (N_9023,N_8559,N_8587);
or U9024 (N_9024,N_8932,N_8562);
or U9025 (N_9025,N_8742,N_8795);
xor U9026 (N_9026,N_8998,N_8738);
and U9027 (N_9027,N_8833,N_8804);
nor U9028 (N_9028,N_8667,N_8831);
nand U9029 (N_9029,N_8823,N_8640);
nand U9030 (N_9030,N_8676,N_8914);
nand U9031 (N_9031,N_8544,N_8951);
nand U9032 (N_9032,N_8967,N_8882);
nand U9033 (N_9033,N_8585,N_8776);
xor U9034 (N_9034,N_8898,N_8561);
or U9035 (N_9035,N_8737,N_8568);
nor U9036 (N_9036,N_8856,N_8810);
or U9037 (N_9037,N_8690,N_8606);
or U9038 (N_9038,N_8661,N_8704);
nor U9039 (N_9039,N_8663,N_8834);
or U9040 (N_9040,N_8579,N_8796);
xor U9041 (N_9041,N_8766,N_8582);
or U9042 (N_9042,N_8911,N_8524);
nor U9043 (N_9043,N_8637,N_8603);
xor U9044 (N_9044,N_8794,N_8624);
or U9045 (N_9045,N_8907,N_8725);
or U9046 (N_9046,N_8773,N_8527);
xnor U9047 (N_9047,N_8591,N_8961);
or U9048 (N_9048,N_8801,N_8913);
xor U9049 (N_9049,N_8772,N_8876);
or U9050 (N_9050,N_8761,N_8588);
xnor U9051 (N_9051,N_8741,N_8950);
nor U9052 (N_9052,N_8539,N_8861);
or U9053 (N_9053,N_8540,N_8596);
or U9054 (N_9054,N_8548,N_8505);
xor U9055 (N_9055,N_8726,N_8620);
nor U9056 (N_9056,N_8931,N_8509);
xor U9057 (N_9057,N_8723,N_8662);
nand U9058 (N_9058,N_8857,N_8991);
nor U9059 (N_9059,N_8702,N_8884);
or U9060 (N_9060,N_8530,N_8851);
nor U9061 (N_9061,N_8641,N_8718);
nor U9062 (N_9062,N_8679,N_8930);
and U9063 (N_9063,N_8750,N_8600);
xor U9064 (N_9064,N_8829,N_8827);
xnor U9065 (N_9065,N_8589,N_8675);
or U9066 (N_9066,N_8751,N_8692);
xor U9067 (N_9067,N_8968,N_8992);
xnor U9068 (N_9068,N_8657,N_8982);
or U9069 (N_9069,N_8784,N_8874);
or U9070 (N_9070,N_8729,N_8578);
nor U9071 (N_9071,N_8836,N_8990);
nor U9072 (N_9072,N_8934,N_8634);
xnor U9073 (N_9073,N_8721,N_8607);
and U9074 (N_9074,N_8815,N_8867);
xnor U9075 (N_9075,N_8511,N_8545);
and U9076 (N_9076,N_8939,N_8759);
nor U9077 (N_9077,N_8908,N_8671);
or U9078 (N_9078,N_8863,N_8781);
xnor U9079 (N_9079,N_8611,N_8840);
nor U9080 (N_9080,N_8820,N_8625);
nand U9081 (N_9081,N_8739,N_8959);
nand U9082 (N_9082,N_8736,N_8631);
nor U9083 (N_9083,N_8639,N_8976);
xor U9084 (N_9084,N_8848,N_8563);
nand U9085 (N_9085,N_8915,N_8979);
nor U9086 (N_9086,N_8849,N_8685);
nor U9087 (N_9087,N_8668,N_8858);
nand U9088 (N_9088,N_8871,N_8984);
nor U9089 (N_9089,N_8933,N_8712);
and U9090 (N_9090,N_8733,N_8745);
and U9091 (N_9091,N_8988,N_8828);
nand U9092 (N_9092,N_8852,N_8541);
nand U9093 (N_9093,N_8709,N_8760);
or U9094 (N_9094,N_8888,N_8799);
nor U9095 (N_9095,N_8633,N_8521);
xnor U9096 (N_9096,N_8658,N_8552);
nand U9097 (N_9097,N_8672,N_8886);
nand U9098 (N_9098,N_8522,N_8821);
nand U9099 (N_9099,N_8728,N_8698);
or U9100 (N_9100,N_8779,N_8654);
nor U9101 (N_9101,N_8782,N_8972);
nand U9102 (N_9102,N_8706,N_8916);
nand U9103 (N_9103,N_8614,N_8843);
and U9104 (N_9104,N_8792,N_8807);
xnor U9105 (N_9105,N_8512,N_8610);
nor U9106 (N_9106,N_8978,N_8935);
and U9107 (N_9107,N_8920,N_8564);
nor U9108 (N_9108,N_8627,N_8774);
and U9109 (N_9109,N_8575,N_8878);
and U9110 (N_9110,N_8746,N_8910);
nor U9111 (N_9111,N_8550,N_8812);
or U9112 (N_9112,N_8525,N_8743);
or U9113 (N_9113,N_8553,N_8700);
or U9114 (N_9114,N_8626,N_8785);
or U9115 (N_9115,N_8532,N_8534);
and U9116 (N_9116,N_8598,N_8803);
nor U9117 (N_9117,N_8789,N_8649);
nor U9118 (N_9118,N_8981,N_8638);
or U9119 (N_9119,N_8621,N_8520);
and U9120 (N_9120,N_8713,N_8818);
and U9121 (N_9121,N_8885,N_8847);
nand U9122 (N_9122,N_8909,N_8921);
xnor U9123 (N_9123,N_8705,N_8513);
xor U9124 (N_9124,N_8752,N_8680);
nor U9125 (N_9125,N_8653,N_8928);
nor U9126 (N_9126,N_8595,N_8983);
nand U9127 (N_9127,N_8536,N_8875);
or U9128 (N_9128,N_8724,N_8684);
nand U9129 (N_9129,N_8943,N_8594);
xnor U9130 (N_9130,N_8632,N_8922);
and U9131 (N_9131,N_8899,N_8865);
nand U9132 (N_9132,N_8945,N_8980);
nand U9133 (N_9133,N_8516,N_8515);
nand U9134 (N_9134,N_8678,N_8997);
xnor U9135 (N_9135,N_8608,N_8659);
xor U9136 (N_9136,N_8962,N_8822);
nor U9137 (N_9137,N_8808,N_8566);
or U9138 (N_9138,N_8652,N_8593);
or U9139 (N_9139,N_8686,N_8581);
and U9140 (N_9140,N_8616,N_8629);
xnor U9141 (N_9141,N_8576,N_8583);
xor U9142 (N_9142,N_8956,N_8648);
nor U9143 (N_9143,N_8628,N_8507);
nor U9144 (N_9144,N_8538,N_8565);
and U9145 (N_9145,N_8985,N_8526);
and U9146 (N_9146,N_8879,N_8660);
nand U9147 (N_9147,N_8584,N_8674);
and U9148 (N_9148,N_8805,N_8954);
nor U9149 (N_9149,N_8517,N_8994);
xor U9150 (N_9150,N_8973,N_8906);
nor U9151 (N_9151,N_8842,N_8612);
nor U9152 (N_9152,N_8655,N_8717);
and U9153 (N_9153,N_8740,N_8529);
nor U9154 (N_9154,N_8949,N_8894);
nor U9155 (N_9155,N_8602,N_8716);
or U9156 (N_9156,N_8619,N_8897);
nand U9157 (N_9157,N_8681,N_8866);
nor U9158 (N_9158,N_8868,N_8986);
or U9159 (N_9159,N_8797,N_8669);
or U9160 (N_9160,N_8787,N_8542);
or U9161 (N_9161,N_8960,N_8788);
nor U9162 (N_9162,N_8528,N_8762);
and U9163 (N_9163,N_8941,N_8533);
nand U9164 (N_9164,N_8763,N_8993);
nor U9165 (N_9165,N_8557,N_8798);
and U9166 (N_9166,N_8925,N_8800);
and U9167 (N_9167,N_8775,N_8747);
or U9168 (N_9168,N_8597,N_8757);
and U9169 (N_9169,N_8996,N_8592);
xor U9170 (N_9170,N_8543,N_8708);
and U9171 (N_9171,N_8816,N_8531);
xor U9172 (N_9172,N_8719,N_8549);
or U9173 (N_9173,N_8644,N_8703);
xor U9174 (N_9174,N_8519,N_8720);
and U9175 (N_9175,N_8673,N_8715);
or U9176 (N_9176,N_8891,N_8802);
xnor U9177 (N_9177,N_8710,N_8650);
xnor U9178 (N_9178,N_8854,N_8806);
nand U9179 (N_9179,N_8824,N_8546);
xor U9180 (N_9180,N_8630,N_8510);
and U9181 (N_9181,N_8560,N_8846);
nor U9182 (N_9182,N_8971,N_8501);
xnor U9183 (N_9183,N_8599,N_8790);
or U9184 (N_9184,N_8975,N_8554);
nor U9185 (N_9185,N_8590,N_8577);
nand U9186 (N_9186,N_8735,N_8677);
xnor U9187 (N_9187,N_8845,N_8753);
nand U9188 (N_9188,N_8837,N_8572);
nand U9189 (N_9189,N_8551,N_8605);
xnor U9190 (N_9190,N_8936,N_8555);
nor U9191 (N_9191,N_8514,N_8877);
or U9192 (N_9192,N_8714,N_8647);
and U9193 (N_9193,N_8889,N_8832);
and U9194 (N_9194,N_8707,N_8927);
or U9195 (N_9195,N_8688,N_8838);
xor U9196 (N_9196,N_8571,N_8817);
or U9197 (N_9197,N_8615,N_8937);
and U9198 (N_9198,N_8547,N_8693);
nor U9199 (N_9199,N_8665,N_8892);
and U9200 (N_9200,N_8995,N_8813);
xor U9201 (N_9201,N_8903,N_8502);
nor U9202 (N_9202,N_8952,N_8645);
xnor U9203 (N_9203,N_8953,N_8786);
or U9204 (N_9204,N_8958,N_8793);
nor U9205 (N_9205,N_8567,N_8651);
xnor U9206 (N_9206,N_8523,N_8642);
or U9207 (N_9207,N_8727,N_8691);
nand U9208 (N_9208,N_8814,N_8722);
nand U9209 (N_9209,N_8918,N_8901);
xor U9210 (N_9210,N_8636,N_8791);
xor U9211 (N_9211,N_8944,N_8754);
and U9212 (N_9212,N_8744,N_8844);
nand U9213 (N_9213,N_8841,N_8689);
nand U9214 (N_9214,N_8923,N_8732);
xor U9215 (N_9215,N_8963,N_8643);
xnor U9216 (N_9216,N_8881,N_8503);
nor U9217 (N_9217,N_8687,N_8859);
or U9218 (N_9218,N_8880,N_8570);
or U9219 (N_9219,N_8768,N_8825);
and U9220 (N_9220,N_8756,N_8749);
or U9221 (N_9221,N_8504,N_8617);
nand U9222 (N_9222,N_8569,N_8618);
and U9223 (N_9223,N_8853,N_8987);
xnor U9224 (N_9224,N_8609,N_8942);
and U9225 (N_9225,N_8778,N_8500);
nor U9226 (N_9226,N_8900,N_8890);
xor U9227 (N_9227,N_8696,N_8839);
nand U9228 (N_9228,N_8535,N_8767);
xnor U9229 (N_9229,N_8917,N_8924);
xor U9230 (N_9230,N_8883,N_8695);
nor U9231 (N_9231,N_8670,N_8974);
nor U9232 (N_9232,N_8965,N_8656);
or U9233 (N_9233,N_8895,N_8604);
or U9234 (N_9234,N_8755,N_8758);
nand U9235 (N_9235,N_8919,N_8731);
nand U9236 (N_9236,N_8826,N_8601);
and U9237 (N_9237,N_8664,N_8730);
xor U9238 (N_9238,N_8893,N_8860);
nand U9239 (N_9239,N_8977,N_8770);
nand U9240 (N_9240,N_8864,N_8896);
nor U9241 (N_9241,N_8969,N_8966);
and U9242 (N_9242,N_8586,N_8999);
nand U9243 (N_9243,N_8830,N_8783);
xor U9244 (N_9244,N_8970,N_8580);
nor U9245 (N_9245,N_8613,N_8622);
nand U9246 (N_9246,N_8780,N_8835);
nand U9247 (N_9247,N_8623,N_8887);
and U9248 (N_9248,N_8771,N_8855);
nor U9249 (N_9249,N_8850,N_8748);
nand U9250 (N_9250,N_8534,N_8850);
xor U9251 (N_9251,N_8879,N_8621);
or U9252 (N_9252,N_8741,N_8825);
or U9253 (N_9253,N_8511,N_8565);
nand U9254 (N_9254,N_8667,N_8640);
or U9255 (N_9255,N_8749,N_8689);
nand U9256 (N_9256,N_8683,N_8798);
or U9257 (N_9257,N_8932,N_8563);
and U9258 (N_9258,N_8635,N_8517);
or U9259 (N_9259,N_8552,N_8604);
and U9260 (N_9260,N_8977,N_8991);
or U9261 (N_9261,N_8891,N_8716);
nand U9262 (N_9262,N_8797,N_8926);
nand U9263 (N_9263,N_8871,N_8769);
or U9264 (N_9264,N_8657,N_8511);
nor U9265 (N_9265,N_8725,N_8978);
or U9266 (N_9266,N_8647,N_8513);
nor U9267 (N_9267,N_8617,N_8879);
nor U9268 (N_9268,N_8659,N_8607);
nor U9269 (N_9269,N_8897,N_8658);
nor U9270 (N_9270,N_8760,N_8671);
nand U9271 (N_9271,N_8937,N_8967);
nor U9272 (N_9272,N_8780,N_8689);
xor U9273 (N_9273,N_8978,N_8762);
xnor U9274 (N_9274,N_8876,N_8624);
or U9275 (N_9275,N_8553,N_8934);
and U9276 (N_9276,N_8568,N_8987);
and U9277 (N_9277,N_8798,N_8757);
nand U9278 (N_9278,N_8757,N_8756);
xor U9279 (N_9279,N_8938,N_8871);
xnor U9280 (N_9280,N_8524,N_8622);
nand U9281 (N_9281,N_8509,N_8526);
or U9282 (N_9282,N_8699,N_8961);
xor U9283 (N_9283,N_8729,N_8704);
nor U9284 (N_9284,N_8956,N_8946);
nand U9285 (N_9285,N_8919,N_8839);
and U9286 (N_9286,N_8655,N_8801);
or U9287 (N_9287,N_8586,N_8849);
or U9288 (N_9288,N_8953,N_8655);
nor U9289 (N_9289,N_8833,N_8979);
nor U9290 (N_9290,N_8807,N_8905);
xor U9291 (N_9291,N_8592,N_8624);
nand U9292 (N_9292,N_8953,N_8751);
and U9293 (N_9293,N_8707,N_8710);
nand U9294 (N_9294,N_8860,N_8773);
or U9295 (N_9295,N_8543,N_8789);
nor U9296 (N_9296,N_8662,N_8994);
nand U9297 (N_9297,N_8580,N_8798);
or U9298 (N_9298,N_8713,N_8872);
xor U9299 (N_9299,N_8715,N_8869);
nand U9300 (N_9300,N_8969,N_8853);
xnor U9301 (N_9301,N_8933,N_8819);
nor U9302 (N_9302,N_8874,N_8665);
nor U9303 (N_9303,N_8795,N_8953);
nand U9304 (N_9304,N_8915,N_8632);
and U9305 (N_9305,N_8678,N_8707);
xnor U9306 (N_9306,N_8760,N_8643);
nor U9307 (N_9307,N_8509,N_8891);
nor U9308 (N_9308,N_8506,N_8820);
or U9309 (N_9309,N_8698,N_8963);
and U9310 (N_9310,N_8906,N_8705);
or U9311 (N_9311,N_8814,N_8871);
nand U9312 (N_9312,N_8985,N_8704);
or U9313 (N_9313,N_8560,N_8555);
or U9314 (N_9314,N_8822,N_8598);
or U9315 (N_9315,N_8693,N_8935);
nor U9316 (N_9316,N_8604,N_8559);
nor U9317 (N_9317,N_8859,N_8662);
and U9318 (N_9318,N_8802,N_8680);
nand U9319 (N_9319,N_8819,N_8525);
and U9320 (N_9320,N_8997,N_8623);
nor U9321 (N_9321,N_8648,N_8963);
or U9322 (N_9322,N_8518,N_8854);
or U9323 (N_9323,N_8959,N_8547);
xor U9324 (N_9324,N_8788,N_8920);
or U9325 (N_9325,N_8529,N_8631);
nor U9326 (N_9326,N_8628,N_8843);
nor U9327 (N_9327,N_8630,N_8691);
xor U9328 (N_9328,N_8634,N_8548);
nor U9329 (N_9329,N_8871,N_8915);
and U9330 (N_9330,N_8937,N_8906);
or U9331 (N_9331,N_8846,N_8674);
xnor U9332 (N_9332,N_8995,N_8598);
nand U9333 (N_9333,N_8952,N_8971);
nand U9334 (N_9334,N_8965,N_8672);
xnor U9335 (N_9335,N_8746,N_8879);
nor U9336 (N_9336,N_8916,N_8728);
and U9337 (N_9337,N_8829,N_8980);
or U9338 (N_9338,N_8933,N_8716);
xnor U9339 (N_9339,N_8756,N_8907);
nor U9340 (N_9340,N_8778,N_8927);
nor U9341 (N_9341,N_8726,N_8990);
nor U9342 (N_9342,N_8947,N_8501);
and U9343 (N_9343,N_8978,N_8556);
or U9344 (N_9344,N_8905,N_8684);
nor U9345 (N_9345,N_8519,N_8557);
xnor U9346 (N_9346,N_8739,N_8902);
nor U9347 (N_9347,N_8878,N_8768);
xor U9348 (N_9348,N_8599,N_8516);
xnor U9349 (N_9349,N_8577,N_8847);
xnor U9350 (N_9350,N_8798,N_8887);
or U9351 (N_9351,N_8878,N_8617);
and U9352 (N_9352,N_8736,N_8560);
xor U9353 (N_9353,N_8740,N_8799);
and U9354 (N_9354,N_8572,N_8505);
nand U9355 (N_9355,N_8606,N_8517);
xor U9356 (N_9356,N_8737,N_8989);
nor U9357 (N_9357,N_8654,N_8757);
and U9358 (N_9358,N_8690,N_8843);
nor U9359 (N_9359,N_8749,N_8591);
and U9360 (N_9360,N_8829,N_8614);
nand U9361 (N_9361,N_8915,N_8734);
nor U9362 (N_9362,N_8845,N_8514);
xnor U9363 (N_9363,N_8605,N_8533);
nand U9364 (N_9364,N_8796,N_8895);
or U9365 (N_9365,N_8719,N_8500);
nand U9366 (N_9366,N_8689,N_8531);
xor U9367 (N_9367,N_8977,N_8946);
nand U9368 (N_9368,N_8561,N_8980);
nor U9369 (N_9369,N_8604,N_8692);
nand U9370 (N_9370,N_8574,N_8518);
nor U9371 (N_9371,N_8727,N_8546);
nor U9372 (N_9372,N_8625,N_8504);
nand U9373 (N_9373,N_8591,N_8899);
or U9374 (N_9374,N_8780,N_8828);
nand U9375 (N_9375,N_8726,N_8659);
xor U9376 (N_9376,N_8911,N_8883);
and U9377 (N_9377,N_8724,N_8548);
nand U9378 (N_9378,N_8568,N_8531);
nand U9379 (N_9379,N_8621,N_8791);
and U9380 (N_9380,N_8961,N_8634);
xor U9381 (N_9381,N_8674,N_8992);
nor U9382 (N_9382,N_8947,N_8586);
nand U9383 (N_9383,N_8654,N_8813);
nand U9384 (N_9384,N_8744,N_8505);
and U9385 (N_9385,N_8864,N_8738);
or U9386 (N_9386,N_8506,N_8575);
nand U9387 (N_9387,N_8896,N_8995);
nand U9388 (N_9388,N_8770,N_8718);
xor U9389 (N_9389,N_8519,N_8781);
and U9390 (N_9390,N_8913,N_8895);
nand U9391 (N_9391,N_8999,N_8501);
or U9392 (N_9392,N_8671,N_8998);
nand U9393 (N_9393,N_8886,N_8949);
and U9394 (N_9394,N_8521,N_8789);
or U9395 (N_9395,N_8938,N_8892);
xnor U9396 (N_9396,N_8939,N_8805);
xnor U9397 (N_9397,N_8500,N_8604);
nor U9398 (N_9398,N_8678,N_8806);
nand U9399 (N_9399,N_8788,N_8554);
nand U9400 (N_9400,N_8864,N_8616);
xnor U9401 (N_9401,N_8848,N_8512);
xor U9402 (N_9402,N_8657,N_8927);
nor U9403 (N_9403,N_8560,N_8896);
or U9404 (N_9404,N_8832,N_8903);
xor U9405 (N_9405,N_8834,N_8706);
and U9406 (N_9406,N_8922,N_8659);
and U9407 (N_9407,N_8521,N_8716);
nor U9408 (N_9408,N_8609,N_8895);
nor U9409 (N_9409,N_8717,N_8657);
or U9410 (N_9410,N_8705,N_8700);
nor U9411 (N_9411,N_8748,N_8756);
xor U9412 (N_9412,N_8812,N_8678);
nor U9413 (N_9413,N_8950,N_8685);
and U9414 (N_9414,N_8592,N_8533);
nor U9415 (N_9415,N_8874,N_8663);
nand U9416 (N_9416,N_8542,N_8804);
or U9417 (N_9417,N_8829,N_8580);
or U9418 (N_9418,N_8543,N_8688);
and U9419 (N_9419,N_8930,N_8835);
and U9420 (N_9420,N_8925,N_8547);
nor U9421 (N_9421,N_8738,N_8638);
nand U9422 (N_9422,N_8662,N_8560);
nand U9423 (N_9423,N_8503,N_8575);
or U9424 (N_9424,N_8635,N_8841);
or U9425 (N_9425,N_8931,N_8513);
and U9426 (N_9426,N_8792,N_8564);
nand U9427 (N_9427,N_8868,N_8651);
and U9428 (N_9428,N_8593,N_8949);
nand U9429 (N_9429,N_8886,N_8780);
or U9430 (N_9430,N_8807,N_8877);
nor U9431 (N_9431,N_8956,N_8921);
nor U9432 (N_9432,N_8745,N_8868);
and U9433 (N_9433,N_8911,N_8724);
nand U9434 (N_9434,N_8764,N_8875);
xor U9435 (N_9435,N_8974,N_8814);
and U9436 (N_9436,N_8855,N_8680);
xor U9437 (N_9437,N_8766,N_8818);
nand U9438 (N_9438,N_8738,N_8811);
xor U9439 (N_9439,N_8554,N_8515);
xnor U9440 (N_9440,N_8601,N_8587);
and U9441 (N_9441,N_8584,N_8529);
or U9442 (N_9442,N_8998,N_8714);
nand U9443 (N_9443,N_8782,N_8845);
nand U9444 (N_9444,N_8941,N_8823);
and U9445 (N_9445,N_8559,N_8840);
nor U9446 (N_9446,N_8781,N_8846);
or U9447 (N_9447,N_8649,N_8926);
nand U9448 (N_9448,N_8671,N_8698);
nand U9449 (N_9449,N_8941,N_8798);
and U9450 (N_9450,N_8828,N_8648);
or U9451 (N_9451,N_8531,N_8801);
and U9452 (N_9452,N_8852,N_8874);
and U9453 (N_9453,N_8551,N_8873);
nand U9454 (N_9454,N_8732,N_8882);
nor U9455 (N_9455,N_8507,N_8898);
and U9456 (N_9456,N_8992,N_8908);
xor U9457 (N_9457,N_8534,N_8546);
nor U9458 (N_9458,N_8650,N_8706);
or U9459 (N_9459,N_8927,N_8774);
xor U9460 (N_9460,N_8513,N_8782);
or U9461 (N_9461,N_8651,N_8855);
nor U9462 (N_9462,N_8585,N_8957);
xor U9463 (N_9463,N_8931,N_8551);
and U9464 (N_9464,N_8932,N_8904);
or U9465 (N_9465,N_8720,N_8948);
xnor U9466 (N_9466,N_8730,N_8620);
or U9467 (N_9467,N_8746,N_8504);
and U9468 (N_9468,N_8710,N_8785);
nor U9469 (N_9469,N_8530,N_8933);
and U9470 (N_9470,N_8945,N_8860);
or U9471 (N_9471,N_8867,N_8642);
nand U9472 (N_9472,N_8787,N_8753);
xor U9473 (N_9473,N_8705,N_8927);
or U9474 (N_9474,N_8823,N_8668);
nor U9475 (N_9475,N_8856,N_8600);
and U9476 (N_9476,N_8971,N_8566);
xor U9477 (N_9477,N_8690,N_8501);
or U9478 (N_9478,N_8661,N_8883);
xor U9479 (N_9479,N_8645,N_8624);
and U9480 (N_9480,N_8746,N_8968);
nor U9481 (N_9481,N_8840,N_8875);
and U9482 (N_9482,N_8991,N_8552);
nand U9483 (N_9483,N_8747,N_8973);
and U9484 (N_9484,N_8681,N_8532);
nand U9485 (N_9485,N_8715,N_8798);
nand U9486 (N_9486,N_8928,N_8616);
and U9487 (N_9487,N_8570,N_8518);
or U9488 (N_9488,N_8598,N_8657);
and U9489 (N_9489,N_8886,N_8658);
and U9490 (N_9490,N_8987,N_8644);
nand U9491 (N_9491,N_8917,N_8565);
or U9492 (N_9492,N_8781,N_8721);
nand U9493 (N_9493,N_8735,N_8707);
or U9494 (N_9494,N_8574,N_8779);
xor U9495 (N_9495,N_8969,N_8736);
nor U9496 (N_9496,N_8526,N_8945);
or U9497 (N_9497,N_8626,N_8849);
nor U9498 (N_9498,N_8912,N_8841);
nor U9499 (N_9499,N_8924,N_8608);
nand U9500 (N_9500,N_9403,N_9048);
or U9501 (N_9501,N_9233,N_9429);
or U9502 (N_9502,N_9019,N_9176);
nor U9503 (N_9503,N_9236,N_9266);
and U9504 (N_9504,N_9410,N_9439);
or U9505 (N_9505,N_9270,N_9042);
nand U9506 (N_9506,N_9199,N_9011);
nand U9507 (N_9507,N_9254,N_9095);
nor U9508 (N_9508,N_9475,N_9278);
xnor U9509 (N_9509,N_9044,N_9295);
and U9510 (N_9510,N_9096,N_9417);
or U9511 (N_9511,N_9074,N_9099);
xor U9512 (N_9512,N_9306,N_9238);
xor U9513 (N_9513,N_9210,N_9000);
nor U9514 (N_9514,N_9024,N_9496);
nand U9515 (N_9515,N_9376,N_9373);
nand U9516 (N_9516,N_9068,N_9018);
xnor U9517 (N_9517,N_9331,N_9123);
nand U9518 (N_9518,N_9089,N_9262);
or U9519 (N_9519,N_9397,N_9250);
nor U9520 (N_9520,N_9005,N_9126);
nor U9521 (N_9521,N_9460,N_9457);
nand U9522 (N_9522,N_9235,N_9259);
or U9523 (N_9523,N_9052,N_9327);
nor U9524 (N_9524,N_9418,N_9187);
or U9525 (N_9525,N_9047,N_9401);
nor U9526 (N_9526,N_9161,N_9225);
and U9527 (N_9527,N_9001,N_9043);
nor U9528 (N_9528,N_9487,N_9413);
nor U9529 (N_9529,N_9125,N_9078);
nand U9530 (N_9530,N_9166,N_9049);
nor U9531 (N_9531,N_9313,N_9408);
or U9532 (N_9532,N_9300,N_9114);
and U9533 (N_9533,N_9085,N_9175);
nor U9534 (N_9534,N_9389,N_9084);
nand U9535 (N_9535,N_9255,N_9363);
nor U9536 (N_9536,N_9347,N_9423);
nand U9537 (N_9537,N_9207,N_9360);
xor U9538 (N_9538,N_9190,N_9141);
nand U9539 (N_9539,N_9346,N_9385);
or U9540 (N_9540,N_9356,N_9222);
xnor U9541 (N_9541,N_9230,N_9058);
and U9542 (N_9542,N_9063,N_9107);
xor U9543 (N_9543,N_9234,N_9372);
nand U9544 (N_9544,N_9223,N_9243);
nand U9545 (N_9545,N_9139,N_9458);
or U9546 (N_9546,N_9064,N_9265);
xnor U9547 (N_9547,N_9100,N_9104);
and U9548 (N_9548,N_9159,N_9289);
or U9549 (N_9549,N_9328,N_9402);
nor U9550 (N_9550,N_9424,N_9076);
nand U9551 (N_9551,N_9256,N_9459);
nand U9552 (N_9552,N_9248,N_9163);
xor U9553 (N_9553,N_9033,N_9274);
and U9554 (N_9554,N_9038,N_9209);
nand U9555 (N_9555,N_9465,N_9387);
and U9556 (N_9556,N_9381,N_9312);
or U9557 (N_9557,N_9258,N_9196);
nand U9558 (N_9558,N_9368,N_9462);
or U9559 (N_9559,N_9437,N_9013);
or U9560 (N_9560,N_9362,N_9276);
nand U9561 (N_9561,N_9473,N_9415);
nand U9562 (N_9562,N_9152,N_9399);
or U9563 (N_9563,N_9380,N_9030);
nand U9564 (N_9564,N_9169,N_9307);
and U9565 (N_9565,N_9371,N_9212);
nand U9566 (N_9566,N_9110,N_9446);
xnor U9567 (N_9567,N_9111,N_9349);
or U9568 (N_9568,N_9338,N_9020);
or U9569 (N_9569,N_9133,N_9476);
xor U9570 (N_9570,N_9390,N_9037);
or U9571 (N_9571,N_9370,N_9193);
xor U9572 (N_9572,N_9442,N_9291);
nor U9573 (N_9573,N_9260,N_9173);
nand U9574 (N_9574,N_9318,N_9112);
or U9575 (N_9575,N_9392,N_9155);
xnor U9576 (N_9576,N_9298,N_9066);
or U9577 (N_9577,N_9148,N_9286);
nor U9578 (N_9578,N_9438,N_9321);
nand U9579 (N_9579,N_9051,N_9131);
xnor U9580 (N_9580,N_9119,N_9087);
xnor U9581 (N_9581,N_9065,N_9178);
xnor U9582 (N_9582,N_9361,N_9201);
nor U9583 (N_9583,N_9088,N_9061);
and U9584 (N_9584,N_9070,N_9191);
xnor U9585 (N_9585,N_9471,N_9086);
or U9586 (N_9586,N_9309,N_9140);
nor U9587 (N_9587,N_9264,N_9241);
or U9588 (N_9588,N_9434,N_9105);
or U9589 (N_9589,N_9228,N_9172);
and U9590 (N_9590,N_9009,N_9326);
nand U9591 (N_9591,N_9257,N_9145);
nand U9592 (N_9592,N_9028,N_9488);
or U9593 (N_9593,N_9467,N_9080);
xnor U9594 (N_9594,N_9345,N_9333);
or U9595 (N_9595,N_9211,N_9025);
and U9596 (N_9596,N_9484,N_9367);
or U9597 (N_9597,N_9229,N_9146);
and U9598 (N_9598,N_9232,N_9436);
or U9599 (N_9599,N_9184,N_9366);
or U9600 (N_9600,N_9046,N_9185);
xor U9601 (N_9601,N_9409,N_9269);
or U9602 (N_9602,N_9314,N_9040);
nand U9603 (N_9603,N_9287,N_9205);
nor U9604 (N_9604,N_9012,N_9383);
or U9605 (N_9605,N_9217,N_9422);
nand U9606 (N_9606,N_9456,N_9128);
nand U9607 (N_9607,N_9451,N_9281);
nor U9608 (N_9608,N_9004,N_9292);
or U9609 (N_9609,N_9160,N_9369);
and U9610 (N_9610,N_9015,N_9059);
and U9611 (N_9611,N_9454,N_9151);
or U9612 (N_9612,N_9108,N_9214);
and U9613 (N_9613,N_9053,N_9393);
and U9614 (N_9614,N_9034,N_9027);
nor U9615 (N_9615,N_9341,N_9204);
xor U9616 (N_9616,N_9419,N_9029);
or U9617 (N_9617,N_9157,N_9247);
nor U9618 (N_9618,N_9103,N_9072);
nor U9619 (N_9619,N_9090,N_9147);
xnor U9620 (N_9620,N_9272,N_9219);
xnor U9621 (N_9621,N_9261,N_9036);
xor U9622 (N_9622,N_9116,N_9472);
nor U9623 (N_9623,N_9069,N_9365);
nand U9624 (N_9624,N_9448,N_9299);
xnor U9625 (N_9625,N_9358,N_9468);
and U9626 (N_9626,N_9240,N_9337);
or U9627 (N_9627,N_9153,N_9324);
and U9628 (N_9628,N_9138,N_9073);
xor U9629 (N_9629,N_9246,N_9118);
or U9630 (N_9630,N_9055,N_9224);
and U9631 (N_9631,N_9433,N_9490);
xor U9632 (N_9632,N_9197,N_9310);
and U9633 (N_9633,N_9395,N_9407);
or U9634 (N_9634,N_9057,N_9198);
xnor U9635 (N_9635,N_9329,N_9242);
xnor U9636 (N_9636,N_9032,N_9091);
and U9637 (N_9637,N_9093,N_9041);
or U9638 (N_9638,N_9227,N_9267);
and U9639 (N_9639,N_9271,N_9453);
or U9640 (N_9640,N_9297,N_9106);
nand U9641 (N_9641,N_9440,N_9355);
xor U9642 (N_9642,N_9294,N_9497);
nor U9643 (N_9643,N_9293,N_9174);
and U9644 (N_9644,N_9102,N_9412);
nor U9645 (N_9645,N_9282,N_9277);
nand U9646 (N_9646,N_9213,N_9319);
nor U9647 (N_9647,N_9014,N_9315);
nor U9648 (N_9648,N_9189,N_9474);
or U9649 (N_9649,N_9249,N_9351);
nor U9650 (N_9650,N_9135,N_9251);
xor U9651 (N_9651,N_9498,N_9283);
or U9652 (N_9652,N_9268,N_9092);
xnor U9653 (N_9653,N_9461,N_9301);
or U9654 (N_9654,N_9342,N_9098);
nand U9655 (N_9655,N_9316,N_9192);
or U9656 (N_9656,N_9414,N_9122);
and U9657 (N_9657,N_9317,N_9127);
or U9658 (N_9658,N_9144,N_9186);
xor U9659 (N_9659,N_9023,N_9167);
or U9660 (N_9660,N_9124,N_9343);
and U9661 (N_9661,N_9352,N_9182);
and U9662 (N_9662,N_9404,N_9374);
xor U9663 (N_9663,N_9480,N_9206);
or U9664 (N_9664,N_9377,N_9179);
nor U9665 (N_9665,N_9117,N_9405);
nand U9666 (N_9666,N_9335,N_9428);
nand U9667 (N_9667,N_9320,N_9493);
xor U9668 (N_9668,N_9334,N_9447);
xor U9669 (N_9669,N_9109,N_9003);
and U9670 (N_9670,N_9452,N_9177);
or U9671 (N_9671,N_9411,N_9077);
nor U9672 (N_9672,N_9168,N_9008);
and U9673 (N_9673,N_9290,N_9245);
xor U9674 (N_9674,N_9220,N_9071);
nor U9675 (N_9675,N_9466,N_9181);
xor U9676 (N_9676,N_9379,N_9489);
and U9677 (N_9677,N_9455,N_9007);
and U9678 (N_9678,N_9406,N_9056);
and U9679 (N_9679,N_9464,N_9171);
xnor U9680 (N_9680,N_9162,N_9323);
nor U9681 (N_9681,N_9026,N_9304);
and U9682 (N_9682,N_9378,N_9142);
xor U9683 (N_9683,N_9398,N_9216);
or U9684 (N_9684,N_9021,N_9357);
xnor U9685 (N_9685,N_9325,N_9344);
nand U9686 (N_9686,N_9280,N_9285);
and U9687 (N_9687,N_9425,N_9330);
or U9688 (N_9688,N_9400,N_9477);
nor U9689 (N_9689,N_9444,N_9195);
xor U9690 (N_9690,N_9031,N_9083);
or U9691 (N_9691,N_9253,N_9483);
nand U9692 (N_9692,N_9010,N_9132);
xnor U9693 (N_9693,N_9188,N_9002);
xor U9694 (N_9694,N_9156,N_9226);
nor U9695 (N_9695,N_9113,N_9200);
xnor U9696 (N_9696,N_9396,N_9391);
xnor U9697 (N_9697,N_9482,N_9486);
and U9698 (N_9698,N_9420,N_9339);
or U9699 (N_9699,N_9495,N_9311);
xnor U9700 (N_9700,N_9441,N_9129);
nand U9701 (N_9701,N_9039,N_9165);
and U9702 (N_9702,N_9237,N_9231);
xor U9703 (N_9703,N_9499,N_9354);
and U9704 (N_9704,N_9180,N_9359);
or U9705 (N_9705,N_9308,N_9121);
or U9706 (N_9706,N_9094,N_9244);
nand U9707 (N_9707,N_9134,N_9375);
or U9708 (N_9708,N_9252,N_9394);
xnor U9709 (N_9709,N_9202,N_9426);
nand U9710 (N_9710,N_9485,N_9340);
and U9711 (N_9711,N_9443,N_9494);
nand U9712 (N_9712,N_9445,N_9416);
xor U9713 (N_9713,N_9164,N_9491);
or U9714 (N_9714,N_9364,N_9353);
or U9715 (N_9715,N_9062,N_9275);
nand U9716 (N_9716,N_9075,N_9203);
nor U9717 (N_9717,N_9421,N_9045);
nand U9718 (N_9718,N_9382,N_9470);
and U9719 (N_9719,N_9183,N_9081);
nor U9720 (N_9720,N_9035,N_9194);
nand U9721 (N_9721,N_9430,N_9386);
nand U9722 (N_9722,N_9432,N_9022);
and U9723 (N_9723,N_9016,N_9449);
and U9724 (N_9724,N_9149,N_9279);
nor U9725 (N_9725,N_9221,N_9332);
nor U9726 (N_9726,N_9158,N_9101);
nor U9727 (N_9727,N_9067,N_9481);
or U9728 (N_9728,N_9170,N_9303);
nor U9729 (N_9729,N_9006,N_9215);
and U9730 (N_9730,N_9284,N_9154);
nand U9731 (N_9731,N_9150,N_9427);
or U9732 (N_9732,N_9435,N_9348);
and U9733 (N_9733,N_9463,N_9079);
or U9734 (N_9734,N_9336,N_9273);
xor U9735 (N_9735,N_9492,N_9479);
nor U9736 (N_9736,N_9136,N_9305);
nand U9737 (N_9737,N_9478,N_9130);
xnor U9738 (N_9738,N_9350,N_9017);
nand U9739 (N_9739,N_9082,N_9322);
nand U9740 (N_9740,N_9450,N_9120);
nor U9741 (N_9741,N_9054,N_9097);
nand U9742 (N_9742,N_9296,N_9388);
nand U9743 (N_9743,N_9431,N_9115);
xor U9744 (N_9744,N_9384,N_9208);
and U9745 (N_9745,N_9239,N_9143);
nand U9746 (N_9746,N_9288,N_9469);
xor U9747 (N_9747,N_9263,N_9137);
xnor U9748 (N_9748,N_9050,N_9218);
nand U9749 (N_9749,N_9060,N_9302);
or U9750 (N_9750,N_9057,N_9070);
and U9751 (N_9751,N_9327,N_9020);
or U9752 (N_9752,N_9454,N_9067);
or U9753 (N_9753,N_9030,N_9288);
nand U9754 (N_9754,N_9069,N_9480);
xor U9755 (N_9755,N_9126,N_9249);
nor U9756 (N_9756,N_9210,N_9139);
xnor U9757 (N_9757,N_9326,N_9353);
or U9758 (N_9758,N_9002,N_9414);
nand U9759 (N_9759,N_9263,N_9061);
or U9760 (N_9760,N_9359,N_9421);
and U9761 (N_9761,N_9176,N_9134);
nor U9762 (N_9762,N_9154,N_9429);
nor U9763 (N_9763,N_9356,N_9255);
and U9764 (N_9764,N_9343,N_9265);
and U9765 (N_9765,N_9140,N_9181);
nand U9766 (N_9766,N_9251,N_9302);
nor U9767 (N_9767,N_9335,N_9069);
nand U9768 (N_9768,N_9211,N_9109);
and U9769 (N_9769,N_9212,N_9004);
xnor U9770 (N_9770,N_9287,N_9361);
nand U9771 (N_9771,N_9113,N_9115);
nand U9772 (N_9772,N_9427,N_9379);
nand U9773 (N_9773,N_9146,N_9056);
nor U9774 (N_9774,N_9011,N_9283);
nor U9775 (N_9775,N_9407,N_9471);
nand U9776 (N_9776,N_9317,N_9214);
and U9777 (N_9777,N_9228,N_9277);
xnor U9778 (N_9778,N_9123,N_9316);
xnor U9779 (N_9779,N_9047,N_9460);
nor U9780 (N_9780,N_9339,N_9374);
nor U9781 (N_9781,N_9316,N_9169);
or U9782 (N_9782,N_9458,N_9013);
or U9783 (N_9783,N_9150,N_9013);
or U9784 (N_9784,N_9023,N_9019);
and U9785 (N_9785,N_9023,N_9132);
nand U9786 (N_9786,N_9235,N_9438);
and U9787 (N_9787,N_9305,N_9171);
nor U9788 (N_9788,N_9342,N_9463);
xnor U9789 (N_9789,N_9174,N_9391);
nor U9790 (N_9790,N_9112,N_9048);
nor U9791 (N_9791,N_9339,N_9182);
nor U9792 (N_9792,N_9278,N_9415);
xor U9793 (N_9793,N_9151,N_9061);
nand U9794 (N_9794,N_9121,N_9276);
nand U9795 (N_9795,N_9365,N_9027);
nor U9796 (N_9796,N_9316,N_9311);
nand U9797 (N_9797,N_9051,N_9270);
xnor U9798 (N_9798,N_9337,N_9078);
or U9799 (N_9799,N_9153,N_9077);
and U9800 (N_9800,N_9084,N_9285);
nand U9801 (N_9801,N_9231,N_9191);
nand U9802 (N_9802,N_9449,N_9238);
or U9803 (N_9803,N_9108,N_9391);
nand U9804 (N_9804,N_9013,N_9118);
nor U9805 (N_9805,N_9162,N_9375);
or U9806 (N_9806,N_9355,N_9258);
and U9807 (N_9807,N_9279,N_9207);
nand U9808 (N_9808,N_9274,N_9495);
xnor U9809 (N_9809,N_9273,N_9102);
or U9810 (N_9810,N_9380,N_9378);
nor U9811 (N_9811,N_9002,N_9299);
nor U9812 (N_9812,N_9240,N_9133);
nor U9813 (N_9813,N_9462,N_9189);
nand U9814 (N_9814,N_9354,N_9285);
and U9815 (N_9815,N_9376,N_9449);
xor U9816 (N_9816,N_9043,N_9497);
nand U9817 (N_9817,N_9237,N_9397);
xnor U9818 (N_9818,N_9390,N_9008);
nand U9819 (N_9819,N_9344,N_9082);
nand U9820 (N_9820,N_9265,N_9189);
or U9821 (N_9821,N_9190,N_9449);
xor U9822 (N_9822,N_9124,N_9336);
nand U9823 (N_9823,N_9454,N_9165);
or U9824 (N_9824,N_9383,N_9204);
xor U9825 (N_9825,N_9486,N_9374);
nand U9826 (N_9826,N_9493,N_9083);
nor U9827 (N_9827,N_9097,N_9233);
nor U9828 (N_9828,N_9244,N_9007);
and U9829 (N_9829,N_9402,N_9115);
xnor U9830 (N_9830,N_9367,N_9296);
nor U9831 (N_9831,N_9469,N_9077);
xnor U9832 (N_9832,N_9228,N_9403);
nand U9833 (N_9833,N_9210,N_9081);
xor U9834 (N_9834,N_9053,N_9068);
nand U9835 (N_9835,N_9047,N_9210);
nand U9836 (N_9836,N_9079,N_9242);
nor U9837 (N_9837,N_9370,N_9032);
xor U9838 (N_9838,N_9256,N_9200);
and U9839 (N_9839,N_9121,N_9224);
nor U9840 (N_9840,N_9455,N_9026);
nor U9841 (N_9841,N_9375,N_9042);
or U9842 (N_9842,N_9071,N_9394);
or U9843 (N_9843,N_9010,N_9056);
nand U9844 (N_9844,N_9226,N_9316);
or U9845 (N_9845,N_9245,N_9433);
nor U9846 (N_9846,N_9393,N_9278);
or U9847 (N_9847,N_9042,N_9061);
and U9848 (N_9848,N_9447,N_9425);
and U9849 (N_9849,N_9183,N_9127);
nor U9850 (N_9850,N_9091,N_9092);
or U9851 (N_9851,N_9249,N_9041);
xnor U9852 (N_9852,N_9314,N_9206);
nand U9853 (N_9853,N_9492,N_9487);
nand U9854 (N_9854,N_9411,N_9227);
nor U9855 (N_9855,N_9242,N_9279);
xnor U9856 (N_9856,N_9049,N_9343);
and U9857 (N_9857,N_9451,N_9020);
or U9858 (N_9858,N_9432,N_9321);
xor U9859 (N_9859,N_9127,N_9326);
and U9860 (N_9860,N_9437,N_9221);
nor U9861 (N_9861,N_9078,N_9131);
or U9862 (N_9862,N_9094,N_9025);
or U9863 (N_9863,N_9033,N_9425);
and U9864 (N_9864,N_9154,N_9004);
nor U9865 (N_9865,N_9159,N_9452);
nor U9866 (N_9866,N_9482,N_9011);
nand U9867 (N_9867,N_9416,N_9196);
nand U9868 (N_9868,N_9216,N_9383);
nand U9869 (N_9869,N_9404,N_9218);
nand U9870 (N_9870,N_9208,N_9140);
and U9871 (N_9871,N_9396,N_9489);
nand U9872 (N_9872,N_9027,N_9465);
nand U9873 (N_9873,N_9144,N_9044);
nand U9874 (N_9874,N_9017,N_9054);
nand U9875 (N_9875,N_9035,N_9089);
xnor U9876 (N_9876,N_9003,N_9086);
xnor U9877 (N_9877,N_9037,N_9328);
xnor U9878 (N_9878,N_9222,N_9371);
nor U9879 (N_9879,N_9396,N_9417);
nor U9880 (N_9880,N_9288,N_9441);
xnor U9881 (N_9881,N_9137,N_9462);
xor U9882 (N_9882,N_9282,N_9250);
and U9883 (N_9883,N_9272,N_9281);
nor U9884 (N_9884,N_9310,N_9236);
nor U9885 (N_9885,N_9090,N_9236);
nor U9886 (N_9886,N_9009,N_9384);
and U9887 (N_9887,N_9147,N_9123);
nor U9888 (N_9888,N_9236,N_9143);
xor U9889 (N_9889,N_9367,N_9132);
nand U9890 (N_9890,N_9387,N_9273);
xor U9891 (N_9891,N_9335,N_9376);
and U9892 (N_9892,N_9146,N_9029);
nor U9893 (N_9893,N_9357,N_9139);
and U9894 (N_9894,N_9037,N_9481);
and U9895 (N_9895,N_9464,N_9354);
nor U9896 (N_9896,N_9222,N_9113);
and U9897 (N_9897,N_9206,N_9186);
nand U9898 (N_9898,N_9020,N_9162);
xor U9899 (N_9899,N_9402,N_9042);
nand U9900 (N_9900,N_9390,N_9125);
or U9901 (N_9901,N_9104,N_9329);
xor U9902 (N_9902,N_9090,N_9485);
nand U9903 (N_9903,N_9396,N_9286);
nor U9904 (N_9904,N_9268,N_9048);
nand U9905 (N_9905,N_9327,N_9445);
nand U9906 (N_9906,N_9037,N_9381);
or U9907 (N_9907,N_9337,N_9242);
and U9908 (N_9908,N_9456,N_9307);
xor U9909 (N_9909,N_9015,N_9244);
and U9910 (N_9910,N_9494,N_9040);
and U9911 (N_9911,N_9187,N_9155);
xor U9912 (N_9912,N_9006,N_9412);
nand U9913 (N_9913,N_9445,N_9311);
and U9914 (N_9914,N_9206,N_9363);
and U9915 (N_9915,N_9044,N_9338);
nor U9916 (N_9916,N_9346,N_9074);
xnor U9917 (N_9917,N_9023,N_9210);
nor U9918 (N_9918,N_9398,N_9211);
nor U9919 (N_9919,N_9210,N_9373);
or U9920 (N_9920,N_9269,N_9336);
or U9921 (N_9921,N_9113,N_9359);
or U9922 (N_9922,N_9396,N_9365);
xnor U9923 (N_9923,N_9494,N_9098);
nand U9924 (N_9924,N_9111,N_9393);
nor U9925 (N_9925,N_9047,N_9330);
or U9926 (N_9926,N_9278,N_9299);
or U9927 (N_9927,N_9132,N_9127);
xor U9928 (N_9928,N_9199,N_9175);
nor U9929 (N_9929,N_9064,N_9104);
nor U9930 (N_9930,N_9046,N_9214);
or U9931 (N_9931,N_9344,N_9367);
nand U9932 (N_9932,N_9043,N_9268);
nor U9933 (N_9933,N_9430,N_9100);
or U9934 (N_9934,N_9410,N_9174);
and U9935 (N_9935,N_9207,N_9050);
nand U9936 (N_9936,N_9085,N_9463);
or U9937 (N_9937,N_9429,N_9499);
or U9938 (N_9938,N_9318,N_9478);
nor U9939 (N_9939,N_9314,N_9122);
or U9940 (N_9940,N_9074,N_9457);
nand U9941 (N_9941,N_9196,N_9205);
nor U9942 (N_9942,N_9069,N_9317);
nand U9943 (N_9943,N_9018,N_9126);
nor U9944 (N_9944,N_9236,N_9316);
and U9945 (N_9945,N_9390,N_9104);
nand U9946 (N_9946,N_9040,N_9233);
or U9947 (N_9947,N_9308,N_9439);
nor U9948 (N_9948,N_9067,N_9158);
nand U9949 (N_9949,N_9492,N_9184);
nand U9950 (N_9950,N_9023,N_9265);
and U9951 (N_9951,N_9419,N_9477);
or U9952 (N_9952,N_9268,N_9053);
nor U9953 (N_9953,N_9356,N_9384);
nor U9954 (N_9954,N_9326,N_9159);
xor U9955 (N_9955,N_9218,N_9352);
nand U9956 (N_9956,N_9208,N_9202);
nand U9957 (N_9957,N_9175,N_9388);
xor U9958 (N_9958,N_9152,N_9165);
nor U9959 (N_9959,N_9017,N_9256);
and U9960 (N_9960,N_9497,N_9136);
xnor U9961 (N_9961,N_9073,N_9128);
xor U9962 (N_9962,N_9176,N_9046);
xnor U9963 (N_9963,N_9371,N_9248);
nand U9964 (N_9964,N_9106,N_9199);
xor U9965 (N_9965,N_9138,N_9401);
xor U9966 (N_9966,N_9006,N_9005);
or U9967 (N_9967,N_9011,N_9230);
nand U9968 (N_9968,N_9449,N_9439);
nor U9969 (N_9969,N_9460,N_9402);
nand U9970 (N_9970,N_9196,N_9097);
nor U9971 (N_9971,N_9317,N_9295);
nand U9972 (N_9972,N_9243,N_9364);
xnor U9973 (N_9973,N_9127,N_9294);
xor U9974 (N_9974,N_9230,N_9294);
xor U9975 (N_9975,N_9342,N_9185);
xor U9976 (N_9976,N_9132,N_9440);
and U9977 (N_9977,N_9457,N_9490);
xnor U9978 (N_9978,N_9499,N_9134);
nand U9979 (N_9979,N_9207,N_9321);
or U9980 (N_9980,N_9090,N_9360);
xor U9981 (N_9981,N_9001,N_9058);
nor U9982 (N_9982,N_9190,N_9079);
nor U9983 (N_9983,N_9357,N_9492);
and U9984 (N_9984,N_9095,N_9363);
xor U9985 (N_9985,N_9134,N_9075);
and U9986 (N_9986,N_9267,N_9330);
and U9987 (N_9987,N_9082,N_9476);
xor U9988 (N_9988,N_9045,N_9326);
xor U9989 (N_9989,N_9012,N_9211);
xor U9990 (N_9990,N_9329,N_9177);
nor U9991 (N_9991,N_9475,N_9257);
nor U9992 (N_9992,N_9164,N_9141);
nor U9993 (N_9993,N_9406,N_9083);
or U9994 (N_9994,N_9347,N_9273);
and U9995 (N_9995,N_9461,N_9268);
or U9996 (N_9996,N_9055,N_9463);
and U9997 (N_9997,N_9178,N_9155);
or U9998 (N_9998,N_9241,N_9418);
nand U9999 (N_9999,N_9088,N_9072);
xor U10000 (N_10000,N_9776,N_9888);
nor U10001 (N_10001,N_9681,N_9691);
xnor U10002 (N_10002,N_9634,N_9794);
nand U10003 (N_10003,N_9677,N_9511);
xor U10004 (N_10004,N_9775,N_9639);
or U10005 (N_10005,N_9865,N_9756);
nand U10006 (N_10006,N_9971,N_9597);
xnor U10007 (N_10007,N_9805,N_9978);
nor U10008 (N_10008,N_9539,N_9549);
or U10009 (N_10009,N_9766,N_9771);
or U10010 (N_10010,N_9531,N_9937);
xor U10011 (N_10011,N_9813,N_9907);
and U10012 (N_10012,N_9855,N_9747);
xnor U10013 (N_10013,N_9544,N_9972);
nand U10014 (N_10014,N_9891,N_9802);
and U10015 (N_10015,N_9648,N_9583);
nand U10016 (N_10016,N_9698,N_9986);
nand U10017 (N_10017,N_9595,N_9717);
and U10018 (N_10018,N_9750,N_9574);
or U10019 (N_10019,N_9850,N_9926);
or U10020 (N_10020,N_9998,N_9719);
and U10021 (N_10021,N_9724,N_9685);
nand U10022 (N_10022,N_9633,N_9697);
or U10023 (N_10023,N_9577,N_9992);
xnor U10024 (N_10024,N_9786,N_9552);
and U10025 (N_10025,N_9751,N_9638);
xor U10026 (N_10026,N_9694,N_9692);
nand U10027 (N_10027,N_9790,N_9812);
or U10028 (N_10028,N_9836,N_9586);
xor U10029 (N_10029,N_9565,N_9592);
and U10030 (N_10030,N_9554,N_9535);
nor U10031 (N_10031,N_9791,N_9861);
and U10032 (N_10032,N_9948,N_9584);
nand U10033 (N_10033,N_9754,N_9914);
nor U10034 (N_10034,N_9875,N_9570);
nor U10035 (N_10035,N_9566,N_9752);
xor U10036 (N_10036,N_9989,N_9748);
or U10037 (N_10037,N_9927,N_9817);
nand U10038 (N_10038,N_9938,N_9506);
nand U10039 (N_10039,N_9821,N_9516);
xor U10040 (N_10040,N_9843,N_9596);
and U10041 (N_10041,N_9670,N_9830);
xnor U10042 (N_10042,N_9587,N_9886);
nor U10043 (N_10043,N_9841,N_9857);
and U10044 (N_10044,N_9848,N_9662);
or U10045 (N_10045,N_9915,N_9921);
nor U10046 (N_10046,N_9782,N_9645);
and U10047 (N_10047,N_9520,N_9933);
nor U10048 (N_10048,N_9952,N_9684);
and U10049 (N_10049,N_9962,N_9970);
xor U10050 (N_10050,N_9873,N_9551);
nand U10051 (N_10051,N_9661,N_9930);
nand U10052 (N_10052,N_9718,N_9576);
and U10053 (N_10053,N_9810,N_9897);
nand U10054 (N_10054,N_9669,N_9777);
xnor U10055 (N_10055,N_9627,N_9612);
and U10056 (N_10056,N_9616,N_9950);
or U10057 (N_10057,N_9580,N_9729);
and U10058 (N_10058,N_9735,N_9779);
and U10059 (N_10059,N_9600,N_9668);
nor U10060 (N_10060,N_9797,N_9528);
or U10061 (N_10061,N_9940,N_9715);
nor U10062 (N_10062,N_9792,N_9993);
nand U10063 (N_10063,N_9558,N_9730);
or U10064 (N_10064,N_9517,N_9975);
and U10065 (N_10065,N_9828,N_9568);
nand U10066 (N_10066,N_9780,N_9579);
xnor U10067 (N_10067,N_9740,N_9667);
or U10068 (N_10068,N_9696,N_9538);
and U10069 (N_10069,N_9679,N_9868);
nor U10070 (N_10070,N_9611,N_9949);
nand U10071 (N_10071,N_9778,N_9932);
xor U10072 (N_10072,N_9653,N_9977);
nor U10073 (N_10073,N_9723,N_9936);
or U10074 (N_10074,N_9901,N_9762);
or U10075 (N_10075,N_9641,N_9708);
xor U10076 (N_10076,N_9967,N_9659);
nand U10077 (N_10077,N_9621,N_9716);
nand U10078 (N_10078,N_9593,N_9822);
and U10079 (N_10079,N_9755,N_9683);
xor U10080 (N_10080,N_9884,N_9935);
nor U10081 (N_10081,N_9690,N_9562);
or U10082 (N_10082,N_9500,N_9877);
and U10083 (N_10083,N_9628,N_9675);
or U10084 (N_10084,N_9845,N_9655);
and U10085 (N_10085,N_9749,N_9642);
xor U10086 (N_10086,N_9705,N_9969);
and U10087 (N_10087,N_9557,N_9991);
and U10088 (N_10088,N_9687,N_9847);
xor U10089 (N_10089,N_9602,N_9573);
nor U10090 (N_10090,N_9546,N_9869);
xnor U10091 (N_10091,N_9688,N_9644);
and U10092 (N_10092,N_9745,N_9806);
xor U10093 (N_10093,N_9783,N_9793);
and U10094 (N_10094,N_9731,N_9713);
nand U10095 (N_10095,N_9686,N_9931);
and U10096 (N_10096,N_9711,N_9739);
or U10097 (N_10097,N_9827,N_9966);
xor U10098 (N_10098,N_9706,N_9519);
nand U10099 (N_10099,N_9957,N_9689);
nand U10100 (N_10100,N_9825,N_9823);
nor U10101 (N_10101,N_9656,N_9714);
and U10102 (N_10102,N_9997,N_9878);
xnor U10103 (N_10103,N_9981,N_9728);
or U10104 (N_10104,N_9742,N_9571);
or U10105 (N_10105,N_9614,N_9814);
and U10106 (N_10106,N_9879,N_9922);
and U10107 (N_10107,N_9701,N_9807);
or U10108 (N_10108,N_9693,N_9598);
or U10109 (N_10109,N_9764,N_9615);
nor U10110 (N_10110,N_9798,N_9959);
xnor U10111 (N_10111,N_9818,N_9504);
xor U10112 (N_10112,N_9856,N_9547);
xnor U10113 (N_10113,N_9533,N_9840);
or U10114 (N_10114,N_9946,N_9703);
and U10115 (N_10115,N_9550,N_9974);
xnor U10116 (N_10116,N_9965,N_9839);
xor U10117 (N_10117,N_9890,N_9833);
or U10118 (N_10118,N_9918,N_9899);
xnor U10119 (N_10119,N_9522,N_9738);
nor U10120 (N_10120,N_9800,N_9909);
and U10121 (N_10121,N_9556,N_9893);
nand U10122 (N_10122,N_9736,N_9502);
and U10123 (N_10123,N_9503,N_9976);
and U10124 (N_10124,N_9725,N_9956);
nor U10125 (N_10125,N_9673,N_9999);
nor U10126 (N_10126,N_9536,N_9955);
xor U10127 (N_10127,N_9575,N_9852);
xor U10128 (N_10128,N_9758,N_9788);
nand U10129 (N_10129,N_9934,N_9514);
xnor U10130 (N_10130,N_9760,N_9996);
xnor U10131 (N_10131,N_9529,N_9954);
nand U10132 (N_10132,N_9676,N_9892);
nand U10133 (N_10133,N_9874,N_9560);
nor U10134 (N_10134,N_9682,N_9829);
xor U10135 (N_10135,N_9590,N_9796);
and U10136 (N_10136,N_9635,N_9545);
nand U10137 (N_10137,N_9636,N_9649);
xor U10138 (N_10138,N_9647,N_9548);
or U10139 (N_10139,N_9985,N_9744);
nand U10140 (N_10140,N_9980,N_9880);
nand U10141 (N_10141,N_9815,N_9663);
xor U10142 (N_10142,N_9983,N_9911);
nor U10143 (N_10143,N_9809,N_9524);
and U10144 (N_10144,N_9942,N_9619);
and U10145 (N_10145,N_9505,N_9862);
and U10146 (N_10146,N_9664,N_9789);
nor U10147 (N_10147,N_9671,N_9808);
or U10148 (N_10148,N_9559,N_9924);
xnor U10149 (N_10149,N_9913,N_9772);
or U10150 (N_10150,N_9555,N_9678);
xnor U10151 (N_10151,N_9553,N_9526);
xor U10152 (N_10152,N_9885,N_9640);
nand U10153 (N_10153,N_9900,N_9785);
xor U10154 (N_10154,N_9801,N_9660);
nor U10155 (N_10155,N_9702,N_9943);
or U10156 (N_10156,N_9905,N_9824);
and U10157 (N_10157,N_9737,N_9844);
nand U10158 (N_10158,N_9721,N_9518);
nand U10159 (N_10159,N_9510,N_9707);
nor U10160 (N_10160,N_9581,N_9695);
nand U10161 (N_10161,N_9923,N_9819);
nand U10162 (N_10162,N_9838,N_9532);
and U10163 (N_10163,N_9629,N_9811);
xnor U10164 (N_10164,N_9854,N_9871);
and U10165 (N_10165,N_9968,N_9994);
or U10166 (N_10166,N_9525,N_9567);
nand U10167 (N_10167,N_9534,N_9889);
nor U10168 (N_10168,N_9606,N_9902);
and U10169 (N_10169,N_9607,N_9781);
and U10170 (N_10170,N_9872,N_9672);
nor U10171 (N_10171,N_9761,N_9773);
and U10172 (N_10172,N_9508,N_9853);
and U10173 (N_10173,N_9906,N_9987);
nor U10174 (N_10174,N_9515,N_9563);
or U10175 (N_10175,N_9620,N_9582);
xnor U10176 (N_10176,N_9765,N_9609);
xor U10177 (N_10177,N_9753,N_9643);
nor U10178 (N_10178,N_9700,N_9929);
and U10179 (N_10179,N_9720,N_9908);
xnor U10180 (N_10180,N_9882,N_9646);
xor U10181 (N_10181,N_9572,N_9832);
nand U10182 (N_10182,N_9658,N_9887);
and U10183 (N_10183,N_9680,N_9953);
xor U10184 (N_10184,N_9916,N_9842);
and U10185 (N_10185,N_9919,N_9608);
xnor U10186 (N_10186,N_9904,N_9804);
or U10187 (N_10187,N_9896,N_9917);
nand U10188 (N_10188,N_9637,N_9599);
xnor U10189 (N_10189,N_9757,N_9803);
nand U10190 (N_10190,N_9537,N_9864);
xor U10191 (N_10191,N_9799,N_9589);
nand U10192 (N_10192,N_9540,N_9951);
or U10193 (N_10193,N_9837,N_9939);
and U10194 (N_10194,N_9578,N_9709);
or U10195 (N_10195,N_9604,N_9973);
and U10196 (N_10196,N_9851,N_9654);
xor U10197 (N_10197,N_9944,N_9831);
xor U10198 (N_10198,N_9945,N_9866);
nor U10199 (N_10199,N_9910,N_9617);
nor U10200 (N_10200,N_9541,N_9834);
xnor U10201 (N_10201,N_9767,N_9903);
nand U10202 (N_10202,N_9501,N_9613);
nor U10203 (N_10203,N_9591,N_9603);
xnor U10204 (N_10204,N_9849,N_9770);
or U10205 (N_10205,N_9759,N_9523);
and U10206 (N_10206,N_9521,N_9623);
or U10207 (N_10207,N_9601,N_9542);
nand U10208 (N_10208,N_9704,N_9513);
and U10209 (N_10209,N_9795,N_9746);
nand U10210 (N_10210,N_9995,N_9963);
nand U10211 (N_10211,N_9727,N_9733);
or U10212 (N_10212,N_9666,N_9961);
and U10213 (N_10213,N_9988,N_9769);
or U10214 (N_10214,N_9622,N_9712);
and U10215 (N_10215,N_9763,N_9650);
nand U10216 (N_10216,N_9741,N_9990);
and U10217 (N_10217,N_9631,N_9674);
and U10218 (N_10218,N_9632,N_9816);
nand U10219 (N_10219,N_9665,N_9512);
or U10220 (N_10220,N_9585,N_9820);
nand U10221 (N_10221,N_9564,N_9870);
nor U10222 (N_10222,N_9883,N_9895);
xnor U10223 (N_10223,N_9734,N_9835);
nand U10224 (N_10224,N_9618,N_9594);
xor U10225 (N_10225,N_9624,N_9710);
or U10226 (N_10226,N_9898,N_9561);
or U10227 (N_10227,N_9826,N_9958);
and U10228 (N_10228,N_9657,N_9732);
xor U10229 (N_10229,N_9964,N_9881);
nor U10230 (N_10230,N_9859,N_9984);
nor U10231 (N_10231,N_9894,N_9588);
or U10232 (N_10232,N_9858,N_9787);
or U10233 (N_10233,N_9960,N_9630);
xor U10234 (N_10234,N_9543,N_9652);
and U10235 (N_10235,N_9610,N_9876);
or U10236 (N_10236,N_9726,N_9626);
nor U10237 (N_10237,N_9530,N_9912);
xor U10238 (N_10238,N_9860,N_9928);
nor U10239 (N_10239,N_9846,N_9784);
xnor U10240 (N_10240,N_9979,N_9920);
and U10241 (N_10241,N_9925,N_9699);
or U10242 (N_10242,N_9605,N_9941);
and U10243 (N_10243,N_9982,N_9774);
or U10244 (N_10244,N_9625,N_9507);
nand U10245 (N_10245,N_9867,N_9527);
and U10246 (N_10246,N_9743,N_9863);
nor U10247 (N_10247,N_9768,N_9722);
and U10248 (N_10248,N_9947,N_9569);
nand U10249 (N_10249,N_9651,N_9509);
nand U10250 (N_10250,N_9990,N_9539);
nor U10251 (N_10251,N_9930,N_9643);
xor U10252 (N_10252,N_9951,N_9954);
xnor U10253 (N_10253,N_9509,N_9503);
xnor U10254 (N_10254,N_9683,N_9976);
nand U10255 (N_10255,N_9748,N_9688);
and U10256 (N_10256,N_9556,N_9679);
nor U10257 (N_10257,N_9830,N_9672);
or U10258 (N_10258,N_9559,N_9500);
xnor U10259 (N_10259,N_9705,N_9521);
xor U10260 (N_10260,N_9885,N_9981);
or U10261 (N_10261,N_9891,N_9571);
xor U10262 (N_10262,N_9772,N_9976);
xor U10263 (N_10263,N_9713,N_9956);
nand U10264 (N_10264,N_9792,N_9694);
nor U10265 (N_10265,N_9980,N_9938);
xor U10266 (N_10266,N_9724,N_9719);
nor U10267 (N_10267,N_9665,N_9558);
nor U10268 (N_10268,N_9627,N_9855);
and U10269 (N_10269,N_9613,N_9904);
xor U10270 (N_10270,N_9913,N_9885);
xnor U10271 (N_10271,N_9900,N_9531);
nand U10272 (N_10272,N_9919,N_9829);
or U10273 (N_10273,N_9749,N_9697);
nand U10274 (N_10274,N_9757,N_9945);
nand U10275 (N_10275,N_9740,N_9677);
nand U10276 (N_10276,N_9657,N_9600);
xnor U10277 (N_10277,N_9711,N_9880);
xnor U10278 (N_10278,N_9724,N_9603);
nand U10279 (N_10279,N_9574,N_9709);
xnor U10280 (N_10280,N_9848,N_9607);
and U10281 (N_10281,N_9659,N_9753);
nor U10282 (N_10282,N_9814,N_9650);
nand U10283 (N_10283,N_9938,N_9822);
xnor U10284 (N_10284,N_9520,N_9685);
and U10285 (N_10285,N_9877,N_9777);
xor U10286 (N_10286,N_9636,N_9907);
xnor U10287 (N_10287,N_9827,N_9773);
xor U10288 (N_10288,N_9843,N_9893);
nand U10289 (N_10289,N_9984,N_9598);
xnor U10290 (N_10290,N_9788,N_9995);
and U10291 (N_10291,N_9900,N_9909);
or U10292 (N_10292,N_9547,N_9949);
or U10293 (N_10293,N_9871,N_9827);
and U10294 (N_10294,N_9691,N_9511);
xnor U10295 (N_10295,N_9558,N_9547);
nand U10296 (N_10296,N_9779,N_9597);
nor U10297 (N_10297,N_9611,N_9713);
and U10298 (N_10298,N_9519,N_9567);
and U10299 (N_10299,N_9532,N_9554);
or U10300 (N_10300,N_9997,N_9653);
xor U10301 (N_10301,N_9878,N_9811);
nor U10302 (N_10302,N_9764,N_9909);
or U10303 (N_10303,N_9960,N_9592);
or U10304 (N_10304,N_9736,N_9509);
or U10305 (N_10305,N_9958,N_9978);
and U10306 (N_10306,N_9722,N_9822);
or U10307 (N_10307,N_9607,N_9660);
nor U10308 (N_10308,N_9761,N_9905);
or U10309 (N_10309,N_9973,N_9877);
or U10310 (N_10310,N_9779,N_9968);
or U10311 (N_10311,N_9852,N_9506);
nor U10312 (N_10312,N_9635,N_9622);
xor U10313 (N_10313,N_9746,N_9895);
xnor U10314 (N_10314,N_9757,N_9742);
nor U10315 (N_10315,N_9642,N_9584);
xor U10316 (N_10316,N_9984,N_9804);
nand U10317 (N_10317,N_9993,N_9846);
nor U10318 (N_10318,N_9854,N_9750);
nor U10319 (N_10319,N_9893,N_9507);
nand U10320 (N_10320,N_9820,N_9741);
nand U10321 (N_10321,N_9994,N_9593);
nand U10322 (N_10322,N_9832,N_9875);
nor U10323 (N_10323,N_9605,N_9641);
and U10324 (N_10324,N_9878,N_9630);
and U10325 (N_10325,N_9584,N_9998);
nor U10326 (N_10326,N_9975,N_9573);
or U10327 (N_10327,N_9524,N_9838);
or U10328 (N_10328,N_9994,N_9611);
nor U10329 (N_10329,N_9690,N_9778);
nand U10330 (N_10330,N_9985,N_9530);
xor U10331 (N_10331,N_9919,N_9904);
nor U10332 (N_10332,N_9981,N_9919);
or U10333 (N_10333,N_9652,N_9707);
or U10334 (N_10334,N_9728,N_9558);
and U10335 (N_10335,N_9520,N_9522);
xor U10336 (N_10336,N_9874,N_9518);
xnor U10337 (N_10337,N_9523,N_9970);
and U10338 (N_10338,N_9553,N_9794);
xor U10339 (N_10339,N_9839,N_9819);
nor U10340 (N_10340,N_9809,N_9521);
or U10341 (N_10341,N_9599,N_9787);
nand U10342 (N_10342,N_9587,N_9594);
or U10343 (N_10343,N_9799,N_9507);
and U10344 (N_10344,N_9760,N_9501);
nor U10345 (N_10345,N_9923,N_9657);
or U10346 (N_10346,N_9967,N_9513);
and U10347 (N_10347,N_9840,N_9697);
and U10348 (N_10348,N_9872,N_9617);
or U10349 (N_10349,N_9670,N_9791);
nand U10350 (N_10350,N_9676,N_9635);
nor U10351 (N_10351,N_9901,N_9534);
or U10352 (N_10352,N_9823,N_9801);
nand U10353 (N_10353,N_9572,N_9776);
or U10354 (N_10354,N_9532,N_9945);
xnor U10355 (N_10355,N_9552,N_9931);
or U10356 (N_10356,N_9843,N_9751);
nor U10357 (N_10357,N_9650,N_9872);
nor U10358 (N_10358,N_9773,N_9937);
nor U10359 (N_10359,N_9842,N_9605);
nand U10360 (N_10360,N_9613,N_9873);
and U10361 (N_10361,N_9648,N_9594);
or U10362 (N_10362,N_9861,N_9866);
and U10363 (N_10363,N_9923,N_9607);
or U10364 (N_10364,N_9822,N_9561);
nor U10365 (N_10365,N_9888,N_9981);
and U10366 (N_10366,N_9686,N_9589);
nand U10367 (N_10367,N_9562,N_9760);
nand U10368 (N_10368,N_9650,N_9935);
and U10369 (N_10369,N_9522,N_9926);
nand U10370 (N_10370,N_9983,N_9727);
or U10371 (N_10371,N_9524,N_9815);
or U10372 (N_10372,N_9618,N_9617);
nand U10373 (N_10373,N_9842,N_9992);
and U10374 (N_10374,N_9916,N_9711);
nand U10375 (N_10375,N_9654,N_9568);
nor U10376 (N_10376,N_9918,N_9607);
nand U10377 (N_10377,N_9696,N_9880);
nand U10378 (N_10378,N_9723,N_9538);
and U10379 (N_10379,N_9513,N_9998);
nand U10380 (N_10380,N_9886,N_9727);
nor U10381 (N_10381,N_9797,N_9573);
and U10382 (N_10382,N_9920,N_9588);
xnor U10383 (N_10383,N_9851,N_9870);
or U10384 (N_10384,N_9877,N_9606);
and U10385 (N_10385,N_9947,N_9980);
xnor U10386 (N_10386,N_9805,N_9772);
or U10387 (N_10387,N_9891,N_9501);
or U10388 (N_10388,N_9573,N_9721);
or U10389 (N_10389,N_9628,N_9903);
nor U10390 (N_10390,N_9867,N_9755);
xor U10391 (N_10391,N_9915,N_9500);
and U10392 (N_10392,N_9696,N_9536);
xor U10393 (N_10393,N_9509,N_9947);
and U10394 (N_10394,N_9584,N_9731);
nor U10395 (N_10395,N_9604,N_9818);
nor U10396 (N_10396,N_9685,N_9810);
nand U10397 (N_10397,N_9873,N_9850);
nand U10398 (N_10398,N_9547,N_9908);
or U10399 (N_10399,N_9766,N_9970);
nor U10400 (N_10400,N_9915,N_9843);
and U10401 (N_10401,N_9531,N_9760);
or U10402 (N_10402,N_9872,N_9616);
and U10403 (N_10403,N_9856,N_9954);
or U10404 (N_10404,N_9540,N_9743);
or U10405 (N_10405,N_9962,N_9828);
and U10406 (N_10406,N_9682,N_9749);
or U10407 (N_10407,N_9549,N_9738);
nor U10408 (N_10408,N_9578,N_9548);
nor U10409 (N_10409,N_9687,N_9633);
xnor U10410 (N_10410,N_9678,N_9572);
xnor U10411 (N_10411,N_9868,N_9890);
nand U10412 (N_10412,N_9641,N_9934);
and U10413 (N_10413,N_9897,N_9818);
or U10414 (N_10414,N_9779,N_9574);
or U10415 (N_10415,N_9732,N_9694);
nand U10416 (N_10416,N_9839,N_9503);
xor U10417 (N_10417,N_9944,N_9724);
or U10418 (N_10418,N_9682,N_9571);
or U10419 (N_10419,N_9598,N_9614);
or U10420 (N_10420,N_9556,N_9569);
or U10421 (N_10421,N_9876,N_9520);
and U10422 (N_10422,N_9984,N_9579);
and U10423 (N_10423,N_9751,N_9948);
nand U10424 (N_10424,N_9551,N_9571);
xor U10425 (N_10425,N_9627,N_9941);
nand U10426 (N_10426,N_9748,N_9647);
and U10427 (N_10427,N_9754,N_9823);
or U10428 (N_10428,N_9543,N_9894);
nand U10429 (N_10429,N_9797,N_9810);
nand U10430 (N_10430,N_9795,N_9661);
nand U10431 (N_10431,N_9965,N_9760);
xor U10432 (N_10432,N_9977,N_9765);
and U10433 (N_10433,N_9857,N_9677);
and U10434 (N_10434,N_9617,N_9666);
or U10435 (N_10435,N_9568,N_9512);
xnor U10436 (N_10436,N_9757,N_9860);
xnor U10437 (N_10437,N_9928,N_9999);
nand U10438 (N_10438,N_9612,N_9950);
xor U10439 (N_10439,N_9638,N_9722);
nand U10440 (N_10440,N_9900,N_9982);
xnor U10441 (N_10441,N_9745,N_9930);
or U10442 (N_10442,N_9883,N_9550);
xnor U10443 (N_10443,N_9640,N_9628);
nand U10444 (N_10444,N_9933,N_9684);
xnor U10445 (N_10445,N_9931,N_9763);
or U10446 (N_10446,N_9840,N_9949);
and U10447 (N_10447,N_9796,N_9850);
xor U10448 (N_10448,N_9899,N_9701);
xor U10449 (N_10449,N_9514,N_9743);
nor U10450 (N_10450,N_9957,N_9663);
and U10451 (N_10451,N_9817,N_9838);
xor U10452 (N_10452,N_9901,N_9950);
or U10453 (N_10453,N_9935,N_9539);
or U10454 (N_10454,N_9887,N_9721);
or U10455 (N_10455,N_9620,N_9663);
nand U10456 (N_10456,N_9756,N_9525);
nor U10457 (N_10457,N_9653,N_9503);
nor U10458 (N_10458,N_9738,N_9728);
and U10459 (N_10459,N_9980,N_9558);
nand U10460 (N_10460,N_9920,N_9836);
and U10461 (N_10461,N_9848,N_9877);
or U10462 (N_10462,N_9794,N_9691);
and U10463 (N_10463,N_9531,N_9679);
nor U10464 (N_10464,N_9687,N_9751);
nand U10465 (N_10465,N_9997,N_9560);
nor U10466 (N_10466,N_9939,N_9649);
nand U10467 (N_10467,N_9759,N_9531);
and U10468 (N_10468,N_9547,N_9972);
xnor U10469 (N_10469,N_9585,N_9552);
nand U10470 (N_10470,N_9633,N_9503);
nor U10471 (N_10471,N_9747,N_9806);
xor U10472 (N_10472,N_9513,N_9941);
or U10473 (N_10473,N_9942,N_9783);
nand U10474 (N_10474,N_9743,N_9789);
or U10475 (N_10475,N_9890,N_9525);
nor U10476 (N_10476,N_9512,N_9507);
and U10477 (N_10477,N_9986,N_9756);
and U10478 (N_10478,N_9544,N_9899);
nor U10479 (N_10479,N_9687,N_9865);
xnor U10480 (N_10480,N_9670,N_9517);
nand U10481 (N_10481,N_9954,N_9508);
nand U10482 (N_10482,N_9564,N_9873);
nor U10483 (N_10483,N_9778,N_9734);
or U10484 (N_10484,N_9935,N_9698);
nand U10485 (N_10485,N_9677,N_9872);
nand U10486 (N_10486,N_9678,N_9625);
nand U10487 (N_10487,N_9819,N_9554);
or U10488 (N_10488,N_9692,N_9764);
nor U10489 (N_10489,N_9681,N_9596);
nor U10490 (N_10490,N_9604,N_9705);
and U10491 (N_10491,N_9909,N_9860);
nand U10492 (N_10492,N_9813,N_9919);
xnor U10493 (N_10493,N_9732,N_9787);
nor U10494 (N_10494,N_9798,N_9713);
and U10495 (N_10495,N_9623,N_9668);
or U10496 (N_10496,N_9764,N_9810);
nor U10497 (N_10497,N_9612,N_9531);
nor U10498 (N_10498,N_9542,N_9966);
xor U10499 (N_10499,N_9856,N_9665);
or U10500 (N_10500,N_10145,N_10118);
or U10501 (N_10501,N_10492,N_10263);
xor U10502 (N_10502,N_10137,N_10153);
or U10503 (N_10503,N_10243,N_10180);
nor U10504 (N_10504,N_10249,N_10406);
nand U10505 (N_10505,N_10046,N_10291);
or U10506 (N_10506,N_10156,N_10253);
and U10507 (N_10507,N_10054,N_10358);
and U10508 (N_10508,N_10272,N_10318);
nand U10509 (N_10509,N_10193,N_10251);
xor U10510 (N_10510,N_10087,N_10402);
xnor U10511 (N_10511,N_10483,N_10347);
or U10512 (N_10512,N_10383,N_10122);
and U10513 (N_10513,N_10098,N_10250);
or U10514 (N_10514,N_10474,N_10419);
and U10515 (N_10515,N_10240,N_10388);
nor U10516 (N_10516,N_10489,N_10049);
xor U10517 (N_10517,N_10469,N_10051);
or U10518 (N_10518,N_10055,N_10493);
xnor U10519 (N_10519,N_10257,N_10459);
or U10520 (N_10520,N_10177,N_10323);
or U10521 (N_10521,N_10311,N_10297);
or U10522 (N_10522,N_10136,N_10453);
nand U10523 (N_10523,N_10476,N_10024);
xnor U10524 (N_10524,N_10315,N_10305);
nor U10525 (N_10525,N_10467,N_10038);
xnor U10526 (N_10526,N_10352,N_10327);
and U10527 (N_10527,N_10096,N_10446);
and U10528 (N_10528,N_10335,N_10460);
xnor U10529 (N_10529,N_10190,N_10040);
nand U10530 (N_10530,N_10037,N_10435);
and U10531 (N_10531,N_10471,N_10449);
nand U10532 (N_10532,N_10018,N_10094);
nor U10533 (N_10533,N_10058,N_10464);
nor U10534 (N_10534,N_10083,N_10201);
and U10535 (N_10535,N_10060,N_10144);
nor U10536 (N_10536,N_10178,N_10102);
xnor U10537 (N_10537,N_10451,N_10126);
nor U10538 (N_10538,N_10142,N_10203);
xor U10539 (N_10539,N_10226,N_10407);
nand U10540 (N_10540,N_10336,N_10208);
and U10541 (N_10541,N_10248,N_10053);
nor U10542 (N_10542,N_10444,N_10260);
xnor U10543 (N_10543,N_10100,N_10025);
and U10544 (N_10544,N_10438,N_10441);
xnor U10545 (N_10545,N_10070,N_10361);
xor U10546 (N_10546,N_10287,N_10155);
or U10547 (N_10547,N_10472,N_10356);
and U10548 (N_10548,N_10484,N_10465);
nand U10549 (N_10549,N_10187,N_10062);
nor U10550 (N_10550,N_10359,N_10228);
and U10551 (N_10551,N_10017,N_10404);
nand U10552 (N_10552,N_10231,N_10061);
and U10553 (N_10553,N_10007,N_10270);
and U10554 (N_10554,N_10281,N_10277);
nand U10555 (N_10555,N_10215,N_10302);
nor U10556 (N_10556,N_10307,N_10320);
nand U10557 (N_10557,N_10052,N_10322);
xnor U10558 (N_10558,N_10285,N_10463);
nor U10559 (N_10559,N_10105,N_10171);
nand U10560 (N_10560,N_10162,N_10166);
or U10561 (N_10561,N_10282,N_10428);
nand U10562 (N_10562,N_10108,N_10115);
nand U10563 (N_10563,N_10072,N_10418);
nor U10564 (N_10564,N_10275,N_10351);
nand U10565 (N_10565,N_10232,N_10033);
or U10566 (N_10566,N_10084,N_10298);
xnor U10567 (N_10567,N_10043,N_10233);
nand U10568 (N_10568,N_10225,N_10158);
nand U10569 (N_10569,N_10019,N_10041);
nor U10570 (N_10570,N_10132,N_10110);
nand U10571 (N_10571,N_10309,N_10172);
xor U10572 (N_10572,N_10324,N_10238);
and U10573 (N_10573,N_10165,N_10290);
or U10574 (N_10574,N_10169,N_10021);
nand U10575 (N_10575,N_10164,N_10325);
or U10576 (N_10576,N_10246,N_10223);
xnor U10577 (N_10577,N_10380,N_10026);
xor U10578 (N_10578,N_10022,N_10129);
xor U10579 (N_10579,N_10434,N_10095);
and U10580 (N_10580,N_10131,N_10128);
xor U10581 (N_10581,N_10377,N_10384);
xor U10582 (N_10582,N_10280,N_10425);
xor U10583 (N_10583,N_10167,N_10374);
or U10584 (N_10584,N_10445,N_10473);
and U10585 (N_10585,N_10082,N_10152);
nand U10586 (N_10586,N_10135,N_10466);
xor U10587 (N_10587,N_10073,N_10047);
nor U10588 (N_10588,N_10191,N_10316);
xor U10589 (N_10589,N_10278,N_10048);
nor U10590 (N_10590,N_10078,N_10074);
and U10591 (N_10591,N_10068,N_10403);
or U10592 (N_10592,N_10410,N_10218);
nand U10593 (N_10593,N_10076,N_10331);
xor U10594 (N_10594,N_10161,N_10353);
xnor U10595 (N_10595,N_10216,N_10150);
xor U10596 (N_10596,N_10424,N_10371);
nor U10597 (N_10597,N_10414,N_10151);
nor U10598 (N_10598,N_10138,N_10326);
or U10599 (N_10599,N_10234,N_10330);
or U10600 (N_10600,N_10106,N_10396);
nor U10601 (N_10601,N_10420,N_10362);
or U10602 (N_10602,N_10067,N_10259);
and U10603 (N_10603,N_10057,N_10276);
or U10604 (N_10604,N_10141,N_10032);
nand U10605 (N_10605,N_10389,N_10411);
nor U10606 (N_10606,N_10455,N_10485);
nand U10607 (N_10607,N_10173,N_10394);
nor U10608 (N_10608,N_10334,N_10130);
xor U10609 (N_10609,N_10398,N_10342);
nor U10610 (N_10610,N_10273,N_10354);
and U10611 (N_10611,N_10268,N_10099);
and U10612 (N_10612,N_10440,N_10381);
xor U10613 (N_10613,N_10159,N_10056);
nor U10614 (N_10614,N_10480,N_10416);
nor U10615 (N_10615,N_10194,N_10378);
and U10616 (N_10616,N_10303,N_10097);
nor U10617 (N_10617,N_10175,N_10286);
and U10618 (N_10618,N_10478,N_10085);
nand U10619 (N_10619,N_10346,N_10014);
and U10620 (N_10620,N_10399,N_10116);
and U10621 (N_10621,N_10462,N_10321);
xnor U10622 (N_10622,N_10109,N_10317);
or U10623 (N_10623,N_10075,N_10221);
nor U10624 (N_10624,N_10202,N_10468);
nand U10625 (N_10625,N_10345,N_10265);
nor U10626 (N_10626,N_10432,N_10300);
xor U10627 (N_10627,N_10222,N_10196);
or U10628 (N_10628,N_10339,N_10192);
and U10629 (N_10629,N_10034,N_10039);
and U10630 (N_10630,N_10120,N_10429);
nand U10631 (N_10631,N_10134,N_10499);
or U10632 (N_10632,N_10496,N_10284);
nand U10633 (N_10633,N_10020,N_10266);
xor U10634 (N_10634,N_10059,N_10042);
nand U10635 (N_10635,N_10079,N_10003);
nor U10636 (N_10636,N_10123,N_10163);
nand U10637 (N_10637,N_10210,N_10168);
and U10638 (N_10638,N_10200,N_10369);
nor U10639 (N_10639,N_10479,N_10386);
nand U10640 (N_10640,N_10308,N_10413);
nand U10641 (N_10641,N_10147,N_10124);
and U10642 (N_10642,N_10036,N_10385);
nand U10643 (N_10643,N_10387,N_10241);
xor U10644 (N_10644,N_10269,N_10149);
xor U10645 (N_10645,N_10366,N_10350);
nor U10646 (N_10646,N_10490,N_10254);
nor U10647 (N_10647,N_10299,N_10401);
xor U10648 (N_10648,N_10206,N_10329);
nor U10649 (N_10649,N_10319,N_10491);
nand U10650 (N_10650,N_10015,N_10198);
xnor U10651 (N_10651,N_10224,N_10211);
xor U10652 (N_10652,N_10422,N_10008);
xor U10653 (N_10653,N_10475,N_10001);
or U10654 (N_10654,N_10392,N_10368);
nand U10655 (N_10655,N_10113,N_10365);
and U10656 (N_10656,N_10408,N_10332);
xnor U10657 (N_10657,N_10121,N_10117);
or U10658 (N_10658,N_10454,N_10101);
and U10659 (N_10659,N_10355,N_10393);
and U10660 (N_10660,N_10482,N_10439);
xnor U10661 (N_10661,N_10089,N_10065);
or U10662 (N_10662,N_10230,N_10433);
nand U10663 (N_10663,N_10288,N_10093);
xor U10664 (N_10664,N_10183,N_10029);
and U10665 (N_10665,N_10456,N_10044);
xnor U10666 (N_10666,N_10256,N_10376);
or U10667 (N_10667,N_10170,N_10397);
xor U10668 (N_10668,N_10154,N_10426);
nor U10669 (N_10669,N_10214,N_10209);
nor U10670 (N_10670,N_10009,N_10139);
nor U10671 (N_10671,N_10245,N_10066);
nand U10672 (N_10672,N_10333,N_10431);
or U10673 (N_10673,N_10005,N_10091);
or U10674 (N_10674,N_10314,N_10312);
nor U10675 (N_10675,N_10498,N_10373);
nor U10676 (N_10676,N_10304,N_10372);
nand U10677 (N_10677,N_10092,N_10111);
or U10678 (N_10678,N_10069,N_10343);
xor U10679 (N_10679,N_10002,N_10236);
or U10680 (N_10680,N_10195,N_10016);
and U10681 (N_10681,N_10458,N_10370);
nand U10682 (N_10682,N_10086,N_10035);
nor U10683 (N_10683,N_10242,N_10421);
or U10684 (N_10684,N_10495,N_10204);
nor U10685 (N_10685,N_10010,N_10104);
and U10686 (N_10686,N_10258,N_10338);
and U10687 (N_10687,N_10448,N_10450);
nand U10688 (N_10688,N_10283,N_10235);
xor U10689 (N_10689,N_10179,N_10143);
or U10690 (N_10690,N_10488,N_10427);
or U10691 (N_10691,N_10415,N_10205);
or U10692 (N_10692,N_10442,N_10148);
xnor U10693 (N_10693,N_10497,N_10340);
nand U10694 (N_10694,N_10000,N_10012);
or U10695 (N_10695,N_10379,N_10181);
nor U10696 (N_10696,N_10207,N_10364);
nand U10697 (N_10697,N_10264,N_10367);
xnor U10698 (N_10698,N_10470,N_10295);
nor U10699 (N_10699,N_10294,N_10360);
xnor U10700 (N_10700,N_10006,N_10262);
nand U10701 (N_10701,N_10247,N_10400);
nand U10702 (N_10702,N_10244,N_10296);
nand U10703 (N_10703,N_10081,N_10447);
nand U10704 (N_10704,N_10409,N_10292);
nor U10705 (N_10705,N_10313,N_10487);
or U10706 (N_10706,N_10289,N_10064);
nor U10707 (N_10707,N_10160,N_10028);
and U10708 (N_10708,N_10395,N_10213);
nand U10709 (N_10709,N_10185,N_10452);
or U10710 (N_10710,N_10103,N_10229);
nand U10711 (N_10711,N_10461,N_10357);
nor U10712 (N_10712,N_10227,N_10363);
and U10713 (N_10713,N_10239,N_10217);
xnor U10714 (N_10714,N_10310,N_10004);
or U10715 (N_10715,N_10349,N_10417);
or U10716 (N_10716,N_10481,N_10197);
xor U10717 (N_10717,N_10013,N_10405);
xor U10718 (N_10718,N_10031,N_10071);
or U10719 (N_10719,N_10212,N_10457);
and U10720 (N_10720,N_10301,N_10112);
and U10721 (N_10721,N_10477,N_10023);
xor U10722 (N_10722,N_10114,N_10140);
or U10723 (N_10723,N_10050,N_10252);
nor U10724 (N_10724,N_10127,N_10080);
xnor U10725 (N_10725,N_10344,N_10157);
nand U10726 (N_10726,N_10279,N_10146);
nand U10727 (N_10727,N_10219,N_10045);
or U10728 (N_10728,N_10337,N_10090);
xor U10729 (N_10729,N_10436,N_10390);
nand U10730 (N_10730,N_10306,N_10063);
or U10731 (N_10731,N_10119,N_10255);
nand U10732 (N_10732,N_10125,N_10030);
and U10733 (N_10733,N_10189,N_10107);
xor U10734 (N_10734,N_10027,N_10184);
and U10735 (N_10735,N_10271,N_10188);
nor U10736 (N_10736,N_10341,N_10199);
nand U10737 (N_10737,N_10011,N_10261);
nand U10738 (N_10738,N_10077,N_10486);
xor U10739 (N_10739,N_10412,N_10186);
or U10740 (N_10740,N_10443,N_10220);
xnor U10741 (N_10741,N_10182,N_10391);
xor U10742 (N_10742,N_10382,N_10293);
or U10743 (N_10743,N_10423,N_10237);
nor U10744 (N_10744,N_10267,N_10328);
nor U10745 (N_10745,N_10274,N_10494);
xnor U10746 (N_10746,N_10430,N_10176);
and U10747 (N_10747,N_10437,N_10174);
nor U10748 (N_10748,N_10133,N_10375);
nor U10749 (N_10749,N_10088,N_10348);
and U10750 (N_10750,N_10175,N_10238);
nand U10751 (N_10751,N_10387,N_10380);
and U10752 (N_10752,N_10273,N_10480);
or U10753 (N_10753,N_10030,N_10357);
nand U10754 (N_10754,N_10102,N_10345);
nor U10755 (N_10755,N_10015,N_10313);
xor U10756 (N_10756,N_10112,N_10222);
or U10757 (N_10757,N_10319,N_10138);
xnor U10758 (N_10758,N_10015,N_10269);
or U10759 (N_10759,N_10163,N_10387);
or U10760 (N_10760,N_10484,N_10259);
or U10761 (N_10761,N_10215,N_10461);
or U10762 (N_10762,N_10258,N_10101);
xnor U10763 (N_10763,N_10451,N_10074);
and U10764 (N_10764,N_10169,N_10041);
or U10765 (N_10765,N_10429,N_10490);
or U10766 (N_10766,N_10107,N_10316);
or U10767 (N_10767,N_10327,N_10332);
nor U10768 (N_10768,N_10369,N_10432);
or U10769 (N_10769,N_10115,N_10380);
nor U10770 (N_10770,N_10215,N_10399);
nor U10771 (N_10771,N_10183,N_10474);
nand U10772 (N_10772,N_10383,N_10046);
and U10773 (N_10773,N_10174,N_10400);
xor U10774 (N_10774,N_10226,N_10384);
nand U10775 (N_10775,N_10478,N_10081);
nor U10776 (N_10776,N_10481,N_10105);
nand U10777 (N_10777,N_10297,N_10159);
and U10778 (N_10778,N_10328,N_10456);
nor U10779 (N_10779,N_10482,N_10151);
nand U10780 (N_10780,N_10095,N_10054);
nand U10781 (N_10781,N_10159,N_10248);
and U10782 (N_10782,N_10165,N_10490);
nand U10783 (N_10783,N_10472,N_10182);
xor U10784 (N_10784,N_10119,N_10154);
xnor U10785 (N_10785,N_10022,N_10065);
nor U10786 (N_10786,N_10149,N_10466);
xor U10787 (N_10787,N_10361,N_10188);
or U10788 (N_10788,N_10329,N_10250);
or U10789 (N_10789,N_10308,N_10430);
nor U10790 (N_10790,N_10433,N_10413);
or U10791 (N_10791,N_10332,N_10104);
or U10792 (N_10792,N_10494,N_10165);
nor U10793 (N_10793,N_10241,N_10017);
nor U10794 (N_10794,N_10252,N_10070);
nor U10795 (N_10795,N_10105,N_10053);
nor U10796 (N_10796,N_10255,N_10442);
nand U10797 (N_10797,N_10340,N_10288);
nand U10798 (N_10798,N_10285,N_10062);
nand U10799 (N_10799,N_10461,N_10230);
xor U10800 (N_10800,N_10414,N_10486);
xor U10801 (N_10801,N_10250,N_10244);
nand U10802 (N_10802,N_10237,N_10408);
nor U10803 (N_10803,N_10109,N_10188);
or U10804 (N_10804,N_10281,N_10297);
nor U10805 (N_10805,N_10481,N_10117);
nand U10806 (N_10806,N_10185,N_10311);
or U10807 (N_10807,N_10119,N_10087);
or U10808 (N_10808,N_10088,N_10281);
nand U10809 (N_10809,N_10350,N_10161);
nand U10810 (N_10810,N_10091,N_10290);
nor U10811 (N_10811,N_10414,N_10349);
nor U10812 (N_10812,N_10418,N_10359);
and U10813 (N_10813,N_10102,N_10013);
nand U10814 (N_10814,N_10155,N_10396);
nand U10815 (N_10815,N_10017,N_10311);
nor U10816 (N_10816,N_10116,N_10375);
or U10817 (N_10817,N_10397,N_10342);
xor U10818 (N_10818,N_10029,N_10091);
nand U10819 (N_10819,N_10408,N_10467);
nor U10820 (N_10820,N_10013,N_10017);
nand U10821 (N_10821,N_10452,N_10265);
nor U10822 (N_10822,N_10101,N_10160);
and U10823 (N_10823,N_10332,N_10206);
nand U10824 (N_10824,N_10026,N_10498);
nor U10825 (N_10825,N_10168,N_10437);
or U10826 (N_10826,N_10217,N_10452);
or U10827 (N_10827,N_10409,N_10004);
nor U10828 (N_10828,N_10172,N_10037);
and U10829 (N_10829,N_10226,N_10242);
nand U10830 (N_10830,N_10038,N_10486);
and U10831 (N_10831,N_10373,N_10393);
nor U10832 (N_10832,N_10075,N_10321);
nor U10833 (N_10833,N_10004,N_10417);
nor U10834 (N_10834,N_10255,N_10482);
nand U10835 (N_10835,N_10240,N_10418);
nand U10836 (N_10836,N_10349,N_10148);
and U10837 (N_10837,N_10448,N_10137);
xor U10838 (N_10838,N_10473,N_10333);
nand U10839 (N_10839,N_10392,N_10389);
xnor U10840 (N_10840,N_10463,N_10328);
xor U10841 (N_10841,N_10233,N_10471);
xor U10842 (N_10842,N_10004,N_10131);
or U10843 (N_10843,N_10474,N_10281);
nor U10844 (N_10844,N_10471,N_10068);
nor U10845 (N_10845,N_10415,N_10291);
and U10846 (N_10846,N_10090,N_10000);
nor U10847 (N_10847,N_10283,N_10447);
or U10848 (N_10848,N_10180,N_10168);
and U10849 (N_10849,N_10335,N_10269);
nand U10850 (N_10850,N_10134,N_10265);
nor U10851 (N_10851,N_10285,N_10418);
and U10852 (N_10852,N_10441,N_10341);
or U10853 (N_10853,N_10352,N_10324);
nand U10854 (N_10854,N_10113,N_10103);
and U10855 (N_10855,N_10001,N_10493);
xor U10856 (N_10856,N_10439,N_10444);
nand U10857 (N_10857,N_10072,N_10335);
nor U10858 (N_10858,N_10183,N_10047);
and U10859 (N_10859,N_10478,N_10090);
and U10860 (N_10860,N_10038,N_10331);
nor U10861 (N_10861,N_10107,N_10248);
and U10862 (N_10862,N_10356,N_10446);
and U10863 (N_10863,N_10425,N_10488);
nand U10864 (N_10864,N_10402,N_10144);
nand U10865 (N_10865,N_10150,N_10120);
or U10866 (N_10866,N_10139,N_10318);
and U10867 (N_10867,N_10181,N_10335);
and U10868 (N_10868,N_10144,N_10298);
nor U10869 (N_10869,N_10078,N_10329);
xor U10870 (N_10870,N_10281,N_10425);
nand U10871 (N_10871,N_10212,N_10071);
nand U10872 (N_10872,N_10258,N_10296);
and U10873 (N_10873,N_10339,N_10287);
nand U10874 (N_10874,N_10223,N_10250);
nor U10875 (N_10875,N_10037,N_10268);
xor U10876 (N_10876,N_10036,N_10328);
or U10877 (N_10877,N_10165,N_10102);
nand U10878 (N_10878,N_10314,N_10183);
and U10879 (N_10879,N_10362,N_10135);
and U10880 (N_10880,N_10113,N_10468);
xor U10881 (N_10881,N_10289,N_10083);
and U10882 (N_10882,N_10434,N_10120);
xnor U10883 (N_10883,N_10109,N_10235);
nand U10884 (N_10884,N_10105,N_10080);
xor U10885 (N_10885,N_10016,N_10097);
nand U10886 (N_10886,N_10026,N_10343);
nand U10887 (N_10887,N_10296,N_10138);
nor U10888 (N_10888,N_10288,N_10122);
xnor U10889 (N_10889,N_10262,N_10357);
nor U10890 (N_10890,N_10408,N_10188);
and U10891 (N_10891,N_10100,N_10416);
and U10892 (N_10892,N_10392,N_10487);
xor U10893 (N_10893,N_10046,N_10245);
and U10894 (N_10894,N_10147,N_10255);
nor U10895 (N_10895,N_10309,N_10223);
nand U10896 (N_10896,N_10457,N_10415);
xnor U10897 (N_10897,N_10449,N_10282);
nand U10898 (N_10898,N_10323,N_10126);
xnor U10899 (N_10899,N_10016,N_10047);
and U10900 (N_10900,N_10252,N_10111);
nor U10901 (N_10901,N_10314,N_10479);
nor U10902 (N_10902,N_10325,N_10225);
or U10903 (N_10903,N_10259,N_10463);
or U10904 (N_10904,N_10262,N_10236);
xor U10905 (N_10905,N_10333,N_10088);
and U10906 (N_10906,N_10089,N_10408);
xnor U10907 (N_10907,N_10493,N_10370);
or U10908 (N_10908,N_10070,N_10221);
or U10909 (N_10909,N_10047,N_10305);
xor U10910 (N_10910,N_10154,N_10099);
or U10911 (N_10911,N_10057,N_10210);
or U10912 (N_10912,N_10229,N_10200);
nand U10913 (N_10913,N_10324,N_10439);
xnor U10914 (N_10914,N_10168,N_10138);
or U10915 (N_10915,N_10391,N_10150);
xnor U10916 (N_10916,N_10127,N_10383);
nand U10917 (N_10917,N_10284,N_10487);
nand U10918 (N_10918,N_10492,N_10473);
nor U10919 (N_10919,N_10296,N_10243);
xnor U10920 (N_10920,N_10317,N_10237);
nand U10921 (N_10921,N_10430,N_10121);
nor U10922 (N_10922,N_10238,N_10308);
and U10923 (N_10923,N_10254,N_10283);
or U10924 (N_10924,N_10131,N_10428);
nor U10925 (N_10925,N_10311,N_10419);
xor U10926 (N_10926,N_10039,N_10119);
nand U10927 (N_10927,N_10364,N_10276);
and U10928 (N_10928,N_10327,N_10108);
nor U10929 (N_10929,N_10236,N_10188);
xnor U10930 (N_10930,N_10382,N_10391);
nor U10931 (N_10931,N_10447,N_10133);
or U10932 (N_10932,N_10306,N_10230);
and U10933 (N_10933,N_10040,N_10168);
nand U10934 (N_10934,N_10208,N_10350);
or U10935 (N_10935,N_10053,N_10266);
and U10936 (N_10936,N_10384,N_10034);
xnor U10937 (N_10937,N_10397,N_10012);
nand U10938 (N_10938,N_10034,N_10332);
nor U10939 (N_10939,N_10334,N_10491);
nand U10940 (N_10940,N_10293,N_10227);
xnor U10941 (N_10941,N_10047,N_10097);
nand U10942 (N_10942,N_10243,N_10274);
nor U10943 (N_10943,N_10450,N_10485);
and U10944 (N_10944,N_10411,N_10208);
or U10945 (N_10945,N_10036,N_10275);
nand U10946 (N_10946,N_10261,N_10043);
nand U10947 (N_10947,N_10457,N_10235);
and U10948 (N_10948,N_10324,N_10410);
xor U10949 (N_10949,N_10253,N_10010);
nor U10950 (N_10950,N_10391,N_10258);
nor U10951 (N_10951,N_10314,N_10184);
and U10952 (N_10952,N_10392,N_10306);
nor U10953 (N_10953,N_10006,N_10332);
xor U10954 (N_10954,N_10116,N_10221);
nand U10955 (N_10955,N_10451,N_10280);
and U10956 (N_10956,N_10458,N_10115);
or U10957 (N_10957,N_10134,N_10177);
and U10958 (N_10958,N_10343,N_10498);
xnor U10959 (N_10959,N_10138,N_10300);
nor U10960 (N_10960,N_10087,N_10391);
and U10961 (N_10961,N_10311,N_10331);
nand U10962 (N_10962,N_10178,N_10486);
and U10963 (N_10963,N_10338,N_10046);
and U10964 (N_10964,N_10087,N_10349);
xor U10965 (N_10965,N_10118,N_10169);
xnor U10966 (N_10966,N_10446,N_10190);
or U10967 (N_10967,N_10312,N_10081);
nand U10968 (N_10968,N_10363,N_10318);
and U10969 (N_10969,N_10369,N_10378);
or U10970 (N_10970,N_10469,N_10235);
and U10971 (N_10971,N_10402,N_10027);
or U10972 (N_10972,N_10447,N_10033);
xor U10973 (N_10973,N_10132,N_10186);
xor U10974 (N_10974,N_10371,N_10450);
nand U10975 (N_10975,N_10313,N_10339);
xnor U10976 (N_10976,N_10131,N_10104);
nand U10977 (N_10977,N_10083,N_10152);
nor U10978 (N_10978,N_10138,N_10315);
nor U10979 (N_10979,N_10318,N_10267);
nand U10980 (N_10980,N_10211,N_10194);
nor U10981 (N_10981,N_10087,N_10371);
xnor U10982 (N_10982,N_10291,N_10401);
and U10983 (N_10983,N_10380,N_10255);
or U10984 (N_10984,N_10470,N_10070);
and U10985 (N_10985,N_10182,N_10241);
nor U10986 (N_10986,N_10116,N_10295);
nand U10987 (N_10987,N_10271,N_10130);
nand U10988 (N_10988,N_10270,N_10380);
and U10989 (N_10989,N_10140,N_10435);
and U10990 (N_10990,N_10278,N_10400);
and U10991 (N_10991,N_10283,N_10360);
and U10992 (N_10992,N_10235,N_10084);
and U10993 (N_10993,N_10001,N_10049);
xor U10994 (N_10994,N_10164,N_10452);
or U10995 (N_10995,N_10269,N_10230);
xnor U10996 (N_10996,N_10029,N_10152);
and U10997 (N_10997,N_10343,N_10449);
or U10998 (N_10998,N_10051,N_10439);
nor U10999 (N_10999,N_10093,N_10404);
or U11000 (N_11000,N_10790,N_10546);
nor U11001 (N_11001,N_10621,N_10788);
nand U11002 (N_11002,N_10797,N_10658);
nor U11003 (N_11003,N_10698,N_10535);
and U11004 (N_11004,N_10666,N_10518);
xor U11005 (N_11005,N_10956,N_10896);
xor U11006 (N_11006,N_10601,N_10882);
nand U11007 (N_11007,N_10954,N_10857);
nand U11008 (N_11008,N_10655,N_10555);
nor U11009 (N_11009,N_10708,N_10829);
or U11010 (N_11010,N_10683,N_10736);
nand U11011 (N_11011,N_10766,N_10802);
nand U11012 (N_11012,N_10938,N_10914);
xor U11013 (N_11013,N_10504,N_10691);
nand U11014 (N_11014,N_10791,N_10558);
or U11015 (N_11015,N_10606,N_10512);
xnor U11016 (N_11016,N_10822,N_10587);
xor U11017 (N_11017,N_10677,N_10984);
or U11018 (N_11018,N_10521,N_10975);
nand U11019 (N_11019,N_10687,N_10615);
nor U11020 (N_11020,N_10780,N_10685);
nor U11021 (N_11021,N_10554,N_10697);
nand U11022 (N_11022,N_10924,N_10508);
nand U11023 (N_11023,N_10837,N_10955);
nor U11024 (N_11024,N_10622,N_10978);
and U11025 (N_11025,N_10915,N_10891);
or U11026 (N_11026,N_10648,N_10541);
nor U11027 (N_11027,N_10646,N_10865);
or U11028 (N_11028,N_10560,N_10787);
xnor U11029 (N_11029,N_10534,N_10653);
nand U11030 (N_11030,N_10768,N_10823);
or U11031 (N_11031,N_10721,N_10966);
or U11032 (N_11032,N_10819,N_10809);
nand U11033 (N_11033,N_10796,N_10827);
xnor U11034 (N_11034,N_10593,N_10784);
xnor U11035 (N_11035,N_10961,N_10644);
nand U11036 (N_11036,N_10573,N_10812);
nor U11037 (N_11037,N_10623,N_10502);
nor U11038 (N_11038,N_10886,N_10759);
and U11039 (N_11039,N_10547,N_10939);
or U11040 (N_11040,N_10716,N_10761);
or U11041 (N_11041,N_10755,N_10572);
nor U11042 (N_11042,N_10597,N_10507);
xnor U11043 (N_11043,N_10964,N_10866);
and U11044 (N_11044,N_10634,N_10556);
nand U11045 (N_11045,N_10569,N_10859);
nand U11046 (N_11046,N_10673,N_10997);
nor U11047 (N_11047,N_10808,N_10847);
and U11048 (N_11048,N_10717,N_10795);
or U11049 (N_11049,N_10506,N_10968);
and U11050 (N_11050,N_10663,N_10722);
or U11051 (N_11051,N_10920,N_10878);
xor U11052 (N_11052,N_10962,N_10856);
nor U11053 (N_11053,N_10540,N_10725);
and U11054 (N_11054,N_10636,N_10945);
xnor U11055 (N_11055,N_10603,N_10758);
nor U11056 (N_11056,N_10906,N_10999);
or U11057 (N_11057,N_10583,N_10713);
or U11058 (N_11058,N_10927,N_10699);
and U11059 (N_11059,N_10660,N_10563);
xor U11060 (N_11060,N_10596,N_10979);
and U11061 (N_11061,N_10779,N_10963);
nand U11062 (N_11062,N_10833,N_10749);
and U11063 (N_11063,N_10888,N_10638);
nor U11064 (N_11064,N_10575,N_10907);
and U11065 (N_11065,N_10625,N_10935);
and U11066 (N_11066,N_10537,N_10574);
or U11067 (N_11067,N_10930,N_10928);
and U11068 (N_11068,N_10871,N_10519);
nor U11069 (N_11069,N_10618,N_10855);
nor U11070 (N_11070,N_10689,N_10885);
nand U11071 (N_11071,N_10799,N_10510);
and U11072 (N_11072,N_10937,N_10843);
nor U11073 (N_11073,N_10582,N_10899);
or U11074 (N_11074,N_10592,N_10693);
nand U11075 (N_11075,N_10501,N_10738);
and U11076 (N_11076,N_10951,N_10835);
or U11077 (N_11077,N_10821,N_10652);
and U11078 (N_11078,N_10694,N_10913);
and U11079 (N_11079,N_10514,N_10986);
xor U11080 (N_11080,N_10630,N_10853);
nand U11081 (N_11081,N_10810,N_10971);
xnor U11082 (N_11082,N_10626,N_10988);
and U11083 (N_11083,N_10728,N_10604);
and U11084 (N_11084,N_10500,N_10909);
nand U11085 (N_11085,N_10958,N_10741);
nor U11086 (N_11086,N_10861,N_10633);
and U11087 (N_11087,N_10996,N_10839);
nor U11088 (N_11088,N_10676,N_10711);
or U11089 (N_11089,N_10820,N_10789);
nand U11090 (N_11090,N_10849,N_10523);
nand U11091 (N_11091,N_10900,N_10680);
nand U11092 (N_11092,N_10854,N_10774);
nand U11093 (N_11093,N_10602,N_10911);
and U11094 (N_11094,N_10559,N_10726);
or U11095 (N_11095,N_10753,N_10760);
and U11096 (N_11096,N_10584,N_10884);
nor U11097 (N_11097,N_10794,N_10917);
nor U11098 (N_11098,N_10511,N_10730);
and U11099 (N_11099,N_10792,N_10723);
xor U11100 (N_11100,N_10664,N_10752);
xnor U11101 (N_11101,N_10724,N_10629);
and U11102 (N_11102,N_10991,N_10897);
or U11103 (N_11103,N_10645,N_10929);
and U11104 (N_11104,N_10684,N_10674);
nor U11105 (N_11105,N_10959,N_10804);
nor U11106 (N_11106,N_10903,N_10588);
or U11107 (N_11107,N_10834,N_10826);
xnor U11108 (N_11108,N_10515,N_10887);
or U11109 (N_11109,N_10750,N_10931);
nor U11110 (N_11110,N_10870,N_10719);
and U11111 (N_11111,N_10651,N_10895);
and U11112 (N_11112,N_10943,N_10889);
xnor U11113 (N_11113,N_10513,N_10776);
and U11114 (N_11114,N_10894,N_10946);
or U11115 (N_11115,N_10967,N_10902);
nor U11116 (N_11116,N_10585,N_10985);
nand U11117 (N_11117,N_10960,N_10934);
nor U11118 (N_11118,N_10570,N_10990);
nand U11119 (N_11119,N_10543,N_10591);
and U11120 (N_11120,N_10881,N_10922);
and U11121 (N_11121,N_10817,N_10539);
xor U11122 (N_11122,N_10702,N_10754);
and U11123 (N_11123,N_10912,N_10505);
or U11124 (N_11124,N_10748,N_10608);
or U11125 (N_11125,N_10670,N_10764);
nand U11126 (N_11126,N_10864,N_10745);
nand U11127 (N_11127,N_10973,N_10667);
nor U11128 (N_11128,N_10781,N_10631);
nor U11129 (N_11129,N_10987,N_10976);
xnor U11130 (N_11130,N_10824,N_10654);
xnor U11131 (N_11131,N_10714,N_10650);
nand U11132 (N_11132,N_10607,N_10688);
nor U11133 (N_11133,N_10747,N_10552);
or U11134 (N_11134,N_10969,N_10579);
nand U11135 (N_11135,N_10800,N_10798);
nor U11136 (N_11136,N_10877,N_10614);
nand U11137 (N_11137,N_10948,N_10825);
nand U11138 (N_11138,N_10947,N_10957);
nor U11139 (N_11139,N_10977,N_10517);
nor U11140 (N_11140,N_10844,N_10994);
and U11141 (N_11141,N_10710,N_10757);
or U11142 (N_11142,N_10709,N_10706);
nand U11143 (N_11143,N_10720,N_10628);
or U11144 (N_11144,N_10732,N_10617);
or U11145 (N_11145,N_10814,N_10801);
nand U11146 (N_11146,N_10503,N_10734);
or U11147 (N_11147,N_10594,N_10863);
xor U11148 (N_11148,N_10729,N_10549);
nor U11149 (N_11149,N_10918,N_10611);
or U11150 (N_11150,N_10568,N_10828);
xor U11151 (N_11151,N_10703,N_10940);
and U11152 (N_11152,N_10530,N_10692);
xnor U11153 (N_11153,N_10845,N_10551);
and U11154 (N_11154,N_10769,N_10662);
nor U11155 (N_11155,N_10590,N_10620);
and U11156 (N_11156,N_10532,N_10923);
and U11157 (N_11157,N_10657,N_10767);
nand U11158 (N_11158,N_10793,N_10893);
nand U11159 (N_11159,N_10671,N_10803);
or U11160 (N_11160,N_10580,N_10612);
nand U11161 (N_11161,N_10553,N_10740);
nor U11162 (N_11162,N_10735,N_10525);
xor U11163 (N_11163,N_10995,N_10522);
or U11164 (N_11164,N_10850,N_10815);
or U11165 (N_11165,N_10727,N_10531);
xnor U11166 (N_11166,N_10528,N_10883);
xor U11167 (N_11167,N_10647,N_10936);
nand U11168 (N_11168,N_10869,N_10542);
or U11169 (N_11169,N_10974,N_10679);
nand U11170 (N_11170,N_10805,N_10695);
nor U11171 (N_11171,N_10571,N_10981);
or U11172 (N_11172,N_10944,N_10840);
nand U11173 (N_11173,N_10953,N_10627);
nand U11174 (N_11174,N_10763,N_10661);
nand U11175 (N_11175,N_10529,N_10851);
xor U11176 (N_11176,N_10970,N_10682);
nand U11177 (N_11177,N_10609,N_10905);
and U11178 (N_11178,N_10635,N_10785);
nand U11179 (N_11179,N_10875,N_10595);
xnor U11180 (N_11180,N_10678,N_10743);
and U11181 (N_11181,N_10783,N_10831);
or U11182 (N_11182,N_10860,N_10901);
nand U11183 (N_11183,N_10696,N_10868);
nand U11184 (N_11184,N_10756,N_10830);
nor U11185 (N_11185,N_10811,N_10807);
or U11186 (N_11186,N_10538,N_10898);
or U11187 (N_11187,N_10516,N_10562);
or U11188 (N_11188,N_10919,N_10576);
and U11189 (N_11189,N_10933,N_10715);
or U11190 (N_11190,N_10567,N_10941);
nor U11191 (N_11191,N_10704,N_10656);
and U11192 (N_11192,N_10848,N_10565);
or U11193 (N_11193,N_10545,N_10643);
and U11194 (N_11194,N_10925,N_10952);
nand U11195 (N_11195,N_10642,N_10548);
xor U11196 (N_11196,N_10700,N_10782);
and U11197 (N_11197,N_10578,N_10733);
nor U11198 (N_11198,N_10520,N_10813);
or U11199 (N_11199,N_10838,N_10841);
nor U11200 (N_11200,N_10836,N_10904);
and U11201 (N_11201,N_10862,N_10600);
nand U11202 (N_11202,N_10874,N_10605);
and U11203 (N_11203,N_10916,N_10557);
or U11204 (N_11204,N_10533,N_10775);
nand U11205 (N_11205,N_10806,N_10598);
or U11206 (N_11206,N_10846,N_10950);
nand U11207 (N_11207,N_10873,N_10589);
xor U11208 (N_11208,N_10972,N_10942);
or U11209 (N_11209,N_10564,N_10773);
xnor U11210 (N_11210,N_10737,N_10949);
or U11211 (N_11211,N_10852,N_10669);
nor U11212 (N_11212,N_10739,N_10993);
xor U11213 (N_11213,N_10982,N_10526);
and U11214 (N_11214,N_10867,N_10613);
or U11215 (N_11215,N_10816,N_10842);
nand U11216 (N_11216,N_10639,N_10998);
or U11217 (N_11217,N_10610,N_10980);
and U11218 (N_11218,N_10765,N_10705);
nor U11219 (N_11219,N_10672,N_10778);
and U11220 (N_11220,N_10879,N_10632);
nor U11221 (N_11221,N_10983,N_10599);
and U11222 (N_11222,N_10762,N_10675);
nand U11223 (N_11223,N_10637,N_10744);
xnor U11224 (N_11224,N_10659,N_10908);
or U11225 (N_11225,N_10832,N_10681);
nand U11226 (N_11226,N_10771,N_10932);
nor U11227 (N_11227,N_10640,N_10524);
or U11228 (N_11228,N_10561,N_10581);
nand U11229 (N_11229,N_10668,N_10921);
or U11230 (N_11230,N_10786,N_10772);
or U11231 (N_11231,N_10777,N_10690);
xnor U11232 (N_11232,N_10619,N_10649);
or U11233 (N_11233,N_10872,N_10665);
nand U11234 (N_11234,N_10536,N_10858);
nand U11235 (N_11235,N_10926,N_10707);
or U11236 (N_11236,N_10624,N_10686);
xor U11237 (N_11237,N_10577,N_10770);
or U11238 (N_11238,N_10731,N_10880);
nor U11239 (N_11239,N_10989,N_10616);
or U11240 (N_11240,N_10712,N_10701);
and U11241 (N_11241,N_10746,N_10742);
nor U11242 (N_11242,N_10876,N_10892);
nor U11243 (N_11243,N_10544,N_10566);
xor U11244 (N_11244,N_10509,N_10527);
xor U11245 (N_11245,N_10910,N_10751);
xnor U11246 (N_11246,N_10586,N_10890);
xnor U11247 (N_11247,N_10818,N_10965);
and U11248 (N_11248,N_10641,N_10992);
nand U11249 (N_11249,N_10550,N_10718);
and U11250 (N_11250,N_10848,N_10669);
xor U11251 (N_11251,N_10932,N_10930);
nor U11252 (N_11252,N_10523,N_10823);
xor U11253 (N_11253,N_10842,N_10549);
and U11254 (N_11254,N_10605,N_10776);
and U11255 (N_11255,N_10642,N_10601);
or U11256 (N_11256,N_10796,N_10793);
or U11257 (N_11257,N_10563,N_10601);
or U11258 (N_11258,N_10935,N_10992);
xor U11259 (N_11259,N_10509,N_10837);
nor U11260 (N_11260,N_10660,N_10514);
and U11261 (N_11261,N_10624,N_10983);
xor U11262 (N_11262,N_10903,N_10574);
and U11263 (N_11263,N_10756,N_10670);
nand U11264 (N_11264,N_10569,N_10751);
or U11265 (N_11265,N_10725,N_10787);
nand U11266 (N_11266,N_10825,N_10802);
or U11267 (N_11267,N_10757,N_10652);
xor U11268 (N_11268,N_10914,N_10937);
and U11269 (N_11269,N_10935,N_10907);
xor U11270 (N_11270,N_10741,N_10781);
nand U11271 (N_11271,N_10643,N_10584);
nand U11272 (N_11272,N_10631,N_10841);
or U11273 (N_11273,N_10748,N_10629);
nand U11274 (N_11274,N_10702,N_10874);
and U11275 (N_11275,N_10938,N_10899);
nand U11276 (N_11276,N_10860,N_10834);
nor U11277 (N_11277,N_10861,N_10785);
nor U11278 (N_11278,N_10747,N_10766);
nand U11279 (N_11279,N_10985,N_10721);
or U11280 (N_11280,N_10504,N_10762);
nand U11281 (N_11281,N_10547,N_10856);
nand U11282 (N_11282,N_10743,N_10835);
nand U11283 (N_11283,N_10921,N_10621);
nor U11284 (N_11284,N_10819,N_10605);
nand U11285 (N_11285,N_10754,N_10872);
nand U11286 (N_11286,N_10999,N_10641);
nor U11287 (N_11287,N_10625,N_10731);
nand U11288 (N_11288,N_10665,N_10577);
or U11289 (N_11289,N_10630,N_10813);
xor U11290 (N_11290,N_10773,N_10552);
or U11291 (N_11291,N_10543,N_10857);
or U11292 (N_11292,N_10726,N_10988);
xnor U11293 (N_11293,N_10690,N_10907);
xnor U11294 (N_11294,N_10857,N_10911);
xnor U11295 (N_11295,N_10846,N_10839);
nand U11296 (N_11296,N_10627,N_10529);
nor U11297 (N_11297,N_10686,N_10890);
xnor U11298 (N_11298,N_10552,N_10520);
xor U11299 (N_11299,N_10954,N_10945);
nor U11300 (N_11300,N_10500,N_10509);
nand U11301 (N_11301,N_10665,N_10978);
nand U11302 (N_11302,N_10833,N_10699);
xor U11303 (N_11303,N_10528,N_10957);
nand U11304 (N_11304,N_10528,N_10524);
nor U11305 (N_11305,N_10510,N_10702);
or U11306 (N_11306,N_10816,N_10659);
xor U11307 (N_11307,N_10502,N_10781);
and U11308 (N_11308,N_10839,N_10885);
nor U11309 (N_11309,N_10865,N_10527);
nand U11310 (N_11310,N_10833,N_10751);
nand U11311 (N_11311,N_10920,N_10887);
nor U11312 (N_11312,N_10518,N_10815);
nor U11313 (N_11313,N_10749,N_10711);
nand U11314 (N_11314,N_10810,N_10978);
nor U11315 (N_11315,N_10639,N_10852);
or U11316 (N_11316,N_10764,N_10831);
and U11317 (N_11317,N_10537,N_10984);
nor U11318 (N_11318,N_10728,N_10796);
or U11319 (N_11319,N_10582,N_10611);
and U11320 (N_11320,N_10647,N_10967);
xnor U11321 (N_11321,N_10975,N_10810);
xor U11322 (N_11322,N_10984,N_10691);
xor U11323 (N_11323,N_10695,N_10953);
nand U11324 (N_11324,N_10705,N_10525);
and U11325 (N_11325,N_10893,N_10644);
nand U11326 (N_11326,N_10909,N_10633);
nor U11327 (N_11327,N_10808,N_10897);
nor U11328 (N_11328,N_10731,N_10741);
nand U11329 (N_11329,N_10598,N_10708);
nor U11330 (N_11330,N_10695,N_10976);
xor U11331 (N_11331,N_10807,N_10736);
and U11332 (N_11332,N_10829,N_10839);
nor U11333 (N_11333,N_10956,N_10943);
or U11334 (N_11334,N_10556,N_10820);
nand U11335 (N_11335,N_10598,N_10572);
and U11336 (N_11336,N_10918,N_10594);
nor U11337 (N_11337,N_10832,N_10528);
and U11338 (N_11338,N_10526,N_10709);
xnor U11339 (N_11339,N_10566,N_10508);
nor U11340 (N_11340,N_10586,N_10637);
or U11341 (N_11341,N_10569,N_10864);
nor U11342 (N_11342,N_10908,N_10705);
or U11343 (N_11343,N_10669,N_10989);
and U11344 (N_11344,N_10646,N_10531);
nand U11345 (N_11345,N_10941,N_10618);
nor U11346 (N_11346,N_10713,N_10764);
nor U11347 (N_11347,N_10586,N_10546);
xnor U11348 (N_11348,N_10630,N_10733);
xor U11349 (N_11349,N_10650,N_10760);
and U11350 (N_11350,N_10861,N_10768);
xor U11351 (N_11351,N_10652,N_10707);
nand U11352 (N_11352,N_10617,N_10769);
or U11353 (N_11353,N_10665,N_10938);
nor U11354 (N_11354,N_10572,N_10697);
or U11355 (N_11355,N_10552,N_10782);
or U11356 (N_11356,N_10582,N_10981);
nand U11357 (N_11357,N_10898,N_10612);
or U11358 (N_11358,N_10932,N_10602);
xor U11359 (N_11359,N_10877,N_10650);
nand U11360 (N_11360,N_10907,N_10872);
and U11361 (N_11361,N_10792,N_10503);
xnor U11362 (N_11362,N_10547,N_10731);
xnor U11363 (N_11363,N_10675,N_10898);
nor U11364 (N_11364,N_10845,N_10908);
xnor U11365 (N_11365,N_10529,N_10533);
xor U11366 (N_11366,N_10859,N_10870);
or U11367 (N_11367,N_10724,N_10570);
and U11368 (N_11368,N_10655,N_10743);
xor U11369 (N_11369,N_10526,N_10731);
or U11370 (N_11370,N_10721,N_10725);
and U11371 (N_11371,N_10506,N_10611);
nor U11372 (N_11372,N_10985,N_10694);
nor U11373 (N_11373,N_10717,N_10733);
nand U11374 (N_11374,N_10501,N_10571);
or U11375 (N_11375,N_10507,N_10902);
nand U11376 (N_11376,N_10624,N_10945);
or U11377 (N_11377,N_10769,N_10534);
and U11378 (N_11378,N_10541,N_10777);
or U11379 (N_11379,N_10798,N_10753);
or U11380 (N_11380,N_10960,N_10571);
and U11381 (N_11381,N_10767,N_10874);
or U11382 (N_11382,N_10632,N_10728);
nand U11383 (N_11383,N_10657,N_10748);
nand U11384 (N_11384,N_10703,N_10668);
or U11385 (N_11385,N_10944,N_10821);
nor U11386 (N_11386,N_10535,N_10757);
nor U11387 (N_11387,N_10753,N_10738);
and U11388 (N_11388,N_10689,N_10862);
nand U11389 (N_11389,N_10672,N_10708);
nor U11390 (N_11390,N_10756,N_10944);
and U11391 (N_11391,N_10813,N_10725);
or U11392 (N_11392,N_10525,N_10561);
and U11393 (N_11393,N_10969,N_10755);
or U11394 (N_11394,N_10990,N_10805);
or U11395 (N_11395,N_10767,N_10555);
or U11396 (N_11396,N_10817,N_10934);
nand U11397 (N_11397,N_10653,N_10960);
and U11398 (N_11398,N_10681,N_10828);
xnor U11399 (N_11399,N_10756,N_10695);
nand U11400 (N_11400,N_10761,N_10756);
nand U11401 (N_11401,N_10735,N_10981);
xnor U11402 (N_11402,N_10652,N_10655);
nand U11403 (N_11403,N_10790,N_10818);
or U11404 (N_11404,N_10633,N_10851);
and U11405 (N_11405,N_10722,N_10583);
xnor U11406 (N_11406,N_10589,N_10888);
xor U11407 (N_11407,N_10990,N_10639);
nor U11408 (N_11408,N_10630,N_10719);
xnor U11409 (N_11409,N_10712,N_10678);
or U11410 (N_11410,N_10772,N_10753);
and U11411 (N_11411,N_10832,N_10745);
nor U11412 (N_11412,N_10509,N_10770);
nor U11413 (N_11413,N_10650,N_10672);
nor U11414 (N_11414,N_10917,N_10652);
or U11415 (N_11415,N_10648,N_10926);
and U11416 (N_11416,N_10597,N_10870);
nor U11417 (N_11417,N_10662,N_10539);
and U11418 (N_11418,N_10746,N_10830);
nor U11419 (N_11419,N_10583,N_10799);
or U11420 (N_11420,N_10513,N_10770);
and U11421 (N_11421,N_10813,N_10608);
or U11422 (N_11422,N_10740,N_10708);
or U11423 (N_11423,N_10797,N_10669);
nand U11424 (N_11424,N_10925,N_10685);
or U11425 (N_11425,N_10965,N_10595);
nand U11426 (N_11426,N_10909,N_10678);
or U11427 (N_11427,N_10820,N_10782);
or U11428 (N_11428,N_10882,N_10589);
and U11429 (N_11429,N_10761,N_10776);
nor U11430 (N_11430,N_10595,N_10936);
and U11431 (N_11431,N_10955,N_10662);
and U11432 (N_11432,N_10827,N_10655);
nor U11433 (N_11433,N_10940,N_10688);
or U11434 (N_11434,N_10920,N_10617);
and U11435 (N_11435,N_10880,N_10660);
or U11436 (N_11436,N_10669,N_10788);
nand U11437 (N_11437,N_10805,N_10669);
nor U11438 (N_11438,N_10804,N_10680);
nand U11439 (N_11439,N_10803,N_10972);
nor U11440 (N_11440,N_10772,N_10639);
or U11441 (N_11441,N_10579,N_10530);
nand U11442 (N_11442,N_10739,N_10504);
nor U11443 (N_11443,N_10966,N_10584);
or U11444 (N_11444,N_10969,N_10591);
xnor U11445 (N_11445,N_10901,N_10853);
nand U11446 (N_11446,N_10583,N_10850);
nor U11447 (N_11447,N_10577,N_10698);
or U11448 (N_11448,N_10844,N_10607);
nor U11449 (N_11449,N_10943,N_10722);
nor U11450 (N_11450,N_10552,N_10752);
or U11451 (N_11451,N_10865,N_10538);
nor U11452 (N_11452,N_10639,N_10736);
nor U11453 (N_11453,N_10891,N_10948);
xor U11454 (N_11454,N_10610,N_10856);
and U11455 (N_11455,N_10967,N_10696);
xnor U11456 (N_11456,N_10958,N_10633);
xor U11457 (N_11457,N_10830,N_10577);
and U11458 (N_11458,N_10562,N_10737);
or U11459 (N_11459,N_10634,N_10670);
nand U11460 (N_11460,N_10558,N_10895);
and U11461 (N_11461,N_10865,N_10924);
or U11462 (N_11462,N_10758,N_10647);
nand U11463 (N_11463,N_10619,N_10772);
and U11464 (N_11464,N_10859,N_10502);
or U11465 (N_11465,N_10944,N_10564);
or U11466 (N_11466,N_10700,N_10953);
or U11467 (N_11467,N_10583,N_10650);
nor U11468 (N_11468,N_10793,N_10655);
xor U11469 (N_11469,N_10857,N_10517);
nor U11470 (N_11470,N_10704,N_10727);
nand U11471 (N_11471,N_10534,N_10926);
and U11472 (N_11472,N_10515,N_10994);
and U11473 (N_11473,N_10882,N_10583);
xor U11474 (N_11474,N_10563,N_10655);
nand U11475 (N_11475,N_10573,N_10810);
nor U11476 (N_11476,N_10676,N_10675);
or U11477 (N_11477,N_10744,N_10812);
and U11478 (N_11478,N_10738,N_10697);
and U11479 (N_11479,N_10671,N_10557);
nand U11480 (N_11480,N_10953,N_10917);
and U11481 (N_11481,N_10986,N_10547);
nor U11482 (N_11482,N_10879,N_10687);
nand U11483 (N_11483,N_10591,N_10892);
or U11484 (N_11484,N_10596,N_10903);
xor U11485 (N_11485,N_10867,N_10519);
xnor U11486 (N_11486,N_10502,N_10666);
or U11487 (N_11487,N_10814,N_10824);
and U11488 (N_11488,N_10535,N_10798);
nor U11489 (N_11489,N_10976,N_10735);
nand U11490 (N_11490,N_10984,N_10889);
and U11491 (N_11491,N_10911,N_10964);
or U11492 (N_11492,N_10913,N_10640);
xor U11493 (N_11493,N_10784,N_10613);
nor U11494 (N_11494,N_10814,N_10761);
nor U11495 (N_11495,N_10626,N_10877);
and U11496 (N_11496,N_10514,N_10502);
and U11497 (N_11497,N_10900,N_10904);
xnor U11498 (N_11498,N_10926,N_10718);
nor U11499 (N_11499,N_10721,N_10694);
xor U11500 (N_11500,N_11040,N_11039);
and U11501 (N_11501,N_11162,N_11445);
nor U11502 (N_11502,N_11411,N_11433);
xor U11503 (N_11503,N_11163,N_11158);
nand U11504 (N_11504,N_11448,N_11356);
xnor U11505 (N_11505,N_11154,N_11145);
or U11506 (N_11506,N_11498,N_11200);
nor U11507 (N_11507,N_11443,N_11206);
or U11508 (N_11508,N_11314,N_11463);
nand U11509 (N_11509,N_11002,N_11435);
and U11510 (N_11510,N_11344,N_11102);
or U11511 (N_11511,N_11101,N_11143);
xnor U11512 (N_11512,N_11460,N_11149);
and U11513 (N_11513,N_11345,N_11017);
nand U11514 (N_11514,N_11380,N_11168);
xor U11515 (N_11515,N_11268,N_11115);
or U11516 (N_11516,N_11100,N_11399);
nand U11517 (N_11517,N_11376,N_11370);
and U11518 (N_11518,N_11069,N_11247);
or U11519 (N_11519,N_11263,N_11325);
and U11520 (N_11520,N_11064,N_11486);
nand U11521 (N_11521,N_11060,N_11201);
nand U11522 (N_11522,N_11442,N_11082);
nand U11523 (N_11523,N_11042,N_11419);
or U11524 (N_11524,N_11093,N_11205);
and U11525 (N_11525,N_11262,N_11342);
xnor U11526 (N_11526,N_11490,N_11131);
nor U11527 (N_11527,N_11312,N_11138);
and U11528 (N_11528,N_11241,N_11333);
or U11529 (N_11529,N_11006,N_11186);
nand U11530 (N_11530,N_11192,N_11375);
and U11531 (N_11531,N_11235,N_11140);
xor U11532 (N_11532,N_11382,N_11352);
nand U11533 (N_11533,N_11215,N_11364);
nor U11534 (N_11534,N_11030,N_11329);
nand U11535 (N_11535,N_11033,N_11450);
nand U11536 (N_11536,N_11198,N_11425);
nor U11537 (N_11537,N_11381,N_11407);
nor U11538 (N_11538,N_11056,N_11146);
and U11539 (N_11539,N_11000,N_11288);
and U11540 (N_11540,N_11319,N_11071);
or U11541 (N_11541,N_11353,N_11208);
nand U11542 (N_11542,N_11103,N_11219);
xnor U11543 (N_11543,N_11127,N_11293);
nor U11544 (N_11544,N_11156,N_11469);
nor U11545 (N_11545,N_11294,N_11456);
xnor U11546 (N_11546,N_11484,N_11067);
nand U11547 (N_11547,N_11359,N_11108);
or U11548 (N_11548,N_11087,N_11479);
nor U11549 (N_11549,N_11130,N_11091);
or U11550 (N_11550,N_11434,N_11080);
xor U11551 (N_11551,N_11045,N_11281);
nor U11552 (N_11552,N_11270,N_11323);
xor U11553 (N_11553,N_11144,N_11259);
and U11554 (N_11554,N_11112,N_11257);
or U11555 (N_11555,N_11298,N_11466);
nor U11556 (N_11556,N_11349,N_11409);
nor U11557 (N_11557,N_11015,N_11309);
nor U11558 (N_11558,N_11034,N_11326);
or U11559 (N_11559,N_11487,N_11141);
xor U11560 (N_11560,N_11142,N_11021);
or U11561 (N_11561,N_11014,N_11222);
or U11562 (N_11562,N_11454,N_11003);
nand U11563 (N_11563,N_11491,N_11134);
nor U11564 (N_11564,N_11387,N_11343);
nand U11565 (N_11565,N_11306,N_11165);
or U11566 (N_11566,N_11248,N_11438);
or U11567 (N_11567,N_11070,N_11077);
or U11568 (N_11568,N_11052,N_11148);
nand U11569 (N_11569,N_11055,N_11078);
nand U11570 (N_11570,N_11444,N_11427);
xnor U11571 (N_11571,N_11389,N_11386);
xor U11572 (N_11572,N_11255,N_11347);
xnor U11573 (N_11573,N_11124,N_11280);
xnor U11574 (N_11574,N_11350,N_11360);
nand U11575 (N_11575,N_11265,N_11129);
and U11576 (N_11576,N_11308,N_11106);
and U11577 (N_11577,N_11458,N_11170);
nor U11578 (N_11578,N_11310,N_11008);
or U11579 (N_11579,N_11098,N_11218);
xnor U11580 (N_11580,N_11181,N_11011);
nand U11581 (N_11581,N_11239,N_11079);
nand U11582 (N_11582,N_11053,N_11361);
nor U11583 (N_11583,N_11446,N_11249);
and U11584 (N_11584,N_11373,N_11049);
nand U11585 (N_11585,N_11429,N_11467);
and U11586 (N_11586,N_11275,N_11152);
and U11587 (N_11587,N_11047,N_11114);
xor U11588 (N_11588,N_11245,N_11224);
nor U11589 (N_11589,N_11461,N_11048);
nand U11590 (N_11590,N_11377,N_11202);
xnor U11591 (N_11591,N_11197,N_11276);
nand U11592 (N_11592,N_11118,N_11385);
nand U11593 (N_11593,N_11324,N_11203);
or U11594 (N_11594,N_11366,N_11475);
and U11595 (N_11595,N_11372,N_11105);
or U11596 (N_11596,N_11032,N_11299);
nand U11597 (N_11597,N_11256,N_11358);
nor U11598 (N_11598,N_11151,N_11439);
or U11599 (N_11599,N_11404,N_11187);
xnor U11600 (N_11600,N_11395,N_11421);
nand U11601 (N_11601,N_11405,N_11004);
and U11602 (N_11602,N_11190,N_11279);
and U11603 (N_11603,N_11258,N_11212);
and U11604 (N_11604,N_11174,N_11044);
nand U11605 (N_11605,N_11058,N_11150);
and U11606 (N_11606,N_11242,N_11043);
nand U11607 (N_11607,N_11182,N_11328);
nor U11608 (N_11608,N_11195,N_11408);
nand U11609 (N_11609,N_11173,N_11396);
nor U11610 (N_11610,N_11228,N_11213);
xnor U11611 (N_11611,N_11357,N_11261);
nand U11612 (N_11612,N_11133,N_11217);
nor U11613 (N_11613,N_11313,N_11413);
xnor U11614 (N_11614,N_11188,N_11480);
nor U11615 (N_11615,N_11172,N_11063);
or U11616 (N_11616,N_11121,N_11009);
or U11617 (N_11617,N_11481,N_11013);
xor U11618 (N_11618,N_11365,N_11311);
and U11619 (N_11619,N_11379,N_11492);
nand U11620 (N_11620,N_11171,N_11119);
and U11621 (N_11621,N_11096,N_11416);
xor U11622 (N_11622,N_11430,N_11295);
and U11623 (N_11623,N_11453,N_11391);
nand U11624 (N_11624,N_11305,N_11022);
nor U11625 (N_11625,N_11059,N_11126);
nand U11626 (N_11626,N_11081,N_11230);
or U11627 (N_11627,N_11260,N_11488);
or U11628 (N_11628,N_11493,N_11199);
nand U11629 (N_11629,N_11403,N_11337);
nor U11630 (N_11630,N_11083,N_11193);
xnor U11631 (N_11631,N_11234,N_11483);
nand U11632 (N_11632,N_11051,N_11169);
nand U11633 (N_11633,N_11191,N_11135);
xnor U11634 (N_11634,N_11465,N_11076);
nor U11635 (N_11635,N_11335,N_11220);
or U11636 (N_11636,N_11354,N_11164);
nor U11637 (N_11637,N_11016,N_11406);
nor U11638 (N_11638,N_11027,N_11420);
nand U11639 (N_11639,N_11029,N_11336);
nand U11640 (N_11640,N_11147,N_11497);
nand U11641 (N_11641,N_11046,N_11287);
or U11642 (N_11642,N_11473,N_11316);
nand U11643 (N_11643,N_11074,N_11010);
nor U11644 (N_11644,N_11221,N_11179);
nor U11645 (N_11645,N_11153,N_11332);
nand U11646 (N_11646,N_11291,N_11412);
or U11647 (N_11647,N_11159,N_11116);
or U11648 (N_11648,N_11274,N_11072);
nand U11649 (N_11649,N_11303,N_11068);
and U11650 (N_11650,N_11225,N_11401);
xnor U11651 (N_11651,N_11334,N_11400);
nand U11652 (N_11652,N_11289,N_11246);
xor U11653 (N_11653,N_11297,N_11229);
or U11654 (N_11654,N_11478,N_11318);
xor U11655 (N_11655,N_11322,N_11415);
xnor U11656 (N_11656,N_11424,N_11211);
xor U11657 (N_11657,N_11264,N_11099);
nor U11658 (N_11658,N_11054,N_11066);
nor U11659 (N_11659,N_11273,N_11041);
xnor U11660 (N_11660,N_11038,N_11109);
xor U11661 (N_11661,N_11455,N_11175);
nand U11662 (N_11662,N_11378,N_11494);
or U11663 (N_11663,N_11167,N_11183);
or U11664 (N_11664,N_11431,N_11094);
nand U11665 (N_11665,N_11123,N_11339);
xnor U11666 (N_11666,N_11307,N_11237);
xnor U11667 (N_11667,N_11452,N_11477);
or U11668 (N_11668,N_11457,N_11132);
or U11669 (N_11669,N_11338,N_11184);
nand U11670 (N_11670,N_11346,N_11271);
nand U11671 (N_11671,N_11436,N_11062);
nand U11672 (N_11672,N_11292,N_11253);
or U11673 (N_11673,N_11089,N_11423);
or U11674 (N_11674,N_11111,N_11459);
nand U11675 (N_11675,N_11428,N_11110);
or U11676 (N_11676,N_11223,N_11231);
nor U11677 (N_11677,N_11464,N_11470);
xor U11678 (N_11678,N_11384,N_11474);
nor U11679 (N_11679,N_11422,N_11166);
nand U11680 (N_11680,N_11296,N_11180);
xor U11681 (N_11681,N_11057,N_11398);
nor U11682 (N_11682,N_11236,N_11432);
or U11683 (N_11683,N_11269,N_11496);
xor U11684 (N_11684,N_11402,N_11018);
xor U11685 (N_11685,N_11449,N_11240);
nor U11686 (N_11686,N_11252,N_11489);
and U11687 (N_11687,N_11113,N_11390);
or U11688 (N_11688,N_11250,N_11209);
nor U11689 (N_11689,N_11025,N_11177);
and U11690 (N_11690,N_11414,N_11161);
xor U11691 (N_11691,N_11315,N_11272);
nand U11692 (N_11692,N_11128,N_11086);
or U11693 (N_11693,N_11383,N_11023);
or U11694 (N_11694,N_11207,N_11254);
nor U11695 (N_11695,N_11330,N_11176);
nor U11696 (N_11696,N_11036,N_11251);
xor U11697 (N_11697,N_11160,N_11302);
and U11698 (N_11698,N_11085,N_11001);
nor U11699 (N_11699,N_11019,N_11088);
xor U11700 (N_11700,N_11117,N_11495);
xor U11701 (N_11701,N_11061,N_11290);
xnor U11702 (N_11702,N_11031,N_11196);
and U11703 (N_11703,N_11351,N_11304);
xnor U11704 (N_11704,N_11341,N_11139);
or U11705 (N_11705,N_11194,N_11283);
nand U11706 (N_11706,N_11363,N_11320);
nand U11707 (N_11707,N_11050,N_11122);
nand U11708 (N_11708,N_11472,N_11227);
nand U11709 (N_11709,N_11233,N_11035);
or U11710 (N_11710,N_11369,N_11482);
or U11711 (N_11711,N_11210,N_11348);
xor U11712 (N_11712,N_11185,N_11485);
xnor U11713 (N_11713,N_11028,N_11084);
nor U11714 (N_11714,N_11286,N_11095);
nand U11715 (N_11715,N_11092,N_11285);
xnor U11716 (N_11716,N_11317,N_11120);
and U11717 (N_11717,N_11266,N_11499);
xnor U11718 (N_11718,N_11417,N_11073);
and U11719 (N_11719,N_11178,N_11090);
and U11720 (N_11720,N_11440,N_11392);
or U11721 (N_11721,N_11284,N_11410);
nor U11722 (N_11722,N_11216,N_11267);
and U11723 (N_11723,N_11214,N_11238);
and U11724 (N_11724,N_11277,N_11026);
xor U11725 (N_11725,N_11471,N_11097);
xor U11726 (N_11726,N_11012,N_11374);
nor U11727 (N_11727,N_11388,N_11037);
or U11728 (N_11728,N_11355,N_11278);
and U11729 (N_11729,N_11204,N_11394);
nor U11730 (N_11730,N_11331,N_11155);
nor U11731 (N_11731,N_11340,N_11300);
nor U11732 (N_11732,N_11282,N_11367);
xnor U11733 (N_11733,N_11137,N_11437);
nor U11734 (N_11734,N_11020,N_11397);
nand U11735 (N_11735,N_11136,N_11321);
nand U11736 (N_11736,N_11426,N_11451);
nand U11737 (N_11737,N_11232,N_11468);
xnor U11738 (N_11738,N_11157,N_11368);
xnor U11739 (N_11739,N_11189,N_11393);
nor U11740 (N_11740,N_11301,N_11441);
and U11741 (N_11741,N_11362,N_11418);
and U11742 (N_11742,N_11075,N_11065);
and U11743 (N_11743,N_11005,N_11462);
and U11744 (N_11744,N_11447,N_11476);
or U11745 (N_11745,N_11371,N_11007);
and U11746 (N_11746,N_11226,N_11244);
and U11747 (N_11747,N_11125,N_11104);
nand U11748 (N_11748,N_11327,N_11243);
nand U11749 (N_11749,N_11107,N_11024);
nor U11750 (N_11750,N_11459,N_11195);
xor U11751 (N_11751,N_11330,N_11132);
nor U11752 (N_11752,N_11266,N_11076);
nand U11753 (N_11753,N_11465,N_11289);
xor U11754 (N_11754,N_11084,N_11196);
or U11755 (N_11755,N_11441,N_11458);
xnor U11756 (N_11756,N_11494,N_11054);
nand U11757 (N_11757,N_11315,N_11056);
xnor U11758 (N_11758,N_11209,N_11054);
nand U11759 (N_11759,N_11139,N_11162);
nand U11760 (N_11760,N_11073,N_11155);
nor U11761 (N_11761,N_11275,N_11433);
and U11762 (N_11762,N_11443,N_11362);
nor U11763 (N_11763,N_11125,N_11143);
or U11764 (N_11764,N_11020,N_11481);
nor U11765 (N_11765,N_11007,N_11312);
nor U11766 (N_11766,N_11469,N_11319);
xor U11767 (N_11767,N_11304,N_11407);
nand U11768 (N_11768,N_11330,N_11140);
xor U11769 (N_11769,N_11278,N_11291);
and U11770 (N_11770,N_11429,N_11075);
nor U11771 (N_11771,N_11242,N_11385);
xnor U11772 (N_11772,N_11166,N_11438);
nand U11773 (N_11773,N_11487,N_11356);
and U11774 (N_11774,N_11346,N_11415);
and U11775 (N_11775,N_11319,N_11401);
nor U11776 (N_11776,N_11484,N_11175);
or U11777 (N_11777,N_11283,N_11129);
nor U11778 (N_11778,N_11393,N_11303);
nor U11779 (N_11779,N_11263,N_11097);
or U11780 (N_11780,N_11016,N_11317);
and U11781 (N_11781,N_11265,N_11053);
or U11782 (N_11782,N_11057,N_11270);
or U11783 (N_11783,N_11461,N_11336);
xor U11784 (N_11784,N_11434,N_11445);
or U11785 (N_11785,N_11287,N_11453);
or U11786 (N_11786,N_11497,N_11454);
and U11787 (N_11787,N_11475,N_11477);
xor U11788 (N_11788,N_11045,N_11199);
nand U11789 (N_11789,N_11271,N_11233);
or U11790 (N_11790,N_11029,N_11098);
nand U11791 (N_11791,N_11349,N_11469);
xor U11792 (N_11792,N_11254,N_11099);
xor U11793 (N_11793,N_11465,N_11085);
nor U11794 (N_11794,N_11365,N_11298);
or U11795 (N_11795,N_11407,N_11488);
nand U11796 (N_11796,N_11194,N_11070);
nand U11797 (N_11797,N_11043,N_11112);
xnor U11798 (N_11798,N_11085,N_11029);
nor U11799 (N_11799,N_11024,N_11457);
nor U11800 (N_11800,N_11106,N_11126);
nand U11801 (N_11801,N_11359,N_11192);
nor U11802 (N_11802,N_11198,N_11465);
or U11803 (N_11803,N_11008,N_11490);
nor U11804 (N_11804,N_11384,N_11271);
xnor U11805 (N_11805,N_11022,N_11441);
nor U11806 (N_11806,N_11309,N_11122);
or U11807 (N_11807,N_11385,N_11030);
and U11808 (N_11808,N_11243,N_11098);
or U11809 (N_11809,N_11185,N_11059);
nand U11810 (N_11810,N_11049,N_11089);
nor U11811 (N_11811,N_11029,N_11287);
nor U11812 (N_11812,N_11194,N_11476);
nor U11813 (N_11813,N_11334,N_11058);
xnor U11814 (N_11814,N_11025,N_11054);
xor U11815 (N_11815,N_11247,N_11319);
and U11816 (N_11816,N_11073,N_11493);
nand U11817 (N_11817,N_11291,N_11056);
and U11818 (N_11818,N_11228,N_11387);
nor U11819 (N_11819,N_11445,N_11366);
xnor U11820 (N_11820,N_11045,N_11043);
nor U11821 (N_11821,N_11194,N_11444);
and U11822 (N_11822,N_11119,N_11350);
nand U11823 (N_11823,N_11028,N_11160);
nand U11824 (N_11824,N_11423,N_11402);
xnor U11825 (N_11825,N_11209,N_11225);
xnor U11826 (N_11826,N_11498,N_11311);
nor U11827 (N_11827,N_11395,N_11036);
and U11828 (N_11828,N_11447,N_11383);
and U11829 (N_11829,N_11303,N_11183);
xnor U11830 (N_11830,N_11031,N_11345);
xnor U11831 (N_11831,N_11227,N_11123);
nand U11832 (N_11832,N_11077,N_11446);
or U11833 (N_11833,N_11219,N_11302);
and U11834 (N_11834,N_11226,N_11007);
xnor U11835 (N_11835,N_11225,N_11105);
nand U11836 (N_11836,N_11221,N_11000);
and U11837 (N_11837,N_11035,N_11450);
xnor U11838 (N_11838,N_11330,N_11154);
nand U11839 (N_11839,N_11399,N_11421);
or U11840 (N_11840,N_11385,N_11391);
xor U11841 (N_11841,N_11134,N_11211);
or U11842 (N_11842,N_11480,N_11151);
and U11843 (N_11843,N_11406,N_11478);
nor U11844 (N_11844,N_11044,N_11233);
and U11845 (N_11845,N_11074,N_11089);
or U11846 (N_11846,N_11323,N_11283);
and U11847 (N_11847,N_11217,N_11281);
or U11848 (N_11848,N_11093,N_11396);
and U11849 (N_11849,N_11179,N_11156);
or U11850 (N_11850,N_11112,N_11099);
or U11851 (N_11851,N_11292,N_11315);
nand U11852 (N_11852,N_11402,N_11496);
nand U11853 (N_11853,N_11117,N_11317);
or U11854 (N_11854,N_11276,N_11350);
and U11855 (N_11855,N_11436,N_11206);
nand U11856 (N_11856,N_11318,N_11371);
nand U11857 (N_11857,N_11384,N_11096);
nor U11858 (N_11858,N_11064,N_11235);
or U11859 (N_11859,N_11318,N_11115);
xor U11860 (N_11860,N_11392,N_11314);
nor U11861 (N_11861,N_11225,N_11219);
or U11862 (N_11862,N_11315,N_11407);
nand U11863 (N_11863,N_11262,N_11097);
nor U11864 (N_11864,N_11155,N_11408);
nor U11865 (N_11865,N_11226,N_11431);
and U11866 (N_11866,N_11136,N_11484);
or U11867 (N_11867,N_11248,N_11489);
nor U11868 (N_11868,N_11063,N_11234);
xnor U11869 (N_11869,N_11401,N_11248);
nor U11870 (N_11870,N_11074,N_11433);
xnor U11871 (N_11871,N_11137,N_11491);
and U11872 (N_11872,N_11221,N_11014);
nor U11873 (N_11873,N_11450,N_11240);
nand U11874 (N_11874,N_11098,N_11494);
and U11875 (N_11875,N_11071,N_11096);
nand U11876 (N_11876,N_11023,N_11156);
nor U11877 (N_11877,N_11328,N_11189);
and U11878 (N_11878,N_11106,N_11329);
nor U11879 (N_11879,N_11201,N_11067);
and U11880 (N_11880,N_11205,N_11035);
xor U11881 (N_11881,N_11407,N_11325);
and U11882 (N_11882,N_11096,N_11309);
nand U11883 (N_11883,N_11308,N_11451);
nand U11884 (N_11884,N_11235,N_11200);
and U11885 (N_11885,N_11275,N_11063);
and U11886 (N_11886,N_11436,N_11003);
or U11887 (N_11887,N_11243,N_11279);
nor U11888 (N_11888,N_11474,N_11096);
or U11889 (N_11889,N_11053,N_11413);
and U11890 (N_11890,N_11365,N_11491);
and U11891 (N_11891,N_11183,N_11190);
xor U11892 (N_11892,N_11099,N_11113);
nor U11893 (N_11893,N_11292,N_11346);
xor U11894 (N_11894,N_11165,N_11015);
or U11895 (N_11895,N_11276,N_11120);
xor U11896 (N_11896,N_11156,N_11243);
xor U11897 (N_11897,N_11260,N_11430);
nor U11898 (N_11898,N_11269,N_11341);
xor U11899 (N_11899,N_11275,N_11420);
nand U11900 (N_11900,N_11218,N_11332);
nand U11901 (N_11901,N_11026,N_11131);
xor U11902 (N_11902,N_11414,N_11072);
or U11903 (N_11903,N_11429,N_11133);
nand U11904 (N_11904,N_11351,N_11442);
nand U11905 (N_11905,N_11281,N_11377);
or U11906 (N_11906,N_11224,N_11461);
and U11907 (N_11907,N_11179,N_11146);
xor U11908 (N_11908,N_11326,N_11491);
or U11909 (N_11909,N_11074,N_11461);
xor U11910 (N_11910,N_11381,N_11011);
xnor U11911 (N_11911,N_11270,N_11281);
nor U11912 (N_11912,N_11038,N_11059);
nand U11913 (N_11913,N_11096,N_11046);
or U11914 (N_11914,N_11200,N_11009);
and U11915 (N_11915,N_11063,N_11427);
nor U11916 (N_11916,N_11042,N_11021);
and U11917 (N_11917,N_11086,N_11038);
xnor U11918 (N_11918,N_11095,N_11353);
and U11919 (N_11919,N_11231,N_11362);
xor U11920 (N_11920,N_11011,N_11497);
xor U11921 (N_11921,N_11114,N_11416);
nor U11922 (N_11922,N_11017,N_11231);
and U11923 (N_11923,N_11416,N_11492);
and U11924 (N_11924,N_11183,N_11401);
and U11925 (N_11925,N_11303,N_11268);
xnor U11926 (N_11926,N_11482,N_11133);
or U11927 (N_11927,N_11317,N_11436);
nand U11928 (N_11928,N_11489,N_11237);
and U11929 (N_11929,N_11445,N_11357);
or U11930 (N_11930,N_11127,N_11215);
xnor U11931 (N_11931,N_11265,N_11499);
and U11932 (N_11932,N_11079,N_11000);
nand U11933 (N_11933,N_11054,N_11168);
nand U11934 (N_11934,N_11182,N_11474);
or U11935 (N_11935,N_11092,N_11475);
nand U11936 (N_11936,N_11334,N_11140);
xnor U11937 (N_11937,N_11433,N_11341);
xor U11938 (N_11938,N_11045,N_11463);
or U11939 (N_11939,N_11132,N_11451);
or U11940 (N_11940,N_11090,N_11285);
nand U11941 (N_11941,N_11229,N_11483);
or U11942 (N_11942,N_11230,N_11485);
xnor U11943 (N_11943,N_11212,N_11056);
nand U11944 (N_11944,N_11208,N_11175);
or U11945 (N_11945,N_11014,N_11402);
or U11946 (N_11946,N_11199,N_11284);
or U11947 (N_11947,N_11298,N_11415);
nand U11948 (N_11948,N_11325,N_11374);
and U11949 (N_11949,N_11111,N_11247);
xor U11950 (N_11950,N_11025,N_11316);
nor U11951 (N_11951,N_11296,N_11064);
xor U11952 (N_11952,N_11377,N_11016);
xnor U11953 (N_11953,N_11397,N_11400);
xor U11954 (N_11954,N_11122,N_11281);
nor U11955 (N_11955,N_11200,N_11092);
and U11956 (N_11956,N_11442,N_11053);
and U11957 (N_11957,N_11310,N_11133);
xor U11958 (N_11958,N_11318,N_11460);
nand U11959 (N_11959,N_11237,N_11186);
or U11960 (N_11960,N_11305,N_11201);
xor U11961 (N_11961,N_11395,N_11351);
xor U11962 (N_11962,N_11019,N_11114);
nand U11963 (N_11963,N_11004,N_11054);
and U11964 (N_11964,N_11237,N_11005);
and U11965 (N_11965,N_11111,N_11185);
and U11966 (N_11966,N_11028,N_11451);
and U11967 (N_11967,N_11323,N_11004);
nor U11968 (N_11968,N_11117,N_11087);
and U11969 (N_11969,N_11494,N_11176);
xnor U11970 (N_11970,N_11204,N_11376);
nor U11971 (N_11971,N_11226,N_11137);
xnor U11972 (N_11972,N_11014,N_11258);
xnor U11973 (N_11973,N_11027,N_11475);
and U11974 (N_11974,N_11151,N_11259);
or U11975 (N_11975,N_11384,N_11211);
or U11976 (N_11976,N_11107,N_11283);
nor U11977 (N_11977,N_11230,N_11114);
nor U11978 (N_11978,N_11312,N_11101);
nor U11979 (N_11979,N_11254,N_11471);
or U11980 (N_11980,N_11363,N_11368);
nand U11981 (N_11981,N_11474,N_11311);
or U11982 (N_11982,N_11157,N_11017);
nor U11983 (N_11983,N_11235,N_11344);
xnor U11984 (N_11984,N_11067,N_11134);
and U11985 (N_11985,N_11377,N_11105);
nor U11986 (N_11986,N_11118,N_11238);
or U11987 (N_11987,N_11382,N_11362);
and U11988 (N_11988,N_11235,N_11382);
and U11989 (N_11989,N_11139,N_11048);
nand U11990 (N_11990,N_11122,N_11214);
or U11991 (N_11991,N_11296,N_11058);
xor U11992 (N_11992,N_11257,N_11424);
nand U11993 (N_11993,N_11155,N_11388);
nand U11994 (N_11994,N_11265,N_11187);
or U11995 (N_11995,N_11351,N_11197);
nand U11996 (N_11996,N_11180,N_11061);
nor U11997 (N_11997,N_11460,N_11445);
xnor U11998 (N_11998,N_11274,N_11195);
xnor U11999 (N_11999,N_11363,N_11010);
nor U12000 (N_12000,N_11554,N_11714);
and U12001 (N_12001,N_11608,N_11767);
and U12002 (N_12002,N_11669,N_11974);
or U12003 (N_12003,N_11566,N_11986);
nor U12004 (N_12004,N_11754,N_11826);
or U12005 (N_12005,N_11970,N_11645);
and U12006 (N_12006,N_11635,N_11910);
or U12007 (N_12007,N_11958,N_11768);
nand U12008 (N_12008,N_11618,N_11581);
xor U12009 (N_12009,N_11877,N_11980);
and U12010 (N_12010,N_11903,N_11819);
and U12011 (N_12011,N_11967,N_11579);
xor U12012 (N_12012,N_11756,N_11926);
xor U12013 (N_12013,N_11884,N_11510);
nand U12014 (N_12014,N_11898,N_11622);
xnor U12015 (N_12015,N_11874,N_11744);
nand U12016 (N_12016,N_11842,N_11868);
nand U12017 (N_12017,N_11969,N_11503);
xnor U12018 (N_12018,N_11987,N_11782);
nand U12019 (N_12019,N_11586,N_11611);
or U12020 (N_12020,N_11810,N_11585);
nor U12021 (N_12021,N_11869,N_11847);
and U12022 (N_12022,N_11808,N_11989);
nor U12023 (N_12023,N_11929,N_11781);
and U12024 (N_12024,N_11730,N_11706);
or U12025 (N_12025,N_11905,N_11511);
nor U12026 (N_12026,N_11801,N_11515);
and U12027 (N_12027,N_11615,N_11594);
and U12028 (N_12028,N_11569,N_11994);
xor U12029 (N_12029,N_11843,N_11512);
nor U12030 (N_12030,N_11750,N_11889);
nand U12031 (N_12031,N_11549,N_11770);
nand U12032 (N_12032,N_11933,N_11671);
xnor U12033 (N_12033,N_11794,N_11605);
nor U12034 (N_12034,N_11942,N_11673);
and U12035 (N_12035,N_11733,N_11598);
or U12036 (N_12036,N_11923,N_11651);
nor U12037 (N_12037,N_11878,N_11500);
nor U12038 (N_12038,N_11864,N_11590);
nand U12039 (N_12039,N_11735,N_11901);
nand U12040 (N_12040,N_11865,N_11725);
nor U12041 (N_12041,N_11998,N_11678);
and U12042 (N_12042,N_11906,N_11856);
nor U12043 (N_12043,N_11857,N_11659);
xor U12044 (N_12044,N_11961,N_11576);
or U12045 (N_12045,N_11976,N_11666);
nor U12046 (N_12046,N_11711,N_11578);
xor U12047 (N_12047,N_11891,N_11621);
or U12048 (N_12048,N_11841,N_11792);
and U12049 (N_12049,N_11939,N_11979);
and U12050 (N_12050,N_11649,N_11648);
or U12051 (N_12051,N_11936,N_11596);
xnor U12052 (N_12052,N_11778,N_11944);
or U12053 (N_12053,N_11997,N_11604);
nand U12054 (N_12054,N_11551,N_11981);
xor U12055 (N_12055,N_11812,N_11928);
or U12056 (N_12056,N_11930,N_11881);
nand U12057 (N_12057,N_11860,N_11769);
nor U12058 (N_12058,N_11946,N_11716);
nor U12059 (N_12059,N_11544,N_11802);
nor U12060 (N_12060,N_11836,N_11825);
or U12061 (N_12061,N_11813,N_11971);
and U12062 (N_12062,N_11870,N_11624);
nor U12063 (N_12063,N_11740,N_11727);
nor U12064 (N_12064,N_11720,N_11952);
nor U12065 (N_12065,N_11527,N_11589);
or U12066 (N_12066,N_11831,N_11746);
and U12067 (N_12067,N_11811,N_11762);
or U12068 (N_12068,N_11751,N_11823);
and U12069 (N_12069,N_11888,N_11682);
xor U12070 (N_12070,N_11504,N_11924);
or U12071 (N_12071,N_11820,N_11885);
or U12072 (N_12072,N_11815,N_11827);
or U12073 (N_12073,N_11690,N_11887);
nand U12074 (N_12074,N_11845,N_11630);
nand U12075 (N_12075,N_11873,N_11797);
or U12076 (N_12076,N_11639,N_11966);
nor U12077 (N_12077,N_11691,N_11636);
nand U12078 (N_12078,N_11695,N_11776);
xnor U12079 (N_12079,N_11814,N_11684);
or U12080 (N_12080,N_11713,N_11851);
or U12081 (N_12081,N_11916,N_11686);
and U12082 (N_12082,N_11542,N_11818);
nor U12083 (N_12083,N_11940,N_11859);
nand U12084 (N_12084,N_11817,N_11988);
xnor U12085 (N_12085,N_11623,N_11644);
and U12086 (N_12086,N_11722,N_11795);
nor U12087 (N_12087,N_11900,N_11600);
nand U12088 (N_12088,N_11753,N_11726);
xor U12089 (N_12089,N_11652,N_11657);
or U12090 (N_12090,N_11588,N_11587);
nand U12091 (N_12091,N_11517,N_11546);
nand U12092 (N_12092,N_11743,N_11862);
xor U12093 (N_12093,N_11573,N_11556);
nor U12094 (N_12094,N_11632,N_11591);
xnor U12095 (N_12095,N_11800,N_11915);
xnor U12096 (N_12096,N_11687,N_11723);
and U12097 (N_12097,N_11634,N_11766);
or U12098 (N_12098,N_11833,N_11858);
xor U12099 (N_12099,N_11890,N_11736);
xnor U12100 (N_12100,N_11982,N_11922);
or U12101 (N_12101,N_11852,N_11925);
or U12102 (N_12102,N_11934,N_11755);
nor U12103 (N_12103,N_11559,N_11627);
and U12104 (N_12104,N_11734,N_11547);
nor U12105 (N_12105,N_11675,N_11731);
nor U12106 (N_12106,N_11507,N_11646);
or U12107 (N_12107,N_11995,N_11724);
and U12108 (N_12108,N_11759,N_11880);
nor U12109 (N_12109,N_11583,N_11502);
and U12110 (N_12110,N_11879,N_11777);
nor U12111 (N_12111,N_11528,N_11564);
nand U12112 (N_12112,N_11787,N_11533);
xnor U12113 (N_12113,N_11899,N_11747);
or U12114 (N_12114,N_11863,N_11830);
and U12115 (N_12115,N_11990,N_11592);
nor U12116 (N_12116,N_11702,N_11893);
or U12117 (N_12117,N_11809,N_11530);
and U12118 (N_12118,N_11543,N_11805);
xor U12119 (N_12119,N_11670,N_11892);
and U12120 (N_12120,N_11793,N_11718);
or U12121 (N_12121,N_11577,N_11558);
or U12122 (N_12122,N_11665,N_11779);
nor U12123 (N_12123,N_11717,N_11653);
nor U12124 (N_12124,N_11571,N_11699);
and U12125 (N_12125,N_11949,N_11532);
or U12126 (N_12126,N_11774,N_11513);
or U12127 (N_12127,N_11752,N_11927);
and U12128 (N_12128,N_11791,N_11835);
xor U12129 (N_12129,N_11745,N_11919);
or U12130 (N_12130,N_11710,N_11701);
or U12131 (N_12131,N_11999,N_11692);
xnor U12132 (N_12132,N_11932,N_11968);
or U12133 (N_12133,N_11786,N_11957);
xnor U12134 (N_12134,N_11975,N_11696);
or U12135 (N_12135,N_11937,N_11788);
xor U12136 (N_12136,N_11822,N_11943);
or U12137 (N_12137,N_11790,N_11620);
and U12138 (N_12138,N_11655,N_11662);
and U12139 (N_12139,N_11693,N_11563);
nand U12140 (N_12140,N_11954,N_11575);
nand U12141 (N_12141,N_11894,N_11535);
and U12142 (N_12142,N_11829,N_11896);
or U12143 (N_12143,N_11629,N_11626);
and U12144 (N_12144,N_11610,N_11920);
and U12145 (N_12145,N_11522,N_11738);
nor U12146 (N_12146,N_11828,N_11694);
nand U12147 (N_12147,N_11850,N_11667);
and U12148 (N_12148,N_11789,N_11548);
nand U12149 (N_12149,N_11509,N_11647);
or U12150 (N_12150,N_11561,N_11913);
or U12151 (N_12151,N_11712,N_11875);
and U12152 (N_12152,N_11601,N_11703);
xnor U12153 (N_12153,N_11617,N_11984);
or U12154 (N_12154,N_11628,N_11876);
or U12155 (N_12155,N_11978,N_11848);
xnor U12156 (N_12156,N_11908,N_11992);
nor U12157 (N_12157,N_11796,N_11947);
or U12158 (N_12158,N_11593,N_11758);
and U12159 (N_12159,N_11640,N_11807);
and U12160 (N_12160,N_11824,N_11973);
or U12161 (N_12161,N_11541,N_11506);
nand U12162 (N_12162,N_11685,N_11698);
nand U12163 (N_12163,N_11965,N_11638);
nand U12164 (N_12164,N_11689,N_11519);
or U12165 (N_12165,N_11945,N_11902);
nor U12166 (N_12166,N_11516,N_11853);
nand U12167 (N_12167,N_11705,N_11839);
and U12168 (N_12168,N_11572,N_11545);
or U12169 (N_12169,N_11721,N_11804);
nor U12170 (N_12170,N_11597,N_11505);
xor U12171 (N_12171,N_11911,N_11642);
nand U12172 (N_12172,N_11524,N_11763);
and U12173 (N_12173,N_11964,N_11707);
nand U12174 (N_12174,N_11668,N_11904);
nand U12175 (N_12175,N_11501,N_11637);
xor U12176 (N_12176,N_11658,N_11799);
and U12177 (N_12177,N_11606,N_11948);
or U12178 (N_12178,N_11959,N_11536);
xnor U12179 (N_12179,N_11508,N_11538);
and U12180 (N_12180,N_11709,N_11599);
nand U12181 (N_12181,N_11914,N_11977);
nor U12182 (N_12182,N_11681,N_11614);
nand U12183 (N_12183,N_11676,N_11663);
nand U12184 (N_12184,N_11855,N_11708);
xor U12185 (N_12185,N_11729,N_11951);
xor U12186 (N_12186,N_11909,N_11895);
nor U12187 (N_12187,N_11741,N_11938);
and U12188 (N_12188,N_11785,N_11749);
nor U12189 (N_12189,N_11531,N_11772);
nand U12190 (N_12190,N_11872,N_11775);
and U12191 (N_12191,N_11907,N_11764);
and U12192 (N_12192,N_11540,N_11742);
and U12193 (N_12193,N_11560,N_11631);
or U12194 (N_12194,N_11567,N_11683);
and U12195 (N_12195,N_11871,N_11866);
or U12196 (N_12196,N_11521,N_11941);
or U12197 (N_12197,N_11518,N_11897);
and U12198 (N_12198,N_11595,N_11837);
nand U12199 (N_12199,N_11728,N_11867);
nand U12200 (N_12200,N_11704,N_11565);
xor U12201 (N_12201,N_11960,N_11529);
xor U12202 (N_12202,N_11962,N_11921);
xor U12203 (N_12203,N_11650,N_11854);
xnor U12204 (N_12204,N_11672,N_11955);
xnor U12205 (N_12205,N_11570,N_11643);
or U12206 (N_12206,N_11582,N_11816);
nand U12207 (N_12207,N_11514,N_11568);
and U12208 (N_12208,N_11846,N_11553);
nor U12209 (N_12209,N_11688,N_11613);
or U12210 (N_12210,N_11539,N_11748);
or U12211 (N_12211,N_11771,N_11537);
nor U12212 (N_12212,N_11654,N_11803);
xnor U12213 (N_12213,N_11765,N_11950);
or U12214 (N_12214,N_11523,N_11983);
nor U12215 (N_12215,N_11991,N_11562);
xor U12216 (N_12216,N_11520,N_11737);
or U12217 (N_12217,N_11773,N_11840);
nor U12218 (N_12218,N_11534,N_11660);
nor U12219 (N_12219,N_11700,N_11739);
or U12220 (N_12220,N_11918,N_11697);
or U12221 (N_12221,N_11580,N_11732);
or U12222 (N_12222,N_11935,N_11844);
xnor U12223 (N_12223,N_11761,N_11525);
xnor U12224 (N_12224,N_11757,N_11719);
or U12225 (N_12225,N_11607,N_11625);
nor U12226 (N_12226,N_11526,N_11886);
nand U12227 (N_12227,N_11806,N_11832);
nor U12228 (N_12228,N_11656,N_11555);
and U12229 (N_12229,N_11760,N_11674);
nand U12230 (N_12230,N_11912,N_11963);
xnor U12231 (N_12231,N_11633,N_11882);
nor U12232 (N_12232,N_11609,N_11784);
nor U12233 (N_12233,N_11616,N_11641);
or U12234 (N_12234,N_11550,N_11552);
nand U12235 (N_12235,N_11996,N_11783);
and U12236 (N_12236,N_11664,N_11677);
or U12237 (N_12237,N_11849,N_11993);
nand U12238 (N_12238,N_11557,N_11715);
nand U12239 (N_12239,N_11953,N_11680);
nand U12240 (N_12240,N_11834,N_11619);
nand U12241 (N_12241,N_11956,N_11584);
and U12242 (N_12242,N_11780,N_11603);
or U12243 (N_12243,N_11821,N_11917);
nand U12244 (N_12244,N_11838,N_11602);
and U12245 (N_12245,N_11612,N_11861);
and U12246 (N_12246,N_11661,N_11574);
or U12247 (N_12247,N_11972,N_11931);
nor U12248 (N_12248,N_11679,N_11798);
xor U12249 (N_12249,N_11883,N_11985);
nand U12250 (N_12250,N_11929,N_11941);
nand U12251 (N_12251,N_11807,N_11596);
xor U12252 (N_12252,N_11566,N_11625);
or U12253 (N_12253,N_11510,N_11667);
or U12254 (N_12254,N_11756,N_11750);
and U12255 (N_12255,N_11514,N_11639);
xor U12256 (N_12256,N_11558,N_11991);
nand U12257 (N_12257,N_11729,N_11589);
and U12258 (N_12258,N_11546,N_11763);
or U12259 (N_12259,N_11827,N_11874);
nand U12260 (N_12260,N_11555,N_11536);
or U12261 (N_12261,N_11749,N_11730);
or U12262 (N_12262,N_11583,N_11558);
or U12263 (N_12263,N_11672,N_11751);
nor U12264 (N_12264,N_11626,N_11896);
nor U12265 (N_12265,N_11886,N_11950);
or U12266 (N_12266,N_11874,N_11701);
nand U12267 (N_12267,N_11763,N_11843);
or U12268 (N_12268,N_11835,N_11508);
and U12269 (N_12269,N_11696,N_11785);
and U12270 (N_12270,N_11689,N_11543);
xnor U12271 (N_12271,N_11924,N_11936);
xnor U12272 (N_12272,N_11949,N_11685);
or U12273 (N_12273,N_11664,N_11943);
and U12274 (N_12274,N_11828,N_11653);
nand U12275 (N_12275,N_11914,N_11894);
nor U12276 (N_12276,N_11584,N_11854);
or U12277 (N_12277,N_11614,N_11536);
xnor U12278 (N_12278,N_11983,N_11532);
and U12279 (N_12279,N_11503,N_11570);
or U12280 (N_12280,N_11979,N_11502);
and U12281 (N_12281,N_11861,N_11740);
xor U12282 (N_12282,N_11764,N_11560);
nand U12283 (N_12283,N_11942,N_11513);
and U12284 (N_12284,N_11500,N_11550);
nor U12285 (N_12285,N_11970,N_11848);
nand U12286 (N_12286,N_11681,N_11941);
nor U12287 (N_12287,N_11626,N_11715);
nand U12288 (N_12288,N_11637,N_11705);
nor U12289 (N_12289,N_11654,N_11728);
nor U12290 (N_12290,N_11692,N_11983);
nor U12291 (N_12291,N_11820,N_11863);
nand U12292 (N_12292,N_11701,N_11628);
nand U12293 (N_12293,N_11653,N_11997);
xor U12294 (N_12294,N_11664,N_11583);
nand U12295 (N_12295,N_11969,N_11625);
and U12296 (N_12296,N_11986,N_11665);
xnor U12297 (N_12297,N_11939,N_11585);
or U12298 (N_12298,N_11851,N_11561);
nor U12299 (N_12299,N_11608,N_11805);
or U12300 (N_12300,N_11746,N_11689);
xnor U12301 (N_12301,N_11727,N_11826);
and U12302 (N_12302,N_11782,N_11543);
nand U12303 (N_12303,N_11895,N_11814);
nand U12304 (N_12304,N_11839,N_11764);
xnor U12305 (N_12305,N_11526,N_11586);
xnor U12306 (N_12306,N_11643,N_11773);
nand U12307 (N_12307,N_11994,N_11879);
and U12308 (N_12308,N_11822,N_11635);
and U12309 (N_12309,N_11603,N_11524);
xnor U12310 (N_12310,N_11848,N_11836);
nor U12311 (N_12311,N_11988,N_11720);
or U12312 (N_12312,N_11764,N_11589);
nor U12313 (N_12313,N_11621,N_11553);
and U12314 (N_12314,N_11662,N_11835);
nor U12315 (N_12315,N_11873,N_11670);
xor U12316 (N_12316,N_11925,N_11709);
and U12317 (N_12317,N_11811,N_11851);
nand U12318 (N_12318,N_11979,N_11840);
or U12319 (N_12319,N_11891,N_11836);
nand U12320 (N_12320,N_11545,N_11863);
nand U12321 (N_12321,N_11675,N_11501);
or U12322 (N_12322,N_11773,N_11609);
xnor U12323 (N_12323,N_11913,N_11865);
or U12324 (N_12324,N_11699,N_11723);
and U12325 (N_12325,N_11798,N_11781);
xor U12326 (N_12326,N_11636,N_11876);
or U12327 (N_12327,N_11979,N_11500);
nor U12328 (N_12328,N_11749,N_11739);
xnor U12329 (N_12329,N_11514,N_11742);
or U12330 (N_12330,N_11667,N_11880);
or U12331 (N_12331,N_11573,N_11546);
nand U12332 (N_12332,N_11943,N_11614);
xor U12333 (N_12333,N_11933,N_11635);
and U12334 (N_12334,N_11551,N_11806);
or U12335 (N_12335,N_11634,N_11723);
xnor U12336 (N_12336,N_11790,N_11776);
nand U12337 (N_12337,N_11775,N_11802);
nand U12338 (N_12338,N_11541,N_11861);
and U12339 (N_12339,N_11686,N_11524);
and U12340 (N_12340,N_11930,N_11935);
xor U12341 (N_12341,N_11736,N_11620);
nor U12342 (N_12342,N_11571,N_11755);
nor U12343 (N_12343,N_11714,N_11812);
nor U12344 (N_12344,N_11508,N_11713);
nand U12345 (N_12345,N_11581,N_11823);
nand U12346 (N_12346,N_11816,N_11796);
nand U12347 (N_12347,N_11921,N_11844);
nor U12348 (N_12348,N_11504,N_11506);
and U12349 (N_12349,N_11922,N_11861);
xor U12350 (N_12350,N_11588,N_11510);
xor U12351 (N_12351,N_11606,N_11785);
nand U12352 (N_12352,N_11508,N_11624);
nand U12353 (N_12353,N_11667,N_11644);
and U12354 (N_12354,N_11802,N_11567);
nor U12355 (N_12355,N_11600,N_11505);
nor U12356 (N_12356,N_11861,N_11834);
nand U12357 (N_12357,N_11951,N_11507);
xor U12358 (N_12358,N_11677,N_11631);
nor U12359 (N_12359,N_11851,N_11723);
and U12360 (N_12360,N_11926,N_11572);
and U12361 (N_12361,N_11742,N_11907);
xor U12362 (N_12362,N_11568,N_11774);
and U12363 (N_12363,N_11645,N_11912);
xor U12364 (N_12364,N_11565,N_11699);
xnor U12365 (N_12365,N_11991,N_11755);
and U12366 (N_12366,N_11959,N_11574);
and U12367 (N_12367,N_11870,N_11750);
and U12368 (N_12368,N_11967,N_11551);
xnor U12369 (N_12369,N_11956,N_11560);
nand U12370 (N_12370,N_11973,N_11857);
or U12371 (N_12371,N_11808,N_11691);
nand U12372 (N_12372,N_11999,N_11804);
or U12373 (N_12373,N_11623,N_11942);
nand U12374 (N_12374,N_11629,N_11980);
or U12375 (N_12375,N_11786,N_11790);
or U12376 (N_12376,N_11904,N_11966);
and U12377 (N_12377,N_11920,N_11536);
xor U12378 (N_12378,N_11831,N_11850);
xnor U12379 (N_12379,N_11763,N_11620);
nand U12380 (N_12380,N_11918,N_11635);
or U12381 (N_12381,N_11822,N_11574);
nand U12382 (N_12382,N_11916,N_11895);
or U12383 (N_12383,N_11844,N_11636);
nand U12384 (N_12384,N_11838,N_11946);
nor U12385 (N_12385,N_11871,N_11569);
nand U12386 (N_12386,N_11788,N_11986);
or U12387 (N_12387,N_11828,N_11832);
or U12388 (N_12388,N_11976,N_11834);
nor U12389 (N_12389,N_11790,N_11506);
nand U12390 (N_12390,N_11902,N_11869);
nor U12391 (N_12391,N_11586,N_11857);
and U12392 (N_12392,N_11676,N_11922);
nand U12393 (N_12393,N_11551,N_11886);
nor U12394 (N_12394,N_11841,N_11668);
nand U12395 (N_12395,N_11505,N_11634);
xor U12396 (N_12396,N_11951,N_11975);
or U12397 (N_12397,N_11781,N_11502);
and U12398 (N_12398,N_11909,N_11894);
nor U12399 (N_12399,N_11939,N_11844);
nor U12400 (N_12400,N_11695,N_11574);
xnor U12401 (N_12401,N_11534,N_11804);
and U12402 (N_12402,N_11984,N_11915);
nand U12403 (N_12403,N_11814,N_11778);
or U12404 (N_12404,N_11635,N_11860);
nand U12405 (N_12405,N_11526,N_11756);
nand U12406 (N_12406,N_11728,N_11896);
xor U12407 (N_12407,N_11758,N_11608);
nor U12408 (N_12408,N_11631,N_11691);
xnor U12409 (N_12409,N_11715,N_11813);
xor U12410 (N_12410,N_11865,N_11763);
or U12411 (N_12411,N_11891,N_11945);
or U12412 (N_12412,N_11848,N_11742);
and U12413 (N_12413,N_11971,N_11966);
and U12414 (N_12414,N_11927,N_11517);
and U12415 (N_12415,N_11740,N_11519);
nand U12416 (N_12416,N_11805,N_11581);
nor U12417 (N_12417,N_11623,N_11996);
or U12418 (N_12418,N_11800,N_11775);
or U12419 (N_12419,N_11912,N_11734);
xor U12420 (N_12420,N_11902,N_11694);
and U12421 (N_12421,N_11889,N_11584);
and U12422 (N_12422,N_11904,N_11586);
nand U12423 (N_12423,N_11687,N_11565);
nand U12424 (N_12424,N_11851,N_11518);
nand U12425 (N_12425,N_11994,N_11792);
nor U12426 (N_12426,N_11919,N_11823);
or U12427 (N_12427,N_11594,N_11701);
nor U12428 (N_12428,N_11903,N_11747);
nor U12429 (N_12429,N_11923,N_11695);
nand U12430 (N_12430,N_11740,N_11922);
or U12431 (N_12431,N_11601,N_11794);
or U12432 (N_12432,N_11960,N_11586);
and U12433 (N_12433,N_11793,N_11897);
or U12434 (N_12434,N_11898,N_11700);
and U12435 (N_12435,N_11546,N_11883);
nand U12436 (N_12436,N_11789,N_11792);
and U12437 (N_12437,N_11756,N_11920);
xnor U12438 (N_12438,N_11703,N_11953);
xnor U12439 (N_12439,N_11580,N_11747);
and U12440 (N_12440,N_11556,N_11671);
or U12441 (N_12441,N_11958,N_11579);
nor U12442 (N_12442,N_11829,N_11855);
xnor U12443 (N_12443,N_11801,N_11708);
nor U12444 (N_12444,N_11920,N_11749);
xor U12445 (N_12445,N_11805,N_11975);
xnor U12446 (N_12446,N_11917,N_11584);
and U12447 (N_12447,N_11942,N_11616);
or U12448 (N_12448,N_11777,N_11900);
nor U12449 (N_12449,N_11707,N_11989);
and U12450 (N_12450,N_11758,N_11780);
and U12451 (N_12451,N_11674,N_11912);
xor U12452 (N_12452,N_11895,N_11775);
and U12453 (N_12453,N_11628,N_11845);
and U12454 (N_12454,N_11764,N_11629);
xor U12455 (N_12455,N_11918,N_11649);
or U12456 (N_12456,N_11773,N_11660);
nand U12457 (N_12457,N_11996,N_11630);
and U12458 (N_12458,N_11618,N_11749);
or U12459 (N_12459,N_11655,N_11809);
nor U12460 (N_12460,N_11716,N_11781);
and U12461 (N_12461,N_11734,N_11676);
xnor U12462 (N_12462,N_11800,N_11553);
and U12463 (N_12463,N_11802,N_11816);
nand U12464 (N_12464,N_11914,N_11834);
or U12465 (N_12465,N_11542,N_11846);
or U12466 (N_12466,N_11645,N_11980);
nand U12467 (N_12467,N_11883,N_11927);
nand U12468 (N_12468,N_11934,N_11581);
and U12469 (N_12469,N_11774,N_11523);
nand U12470 (N_12470,N_11568,N_11635);
xnor U12471 (N_12471,N_11821,N_11705);
or U12472 (N_12472,N_11671,N_11996);
and U12473 (N_12473,N_11929,N_11764);
nor U12474 (N_12474,N_11738,N_11893);
or U12475 (N_12475,N_11629,N_11608);
nor U12476 (N_12476,N_11728,N_11606);
nand U12477 (N_12477,N_11632,N_11737);
xnor U12478 (N_12478,N_11925,N_11986);
and U12479 (N_12479,N_11781,N_11743);
and U12480 (N_12480,N_11652,N_11722);
and U12481 (N_12481,N_11682,N_11533);
nand U12482 (N_12482,N_11667,N_11638);
and U12483 (N_12483,N_11753,N_11618);
or U12484 (N_12484,N_11951,N_11956);
or U12485 (N_12485,N_11773,N_11784);
nor U12486 (N_12486,N_11707,N_11547);
or U12487 (N_12487,N_11646,N_11953);
nor U12488 (N_12488,N_11774,N_11566);
or U12489 (N_12489,N_11712,N_11983);
xor U12490 (N_12490,N_11829,N_11740);
xor U12491 (N_12491,N_11971,N_11973);
and U12492 (N_12492,N_11668,N_11634);
and U12493 (N_12493,N_11823,N_11856);
xor U12494 (N_12494,N_11825,N_11923);
and U12495 (N_12495,N_11896,N_11584);
and U12496 (N_12496,N_11527,N_11978);
and U12497 (N_12497,N_11900,N_11955);
or U12498 (N_12498,N_11668,N_11769);
or U12499 (N_12499,N_11841,N_11900);
nand U12500 (N_12500,N_12293,N_12497);
and U12501 (N_12501,N_12418,N_12439);
and U12502 (N_12502,N_12208,N_12124);
and U12503 (N_12503,N_12481,N_12441);
or U12504 (N_12504,N_12318,N_12472);
or U12505 (N_12505,N_12456,N_12374);
and U12506 (N_12506,N_12494,N_12491);
or U12507 (N_12507,N_12368,N_12363);
xnor U12508 (N_12508,N_12273,N_12409);
or U12509 (N_12509,N_12181,N_12437);
xor U12510 (N_12510,N_12218,N_12005);
nor U12511 (N_12511,N_12394,N_12285);
and U12512 (N_12512,N_12268,N_12291);
and U12513 (N_12513,N_12463,N_12028);
or U12514 (N_12514,N_12294,N_12036);
nand U12515 (N_12515,N_12246,N_12050);
or U12516 (N_12516,N_12261,N_12323);
nor U12517 (N_12517,N_12142,N_12446);
nor U12518 (N_12518,N_12077,N_12373);
and U12519 (N_12519,N_12249,N_12467);
xor U12520 (N_12520,N_12328,N_12111);
and U12521 (N_12521,N_12358,N_12371);
nand U12522 (N_12522,N_12041,N_12287);
and U12523 (N_12523,N_12498,N_12023);
nand U12524 (N_12524,N_12019,N_12448);
and U12525 (N_12525,N_12134,N_12252);
nor U12526 (N_12526,N_12243,N_12039);
and U12527 (N_12527,N_12244,N_12392);
nor U12528 (N_12528,N_12359,N_12033);
or U12529 (N_12529,N_12277,N_12232);
xor U12530 (N_12530,N_12308,N_12049);
and U12531 (N_12531,N_12251,N_12304);
nand U12532 (N_12532,N_12337,N_12065);
nor U12533 (N_12533,N_12402,N_12298);
nor U12534 (N_12534,N_12344,N_12151);
and U12535 (N_12535,N_12201,N_12025);
and U12536 (N_12536,N_12235,N_12078);
nor U12537 (N_12537,N_12169,N_12297);
nand U12538 (N_12538,N_12132,N_12204);
nor U12539 (N_12539,N_12457,N_12450);
nand U12540 (N_12540,N_12461,N_12109);
and U12541 (N_12541,N_12495,N_12114);
nand U12542 (N_12542,N_12051,N_12205);
nor U12543 (N_12543,N_12014,N_12464);
nand U12544 (N_12544,N_12335,N_12168);
or U12545 (N_12545,N_12302,N_12061);
nand U12546 (N_12546,N_12037,N_12279);
and U12547 (N_12547,N_12237,N_12177);
and U12548 (N_12548,N_12343,N_12339);
and U12549 (N_12549,N_12329,N_12125);
nand U12550 (N_12550,N_12044,N_12367);
xnor U12551 (N_12551,N_12180,N_12471);
or U12552 (N_12552,N_12118,N_12390);
or U12553 (N_12553,N_12197,N_12216);
xor U12554 (N_12554,N_12121,N_12231);
nor U12555 (N_12555,N_12338,N_12452);
nor U12556 (N_12556,N_12191,N_12032);
and U12557 (N_12557,N_12454,N_12375);
nor U12558 (N_12558,N_12492,N_12012);
nand U12559 (N_12559,N_12095,N_12101);
nand U12560 (N_12560,N_12211,N_12444);
and U12561 (N_12561,N_12143,N_12021);
and U12562 (N_12562,N_12000,N_12099);
nor U12563 (N_12563,N_12364,N_12167);
xnor U12564 (N_12564,N_12391,N_12082);
xnor U12565 (N_12565,N_12440,N_12489);
nand U12566 (N_12566,N_12352,N_12372);
nor U12567 (N_12567,N_12434,N_12406);
xor U12568 (N_12568,N_12206,N_12228);
and U12569 (N_12569,N_12257,N_12163);
or U12570 (N_12570,N_12426,N_12160);
xnor U12571 (N_12571,N_12193,N_12239);
and U12572 (N_12572,N_12397,N_12284);
nand U12573 (N_12573,N_12320,N_12070);
nand U12574 (N_12574,N_12145,N_12186);
or U12575 (N_12575,N_12084,N_12135);
or U12576 (N_12576,N_12360,N_12350);
nand U12577 (N_12577,N_12332,N_12148);
nor U12578 (N_12578,N_12092,N_12274);
nor U12579 (N_12579,N_12477,N_12089);
or U12580 (N_12580,N_12133,N_12306);
nand U12581 (N_12581,N_12403,N_12241);
and U12582 (N_12582,N_12378,N_12140);
xnor U12583 (N_12583,N_12153,N_12131);
and U12584 (N_12584,N_12020,N_12264);
nand U12585 (N_12585,N_12333,N_12215);
nor U12586 (N_12586,N_12316,N_12233);
xnor U12587 (N_12587,N_12146,N_12071);
xnor U12588 (N_12588,N_12056,N_12093);
nand U12589 (N_12589,N_12183,N_12230);
xnor U12590 (N_12590,N_12016,N_12017);
or U12591 (N_12591,N_12399,N_12288);
xnor U12592 (N_12592,N_12433,N_12354);
nand U12593 (N_12593,N_12068,N_12384);
or U12594 (N_12594,N_12048,N_12010);
xnor U12595 (N_12595,N_12419,N_12485);
xor U12596 (N_12596,N_12415,N_12198);
nor U12597 (N_12597,N_12194,N_12057);
nor U12598 (N_12598,N_12094,N_12324);
nand U12599 (N_12599,N_12427,N_12214);
nand U12600 (N_12600,N_12238,N_12383);
nor U12601 (N_12601,N_12266,N_12296);
nand U12602 (N_12602,N_12362,N_12436);
xnor U12603 (N_12603,N_12240,N_12482);
nor U12604 (N_12604,N_12009,N_12468);
or U12605 (N_12605,N_12090,N_12281);
and U12606 (N_12606,N_12159,N_12203);
nor U12607 (N_12607,N_12270,N_12086);
and U12608 (N_12608,N_12120,N_12008);
or U12609 (N_12609,N_12263,N_12018);
nor U12610 (N_12610,N_12129,N_12073);
nor U12611 (N_12611,N_12227,N_12462);
or U12612 (N_12612,N_12007,N_12052);
nand U12613 (N_12613,N_12484,N_12283);
xnor U12614 (N_12614,N_12207,N_12262);
or U12615 (N_12615,N_12200,N_12490);
nand U12616 (N_12616,N_12024,N_12331);
or U12617 (N_12617,N_12040,N_12108);
and U12618 (N_12618,N_12385,N_12149);
nand U12619 (N_12619,N_12376,N_12002);
nor U12620 (N_12620,N_12387,N_12171);
nor U12621 (N_12621,N_12380,N_12189);
nor U12622 (N_12622,N_12496,N_12336);
xnor U12623 (N_12623,N_12074,N_12079);
xor U12624 (N_12624,N_12369,N_12414);
or U12625 (N_12625,N_12348,N_12217);
or U12626 (N_12626,N_12199,N_12451);
nand U12627 (N_12627,N_12345,N_12395);
nor U12628 (N_12628,N_12405,N_12098);
nor U12629 (N_12629,N_12123,N_12488);
or U12630 (N_12630,N_12001,N_12442);
xnor U12631 (N_12631,N_12493,N_12187);
or U12632 (N_12632,N_12110,N_12416);
nand U12633 (N_12633,N_12224,N_12299);
nand U12634 (N_12634,N_12470,N_12046);
nand U12635 (N_12635,N_12034,N_12213);
xor U12636 (N_12636,N_12340,N_12139);
nor U12637 (N_12637,N_12147,N_12280);
or U12638 (N_12638,N_12389,N_12355);
xor U12639 (N_12639,N_12478,N_12130);
nand U12640 (N_12640,N_12113,N_12062);
nor U12641 (N_12641,N_12404,N_12386);
or U12642 (N_12642,N_12388,N_12100);
or U12643 (N_12643,N_12413,N_12322);
nor U12644 (N_12644,N_12196,N_12236);
xnor U12645 (N_12645,N_12247,N_12043);
nand U12646 (N_12646,N_12072,N_12282);
nand U12647 (N_12647,N_12310,N_12104);
nand U12648 (N_12648,N_12253,N_12401);
and U12649 (N_12649,N_12170,N_12286);
or U12650 (N_12650,N_12311,N_12223);
xor U12651 (N_12651,N_12161,N_12222);
nand U12652 (N_12652,N_12487,N_12122);
nand U12653 (N_12653,N_12410,N_12212);
or U12654 (N_12654,N_12027,N_12267);
nand U12655 (N_12655,N_12116,N_12435);
or U12656 (N_12656,N_12141,N_12469);
nor U12657 (N_12657,N_12424,N_12379);
and U12658 (N_12658,N_12309,N_12102);
nor U12659 (N_12659,N_12081,N_12192);
xor U12660 (N_12660,N_12155,N_12075);
and U12661 (N_12661,N_12221,N_12476);
xor U12662 (N_12662,N_12172,N_12256);
xor U12663 (N_12663,N_12301,N_12229);
or U12664 (N_12664,N_12429,N_12269);
or U12665 (N_12665,N_12096,N_12449);
nor U12666 (N_12666,N_12030,N_12420);
nor U12667 (N_12667,N_12085,N_12432);
xnor U12668 (N_12668,N_12382,N_12174);
nor U12669 (N_12669,N_12209,N_12321);
or U12670 (N_12670,N_12254,N_12412);
or U12671 (N_12671,N_12076,N_12083);
or U12672 (N_12672,N_12453,N_12091);
nand U12673 (N_12673,N_12447,N_12317);
and U12674 (N_12674,N_12271,N_12346);
xnor U12675 (N_12675,N_12066,N_12097);
nand U12676 (N_12676,N_12045,N_12087);
or U12677 (N_12677,N_12265,N_12353);
and U12678 (N_12678,N_12054,N_12053);
nor U12679 (N_12679,N_12220,N_12455);
or U12680 (N_12680,N_12158,N_12138);
nor U12681 (N_12681,N_12474,N_12105);
nand U12682 (N_12682,N_12176,N_12226);
xnor U12683 (N_12683,N_12080,N_12377);
xnor U12684 (N_12684,N_12443,N_12136);
nor U12685 (N_12685,N_12119,N_12144);
or U12686 (N_12686,N_12365,N_12258);
xor U12687 (N_12687,N_12055,N_12107);
nand U12688 (N_12688,N_12276,N_12466);
nand U12689 (N_12689,N_12004,N_12421);
nand U12690 (N_12690,N_12067,N_12210);
nand U12691 (N_12691,N_12022,N_12341);
and U12692 (N_12692,N_12393,N_12015);
nand U12693 (N_12693,N_12188,N_12425);
nand U12694 (N_12694,N_12165,N_12115);
or U12695 (N_12695,N_12438,N_12255);
or U12696 (N_12696,N_12351,N_12003);
or U12697 (N_12697,N_12361,N_12295);
nor U12698 (N_12698,N_12417,N_12202);
nand U12699 (N_12699,N_12250,N_12064);
and U12700 (N_12700,N_12325,N_12225);
xnor U12701 (N_12701,N_12166,N_12423);
or U12702 (N_12702,N_12112,N_12342);
nor U12703 (N_12703,N_12127,N_12059);
nor U12704 (N_12704,N_12026,N_12031);
and U12705 (N_12705,N_12408,N_12242);
xor U12706 (N_12706,N_12088,N_12182);
nand U12707 (N_12707,N_12173,N_12319);
nand U12708 (N_12708,N_12305,N_12473);
nand U12709 (N_12709,N_12234,N_12303);
and U12710 (N_12710,N_12396,N_12128);
nor U12711 (N_12711,N_12219,N_12035);
and U12712 (N_12712,N_12117,N_12013);
xnor U12713 (N_12713,N_12190,N_12275);
xor U12714 (N_12714,N_12058,N_12486);
nor U12715 (N_12715,N_12465,N_12154);
xnor U12716 (N_12716,N_12458,N_12400);
nor U12717 (N_12717,N_12184,N_12422);
nor U12718 (N_12718,N_12398,N_12069);
and U12719 (N_12719,N_12103,N_12411);
nor U12720 (N_12720,N_12152,N_12060);
nand U12721 (N_12721,N_12480,N_12356);
nand U12722 (N_12722,N_12349,N_12042);
nand U12723 (N_12723,N_12106,N_12334);
nor U12724 (N_12724,N_12483,N_12179);
or U12725 (N_12725,N_12330,N_12248);
or U12726 (N_12726,N_12381,N_12038);
and U12727 (N_12727,N_12499,N_12407);
nand U12728 (N_12728,N_12278,N_12260);
nor U12729 (N_12729,N_12047,N_12460);
xnor U12730 (N_12730,N_12290,N_12428);
xnor U12731 (N_12731,N_12312,N_12259);
and U12732 (N_12732,N_12157,N_12195);
xor U12733 (N_12733,N_12289,N_12327);
and U12734 (N_12734,N_12314,N_12011);
xnor U12735 (N_12735,N_12156,N_12185);
xnor U12736 (N_12736,N_12137,N_12445);
or U12737 (N_12737,N_12479,N_12475);
and U12738 (N_12738,N_12164,N_12162);
xor U12739 (N_12739,N_12366,N_12292);
and U12740 (N_12740,N_12315,N_12300);
xor U12741 (N_12741,N_12431,N_12430);
and U12742 (N_12742,N_12326,N_12150);
nand U12743 (N_12743,N_12175,N_12126);
xor U12744 (N_12744,N_12272,N_12357);
xor U12745 (N_12745,N_12459,N_12245);
nand U12746 (N_12746,N_12370,N_12006);
and U12747 (N_12747,N_12178,N_12029);
xnor U12748 (N_12748,N_12347,N_12307);
xor U12749 (N_12749,N_12063,N_12313);
and U12750 (N_12750,N_12182,N_12478);
and U12751 (N_12751,N_12131,N_12339);
or U12752 (N_12752,N_12426,N_12187);
nor U12753 (N_12753,N_12434,N_12089);
nand U12754 (N_12754,N_12007,N_12291);
or U12755 (N_12755,N_12368,N_12455);
and U12756 (N_12756,N_12427,N_12440);
xor U12757 (N_12757,N_12270,N_12413);
nor U12758 (N_12758,N_12462,N_12335);
and U12759 (N_12759,N_12291,N_12390);
nor U12760 (N_12760,N_12226,N_12040);
nand U12761 (N_12761,N_12452,N_12336);
xor U12762 (N_12762,N_12079,N_12137);
xor U12763 (N_12763,N_12010,N_12429);
and U12764 (N_12764,N_12327,N_12145);
nor U12765 (N_12765,N_12193,N_12161);
nand U12766 (N_12766,N_12037,N_12331);
or U12767 (N_12767,N_12172,N_12451);
nor U12768 (N_12768,N_12161,N_12420);
and U12769 (N_12769,N_12410,N_12374);
nor U12770 (N_12770,N_12117,N_12011);
or U12771 (N_12771,N_12435,N_12337);
nor U12772 (N_12772,N_12419,N_12368);
and U12773 (N_12773,N_12299,N_12284);
and U12774 (N_12774,N_12208,N_12170);
xor U12775 (N_12775,N_12111,N_12266);
nand U12776 (N_12776,N_12314,N_12162);
and U12777 (N_12777,N_12187,N_12353);
nor U12778 (N_12778,N_12126,N_12162);
nand U12779 (N_12779,N_12111,N_12246);
xor U12780 (N_12780,N_12007,N_12060);
nand U12781 (N_12781,N_12322,N_12128);
and U12782 (N_12782,N_12385,N_12273);
nand U12783 (N_12783,N_12462,N_12061);
nand U12784 (N_12784,N_12182,N_12225);
xnor U12785 (N_12785,N_12382,N_12006);
nand U12786 (N_12786,N_12421,N_12329);
nor U12787 (N_12787,N_12046,N_12017);
or U12788 (N_12788,N_12244,N_12427);
nand U12789 (N_12789,N_12043,N_12486);
nand U12790 (N_12790,N_12296,N_12241);
and U12791 (N_12791,N_12012,N_12190);
nor U12792 (N_12792,N_12171,N_12421);
xnor U12793 (N_12793,N_12245,N_12226);
nand U12794 (N_12794,N_12022,N_12227);
nand U12795 (N_12795,N_12383,N_12441);
and U12796 (N_12796,N_12202,N_12095);
nor U12797 (N_12797,N_12487,N_12224);
nand U12798 (N_12798,N_12150,N_12118);
or U12799 (N_12799,N_12312,N_12137);
or U12800 (N_12800,N_12240,N_12378);
nor U12801 (N_12801,N_12413,N_12084);
nor U12802 (N_12802,N_12446,N_12491);
nand U12803 (N_12803,N_12133,N_12143);
and U12804 (N_12804,N_12166,N_12381);
nand U12805 (N_12805,N_12044,N_12016);
nand U12806 (N_12806,N_12126,N_12183);
xnor U12807 (N_12807,N_12398,N_12043);
xor U12808 (N_12808,N_12435,N_12027);
xor U12809 (N_12809,N_12383,N_12469);
and U12810 (N_12810,N_12250,N_12218);
xor U12811 (N_12811,N_12353,N_12158);
xnor U12812 (N_12812,N_12356,N_12141);
or U12813 (N_12813,N_12220,N_12255);
nor U12814 (N_12814,N_12086,N_12364);
nand U12815 (N_12815,N_12247,N_12122);
nor U12816 (N_12816,N_12111,N_12273);
xnor U12817 (N_12817,N_12019,N_12117);
or U12818 (N_12818,N_12181,N_12032);
nor U12819 (N_12819,N_12164,N_12427);
nand U12820 (N_12820,N_12365,N_12395);
nand U12821 (N_12821,N_12062,N_12203);
or U12822 (N_12822,N_12429,N_12057);
or U12823 (N_12823,N_12198,N_12060);
and U12824 (N_12824,N_12326,N_12010);
or U12825 (N_12825,N_12192,N_12098);
xnor U12826 (N_12826,N_12389,N_12059);
nand U12827 (N_12827,N_12478,N_12016);
or U12828 (N_12828,N_12071,N_12083);
xnor U12829 (N_12829,N_12121,N_12204);
xor U12830 (N_12830,N_12480,N_12050);
xor U12831 (N_12831,N_12288,N_12128);
and U12832 (N_12832,N_12033,N_12311);
and U12833 (N_12833,N_12004,N_12108);
xor U12834 (N_12834,N_12131,N_12017);
nand U12835 (N_12835,N_12352,N_12058);
nor U12836 (N_12836,N_12453,N_12429);
xor U12837 (N_12837,N_12232,N_12498);
and U12838 (N_12838,N_12176,N_12133);
and U12839 (N_12839,N_12423,N_12243);
or U12840 (N_12840,N_12235,N_12338);
or U12841 (N_12841,N_12003,N_12078);
xor U12842 (N_12842,N_12433,N_12180);
or U12843 (N_12843,N_12245,N_12438);
or U12844 (N_12844,N_12250,N_12242);
nor U12845 (N_12845,N_12432,N_12399);
or U12846 (N_12846,N_12459,N_12395);
or U12847 (N_12847,N_12148,N_12334);
or U12848 (N_12848,N_12400,N_12179);
nand U12849 (N_12849,N_12052,N_12293);
xnor U12850 (N_12850,N_12497,N_12155);
xnor U12851 (N_12851,N_12210,N_12103);
and U12852 (N_12852,N_12433,N_12330);
or U12853 (N_12853,N_12127,N_12440);
nor U12854 (N_12854,N_12454,N_12429);
xnor U12855 (N_12855,N_12036,N_12090);
or U12856 (N_12856,N_12334,N_12316);
and U12857 (N_12857,N_12211,N_12317);
nor U12858 (N_12858,N_12422,N_12233);
nor U12859 (N_12859,N_12083,N_12231);
and U12860 (N_12860,N_12335,N_12371);
or U12861 (N_12861,N_12283,N_12150);
nand U12862 (N_12862,N_12056,N_12008);
or U12863 (N_12863,N_12372,N_12412);
xor U12864 (N_12864,N_12424,N_12119);
nor U12865 (N_12865,N_12205,N_12267);
or U12866 (N_12866,N_12158,N_12377);
and U12867 (N_12867,N_12259,N_12435);
and U12868 (N_12868,N_12352,N_12156);
nor U12869 (N_12869,N_12270,N_12462);
and U12870 (N_12870,N_12223,N_12357);
and U12871 (N_12871,N_12031,N_12161);
xnor U12872 (N_12872,N_12346,N_12285);
xnor U12873 (N_12873,N_12224,N_12042);
xnor U12874 (N_12874,N_12196,N_12459);
nand U12875 (N_12875,N_12057,N_12463);
nor U12876 (N_12876,N_12457,N_12122);
or U12877 (N_12877,N_12007,N_12183);
or U12878 (N_12878,N_12444,N_12283);
and U12879 (N_12879,N_12357,N_12338);
nor U12880 (N_12880,N_12342,N_12087);
or U12881 (N_12881,N_12442,N_12103);
nor U12882 (N_12882,N_12148,N_12499);
and U12883 (N_12883,N_12193,N_12375);
xnor U12884 (N_12884,N_12152,N_12127);
nand U12885 (N_12885,N_12218,N_12204);
xor U12886 (N_12886,N_12423,N_12244);
or U12887 (N_12887,N_12103,N_12058);
xnor U12888 (N_12888,N_12376,N_12119);
and U12889 (N_12889,N_12335,N_12488);
xor U12890 (N_12890,N_12126,N_12268);
nor U12891 (N_12891,N_12302,N_12464);
nand U12892 (N_12892,N_12319,N_12063);
and U12893 (N_12893,N_12150,N_12085);
or U12894 (N_12894,N_12462,N_12138);
and U12895 (N_12895,N_12497,N_12440);
or U12896 (N_12896,N_12193,N_12267);
and U12897 (N_12897,N_12075,N_12201);
or U12898 (N_12898,N_12158,N_12154);
nor U12899 (N_12899,N_12135,N_12103);
xnor U12900 (N_12900,N_12077,N_12094);
or U12901 (N_12901,N_12101,N_12317);
or U12902 (N_12902,N_12320,N_12419);
xor U12903 (N_12903,N_12404,N_12115);
and U12904 (N_12904,N_12299,N_12148);
and U12905 (N_12905,N_12038,N_12403);
and U12906 (N_12906,N_12470,N_12288);
nand U12907 (N_12907,N_12224,N_12400);
nand U12908 (N_12908,N_12122,N_12194);
nor U12909 (N_12909,N_12420,N_12266);
or U12910 (N_12910,N_12076,N_12460);
nand U12911 (N_12911,N_12002,N_12488);
nor U12912 (N_12912,N_12242,N_12260);
or U12913 (N_12913,N_12347,N_12231);
xor U12914 (N_12914,N_12291,N_12260);
xor U12915 (N_12915,N_12432,N_12192);
nand U12916 (N_12916,N_12006,N_12059);
and U12917 (N_12917,N_12034,N_12038);
nor U12918 (N_12918,N_12214,N_12403);
nor U12919 (N_12919,N_12224,N_12312);
nor U12920 (N_12920,N_12024,N_12318);
xor U12921 (N_12921,N_12318,N_12499);
and U12922 (N_12922,N_12419,N_12003);
nor U12923 (N_12923,N_12134,N_12399);
or U12924 (N_12924,N_12059,N_12052);
nand U12925 (N_12925,N_12027,N_12110);
xor U12926 (N_12926,N_12327,N_12104);
or U12927 (N_12927,N_12406,N_12288);
xnor U12928 (N_12928,N_12151,N_12134);
or U12929 (N_12929,N_12462,N_12250);
and U12930 (N_12930,N_12253,N_12465);
nor U12931 (N_12931,N_12483,N_12225);
nor U12932 (N_12932,N_12069,N_12068);
nor U12933 (N_12933,N_12153,N_12193);
nand U12934 (N_12934,N_12363,N_12309);
nor U12935 (N_12935,N_12463,N_12425);
or U12936 (N_12936,N_12332,N_12050);
nor U12937 (N_12937,N_12112,N_12383);
nor U12938 (N_12938,N_12011,N_12185);
nand U12939 (N_12939,N_12056,N_12171);
xnor U12940 (N_12940,N_12165,N_12121);
or U12941 (N_12941,N_12188,N_12095);
or U12942 (N_12942,N_12396,N_12023);
and U12943 (N_12943,N_12180,N_12359);
xnor U12944 (N_12944,N_12286,N_12444);
or U12945 (N_12945,N_12244,N_12199);
nand U12946 (N_12946,N_12063,N_12139);
and U12947 (N_12947,N_12398,N_12430);
xor U12948 (N_12948,N_12380,N_12376);
xor U12949 (N_12949,N_12428,N_12296);
nand U12950 (N_12950,N_12320,N_12498);
xnor U12951 (N_12951,N_12044,N_12226);
and U12952 (N_12952,N_12064,N_12075);
xnor U12953 (N_12953,N_12259,N_12381);
or U12954 (N_12954,N_12384,N_12463);
or U12955 (N_12955,N_12312,N_12424);
xor U12956 (N_12956,N_12157,N_12122);
nor U12957 (N_12957,N_12195,N_12323);
or U12958 (N_12958,N_12345,N_12142);
xor U12959 (N_12959,N_12452,N_12255);
nor U12960 (N_12960,N_12251,N_12399);
xor U12961 (N_12961,N_12326,N_12093);
or U12962 (N_12962,N_12314,N_12333);
xor U12963 (N_12963,N_12356,N_12142);
nand U12964 (N_12964,N_12193,N_12379);
nor U12965 (N_12965,N_12382,N_12139);
nand U12966 (N_12966,N_12448,N_12049);
nand U12967 (N_12967,N_12277,N_12416);
and U12968 (N_12968,N_12146,N_12195);
xnor U12969 (N_12969,N_12098,N_12327);
xor U12970 (N_12970,N_12000,N_12271);
nor U12971 (N_12971,N_12276,N_12087);
or U12972 (N_12972,N_12257,N_12014);
nand U12973 (N_12973,N_12115,N_12324);
nor U12974 (N_12974,N_12443,N_12254);
nand U12975 (N_12975,N_12339,N_12027);
xor U12976 (N_12976,N_12001,N_12350);
xor U12977 (N_12977,N_12301,N_12385);
xor U12978 (N_12978,N_12230,N_12245);
nand U12979 (N_12979,N_12326,N_12166);
nand U12980 (N_12980,N_12218,N_12036);
xnor U12981 (N_12981,N_12007,N_12133);
and U12982 (N_12982,N_12134,N_12373);
nand U12983 (N_12983,N_12043,N_12374);
and U12984 (N_12984,N_12196,N_12052);
nor U12985 (N_12985,N_12287,N_12022);
xor U12986 (N_12986,N_12164,N_12389);
or U12987 (N_12987,N_12465,N_12092);
or U12988 (N_12988,N_12131,N_12204);
nand U12989 (N_12989,N_12046,N_12419);
and U12990 (N_12990,N_12200,N_12324);
xor U12991 (N_12991,N_12217,N_12079);
nand U12992 (N_12992,N_12493,N_12266);
nor U12993 (N_12993,N_12129,N_12117);
or U12994 (N_12994,N_12130,N_12493);
nand U12995 (N_12995,N_12173,N_12063);
and U12996 (N_12996,N_12173,N_12212);
and U12997 (N_12997,N_12430,N_12428);
nand U12998 (N_12998,N_12487,N_12456);
nand U12999 (N_12999,N_12105,N_12131);
or U13000 (N_13000,N_12675,N_12936);
nor U13001 (N_13001,N_12543,N_12997);
xnor U13002 (N_13002,N_12663,N_12837);
nand U13003 (N_13003,N_12773,N_12798);
xnor U13004 (N_13004,N_12963,N_12615);
and U13005 (N_13005,N_12737,N_12525);
nand U13006 (N_13006,N_12602,N_12645);
nor U13007 (N_13007,N_12589,N_12971);
xnor U13008 (N_13008,N_12641,N_12574);
and U13009 (N_13009,N_12923,N_12839);
xnor U13010 (N_13010,N_12551,N_12616);
xnor U13011 (N_13011,N_12863,N_12503);
and U13012 (N_13012,N_12911,N_12517);
nor U13013 (N_13013,N_12665,N_12850);
or U13014 (N_13014,N_12873,N_12741);
nand U13015 (N_13015,N_12921,N_12766);
nand U13016 (N_13016,N_12761,N_12989);
and U13017 (N_13017,N_12701,N_12662);
and U13018 (N_13018,N_12804,N_12985);
xnor U13019 (N_13019,N_12747,N_12678);
xor U13020 (N_13020,N_12995,N_12550);
or U13021 (N_13021,N_12728,N_12890);
nand U13022 (N_13022,N_12639,N_12722);
xnor U13023 (N_13023,N_12729,N_12857);
xor U13024 (N_13024,N_12870,N_12607);
nor U13025 (N_13025,N_12751,N_12868);
xnor U13026 (N_13026,N_12869,N_12695);
or U13027 (N_13027,N_12820,N_12768);
xnor U13028 (N_13028,N_12875,N_12745);
or U13029 (N_13029,N_12955,N_12774);
xor U13030 (N_13030,N_12805,N_12946);
nor U13031 (N_13031,N_12933,N_12530);
xnor U13032 (N_13032,N_12723,N_12548);
or U13033 (N_13033,N_12860,N_12852);
or U13034 (N_13034,N_12735,N_12856);
or U13035 (N_13035,N_12784,N_12508);
and U13036 (N_13036,N_12902,N_12754);
or U13037 (N_13037,N_12789,N_12585);
xor U13038 (N_13038,N_12840,N_12811);
nor U13039 (N_13039,N_12898,N_12590);
nand U13040 (N_13040,N_12785,N_12769);
nor U13041 (N_13041,N_12521,N_12601);
or U13042 (N_13042,N_12622,N_12793);
and U13043 (N_13043,N_12709,N_12760);
xor U13044 (N_13044,N_12649,N_12644);
xnor U13045 (N_13045,N_12549,N_12648);
xnor U13046 (N_13046,N_12986,N_12726);
nor U13047 (N_13047,N_12818,N_12948);
nand U13048 (N_13048,N_12515,N_12573);
or U13049 (N_13049,N_12755,N_12881);
and U13050 (N_13050,N_12600,N_12762);
xor U13051 (N_13051,N_12894,N_12721);
or U13052 (N_13052,N_12579,N_12987);
or U13053 (N_13053,N_12611,N_12799);
nand U13054 (N_13054,N_12795,N_12929);
or U13055 (N_13055,N_12567,N_12674);
and U13056 (N_13056,N_12779,N_12738);
or U13057 (N_13057,N_12560,N_12966);
nand U13058 (N_13058,N_12536,N_12512);
nand U13059 (N_13059,N_12927,N_12564);
or U13060 (N_13060,N_12937,N_12866);
nand U13061 (N_13061,N_12896,N_12900);
and U13062 (N_13062,N_12862,N_12878);
nor U13063 (N_13063,N_12834,N_12913);
and U13064 (N_13064,N_12719,N_12990);
or U13065 (N_13065,N_12786,N_12707);
nand U13066 (N_13066,N_12667,N_12706);
xnor U13067 (N_13067,N_12874,N_12630);
xnor U13068 (N_13068,N_12893,N_12565);
xnor U13069 (N_13069,N_12808,N_12651);
or U13070 (N_13070,N_12626,N_12570);
xor U13071 (N_13071,N_12578,N_12715);
or U13072 (N_13072,N_12671,N_12800);
nor U13073 (N_13073,N_12920,N_12625);
and U13074 (N_13074,N_12531,N_12988);
or U13075 (N_13075,N_12539,N_12711);
or U13076 (N_13076,N_12770,N_12763);
nor U13077 (N_13077,N_12838,N_12960);
or U13078 (N_13078,N_12664,N_12841);
xnor U13079 (N_13079,N_12702,N_12813);
or U13080 (N_13080,N_12858,N_12951);
nand U13081 (N_13081,N_12764,N_12712);
or U13082 (N_13082,N_12572,N_12757);
and U13083 (N_13083,N_12608,N_12912);
or U13084 (N_13084,N_12859,N_12683);
and U13085 (N_13085,N_12851,N_12931);
and U13086 (N_13086,N_12733,N_12756);
and U13087 (N_13087,N_12928,N_12734);
xnor U13088 (N_13088,N_12666,N_12825);
nor U13089 (N_13089,N_12584,N_12610);
xor U13090 (N_13090,N_12516,N_12624);
and U13091 (N_13091,N_12593,N_12716);
and U13092 (N_13092,N_12545,N_12821);
nor U13093 (N_13093,N_12872,N_12970);
xor U13094 (N_13094,N_12725,N_12887);
nand U13095 (N_13095,N_12563,N_12807);
and U13096 (N_13096,N_12926,N_12705);
or U13097 (N_13097,N_12953,N_12700);
nor U13098 (N_13098,N_12500,N_12999);
and U13099 (N_13099,N_12698,N_12778);
xnor U13100 (N_13100,N_12771,N_12681);
and U13101 (N_13101,N_12680,N_12682);
xor U13102 (N_13102,N_12861,N_12659);
xnor U13103 (N_13103,N_12520,N_12653);
or U13104 (N_13104,N_12930,N_12606);
nor U13105 (N_13105,N_12583,N_12886);
nor U13106 (N_13106,N_12686,N_12958);
nor U13107 (N_13107,N_12802,N_12777);
or U13108 (N_13108,N_12961,N_12855);
nor U13109 (N_13109,N_12504,N_12910);
or U13110 (N_13110,N_12993,N_12612);
xor U13111 (N_13111,N_12720,N_12914);
xor U13112 (N_13112,N_12591,N_12758);
and U13113 (N_13113,N_12724,N_12978);
nor U13114 (N_13114,N_12984,N_12628);
nor U13115 (N_13115,N_12824,N_12580);
and U13116 (N_13116,N_12939,N_12919);
nand U13117 (N_13117,N_12979,N_12907);
or U13118 (N_13118,N_12934,N_12740);
nor U13119 (N_13119,N_12957,N_12638);
or U13120 (N_13120,N_12688,N_12782);
and U13121 (N_13121,N_12609,N_12621);
nand U13122 (N_13122,N_12915,N_12592);
and U13123 (N_13123,N_12830,N_12952);
xor U13124 (N_13124,N_12932,N_12627);
nand U13125 (N_13125,N_12561,N_12901);
and U13126 (N_13126,N_12876,N_12569);
and U13127 (N_13127,N_12614,N_12581);
nand U13128 (N_13128,N_12540,N_12604);
nand U13129 (N_13129,N_12636,N_12947);
nor U13130 (N_13130,N_12699,N_12884);
and U13131 (N_13131,N_12708,N_12642);
nand U13132 (N_13132,N_12596,N_12534);
nor U13133 (N_13133,N_12750,N_12677);
nand U13134 (N_13134,N_12513,N_12511);
and U13135 (N_13135,N_12576,N_12619);
nor U13136 (N_13136,N_12657,N_12658);
nor U13137 (N_13137,N_12836,N_12996);
nor U13138 (N_13138,N_12618,N_12742);
and U13139 (N_13139,N_12817,N_12991);
nand U13140 (N_13140,N_12787,N_12822);
nand U13141 (N_13141,N_12949,N_12599);
or U13142 (N_13142,N_12848,N_12917);
nand U13143 (N_13143,N_12660,N_12823);
nor U13144 (N_13144,N_12588,N_12739);
or U13145 (N_13145,N_12577,N_12717);
nand U13146 (N_13146,N_12690,N_12629);
or U13147 (N_13147,N_12803,N_12692);
xor U13148 (N_13148,N_12633,N_12810);
nand U13149 (N_13149,N_12522,N_12746);
nor U13150 (N_13150,N_12586,N_12555);
or U13151 (N_13151,N_12670,N_12637);
nor U13152 (N_13152,N_12714,N_12865);
xnor U13153 (N_13153,N_12544,N_12964);
nand U13154 (N_13154,N_12956,N_12704);
nand U13155 (N_13155,N_12781,N_12634);
nand U13156 (N_13156,N_12689,N_12788);
nor U13157 (N_13157,N_12526,N_12767);
nor U13158 (N_13158,N_12832,N_12983);
and U13159 (N_13159,N_12973,N_12967);
xnor U13160 (N_13160,N_12968,N_12542);
or U13161 (N_13161,N_12879,N_12847);
nand U13162 (N_13162,N_12685,N_12655);
and U13163 (N_13163,N_12669,N_12944);
or U13164 (N_13164,N_12814,N_12546);
nand U13165 (N_13165,N_12980,N_12713);
or U13166 (N_13166,N_12864,N_12994);
xnor U13167 (N_13167,N_12889,N_12552);
nor U13168 (N_13168,N_12965,N_12587);
or U13169 (N_13169,N_12909,N_12916);
nand U13170 (N_13170,N_12918,N_12620);
and U13171 (N_13171,N_12595,N_12790);
nor U13172 (N_13172,N_12730,N_12752);
or U13173 (N_13173,N_12892,N_12753);
and U13174 (N_13174,N_12718,N_12582);
and U13175 (N_13175,N_12679,N_12528);
nand U13176 (N_13176,N_12553,N_12696);
nor U13177 (N_13177,N_12833,N_12831);
or U13178 (N_13178,N_12535,N_12977);
nor U13179 (N_13179,N_12661,N_12849);
nand U13180 (N_13180,N_12732,N_12940);
nand U13181 (N_13181,N_12815,N_12806);
nor U13182 (N_13182,N_12812,N_12883);
nand U13183 (N_13183,N_12668,N_12791);
and U13184 (N_13184,N_12826,N_12974);
and U13185 (N_13185,N_12853,N_12623);
or U13186 (N_13186,N_12976,N_12827);
and U13187 (N_13187,N_12556,N_12731);
nand U13188 (N_13188,N_12532,N_12801);
or U13189 (N_13189,N_12575,N_12809);
nand U13190 (N_13190,N_12505,N_12597);
nor U13191 (N_13191,N_12643,N_12506);
and U13192 (N_13192,N_12906,N_12935);
nor U13193 (N_13193,N_12529,N_12524);
xor U13194 (N_13194,N_12835,N_12509);
and U13195 (N_13195,N_12537,N_12945);
or U13196 (N_13196,N_12558,N_12672);
or U13197 (N_13197,N_12559,N_12962);
or U13198 (N_13198,N_12571,N_12744);
xor U13199 (N_13199,N_12891,N_12897);
and U13200 (N_13200,N_12693,N_12650);
and U13201 (N_13201,N_12829,N_12647);
or U13202 (N_13202,N_12603,N_12568);
nor U13203 (N_13203,N_12938,N_12792);
nor U13204 (N_13204,N_12523,N_12941);
nand U13205 (N_13205,N_12950,N_12518);
xor U13206 (N_13206,N_12888,N_12924);
nand U13207 (N_13207,N_12903,N_12710);
or U13208 (N_13208,N_12594,N_12640);
nand U13209 (N_13209,N_12783,N_12765);
or U13210 (N_13210,N_12527,N_12703);
nand U13211 (N_13211,N_12736,N_12877);
nor U13212 (N_13212,N_12656,N_12882);
xor U13213 (N_13213,N_12519,N_12538);
nand U13214 (N_13214,N_12794,N_12727);
and U13215 (N_13215,N_12796,N_12981);
and U13216 (N_13216,N_12652,N_12842);
nor U13217 (N_13217,N_12880,N_12871);
nand U13218 (N_13218,N_12844,N_12748);
nand U13219 (N_13219,N_12691,N_12514);
nor U13220 (N_13220,N_12843,N_12885);
nor U13221 (N_13221,N_12502,N_12566);
nor U13222 (N_13222,N_12959,N_12972);
xnor U13223 (N_13223,N_12943,N_12776);
and U13224 (N_13224,N_12925,N_12816);
xor U13225 (N_13225,N_12613,N_12510);
nand U13226 (N_13226,N_12895,N_12687);
nand U13227 (N_13227,N_12905,N_12541);
and U13228 (N_13228,N_12557,N_12547);
and U13229 (N_13229,N_12759,N_12904);
or U13230 (N_13230,N_12975,N_12632);
nor U13231 (N_13231,N_12673,N_12954);
nand U13232 (N_13232,N_12605,N_12780);
xnor U13233 (N_13233,N_12867,N_12697);
and U13234 (N_13234,N_12922,N_12797);
and U13235 (N_13235,N_12684,N_12743);
and U13236 (N_13236,N_12775,N_12772);
and U13237 (N_13237,N_12846,N_12562);
and U13238 (N_13238,N_12749,N_12694);
nor U13239 (N_13239,N_12635,N_12992);
nor U13240 (N_13240,N_12654,N_12554);
nor U13241 (N_13241,N_12646,N_12828);
nor U13242 (N_13242,N_12845,N_12617);
nand U13243 (N_13243,N_12676,N_12998);
nand U13244 (N_13244,N_12908,N_12819);
or U13245 (N_13245,N_12598,N_12899);
nor U13246 (N_13246,N_12631,N_12969);
or U13247 (N_13247,N_12854,N_12982);
nor U13248 (N_13248,N_12533,N_12501);
nand U13249 (N_13249,N_12942,N_12507);
or U13250 (N_13250,N_12986,N_12553);
nor U13251 (N_13251,N_12875,N_12692);
or U13252 (N_13252,N_12893,N_12799);
nand U13253 (N_13253,N_12829,N_12933);
or U13254 (N_13254,N_12726,N_12638);
nand U13255 (N_13255,N_12737,N_12894);
nor U13256 (N_13256,N_12750,N_12622);
and U13257 (N_13257,N_12591,N_12808);
and U13258 (N_13258,N_12640,N_12617);
nor U13259 (N_13259,N_12899,N_12619);
nand U13260 (N_13260,N_12934,N_12708);
nand U13261 (N_13261,N_12526,N_12965);
nand U13262 (N_13262,N_12804,N_12753);
nand U13263 (N_13263,N_12758,N_12893);
and U13264 (N_13264,N_12750,N_12686);
and U13265 (N_13265,N_12709,N_12971);
and U13266 (N_13266,N_12646,N_12570);
xor U13267 (N_13267,N_12677,N_12568);
nor U13268 (N_13268,N_12594,N_12638);
nand U13269 (N_13269,N_12591,N_12859);
and U13270 (N_13270,N_12911,N_12928);
xor U13271 (N_13271,N_12668,N_12561);
and U13272 (N_13272,N_12978,N_12520);
nor U13273 (N_13273,N_12592,N_12902);
xor U13274 (N_13274,N_12875,N_12907);
nand U13275 (N_13275,N_12681,N_12951);
nor U13276 (N_13276,N_12577,N_12941);
nor U13277 (N_13277,N_12797,N_12694);
or U13278 (N_13278,N_12788,N_12789);
or U13279 (N_13279,N_12746,N_12873);
xnor U13280 (N_13280,N_12763,N_12739);
nand U13281 (N_13281,N_12728,N_12962);
xor U13282 (N_13282,N_12859,N_12793);
or U13283 (N_13283,N_12821,N_12764);
xnor U13284 (N_13284,N_12857,N_12847);
or U13285 (N_13285,N_12746,N_12974);
nand U13286 (N_13286,N_12805,N_12938);
nor U13287 (N_13287,N_12902,N_12833);
xor U13288 (N_13288,N_12736,N_12830);
or U13289 (N_13289,N_12757,N_12839);
xnor U13290 (N_13290,N_12776,N_12593);
and U13291 (N_13291,N_12563,N_12718);
xnor U13292 (N_13292,N_12857,N_12569);
or U13293 (N_13293,N_12788,N_12893);
xnor U13294 (N_13294,N_12701,N_12571);
or U13295 (N_13295,N_12957,N_12725);
nor U13296 (N_13296,N_12669,N_12870);
or U13297 (N_13297,N_12621,N_12614);
and U13298 (N_13298,N_12833,N_12599);
or U13299 (N_13299,N_12944,N_12979);
or U13300 (N_13300,N_12800,N_12536);
and U13301 (N_13301,N_12829,N_12964);
and U13302 (N_13302,N_12638,N_12822);
nand U13303 (N_13303,N_12577,N_12653);
xor U13304 (N_13304,N_12784,N_12956);
and U13305 (N_13305,N_12508,N_12562);
nor U13306 (N_13306,N_12987,N_12921);
nand U13307 (N_13307,N_12936,N_12912);
nor U13308 (N_13308,N_12516,N_12984);
and U13309 (N_13309,N_12990,N_12702);
nand U13310 (N_13310,N_12636,N_12908);
nor U13311 (N_13311,N_12949,N_12593);
nand U13312 (N_13312,N_12568,N_12896);
xnor U13313 (N_13313,N_12860,N_12644);
nand U13314 (N_13314,N_12627,N_12940);
or U13315 (N_13315,N_12968,N_12697);
xnor U13316 (N_13316,N_12988,N_12907);
xor U13317 (N_13317,N_12501,N_12837);
xor U13318 (N_13318,N_12966,N_12736);
nand U13319 (N_13319,N_12823,N_12593);
nand U13320 (N_13320,N_12960,N_12528);
or U13321 (N_13321,N_12539,N_12706);
nor U13322 (N_13322,N_12613,N_12939);
xnor U13323 (N_13323,N_12544,N_12972);
or U13324 (N_13324,N_12770,N_12573);
xor U13325 (N_13325,N_12698,N_12989);
or U13326 (N_13326,N_12637,N_12829);
nand U13327 (N_13327,N_12584,N_12781);
and U13328 (N_13328,N_12961,N_12542);
nand U13329 (N_13329,N_12994,N_12900);
and U13330 (N_13330,N_12763,N_12674);
xor U13331 (N_13331,N_12947,N_12694);
and U13332 (N_13332,N_12884,N_12551);
and U13333 (N_13333,N_12780,N_12756);
xnor U13334 (N_13334,N_12935,N_12611);
or U13335 (N_13335,N_12853,N_12846);
or U13336 (N_13336,N_12518,N_12906);
nor U13337 (N_13337,N_12748,N_12775);
and U13338 (N_13338,N_12789,N_12548);
or U13339 (N_13339,N_12784,N_12592);
or U13340 (N_13340,N_12734,N_12673);
nor U13341 (N_13341,N_12952,N_12743);
or U13342 (N_13342,N_12844,N_12533);
nand U13343 (N_13343,N_12579,N_12978);
xor U13344 (N_13344,N_12836,N_12603);
nand U13345 (N_13345,N_12516,N_12956);
and U13346 (N_13346,N_12923,N_12883);
or U13347 (N_13347,N_12532,N_12507);
or U13348 (N_13348,N_12515,N_12611);
xor U13349 (N_13349,N_12792,N_12642);
nor U13350 (N_13350,N_12502,N_12942);
nor U13351 (N_13351,N_12750,N_12649);
nand U13352 (N_13352,N_12987,N_12850);
xor U13353 (N_13353,N_12761,N_12672);
nand U13354 (N_13354,N_12795,N_12675);
nand U13355 (N_13355,N_12655,N_12972);
nor U13356 (N_13356,N_12783,N_12503);
xor U13357 (N_13357,N_12884,N_12623);
nand U13358 (N_13358,N_12558,N_12619);
nor U13359 (N_13359,N_12708,N_12649);
nor U13360 (N_13360,N_12778,N_12624);
or U13361 (N_13361,N_12558,N_12865);
xor U13362 (N_13362,N_12805,N_12825);
or U13363 (N_13363,N_12670,N_12755);
or U13364 (N_13364,N_12814,N_12951);
nand U13365 (N_13365,N_12790,N_12585);
xnor U13366 (N_13366,N_12747,N_12593);
nand U13367 (N_13367,N_12672,N_12566);
xor U13368 (N_13368,N_12535,N_12516);
xor U13369 (N_13369,N_12941,N_12701);
or U13370 (N_13370,N_12872,N_12709);
nor U13371 (N_13371,N_12524,N_12525);
or U13372 (N_13372,N_12829,N_12773);
and U13373 (N_13373,N_12909,N_12657);
nand U13374 (N_13374,N_12982,N_12797);
nor U13375 (N_13375,N_12823,N_12942);
nand U13376 (N_13376,N_12869,N_12792);
nand U13377 (N_13377,N_12550,N_12912);
nor U13378 (N_13378,N_12573,N_12759);
or U13379 (N_13379,N_12525,N_12691);
nor U13380 (N_13380,N_12613,N_12807);
nor U13381 (N_13381,N_12820,N_12539);
nor U13382 (N_13382,N_12694,N_12669);
nand U13383 (N_13383,N_12911,N_12612);
xnor U13384 (N_13384,N_12604,N_12690);
or U13385 (N_13385,N_12900,N_12612);
and U13386 (N_13386,N_12825,N_12500);
xnor U13387 (N_13387,N_12760,N_12547);
xor U13388 (N_13388,N_12913,N_12950);
and U13389 (N_13389,N_12560,N_12848);
and U13390 (N_13390,N_12554,N_12780);
or U13391 (N_13391,N_12816,N_12856);
xnor U13392 (N_13392,N_12747,N_12887);
or U13393 (N_13393,N_12967,N_12553);
or U13394 (N_13394,N_12960,N_12583);
nor U13395 (N_13395,N_12560,N_12802);
nand U13396 (N_13396,N_12772,N_12564);
nor U13397 (N_13397,N_12778,N_12898);
and U13398 (N_13398,N_12789,N_12664);
or U13399 (N_13399,N_12710,N_12836);
and U13400 (N_13400,N_12643,N_12859);
xor U13401 (N_13401,N_12892,N_12675);
xor U13402 (N_13402,N_12827,N_12658);
nand U13403 (N_13403,N_12832,N_12951);
nor U13404 (N_13404,N_12592,N_12557);
xnor U13405 (N_13405,N_12819,N_12890);
nor U13406 (N_13406,N_12575,N_12614);
and U13407 (N_13407,N_12762,N_12936);
nor U13408 (N_13408,N_12829,N_12564);
and U13409 (N_13409,N_12746,N_12764);
and U13410 (N_13410,N_12552,N_12668);
xnor U13411 (N_13411,N_12662,N_12966);
or U13412 (N_13412,N_12754,N_12623);
nand U13413 (N_13413,N_12576,N_12910);
nor U13414 (N_13414,N_12980,N_12939);
and U13415 (N_13415,N_12878,N_12798);
nor U13416 (N_13416,N_12517,N_12566);
xnor U13417 (N_13417,N_12585,N_12963);
nor U13418 (N_13418,N_12901,N_12912);
nand U13419 (N_13419,N_12727,N_12948);
xnor U13420 (N_13420,N_12623,N_12947);
nand U13421 (N_13421,N_12646,N_12500);
and U13422 (N_13422,N_12844,N_12723);
nand U13423 (N_13423,N_12626,N_12855);
and U13424 (N_13424,N_12563,N_12540);
nand U13425 (N_13425,N_12887,N_12729);
and U13426 (N_13426,N_12842,N_12804);
or U13427 (N_13427,N_12526,N_12766);
xor U13428 (N_13428,N_12616,N_12739);
or U13429 (N_13429,N_12932,N_12863);
nor U13430 (N_13430,N_12790,N_12649);
and U13431 (N_13431,N_12778,N_12925);
or U13432 (N_13432,N_12569,N_12849);
nor U13433 (N_13433,N_12542,N_12601);
xnor U13434 (N_13434,N_12509,N_12994);
nand U13435 (N_13435,N_12691,N_12581);
nor U13436 (N_13436,N_12638,N_12646);
and U13437 (N_13437,N_12685,N_12812);
and U13438 (N_13438,N_12847,N_12621);
and U13439 (N_13439,N_12875,N_12525);
nor U13440 (N_13440,N_12629,N_12644);
nor U13441 (N_13441,N_12597,N_12733);
nand U13442 (N_13442,N_12963,N_12921);
nor U13443 (N_13443,N_12911,N_12539);
and U13444 (N_13444,N_12982,N_12671);
and U13445 (N_13445,N_12760,N_12990);
and U13446 (N_13446,N_12783,N_12610);
and U13447 (N_13447,N_12752,N_12854);
nor U13448 (N_13448,N_12964,N_12958);
and U13449 (N_13449,N_12815,N_12745);
nand U13450 (N_13450,N_12609,N_12969);
nand U13451 (N_13451,N_12699,N_12713);
or U13452 (N_13452,N_12991,N_12851);
and U13453 (N_13453,N_12957,N_12947);
or U13454 (N_13454,N_12512,N_12933);
xnor U13455 (N_13455,N_12581,N_12918);
and U13456 (N_13456,N_12684,N_12923);
or U13457 (N_13457,N_12640,N_12932);
nand U13458 (N_13458,N_12896,N_12978);
nor U13459 (N_13459,N_12814,N_12788);
nor U13460 (N_13460,N_12511,N_12755);
nand U13461 (N_13461,N_12997,N_12643);
or U13462 (N_13462,N_12555,N_12934);
and U13463 (N_13463,N_12742,N_12989);
nand U13464 (N_13464,N_12887,N_12898);
or U13465 (N_13465,N_12796,N_12917);
or U13466 (N_13466,N_12832,N_12797);
nor U13467 (N_13467,N_12560,N_12756);
or U13468 (N_13468,N_12993,N_12717);
nand U13469 (N_13469,N_12604,N_12511);
nor U13470 (N_13470,N_12585,N_12869);
and U13471 (N_13471,N_12791,N_12954);
xor U13472 (N_13472,N_12978,N_12832);
xnor U13473 (N_13473,N_12613,N_12838);
and U13474 (N_13474,N_12750,N_12578);
xor U13475 (N_13475,N_12589,N_12651);
and U13476 (N_13476,N_12501,N_12891);
xor U13477 (N_13477,N_12795,N_12608);
or U13478 (N_13478,N_12584,N_12643);
nor U13479 (N_13479,N_12654,N_12942);
nor U13480 (N_13480,N_12954,N_12989);
nor U13481 (N_13481,N_12515,N_12843);
nor U13482 (N_13482,N_12765,N_12535);
nor U13483 (N_13483,N_12728,N_12977);
nor U13484 (N_13484,N_12905,N_12816);
nand U13485 (N_13485,N_12567,N_12751);
nor U13486 (N_13486,N_12822,N_12916);
xor U13487 (N_13487,N_12587,N_12653);
or U13488 (N_13488,N_12892,N_12652);
and U13489 (N_13489,N_12787,N_12621);
and U13490 (N_13490,N_12913,N_12624);
and U13491 (N_13491,N_12946,N_12998);
and U13492 (N_13492,N_12948,N_12638);
and U13493 (N_13493,N_12853,N_12614);
nor U13494 (N_13494,N_12617,N_12886);
xnor U13495 (N_13495,N_12867,N_12760);
or U13496 (N_13496,N_12889,N_12815);
nand U13497 (N_13497,N_12736,N_12783);
nand U13498 (N_13498,N_12682,N_12938);
nor U13499 (N_13499,N_12601,N_12951);
or U13500 (N_13500,N_13401,N_13473);
xor U13501 (N_13501,N_13020,N_13194);
nand U13502 (N_13502,N_13129,N_13202);
or U13503 (N_13503,N_13170,N_13210);
nor U13504 (N_13504,N_13387,N_13152);
xnor U13505 (N_13505,N_13464,N_13304);
nand U13506 (N_13506,N_13485,N_13320);
xnor U13507 (N_13507,N_13157,N_13144);
and U13508 (N_13508,N_13119,N_13084);
and U13509 (N_13509,N_13469,N_13021);
and U13510 (N_13510,N_13291,N_13322);
xnor U13511 (N_13511,N_13372,N_13145);
nor U13512 (N_13512,N_13420,N_13406);
or U13513 (N_13513,N_13236,N_13013);
nand U13514 (N_13514,N_13216,N_13318);
or U13515 (N_13515,N_13112,N_13288);
nand U13516 (N_13516,N_13051,N_13414);
nor U13517 (N_13517,N_13223,N_13100);
nand U13518 (N_13518,N_13371,N_13150);
nand U13519 (N_13519,N_13040,N_13085);
xor U13520 (N_13520,N_13249,N_13224);
xor U13521 (N_13521,N_13275,N_13008);
xor U13522 (N_13522,N_13125,N_13063);
nand U13523 (N_13523,N_13234,N_13491);
nor U13524 (N_13524,N_13128,N_13316);
nand U13525 (N_13525,N_13427,N_13199);
nor U13526 (N_13526,N_13358,N_13294);
xor U13527 (N_13527,N_13321,N_13001);
and U13528 (N_13528,N_13036,N_13292);
xor U13529 (N_13529,N_13211,N_13400);
xor U13530 (N_13530,N_13277,N_13446);
xor U13531 (N_13531,N_13107,N_13424);
nor U13532 (N_13532,N_13383,N_13127);
nor U13533 (N_13533,N_13237,N_13088);
and U13534 (N_13534,N_13094,N_13432);
xnor U13535 (N_13535,N_13189,N_13232);
and U13536 (N_13536,N_13488,N_13238);
or U13537 (N_13537,N_13208,N_13384);
nand U13538 (N_13538,N_13311,N_13258);
xnor U13539 (N_13539,N_13395,N_13018);
xnor U13540 (N_13540,N_13142,N_13172);
nor U13541 (N_13541,N_13156,N_13255);
xor U13542 (N_13542,N_13069,N_13350);
nand U13543 (N_13543,N_13265,N_13066);
and U13544 (N_13544,N_13283,N_13264);
nor U13545 (N_13545,N_13435,N_13287);
or U13546 (N_13546,N_13442,N_13022);
xnor U13547 (N_13547,N_13204,N_13039);
and U13548 (N_13548,N_13086,N_13334);
or U13549 (N_13549,N_13399,N_13391);
xor U13550 (N_13550,N_13183,N_13028);
nand U13551 (N_13551,N_13072,N_13034);
and U13552 (N_13552,N_13148,N_13062);
or U13553 (N_13553,N_13184,N_13165);
or U13554 (N_13554,N_13413,N_13181);
and U13555 (N_13555,N_13076,N_13425);
and U13556 (N_13556,N_13380,N_13226);
or U13557 (N_13557,N_13359,N_13059);
or U13558 (N_13558,N_13079,N_13466);
and U13559 (N_13559,N_13201,N_13138);
and U13560 (N_13560,N_13071,N_13168);
xnor U13561 (N_13561,N_13389,N_13332);
xor U13562 (N_13562,N_13467,N_13324);
nor U13563 (N_13563,N_13319,N_13045);
and U13564 (N_13564,N_13049,N_13106);
and U13565 (N_13565,N_13483,N_13019);
nor U13566 (N_13566,N_13038,N_13227);
nand U13567 (N_13567,N_13115,N_13489);
xnor U13568 (N_13568,N_13303,N_13460);
or U13569 (N_13569,N_13269,N_13012);
nand U13570 (N_13570,N_13338,N_13381);
or U13571 (N_13571,N_13271,N_13472);
xor U13572 (N_13572,N_13171,N_13477);
or U13573 (N_13573,N_13445,N_13360);
nand U13574 (N_13574,N_13180,N_13123);
xnor U13575 (N_13575,N_13465,N_13447);
and U13576 (N_13576,N_13176,N_13299);
and U13577 (N_13577,N_13197,N_13124);
nor U13578 (N_13578,N_13159,N_13101);
and U13579 (N_13579,N_13089,N_13367);
and U13580 (N_13580,N_13033,N_13354);
nand U13581 (N_13581,N_13268,N_13104);
or U13582 (N_13582,N_13476,N_13459);
nor U13583 (N_13583,N_13035,N_13468);
xnor U13584 (N_13584,N_13209,N_13300);
nor U13585 (N_13585,N_13370,N_13245);
nor U13586 (N_13586,N_13130,N_13247);
xor U13587 (N_13587,N_13498,N_13212);
xor U13588 (N_13588,N_13011,N_13302);
or U13589 (N_13589,N_13002,N_13060);
xor U13590 (N_13590,N_13274,N_13487);
or U13591 (N_13591,N_13133,N_13331);
nor U13592 (N_13592,N_13496,N_13290);
xor U13593 (N_13593,N_13207,N_13481);
nand U13594 (N_13594,N_13080,N_13217);
nor U13595 (N_13595,N_13047,N_13041);
or U13596 (N_13596,N_13032,N_13270);
xor U13597 (N_13597,N_13286,N_13024);
xor U13598 (N_13598,N_13281,N_13110);
nand U13599 (N_13599,N_13365,N_13014);
nand U13600 (N_13600,N_13355,N_13139);
or U13601 (N_13601,N_13273,N_13474);
nand U13602 (N_13602,N_13308,N_13193);
xor U13603 (N_13603,N_13221,N_13007);
or U13604 (N_13604,N_13105,N_13437);
or U13605 (N_13605,N_13376,N_13462);
xnor U13606 (N_13606,N_13453,N_13261);
and U13607 (N_13607,N_13449,N_13305);
and U13608 (N_13608,N_13337,N_13187);
and U13609 (N_13609,N_13393,N_13064);
nor U13610 (N_13610,N_13048,N_13402);
or U13611 (N_13611,N_13450,N_13225);
nor U13612 (N_13612,N_13251,N_13284);
nand U13613 (N_13613,N_13412,N_13254);
and U13614 (N_13614,N_13031,N_13361);
nor U13615 (N_13615,N_13407,N_13117);
and U13616 (N_13616,N_13233,N_13428);
or U13617 (N_13617,N_13423,N_13073);
nand U13618 (N_13618,N_13030,N_13392);
and U13619 (N_13619,N_13443,N_13158);
or U13620 (N_13620,N_13253,N_13307);
nor U13621 (N_13621,N_13009,N_13050);
or U13622 (N_13622,N_13075,N_13377);
nor U13623 (N_13623,N_13135,N_13298);
nor U13624 (N_13624,N_13114,N_13352);
xor U13625 (N_13625,N_13140,N_13186);
xor U13626 (N_13626,N_13102,N_13192);
or U13627 (N_13627,N_13146,N_13058);
nor U13628 (N_13628,N_13454,N_13494);
xor U13629 (N_13629,N_13043,N_13369);
nand U13630 (N_13630,N_13364,N_13357);
and U13631 (N_13631,N_13082,N_13067);
xnor U13632 (N_13632,N_13242,N_13235);
nand U13633 (N_13633,N_13341,N_13200);
nor U13634 (N_13634,N_13055,N_13163);
xor U13635 (N_13635,N_13241,N_13218);
and U13636 (N_13636,N_13083,N_13325);
nand U13637 (N_13637,N_13220,N_13153);
nand U13638 (N_13638,N_13004,N_13042);
and U13639 (N_13639,N_13132,N_13044);
nand U13640 (N_13640,N_13185,N_13351);
and U13641 (N_13641,N_13052,N_13312);
nor U13642 (N_13642,N_13342,N_13074);
and U13643 (N_13643,N_13065,N_13214);
xor U13644 (N_13644,N_13025,N_13166);
nand U13645 (N_13645,N_13482,N_13077);
xor U13646 (N_13646,N_13203,N_13182);
or U13647 (N_13647,N_13431,N_13396);
nand U13648 (N_13648,N_13314,N_13098);
and U13649 (N_13649,N_13382,N_13090);
nor U13650 (N_13650,N_13243,N_13154);
and U13651 (N_13651,N_13285,N_13417);
and U13652 (N_13652,N_13103,N_13160);
xor U13653 (N_13653,N_13313,N_13409);
nand U13654 (N_13654,N_13289,N_13346);
xnor U13655 (N_13655,N_13239,N_13000);
nand U13656 (N_13656,N_13344,N_13081);
or U13657 (N_13657,N_13260,N_13282);
or U13658 (N_13658,N_13246,N_13326);
and U13659 (N_13659,N_13143,N_13419);
xnor U13660 (N_13660,N_13456,N_13295);
and U13661 (N_13661,N_13070,N_13177);
xnor U13662 (N_13662,N_13256,N_13330);
nor U13663 (N_13663,N_13374,N_13109);
nand U13664 (N_13664,N_13141,N_13398);
or U13665 (N_13665,N_13458,N_13175);
and U13666 (N_13666,N_13134,N_13056);
xnor U13667 (N_13667,N_13348,N_13345);
and U13668 (N_13668,N_13126,N_13015);
nand U13669 (N_13669,N_13252,N_13244);
and U13670 (N_13670,N_13333,N_13276);
nor U13671 (N_13671,N_13099,N_13068);
and U13672 (N_13672,N_13385,N_13497);
nor U13673 (N_13673,N_13309,N_13188);
nand U13674 (N_13674,N_13301,N_13388);
xor U13675 (N_13675,N_13404,N_13167);
and U13676 (N_13676,N_13495,N_13444);
or U13677 (N_13677,N_13478,N_13433);
nor U13678 (N_13678,N_13457,N_13122);
or U13679 (N_13679,N_13092,N_13023);
or U13680 (N_13680,N_13339,N_13149);
nand U13681 (N_13681,N_13113,N_13215);
nor U13682 (N_13682,N_13147,N_13492);
and U13683 (N_13683,N_13335,N_13196);
nand U13684 (N_13684,N_13362,N_13178);
and U13685 (N_13685,N_13272,N_13087);
nand U13686 (N_13686,N_13230,N_13415);
and U13687 (N_13687,N_13164,N_13231);
nor U13688 (N_13688,N_13250,N_13373);
and U13689 (N_13689,N_13328,N_13219);
xor U13690 (N_13690,N_13190,N_13418);
nor U13691 (N_13691,N_13093,N_13279);
and U13692 (N_13692,N_13349,N_13195);
nand U13693 (N_13693,N_13027,N_13347);
or U13694 (N_13694,N_13343,N_13297);
or U13695 (N_13695,N_13280,N_13451);
and U13696 (N_13696,N_13259,N_13356);
xnor U13697 (N_13697,N_13054,N_13317);
nor U13698 (N_13698,N_13037,N_13179);
nor U13699 (N_13699,N_13296,N_13240);
nor U13700 (N_13700,N_13029,N_13394);
nor U13701 (N_13701,N_13390,N_13368);
or U13702 (N_13702,N_13430,N_13078);
nand U13703 (N_13703,N_13191,N_13440);
nand U13704 (N_13704,N_13327,N_13475);
nand U13705 (N_13705,N_13486,N_13108);
nand U13706 (N_13706,N_13206,N_13379);
nor U13707 (N_13707,N_13293,N_13329);
nor U13708 (N_13708,N_13353,N_13174);
and U13709 (N_13709,N_13111,N_13405);
nand U13710 (N_13710,N_13248,N_13323);
or U13711 (N_13711,N_13151,N_13436);
nand U13712 (N_13712,N_13131,N_13120);
xnor U13713 (N_13713,N_13490,N_13421);
nand U13714 (N_13714,N_13375,N_13278);
nor U13715 (N_13715,N_13137,N_13416);
nand U13716 (N_13716,N_13162,N_13169);
xnor U13717 (N_13717,N_13429,N_13026);
xnor U13718 (N_13718,N_13003,N_13205);
xnor U13719 (N_13719,N_13470,N_13439);
and U13720 (N_13720,N_13448,N_13336);
and U13721 (N_13721,N_13479,N_13471);
nor U13722 (N_13722,N_13046,N_13262);
nor U13723 (N_13723,N_13155,N_13306);
nand U13724 (N_13724,N_13006,N_13403);
and U13725 (N_13725,N_13455,N_13222);
nor U13726 (N_13726,N_13213,N_13096);
and U13727 (N_13727,N_13016,N_13366);
xnor U13728 (N_13728,N_13263,N_13493);
nor U13729 (N_13729,N_13484,N_13118);
xnor U13730 (N_13730,N_13438,N_13017);
or U13731 (N_13731,N_13340,N_13461);
xnor U13732 (N_13732,N_13410,N_13091);
xnor U13733 (N_13733,N_13499,N_13257);
nor U13734 (N_13734,N_13363,N_13116);
nand U13735 (N_13735,N_13010,N_13434);
xnor U13736 (N_13736,N_13097,N_13005);
and U13737 (N_13737,N_13228,N_13267);
or U13738 (N_13738,N_13136,N_13198);
nand U13739 (N_13739,N_13229,N_13397);
nor U13740 (N_13740,N_13378,N_13441);
nor U13741 (N_13741,N_13463,N_13480);
or U13742 (N_13742,N_13411,N_13310);
or U13743 (N_13743,N_13426,N_13161);
xor U13744 (N_13744,N_13121,N_13095);
xnor U13745 (N_13745,N_13266,N_13315);
or U13746 (N_13746,N_13053,N_13061);
or U13747 (N_13747,N_13422,N_13408);
nor U13748 (N_13748,N_13386,N_13452);
and U13749 (N_13749,N_13057,N_13173);
xnor U13750 (N_13750,N_13062,N_13260);
nand U13751 (N_13751,N_13205,N_13200);
nor U13752 (N_13752,N_13391,N_13485);
nor U13753 (N_13753,N_13128,N_13052);
or U13754 (N_13754,N_13447,N_13493);
nand U13755 (N_13755,N_13139,N_13190);
or U13756 (N_13756,N_13282,N_13286);
nand U13757 (N_13757,N_13193,N_13156);
and U13758 (N_13758,N_13496,N_13458);
and U13759 (N_13759,N_13116,N_13219);
xnor U13760 (N_13760,N_13325,N_13349);
and U13761 (N_13761,N_13186,N_13337);
xnor U13762 (N_13762,N_13336,N_13182);
or U13763 (N_13763,N_13257,N_13165);
and U13764 (N_13764,N_13067,N_13397);
or U13765 (N_13765,N_13009,N_13018);
or U13766 (N_13766,N_13346,N_13306);
or U13767 (N_13767,N_13306,N_13300);
xnor U13768 (N_13768,N_13481,N_13306);
nand U13769 (N_13769,N_13008,N_13152);
nor U13770 (N_13770,N_13042,N_13399);
and U13771 (N_13771,N_13433,N_13174);
nand U13772 (N_13772,N_13481,N_13214);
and U13773 (N_13773,N_13483,N_13490);
or U13774 (N_13774,N_13284,N_13279);
nand U13775 (N_13775,N_13235,N_13332);
nand U13776 (N_13776,N_13461,N_13257);
xnor U13777 (N_13777,N_13171,N_13475);
or U13778 (N_13778,N_13486,N_13487);
or U13779 (N_13779,N_13329,N_13050);
and U13780 (N_13780,N_13107,N_13317);
nand U13781 (N_13781,N_13258,N_13454);
or U13782 (N_13782,N_13289,N_13034);
nor U13783 (N_13783,N_13021,N_13465);
or U13784 (N_13784,N_13465,N_13134);
and U13785 (N_13785,N_13367,N_13052);
or U13786 (N_13786,N_13057,N_13436);
and U13787 (N_13787,N_13466,N_13468);
xnor U13788 (N_13788,N_13357,N_13422);
and U13789 (N_13789,N_13219,N_13405);
xnor U13790 (N_13790,N_13010,N_13287);
or U13791 (N_13791,N_13079,N_13231);
or U13792 (N_13792,N_13007,N_13093);
nor U13793 (N_13793,N_13236,N_13302);
nand U13794 (N_13794,N_13238,N_13279);
nand U13795 (N_13795,N_13353,N_13225);
or U13796 (N_13796,N_13120,N_13070);
xnor U13797 (N_13797,N_13157,N_13348);
xor U13798 (N_13798,N_13027,N_13367);
nand U13799 (N_13799,N_13217,N_13380);
and U13800 (N_13800,N_13353,N_13056);
and U13801 (N_13801,N_13259,N_13387);
or U13802 (N_13802,N_13155,N_13045);
xor U13803 (N_13803,N_13370,N_13018);
or U13804 (N_13804,N_13444,N_13318);
nor U13805 (N_13805,N_13082,N_13231);
xor U13806 (N_13806,N_13025,N_13114);
nor U13807 (N_13807,N_13471,N_13189);
nor U13808 (N_13808,N_13036,N_13043);
nand U13809 (N_13809,N_13073,N_13477);
and U13810 (N_13810,N_13390,N_13214);
nand U13811 (N_13811,N_13379,N_13020);
xor U13812 (N_13812,N_13123,N_13343);
nor U13813 (N_13813,N_13186,N_13131);
xnor U13814 (N_13814,N_13269,N_13056);
or U13815 (N_13815,N_13463,N_13421);
xnor U13816 (N_13816,N_13084,N_13142);
nand U13817 (N_13817,N_13171,N_13334);
nand U13818 (N_13818,N_13354,N_13240);
xor U13819 (N_13819,N_13110,N_13497);
and U13820 (N_13820,N_13191,N_13451);
xor U13821 (N_13821,N_13453,N_13447);
or U13822 (N_13822,N_13200,N_13037);
or U13823 (N_13823,N_13244,N_13185);
xor U13824 (N_13824,N_13337,N_13417);
xnor U13825 (N_13825,N_13244,N_13112);
or U13826 (N_13826,N_13492,N_13131);
and U13827 (N_13827,N_13190,N_13040);
or U13828 (N_13828,N_13185,N_13050);
nand U13829 (N_13829,N_13104,N_13300);
nand U13830 (N_13830,N_13250,N_13193);
and U13831 (N_13831,N_13099,N_13173);
nand U13832 (N_13832,N_13375,N_13464);
nor U13833 (N_13833,N_13029,N_13281);
nand U13834 (N_13834,N_13441,N_13439);
nor U13835 (N_13835,N_13420,N_13106);
and U13836 (N_13836,N_13210,N_13195);
nand U13837 (N_13837,N_13318,N_13276);
nor U13838 (N_13838,N_13136,N_13484);
nand U13839 (N_13839,N_13332,N_13383);
xor U13840 (N_13840,N_13455,N_13058);
or U13841 (N_13841,N_13279,N_13175);
and U13842 (N_13842,N_13175,N_13249);
nand U13843 (N_13843,N_13106,N_13252);
nor U13844 (N_13844,N_13417,N_13499);
xor U13845 (N_13845,N_13089,N_13347);
nand U13846 (N_13846,N_13051,N_13386);
xnor U13847 (N_13847,N_13491,N_13239);
nand U13848 (N_13848,N_13324,N_13419);
nand U13849 (N_13849,N_13066,N_13208);
or U13850 (N_13850,N_13112,N_13400);
or U13851 (N_13851,N_13174,N_13120);
nand U13852 (N_13852,N_13456,N_13349);
and U13853 (N_13853,N_13272,N_13215);
and U13854 (N_13854,N_13244,N_13350);
xnor U13855 (N_13855,N_13280,N_13494);
nor U13856 (N_13856,N_13346,N_13431);
nor U13857 (N_13857,N_13358,N_13495);
and U13858 (N_13858,N_13252,N_13468);
nand U13859 (N_13859,N_13448,N_13493);
xor U13860 (N_13860,N_13322,N_13047);
xnor U13861 (N_13861,N_13176,N_13130);
and U13862 (N_13862,N_13310,N_13104);
and U13863 (N_13863,N_13234,N_13478);
and U13864 (N_13864,N_13351,N_13003);
nor U13865 (N_13865,N_13294,N_13139);
or U13866 (N_13866,N_13195,N_13380);
or U13867 (N_13867,N_13272,N_13234);
xnor U13868 (N_13868,N_13495,N_13481);
xnor U13869 (N_13869,N_13135,N_13306);
nand U13870 (N_13870,N_13031,N_13131);
or U13871 (N_13871,N_13380,N_13450);
and U13872 (N_13872,N_13490,N_13002);
or U13873 (N_13873,N_13470,N_13458);
or U13874 (N_13874,N_13037,N_13381);
nand U13875 (N_13875,N_13226,N_13179);
nand U13876 (N_13876,N_13095,N_13304);
xnor U13877 (N_13877,N_13275,N_13285);
nand U13878 (N_13878,N_13259,N_13480);
xor U13879 (N_13879,N_13155,N_13404);
nor U13880 (N_13880,N_13367,N_13303);
xor U13881 (N_13881,N_13270,N_13396);
nand U13882 (N_13882,N_13044,N_13329);
nor U13883 (N_13883,N_13184,N_13473);
xor U13884 (N_13884,N_13251,N_13145);
or U13885 (N_13885,N_13372,N_13425);
or U13886 (N_13886,N_13327,N_13182);
xnor U13887 (N_13887,N_13089,N_13103);
xnor U13888 (N_13888,N_13349,N_13035);
xor U13889 (N_13889,N_13314,N_13096);
nand U13890 (N_13890,N_13384,N_13083);
xor U13891 (N_13891,N_13244,N_13264);
nand U13892 (N_13892,N_13022,N_13462);
nor U13893 (N_13893,N_13368,N_13383);
or U13894 (N_13894,N_13310,N_13350);
or U13895 (N_13895,N_13198,N_13000);
or U13896 (N_13896,N_13366,N_13400);
or U13897 (N_13897,N_13468,N_13328);
or U13898 (N_13898,N_13346,N_13031);
nor U13899 (N_13899,N_13341,N_13085);
nand U13900 (N_13900,N_13338,N_13297);
or U13901 (N_13901,N_13493,N_13086);
or U13902 (N_13902,N_13199,N_13310);
nand U13903 (N_13903,N_13012,N_13041);
and U13904 (N_13904,N_13261,N_13164);
xor U13905 (N_13905,N_13121,N_13050);
or U13906 (N_13906,N_13055,N_13344);
nand U13907 (N_13907,N_13344,N_13257);
and U13908 (N_13908,N_13191,N_13495);
xor U13909 (N_13909,N_13291,N_13177);
nor U13910 (N_13910,N_13497,N_13253);
nand U13911 (N_13911,N_13192,N_13183);
nand U13912 (N_13912,N_13376,N_13074);
nand U13913 (N_13913,N_13200,N_13160);
or U13914 (N_13914,N_13095,N_13472);
or U13915 (N_13915,N_13281,N_13461);
nand U13916 (N_13916,N_13087,N_13117);
and U13917 (N_13917,N_13275,N_13099);
nand U13918 (N_13918,N_13186,N_13349);
xnor U13919 (N_13919,N_13100,N_13433);
nor U13920 (N_13920,N_13321,N_13230);
xor U13921 (N_13921,N_13200,N_13172);
or U13922 (N_13922,N_13327,N_13426);
nand U13923 (N_13923,N_13031,N_13259);
nand U13924 (N_13924,N_13049,N_13060);
nor U13925 (N_13925,N_13391,N_13142);
or U13926 (N_13926,N_13228,N_13493);
xnor U13927 (N_13927,N_13112,N_13193);
nor U13928 (N_13928,N_13258,N_13447);
nand U13929 (N_13929,N_13224,N_13455);
nor U13930 (N_13930,N_13019,N_13129);
and U13931 (N_13931,N_13166,N_13217);
xor U13932 (N_13932,N_13222,N_13396);
or U13933 (N_13933,N_13045,N_13091);
nand U13934 (N_13934,N_13301,N_13287);
and U13935 (N_13935,N_13311,N_13147);
xnor U13936 (N_13936,N_13168,N_13486);
nor U13937 (N_13937,N_13430,N_13282);
xor U13938 (N_13938,N_13217,N_13183);
nand U13939 (N_13939,N_13057,N_13416);
nand U13940 (N_13940,N_13184,N_13293);
xor U13941 (N_13941,N_13233,N_13346);
nor U13942 (N_13942,N_13207,N_13404);
or U13943 (N_13943,N_13124,N_13350);
nand U13944 (N_13944,N_13133,N_13050);
and U13945 (N_13945,N_13276,N_13207);
xor U13946 (N_13946,N_13481,N_13477);
or U13947 (N_13947,N_13400,N_13134);
nor U13948 (N_13948,N_13361,N_13321);
nand U13949 (N_13949,N_13252,N_13248);
or U13950 (N_13950,N_13127,N_13309);
and U13951 (N_13951,N_13425,N_13116);
and U13952 (N_13952,N_13435,N_13160);
nand U13953 (N_13953,N_13120,N_13315);
or U13954 (N_13954,N_13094,N_13341);
and U13955 (N_13955,N_13162,N_13013);
or U13956 (N_13956,N_13264,N_13332);
nand U13957 (N_13957,N_13327,N_13384);
xor U13958 (N_13958,N_13137,N_13156);
or U13959 (N_13959,N_13216,N_13256);
xor U13960 (N_13960,N_13446,N_13297);
and U13961 (N_13961,N_13370,N_13050);
xnor U13962 (N_13962,N_13029,N_13010);
or U13963 (N_13963,N_13372,N_13350);
xnor U13964 (N_13964,N_13310,N_13464);
or U13965 (N_13965,N_13129,N_13056);
nand U13966 (N_13966,N_13373,N_13217);
xor U13967 (N_13967,N_13274,N_13066);
and U13968 (N_13968,N_13444,N_13374);
nand U13969 (N_13969,N_13474,N_13373);
nand U13970 (N_13970,N_13382,N_13113);
nor U13971 (N_13971,N_13421,N_13397);
xnor U13972 (N_13972,N_13420,N_13343);
xor U13973 (N_13973,N_13266,N_13189);
nand U13974 (N_13974,N_13407,N_13316);
xor U13975 (N_13975,N_13062,N_13322);
nor U13976 (N_13976,N_13113,N_13338);
or U13977 (N_13977,N_13154,N_13003);
xnor U13978 (N_13978,N_13307,N_13385);
nor U13979 (N_13979,N_13296,N_13404);
nand U13980 (N_13980,N_13357,N_13345);
nor U13981 (N_13981,N_13177,N_13122);
nor U13982 (N_13982,N_13088,N_13246);
or U13983 (N_13983,N_13428,N_13001);
or U13984 (N_13984,N_13418,N_13312);
and U13985 (N_13985,N_13354,N_13498);
or U13986 (N_13986,N_13070,N_13332);
and U13987 (N_13987,N_13220,N_13382);
or U13988 (N_13988,N_13138,N_13319);
xor U13989 (N_13989,N_13416,N_13452);
nor U13990 (N_13990,N_13207,N_13358);
or U13991 (N_13991,N_13142,N_13319);
or U13992 (N_13992,N_13291,N_13020);
nor U13993 (N_13993,N_13107,N_13484);
nand U13994 (N_13994,N_13049,N_13495);
xnor U13995 (N_13995,N_13054,N_13365);
and U13996 (N_13996,N_13138,N_13305);
nor U13997 (N_13997,N_13484,N_13259);
nand U13998 (N_13998,N_13111,N_13446);
nor U13999 (N_13999,N_13080,N_13301);
and U14000 (N_14000,N_13859,N_13624);
nand U14001 (N_14001,N_13844,N_13960);
or U14002 (N_14002,N_13838,N_13807);
and U14003 (N_14003,N_13784,N_13634);
nor U14004 (N_14004,N_13720,N_13598);
and U14005 (N_14005,N_13576,N_13904);
nor U14006 (N_14006,N_13951,N_13759);
or U14007 (N_14007,N_13950,N_13564);
nor U14008 (N_14008,N_13845,N_13881);
or U14009 (N_14009,N_13637,N_13919);
nor U14010 (N_14010,N_13908,N_13544);
xor U14011 (N_14011,N_13945,N_13780);
or U14012 (N_14012,N_13627,N_13548);
nor U14013 (N_14013,N_13873,N_13650);
xnor U14014 (N_14014,N_13591,N_13840);
xnor U14015 (N_14015,N_13594,N_13600);
nand U14016 (N_14016,N_13897,N_13708);
and U14017 (N_14017,N_13741,N_13651);
xnor U14018 (N_14018,N_13864,N_13788);
xnor U14019 (N_14019,N_13882,N_13753);
nor U14020 (N_14020,N_13682,N_13517);
xnor U14021 (N_14021,N_13734,N_13957);
and U14022 (N_14022,N_13641,N_13520);
or U14023 (N_14023,N_13891,N_13901);
nor U14024 (N_14024,N_13586,N_13746);
or U14025 (N_14025,N_13542,N_13553);
xnor U14026 (N_14026,N_13642,N_13690);
nor U14027 (N_14027,N_13561,N_13927);
and U14028 (N_14028,N_13604,N_13850);
xnor U14029 (N_14029,N_13767,N_13718);
or U14030 (N_14030,N_13981,N_13535);
nand U14031 (N_14031,N_13851,N_13810);
nor U14032 (N_14032,N_13808,N_13735);
nand U14033 (N_14033,N_13843,N_13875);
or U14034 (N_14034,N_13648,N_13670);
nor U14035 (N_14035,N_13939,N_13511);
and U14036 (N_14036,N_13884,N_13785);
xor U14037 (N_14037,N_13774,N_13958);
xor U14038 (N_14038,N_13660,N_13584);
nor U14039 (N_14039,N_13905,N_13763);
and U14040 (N_14040,N_13538,N_13698);
nand U14041 (N_14041,N_13953,N_13892);
and U14042 (N_14042,N_13654,N_13940);
nand U14043 (N_14043,N_13912,N_13679);
or U14044 (N_14044,N_13809,N_13828);
or U14045 (N_14045,N_13988,N_13854);
nor U14046 (N_14046,N_13579,N_13781);
nor U14047 (N_14047,N_13563,N_13583);
nor U14048 (N_14048,N_13874,N_13692);
nand U14049 (N_14049,N_13727,N_13573);
nor U14050 (N_14050,N_13929,N_13920);
and U14051 (N_14051,N_13500,N_13972);
xor U14052 (N_14052,N_13688,N_13695);
xnor U14053 (N_14053,N_13524,N_13932);
nand U14054 (N_14054,N_13914,N_13508);
and U14055 (N_14055,N_13903,N_13885);
nor U14056 (N_14056,N_13707,N_13525);
xor U14057 (N_14057,N_13684,N_13752);
xnor U14058 (N_14058,N_13986,N_13714);
nor U14059 (N_14059,N_13536,N_13612);
or U14060 (N_14060,N_13996,N_13628);
nor U14061 (N_14061,N_13504,N_13539);
or U14062 (N_14062,N_13603,N_13755);
and U14063 (N_14063,N_13693,N_13775);
nand U14064 (N_14064,N_13878,N_13963);
nand U14065 (N_14065,N_13617,N_13622);
and U14066 (N_14066,N_13805,N_13938);
nand U14067 (N_14067,N_13546,N_13537);
xor U14068 (N_14068,N_13956,N_13609);
and U14069 (N_14069,N_13635,N_13893);
xor U14070 (N_14070,N_13765,N_13822);
and U14071 (N_14071,N_13747,N_13979);
nor U14072 (N_14072,N_13502,N_13771);
xor U14073 (N_14073,N_13991,N_13769);
or U14074 (N_14074,N_13661,N_13918);
xnor U14075 (N_14075,N_13976,N_13970);
xnor U14076 (N_14076,N_13751,N_13614);
and U14077 (N_14077,N_13899,N_13709);
nand U14078 (N_14078,N_13526,N_13801);
or U14079 (N_14079,N_13619,N_13968);
nor U14080 (N_14080,N_13889,N_13560);
and U14081 (N_14081,N_13719,N_13566);
or U14082 (N_14082,N_13944,N_13620);
and U14083 (N_14083,N_13898,N_13621);
xor U14084 (N_14084,N_13832,N_13866);
xor U14085 (N_14085,N_13954,N_13795);
nand U14086 (N_14086,N_13552,N_13570);
or U14087 (N_14087,N_13503,N_13978);
or U14088 (N_14088,N_13772,N_13662);
nor U14089 (N_14089,N_13501,N_13879);
nand U14090 (N_14090,N_13565,N_13597);
xnor U14091 (N_14091,N_13923,N_13649);
xnor U14092 (N_14092,N_13916,N_13791);
and U14093 (N_14093,N_13802,N_13992);
nand U14094 (N_14094,N_13855,N_13729);
nand U14095 (N_14095,N_13962,N_13982);
or U14096 (N_14096,N_13626,N_13789);
nor U14097 (N_14097,N_13636,N_13611);
or U14098 (N_14098,N_13578,N_13607);
nand U14099 (N_14099,N_13739,N_13925);
or U14100 (N_14100,N_13815,N_13906);
and U14101 (N_14101,N_13625,N_13750);
nor U14102 (N_14102,N_13724,N_13588);
xor U14103 (N_14103,N_13702,N_13645);
xnor U14104 (N_14104,N_13581,N_13616);
or U14105 (N_14105,N_13731,N_13993);
nand U14106 (N_14106,N_13744,N_13847);
or U14107 (N_14107,N_13715,N_13639);
nand U14108 (N_14108,N_13704,N_13575);
xnor U14109 (N_14109,N_13913,N_13673);
nand U14110 (N_14110,N_13778,N_13915);
xnor U14111 (N_14111,N_13934,N_13936);
or U14112 (N_14112,N_13999,N_13605);
nand U14113 (N_14113,N_13506,N_13608);
nand U14114 (N_14114,N_13694,N_13633);
or U14115 (N_14115,N_13726,N_13928);
nand U14116 (N_14116,N_13745,N_13658);
or U14117 (N_14117,N_13532,N_13521);
nand U14118 (N_14118,N_13687,N_13852);
nor U14119 (N_14119,N_13700,N_13768);
xnor U14120 (N_14120,N_13568,N_13530);
or U14121 (N_14121,N_13678,N_13967);
xor U14122 (N_14122,N_13665,N_13623);
and U14123 (N_14123,N_13722,N_13712);
nand U14124 (N_14124,N_13868,N_13723);
or U14125 (N_14125,N_13937,N_13857);
nor U14126 (N_14126,N_13887,N_13653);
and U14127 (N_14127,N_13652,N_13699);
nor U14128 (N_14128,N_13748,N_13933);
and U14129 (N_14129,N_13816,N_13827);
nand U14130 (N_14130,N_13674,N_13531);
and U14131 (N_14131,N_13518,N_13523);
or U14132 (N_14132,N_13860,N_13743);
or U14133 (N_14133,N_13580,N_13942);
nor U14134 (N_14134,N_13514,N_13814);
nand U14135 (N_14135,N_13691,N_13762);
nand U14136 (N_14136,N_13717,N_13921);
and U14137 (N_14137,N_13592,N_13664);
nor U14138 (N_14138,N_13911,N_13671);
nor U14139 (N_14139,N_13959,N_13812);
or U14140 (N_14140,N_13629,N_13640);
or U14141 (N_14141,N_13943,N_13711);
nand U14142 (N_14142,N_13596,N_13948);
nand U14143 (N_14143,N_13754,N_13657);
xnor U14144 (N_14144,N_13835,N_13736);
nand U14145 (N_14145,N_13955,N_13819);
and U14146 (N_14146,N_13601,N_13764);
and U14147 (N_14147,N_13541,N_13632);
nor U14148 (N_14148,N_13522,N_13817);
nor U14149 (N_14149,N_13585,N_13783);
xor U14150 (N_14150,N_13766,N_13924);
or U14151 (N_14151,N_13848,N_13556);
or U14152 (N_14152,N_13610,N_13683);
or U14153 (N_14153,N_13703,N_13829);
and U14154 (N_14154,N_13527,N_13836);
xnor U14155 (N_14155,N_13572,N_13900);
nand U14156 (N_14156,N_13862,N_13550);
and U14157 (N_14157,N_13985,N_13760);
nor U14158 (N_14158,N_13567,N_13888);
or U14159 (N_14159,N_13587,N_13507);
nand U14160 (N_14160,N_13926,N_13883);
nor U14161 (N_14161,N_13738,N_13730);
xnor U14162 (N_14162,N_13890,N_13515);
nand U14163 (N_14163,N_13902,N_13757);
and U14164 (N_14164,N_13895,N_13706);
nand U14165 (N_14165,N_13630,N_13554);
or U14166 (N_14166,N_13680,N_13713);
nor U14167 (N_14167,N_13803,N_13725);
xnor U14168 (N_14168,N_13646,N_13681);
xnor U14169 (N_14169,N_13797,N_13677);
nand U14170 (N_14170,N_13533,N_13647);
or U14171 (N_14171,N_13540,N_13615);
xnor U14172 (N_14172,N_13577,N_13510);
nor U14173 (N_14173,N_13995,N_13589);
nand U14174 (N_14174,N_13973,N_13742);
and U14175 (N_14175,N_13672,N_13790);
or U14176 (N_14176,N_13606,N_13971);
and U14177 (N_14177,N_13994,N_13872);
and U14178 (N_14178,N_13952,N_13516);
and U14179 (N_14179,N_13716,N_13728);
xnor U14180 (N_14180,N_13941,N_13831);
nor U14181 (N_14181,N_13770,N_13909);
nand U14182 (N_14182,N_13974,N_13977);
or U14183 (N_14183,N_13989,N_13799);
nand U14184 (N_14184,N_13946,N_13761);
nor U14185 (N_14185,N_13798,N_13867);
or U14186 (N_14186,N_13569,N_13666);
and U14187 (N_14187,N_13964,N_13571);
or U14188 (N_14188,N_13935,N_13787);
and U14189 (N_14189,N_13907,N_13710);
xor U14190 (N_14190,N_13701,N_13930);
nand U14191 (N_14191,N_13830,N_13676);
or U14192 (N_14192,N_13837,N_13667);
and U14193 (N_14193,N_13846,N_13547);
xor U14194 (N_14194,N_13794,N_13998);
nand U14195 (N_14195,N_13777,N_13980);
and U14196 (N_14196,N_13689,N_13910);
and U14197 (N_14197,N_13821,N_13732);
nand U14198 (N_14198,N_13758,N_13749);
or U14199 (N_14199,N_13686,N_13824);
nor U14200 (N_14200,N_13969,N_13559);
or U14201 (N_14201,N_13655,N_13638);
and U14202 (N_14202,N_13590,N_13593);
nand U14203 (N_14203,N_13792,N_13644);
or U14204 (N_14204,N_13669,N_13631);
xnor U14205 (N_14205,N_13705,N_13733);
xor U14206 (N_14206,N_13782,N_13618);
and U14207 (N_14207,N_13833,N_13856);
nor U14208 (N_14208,N_13820,N_13549);
xnor U14209 (N_14209,N_13534,N_13961);
and U14210 (N_14210,N_13543,N_13779);
and U14211 (N_14211,N_13786,N_13990);
nand U14212 (N_14212,N_13965,N_13551);
or U14213 (N_14213,N_13613,N_13931);
or U14214 (N_14214,N_13825,N_13894);
and U14215 (N_14215,N_13839,N_13853);
xor U14216 (N_14216,N_13983,N_13505);
nand U14217 (N_14217,N_13582,N_13917);
or U14218 (N_14218,N_13877,N_13984);
and U14219 (N_14219,N_13737,N_13555);
nor U14220 (N_14220,N_13513,N_13826);
nand U14221 (N_14221,N_13880,N_13796);
xnor U14222 (N_14222,N_13813,N_13886);
or U14223 (N_14223,N_13922,N_13599);
or U14224 (N_14224,N_13557,N_13756);
or U14225 (N_14225,N_13602,N_13947);
nand U14226 (N_14226,N_13528,N_13987);
or U14227 (N_14227,N_13776,N_13834);
and U14228 (N_14228,N_13818,N_13849);
or U14229 (N_14229,N_13806,N_13800);
xnor U14230 (N_14230,N_13870,N_13869);
nor U14231 (N_14231,N_13842,N_13793);
nor U14232 (N_14232,N_13519,N_13896);
or U14233 (N_14233,N_13858,N_13966);
or U14234 (N_14234,N_13975,N_13529);
nand U14235 (N_14235,N_13663,N_13656);
nor U14236 (N_14236,N_13696,N_13740);
or U14237 (N_14237,N_13823,N_13997);
nor U14238 (N_14238,N_13949,N_13643);
and U14239 (N_14239,N_13512,N_13871);
or U14240 (N_14240,N_13773,N_13697);
or U14241 (N_14241,N_13558,N_13545);
xnor U14242 (N_14242,N_13562,N_13574);
and U14243 (N_14243,N_13876,N_13861);
nand U14244 (N_14244,N_13509,N_13863);
nand U14245 (N_14245,N_13841,N_13685);
xnor U14246 (N_14246,N_13595,N_13865);
or U14247 (N_14247,N_13721,N_13811);
nor U14248 (N_14248,N_13804,N_13668);
nor U14249 (N_14249,N_13675,N_13659);
xnor U14250 (N_14250,N_13522,N_13693);
nor U14251 (N_14251,N_13620,N_13873);
or U14252 (N_14252,N_13520,N_13777);
xnor U14253 (N_14253,N_13675,N_13507);
or U14254 (N_14254,N_13844,N_13780);
nand U14255 (N_14255,N_13786,N_13704);
and U14256 (N_14256,N_13652,N_13910);
nor U14257 (N_14257,N_13674,N_13992);
nand U14258 (N_14258,N_13910,N_13916);
or U14259 (N_14259,N_13705,N_13970);
and U14260 (N_14260,N_13949,N_13850);
nand U14261 (N_14261,N_13851,N_13825);
or U14262 (N_14262,N_13569,N_13546);
nor U14263 (N_14263,N_13729,N_13926);
nor U14264 (N_14264,N_13581,N_13670);
or U14265 (N_14265,N_13845,N_13627);
or U14266 (N_14266,N_13803,N_13614);
xor U14267 (N_14267,N_13956,N_13506);
xor U14268 (N_14268,N_13681,N_13701);
nand U14269 (N_14269,N_13853,N_13889);
nor U14270 (N_14270,N_13612,N_13531);
nand U14271 (N_14271,N_13883,N_13861);
nor U14272 (N_14272,N_13572,N_13884);
xnor U14273 (N_14273,N_13761,N_13650);
nand U14274 (N_14274,N_13535,N_13686);
and U14275 (N_14275,N_13818,N_13535);
nand U14276 (N_14276,N_13594,N_13659);
xor U14277 (N_14277,N_13720,N_13663);
nor U14278 (N_14278,N_13930,N_13756);
nand U14279 (N_14279,N_13910,N_13590);
and U14280 (N_14280,N_13966,N_13667);
nor U14281 (N_14281,N_13610,N_13547);
xor U14282 (N_14282,N_13715,N_13559);
nor U14283 (N_14283,N_13506,N_13714);
nor U14284 (N_14284,N_13624,N_13536);
xor U14285 (N_14285,N_13837,N_13546);
xor U14286 (N_14286,N_13618,N_13979);
xnor U14287 (N_14287,N_13909,N_13874);
nor U14288 (N_14288,N_13900,N_13664);
or U14289 (N_14289,N_13823,N_13660);
or U14290 (N_14290,N_13599,N_13920);
or U14291 (N_14291,N_13737,N_13738);
nor U14292 (N_14292,N_13959,N_13940);
or U14293 (N_14293,N_13595,N_13858);
and U14294 (N_14294,N_13857,N_13887);
xor U14295 (N_14295,N_13740,N_13797);
nor U14296 (N_14296,N_13541,N_13918);
or U14297 (N_14297,N_13752,N_13799);
xnor U14298 (N_14298,N_13772,N_13656);
and U14299 (N_14299,N_13579,N_13562);
xnor U14300 (N_14300,N_13979,N_13973);
nor U14301 (N_14301,N_13565,N_13919);
nor U14302 (N_14302,N_13598,N_13708);
xor U14303 (N_14303,N_13983,N_13657);
nand U14304 (N_14304,N_13802,N_13664);
nand U14305 (N_14305,N_13533,N_13922);
nor U14306 (N_14306,N_13854,N_13935);
nand U14307 (N_14307,N_13882,N_13547);
and U14308 (N_14308,N_13979,N_13514);
nor U14309 (N_14309,N_13938,N_13674);
and U14310 (N_14310,N_13883,N_13648);
and U14311 (N_14311,N_13630,N_13584);
and U14312 (N_14312,N_13991,N_13973);
nor U14313 (N_14313,N_13936,N_13975);
nor U14314 (N_14314,N_13551,N_13891);
and U14315 (N_14315,N_13875,N_13783);
xnor U14316 (N_14316,N_13690,N_13500);
and U14317 (N_14317,N_13930,N_13557);
xor U14318 (N_14318,N_13987,N_13919);
nor U14319 (N_14319,N_13920,N_13702);
and U14320 (N_14320,N_13958,N_13538);
or U14321 (N_14321,N_13797,N_13991);
and U14322 (N_14322,N_13640,N_13677);
and U14323 (N_14323,N_13940,N_13592);
xnor U14324 (N_14324,N_13849,N_13509);
nand U14325 (N_14325,N_13659,N_13948);
or U14326 (N_14326,N_13882,N_13861);
nand U14327 (N_14327,N_13625,N_13984);
nand U14328 (N_14328,N_13575,N_13965);
and U14329 (N_14329,N_13722,N_13794);
or U14330 (N_14330,N_13945,N_13938);
and U14331 (N_14331,N_13658,N_13607);
nor U14332 (N_14332,N_13834,N_13908);
xnor U14333 (N_14333,N_13916,N_13948);
or U14334 (N_14334,N_13519,N_13989);
nand U14335 (N_14335,N_13974,N_13616);
and U14336 (N_14336,N_13621,N_13730);
or U14337 (N_14337,N_13811,N_13642);
and U14338 (N_14338,N_13948,N_13811);
nand U14339 (N_14339,N_13777,N_13664);
nor U14340 (N_14340,N_13513,N_13862);
nand U14341 (N_14341,N_13805,N_13708);
nor U14342 (N_14342,N_13524,N_13806);
or U14343 (N_14343,N_13773,N_13502);
or U14344 (N_14344,N_13753,N_13942);
or U14345 (N_14345,N_13879,N_13816);
nor U14346 (N_14346,N_13717,N_13779);
nor U14347 (N_14347,N_13570,N_13594);
nor U14348 (N_14348,N_13763,N_13677);
and U14349 (N_14349,N_13963,N_13911);
nor U14350 (N_14350,N_13738,N_13868);
and U14351 (N_14351,N_13666,N_13860);
nand U14352 (N_14352,N_13551,N_13738);
or U14353 (N_14353,N_13810,N_13717);
and U14354 (N_14354,N_13696,N_13545);
nor U14355 (N_14355,N_13520,N_13563);
and U14356 (N_14356,N_13754,N_13615);
xor U14357 (N_14357,N_13631,N_13556);
xor U14358 (N_14358,N_13530,N_13679);
xnor U14359 (N_14359,N_13951,N_13950);
nor U14360 (N_14360,N_13977,N_13693);
xnor U14361 (N_14361,N_13614,N_13801);
or U14362 (N_14362,N_13947,N_13603);
xnor U14363 (N_14363,N_13932,N_13545);
nor U14364 (N_14364,N_13601,N_13977);
nand U14365 (N_14365,N_13785,N_13555);
and U14366 (N_14366,N_13627,N_13729);
and U14367 (N_14367,N_13998,N_13523);
or U14368 (N_14368,N_13739,N_13841);
or U14369 (N_14369,N_13904,N_13617);
xor U14370 (N_14370,N_13787,N_13992);
nor U14371 (N_14371,N_13827,N_13725);
or U14372 (N_14372,N_13655,N_13737);
or U14373 (N_14373,N_13942,N_13988);
and U14374 (N_14374,N_13995,N_13614);
nor U14375 (N_14375,N_13543,N_13816);
or U14376 (N_14376,N_13699,N_13555);
nand U14377 (N_14377,N_13614,N_13930);
nor U14378 (N_14378,N_13636,N_13536);
nor U14379 (N_14379,N_13903,N_13982);
and U14380 (N_14380,N_13935,N_13691);
or U14381 (N_14381,N_13775,N_13544);
and U14382 (N_14382,N_13921,N_13531);
and U14383 (N_14383,N_13545,N_13793);
or U14384 (N_14384,N_13634,N_13972);
nand U14385 (N_14385,N_13941,N_13652);
nand U14386 (N_14386,N_13867,N_13528);
nand U14387 (N_14387,N_13994,N_13771);
and U14388 (N_14388,N_13946,N_13892);
nor U14389 (N_14389,N_13637,N_13947);
xor U14390 (N_14390,N_13590,N_13746);
xnor U14391 (N_14391,N_13528,N_13787);
nor U14392 (N_14392,N_13946,N_13704);
or U14393 (N_14393,N_13508,N_13911);
or U14394 (N_14394,N_13612,N_13518);
xor U14395 (N_14395,N_13789,N_13587);
and U14396 (N_14396,N_13926,N_13708);
or U14397 (N_14397,N_13651,N_13601);
or U14398 (N_14398,N_13629,N_13978);
or U14399 (N_14399,N_13707,N_13629);
nor U14400 (N_14400,N_13569,N_13820);
nand U14401 (N_14401,N_13556,N_13593);
nand U14402 (N_14402,N_13901,N_13538);
nand U14403 (N_14403,N_13656,N_13931);
nand U14404 (N_14404,N_13882,N_13647);
xnor U14405 (N_14405,N_13560,N_13654);
or U14406 (N_14406,N_13983,N_13626);
nor U14407 (N_14407,N_13649,N_13963);
or U14408 (N_14408,N_13866,N_13907);
xor U14409 (N_14409,N_13981,N_13506);
and U14410 (N_14410,N_13634,N_13753);
xor U14411 (N_14411,N_13561,N_13518);
xnor U14412 (N_14412,N_13727,N_13664);
or U14413 (N_14413,N_13877,N_13965);
and U14414 (N_14414,N_13846,N_13665);
or U14415 (N_14415,N_13862,N_13610);
xnor U14416 (N_14416,N_13774,N_13596);
and U14417 (N_14417,N_13595,N_13583);
and U14418 (N_14418,N_13671,N_13734);
nor U14419 (N_14419,N_13912,N_13654);
xor U14420 (N_14420,N_13726,N_13607);
xor U14421 (N_14421,N_13878,N_13944);
xor U14422 (N_14422,N_13607,N_13840);
or U14423 (N_14423,N_13739,N_13746);
xor U14424 (N_14424,N_13878,N_13964);
xor U14425 (N_14425,N_13849,N_13584);
and U14426 (N_14426,N_13763,N_13860);
and U14427 (N_14427,N_13750,N_13937);
xor U14428 (N_14428,N_13618,N_13666);
xor U14429 (N_14429,N_13964,N_13580);
nand U14430 (N_14430,N_13704,N_13647);
and U14431 (N_14431,N_13655,N_13713);
and U14432 (N_14432,N_13592,N_13856);
nand U14433 (N_14433,N_13729,N_13678);
and U14434 (N_14434,N_13937,N_13631);
or U14435 (N_14435,N_13561,N_13953);
nor U14436 (N_14436,N_13816,N_13652);
or U14437 (N_14437,N_13897,N_13537);
nand U14438 (N_14438,N_13963,N_13992);
xnor U14439 (N_14439,N_13585,N_13929);
xnor U14440 (N_14440,N_13657,N_13664);
nand U14441 (N_14441,N_13788,N_13922);
or U14442 (N_14442,N_13999,N_13652);
or U14443 (N_14443,N_13838,N_13560);
or U14444 (N_14444,N_13951,N_13736);
or U14445 (N_14445,N_13538,N_13709);
nor U14446 (N_14446,N_13509,N_13728);
xnor U14447 (N_14447,N_13965,N_13678);
nor U14448 (N_14448,N_13915,N_13933);
nor U14449 (N_14449,N_13948,N_13910);
nor U14450 (N_14450,N_13639,N_13528);
or U14451 (N_14451,N_13536,N_13725);
nor U14452 (N_14452,N_13617,N_13832);
xnor U14453 (N_14453,N_13896,N_13761);
and U14454 (N_14454,N_13507,N_13767);
or U14455 (N_14455,N_13757,N_13626);
or U14456 (N_14456,N_13868,N_13853);
or U14457 (N_14457,N_13692,N_13614);
or U14458 (N_14458,N_13942,N_13522);
or U14459 (N_14459,N_13953,N_13606);
and U14460 (N_14460,N_13745,N_13520);
nand U14461 (N_14461,N_13679,N_13972);
or U14462 (N_14462,N_13541,N_13858);
or U14463 (N_14463,N_13526,N_13667);
xor U14464 (N_14464,N_13565,N_13500);
xnor U14465 (N_14465,N_13969,N_13978);
xor U14466 (N_14466,N_13582,N_13745);
or U14467 (N_14467,N_13701,N_13944);
xor U14468 (N_14468,N_13787,N_13519);
and U14469 (N_14469,N_13908,N_13718);
or U14470 (N_14470,N_13519,N_13502);
or U14471 (N_14471,N_13835,N_13772);
xor U14472 (N_14472,N_13842,N_13853);
nor U14473 (N_14473,N_13868,N_13990);
nor U14474 (N_14474,N_13826,N_13552);
nand U14475 (N_14475,N_13823,N_13871);
or U14476 (N_14476,N_13722,N_13825);
and U14477 (N_14477,N_13841,N_13831);
nand U14478 (N_14478,N_13872,N_13680);
nand U14479 (N_14479,N_13699,N_13858);
and U14480 (N_14480,N_13816,N_13500);
or U14481 (N_14481,N_13602,N_13607);
nand U14482 (N_14482,N_13987,N_13719);
nand U14483 (N_14483,N_13531,N_13557);
nor U14484 (N_14484,N_13500,N_13867);
nand U14485 (N_14485,N_13721,N_13943);
xor U14486 (N_14486,N_13546,N_13824);
and U14487 (N_14487,N_13868,N_13741);
xor U14488 (N_14488,N_13883,N_13754);
and U14489 (N_14489,N_13645,N_13501);
xor U14490 (N_14490,N_13534,N_13738);
xor U14491 (N_14491,N_13844,N_13618);
or U14492 (N_14492,N_13626,N_13645);
nor U14493 (N_14493,N_13819,N_13531);
and U14494 (N_14494,N_13854,N_13653);
or U14495 (N_14495,N_13903,N_13806);
nor U14496 (N_14496,N_13732,N_13988);
and U14497 (N_14497,N_13945,N_13951);
nor U14498 (N_14498,N_13569,N_13866);
or U14499 (N_14499,N_13780,N_13831);
or U14500 (N_14500,N_14260,N_14414);
nor U14501 (N_14501,N_14055,N_14274);
nor U14502 (N_14502,N_14167,N_14486);
nor U14503 (N_14503,N_14023,N_14233);
or U14504 (N_14504,N_14273,N_14460);
or U14505 (N_14505,N_14066,N_14162);
and U14506 (N_14506,N_14223,N_14176);
or U14507 (N_14507,N_14391,N_14296);
xnor U14508 (N_14508,N_14267,N_14427);
nor U14509 (N_14509,N_14089,N_14229);
or U14510 (N_14510,N_14006,N_14417);
nor U14511 (N_14511,N_14111,N_14234);
and U14512 (N_14512,N_14336,N_14333);
and U14513 (N_14513,N_14377,N_14413);
nand U14514 (N_14514,N_14497,N_14283);
and U14515 (N_14515,N_14096,N_14416);
nor U14516 (N_14516,N_14489,N_14115);
and U14517 (N_14517,N_14249,N_14094);
xor U14518 (N_14518,N_14087,N_14065);
nand U14519 (N_14519,N_14280,N_14491);
or U14520 (N_14520,N_14330,N_14247);
nand U14521 (N_14521,N_14258,N_14105);
xor U14522 (N_14522,N_14161,N_14129);
and U14523 (N_14523,N_14194,N_14048);
nor U14524 (N_14524,N_14085,N_14300);
nor U14525 (N_14525,N_14043,N_14073);
and U14526 (N_14526,N_14181,N_14084);
nor U14527 (N_14527,N_14057,N_14356);
xnor U14528 (N_14528,N_14437,N_14131);
or U14529 (N_14529,N_14360,N_14468);
and U14530 (N_14530,N_14086,N_14464);
nand U14531 (N_14531,N_14415,N_14425);
xor U14532 (N_14532,N_14494,N_14294);
nor U14533 (N_14533,N_14047,N_14244);
or U14534 (N_14534,N_14466,N_14275);
nand U14535 (N_14535,N_14319,N_14257);
and U14536 (N_14536,N_14371,N_14216);
and U14537 (N_14537,N_14374,N_14357);
xor U14538 (N_14538,N_14403,N_14237);
xnor U14539 (N_14539,N_14235,N_14017);
or U14540 (N_14540,N_14116,N_14003);
nand U14541 (N_14541,N_14386,N_14035);
and U14542 (N_14542,N_14350,N_14384);
nor U14543 (N_14543,N_14262,N_14240);
nand U14544 (N_14544,N_14304,N_14478);
and U14545 (N_14545,N_14245,N_14124);
nand U14546 (N_14546,N_14156,N_14232);
and U14547 (N_14547,N_14355,N_14075);
xnor U14548 (N_14548,N_14447,N_14405);
nand U14549 (N_14549,N_14288,N_14038);
nand U14550 (N_14550,N_14496,N_14482);
and U14551 (N_14551,N_14428,N_14099);
and U14552 (N_14552,N_14469,N_14007);
nand U14553 (N_14553,N_14198,N_14227);
or U14554 (N_14554,N_14254,N_14297);
nor U14555 (N_14555,N_14163,N_14347);
xnor U14556 (N_14556,N_14081,N_14343);
nor U14557 (N_14557,N_14175,N_14338);
xnor U14558 (N_14558,N_14327,N_14404);
nor U14559 (N_14559,N_14207,N_14430);
nor U14560 (N_14560,N_14444,N_14074);
nand U14561 (N_14561,N_14160,N_14222);
or U14562 (N_14562,N_14445,N_14465);
nand U14563 (N_14563,N_14044,N_14231);
nor U14564 (N_14564,N_14368,N_14166);
nand U14565 (N_14565,N_14461,N_14359);
or U14566 (N_14566,N_14046,N_14266);
xor U14567 (N_14567,N_14100,N_14412);
xor U14568 (N_14568,N_14389,N_14120);
nand U14569 (N_14569,N_14097,N_14189);
or U14570 (N_14570,N_14011,N_14353);
nand U14571 (N_14571,N_14316,N_14031);
xnor U14572 (N_14572,N_14130,N_14248);
nand U14573 (N_14573,N_14209,N_14337);
or U14574 (N_14574,N_14381,N_14481);
nor U14575 (N_14575,N_14148,N_14400);
nor U14576 (N_14576,N_14424,N_14242);
or U14577 (N_14577,N_14180,N_14383);
and U14578 (N_14578,N_14463,N_14206);
nand U14579 (N_14579,N_14341,N_14291);
xor U14580 (N_14580,N_14236,N_14265);
and U14581 (N_14581,N_14268,N_14184);
and U14582 (N_14582,N_14168,N_14363);
and U14583 (N_14583,N_14070,N_14431);
or U14584 (N_14584,N_14433,N_14448);
nand U14585 (N_14585,N_14002,N_14113);
nor U14586 (N_14586,N_14018,N_14078);
nand U14587 (N_14587,N_14419,N_14495);
nor U14588 (N_14588,N_14479,N_14451);
or U14589 (N_14589,N_14118,N_14421);
and U14590 (N_14590,N_14058,N_14332);
xor U14591 (N_14591,N_14467,N_14435);
nand U14592 (N_14592,N_14345,N_14201);
or U14593 (N_14593,N_14178,N_14114);
nor U14594 (N_14594,N_14393,N_14107);
xnor U14595 (N_14595,N_14224,N_14325);
nand U14596 (N_14596,N_14348,N_14193);
or U14597 (N_14597,N_14137,N_14072);
nand U14598 (N_14598,N_14225,N_14128);
and U14599 (N_14599,N_14269,N_14033);
or U14600 (N_14600,N_14351,N_14387);
nand U14601 (N_14601,N_14364,N_14378);
and U14602 (N_14602,N_14195,N_14256);
or U14603 (N_14603,N_14082,N_14395);
and U14604 (N_14604,N_14090,N_14152);
nand U14605 (N_14605,N_14052,N_14138);
and U14606 (N_14606,N_14213,N_14077);
or U14607 (N_14607,N_14487,N_14014);
and U14608 (N_14608,N_14476,N_14230);
or U14609 (N_14609,N_14191,N_14239);
nand U14610 (N_14610,N_14165,N_14313);
xor U14611 (N_14611,N_14335,N_14408);
and U14612 (N_14612,N_14020,N_14289);
or U14613 (N_14613,N_14396,N_14228);
nor U14614 (N_14614,N_14310,N_14443);
and U14615 (N_14615,N_14358,N_14344);
and U14616 (N_14616,N_14346,N_14342);
or U14617 (N_14617,N_14025,N_14446);
and U14618 (N_14618,N_14001,N_14205);
nor U14619 (N_14619,N_14154,N_14170);
or U14620 (N_14620,N_14314,N_14411);
xor U14621 (N_14621,N_14136,N_14286);
nand U14622 (N_14622,N_14034,N_14454);
or U14623 (N_14623,N_14027,N_14320);
nand U14624 (N_14624,N_14158,N_14135);
or U14625 (N_14625,N_14188,N_14270);
or U14626 (N_14626,N_14369,N_14423);
or U14627 (N_14627,N_14076,N_14329);
nand U14628 (N_14628,N_14155,N_14362);
or U14629 (N_14629,N_14040,N_14054);
xnor U14630 (N_14630,N_14109,N_14009);
nor U14631 (N_14631,N_14410,N_14452);
xor U14632 (N_14632,N_14302,N_14303);
nor U14633 (N_14633,N_14484,N_14474);
nand U14634 (N_14634,N_14261,N_14279);
nand U14635 (N_14635,N_14490,N_14071);
nand U14636 (N_14636,N_14278,N_14005);
or U14637 (N_14637,N_14305,N_14104);
nor U14638 (N_14638,N_14241,N_14331);
nand U14639 (N_14639,N_14064,N_14141);
xor U14640 (N_14640,N_14068,N_14293);
and U14641 (N_14641,N_14264,N_14488);
nand U14642 (N_14642,N_14028,N_14015);
xnor U14643 (N_14643,N_14458,N_14106);
xnor U14644 (N_14644,N_14203,N_14485);
nand U14645 (N_14645,N_14311,N_14470);
or U14646 (N_14646,N_14016,N_14182);
or U14647 (N_14647,N_14091,N_14441);
xor U14648 (N_14648,N_14146,N_14164);
or U14649 (N_14649,N_14409,N_14063);
nand U14650 (N_14650,N_14008,N_14246);
xor U14651 (N_14651,N_14051,N_14185);
xnor U14652 (N_14652,N_14093,N_14208);
and U14653 (N_14653,N_14459,N_14127);
nand U14654 (N_14654,N_14322,N_14402);
nor U14655 (N_14655,N_14036,N_14455);
or U14656 (N_14656,N_14492,N_14462);
nor U14657 (N_14657,N_14321,N_14438);
and U14658 (N_14658,N_14143,N_14498);
and U14659 (N_14659,N_14112,N_14376);
xor U14660 (N_14660,N_14049,N_14149);
nand U14661 (N_14661,N_14394,N_14295);
or U14662 (N_14662,N_14108,N_14010);
and U14663 (N_14663,N_14039,N_14192);
xor U14664 (N_14664,N_14315,N_14067);
and U14665 (N_14665,N_14339,N_14250);
xor U14666 (N_14666,N_14281,N_14217);
and U14667 (N_14667,N_14019,N_14285);
nand U14668 (N_14668,N_14397,N_14179);
nand U14669 (N_14669,N_14432,N_14282);
or U14670 (N_14670,N_14110,N_14334);
nand U14671 (N_14671,N_14436,N_14069);
xnor U14672 (N_14672,N_14349,N_14379);
xor U14673 (N_14673,N_14226,N_14151);
and U14674 (N_14674,N_14183,N_14398);
or U14675 (N_14675,N_14061,N_14045);
xnor U14676 (N_14676,N_14050,N_14126);
xnor U14677 (N_14677,N_14053,N_14317);
and U14678 (N_14678,N_14062,N_14060);
xor U14679 (N_14679,N_14101,N_14340);
or U14680 (N_14680,N_14290,N_14292);
and U14681 (N_14681,N_14312,N_14453);
nor U14682 (N_14682,N_14032,N_14287);
or U14683 (N_14683,N_14238,N_14449);
or U14684 (N_14684,N_14121,N_14095);
or U14685 (N_14685,N_14259,N_14041);
and U14686 (N_14686,N_14480,N_14299);
or U14687 (N_14687,N_14388,N_14399);
and U14688 (N_14688,N_14243,N_14134);
nand U14689 (N_14689,N_14493,N_14221);
and U14690 (N_14690,N_14380,N_14373);
nand U14691 (N_14691,N_14471,N_14171);
nor U14692 (N_14692,N_14307,N_14122);
xor U14693 (N_14693,N_14326,N_14169);
or U14694 (N_14694,N_14210,N_14301);
xnor U14695 (N_14695,N_14390,N_14277);
or U14696 (N_14696,N_14150,N_14013);
xor U14697 (N_14697,N_14123,N_14361);
and U14698 (N_14698,N_14098,N_14026);
nor U14699 (N_14699,N_14024,N_14103);
nand U14700 (N_14700,N_14457,N_14215);
nand U14701 (N_14701,N_14092,N_14173);
nand U14702 (N_14702,N_14426,N_14139);
nand U14703 (N_14703,N_14144,N_14407);
or U14704 (N_14704,N_14088,N_14477);
xor U14705 (N_14705,N_14372,N_14367);
xnor U14706 (N_14706,N_14125,N_14174);
nand U14707 (N_14707,N_14132,N_14366);
nor U14708 (N_14708,N_14142,N_14153);
and U14709 (N_14709,N_14197,N_14187);
nand U14710 (N_14710,N_14420,N_14177);
nor U14711 (N_14711,N_14418,N_14204);
nor U14712 (N_14712,N_14309,N_14080);
nand U14713 (N_14713,N_14255,N_14021);
xnor U14714 (N_14714,N_14251,N_14429);
nor U14715 (N_14715,N_14472,N_14196);
and U14716 (N_14716,N_14252,N_14199);
xor U14717 (N_14717,N_14133,N_14172);
nor U14718 (N_14718,N_14499,N_14083);
or U14719 (N_14719,N_14079,N_14220);
xor U14720 (N_14720,N_14059,N_14406);
nand U14721 (N_14721,N_14365,N_14214);
nand U14722 (N_14722,N_14352,N_14306);
xor U14723 (N_14723,N_14422,N_14440);
xnor U14724 (N_14724,N_14442,N_14004);
and U14725 (N_14725,N_14475,N_14190);
nor U14726 (N_14726,N_14145,N_14219);
xor U14727 (N_14727,N_14253,N_14434);
nor U14728 (N_14728,N_14450,N_14370);
nor U14729 (N_14729,N_14298,N_14029);
nand U14730 (N_14730,N_14140,N_14284);
and U14731 (N_14731,N_14211,N_14117);
nor U14732 (N_14732,N_14456,N_14037);
and U14733 (N_14733,N_14200,N_14272);
or U14734 (N_14734,N_14147,N_14308);
nand U14735 (N_14735,N_14271,N_14392);
and U14736 (N_14736,N_14375,N_14157);
or U14737 (N_14737,N_14022,N_14328);
nand U14738 (N_14738,N_14012,N_14102);
xnor U14739 (N_14739,N_14483,N_14263);
and U14740 (N_14740,N_14212,N_14401);
nor U14741 (N_14741,N_14324,N_14000);
nand U14742 (N_14742,N_14056,N_14042);
and U14743 (N_14743,N_14473,N_14382);
or U14744 (N_14744,N_14323,N_14439);
or U14745 (N_14745,N_14119,N_14385);
xor U14746 (N_14746,N_14186,N_14318);
nor U14747 (N_14747,N_14030,N_14159);
or U14748 (N_14748,N_14202,N_14218);
or U14749 (N_14749,N_14354,N_14276);
nand U14750 (N_14750,N_14332,N_14252);
or U14751 (N_14751,N_14369,N_14444);
or U14752 (N_14752,N_14286,N_14472);
or U14753 (N_14753,N_14272,N_14001);
xor U14754 (N_14754,N_14243,N_14491);
nand U14755 (N_14755,N_14161,N_14242);
and U14756 (N_14756,N_14194,N_14368);
nor U14757 (N_14757,N_14114,N_14013);
or U14758 (N_14758,N_14304,N_14135);
or U14759 (N_14759,N_14324,N_14250);
or U14760 (N_14760,N_14222,N_14068);
nand U14761 (N_14761,N_14188,N_14375);
nand U14762 (N_14762,N_14218,N_14252);
nand U14763 (N_14763,N_14202,N_14207);
or U14764 (N_14764,N_14303,N_14317);
nand U14765 (N_14765,N_14205,N_14327);
nor U14766 (N_14766,N_14261,N_14320);
or U14767 (N_14767,N_14205,N_14385);
xnor U14768 (N_14768,N_14174,N_14466);
or U14769 (N_14769,N_14094,N_14361);
xnor U14770 (N_14770,N_14064,N_14027);
nand U14771 (N_14771,N_14279,N_14398);
nand U14772 (N_14772,N_14428,N_14300);
nor U14773 (N_14773,N_14378,N_14168);
or U14774 (N_14774,N_14353,N_14358);
nor U14775 (N_14775,N_14096,N_14097);
and U14776 (N_14776,N_14260,N_14429);
or U14777 (N_14777,N_14457,N_14079);
or U14778 (N_14778,N_14067,N_14346);
nor U14779 (N_14779,N_14472,N_14138);
nor U14780 (N_14780,N_14477,N_14043);
nand U14781 (N_14781,N_14377,N_14222);
nand U14782 (N_14782,N_14493,N_14084);
and U14783 (N_14783,N_14474,N_14108);
or U14784 (N_14784,N_14006,N_14137);
or U14785 (N_14785,N_14094,N_14090);
xnor U14786 (N_14786,N_14288,N_14374);
nand U14787 (N_14787,N_14215,N_14416);
xor U14788 (N_14788,N_14410,N_14179);
xor U14789 (N_14789,N_14107,N_14457);
xnor U14790 (N_14790,N_14365,N_14490);
or U14791 (N_14791,N_14019,N_14309);
nor U14792 (N_14792,N_14126,N_14118);
nor U14793 (N_14793,N_14254,N_14130);
nand U14794 (N_14794,N_14277,N_14393);
nand U14795 (N_14795,N_14074,N_14168);
nor U14796 (N_14796,N_14396,N_14044);
nor U14797 (N_14797,N_14355,N_14364);
xnor U14798 (N_14798,N_14124,N_14371);
and U14799 (N_14799,N_14106,N_14235);
or U14800 (N_14800,N_14172,N_14194);
nand U14801 (N_14801,N_14078,N_14115);
and U14802 (N_14802,N_14455,N_14370);
nor U14803 (N_14803,N_14398,N_14499);
xnor U14804 (N_14804,N_14428,N_14285);
nand U14805 (N_14805,N_14413,N_14298);
nand U14806 (N_14806,N_14396,N_14182);
nand U14807 (N_14807,N_14262,N_14052);
and U14808 (N_14808,N_14021,N_14142);
xor U14809 (N_14809,N_14118,N_14323);
or U14810 (N_14810,N_14413,N_14310);
xor U14811 (N_14811,N_14189,N_14382);
and U14812 (N_14812,N_14191,N_14436);
or U14813 (N_14813,N_14306,N_14176);
nor U14814 (N_14814,N_14105,N_14431);
nand U14815 (N_14815,N_14386,N_14391);
xnor U14816 (N_14816,N_14369,N_14084);
or U14817 (N_14817,N_14028,N_14414);
and U14818 (N_14818,N_14369,N_14308);
nor U14819 (N_14819,N_14097,N_14121);
xor U14820 (N_14820,N_14031,N_14431);
xor U14821 (N_14821,N_14113,N_14042);
nand U14822 (N_14822,N_14424,N_14161);
or U14823 (N_14823,N_14492,N_14412);
nand U14824 (N_14824,N_14176,N_14036);
nand U14825 (N_14825,N_14009,N_14432);
nand U14826 (N_14826,N_14320,N_14116);
xor U14827 (N_14827,N_14001,N_14484);
and U14828 (N_14828,N_14220,N_14407);
nor U14829 (N_14829,N_14098,N_14047);
xor U14830 (N_14830,N_14068,N_14326);
xor U14831 (N_14831,N_14105,N_14044);
or U14832 (N_14832,N_14394,N_14282);
nand U14833 (N_14833,N_14037,N_14245);
nor U14834 (N_14834,N_14104,N_14183);
and U14835 (N_14835,N_14069,N_14162);
xnor U14836 (N_14836,N_14037,N_14062);
xor U14837 (N_14837,N_14151,N_14232);
nand U14838 (N_14838,N_14442,N_14365);
and U14839 (N_14839,N_14094,N_14050);
or U14840 (N_14840,N_14101,N_14265);
or U14841 (N_14841,N_14191,N_14295);
and U14842 (N_14842,N_14182,N_14059);
nand U14843 (N_14843,N_14375,N_14096);
or U14844 (N_14844,N_14497,N_14127);
nor U14845 (N_14845,N_14333,N_14006);
and U14846 (N_14846,N_14381,N_14408);
nor U14847 (N_14847,N_14038,N_14495);
and U14848 (N_14848,N_14139,N_14341);
nor U14849 (N_14849,N_14178,N_14296);
xnor U14850 (N_14850,N_14263,N_14402);
nand U14851 (N_14851,N_14222,N_14103);
nand U14852 (N_14852,N_14041,N_14384);
xnor U14853 (N_14853,N_14303,N_14392);
xnor U14854 (N_14854,N_14482,N_14274);
nor U14855 (N_14855,N_14474,N_14264);
or U14856 (N_14856,N_14147,N_14437);
and U14857 (N_14857,N_14221,N_14463);
and U14858 (N_14858,N_14483,N_14073);
nor U14859 (N_14859,N_14458,N_14099);
nor U14860 (N_14860,N_14452,N_14354);
and U14861 (N_14861,N_14160,N_14157);
xor U14862 (N_14862,N_14316,N_14047);
and U14863 (N_14863,N_14251,N_14490);
nor U14864 (N_14864,N_14109,N_14036);
and U14865 (N_14865,N_14440,N_14093);
and U14866 (N_14866,N_14007,N_14289);
or U14867 (N_14867,N_14059,N_14437);
or U14868 (N_14868,N_14428,N_14487);
nand U14869 (N_14869,N_14050,N_14035);
nor U14870 (N_14870,N_14245,N_14341);
or U14871 (N_14871,N_14469,N_14413);
nor U14872 (N_14872,N_14377,N_14411);
nor U14873 (N_14873,N_14201,N_14435);
or U14874 (N_14874,N_14160,N_14009);
or U14875 (N_14875,N_14329,N_14415);
xor U14876 (N_14876,N_14117,N_14082);
nor U14877 (N_14877,N_14461,N_14175);
nor U14878 (N_14878,N_14391,N_14419);
and U14879 (N_14879,N_14356,N_14108);
and U14880 (N_14880,N_14045,N_14031);
xor U14881 (N_14881,N_14140,N_14275);
nor U14882 (N_14882,N_14457,N_14142);
xnor U14883 (N_14883,N_14143,N_14182);
xor U14884 (N_14884,N_14250,N_14214);
nor U14885 (N_14885,N_14244,N_14484);
nor U14886 (N_14886,N_14353,N_14153);
xnor U14887 (N_14887,N_14249,N_14350);
nor U14888 (N_14888,N_14457,N_14012);
nand U14889 (N_14889,N_14421,N_14457);
xor U14890 (N_14890,N_14408,N_14373);
or U14891 (N_14891,N_14386,N_14485);
nor U14892 (N_14892,N_14253,N_14467);
xor U14893 (N_14893,N_14384,N_14482);
nand U14894 (N_14894,N_14052,N_14423);
xnor U14895 (N_14895,N_14233,N_14070);
nand U14896 (N_14896,N_14302,N_14135);
nor U14897 (N_14897,N_14151,N_14463);
or U14898 (N_14898,N_14233,N_14354);
xor U14899 (N_14899,N_14184,N_14095);
xor U14900 (N_14900,N_14190,N_14411);
nand U14901 (N_14901,N_14371,N_14010);
or U14902 (N_14902,N_14293,N_14345);
nand U14903 (N_14903,N_14272,N_14183);
and U14904 (N_14904,N_14230,N_14388);
and U14905 (N_14905,N_14116,N_14477);
xnor U14906 (N_14906,N_14070,N_14292);
nand U14907 (N_14907,N_14358,N_14090);
nor U14908 (N_14908,N_14120,N_14060);
nand U14909 (N_14909,N_14383,N_14194);
or U14910 (N_14910,N_14379,N_14491);
nor U14911 (N_14911,N_14138,N_14234);
nand U14912 (N_14912,N_14193,N_14225);
nand U14913 (N_14913,N_14311,N_14241);
nand U14914 (N_14914,N_14278,N_14302);
and U14915 (N_14915,N_14301,N_14212);
xnor U14916 (N_14916,N_14286,N_14359);
xnor U14917 (N_14917,N_14279,N_14240);
or U14918 (N_14918,N_14312,N_14076);
and U14919 (N_14919,N_14437,N_14475);
and U14920 (N_14920,N_14097,N_14091);
nand U14921 (N_14921,N_14413,N_14458);
or U14922 (N_14922,N_14322,N_14223);
xor U14923 (N_14923,N_14381,N_14009);
or U14924 (N_14924,N_14230,N_14411);
xnor U14925 (N_14925,N_14176,N_14396);
or U14926 (N_14926,N_14244,N_14149);
xor U14927 (N_14927,N_14178,N_14096);
or U14928 (N_14928,N_14016,N_14467);
and U14929 (N_14929,N_14142,N_14235);
nor U14930 (N_14930,N_14043,N_14327);
or U14931 (N_14931,N_14348,N_14488);
nand U14932 (N_14932,N_14470,N_14458);
or U14933 (N_14933,N_14383,N_14360);
nor U14934 (N_14934,N_14411,N_14339);
and U14935 (N_14935,N_14496,N_14305);
nand U14936 (N_14936,N_14036,N_14019);
nand U14937 (N_14937,N_14090,N_14397);
and U14938 (N_14938,N_14170,N_14021);
nor U14939 (N_14939,N_14010,N_14448);
and U14940 (N_14940,N_14190,N_14162);
xor U14941 (N_14941,N_14152,N_14093);
nor U14942 (N_14942,N_14085,N_14238);
and U14943 (N_14943,N_14171,N_14422);
xor U14944 (N_14944,N_14268,N_14075);
nand U14945 (N_14945,N_14367,N_14005);
and U14946 (N_14946,N_14002,N_14347);
nor U14947 (N_14947,N_14203,N_14446);
nor U14948 (N_14948,N_14133,N_14333);
or U14949 (N_14949,N_14440,N_14185);
or U14950 (N_14950,N_14432,N_14395);
or U14951 (N_14951,N_14011,N_14217);
nand U14952 (N_14952,N_14426,N_14113);
or U14953 (N_14953,N_14232,N_14225);
nor U14954 (N_14954,N_14123,N_14371);
nor U14955 (N_14955,N_14188,N_14134);
xor U14956 (N_14956,N_14013,N_14153);
xor U14957 (N_14957,N_14255,N_14317);
nand U14958 (N_14958,N_14339,N_14367);
or U14959 (N_14959,N_14114,N_14229);
xnor U14960 (N_14960,N_14089,N_14495);
and U14961 (N_14961,N_14058,N_14187);
and U14962 (N_14962,N_14406,N_14085);
xor U14963 (N_14963,N_14110,N_14187);
nand U14964 (N_14964,N_14410,N_14371);
nor U14965 (N_14965,N_14309,N_14310);
and U14966 (N_14966,N_14335,N_14490);
nor U14967 (N_14967,N_14228,N_14251);
xnor U14968 (N_14968,N_14281,N_14393);
nand U14969 (N_14969,N_14089,N_14160);
nor U14970 (N_14970,N_14245,N_14281);
nand U14971 (N_14971,N_14376,N_14006);
nand U14972 (N_14972,N_14224,N_14399);
nor U14973 (N_14973,N_14317,N_14314);
nand U14974 (N_14974,N_14499,N_14466);
and U14975 (N_14975,N_14418,N_14066);
nor U14976 (N_14976,N_14412,N_14418);
or U14977 (N_14977,N_14016,N_14100);
nor U14978 (N_14978,N_14311,N_14124);
nand U14979 (N_14979,N_14138,N_14273);
nor U14980 (N_14980,N_14327,N_14148);
nor U14981 (N_14981,N_14382,N_14078);
and U14982 (N_14982,N_14269,N_14439);
xnor U14983 (N_14983,N_14437,N_14461);
or U14984 (N_14984,N_14030,N_14467);
and U14985 (N_14985,N_14179,N_14215);
xnor U14986 (N_14986,N_14220,N_14049);
nand U14987 (N_14987,N_14075,N_14066);
or U14988 (N_14988,N_14336,N_14485);
or U14989 (N_14989,N_14023,N_14104);
xor U14990 (N_14990,N_14019,N_14482);
xnor U14991 (N_14991,N_14112,N_14488);
xnor U14992 (N_14992,N_14378,N_14494);
nand U14993 (N_14993,N_14259,N_14375);
nor U14994 (N_14994,N_14469,N_14412);
or U14995 (N_14995,N_14443,N_14131);
nor U14996 (N_14996,N_14272,N_14355);
nand U14997 (N_14997,N_14131,N_14299);
xor U14998 (N_14998,N_14181,N_14092);
xnor U14999 (N_14999,N_14083,N_14447);
xor UO_0 (O_0,N_14516,N_14946);
nor UO_1 (O_1,N_14553,N_14791);
nand UO_2 (O_2,N_14619,N_14644);
xnor UO_3 (O_3,N_14608,N_14874);
xnor UO_4 (O_4,N_14637,N_14808);
nor UO_5 (O_5,N_14835,N_14910);
or UO_6 (O_6,N_14670,N_14728);
or UO_7 (O_7,N_14536,N_14783);
and UO_8 (O_8,N_14793,N_14603);
or UO_9 (O_9,N_14813,N_14676);
or UO_10 (O_10,N_14502,N_14734);
nor UO_11 (O_11,N_14661,N_14565);
nor UO_12 (O_12,N_14664,N_14669);
and UO_13 (O_13,N_14591,N_14842);
xnor UO_14 (O_14,N_14948,N_14710);
or UO_15 (O_15,N_14537,N_14753);
or UO_16 (O_16,N_14709,N_14823);
xor UO_17 (O_17,N_14902,N_14802);
or UO_18 (O_18,N_14564,N_14784);
xnor UO_19 (O_19,N_14843,N_14764);
nand UO_20 (O_20,N_14872,N_14566);
and UO_21 (O_21,N_14555,N_14697);
or UO_22 (O_22,N_14828,N_14759);
nor UO_23 (O_23,N_14920,N_14853);
and UO_24 (O_24,N_14888,N_14520);
and UO_25 (O_25,N_14579,N_14716);
and UO_26 (O_26,N_14668,N_14826);
nand UO_27 (O_27,N_14798,N_14901);
xnor UO_28 (O_28,N_14940,N_14900);
nor UO_29 (O_29,N_14860,N_14976);
xnor UO_30 (O_30,N_14679,N_14846);
or UO_31 (O_31,N_14725,N_14702);
nand UO_32 (O_32,N_14634,N_14720);
xor UO_33 (O_33,N_14756,N_14656);
xnor UO_34 (O_34,N_14944,N_14941);
and UO_35 (O_35,N_14815,N_14622);
and UO_36 (O_36,N_14769,N_14677);
xor UO_37 (O_37,N_14501,N_14873);
nor UO_38 (O_38,N_14703,N_14535);
and UO_39 (O_39,N_14856,N_14523);
nor UO_40 (O_40,N_14780,N_14561);
or UO_41 (O_41,N_14961,N_14951);
or UO_42 (O_42,N_14527,N_14792);
and UO_43 (O_43,N_14594,N_14840);
and UO_44 (O_44,N_14859,N_14788);
or UO_45 (O_45,N_14576,N_14581);
or UO_46 (O_46,N_14991,N_14767);
nand UO_47 (O_47,N_14949,N_14999);
and UO_48 (O_48,N_14636,N_14510);
or UO_49 (O_49,N_14772,N_14683);
xnor UO_50 (O_50,N_14867,N_14863);
nand UO_51 (O_51,N_14893,N_14947);
and UO_52 (O_52,N_14519,N_14580);
nand UO_53 (O_53,N_14542,N_14620);
and UO_54 (O_54,N_14665,N_14886);
nand UO_55 (O_55,N_14639,N_14795);
nand UO_56 (O_56,N_14800,N_14938);
and UO_57 (O_57,N_14586,N_14575);
nor UO_58 (O_58,N_14610,N_14653);
and UO_59 (O_59,N_14507,N_14917);
xor UO_60 (O_60,N_14629,N_14824);
or UO_61 (O_61,N_14916,N_14547);
xor UO_62 (O_62,N_14680,N_14939);
xor UO_63 (O_63,N_14745,N_14628);
nand UO_64 (O_64,N_14545,N_14965);
nand UO_65 (O_65,N_14666,N_14834);
nand UO_66 (O_66,N_14662,N_14650);
nand UO_67 (O_67,N_14692,N_14771);
nand UO_68 (O_68,N_14922,N_14848);
xor UO_69 (O_69,N_14736,N_14587);
nor UO_70 (O_70,N_14647,N_14562);
nand UO_71 (O_71,N_14616,N_14701);
nor UO_72 (O_72,N_14735,N_14930);
and UO_73 (O_73,N_14796,N_14718);
or UO_74 (O_74,N_14573,N_14583);
and UO_75 (O_75,N_14560,N_14659);
nor UO_76 (O_76,N_14538,N_14567);
nor UO_77 (O_77,N_14915,N_14526);
nor UO_78 (O_78,N_14623,N_14990);
xor UO_79 (O_79,N_14958,N_14604);
and UO_80 (O_80,N_14731,N_14690);
nand UO_81 (O_81,N_14773,N_14762);
nor UO_82 (O_82,N_14751,N_14599);
and UO_83 (O_83,N_14621,N_14631);
xnor UO_84 (O_84,N_14673,N_14998);
and UO_85 (O_85,N_14511,N_14512);
nor UO_86 (O_86,N_14973,N_14651);
nor UO_87 (O_87,N_14908,N_14919);
nor UO_88 (O_88,N_14598,N_14812);
nand UO_89 (O_89,N_14833,N_14879);
or UO_90 (O_90,N_14667,N_14758);
xor UO_91 (O_91,N_14504,N_14768);
nor UO_92 (O_92,N_14766,N_14881);
nor UO_93 (O_93,N_14674,N_14882);
and UO_94 (O_94,N_14984,N_14626);
or UO_95 (O_95,N_14831,N_14929);
nand UO_96 (O_96,N_14817,N_14509);
xnor UO_97 (O_97,N_14832,N_14937);
or UO_98 (O_98,N_14844,N_14557);
and UO_99 (O_99,N_14752,N_14717);
or UO_100 (O_100,N_14827,N_14957);
and UO_101 (O_101,N_14614,N_14524);
nor UO_102 (O_102,N_14529,N_14993);
nand UO_103 (O_103,N_14500,N_14956);
nand UO_104 (O_104,N_14801,N_14714);
and UO_105 (O_105,N_14570,N_14657);
or UO_106 (O_106,N_14803,N_14777);
or UO_107 (O_107,N_14612,N_14508);
and UO_108 (O_108,N_14592,N_14695);
xnor UO_109 (O_109,N_14986,N_14926);
nor UO_110 (O_110,N_14595,N_14515);
and UO_111 (O_111,N_14954,N_14968);
or UO_112 (O_112,N_14606,N_14630);
xnor UO_113 (O_113,N_14871,N_14906);
and UO_114 (O_114,N_14715,N_14593);
or UO_115 (O_115,N_14822,N_14774);
or UO_116 (O_116,N_14989,N_14923);
nand UO_117 (O_117,N_14607,N_14678);
or UO_118 (O_118,N_14672,N_14855);
and UO_119 (O_119,N_14837,N_14521);
nand UO_120 (O_120,N_14503,N_14540);
xor UO_121 (O_121,N_14980,N_14531);
nor UO_122 (O_122,N_14569,N_14546);
and UO_123 (O_123,N_14596,N_14691);
nand UO_124 (O_124,N_14530,N_14790);
nor UO_125 (O_125,N_14825,N_14857);
xor UO_126 (O_126,N_14789,N_14649);
nor UO_127 (O_127,N_14559,N_14694);
nand UO_128 (O_128,N_14601,N_14689);
or UO_129 (O_129,N_14525,N_14894);
nand UO_130 (O_130,N_14979,N_14847);
nand UO_131 (O_131,N_14663,N_14799);
nand UO_132 (O_132,N_14638,N_14988);
or UO_133 (O_133,N_14876,N_14810);
and UO_134 (O_134,N_14642,N_14539);
xnor UO_135 (O_135,N_14605,N_14912);
nand UO_136 (O_136,N_14839,N_14870);
or UO_137 (O_137,N_14978,N_14633);
nor UO_138 (O_138,N_14982,N_14829);
xor UO_139 (O_139,N_14787,N_14821);
nor UO_140 (O_140,N_14913,N_14811);
or UO_141 (O_141,N_14806,N_14786);
and UO_142 (O_142,N_14757,N_14571);
and UO_143 (O_143,N_14804,N_14942);
nand UO_144 (O_144,N_14641,N_14970);
nand UO_145 (O_145,N_14548,N_14866);
nor UO_146 (O_146,N_14646,N_14719);
xnor UO_147 (O_147,N_14864,N_14685);
nor UO_148 (O_148,N_14987,N_14609);
and UO_149 (O_149,N_14549,N_14841);
nor UO_150 (O_150,N_14578,N_14820);
xor UO_151 (O_151,N_14985,N_14883);
nand UO_152 (O_152,N_14624,N_14574);
or UO_153 (O_153,N_14921,N_14618);
or UO_154 (O_154,N_14708,N_14517);
nor UO_155 (O_155,N_14933,N_14747);
and UO_156 (O_156,N_14577,N_14700);
nor UO_157 (O_157,N_14895,N_14640);
or UO_158 (O_158,N_14729,N_14738);
and UO_159 (O_159,N_14746,N_14966);
nor UO_160 (O_160,N_14918,N_14754);
xor UO_161 (O_161,N_14972,N_14563);
or UO_162 (O_162,N_14730,N_14849);
or UO_163 (O_163,N_14974,N_14643);
xnor UO_164 (O_164,N_14588,N_14617);
xor UO_165 (O_165,N_14721,N_14625);
nand UO_166 (O_166,N_14816,N_14878);
xor UO_167 (O_167,N_14967,N_14655);
and UO_168 (O_168,N_14892,N_14505);
nand UO_169 (O_169,N_14550,N_14977);
or UO_170 (O_170,N_14869,N_14955);
or UO_171 (O_171,N_14532,N_14924);
nor UO_172 (O_172,N_14654,N_14763);
nand UO_173 (O_173,N_14931,N_14749);
xor UO_174 (O_174,N_14541,N_14627);
xnor UO_175 (O_175,N_14794,N_14890);
and UO_176 (O_176,N_14880,N_14785);
xor UO_177 (O_177,N_14934,N_14877);
nor UO_178 (O_178,N_14885,N_14687);
nand UO_179 (O_179,N_14558,N_14506);
and UO_180 (O_180,N_14652,N_14554);
or UO_181 (O_181,N_14852,N_14632);
nor UO_182 (O_182,N_14684,N_14600);
xnor UO_183 (O_183,N_14740,N_14962);
nor UO_184 (O_184,N_14838,N_14782);
and UO_185 (O_185,N_14914,N_14865);
nor UO_186 (O_186,N_14907,N_14675);
or UO_187 (O_187,N_14741,N_14615);
and UO_188 (O_188,N_14971,N_14928);
nor UO_189 (O_189,N_14611,N_14693);
nand UO_190 (O_190,N_14585,N_14727);
nand UO_191 (O_191,N_14845,N_14645);
nor UO_192 (O_192,N_14613,N_14770);
nor UO_193 (O_193,N_14994,N_14743);
nor UO_194 (O_194,N_14889,N_14705);
and UO_195 (O_195,N_14713,N_14897);
xor UO_196 (O_196,N_14543,N_14868);
and UO_197 (O_197,N_14589,N_14699);
xor UO_198 (O_198,N_14862,N_14704);
and UO_199 (O_199,N_14513,N_14556);
and UO_200 (O_200,N_14776,N_14836);
or UO_201 (O_201,N_14723,N_14797);
or UO_202 (O_202,N_14744,N_14760);
or UO_203 (O_203,N_14602,N_14935);
nand UO_204 (O_204,N_14875,N_14775);
and UO_205 (O_205,N_14551,N_14960);
or UO_206 (O_206,N_14778,N_14712);
nor UO_207 (O_207,N_14528,N_14706);
nor UO_208 (O_208,N_14995,N_14732);
nand UO_209 (O_209,N_14953,N_14861);
nand UO_210 (O_210,N_14997,N_14805);
and UO_211 (O_211,N_14686,N_14854);
nor UO_212 (O_212,N_14514,N_14896);
nand UO_213 (O_213,N_14830,N_14903);
nor UO_214 (O_214,N_14681,N_14711);
or UO_215 (O_215,N_14818,N_14945);
nor UO_216 (O_216,N_14522,N_14905);
and UO_217 (O_217,N_14544,N_14809);
nor UO_218 (O_218,N_14858,N_14750);
or UO_219 (O_219,N_14964,N_14737);
nand UO_220 (O_220,N_14884,N_14891);
or UO_221 (O_221,N_14733,N_14996);
nor UO_222 (O_222,N_14696,N_14887);
or UO_223 (O_223,N_14726,N_14688);
or UO_224 (O_224,N_14814,N_14648);
nand UO_225 (O_225,N_14936,N_14597);
nor UO_226 (O_226,N_14742,N_14911);
and UO_227 (O_227,N_14698,N_14552);
xor UO_228 (O_228,N_14850,N_14682);
and UO_229 (O_229,N_14952,N_14534);
nor UO_230 (O_230,N_14739,N_14671);
or UO_231 (O_231,N_14983,N_14755);
xor UO_232 (O_232,N_14572,N_14568);
or UO_233 (O_233,N_14975,N_14707);
nand UO_234 (O_234,N_14635,N_14781);
or UO_235 (O_235,N_14533,N_14899);
nand UO_236 (O_236,N_14584,N_14851);
or UO_237 (O_237,N_14590,N_14658);
or UO_238 (O_238,N_14722,N_14969);
and UO_239 (O_239,N_14909,N_14779);
nor UO_240 (O_240,N_14959,N_14761);
or UO_241 (O_241,N_14819,N_14963);
nand UO_242 (O_242,N_14748,N_14898);
or UO_243 (O_243,N_14807,N_14992);
or UO_244 (O_244,N_14724,N_14518);
nor UO_245 (O_245,N_14932,N_14660);
or UO_246 (O_246,N_14943,N_14582);
nand UO_247 (O_247,N_14927,N_14925);
and UO_248 (O_248,N_14981,N_14765);
xnor UO_249 (O_249,N_14950,N_14904);
nand UO_250 (O_250,N_14961,N_14928);
nor UO_251 (O_251,N_14956,N_14755);
xnor UO_252 (O_252,N_14693,N_14976);
or UO_253 (O_253,N_14698,N_14847);
and UO_254 (O_254,N_14733,N_14823);
nand UO_255 (O_255,N_14579,N_14975);
xnor UO_256 (O_256,N_14614,N_14801);
nand UO_257 (O_257,N_14683,N_14671);
or UO_258 (O_258,N_14715,N_14533);
xor UO_259 (O_259,N_14980,N_14969);
nor UO_260 (O_260,N_14930,N_14879);
and UO_261 (O_261,N_14573,N_14723);
and UO_262 (O_262,N_14602,N_14904);
and UO_263 (O_263,N_14577,N_14760);
or UO_264 (O_264,N_14874,N_14585);
and UO_265 (O_265,N_14990,N_14631);
nor UO_266 (O_266,N_14795,N_14806);
nor UO_267 (O_267,N_14815,N_14706);
nor UO_268 (O_268,N_14587,N_14536);
nand UO_269 (O_269,N_14705,N_14734);
or UO_270 (O_270,N_14988,N_14932);
and UO_271 (O_271,N_14946,N_14873);
xor UO_272 (O_272,N_14869,N_14542);
nand UO_273 (O_273,N_14652,N_14787);
nand UO_274 (O_274,N_14769,N_14876);
and UO_275 (O_275,N_14519,N_14690);
nand UO_276 (O_276,N_14664,N_14705);
nor UO_277 (O_277,N_14712,N_14807);
nand UO_278 (O_278,N_14705,N_14761);
and UO_279 (O_279,N_14560,N_14957);
nor UO_280 (O_280,N_14716,N_14793);
and UO_281 (O_281,N_14927,N_14787);
or UO_282 (O_282,N_14898,N_14633);
xnor UO_283 (O_283,N_14684,N_14669);
nand UO_284 (O_284,N_14869,N_14547);
or UO_285 (O_285,N_14925,N_14805);
nand UO_286 (O_286,N_14780,N_14736);
nor UO_287 (O_287,N_14728,N_14797);
nor UO_288 (O_288,N_14715,N_14560);
nand UO_289 (O_289,N_14898,N_14774);
nor UO_290 (O_290,N_14735,N_14664);
nor UO_291 (O_291,N_14945,N_14930);
nand UO_292 (O_292,N_14836,N_14536);
nand UO_293 (O_293,N_14602,N_14541);
and UO_294 (O_294,N_14700,N_14717);
and UO_295 (O_295,N_14635,N_14810);
and UO_296 (O_296,N_14565,N_14961);
xnor UO_297 (O_297,N_14964,N_14992);
or UO_298 (O_298,N_14770,N_14749);
xnor UO_299 (O_299,N_14653,N_14545);
and UO_300 (O_300,N_14951,N_14623);
nor UO_301 (O_301,N_14771,N_14826);
nand UO_302 (O_302,N_14709,N_14860);
nor UO_303 (O_303,N_14961,N_14661);
or UO_304 (O_304,N_14525,N_14731);
nand UO_305 (O_305,N_14580,N_14656);
xnor UO_306 (O_306,N_14884,N_14829);
or UO_307 (O_307,N_14581,N_14998);
or UO_308 (O_308,N_14746,N_14650);
nor UO_309 (O_309,N_14733,N_14545);
nand UO_310 (O_310,N_14975,N_14967);
and UO_311 (O_311,N_14754,N_14550);
or UO_312 (O_312,N_14691,N_14747);
xnor UO_313 (O_313,N_14895,N_14972);
nand UO_314 (O_314,N_14702,N_14709);
nand UO_315 (O_315,N_14977,N_14731);
nand UO_316 (O_316,N_14831,N_14738);
xnor UO_317 (O_317,N_14617,N_14576);
nand UO_318 (O_318,N_14791,N_14870);
xor UO_319 (O_319,N_14851,N_14936);
xnor UO_320 (O_320,N_14972,N_14835);
xnor UO_321 (O_321,N_14510,N_14892);
nand UO_322 (O_322,N_14815,N_14896);
or UO_323 (O_323,N_14794,N_14881);
or UO_324 (O_324,N_14744,N_14831);
nor UO_325 (O_325,N_14585,N_14594);
and UO_326 (O_326,N_14896,N_14989);
or UO_327 (O_327,N_14625,N_14910);
and UO_328 (O_328,N_14723,N_14914);
or UO_329 (O_329,N_14550,N_14865);
or UO_330 (O_330,N_14899,N_14690);
and UO_331 (O_331,N_14890,N_14866);
xnor UO_332 (O_332,N_14573,N_14504);
xnor UO_333 (O_333,N_14943,N_14665);
or UO_334 (O_334,N_14810,N_14714);
and UO_335 (O_335,N_14844,N_14595);
and UO_336 (O_336,N_14942,N_14802);
and UO_337 (O_337,N_14796,N_14783);
nor UO_338 (O_338,N_14563,N_14515);
or UO_339 (O_339,N_14920,N_14842);
or UO_340 (O_340,N_14587,N_14778);
nand UO_341 (O_341,N_14932,N_14714);
or UO_342 (O_342,N_14557,N_14878);
nor UO_343 (O_343,N_14525,N_14877);
and UO_344 (O_344,N_14654,N_14865);
xor UO_345 (O_345,N_14969,N_14686);
nor UO_346 (O_346,N_14520,N_14558);
and UO_347 (O_347,N_14512,N_14953);
xnor UO_348 (O_348,N_14503,N_14707);
nor UO_349 (O_349,N_14566,N_14810);
nand UO_350 (O_350,N_14706,N_14553);
nor UO_351 (O_351,N_14631,N_14921);
or UO_352 (O_352,N_14663,N_14569);
and UO_353 (O_353,N_14546,N_14691);
or UO_354 (O_354,N_14576,N_14695);
and UO_355 (O_355,N_14750,N_14719);
and UO_356 (O_356,N_14808,N_14593);
or UO_357 (O_357,N_14991,N_14911);
nand UO_358 (O_358,N_14659,N_14924);
or UO_359 (O_359,N_14814,N_14902);
xor UO_360 (O_360,N_14575,N_14755);
xnor UO_361 (O_361,N_14547,N_14991);
xor UO_362 (O_362,N_14906,N_14888);
or UO_363 (O_363,N_14670,N_14986);
or UO_364 (O_364,N_14749,N_14630);
nor UO_365 (O_365,N_14918,N_14648);
xor UO_366 (O_366,N_14520,N_14966);
and UO_367 (O_367,N_14597,N_14785);
nor UO_368 (O_368,N_14633,N_14680);
and UO_369 (O_369,N_14892,N_14986);
nor UO_370 (O_370,N_14694,N_14638);
and UO_371 (O_371,N_14701,N_14653);
and UO_372 (O_372,N_14647,N_14758);
nand UO_373 (O_373,N_14898,N_14836);
and UO_374 (O_374,N_14662,N_14786);
or UO_375 (O_375,N_14662,N_14522);
or UO_376 (O_376,N_14989,N_14987);
and UO_377 (O_377,N_14665,N_14733);
nand UO_378 (O_378,N_14777,N_14812);
nor UO_379 (O_379,N_14667,N_14827);
and UO_380 (O_380,N_14799,N_14542);
and UO_381 (O_381,N_14718,N_14988);
and UO_382 (O_382,N_14891,N_14648);
and UO_383 (O_383,N_14859,N_14797);
nand UO_384 (O_384,N_14646,N_14602);
xor UO_385 (O_385,N_14871,N_14720);
nand UO_386 (O_386,N_14814,N_14523);
xor UO_387 (O_387,N_14974,N_14757);
nand UO_388 (O_388,N_14503,N_14714);
nor UO_389 (O_389,N_14503,N_14818);
nand UO_390 (O_390,N_14713,N_14798);
nand UO_391 (O_391,N_14709,N_14508);
xnor UO_392 (O_392,N_14812,N_14865);
nand UO_393 (O_393,N_14743,N_14760);
nor UO_394 (O_394,N_14676,N_14994);
xor UO_395 (O_395,N_14971,N_14824);
nand UO_396 (O_396,N_14826,N_14598);
or UO_397 (O_397,N_14702,N_14569);
xor UO_398 (O_398,N_14828,N_14524);
nor UO_399 (O_399,N_14822,N_14844);
nor UO_400 (O_400,N_14532,N_14597);
nor UO_401 (O_401,N_14718,N_14768);
nor UO_402 (O_402,N_14828,N_14723);
nand UO_403 (O_403,N_14841,N_14832);
nand UO_404 (O_404,N_14695,N_14941);
nor UO_405 (O_405,N_14574,N_14889);
nand UO_406 (O_406,N_14865,N_14965);
xor UO_407 (O_407,N_14921,N_14600);
and UO_408 (O_408,N_14554,N_14896);
nand UO_409 (O_409,N_14963,N_14758);
nand UO_410 (O_410,N_14654,N_14737);
or UO_411 (O_411,N_14797,N_14891);
nand UO_412 (O_412,N_14956,N_14850);
or UO_413 (O_413,N_14677,N_14991);
or UO_414 (O_414,N_14530,N_14559);
or UO_415 (O_415,N_14544,N_14932);
nor UO_416 (O_416,N_14529,N_14744);
xor UO_417 (O_417,N_14818,N_14692);
nand UO_418 (O_418,N_14853,N_14997);
or UO_419 (O_419,N_14838,N_14980);
xor UO_420 (O_420,N_14625,N_14567);
nand UO_421 (O_421,N_14564,N_14641);
and UO_422 (O_422,N_14968,N_14918);
nor UO_423 (O_423,N_14627,N_14759);
xnor UO_424 (O_424,N_14923,N_14572);
nor UO_425 (O_425,N_14645,N_14578);
nor UO_426 (O_426,N_14949,N_14970);
or UO_427 (O_427,N_14787,N_14802);
or UO_428 (O_428,N_14974,N_14577);
nand UO_429 (O_429,N_14567,N_14812);
nor UO_430 (O_430,N_14792,N_14868);
or UO_431 (O_431,N_14888,N_14530);
nor UO_432 (O_432,N_14653,N_14546);
or UO_433 (O_433,N_14980,N_14699);
and UO_434 (O_434,N_14996,N_14566);
nand UO_435 (O_435,N_14589,N_14752);
nand UO_436 (O_436,N_14824,N_14789);
or UO_437 (O_437,N_14738,N_14887);
and UO_438 (O_438,N_14941,N_14629);
nand UO_439 (O_439,N_14885,N_14762);
nand UO_440 (O_440,N_14598,N_14514);
and UO_441 (O_441,N_14591,N_14631);
or UO_442 (O_442,N_14583,N_14910);
nand UO_443 (O_443,N_14670,N_14765);
nand UO_444 (O_444,N_14590,N_14906);
nand UO_445 (O_445,N_14525,N_14745);
xor UO_446 (O_446,N_14804,N_14653);
and UO_447 (O_447,N_14943,N_14815);
nand UO_448 (O_448,N_14512,N_14749);
and UO_449 (O_449,N_14709,N_14941);
or UO_450 (O_450,N_14587,N_14633);
xor UO_451 (O_451,N_14554,N_14918);
nor UO_452 (O_452,N_14985,N_14820);
xnor UO_453 (O_453,N_14563,N_14831);
xnor UO_454 (O_454,N_14996,N_14947);
nand UO_455 (O_455,N_14824,N_14963);
nor UO_456 (O_456,N_14845,N_14613);
and UO_457 (O_457,N_14955,N_14649);
xor UO_458 (O_458,N_14885,N_14683);
nor UO_459 (O_459,N_14500,N_14682);
xnor UO_460 (O_460,N_14876,N_14934);
or UO_461 (O_461,N_14824,N_14856);
xor UO_462 (O_462,N_14712,N_14797);
xnor UO_463 (O_463,N_14884,N_14703);
and UO_464 (O_464,N_14540,N_14898);
and UO_465 (O_465,N_14797,N_14771);
xor UO_466 (O_466,N_14912,N_14519);
nor UO_467 (O_467,N_14713,N_14631);
or UO_468 (O_468,N_14860,N_14883);
xor UO_469 (O_469,N_14566,N_14904);
or UO_470 (O_470,N_14853,N_14554);
and UO_471 (O_471,N_14964,N_14988);
nor UO_472 (O_472,N_14980,N_14953);
or UO_473 (O_473,N_14954,N_14839);
xor UO_474 (O_474,N_14808,N_14736);
or UO_475 (O_475,N_14985,N_14939);
nand UO_476 (O_476,N_14565,N_14536);
and UO_477 (O_477,N_14654,N_14764);
or UO_478 (O_478,N_14924,N_14815);
xor UO_479 (O_479,N_14549,N_14578);
nor UO_480 (O_480,N_14823,N_14573);
xor UO_481 (O_481,N_14611,N_14603);
or UO_482 (O_482,N_14554,N_14521);
nor UO_483 (O_483,N_14932,N_14526);
or UO_484 (O_484,N_14518,N_14627);
xnor UO_485 (O_485,N_14579,N_14629);
or UO_486 (O_486,N_14528,N_14897);
or UO_487 (O_487,N_14970,N_14785);
nor UO_488 (O_488,N_14692,N_14730);
nand UO_489 (O_489,N_14813,N_14547);
nand UO_490 (O_490,N_14650,N_14930);
or UO_491 (O_491,N_14628,N_14864);
nand UO_492 (O_492,N_14816,N_14896);
xor UO_493 (O_493,N_14826,N_14535);
nand UO_494 (O_494,N_14894,N_14857);
nor UO_495 (O_495,N_14753,N_14884);
nor UO_496 (O_496,N_14589,N_14714);
xnor UO_497 (O_497,N_14537,N_14573);
or UO_498 (O_498,N_14555,N_14752);
nor UO_499 (O_499,N_14851,N_14995);
nand UO_500 (O_500,N_14528,N_14978);
nand UO_501 (O_501,N_14679,N_14991);
nor UO_502 (O_502,N_14638,N_14939);
nor UO_503 (O_503,N_14865,N_14578);
nor UO_504 (O_504,N_14547,N_14864);
or UO_505 (O_505,N_14826,N_14707);
and UO_506 (O_506,N_14822,N_14635);
nor UO_507 (O_507,N_14689,N_14713);
nor UO_508 (O_508,N_14517,N_14579);
and UO_509 (O_509,N_14757,N_14833);
and UO_510 (O_510,N_14703,N_14983);
or UO_511 (O_511,N_14594,N_14986);
or UO_512 (O_512,N_14793,N_14942);
nor UO_513 (O_513,N_14994,N_14762);
or UO_514 (O_514,N_14695,N_14525);
and UO_515 (O_515,N_14977,N_14740);
nand UO_516 (O_516,N_14836,N_14514);
nand UO_517 (O_517,N_14878,N_14839);
and UO_518 (O_518,N_14790,N_14769);
or UO_519 (O_519,N_14750,N_14672);
and UO_520 (O_520,N_14774,N_14990);
or UO_521 (O_521,N_14988,N_14598);
nand UO_522 (O_522,N_14968,N_14543);
or UO_523 (O_523,N_14567,N_14617);
and UO_524 (O_524,N_14989,N_14677);
nor UO_525 (O_525,N_14520,N_14878);
nand UO_526 (O_526,N_14540,N_14565);
and UO_527 (O_527,N_14748,N_14845);
nand UO_528 (O_528,N_14979,N_14856);
xnor UO_529 (O_529,N_14776,N_14705);
or UO_530 (O_530,N_14570,N_14756);
or UO_531 (O_531,N_14673,N_14775);
xor UO_532 (O_532,N_14982,N_14955);
xnor UO_533 (O_533,N_14604,N_14808);
and UO_534 (O_534,N_14768,N_14759);
and UO_535 (O_535,N_14918,N_14774);
nor UO_536 (O_536,N_14826,N_14786);
or UO_537 (O_537,N_14663,N_14908);
nand UO_538 (O_538,N_14950,N_14670);
or UO_539 (O_539,N_14591,N_14688);
or UO_540 (O_540,N_14759,N_14788);
and UO_541 (O_541,N_14852,N_14888);
and UO_542 (O_542,N_14866,N_14785);
nand UO_543 (O_543,N_14712,N_14619);
and UO_544 (O_544,N_14866,N_14614);
xnor UO_545 (O_545,N_14775,N_14861);
or UO_546 (O_546,N_14521,N_14625);
nand UO_547 (O_547,N_14933,N_14590);
and UO_548 (O_548,N_14719,N_14668);
or UO_549 (O_549,N_14983,N_14782);
nor UO_550 (O_550,N_14656,N_14848);
nand UO_551 (O_551,N_14664,N_14926);
xnor UO_552 (O_552,N_14979,N_14993);
nor UO_553 (O_553,N_14744,N_14818);
xnor UO_554 (O_554,N_14561,N_14845);
nor UO_555 (O_555,N_14515,N_14576);
and UO_556 (O_556,N_14913,N_14604);
and UO_557 (O_557,N_14859,N_14834);
nor UO_558 (O_558,N_14590,N_14822);
nand UO_559 (O_559,N_14610,N_14531);
nand UO_560 (O_560,N_14968,N_14723);
and UO_561 (O_561,N_14733,N_14969);
nor UO_562 (O_562,N_14634,N_14903);
nor UO_563 (O_563,N_14660,N_14831);
and UO_564 (O_564,N_14981,N_14931);
and UO_565 (O_565,N_14800,N_14515);
or UO_566 (O_566,N_14888,N_14608);
xor UO_567 (O_567,N_14596,N_14687);
xor UO_568 (O_568,N_14528,N_14972);
nand UO_569 (O_569,N_14924,N_14675);
nand UO_570 (O_570,N_14929,N_14769);
xnor UO_571 (O_571,N_14872,N_14817);
nand UO_572 (O_572,N_14897,N_14866);
or UO_573 (O_573,N_14852,N_14686);
and UO_574 (O_574,N_14732,N_14665);
nor UO_575 (O_575,N_14971,N_14780);
or UO_576 (O_576,N_14628,N_14692);
and UO_577 (O_577,N_14769,N_14618);
or UO_578 (O_578,N_14788,N_14842);
nand UO_579 (O_579,N_14709,N_14624);
nand UO_580 (O_580,N_14838,N_14565);
xor UO_581 (O_581,N_14919,N_14644);
nand UO_582 (O_582,N_14714,N_14719);
xor UO_583 (O_583,N_14711,N_14835);
nand UO_584 (O_584,N_14848,N_14762);
nor UO_585 (O_585,N_14674,N_14850);
nor UO_586 (O_586,N_14974,N_14630);
xor UO_587 (O_587,N_14668,N_14709);
and UO_588 (O_588,N_14807,N_14740);
and UO_589 (O_589,N_14688,N_14516);
and UO_590 (O_590,N_14664,N_14850);
nand UO_591 (O_591,N_14614,N_14963);
or UO_592 (O_592,N_14532,N_14955);
or UO_593 (O_593,N_14710,N_14861);
xor UO_594 (O_594,N_14980,N_14826);
and UO_595 (O_595,N_14875,N_14683);
xor UO_596 (O_596,N_14965,N_14641);
xor UO_597 (O_597,N_14986,N_14814);
nor UO_598 (O_598,N_14994,N_14501);
nand UO_599 (O_599,N_14976,N_14915);
or UO_600 (O_600,N_14710,N_14780);
and UO_601 (O_601,N_14588,N_14694);
or UO_602 (O_602,N_14505,N_14768);
nand UO_603 (O_603,N_14613,N_14735);
or UO_604 (O_604,N_14567,N_14735);
or UO_605 (O_605,N_14643,N_14792);
nor UO_606 (O_606,N_14772,N_14806);
nand UO_607 (O_607,N_14796,N_14664);
xnor UO_608 (O_608,N_14691,N_14785);
xnor UO_609 (O_609,N_14744,N_14679);
xnor UO_610 (O_610,N_14537,N_14884);
nor UO_611 (O_611,N_14914,N_14769);
and UO_612 (O_612,N_14784,N_14720);
nand UO_613 (O_613,N_14542,N_14932);
xnor UO_614 (O_614,N_14876,N_14552);
or UO_615 (O_615,N_14948,N_14568);
or UO_616 (O_616,N_14900,N_14868);
nor UO_617 (O_617,N_14956,N_14648);
or UO_618 (O_618,N_14548,N_14531);
and UO_619 (O_619,N_14955,N_14727);
nor UO_620 (O_620,N_14887,N_14806);
nand UO_621 (O_621,N_14616,N_14890);
nand UO_622 (O_622,N_14659,N_14616);
nand UO_623 (O_623,N_14596,N_14809);
xor UO_624 (O_624,N_14586,N_14880);
or UO_625 (O_625,N_14883,N_14901);
xnor UO_626 (O_626,N_14972,N_14579);
nand UO_627 (O_627,N_14515,N_14971);
xor UO_628 (O_628,N_14816,N_14612);
nor UO_629 (O_629,N_14572,N_14629);
and UO_630 (O_630,N_14631,N_14741);
xnor UO_631 (O_631,N_14539,N_14928);
xor UO_632 (O_632,N_14633,N_14968);
xnor UO_633 (O_633,N_14609,N_14880);
nand UO_634 (O_634,N_14615,N_14583);
and UO_635 (O_635,N_14902,N_14710);
xor UO_636 (O_636,N_14650,N_14989);
and UO_637 (O_637,N_14686,N_14772);
nor UO_638 (O_638,N_14879,N_14650);
and UO_639 (O_639,N_14957,N_14702);
or UO_640 (O_640,N_14936,N_14716);
nor UO_641 (O_641,N_14509,N_14632);
nor UO_642 (O_642,N_14733,N_14724);
nor UO_643 (O_643,N_14598,N_14821);
nand UO_644 (O_644,N_14515,N_14571);
nand UO_645 (O_645,N_14863,N_14837);
nand UO_646 (O_646,N_14999,N_14861);
xor UO_647 (O_647,N_14887,N_14634);
nand UO_648 (O_648,N_14565,N_14949);
or UO_649 (O_649,N_14839,N_14590);
or UO_650 (O_650,N_14877,N_14637);
xnor UO_651 (O_651,N_14509,N_14609);
nor UO_652 (O_652,N_14598,N_14832);
nor UO_653 (O_653,N_14531,N_14814);
xnor UO_654 (O_654,N_14505,N_14556);
nand UO_655 (O_655,N_14644,N_14851);
or UO_656 (O_656,N_14899,N_14747);
and UO_657 (O_657,N_14533,N_14949);
nand UO_658 (O_658,N_14629,N_14670);
xnor UO_659 (O_659,N_14501,N_14656);
nand UO_660 (O_660,N_14820,N_14735);
or UO_661 (O_661,N_14950,N_14606);
nand UO_662 (O_662,N_14959,N_14722);
nand UO_663 (O_663,N_14617,N_14705);
nor UO_664 (O_664,N_14664,N_14901);
and UO_665 (O_665,N_14703,N_14736);
nand UO_666 (O_666,N_14742,N_14759);
nand UO_667 (O_667,N_14893,N_14763);
nor UO_668 (O_668,N_14722,N_14981);
nor UO_669 (O_669,N_14939,N_14867);
xnor UO_670 (O_670,N_14911,N_14909);
nand UO_671 (O_671,N_14519,N_14667);
nor UO_672 (O_672,N_14860,N_14734);
and UO_673 (O_673,N_14806,N_14900);
and UO_674 (O_674,N_14570,N_14629);
nand UO_675 (O_675,N_14699,N_14821);
xnor UO_676 (O_676,N_14976,N_14607);
nor UO_677 (O_677,N_14915,N_14504);
or UO_678 (O_678,N_14731,N_14839);
or UO_679 (O_679,N_14696,N_14513);
xnor UO_680 (O_680,N_14821,N_14998);
and UO_681 (O_681,N_14927,N_14671);
nor UO_682 (O_682,N_14502,N_14567);
xor UO_683 (O_683,N_14623,N_14644);
and UO_684 (O_684,N_14982,N_14878);
nand UO_685 (O_685,N_14856,N_14795);
xor UO_686 (O_686,N_14973,N_14522);
xor UO_687 (O_687,N_14633,N_14917);
nor UO_688 (O_688,N_14793,N_14510);
xor UO_689 (O_689,N_14658,N_14579);
nor UO_690 (O_690,N_14562,N_14646);
and UO_691 (O_691,N_14835,N_14677);
nand UO_692 (O_692,N_14693,N_14887);
xnor UO_693 (O_693,N_14745,N_14513);
xnor UO_694 (O_694,N_14961,N_14562);
nand UO_695 (O_695,N_14838,N_14680);
xor UO_696 (O_696,N_14992,N_14916);
or UO_697 (O_697,N_14919,N_14750);
and UO_698 (O_698,N_14890,N_14591);
nor UO_699 (O_699,N_14534,N_14588);
xnor UO_700 (O_700,N_14855,N_14787);
or UO_701 (O_701,N_14799,N_14730);
nand UO_702 (O_702,N_14890,N_14550);
nor UO_703 (O_703,N_14772,N_14701);
nand UO_704 (O_704,N_14973,N_14828);
or UO_705 (O_705,N_14669,N_14575);
or UO_706 (O_706,N_14763,N_14745);
nand UO_707 (O_707,N_14678,N_14914);
or UO_708 (O_708,N_14598,N_14798);
nor UO_709 (O_709,N_14818,N_14843);
and UO_710 (O_710,N_14980,N_14503);
nor UO_711 (O_711,N_14667,N_14651);
and UO_712 (O_712,N_14634,N_14706);
or UO_713 (O_713,N_14620,N_14757);
and UO_714 (O_714,N_14545,N_14728);
xor UO_715 (O_715,N_14677,N_14637);
xnor UO_716 (O_716,N_14657,N_14876);
xor UO_717 (O_717,N_14597,N_14672);
nand UO_718 (O_718,N_14762,N_14526);
xor UO_719 (O_719,N_14765,N_14709);
nand UO_720 (O_720,N_14750,N_14535);
and UO_721 (O_721,N_14648,N_14901);
nand UO_722 (O_722,N_14502,N_14645);
nor UO_723 (O_723,N_14831,N_14822);
xnor UO_724 (O_724,N_14996,N_14675);
nand UO_725 (O_725,N_14629,N_14749);
and UO_726 (O_726,N_14605,N_14822);
nand UO_727 (O_727,N_14708,N_14887);
nand UO_728 (O_728,N_14657,N_14565);
nor UO_729 (O_729,N_14644,N_14545);
nor UO_730 (O_730,N_14787,N_14842);
nand UO_731 (O_731,N_14603,N_14752);
nand UO_732 (O_732,N_14503,N_14854);
nor UO_733 (O_733,N_14688,N_14977);
and UO_734 (O_734,N_14772,N_14593);
xnor UO_735 (O_735,N_14873,N_14785);
nor UO_736 (O_736,N_14634,N_14619);
xnor UO_737 (O_737,N_14808,N_14855);
nor UO_738 (O_738,N_14966,N_14699);
nand UO_739 (O_739,N_14955,N_14553);
xor UO_740 (O_740,N_14664,N_14956);
nor UO_741 (O_741,N_14689,N_14541);
or UO_742 (O_742,N_14939,N_14994);
and UO_743 (O_743,N_14539,N_14580);
xor UO_744 (O_744,N_14856,N_14574);
or UO_745 (O_745,N_14881,N_14563);
nand UO_746 (O_746,N_14888,N_14571);
xnor UO_747 (O_747,N_14827,N_14814);
or UO_748 (O_748,N_14654,N_14516);
and UO_749 (O_749,N_14945,N_14692);
xnor UO_750 (O_750,N_14525,N_14840);
nor UO_751 (O_751,N_14697,N_14715);
and UO_752 (O_752,N_14540,N_14990);
nand UO_753 (O_753,N_14768,N_14611);
or UO_754 (O_754,N_14980,N_14596);
nor UO_755 (O_755,N_14767,N_14580);
xnor UO_756 (O_756,N_14673,N_14565);
nor UO_757 (O_757,N_14998,N_14720);
xnor UO_758 (O_758,N_14788,N_14810);
and UO_759 (O_759,N_14681,N_14665);
nand UO_760 (O_760,N_14931,N_14987);
nor UO_761 (O_761,N_14705,N_14654);
and UO_762 (O_762,N_14667,N_14714);
xnor UO_763 (O_763,N_14786,N_14728);
nand UO_764 (O_764,N_14592,N_14896);
nor UO_765 (O_765,N_14760,N_14996);
or UO_766 (O_766,N_14797,N_14623);
and UO_767 (O_767,N_14670,N_14530);
xnor UO_768 (O_768,N_14986,N_14596);
nand UO_769 (O_769,N_14790,N_14959);
nor UO_770 (O_770,N_14602,N_14897);
nor UO_771 (O_771,N_14903,N_14758);
nor UO_772 (O_772,N_14809,N_14517);
xor UO_773 (O_773,N_14752,N_14604);
xnor UO_774 (O_774,N_14890,N_14708);
and UO_775 (O_775,N_14504,N_14647);
or UO_776 (O_776,N_14748,N_14802);
or UO_777 (O_777,N_14835,N_14743);
nor UO_778 (O_778,N_14782,N_14614);
or UO_779 (O_779,N_14729,N_14911);
xor UO_780 (O_780,N_14844,N_14907);
nand UO_781 (O_781,N_14854,N_14812);
nor UO_782 (O_782,N_14702,N_14528);
and UO_783 (O_783,N_14503,N_14640);
and UO_784 (O_784,N_14694,N_14621);
and UO_785 (O_785,N_14814,N_14846);
or UO_786 (O_786,N_14597,N_14720);
xnor UO_787 (O_787,N_14561,N_14715);
nor UO_788 (O_788,N_14521,N_14595);
or UO_789 (O_789,N_14763,N_14804);
nor UO_790 (O_790,N_14915,N_14533);
xnor UO_791 (O_791,N_14558,N_14810);
and UO_792 (O_792,N_14658,N_14657);
nand UO_793 (O_793,N_14831,N_14969);
xnor UO_794 (O_794,N_14605,N_14649);
nand UO_795 (O_795,N_14924,N_14719);
nor UO_796 (O_796,N_14873,N_14999);
or UO_797 (O_797,N_14993,N_14958);
or UO_798 (O_798,N_14724,N_14991);
xnor UO_799 (O_799,N_14558,N_14817);
xnor UO_800 (O_800,N_14966,N_14501);
or UO_801 (O_801,N_14516,N_14558);
and UO_802 (O_802,N_14749,N_14805);
or UO_803 (O_803,N_14531,N_14630);
or UO_804 (O_804,N_14807,N_14756);
nor UO_805 (O_805,N_14770,N_14924);
xnor UO_806 (O_806,N_14782,N_14902);
and UO_807 (O_807,N_14645,N_14823);
nand UO_808 (O_808,N_14919,N_14814);
nand UO_809 (O_809,N_14907,N_14677);
nor UO_810 (O_810,N_14655,N_14754);
and UO_811 (O_811,N_14935,N_14701);
nand UO_812 (O_812,N_14590,N_14971);
xor UO_813 (O_813,N_14534,N_14676);
and UO_814 (O_814,N_14856,N_14865);
nand UO_815 (O_815,N_14553,N_14567);
nor UO_816 (O_816,N_14864,N_14941);
and UO_817 (O_817,N_14632,N_14633);
xor UO_818 (O_818,N_14552,N_14726);
nor UO_819 (O_819,N_14639,N_14700);
nor UO_820 (O_820,N_14829,N_14730);
nand UO_821 (O_821,N_14906,N_14840);
and UO_822 (O_822,N_14764,N_14970);
xnor UO_823 (O_823,N_14756,N_14645);
or UO_824 (O_824,N_14820,N_14666);
xor UO_825 (O_825,N_14558,N_14725);
nand UO_826 (O_826,N_14610,N_14642);
nand UO_827 (O_827,N_14790,N_14538);
nand UO_828 (O_828,N_14911,N_14871);
and UO_829 (O_829,N_14704,N_14675);
and UO_830 (O_830,N_14632,N_14873);
or UO_831 (O_831,N_14608,N_14739);
or UO_832 (O_832,N_14959,N_14754);
or UO_833 (O_833,N_14783,N_14828);
or UO_834 (O_834,N_14850,N_14949);
xor UO_835 (O_835,N_14707,N_14536);
nand UO_836 (O_836,N_14843,N_14668);
or UO_837 (O_837,N_14838,N_14868);
or UO_838 (O_838,N_14824,N_14667);
xor UO_839 (O_839,N_14531,N_14803);
xnor UO_840 (O_840,N_14545,N_14563);
or UO_841 (O_841,N_14928,N_14702);
or UO_842 (O_842,N_14542,N_14867);
nor UO_843 (O_843,N_14763,N_14710);
and UO_844 (O_844,N_14549,N_14855);
or UO_845 (O_845,N_14763,N_14734);
and UO_846 (O_846,N_14611,N_14877);
nor UO_847 (O_847,N_14986,N_14518);
or UO_848 (O_848,N_14567,N_14839);
or UO_849 (O_849,N_14956,N_14884);
nand UO_850 (O_850,N_14622,N_14563);
xor UO_851 (O_851,N_14594,N_14926);
nand UO_852 (O_852,N_14878,N_14980);
xor UO_853 (O_853,N_14854,N_14673);
xor UO_854 (O_854,N_14888,N_14564);
and UO_855 (O_855,N_14784,N_14661);
nand UO_856 (O_856,N_14605,N_14559);
or UO_857 (O_857,N_14703,N_14501);
xor UO_858 (O_858,N_14763,N_14691);
xnor UO_859 (O_859,N_14613,N_14577);
nor UO_860 (O_860,N_14537,N_14875);
nand UO_861 (O_861,N_14638,N_14992);
nand UO_862 (O_862,N_14575,N_14614);
nand UO_863 (O_863,N_14599,N_14880);
xor UO_864 (O_864,N_14976,N_14871);
or UO_865 (O_865,N_14789,N_14688);
nand UO_866 (O_866,N_14983,N_14925);
or UO_867 (O_867,N_14681,N_14645);
nor UO_868 (O_868,N_14628,N_14879);
xor UO_869 (O_869,N_14595,N_14621);
and UO_870 (O_870,N_14538,N_14612);
and UO_871 (O_871,N_14528,N_14563);
and UO_872 (O_872,N_14550,N_14618);
nor UO_873 (O_873,N_14753,N_14854);
nand UO_874 (O_874,N_14911,N_14691);
or UO_875 (O_875,N_14693,N_14635);
and UO_876 (O_876,N_14952,N_14512);
or UO_877 (O_877,N_14888,N_14672);
or UO_878 (O_878,N_14595,N_14628);
or UO_879 (O_879,N_14579,N_14887);
xnor UO_880 (O_880,N_14720,N_14931);
xnor UO_881 (O_881,N_14687,N_14890);
xor UO_882 (O_882,N_14938,N_14940);
nand UO_883 (O_883,N_14666,N_14813);
xnor UO_884 (O_884,N_14531,N_14895);
nand UO_885 (O_885,N_14715,N_14836);
and UO_886 (O_886,N_14770,N_14753);
xor UO_887 (O_887,N_14621,N_14770);
nand UO_888 (O_888,N_14945,N_14519);
and UO_889 (O_889,N_14780,N_14559);
nor UO_890 (O_890,N_14834,N_14908);
or UO_891 (O_891,N_14523,N_14975);
nor UO_892 (O_892,N_14935,N_14625);
or UO_893 (O_893,N_14994,N_14869);
or UO_894 (O_894,N_14685,N_14536);
and UO_895 (O_895,N_14613,N_14659);
xor UO_896 (O_896,N_14968,N_14738);
and UO_897 (O_897,N_14576,N_14926);
and UO_898 (O_898,N_14896,N_14534);
nor UO_899 (O_899,N_14846,N_14858);
nor UO_900 (O_900,N_14956,N_14982);
and UO_901 (O_901,N_14819,N_14566);
nor UO_902 (O_902,N_14867,N_14768);
nor UO_903 (O_903,N_14742,N_14978);
nor UO_904 (O_904,N_14802,N_14823);
xor UO_905 (O_905,N_14610,N_14708);
and UO_906 (O_906,N_14743,N_14724);
and UO_907 (O_907,N_14772,N_14668);
or UO_908 (O_908,N_14938,N_14582);
nor UO_909 (O_909,N_14538,N_14903);
nand UO_910 (O_910,N_14860,N_14599);
xnor UO_911 (O_911,N_14857,N_14504);
and UO_912 (O_912,N_14762,N_14603);
nor UO_913 (O_913,N_14511,N_14919);
xor UO_914 (O_914,N_14818,N_14731);
or UO_915 (O_915,N_14647,N_14911);
xor UO_916 (O_916,N_14982,N_14852);
nand UO_917 (O_917,N_14503,N_14769);
nor UO_918 (O_918,N_14868,N_14594);
nand UO_919 (O_919,N_14907,N_14730);
xnor UO_920 (O_920,N_14782,N_14539);
nor UO_921 (O_921,N_14671,N_14779);
nor UO_922 (O_922,N_14664,N_14698);
xnor UO_923 (O_923,N_14596,N_14959);
nand UO_924 (O_924,N_14510,N_14532);
nand UO_925 (O_925,N_14793,N_14654);
xor UO_926 (O_926,N_14894,N_14784);
nand UO_927 (O_927,N_14682,N_14727);
or UO_928 (O_928,N_14729,N_14766);
or UO_929 (O_929,N_14526,N_14883);
xnor UO_930 (O_930,N_14690,N_14508);
and UO_931 (O_931,N_14886,N_14776);
nor UO_932 (O_932,N_14754,N_14598);
and UO_933 (O_933,N_14703,N_14969);
nand UO_934 (O_934,N_14723,N_14545);
and UO_935 (O_935,N_14712,N_14750);
nand UO_936 (O_936,N_14833,N_14999);
nand UO_937 (O_937,N_14795,N_14887);
nor UO_938 (O_938,N_14635,N_14689);
nand UO_939 (O_939,N_14517,N_14555);
nor UO_940 (O_940,N_14540,N_14837);
nor UO_941 (O_941,N_14504,N_14888);
xor UO_942 (O_942,N_14503,N_14560);
and UO_943 (O_943,N_14913,N_14641);
nand UO_944 (O_944,N_14789,N_14868);
or UO_945 (O_945,N_14870,N_14672);
and UO_946 (O_946,N_14814,N_14774);
nand UO_947 (O_947,N_14898,N_14883);
and UO_948 (O_948,N_14869,N_14928);
nor UO_949 (O_949,N_14701,N_14951);
nand UO_950 (O_950,N_14797,N_14767);
xnor UO_951 (O_951,N_14506,N_14715);
nor UO_952 (O_952,N_14502,N_14959);
xor UO_953 (O_953,N_14775,N_14630);
or UO_954 (O_954,N_14755,N_14819);
or UO_955 (O_955,N_14657,N_14544);
or UO_956 (O_956,N_14660,N_14883);
nand UO_957 (O_957,N_14782,N_14665);
nand UO_958 (O_958,N_14634,N_14899);
or UO_959 (O_959,N_14877,N_14779);
or UO_960 (O_960,N_14908,N_14510);
and UO_961 (O_961,N_14828,N_14733);
or UO_962 (O_962,N_14734,N_14857);
and UO_963 (O_963,N_14866,N_14542);
and UO_964 (O_964,N_14594,N_14751);
xor UO_965 (O_965,N_14581,N_14532);
and UO_966 (O_966,N_14811,N_14958);
xor UO_967 (O_967,N_14614,N_14627);
nand UO_968 (O_968,N_14913,N_14738);
nor UO_969 (O_969,N_14918,N_14570);
and UO_970 (O_970,N_14817,N_14774);
nand UO_971 (O_971,N_14713,N_14812);
nor UO_972 (O_972,N_14716,N_14530);
and UO_973 (O_973,N_14832,N_14865);
and UO_974 (O_974,N_14513,N_14946);
or UO_975 (O_975,N_14745,N_14769);
and UO_976 (O_976,N_14618,N_14842);
or UO_977 (O_977,N_14847,N_14556);
nor UO_978 (O_978,N_14585,N_14975);
and UO_979 (O_979,N_14690,N_14716);
xor UO_980 (O_980,N_14545,N_14797);
and UO_981 (O_981,N_14805,N_14726);
and UO_982 (O_982,N_14736,N_14525);
xnor UO_983 (O_983,N_14801,N_14871);
xnor UO_984 (O_984,N_14953,N_14889);
and UO_985 (O_985,N_14991,N_14814);
or UO_986 (O_986,N_14769,N_14768);
nand UO_987 (O_987,N_14600,N_14914);
or UO_988 (O_988,N_14532,N_14574);
xnor UO_989 (O_989,N_14579,N_14512);
and UO_990 (O_990,N_14987,N_14942);
and UO_991 (O_991,N_14912,N_14600);
nand UO_992 (O_992,N_14805,N_14708);
or UO_993 (O_993,N_14943,N_14800);
and UO_994 (O_994,N_14722,N_14987);
nand UO_995 (O_995,N_14553,N_14575);
and UO_996 (O_996,N_14815,N_14659);
and UO_997 (O_997,N_14603,N_14764);
and UO_998 (O_998,N_14952,N_14591);
nand UO_999 (O_999,N_14830,N_14636);
nand UO_1000 (O_1000,N_14987,N_14713);
and UO_1001 (O_1001,N_14671,N_14981);
xnor UO_1002 (O_1002,N_14693,N_14889);
xnor UO_1003 (O_1003,N_14674,N_14979);
nand UO_1004 (O_1004,N_14995,N_14981);
nor UO_1005 (O_1005,N_14972,N_14780);
nor UO_1006 (O_1006,N_14513,N_14984);
or UO_1007 (O_1007,N_14576,N_14552);
or UO_1008 (O_1008,N_14628,N_14602);
nor UO_1009 (O_1009,N_14676,N_14983);
nor UO_1010 (O_1010,N_14514,N_14522);
and UO_1011 (O_1011,N_14839,N_14608);
xnor UO_1012 (O_1012,N_14629,N_14695);
and UO_1013 (O_1013,N_14847,N_14681);
and UO_1014 (O_1014,N_14535,N_14540);
nand UO_1015 (O_1015,N_14914,N_14561);
or UO_1016 (O_1016,N_14785,N_14730);
or UO_1017 (O_1017,N_14661,N_14606);
nor UO_1018 (O_1018,N_14569,N_14931);
or UO_1019 (O_1019,N_14740,N_14926);
xnor UO_1020 (O_1020,N_14672,N_14725);
or UO_1021 (O_1021,N_14819,N_14821);
xor UO_1022 (O_1022,N_14792,N_14502);
xor UO_1023 (O_1023,N_14751,N_14788);
nand UO_1024 (O_1024,N_14541,N_14596);
or UO_1025 (O_1025,N_14890,N_14822);
nor UO_1026 (O_1026,N_14750,N_14660);
nand UO_1027 (O_1027,N_14635,N_14922);
or UO_1028 (O_1028,N_14945,N_14638);
nor UO_1029 (O_1029,N_14756,N_14539);
or UO_1030 (O_1030,N_14975,N_14876);
xor UO_1031 (O_1031,N_14678,N_14523);
xor UO_1032 (O_1032,N_14886,N_14703);
xnor UO_1033 (O_1033,N_14804,N_14543);
or UO_1034 (O_1034,N_14767,N_14783);
or UO_1035 (O_1035,N_14588,N_14565);
and UO_1036 (O_1036,N_14764,N_14559);
or UO_1037 (O_1037,N_14754,N_14961);
nor UO_1038 (O_1038,N_14999,N_14649);
xnor UO_1039 (O_1039,N_14513,N_14857);
nand UO_1040 (O_1040,N_14975,N_14580);
xnor UO_1041 (O_1041,N_14803,N_14678);
xnor UO_1042 (O_1042,N_14522,N_14651);
nand UO_1043 (O_1043,N_14585,N_14611);
nor UO_1044 (O_1044,N_14829,N_14617);
nand UO_1045 (O_1045,N_14717,N_14810);
nand UO_1046 (O_1046,N_14835,N_14542);
and UO_1047 (O_1047,N_14560,N_14975);
nand UO_1048 (O_1048,N_14954,N_14603);
or UO_1049 (O_1049,N_14979,N_14901);
nand UO_1050 (O_1050,N_14988,N_14993);
nor UO_1051 (O_1051,N_14506,N_14643);
nand UO_1052 (O_1052,N_14536,N_14743);
nand UO_1053 (O_1053,N_14511,N_14925);
nor UO_1054 (O_1054,N_14716,N_14666);
xor UO_1055 (O_1055,N_14517,N_14823);
nor UO_1056 (O_1056,N_14902,N_14519);
xnor UO_1057 (O_1057,N_14993,N_14548);
nand UO_1058 (O_1058,N_14933,N_14629);
xnor UO_1059 (O_1059,N_14693,N_14736);
xor UO_1060 (O_1060,N_14797,N_14541);
nor UO_1061 (O_1061,N_14931,N_14545);
or UO_1062 (O_1062,N_14900,N_14512);
and UO_1063 (O_1063,N_14780,N_14634);
xnor UO_1064 (O_1064,N_14637,N_14699);
xor UO_1065 (O_1065,N_14529,N_14759);
or UO_1066 (O_1066,N_14808,N_14810);
xnor UO_1067 (O_1067,N_14531,N_14712);
and UO_1068 (O_1068,N_14513,N_14615);
or UO_1069 (O_1069,N_14545,N_14626);
nand UO_1070 (O_1070,N_14776,N_14827);
xnor UO_1071 (O_1071,N_14668,N_14601);
nand UO_1072 (O_1072,N_14808,N_14661);
and UO_1073 (O_1073,N_14667,N_14951);
xnor UO_1074 (O_1074,N_14688,N_14976);
nand UO_1075 (O_1075,N_14803,N_14542);
xor UO_1076 (O_1076,N_14711,N_14908);
or UO_1077 (O_1077,N_14647,N_14727);
nand UO_1078 (O_1078,N_14722,N_14576);
xnor UO_1079 (O_1079,N_14595,N_14578);
nor UO_1080 (O_1080,N_14875,N_14688);
xnor UO_1081 (O_1081,N_14782,N_14751);
nor UO_1082 (O_1082,N_14723,N_14967);
nand UO_1083 (O_1083,N_14771,N_14658);
or UO_1084 (O_1084,N_14940,N_14613);
and UO_1085 (O_1085,N_14512,N_14829);
and UO_1086 (O_1086,N_14642,N_14637);
and UO_1087 (O_1087,N_14868,N_14763);
nand UO_1088 (O_1088,N_14826,N_14838);
xnor UO_1089 (O_1089,N_14921,N_14667);
or UO_1090 (O_1090,N_14605,N_14867);
xnor UO_1091 (O_1091,N_14575,N_14537);
or UO_1092 (O_1092,N_14659,N_14918);
nor UO_1093 (O_1093,N_14795,N_14741);
or UO_1094 (O_1094,N_14572,N_14534);
xnor UO_1095 (O_1095,N_14827,N_14748);
xor UO_1096 (O_1096,N_14814,N_14994);
nand UO_1097 (O_1097,N_14703,N_14620);
xnor UO_1098 (O_1098,N_14696,N_14990);
xor UO_1099 (O_1099,N_14561,N_14822);
or UO_1100 (O_1100,N_14784,N_14978);
and UO_1101 (O_1101,N_14985,N_14794);
or UO_1102 (O_1102,N_14954,N_14901);
nor UO_1103 (O_1103,N_14949,N_14888);
nor UO_1104 (O_1104,N_14977,N_14579);
nand UO_1105 (O_1105,N_14929,N_14611);
and UO_1106 (O_1106,N_14582,N_14751);
nor UO_1107 (O_1107,N_14895,N_14696);
or UO_1108 (O_1108,N_14518,N_14612);
nand UO_1109 (O_1109,N_14956,N_14914);
xor UO_1110 (O_1110,N_14961,N_14793);
nor UO_1111 (O_1111,N_14847,N_14768);
xor UO_1112 (O_1112,N_14695,N_14565);
nand UO_1113 (O_1113,N_14739,N_14784);
xor UO_1114 (O_1114,N_14697,N_14706);
or UO_1115 (O_1115,N_14970,N_14873);
nand UO_1116 (O_1116,N_14699,N_14776);
nor UO_1117 (O_1117,N_14592,N_14563);
xor UO_1118 (O_1118,N_14737,N_14942);
nor UO_1119 (O_1119,N_14962,N_14905);
xnor UO_1120 (O_1120,N_14975,N_14674);
and UO_1121 (O_1121,N_14990,N_14761);
and UO_1122 (O_1122,N_14848,N_14799);
xnor UO_1123 (O_1123,N_14758,N_14898);
xor UO_1124 (O_1124,N_14570,N_14771);
or UO_1125 (O_1125,N_14837,N_14972);
and UO_1126 (O_1126,N_14927,N_14724);
and UO_1127 (O_1127,N_14859,N_14957);
and UO_1128 (O_1128,N_14565,N_14604);
or UO_1129 (O_1129,N_14966,N_14529);
nor UO_1130 (O_1130,N_14557,N_14754);
nor UO_1131 (O_1131,N_14546,N_14857);
and UO_1132 (O_1132,N_14868,N_14685);
nor UO_1133 (O_1133,N_14786,N_14930);
nand UO_1134 (O_1134,N_14660,N_14684);
xor UO_1135 (O_1135,N_14915,N_14706);
xnor UO_1136 (O_1136,N_14768,N_14647);
nor UO_1137 (O_1137,N_14869,N_14621);
nor UO_1138 (O_1138,N_14964,N_14501);
nor UO_1139 (O_1139,N_14857,N_14564);
xor UO_1140 (O_1140,N_14985,N_14829);
nand UO_1141 (O_1141,N_14635,N_14540);
and UO_1142 (O_1142,N_14534,N_14705);
nand UO_1143 (O_1143,N_14730,N_14559);
or UO_1144 (O_1144,N_14742,N_14777);
xnor UO_1145 (O_1145,N_14501,N_14878);
nand UO_1146 (O_1146,N_14774,N_14849);
or UO_1147 (O_1147,N_14522,N_14633);
and UO_1148 (O_1148,N_14901,N_14974);
and UO_1149 (O_1149,N_14907,N_14952);
nor UO_1150 (O_1150,N_14814,N_14918);
or UO_1151 (O_1151,N_14958,N_14505);
nor UO_1152 (O_1152,N_14533,N_14832);
nand UO_1153 (O_1153,N_14912,N_14782);
nor UO_1154 (O_1154,N_14821,N_14927);
or UO_1155 (O_1155,N_14678,N_14957);
or UO_1156 (O_1156,N_14890,N_14990);
and UO_1157 (O_1157,N_14688,N_14907);
or UO_1158 (O_1158,N_14556,N_14815);
nor UO_1159 (O_1159,N_14708,N_14875);
or UO_1160 (O_1160,N_14999,N_14828);
and UO_1161 (O_1161,N_14999,N_14826);
or UO_1162 (O_1162,N_14575,N_14554);
and UO_1163 (O_1163,N_14768,N_14551);
nand UO_1164 (O_1164,N_14934,N_14957);
or UO_1165 (O_1165,N_14867,N_14721);
xnor UO_1166 (O_1166,N_14789,N_14648);
nand UO_1167 (O_1167,N_14547,N_14862);
nand UO_1168 (O_1168,N_14546,N_14516);
nor UO_1169 (O_1169,N_14761,N_14653);
nand UO_1170 (O_1170,N_14745,N_14695);
and UO_1171 (O_1171,N_14970,N_14721);
xor UO_1172 (O_1172,N_14757,N_14630);
or UO_1173 (O_1173,N_14674,N_14916);
nand UO_1174 (O_1174,N_14987,N_14972);
xor UO_1175 (O_1175,N_14644,N_14907);
nor UO_1176 (O_1176,N_14881,N_14679);
or UO_1177 (O_1177,N_14779,N_14642);
nor UO_1178 (O_1178,N_14804,N_14602);
or UO_1179 (O_1179,N_14767,N_14941);
nand UO_1180 (O_1180,N_14787,N_14545);
and UO_1181 (O_1181,N_14561,N_14931);
and UO_1182 (O_1182,N_14801,N_14560);
or UO_1183 (O_1183,N_14865,N_14909);
nor UO_1184 (O_1184,N_14805,N_14950);
or UO_1185 (O_1185,N_14781,N_14617);
or UO_1186 (O_1186,N_14728,N_14952);
xor UO_1187 (O_1187,N_14603,N_14635);
or UO_1188 (O_1188,N_14795,N_14558);
nor UO_1189 (O_1189,N_14523,N_14613);
xnor UO_1190 (O_1190,N_14597,N_14609);
xor UO_1191 (O_1191,N_14758,N_14638);
or UO_1192 (O_1192,N_14756,N_14738);
xor UO_1193 (O_1193,N_14647,N_14683);
xor UO_1194 (O_1194,N_14785,N_14538);
xnor UO_1195 (O_1195,N_14624,N_14623);
or UO_1196 (O_1196,N_14614,N_14777);
nand UO_1197 (O_1197,N_14806,N_14778);
and UO_1198 (O_1198,N_14708,N_14710);
or UO_1199 (O_1199,N_14544,N_14940);
xor UO_1200 (O_1200,N_14542,N_14513);
nand UO_1201 (O_1201,N_14518,N_14963);
nand UO_1202 (O_1202,N_14692,N_14738);
nor UO_1203 (O_1203,N_14795,N_14906);
xor UO_1204 (O_1204,N_14524,N_14971);
and UO_1205 (O_1205,N_14903,N_14749);
xnor UO_1206 (O_1206,N_14739,N_14520);
and UO_1207 (O_1207,N_14702,N_14984);
nand UO_1208 (O_1208,N_14757,N_14654);
or UO_1209 (O_1209,N_14889,N_14900);
nand UO_1210 (O_1210,N_14892,N_14729);
or UO_1211 (O_1211,N_14932,N_14769);
and UO_1212 (O_1212,N_14527,N_14941);
nand UO_1213 (O_1213,N_14785,N_14521);
nand UO_1214 (O_1214,N_14819,N_14929);
nand UO_1215 (O_1215,N_14783,N_14812);
nand UO_1216 (O_1216,N_14948,N_14527);
xnor UO_1217 (O_1217,N_14599,N_14885);
or UO_1218 (O_1218,N_14973,N_14573);
nand UO_1219 (O_1219,N_14967,N_14845);
xor UO_1220 (O_1220,N_14647,N_14935);
nor UO_1221 (O_1221,N_14586,N_14604);
nor UO_1222 (O_1222,N_14798,N_14938);
xor UO_1223 (O_1223,N_14800,N_14607);
nor UO_1224 (O_1224,N_14914,N_14918);
nand UO_1225 (O_1225,N_14980,N_14748);
nand UO_1226 (O_1226,N_14669,N_14548);
nand UO_1227 (O_1227,N_14968,N_14539);
and UO_1228 (O_1228,N_14516,N_14879);
and UO_1229 (O_1229,N_14748,N_14596);
nand UO_1230 (O_1230,N_14657,N_14602);
and UO_1231 (O_1231,N_14579,N_14759);
nor UO_1232 (O_1232,N_14662,N_14945);
and UO_1233 (O_1233,N_14535,N_14756);
nor UO_1234 (O_1234,N_14961,N_14791);
xor UO_1235 (O_1235,N_14651,N_14884);
xnor UO_1236 (O_1236,N_14938,N_14520);
nand UO_1237 (O_1237,N_14756,N_14995);
xnor UO_1238 (O_1238,N_14780,N_14866);
xor UO_1239 (O_1239,N_14907,N_14711);
or UO_1240 (O_1240,N_14911,N_14633);
nand UO_1241 (O_1241,N_14919,N_14755);
nand UO_1242 (O_1242,N_14636,N_14505);
xnor UO_1243 (O_1243,N_14958,N_14968);
nor UO_1244 (O_1244,N_14658,N_14540);
or UO_1245 (O_1245,N_14868,N_14747);
nor UO_1246 (O_1246,N_14928,N_14668);
xnor UO_1247 (O_1247,N_14782,N_14656);
and UO_1248 (O_1248,N_14907,N_14578);
xor UO_1249 (O_1249,N_14880,N_14865);
and UO_1250 (O_1250,N_14705,N_14598);
nand UO_1251 (O_1251,N_14878,N_14549);
xnor UO_1252 (O_1252,N_14891,N_14534);
or UO_1253 (O_1253,N_14637,N_14951);
and UO_1254 (O_1254,N_14923,N_14835);
and UO_1255 (O_1255,N_14974,N_14849);
and UO_1256 (O_1256,N_14647,N_14946);
xor UO_1257 (O_1257,N_14620,N_14675);
xnor UO_1258 (O_1258,N_14561,N_14623);
or UO_1259 (O_1259,N_14748,N_14546);
nand UO_1260 (O_1260,N_14861,N_14939);
nand UO_1261 (O_1261,N_14900,N_14617);
nand UO_1262 (O_1262,N_14792,N_14763);
or UO_1263 (O_1263,N_14921,N_14683);
or UO_1264 (O_1264,N_14883,N_14791);
or UO_1265 (O_1265,N_14997,N_14756);
xnor UO_1266 (O_1266,N_14613,N_14681);
or UO_1267 (O_1267,N_14581,N_14983);
or UO_1268 (O_1268,N_14643,N_14714);
xnor UO_1269 (O_1269,N_14982,N_14914);
xor UO_1270 (O_1270,N_14557,N_14763);
and UO_1271 (O_1271,N_14598,N_14872);
and UO_1272 (O_1272,N_14562,N_14977);
nand UO_1273 (O_1273,N_14628,N_14982);
and UO_1274 (O_1274,N_14696,N_14672);
xor UO_1275 (O_1275,N_14883,N_14759);
and UO_1276 (O_1276,N_14665,N_14741);
nand UO_1277 (O_1277,N_14715,N_14829);
and UO_1278 (O_1278,N_14512,N_14569);
or UO_1279 (O_1279,N_14637,N_14596);
nand UO_1280 (O_1280,N_14856,N_14994);
nor UO_1281 (O_1281,N_14861,N_14545);
xor UO_1282 (O_1282,N_14500,N_14852);
xor UO_1283 (O_1283,N_14671,N_14703);
nor UO_1284 (O_1284,N_14610,N_14963);
xor UO_1285 (O_1285,N_14846,N_14832);
or UO_1286 (O_1286,N_14690,N_14687);
nand UO_1287 (O_1287,N_14542,N_14751);
or UO_1288 (O_1288,N_14568,N_14593);
or UO_1289 (O_1289,N_14939,N_14790);
xnor UO_1290 (O_1290,N_14506,N_14843);
or UO_1291 (O_1291,N_14765,N_14580);
nor UO_1292 (O_1292,N_14946,N_14577);
nor UO_1293 (O_1293,N_14786,N_14905);
nand UO_1294 (O_1294,N_14595,N_14602);
and UO_1295 (O_1295,N_14566,N_14773);
nor UO_1296 (O_1296,N_14615,N_14664);
or UO_1297 (O_1297,N_14816,N_14945);
xor UO_1298 (O_1298,N_14593,N_14950);
or UO_1299 (O_1299,N_14636,N_14535);
or UO_1300 (O_1300,N_14951,N_14552);
or UO_1301 (O_1301,N_14982,N_14570);
and UO_1302 (O_1302,N_14994,N_14750);
nor UO_1303 (O_1303,N_14738,N_14966);
or UO_1304 (O_1304,N_14740,N_14856);
and UO_1305 (O_1305,N_14512,N_14588);
nand UO_1306 (O_1306,N_14864,N_14704);
nand UO_1307 (O_1307,N_14631,N_14627);
nor UO_1308 (O_1308,N_14882,N_14776);
nand UO_1309 (O_1309,N_14819,N_14842);
xor UO_1310 (O_1310,N_14614,N_14728);
xor UO_1311 (O_1311,N_14672,N_14517);
and UO_1312 (O_1312,N_14633,N_14999);
nand UO_1313 (O_1313,N_14852,N_14965);
nand UO_1314 (O_1314,N_14532,N_14577);
or UO_1315 (O_1315,N_14922,N_14699);
xor UO_1316 (O_1316,N_14590,N_14661);
and UO_1317 (O_1317,N_14596,N_14820);
nand UO_1318 (O_1318,N_14751,N_14881);
nand UO_1319 (O_1319,N_14695,N_14671);
or UO_1320 (O_1320,N_14943,N_14817);
or UO_1321 (O_1321,N_14979,N_14868);
nand UO_1322 (O_1322,N_14621,N_14835);
nand UO_1323 (O_1323,N_14929,N_14589);
or UO_1324 (O_1324,N_14810,N_14643);
or UO_1325 (O_1325,N_14595,N_14719);
xor UO_1326 (O_1326,N_14704,N_14693);
nand UO_1327 (O_1327,N_14681,N_14892);
nor UO_1328 (O_1328,N_14687,N_14875);
and UO_1329 (O_1329,N_14754,N_14912);
xnor UO_1330 (O_1330,N_14600,N_14748);
nor UO_1331 (O_1331,N_14599,N_14919);
or UO_1332 (O_1332,N_14673,N_14877);
or UO_1333 (O_1333,N_14727,N_14646);
and UO_1334 (O_1334,N_14571,N_14823);
nor UO_1335 (O_1335,N_14506,N_14664);
nand UO_1336 (O_1336,N_14641,N_14768);
nand UO_1337 (O_1337,N_14746,N_14736);
nand UO_1338 (O_1338,N_14560,N_14923);
xnor UO_1339 (O_1339,N_14996,N_14953);
or UO_1340 (O_1340,N_14920,N_14632);
nand UO_1341 (O_1341,N_14657,N_14895);
nand UO_1342 (O_1342,N_14563,N_14937);
and UO_1343 (O_1343,N_14655,N_14886);
xnor UO_1344 (O_1344,N_14992,N_14607);
nor UO_1345 (O_1345,N_14808,N_14779);
nand UO_1346 (O_1346,N_14936,N_14711);
and UO_1347 (O_1347,N_14666,N_14693);
or UO_1348 (O_1348,N_14977,N_14691);
and UO_1349 (O_1349,N_14872,N_14998);
nor UO_1350 (O_1350,N_14541,N_14536);
xor UO_1351 (O_1351,N_14730,N_14975);
xnor UO_1352 (O_1352,N_14598,N_14749);
xor UO_1353 (O_1353,N_14954,N_14864);
nand UO_1354 (O_1354,N_14585,N_14867);
xnor UO_1355 (O_1355,N_14808,N_14557);
nand UO_1356 (O_1356,N_14656,N_14999);
or UO_1357 (O_1357,N_14800,N_14890);
nor UO_1358 (O_1358,N_14869,N_14853);
xnor UO_1359 (O_1359,N_14852,N_14738);
nor UO_1360 (O_1360,N_14765,N_14739);
or UO_1361 (O_1361,N_14552,N_14683);
nand UO_1362 (O_1362,N_14665,N_14703);
and UO_1363 (O_1363,N_14714,N_14790);
nand UO_1364 (O_1364,N_14850,N_14856);
or UO_1365 (O_1365,N_14589,N_14712);
and UO_1366 (O_1366,N_14936,N_14587);
xnor UO_1367 (O_1367,N_14898,N_14876);
xnor UO_1368 (O_1368,N_14725,N_14600);
nand UO_1369 (O_1369,N_14795,N_14864);
or UO_1370 (O_1370,N_14872,N_14759);
or UO_1371 (O_1371,N_14670,N_14678);
and UO_1372 (O_1372,N_14808,N_14952);
or UO_1373 (O_1373,N_14646,N_14906);
or UO_1374 (O_1374,N_14657,N_14947);
nand UO_1375 (O_1375,N_14621,N_14834);
or UO_1376 (O_1376,N_14953,N_14557);
nand UO_1377 (O_1377,N_14534,N_14638);
xor UO_1378 (O_1378,N_14784,N_14626);
nor UO_1379 (O_1379,N_14701,N_14639);
nor UO_1380 (O_1380,N_14861,N_14703);
xor UO_1381 (O_1381,N_14958,N_14882);
nand UO_1382 (O_1382,N_14921,N_14725);
nor UO_1383 (O_1383,N_14637,N_14890);
nand UO_1384 (O_1384,N_14938,N_14680);
xor UO_1385 (O_1385,N_14954,N_14894);
or UO_1386 (O_1386,N_14638,N_14699);
xnor UO_1387 (O_1387,N_14617,N_14637);
xor UO_1388 (O_1388,N_14573,N_14804);
or UO_1389 (O_1389,N_14793,N_14880);
nor UO_1390 (O_1390,N_14660,N_14898);
xnor UO_1391 (O_1391,N_14738,N_14541);
nor UO_1392 (O_1392,N_14694,N_14645);
and UO_1393 (O_1393,N_14742,N_14809);
xnor UO_1394 (O_1394,N_14806,N_14550);
nor UO_1395 (O_1395,N_14899,N_14641);
and UO_1396 (O_1396,N_14630,N_14995);
xnor UO_1397 (O_1397,N_14858,N_14680);
and UO_1398 (O_1398,N_14809,N_14501);
nand UO_1399 (O_1399,N_14757,N_14501);
nand UO_1400 (O_1400,N_14641,N_14982);
nor UO_1401 (O_1401,N_14789,N_14875);
or UO_1402 (O_1402,N_14607,N_14927);
xor UO_1403 (O_1403,N_14618,N_14896);
xor UO_1404 (O_1404,N_14767,N_14617);
or UO_1405 (O_1405,N_14936,N_14507);
and UO_1406 (O_1406,N_14764,N_14926);
nand UO_1407 (O_1407,N_14587,N_14897);
nand UO_1408 (O_1408,N_14766,N_14792);
nor UO_1409 (O_1409,N_14815,N_14563);
nor UO_1410 (O_1410,N_14503,N_14569);
and UO_1411 (O_1411,N_14729,N_14728);
or UO_1412 (O_1412,N_14716,N_14571);
and UO_1413 (O_1413,N_14563,N_14532);
and UO_1414 (O_1414,N_14565,N_14895);
nor UO_1415 (O_1415,N_14866,N_14862);
xnor UO_1416 (O_1416,N_14674,N_14576);
and UO_1417 (O_1417,N_14901,N_14504);
xor UO_1418 (O_1418,N_14758,N_14835);
nor UO_1419 (O_1419,N_14858,N_14592);
nor UO_1420 (O_1420,N_14661,N_14527);
xor UO_1421 (O_1421,N_14628,N_14717);
and UO_1422 (O_1422,N_14676,N_14949);
xnor UO_1423 (O_1423,N_14814,N_14884);
nor UO_1424 (O_1424,N_14701,N_14593);
xor UO_1425 (O_1425,N_14641,N_14881);
nor UO_1426 (O_1426,N_14915,N_14816);
nor UO_1427 (O_1427,N_14552,N_14831);
and UO_1428 (O_1428,N_14548,N_14553);
and UO_1429 (O_1429,N_14589,N_14770);
nor UO_1430 (O_1430,N_14905,N_14532);
nor UO_1431 (O_1431,N_14908,N_14743);
nor UO_1432 (O_1432,N_14909,N_14835);
nand UO_1433 (O_1433,N_14903,N_14848);
xor UO_1434 (O_1434,N_14823,N_14599);
or UO_1435 (O_1435,N_14828,N_14885);
nor UO_1436 (O_1436,N_14684,N_14621);
xnor UO_1437 (O_1437,N_14663,N_14616);
nand UO_1438 (O_1438,N_14700,N_14932);
nor UO_1439 (O_1439,N_14741,N_14947);
or UO_1440 (O_1440,N_14685,N_14579);
nand UO_1441 (O_1441,N_14839,N_14943);
nor UO_1442 (O_1442,N_14980,N_14651);
nor UO_1443 (O_1443,N_14801,N_14813);
nand UO_1444 (O_1444,N_14548,N_14510);
nor UO_1445 (O_1445,N_14811,N_14962);
nand UO_1446 (O_1446,N_14816,N_14645);
or UO_1447 (O_1447,N_14758,N_14920);
xnor UO_1448 (O_1448,N_14797,N_14881);
and UO_1449 (O_1449,N_14766,N_14775);
xnor UO_1450 (O_1450,N_14968,N_14659);
and UO_1451 (O_1451,N_14567,N_14766);
nor UO_1452 (O_1452,N_14766,N_14811);
xor UO_1453 (O_1453,N_14577,N_14521);
nor UO_1454 (O_1454,N_14733,N_14529);
nand UO_1455 (O_1455,N_14920,N_14736);
nand UO_1456 (O_1456,N_14804,N_14612);
xor UO_1457 (O_1457,N_14770,N_14807);
or UO_1458 (O_1458,N_14732,N_14534);
nor UO_1459 (O_1459,N_14565,N_14529);
nand UO_1460 (O_1460,N_14711,N_14956);
and UO_1461 (O_1461,N_14560,N_14518);
nand UO_1462 (O_1462,N_14698,N_14955);
and UO_1463 (O_1463,N_14871,N_14548);
or UO_1464 (O_1464,N_14537,N_14687);
xnor UO_1465 (O_1465,N_14957,N_14835);
xor UO_1466 (O_1466,N_14671,N_14648);
or UO_1467 (O_1467,N_14555,N_14754);
or UO_1468 (O_1468,N_14898,N_14554);
nor UO_1469 (O_1469,N_14766,N_14632);
and UO_1470 (O_1470,N_14759,N_14708);
and UO_1471 (O_1471,N_14639,N_14999);
or UO_1472 (O_1472,N_14902,N_14662);
and UO_1473 (O_1473,N_14858,N_14672);
nor UO_1474 (O_1474,N_14582,N_14901);
and UO_1475 (O_1475,N_14683,N_14555);
nand UO_1476 (O_1476,N_14616,N_14765);
nor UO_1477 (O_1477,N_14557,N_14822);
nand UO_1478 (O_1478,N_14584,N_14738);
xnor UO_1479 (O_1479,N_14823,N_14595);
xnor UO_1480 (O_1480,N_14820,N_14692);
or UO_1481 (O_1481,N_14606,N_14928);
or UO_1482 (O_1482,N_14515,N_14679);
nand UO_1483 (O_1483,N_14747,N_14956);
xnor UO_1484 (O_1484,N_14667,N_14976);
and UO_1485 (O_1485,N_14962,N_14554);
xor UO_1486 (O_1486,N_14954,N_14949);
xnor UO_1487 (O_1487,N_14626,N_14995);
xnor UO_1488 (O_1488,N_14713,N_14801);
or UO_1489 (O_1489,N_14649,N_14591);
nor UO_1490 (O_1490,N_14734,N_14975);
or UO_1491 (O_1491,N_14622,N_14693);
and UO_1492 (O_1492,N_14829,N_14750);
and UO_1493 (O_1493,N_14816,N_14862);
nor UO_1494 (O_1494,N_14637,N_14840);
or UO_1495 (O_1495,N_14622,N_14665);
or UO_1496 (O_1496,N_14770,N_14964);
nor UO_1497 (O_1497,N_14828,N_14554);
nor UO_1498 (O_1498,N_14815,N_14584);
nor UO_1499 (O_1499,N_14916,N_14949);
and UO_1500 (O_1500,N_14568,N_14907);
nand UO_1501 (O_1501,N_14515,N_14901);
nor UO_1502 (O_1502,N_14684,N_14662);
nand UO_1503 (O_1503,N_14739,N_14583);
nand UO_1504 (O_1504,N_14743,N_14522);
or UO_1505 (O_1505,N_14886,N_14626);
nor UO_1506 (O_1506,N_14982,N_14584);
xnor UO_1507 (O_1507,N_14967,N_14945);
nand UO_1508 (O_1508,N_14542,N_14722);
nand UO_1509 (O_1509,N_14555,N_14595);
nor UO_1510 (O_1510,N_14931,N_14549);
and UO_1511 (O_1511,N_14620,N_14735);
and UO_1512 (O_1512,N_14756,N_14663);
and UO_1513 (O_1513,N_14512,N_14795);
nor UO_1514 (O_1514,N_14806,N_14690);
or UO_1515 (O_1515,N_14848,N_14667);
and UO_1516 (O_1516,N_14674,N_14783);
and UO_1517 (O_1517,N_14730,N_14901);
nor UO_1518 (O_1518,N_14951,N_14705);
and UO_1519 (O_1519,N_14787,N_14929);
nor UO_1520 (O_1520,N_14851,N_14789);
nor UO_1521 (O_1521,N_14781,N_14805);
nor UO_1522 (O_1522,N_14527,N_14509);
nand UO_1523 (O_1523,N_14655,N_14947);
xnor UO_1524 (O_1524,N_14934,N_14729);
or UO_1525 (O_1525,N_14538,N_14937);
nand UO_1526 (O_1526,N_14686,N_14599);
nand UO_1527 (O_1527,N_14908,N_14662);
or UO_1528 (O_1528,N_14736,N_14637);
nor UO_1529 (O_1529,N_14617,N_14984);
and UO_1530 (O_1530,N_14947,N_14569);
or UO_1531 (O_1531,N_14706,N_14985);
xnor UO_1532 (O_1532,N_14605,N_14736);
and UO_1533 (O_1533,N_14874,N_14578);
xor UO_1534 (O_1534,N_14949,N_14982);
or UO_1535 (O_1535,N_14777,N_14910);
xnor UO_1536 (O_1536,N_14568,N_14562);
nor UO_1537 (O_1537,N_14978,N_14960);
nor UO_1538 (O_1538,N_14704,N_14503);
nand UO_1539 (O_1539,N_14847,N_14895);
and UO_1540 (O_1540,N_14669,N_14590);
xnor UO_1541 (O_1541,N_14794,N_14773);
nand UO_1542 (O_1542,N_14799,N_14748);
nor UO_1543 (O_1543,N_14632,N_14864);
nand UO_1544 (O_1544,N_14733,N_14952);
nor UO_1545 (O_1545,N_14541,N_14650);
and UO_1546 (O_1546,N_14944,N_14726);
or UO_1547 (O_1547,N_14932,N_14713);
or UO_1548 (O_1548,N_14843,N_14779);
nor UO_1549 (O_1549,N_14638,N_14855);
nand UO_1550 (O_1550,N_14838,N_14798);
nor UO_1551 (O_1551,N_14616,N_14746);
nor UO_1552 (O_1552,N_14935,N_14794);
xor UO_1553 (O_1553,N_14668,N_14849);
nor UO_1554 (O_1554,N_14607,N_14801);
xor UO_1555 (O_1555,N_14763,N_14802);
and UO_1556 (O_1556,N_14625,N_14750);
and UO_1557 (O_1557,N_14928,N_14557);
nor UO_1558 (O_1558,N_14552,N_14949);
nor UO_1559 (O_1559,N_14572,N_14981);
xor UO_1560 (O_1560,N_14630,N_14689);
xor UO_1561 (O_1561,N_14568,N_14777);
nor UO_1562 (O_1562,N_14669,N_14897);
xnor UO_1563 (O_1563,N_14919,N_14645);
nand UO_1564 (O_1564,N_14954,N_14975);
or UO_1565 (O_1565,N_14902,N_14829);
and UO_1566 (O_1566,N_14518,N_14758);
nand UO_1567 (O_1567,N_14562,N_14949);
nor UO_1568 (O_1568,N_14530,N_14842);
nor UO_1569 (O_1569,N_14964,N_14608);
nand UO_1570 (O_1570,N_14565,N_14688);
xnor UO_1571 (O_1571,N_14894,N_14831);
nand UO_1572 (O_1572,N_14725,N_14895);
or UO_1573 (O_1573,N_14654,N_14769);
xor UO_1574 (O_1574,N_14789,N_14815);
xnor UO_1575 (O_1575,N_14958,N_14723);
nor UO_1576 (O_1576,N_14509,N_14612);
nor UO_1577 (O_1577,N_14645,N_14807);
or UO_1578 (O_1578,N_14722,N_14665);
nand UO_1579 (O_1579,N_14517,N_14747);
nand UO_1580 (O_1580,N_14547,N_14816);
nor UO_1581 (O_1581,N_14660,N_14812);
and UO_1582 (O_1582,N_14736,N_14855);
xor UO_1583 (O_1583,N_14775,N_14770);
and UO_1584 (O_1584,N_14777,N_14853);
nand UO_1585 (O_1585,N_14763,N_14621);
nand UO_1586 (O_1586,N_14533,N_14789);
or UO_1587 (O_1587,N_14599,N_14661);
or UO_1588 (O_1588,N_14705,N_14788);
nand UO_1589 (O_1589,N_14948,N_14643);
nand UO_1590 (O_1590,N_14809,N_14549);
and UO_1591 (O_1591,N_14944,N_14556);
or UO_1592 (O_1592,N_14586,N_14618);
xnor UO_1593 (O_1593,N_14629,N_14575);
nand UO_1594 (O_1594,N_14707,N_14657);
nand UO_1595 (O_1595,N_14570,N_14926);
or UO_1596 (O_1596,N_14525,N_14536);
xor UO_1597 (O_1597,N_14713,N_14989);
xor UO_1598 (O_1598,N_14520,N_14953);
and UO_1599 (O_1599,N_14856,N_14602);
nor UO_1600 (O_1600,N_14671,N_14886);
and UO_1601 (O_1601,N_14610,N_14817);
and UO_1602 (O_1602,N_14850,N_14777);
or UO_1603 (O_1603,N_14868,N_14510);
xnor UO_1604 (O_1604,N_14781,N_14858);
or UO_1605 (O_1605,N_14885,N_14578);
nor UO_1606 (O_1606,N_14883,N_14636);
nor UO_1607 (O_1607,N_14708,N_14829);
nand UO_1608 (O_1608,N_14808,N_14505);
or UO_1609 (O_1609,N_14891,N_14830);
or UO_1610 (O_1610,N_14618,N_14512);
nand UO_1611 (O_1611,N_14516,N_14696);
nand UO_1612 (O_1612,N_14548,N_14543);
nand UO_1613 (O_1613,N_14509,N_14775);
nand UO_1614 (O_1614,N_14700,N_14951);
nand UO_1615 (O_1615,N_14991,N_14579);
or UO_1616 (O_1616,N_14556,N_14735);
nor UO_1617 (O_1617,N_14838,N_14638);
nand UO_1618 (O_1618,N_14692,N_14962);
nor UO_1619 (O_1619,N_14754,N_14815);
and UO_1620 (O_1620,N_14613,N_14744);
and UO_1621 (O_1621,N_14889,N_14820);
xnor UO_1622 (O_1622,N_14882,N_14678);
or UO_1623 (O_1623,N_14577,N_14657);
nor UO_1624 (O_1624,N_14659,N_14603);
or UO_1625 (O_1625,N_14869,N_14949);
or UO_1626 (O_1626,N_14523,N_14889);
and UO_1627 (O_1627,N_14637,N_14923);
or UO_1628 (O_1628,N_14718,N_14745);
nor UO_1629 (O_1629,N_14930,N_14675);
xor UO_1630 (O_1630,N_14532,N_14791);
and UO_1631 (O_1631,N_14856,N_14904);
nor UO_1632 (O_1632,N_14940,N_14558);
or UO_1633 (O_1633,N_14629,N_14505);
xor UO_1634 (O_1634,N_14993,N_14967);
xor UO_1635 (O_1635,N_14547,N_14529);
nand UO_1636 (O_1636,N_14987,N_14539);
nor UO_1637 (O_1637,N_14684,N_14513);
xnor UO_1638 (O_1638,N_14962,N_14584);
or UO_1639 (O_1639,N_14525,N_14763);
nor UO_1640 (O_1640,N_14751,N_14617);
nor UO_1641 (O_1641,N_14691,N_14885);
nor UO_1642 (O_1642,N_14951,N_14510);
nor UO_1643 (O_1643,N_14516,N_14661);
nand UO_1644 (O_1644,N_14911,N_14915);
and UO_1645 (O_1645,N_14626,N_14807);
xnor UO_1646 (O_1646,N_14868,N_14924);
xnor UO_1647 (O_1647,N_14972,N_14772);
and UO_1648 (O_1648,N_14525,N_14618);
xor UO_1649 (O_1649,N_14961,N_14557);
and UO_1650 (O_1650,N_14580,N_14794);
or UO_1651 (O_1651,N_14906,N_14924);
or UO_1652 (O_1652,N_14590,N_14867);
or UO_1653 (O_1653,N_14838,N_14657);
xor UO_1654 (O_1654,N_14793,N_14870);
nor UO_1655 (O_1655,N_14857,N_14783);
nor UO_1656 (O_1656,N_14949,N_14818);
nor UO_1657 (O_1657,N_14524,N_14907);
nand UO_1658 (O_1658,N_14845,N_14554);
and UO_1659 (O_1659,N_14733,N_14591);
xnor UO_1660 (O_1660,N_14838,N_14612);
xnor UO_1661 (O_1661,N_14697,N_14764);
xnor UO_1662 (O_1662,N_14719,N_14902);
or UO_1663 (O_1663,N_14612,N_14906);
nor UO_1664 (O_1664,N_14554,N_14741);
and UO_1665 (O_1665,N_14566,N_14766);
xnor UO_1666 (O_1666,N_14928,N_14665);
and UO_1667 (O_1667,N_14683,N_14546);
or UO_1668 (O_1668,N_14927,N_14544);
and UO_1669 (O_1669,N_14839,N_14771);
and UO_1670 (O_1670,N_14888,N_14726);
nand UO_1671 (O_1671,N_14964,N_14852);
or UO_1672 (O_1672,N_14513,N_14624);
and UO_1673 (O_1673,N_14586,N_14918);
or UO_1674 (O_1674,N_14667,N_14815);
nor UO_1675 (O_1675,N_14752,N_14875);
and UO_1676 (O_1676,N_14847,N_14765);
nand UO_1677 (O_1677,N_14850,N_14808);
nor UO_1678 (O_1678,N_14603,N_14546);
and UO_1679 (O_1679,N_14971,N_14912);
nand UO_1680 (O_1680,N_14779,N_14838);
nor UO_1681 (O_1681,N_14509,N_14790);
and UO_1682 (O_1682,N_14930,N_14911);
nand UO_1683 (O_1683,N_14795,N_14952);
nor UO_1684 (O_1684,N_14502,N_14909);
xor UO_1685 (O_1685,N_14501,N_14658);
or UO_1686 (O_1686,N_14726,N_14710);
nand UO_1687 (O_1687,N_14956,N_14830);
nor UO_1688 (O_1688,N_14691,N_14670);
nor UO_1689 (O_1689,N_14902,N_14643);
or UO_1690 (O_1690,N_14784,N_14532);
xor UO_1691 (O_1691,N_14748,N_14706);
xor UO_1692 (O_1692,N_14692,N_14886);
nor UO_1693 (O_1693,N_14771,N_14547);
nand UO_1694 (O_1694,N_14847,N_14802);
and UO_1695 (O_1695,N_14737,N_14573);
or UO_1696 (O_1696,N_14752,N_14924);
or UO_1697 (O_1697,N_14713,N_14667);
or UO_1698 (O_1698,N_14552,N_14844);
nor UO_1699 (O_1699,N_14776,N_14594);
and UO_1700 (O_1700,N_14630,N_14980);
xnor UO_1701 (O_1701,N_14910,N_14813);
nor UO_1702 (O_1702,N_14588,N_14861);
nand UO_1703 (O_1703,N_14808,N_14981);
xnor UO_1704 (O_1704,N_14826,N_14579);
xnor UO_1705 (O_1705,N_14787,N_14916);
or UO_1706 (O_1706,N_14522,N_14688);
nor UO_1707 (O_1707,N_14503,N_14886);
and UO_1708 (O_1708,N_14675,N_14539);
nor UO_1709 (O_1709,N_14559,N_14513);
or UO_1710 (O_1710,N_14725,N_14684);
and UO_1711 (O_1711,N_14820,N_14710);
or UO_1712 (O_1712,N_14608,N_14835);
nand UO_1713 (O_1713,N_14546,N_14968);
or UO_1714 (O_1714,N_14510,N_14527);
and UO_1715 (O_1715,N_14864,N_14750);
nand UO_1716 (O_1716,N_14666,N_14880);
and UO_1717 (O_1717,N_14984,N_14806);
nor UO_1718 (O_1718,N_14518,N_14989);
xnor UO_1719 (O_1719,N_14550,N_14921);
and UO_1720 (O_1720,N_14942,N_14877);
or UO_1721 (O_1721,N_14891,N_14558);
or UO_1722 (O_1722,N_14972,N_14711);
xor UO_1723 (O_1723,N_14805,N_14829);
xor UO_1724 (O_1724,N_14872,N_14681);
and UO_1725 (O_1725,N_14512,N_14955);
and UO_1726 (O_1726,N_14940,N_14605);
or UO_1727 (O_1727,N_14996,N_14977);
nor UO_1728 (O_1728,N_14861,N_14937);
nand UO_1729 (O_1729,N_14625,N_14660);
and UO_1730 (O_1730,N_14999,N_14515);
nand UO_1731 (O_1731,N_14533,N_14669);
and UO_1732 (O_1732,N_14975,N_14688);
nor UO_1733 (O_1733,N_14928,N_14877);
or UO_1734 (O_1734,N_14974,N_14627);
and UO_1735 (O_1735,N_14781,N_14620);
or UO_1736 (O_1736,N_14689,N_14805);
nand UO_1737 (O_1737,N_14876,N_14819);
nor UO_1738 (O_1738,N_14640,N_14901);
or UO_1739 (O_1739,N_14691,N_14936);
and UO_1740 (O_1740,N_14848,N_14526);
and UO_1741 (O_1741,N_14691,N_14843);
xnor UO_1742 (O_1742,N_14509,N_14743);
and UO_1743 (O_1743,N_14997,N_14546);
nor UO_1744 (O_1744,N_14858,N_14992);
and UO_1745 (O_1745,N_14725,N_14740);
or UO_1746 (O_1746,N_14838,N_14717);
nor UO_1747 (O_1747,N_14600,N_14564);
and UO_1748 (O_1748,N_14960,N_14641);
or UO_1749 (O_1749,N_14552,N_14529);
nand UO_1750 (O_1750,N_14907,N_14630);
xor UO_1751 (O_1751,N_14785,N_14603);
xnor UO_1752 (O_1752,N_14958,N_14894);
nand UO_1753 (O_1753,N_14691,N_14876);
and UO_1754 (O_1754,N_14523,N_14735);
and UO_1755 (O_1755,N_14842,N_14949);
and UO_1756 (O_1756,N_14593,N_14845);
nor UO_1757 (O_1757,N_14842,N_14809);
or UO_1758 (O_1758,N_14741,N_14888);
xnor UO_1759 (O_1759,N_14882,N_14597);
or UO_1760 (O_1760,N_14785,N_14621);
nand UO_1761 (O_1761,N_14784,N_14865);
nand UO_1762 (O_1762,N_14764,N_14551);
nor UO_1763 (O_1763,N_14555,N_14723);
nand UO_1764 (O_1764,N_14885,N_14681);
and UO_1765 (O_1765,N_14599,N_14528);
xnor UO_1766 (O_1766,N_14825,N_14769);
or UO_1767 (O_1767,N_14639,N_14643);
nor UO_1768 (O_1768,N_14928,N_14824);
and UO_1769 (O_1769,N_14806,N_14873);
xnor UO_1770 (O_1770,N_14546,N_14699);
or UO_1771 (O_1771,N_14503,N_14757);
xnor UO_1772 (O_1772,N_14602,N_14591);
and UO_1773 (O_1773,N_14519,N_14959);
and UO_1774 (O_1774,N_14874,N_14821);
xor UO_1775 (O_1775,N_14510,N_14627);
nand UO_1776 (O_1776,N_14682,N_14827);
or UO_1777 (O_1777,N_14895,N_14627);
nand UO_1778 (O_1778,N_14810,N_14524);
nand UO_1779 (O_1779,N_14996,N_14507);
or UO_1780 (O_1780,N_14750,N_14789);
nor UO_1781 (O_1781,N_14993,N_14595);
and UO_1782 (O_1782,N_14862,N_14621);
xor UO_1783 (O_1783,N_14607,N_14555);
nand UO_1784 (O_1784,N_14889,N_14959);
and UO_1785 (O_1785,N_14973,N_14744);
nand UO_1786 (O_1786,N_14848,N_14957);
and UO_1787 (O_1787,N_14741,N_14920);
and UO_1788 (O_1788,N_14826,N_14640);
or UO_1789 (O_1789,N_14893,N_14627);
nand UO_1790 (O_1790,N_14606,N_14579);
xnor UO_1791 (O_1791,N_14869,N_14858);
xnor UO_1792 (O_1792,N_14615,N_14773);
or UO_1793 (O_1793,N_14686,N_14593);
and UO_1794 (O_1794,N_14526,N_14523);
nand UO_1795 (O_1795,N_14685,N_14930);
and UO_1796 (O_1796,N_14732,N_14596);
or UO_1797 (O_1797,N_14915,N_14921);
nor UO_1798 (O_1798,N_14577,N_14892);
xnor UO_1799 (O_1799,N_14849,N_14613);
xor UO_1800 (O_1800,N_14728,N_14655);
nand UO_1801 (O_1801,N_14980,N_14993);
nor UO_1802 (O_1802,N_14981,N_14680);
xnor UO_1803 (O_1803,N_14682,N_14952);
and UO_1804 (O_1804,N_14856,N_14944);
and UO_1805 (O_1805,N_14875,N_14773);
nor UO_1806 (O_1806,N_14594,N_14566);
xor UO_1807 (O_1807,N_14980,N_14538);
and UO_1808 (O_1808,N_14988,N_14810);
nand UO_1809 (O_1809,N_14874,N_14924);
xor UO_1810 (O_1810,N_14591,N_14599);
nor UO_1811 (O_1811,N_14813,N_14705);
xor UO_1812 (O_1812,N_14696,N_14791);
nor UO_1813 (O_1813,N_14595,N_14588);
or UO_1814 (O_1814,N_14895,N_14573);
or UO_1815 (O_1815,N_14614,N_14604);
or UO_1816 (O_1816,N_14620,N_14831);
nand UO_1817 (O_1817,N_14501,N_14806);
nor UO_1818 (O_1818,N_14503,N_14581);
or UO_1819 (O_1819,N_14555,N_14875);
and UO_1820 (O_1820,N_14823,N_14907);
nor UO_1821 (O_1821,N_14639,N_14752);
or UO_1822 (O_1822,N_14774,N_14685);
xor UO_1823 (O_1823,N_14673,N_14658);
or UO_1824 (O_1824,N_14707,N_14774);
xor UO_1825 (O_1825,N_14768,N_14742);
nor UO_1826 (O_1826,N_14723,N_14980);
nand UO_1827 (O_1827,N_14569,N_14765);
xor UO_1828 (O_1828,N_14724,N_14684);
and UO_1829 (O_1829,N_14936,N_14650);
nor UO_1830 (O_1830,N_14501,N_14535);
nand UO_1831 (O_1831,N_14627,N_14979);
nor UO_1832 (O_1832,N_14815,N_14893);
xor UO_1833 (O_1833,N_14601,N_14866);
or UO_1834 (O_1834,N_14992,N_14973);
xor UO_1835 (O_1835,N_14688,N_14731);
or UO_1836 (O_1836,N_14645,N_14593);
or UO_1837 (O_1837,N_14543,N_14607);
or UO_1838 (O_1838,N_14831,N_14819);
or UO_1839 (O_1839,N_14848,N_14934);
xor UO_1840 (O_1840,N_14619,N_14754);
nand UO_1841 (O_1841,N_14730,N_14888);
and UO_1842 (O_1842,N_14828,N_14991);
nor UO_1843 (O_1843,N_14841,N_14899);
or UO_1844 (O_1844,N_14984,N_14700);
or UO_1845 (O_1845,N_14529,N_14985);
and UO_1846 (O_1846,N_14876,N_14705);
and UO_1847 (O_1847,N_14753,N_14538);
and UO_1848 (O_1848,N_14695,N_14892);
nor UO_1849 (O_1849,N_14653,N_14836);
or UO_1850 (O_1850,N_14659,N_14506);
nand UO_1851 (O_1851,N_14774,N_14984);
and UO_1852 (O_1852,N_14918,N_14853);
and UO_1853 (O_1853,N_14672,N_14524);
xnor UO_1854 (O_1854,N_14823,N_14989);
and UO_1855 (O_1855,N_14546,N_14595);
nand UO_1856 (O_1856,N_14939,N_14535);
xnor UO_1857 (O_1857,N_14526,N_14836);
nand UO_1858 (O_1858,N_14895,N_14921);
xor UO_1859 (O_1859,N_14526,N_14847);
xnor UO_1860 (O_1860,N_14574,N_14991);
nor UO_1861 (O_1861,N_14698,N_14914);
xor UO_1862 (O_1862,N_14925,N_14603);
and UO_1863 (O_1863,N_14701,N_14723);
nand UO_1864 (O_1864,N_14870,N_14788);
or UO_1865 (O_1865,N_14907,N_14754);
nand UO_1866 (O_1866,N_14973,N_14543);
nand UO_1867 (O_1867,N_14504,N_14701);
and UO_1868 (O_1868,N_14527,N_14960);
nor UO_1869 (O_1869,N_14782,N_14753);
or UO_1870 (O_1870,N_14999,N_14666);
nand UO_1871 (O_1871,N_14645,N_14780);
nor UO_1872 (O_1872,N_14974,N_14938);
nand UO_1873 (O_1873,N_14948,N_14532);
nand UO_1874 (O_1874,N_14882,N_14520);
and UO_1875 (O_1875,N_14896,N_14603);
nor UO_1876 (O_1876,N_14587,N_14541);
nor UO_1877 (O_1877,N_14607,N_14981);
nor UO_1878 (O_1878,N_14855,N_14591);
and UO_1879 (O_1879,N_14557,N_14980);
or UO_1880 (O_1880,N_14831,N_14972);
or UO_1881 (O_1881,N_14746,N_14740);
nor UO_1882 (O_1882,N_14566,N_14502);
nor UO_1883 (O_1883,N_14951,N_14875);
and UO_1884 (O_1884,N_14912,N_14581);
or UO_1885 (O_1885,N_14822,N_14941);
xor UO_1886 (O_1886,N_14897,N_14689);
nand UO_1887 (O_1887,N_14539,N_14883);
xor UO_1888 (O_1888,N_14536,N_14853);
xor UO_1889 (O_1889,N_14996,N_14531);
nor UO_1890 (O_1890,N_14837,N_14732);
xor UO_1891 (O_1891,N_14970,N_14723);
xor UO_1892 (O_1892,N_14571,N_14585);
and UO_1893 (O_1893,N_14710,N_14641);
nand UO_1894 (O_1894,N_14746,N_14980);
nand UO_1895 (O_1895,N_14736,N_14904);
and UO_1896 (O_1896,N_14864,N_14611);
nor UO_1897 (O_1897,N_14998,N_14766);
and UO_1898 (O_1898,N_14787,N_14869);
nand UO_1899 (O_1899,N_14579,N_14697);
nand UO_1900 (O_1900,N_14840,N_14918);
and UO_1901 (O_1901,N_14650,N_14556);
xnor UO_1902 (O_1902,N_14749,N_14905);
xor UO_1903 (O_1903,N_14501,N_14503);
nor UO_1904 (O_1904,N_14975,N_14508);
xor UO_1905 (O_1905,N_14891,N_14698);
nand UO_1906 (O_1906,N_14641,N_14650);
nor UO_1907 (O_1907,N_14644,N_14573);
nor UO_1908 (O_1908,N_14806,N_14666);
nand UO_1909 (O_1909,N_14825,N_14892);
or UO_1910 (O_1910,N_14600,N_14909);
and UO_1911 (O_1911,N_14767,N_14706);
or UO_1912 (O_1912,N_14709,N_14959);
nand UO_1913 (O_1913,N_14692,N_14642);
and UO_1914 (O_1914,N_14784,N_14614);
or UO_1915 (O_1915,N_14613,N_14687);
or UO_1916 (O_1916,N_14696,N_14730);
and UO_1917 (O_1917,N_14610,N_14785);
and UO_1918 (O_1918,N_14971,N_14827);
and UO_1919 (O_1919,N_14572,N_14687);
nand UO_1920 (O_1920,N_14910,N_14923);
nand UO_1921 (O_1921,N_14607,N_14846);
and UO_1922 (O_1922,N_14979,N_14736);
or UO_1923 (O_1923,N_14708,N_14780);
nor UO_1924 (O_1924,N_14601,N_14980);
and UO_1925 (O_1925,N_14666,N_14816);
nor UO_1926 (O_1926,N_14963,N_14802);
xnor UO_1927 (O_1927,N_14962,N_14933);
or UO_1928 (O_1928,N_14957,N_14510);
and UO_1929 (O_1929,N_14963,N_14835);
xor UO_1930 (O_1930,N_14858,N_14574);
and UO_1931 (O_1931,N_14539,N_14966);
xnor UO_1932 (O_1932,N_14899,N_14635);
nand UO_1933 (O_1933,N_14813,N_14990);
nor UO_1934 (O_1934,N_14807,N_14868);
nand UO_1935 (O_1935,N_14696,N_14615);
and UO_1936 (O_1936,N_14755,N_14681);
or UO_1937 (O_1937,N_14632,N_14792);
nand UO_1938 (O_1938,N_14522,N_14653);
nor UO_1939 (O_1939,N_14602,N_14928);
xor UO_1940 (O_1940,N_14813,N_14611);
and UO_1941 (O_1941,N_14784,N_14539);
nand UO_1942 (O_1942,N_14732,N_14716);
and UO_1943 (O_1943,N_14912,N_14521);
xnor UO_1944 (O_1944,N_14570,N_14789);
and UO_1945 (O_1945,N_14635,N_14816);
nand UO_1946 (O_1946,N_14538,N_14909);
nor UO_1947 (O_1947,N_14527,N_14889);
nor UO_1948 (O_1948,N_14951,N_14513);
or UO_1949 (O_1949,N_14684,N_14795);
and UO_1950 (O_1950,N_14657,N_14633);
nor UO_1951 (O_1951,N_14524,N_14760);
nor UO_1952 (O_1952,N_14542,N_14811);
or UO_1953 (O_1953,N_14747,N_14900);
nor UO_1954 (O_1954,N_14913,N_14552);
nor UO_1955 (O_1955,N_14884,N_14707);
and UO_1956 (O_1956,N_14800,N_14717);
or UO_1957 (O_1957,N_14913,N_14798);
xnor UO_1958 (O_1958,N_14764,N_14859);
nand UO_1959 (O_1959,N_14556,N_14949);
and UO_1960 (O_1960,N_14986,N_14957);
xor UO_1961 (O_1961,N_14888,N_14729);
nor UO_1962 (O_1962,N_14778,N_14921);
nor UO_1963 (O_1963,N_14960,N_14709);
and UO_1964 (O_1964,N_14786,N_14777);
xor UO_1965 (O_1965,N_14989,N_14905);
and UO_1966 (O_1966,N_14901,N_14965);
or UO_1967 (O_1967,N_14644,N_14506);
xor UO_1968 (O_1968,N_14688,N_14969);
or UO_1969 (O_1969,N_14836,N_14517);
xnor UO_1970 (O_1970,N_14867,N_14744);
nor UO_1971 (O_1971,N_14683,N_14996);
and UO_1972 (O_1972,N_14660,N_14896);
nand UO_1973 (O_1973,N_14990,N_14755);
nand UO_1974 (O_1974,N_14533,N_14831);
nor UO_1975 (O_1975,N_14710,N_14520);
or UO_1976 (O_1976,N_14557,N_14973);
or UO_1977 (O_1977,N_14520,N_14694);
nor UO_1978 (O_1978,N_14681,N_14812);
xnor UO_1979 (O_1979,N_14861,N_14716);
or UO_1980 (O_1980,N_14666,N_14853);
xor UO_1981 (O_1981,N_14803,N_14973);
or UO_1982 (O_1982,N_14818,N_14790);
xor UO_1983 (O_1983,N_14768,N_14613);
xor UO_1984 (O_1984,N_14729,N_14609);
nand UO_1985 (O_1985,N_14597,N_14768);
nor UO_1986 (O_1986,N_14810,N_14511);
nand UO_1987 (O_1987,N_14808,N_14673);
or UO_1988 (O_1988,N_14664,N_14502);
nor UO_1989 (O_1989,N_14925,N_14930);
and UO_1990 (O_1990,N_14768,N_14531);
and UO_1991 (O_1991,N_14926,N_14708);
or UO_1992 (O_1992,N_14581,N_14962);
nand UO_1993 (O_1993,N_14634,N_14538);
nor UO_1994 (O_1994,N_14631,N_14503);
or UO_1995 (O_1995,N_14738,N_14879);
nor UO_1996 (O_1996,N_14688,N_14933);
xor UO_1997 (O_1997,N_14750,N_14701);
nor UO_1998 (O_1998,N_14544,N_14581);
nor UO_1999 (O_1999,N_14854,N_14632);
endmodule