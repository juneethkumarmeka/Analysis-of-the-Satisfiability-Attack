module basic_2500_25000_3000_20_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_533,In_1104);
xnor U1 (N_1,In_1727,In_2150);
nor U2 (N_2,In_1566,In_891);
xor U3 (N_3,In_142,In_2182);
or U4 (N_4,In_1294,In_167);
or U5 (N_5,In_488,In_1484);
nand U6 (N_6,In_2280,In_408);
nand U7 (N_7,In_499,In_1542);
or U8 (N_8,In_2498,In_636);
or U9 (N_9,In_1924,In_2096);
and U10 (N_10,In_2416,In_1246);
and U11 (N_11,In_1631,In_725);
or U12 (N_12,In_157,In_972);
nand U13 (N_13,In_1930,In_539);
nor U14 (N_14,In_466,In_1298);
and U15 (N_15,In_1148,In_518);
nor U16 (N_16,In_1256,In_2375);
nor U17 (N_17,In_1705,In_2112);
xor U18 (N_18,In_591,In_17);
and U19 (N_19,In_1910,In_937);
xor U20 (N_20,In_1602,In_1624);
xnor U21 (N_21,In_2013,In_66);
or U22 (N_22,In_1545,In_2148);
xnor U23 (N_23,In_2025,In_387);
xor U24 (N_24,In_240,In_2170);
xnor U25 (N_25,In_267,In_847);
nor U26 (N_26,In_1702,In_2451);
nor U27 (N_27,In_337,In_2484);
or U28 (N_28,In_410,In_249);
nand U29 (N_29,In_1547,In_1959);
xor U30 (N_30,In_122,In_1058);
nor U31 (N_31,In_946,In_1604);
nand U32 (N_32,In_1319,In_346);
or U33 (N_33,In_852,In_182);
xnor U34 (N_34,In_123,In_81);
and U35 (N_35,In_357,In_631);
or U36 (N_36,In_1584,In_235);
nor U37 (N_37,In_1730,In_2360);
or U38 (N_38,In_1769,In_365);
xnor U39 (N_39,In_1474,In_1239);
or U40 (N_40,In_111,In_248);
nand U41 (N_41,In_130,In_2132);
or U42 (N_42,In_84,In_1462);
nor U43 (N_43,In_332,In_2259);
or U44 (N_44,In_40,In_1221);
or U45 (N_45,In_1270,In_379);
nor U46 (N_46,In_798,In_724);
and U47 (N_47,In_1044,In_2341);
or U48 (N_48,In_2100,In_2139);
nor U49 (N_49,In_1269,In_431);
nand U50 (N_50,In_2242,In_160);
nor U51 (N_51,In_817,In_1983);
or U52 (N_52,In_803,In_1353);
nand U53 (N_53,In_510,In_351);
nand U54 (N_54,In_386,In_1621);
and U55 (N_55,In_1312,In_392);
or U56 (N_56,In_1118,In_753);
nor U57 (N_57,In_2345,In_1367);
or U58 (N_58,In_2144,In_537);
xnor U59 (N_59,In_2351,In_287);
nor U60 (N_60,In_1211,In_158);
and U61 (N_61,In_630,In_1093);
and U62 (N_62,In_2338,In_1403);
nor U63 (N_63,In_1160,In_2142);
nand U64 (N_64,In_872,In_399);
nand U65 (N_65,In_1725,In_502);
nor U66 (N_66,In_1635,In_140);
or U67 (N_67,In_1075,In_336);
nor U68 (N_68,In_1709,In_1215);
nand U69 (N_69,In_599,In_886);
or U70 (N_70,In_1579,In_2414);
and U71 (N_71,In_1081,In_796);
or U72 (N_72,In_650,In_290);
xor U73 (N_73,In_821,In_1455);
nor U74 (N_74,In_1751,In_87);
or U75 (N_75,In_1811,In_535);
nor U76 (N_76,In_1210,In_137);
nand U77 (N_77,In_1176,In_2236);
nand U78 (N_78,In_480,In_1423);
or U79 (N_79,In_614,In_540);
xnor U80 (N_80,In_920,In_2077);
or U81 (N_81,In_1563,In_458);
xor U82 (N_82,In_2047,In_294);
xor U83 (N_83,In_475,In_320);
xor U84 (N_84,In_2174,In_1807);
or U85 (N_85,In_1236,In_1864);
nor U86 (N_86,In_1443,In_1140);
and U87 (N_87,In_2040,In_1204);
and U88 (N_88,In_1847,In_2364);
and U89 (N_89,In_1047,In_1684);
or U90 (N_90,In_1736,In_1516);
or U91 (N_91,In_1589,In_93);
nand U92 (N_92,In_2243,In_2283);
or U93 (N_93,In_1653,In_2021);
nand U94 (N_94,In_1626,In_613);
xor U95 (N_95,In_1080,In_401);
and U96 (N_96,In_1143,In_1171);
and U97 (N_97,In_104,In_1486);
nand U98 (N_98,In_1416,In_624);
or U99 (N_99,In_1981,In_1758);
or U100 (N_100,In_1759,In_2445);
nor U101 (N_101,In_1755,In_192);
nand U102 (N_102,In_923,In_51);
nor U103 (N_103,In_1855,In_1374);
nand U104 (N_104,In_1515,In_1955);
nand U105 (N_105,In_1170,In_1028);
nand U106 (N_106,In_1708,In_418);
and U107 (N_107,In_1921,In_1223);
nor U108 (N_108,In_1682,In_1741);
nor U109 (N_109,In_695,In_2463);
nor U110 (N_110,In_2442,In_702);
xor U111 (N_111,In_2298,In_571);
or U112 (N_112,In_378,In_2089);
or U113 (N_113,In_7,In_1393);
or U114 (N_114,In_2293,In_2116);
nand U115 (N_115,In_143,In_2322);
nand U116 (N_116,In_958,In_1217);
xnor U117 (N_117,In_355,In_637);
nor U118 (N_118,In_989,In_1922);
and U119 (N_119,In_1465,In_2146);
and U120 (N_120,In_921,In_1884);
nor U121 (N_121,In_445,In_2129);
and U122 (N_122,In_1501,In_203);
nand U123 (N_123,In_524,In_1259);
or U124 (N_124,In_327,In_1676);
or U125 (N_125,In_2367,In_164);
nor U126 (N_126,In_2453,In_666);
nor U127 (N_127,In_459,In_1664);
xnor U128 (N_128,In_1686,In_992);
and U129 (N_129,In_751,In_1477);
xor U130 (N_130,In_310,In_333);
xnor U131 (N_131,In_2181,In_574);
xnor U132 (N_132,In_1603,In_1527);
nor U133 (N_133,In_1805,In_1371);
nor U134 (N_134,In_1011,In_1095);
xor U135 (N_135,In_1562,In_1601);
nor U136 (N_136,In_397,In_2326);
or U137 (N_137,In_1905,In_2394);
or U138 (N_138,In_146,In_498);
nand U139 (N_139,In_1629,In_1514);
nand U140 (N_140,In_955,In_328);
or U141 (N_141,In_1136,In_2268);
xor U142 (N_142,In_1658,In_693);
and U143 (N_143,In_1744,In_126);
nor U144 (N_144,In_1345,In_727);
nor U145 (N_145,In_1105,In_1100);
xnor U146 (N_146,In_394,In_362);
nor U147 (N_147,In_1652,In_640);
nand U148 (N_148,In_764,In_211);
xor U149 (N_149,In_423,In_1793);
or U150 (N_150,In_712,In_256);
xor U151 (N_151,In_180,In_552);
xnor U152 (N_152,In_1703,In_1853);
and U153 (N_153,In_25,In_1231);
nor U154 (N_154,In_2410,In_471);
and U155 (N_155,In_760,In_348);
nor U156 (N_156,In_787,In_307);
and U157 (N_157,In_1690,In_1369);
nor U158 (N_158,In_2485,In_1972);
xnor U159 (N_159,In_1523,In_324);
or U160 (N_160,In_212,In_437);
xnor U161 (N_161,In_42,In_411);
or U162 (N_162,In_1588,In_846);
nand U163 (N_163,In_2130,In_2422);
nor U164 (N_164,In_2368,In_406);
xnor U165 (N_165,In_2255,In_1957);
nor U166 (N_166,In_2260,In_1863);
xor U167 (N_167,In_987,In_954);
and U168 (N_168,In_1533,In_1030);
or U169 (N_169,In_1732,In_1883);
nor U170 (N_170,In_276,In_1026);
nand U171 (N_171,In_1498,In_1599);
or U172 (N_172,In_2031,In_1908);
and U173 (N_173,In_482,In_67);
xnor U174 (N_174,In_2333,In_2330);
nand U175 (N_175,In_710,In_651);
and U176 (N_176,In_676,In_1489);
nor U177 (N_177,In_628,In_1814);
xnor U178 (N_178,In_2276,In_2003);
nor U179 (N_179,In_2063,In_2018);
and U180 (N_180,In_580,In_79);
and U181 (N_181,In_1000,In_795);
xor U182 (N_182,In_1344,In_762);
nand U183 (N_183,In_1934,In_2434);
or U184 (N_184,In_1913,In_1616);
xor U185 (N_185,In_80,In_49);
xor U186 (N_186,In_1822,In_1359);
or U187 (N_187,In_1154,In_1642);
xnor U188 (N_188,In_2210,In_117);
and U189 (N_189,In_1557,In_363);
nor U190 (N_190,In_2123,In_1409);
xnor U191 (N_191,In_858,In_136);
or U192 (N_192,In_546,In_1340);
nor U193 (N_193,In_2432,In_1130);
xor U194 (N_194,In_2402,In_1268);
and U195 (N_195,In_2151,In_1487);
nand U196 (N_196,In_1398,In_2014);
nor U197 (N_197,In_154,In_4);
xnor U198 (N_198,In_260,In_1321);
and U199 (N_199,In_658,In_739);
and U200 (N_200,In_263,In_1633);
and U201 (N_201,In_494,In_626);
nand U202 (N_202,In_1786,In_85);
nand U203 (N_203,In_1694,In_1421);
xnor U204 (N_204,In_1290,In_664);
nor U205 (N_205,In_1643,In_1045);
nor U206 (N_206,In_1912,In_129);
nor U207 (N_207,In_1789,In_2070);
xnor U208 (N_208,In_1201,In_220);
or U209 (N_209,In_912,In_2385);
nand U210 (N_210,In_1458,In_155);
xor U211 (N_211,In_152,In_2284);
or U212 (N_212,In_2152,In_1795);
xnor U213 (N_213,In_997,In_1552);
and U214 (N_214,In_696,In_2273);
xnor U215 (N_215,In_1561,In_1440);
xor U216 (N_216,In_334,In_934);
nor U217 (N_217,In_918,In_1647);
and U218 (N_218,In_1889,In_1228);
nand U219 (N_219,In_1018,In_807);
or U220 (N_220,In_1932,In_1005);
or U221 (N_221,In_31,In_2468);
nand U222 (N_222,In_2166,In_608);
nor U223 (N_223,In_1851,In_2302);
or U224 (N_224,In_1362,In_2353);
or U225 (N_225,In_1915,In_1608);
or U226 (N_226,In_2127,In_2030);
and U227 (N_227,In_1302,In_90);
or U228 (N_228,In_2004,In_2454);
and U229 (N_229,In_1405,In_1053);
or U230 (N_230,In_1222,In_1150);
nand U231 (N_231,In_2471,In_2167);
nor U232 (N_232,In_2172,In_715);
nand U233 (N_233,In_1146,In_1568);
or U234 (N_234,In_1098,In_2232);
or U235 (N_235,In_1370,In_1989);
xnor U236 (N_236,In_71,In_436);
xor U237 (N_237,In_655,In_1876);
and U238 (N_238,In_1802,In_1101);
xor U239 (N_239,In_930,In_1419);
nor U240 (N_240,In_472,In_1683);
nand U241 (N_241,In_906,In_1059);
or U242 (N_242,In_1559,In_16);
nand U243 (N_243,In_1771,In_456);
and U244 (N_244,In_1004,In_890);
xor U245 (N_245,In_2080,In_2493);
and U246 (N_246,In_2292,In_1351);
or U247 (N_247,In_2046,In_1435);
nand U248 (N_248,In_281,In_583);
nor U249 (N_249,In_848,In_1979);
or U250 (N_250,In_447,In_1110);
nor U251 (N_251,In_162,In_1008);
and U252 (N_252,In_1417,In_174);
nand U253 (N_253,In_828,In_2055);
xnor U254 (N_254,In_802,In_497);
xnor U255 (N_255,In_1704,In_2431);
and U256 (N_256,In_733,In_2008);
xor U257 (N_257,In_295,In_2264);
or U258 (N_258,In_366,In_1133);
nor U259 (N_259,In_582,In_103);
or U260 (N_260,In_780,In_2352);
nor U261 (N_261,In_550,In_2230);
nor U262 (N_262,In_2305,In_1580);
or U263 (N_263,In_519,In_672);
or U264 (N_264,In_959,In_1985);
xnor U265 (N_265,In_2262,In_1511);
and U266 (N_266,In_943,In_826);
nor U267 (N_267,In_549,In_1494);
nand U268 (N_268,In_1733,In_1636);
xor U269 (N_269,In_2479,In_325);
or U270 (N_270,In_46,In_931);
nand U271 (N_271,In_1281,In_24);
or U272 (N_272,In_2098,In_2193);
and U273 (N_273,In_1038,In_545);
or U274 (N_274,In_874,In_206);
or U275 (N_275,In_1036,In_329);
and U276 (N_276,In_187,In_1861);
and U277 (N_277,In_1195,In_496);
nand U278 (N_278,In_264,In_2488);
xor U279 (N_279,In_711,In_1818);
nand U280 (N_280,In_1166,In_1391);
nor U281 (N_281,In_889,In_2334);
or U282 (N_282,In_981,In_2299);
and U283 (N_283,In_1640,In_1969);
nor U284 (N_284,In_1743,In_1890);
and U285 (N_285,In_314,In_928);
nand U286 (N_286,In_1900,In_1078);
and U287 (N_287,In_309,In_88);
xor U288 (N_288,In_561,In_2002);
and U289 (N_289,In_426,In_1243);
or U290 (N_290,In_1114,In_302);
nor U291 (N_291,In_1848,In_1249);
or U292 (N_292,In_2245,In_1939);
nor U293 (N_293,In_1503,In_195);
nand U294 (N_294,In_2229,In_1257);
nor U295 (N_295,In_177,In_347);
or U296 (N_296,In_1179,In_230);
xnor U297 (N_297,In_1553,In_633);
xnor U298 (N_298,In_428,In_1206);
and U299 (N_299,In_1801,In_862);
nor U300 (N_300,In_300,In_107);
or U301 (N_301,In_272,In_2147);
nand U302 (N_302,In_1227,In_790);
or U303 (N_303,In_885,In_1212);
xnor U304 (N_304,In_2094,In_2117);
and U305 (N_305,In_2121,In_770);
or U306 (N_306,In_1071,In_38);
and U307 (N_307,In_1885,In_116);
nand U308 (N_308,In_812,In_217);
nor U309 (N_309,In_1792,In_576);
xnor U310 (N_310,In_442,In_288);
and U311 (N_311,In_1657,In_1823);
nand U312 (N_312,In_1950,In_1685);
nand U313 (N_313,In_377,In_367);
or U314 (N_314,In_1615,In_1549);
nand U315 (N_315,In_2071,In_2291);
xor U316 (N_316,In_1596,In_2029);
or U317 (N_317,In_94,In_2389);
and U318 (N_318,In_880,In_19);
xnor U319 (N_319,In_823,In_2306);
nor U320 (N_320,In_898,In_2495);
or U321 (N_321,In_1035,In_771);
or U322 (N_322,In_686,In_568);
or U323 (N_323,In_1672,In_2176);
and U324 (N_324,In_784,In_448);
nor U325 (N_325,In_528,In_1606);
nor U326 (N_326,In_1010,In_1209);
and U327 (N_327,In_1893,In_1062);
and U328 (N_328,In_1783,In_1055);
and U329 (N_329,In_1200,In_793);
nor U330 (N_330,In_139,In_2424);
nor U331 (N_331,In_2449,In_596);
or U332 (N_332,In_629,In_2043);
or U333 (N_333,In_2024,In_1582);
or U334 (N_334,In_781,In_134);
nor U335 (N_335,In_1128,In_1190);
nor U336 (N_336,In_1453,In_689);
or U337 (N_337,In_274,In_200);
and U338 (N_338,In_1701,In_926);
nand U339 (N_339,In_598,In_1627);
or U340 (N_340,In_2266,In_1479);
or U341 (N_341,In_1226,In_503);
nand U342 (N_342,In_1232,In_1536);
or U343 (N_343,In_2392,In_800);
and U344 (N_344,In_2443,In_2192);
or U345 (N_345,In_477,In_1264);
or U346 (N_346,In_2061,In_945);
nor U347 (N_347,In_967,In_1949);
nand U348 (N_348,In_1082,In_2459);
nor U349 (N_349,In_936,In_1841);
nor U350 (N_350,In_1571,In_1696);
nand U351 (N_351,In_1216,In_2277);
and U352 (N_352,In_2057,In_214);
nand U353 (N_353,In_2418,In_32);
or U354 (N_354,In_383,In_173);
and U355 (N_355,In_1926,In_1670);
and U356 (N_356,In_2331,In_1408);
nor U357 (N_357,In_2474,In_1187);
nor U358 (N_358,In_1585,In_2374);
and U359 (N_359,In_2278,In_515);
nand U360 (N_360,In_638,In_161);
and U361 (N_361,In_856,In_973);
nand U362 (N_362,In_1669,In_754);
nand U363 (N_363,In_1528,In_64);
nand U364 (N_364,In_1966,In_1174);
or U365 (N_365,In_1534,In_1272);
xnor U366 (N_366,In_1878,In_313);
nor U367 (N_367,In_404,In_701);
nor U368 (N_368,In_1961,In_506);
and U369 (N_369,In_1454,In_1001);
xor U370 (N_370,In_2241,In_529);
and U371 (N_371,In_1158,In_2175);
xnor U372 (N_372,In_572,In_884);
xnor U373 (N_373,In_395,In_646);
or U374 (N_374,In_649,In_1806);
xor U375 (N_375,In_900,In_102);
nand U376 (N_376,In_2068,In_2083);
or U377 (N_377,In_1574,In_857);
nand U378 (N_378,In_1329,In_609);
and U379 (N_379,In_755,In_1051);
nand U380 (N_380,In_2058,In_1444);
xor U381 (N_381,In_556,In_625);
xor U382 (N_382,In_1695,In_1586);
nand U383 (N_383,In_1073,In_2075);
or U384 (N_384,In_1247,In_1466);
nand U385 (N_385,In_635,In_2337);
or U386 (N_386,In_1338,In_1524);
and U387 (N_387,In_2009,In_1188);
nand U388 (N_388,In_748,In_2188);
nand U389 (N_389,In_601,In_151);
nand U390 (N_390,In_2282,In_2436);
nand U391 (N_391,In_2135,In_1102);
and U392 (N_392,In_2109,In_184);
xnor U393 (N_393,In_1833,In_425);
nand U394 (N_394,In_2473,In_373);
nor U395 (N_395,In_1826,In_2189);
nand U396 (N_396,In_961,In_2234);
or U397 (N_397,In_1379,In_809);
or U398 (N_398,In_1161,In_2203);
nor U399 (N_399,In_836,In_1040);
and U400 (N_400,In_2218,In_417);
nor U401 (N_401,In_1872,In_2177);
nor U402 (N_402,In_368,In_209);
and U403 (N_403,In_283,In_1343);
and U404 (N_404,In_2339,In_1901);
nor U405 (N_405,In_1753,In_1325);
nor U406 (N_406,In_1844,In_196);
nor U407 (N_407,In_279,In_1012);
nand U408 (N_408,In_132,In_839);
nor U409 (N_409,In_1526,In_2274);
or U410 (N_410,In_1084,In_2373);
nor U411 (N_411,In_2289,In_834);
nand U412 (N_412,In_841,In_1825);
and U413 (N_413,In_743,In_684);
nand U414 (N_414,In_665,In_1386);
xnor U415 (N_415,In_259,In_2154);
nand U416 (N_416,In_1927,In_709);
or U417 (N_417,In_949,In_1903);
xnor U418 (N_418,In_1845,In_2126);
nand U419 (N_419,In_1992,In_602);
nand U420 (N_420,In_1986,In_1407);
and U421 (N_421,In_674,In_866);
nor U422 (N_422,In_424,In_745);
nor U423 (N_423,In_1315,In_1618);
or U424 (N_424,In_618,In_271);
nor U425 (N_425,In_23,In_1718);
nand U426 (N_426,In_2252,In_851);
and U427 (N_427,In_306,In_2429);
nand U428 (N_428,In_963,In_2461);
nor U429 (N_429,In_100,In_1681);
and U430 (N_430,In_737,In_1737);
nand U431 (N_431,In_312,In_1230);
nand U432 (N_432,In_1337,In_1021);
or U433 (N_433,In_1275,In_1445);
xnor U434 (N_434,In_278,In_2141);
nand U435 (N_435,In_1063,In_639);
or U436 (N_436,In_2050,In_777);
xor U437 (N_437,In_2324,In_1997);
and U438 (N_438,In_1122,In_1317);
and U439 (N_439,In_2173,In_258);
nand U440 (N_440,In_354,In_863);
or U441 (N_441,In_2012,In_340);
nand U442 (N_442,In_1581,In_2197);
and U443 (N_443,In_2206,In_893);
or U444 (N_444,In_1491,In_2329);
or U445 (N_445,In_1303,In_621);
nor U446 (N_446,In_1242,In_1224);
nand U447 (N_447,In_1429,In_2240);
and U448 (N_448,In_2244,In_1687);
xnor U449 (N_449,In_1518,In_776);
or U450 (N_450,In_229,In_1335);
nand U451 (N_451,In_1813,In_2048);
and U452 (N_452,In_1892,In_1787);
and U453 (N_453,In_1775,In_2270);
nor U454 (N_454,In_1998,In_204);
or U455 (N_455,In_469,In_1381);
or U456 (N_456,In_2476,In_219);
nor U457 (N_457,In_1425,In_1354);
or U458 (N_458,In_186,In_1456);
or U459 (N_459,In_2209,In_1331);
nor U460 (N_460,In_1449,In_1418);
and U461 (N_461,In_1020,In_1460);
nand U462 (N_462,In_0,In_956);
nand U463 (N_463,In_763,In_1790);
or U464 (N_464,In_382,In_1506);
or U465 (N_465,In_76,In_59);
nand U466 (N_466,In_994,In_297);
and U467 (N_467,In_251,In_1570);
xnor U468 (N_468,In_323,In_1830);
nor U469 (N_469,In_570,In_453);
nor U470 (N_470,In_2257,In_1594);
or U471 (N_471,In_718,In_2428);
and U472 (N_472,In_1390,In_2311);
nor U473 (N_473,In_688,In_1923);
and U474 (N_474,In_564,In_1244);
or U475 (N_475,In_343,In_1121);
or U476 (N_476,In_993,In_1087);
or U477 (N_477,In_716,In_542);
or U478 (N_478,In_2489,In_349);
and U479 (N_479,In_1346,In_1540);
or U480 (N_480,In_1609,In_361);
or U481 (N_481,In_486,In_83);
nand U482 (N_482,In_2064,In_474);
and U483 (N_483,In_603,In_791);
or U484 (N_484,In_818,In_1459);
nand U485 (N_485,In_653,In_2478);
nor U486 (N_486,In_704,In_2145);
nor U487 (N_487,In_223,In_2225);
or U488 (N_488,In_792,In_869);
xnor U489 (N_489,In_590,In_1816);
and U490 (N_490,In_413,In_1083);
and U491 (N_491,In_2059,In_2386);
or U492 (N_492,In_1638,In_96);
and U493 (N_493,In_119,In_756);
nor U494 (N_494,In_1740,In_789);
nor U495 (N_495,In_252,In_13);
and U496 (N_496,In_2470,In_1954);
xnor U497 (N_497,In_284,In_878);
and U498 (N_498,In_648,In_1819);
xor U499 (N_499,In_2134,In_2433);
xnor U500 (N_500,In_319,In_2408);
and U501 (N_501,In_1043,In_2221);
nand U502 (N_502,In_282,In_855);
and U503 (N_503,In_2361,In_507);
nor U504 (N_504,In_1079,In_2288);
xor U505 (N_505,In_671,In_1287);
xor U506 (N_506,In_2001,In_2107);
xnor U507 (N_507,In_1309,In_2336);
nor U508 (N_508,In_159,In_1134);
nor U509 (N_509,In_730,In_2212);
or U510 (N_510,In_1904,In_45);
nand U511 (N_511,In_765,In_1144);
nand U512 (N_512,In_1550,In_2155);
and U513 (N_513,In_1410,In_1070);
nand U514 (N_514,In_516,In_478);
nor U515 (N_515,In_1630,In_72);
or U516 (N_516,In_657,In_1569);
nor U517 (N_517,In_1333,In_619);
or U518 (N_518,In_1760,In_1551);
and U519 (N_519,In_97,In_275);
nor U520 (N_520,In_2310,In_2222);
nor U521 (N_521,In_476,In_1575);
xor U522 (N_522,In_2399,In_534);
and U523 (N_523,In_1448,In_353);
or U524 (N_524,In_1318,In_1308);
nand U525 (N_525,In_298,In_1809);
xor U526 (N_526,In_2359,In_1229);
nor U527 (N_527,In_202,In_911);
and U528 (N_528,In_1015,In_1473);
nand U529 (N_529,In_1761,In_2137);
nand U530 (N_530,In_708,In_1304);
and U531 (N_531,In_1541,In_543);
nor U532 (N_532,In_77,In_190);
xnor U533 (N_533,In_2054,In_1361);
nand U534 (N_534,In_1866,In_2462);
and U535 (N_535,In_1781,In_1131);
xnor U536 (N_536,In_916,In_1086);
nor U537 (N_537,In_2251,In_450);
and U538 (N_538,In_1027,In_1578);
nand U539 (N_539,In_1746,In_1091);
xor U540 (N_540,In_1591,In_2017);
xnor U541 (N_541,In_172,In_683);
or U542 (N_542,In_738,In_396);
and U543 (N_543,In_1914,In_1875);
nand U544 (N_544,In_432,In_138);
nor U545 (N_545,In_1933,In_409);
or U546 (N_546,In_389,In_1538);
and U547 (N_547,In_1387,In_2099);
or U548 (N_548,In_371,In_1646);
and U549 (N_549,In_822,In_415);
xnor U550 (N_550,In_1049,In_1024);
nand U551 (N_551,In_243,In_47);
xnor U552 (N_552,In_227,In_2427);
or U553 (N_553,In_289,In_1472);
and U554 (N_554,In_2430,In_1330);
and U555 (N_555,In_115,In_509);
or U556 (N_556,In_2185,In_786);
and U557 (N_557,In_178,In_109);
nand U558 (N_558,In_1238,In_669);
nand U559 (N_559,In_726,In_1597);
and U560 (N_560,In_1186,In_1525);
nand U561 (N_561,In_145,In_2285);
nand U562 (N_562,In_1659,In_225);
or U563 (N_563,In_1415,In_1461);
and U564 (N_564,In_412,In_1770);
xnor U565 (N_565,In_2049,In_2149);
nor U566 (N_566,In_1724,In_322);
and U567 (N_567,In_2342,In_1797);
or U568 (N_568,In_897,In_1858);
nand U569 (N_569,In_1156,In_1654);
and U570 (N_570,In_2475,In_335);
nor U571 (N_571,In_73,In_2184);
xnor U572 (N_572,In_2477,In_407);
and U573 (N_573,In_460,In_581);
nand U574 (N_574,In_226,In_1567);
or U575 (N_575,In_623,In_1163);
xor U576 (N_576,In_2104,In_679);
nand U577 (N_577,In_1607,In_1535);
or U578 (N_578,In_2235,In_797);
xor U579 (N_579,In_1798,In_1432);
nor U580 (N_580,In_1613,In_2267);
and U581 (N_581,In_2456,In_1810);
nand U582 (N_582,In_2387,In_370);
and U583 (N_583,In_1990,In_2204);
and U584 (N_584,In_2231,In_384);
and U585 (N_585,In_1019,In_1007);
nor U586 (N_586,In_1510,In_68);
xnor U587 (N_587,In_430,In_33);
or U588 (N_588,In_2390,In_662);
nand U589 (N_589,In_929,In_1292);
and U590 (N_590,In_680,In_641);
nor U591 (N_591,In_1911,In_1931);
nand U592 (N_592,In_673,In_1225);
and U593 (N_593,In_1852,In_1155);
or U594 (N_594,In_350,In_767);
nand U595 (N_595,In_586,In_364);
nand U596 (N_596,In_1328,In_1189);
nand U597 (N_597,In_565,In_984);
and U598 (N_598,In_2092,In_2319);
or U599 (N_599,In_1572,In_2346);
nor U600 (N_600,In_14,In_758);
and U601 (N_601,In_1671,In_1031);
xnor U602 (N_602,In_1284,In_1064);
nand U603 (N_603,In_18,In_827);
xor U604 (N_604,In_69,In_113);
or U605 (N_605,In_2397,In_2340);
nand U606 (N_606,In_2090,In_953);
xor U607 (N_607,In_15,In_1879);
xnor U608 (N_608,In_1977,In_2483);
or U609 (N_609,In_2465,In_1288);
or U610 (N_610,In_1859,In_1700);
and U611 (N_611,In_1117,In_1832);
nor U612 (N_612,In_1963,In_805);
and U613 (N_613,In_2419,In_1180);
or U614 (N_614,In_439,In_1940);
nor U615 (N_615,In_1003,In_947);
nor U616 (N_616,In_1721,In_2404);
nand U617 (N_617,In_1363,In_270);
and U618 (N_618,In_2269,In_1617);
or U619 (N_619,In_1973,In_1067);
xnor U620 (N_620,In_311,In_687);
xor U621 (N_621,In_1947,In_722);
and U622 (N_622,In_1632,In_1902);
nand U623 (N_623,In_359,In_1610);
or U624 (N_624,In_919,In_2258);
nand U625 (N_625,In_741,In_1368);
xnor U626 (N_626,In_2085,In_838);
or U627 (N_627,In_1512,In_1764);
or U628 (N_628,In_1214,In_1862);
and U629 (N_629,In_1896,In_971);
nand U630 (N_630,In_1723,In_2247);
nor U631 (N_631,In_1441,In_1348);
nand U632 (N_632,In_419,In_1948);
xor U633 (N_633,In_1280,In_20);
and U634 (N_634,In_241,In_62);
xor U635 (N_635,In_1245,In_1050);
nor U636 (N_636,In_464,In_1248);
nor U637 (N_637,In_1785,In_654);
nor U638 (N_638,In_966,In_1276);
xnor U639 (N_639,In_808,In_1906);
or U640 (N_640,In_1530,In_558);
nand U641 (N_641,In_224,In_1728);
and U642 (N_642,In_1305,In_2163);
xnor U643 (N_643,In_850,In_1048);
and U644 (N_644,In_393,In_2220);
nand U645 (N_645,In_165,In_483);
or U646 (N_646,In_1483,In_1509);
nor U647 (N_647,In_668,In_1220);
xnor U648 (N_648,In_2316,In_2391);
nand U649 (N_649,In_1522,In_1277);
xnor U650 (N_650,In_1447,In_2108);
nand U651 (N_651,In_2393,In_750);
xnor U652 (N_652,In_594,In_1895);
and U653 (N_653,In_321,In_816);
nor U654 (N_654,In_1697,In_421);
xor U655 (N_655,In_1099,In_1469);
or U656 (N_656,In_2406,In_479);
xor U657 (N_657,In_532,In_617);
nand U658 (N_658,In_1046,In_2301);
nand U659 (N_659,In_1316,In_1411);
nand U660 (N_660,In_1749,In_27);
nor U661 (N_661,In_1628,In_1693);
or U662 (N_662,In_887,In_1661);
or U663 (N_663,In_1267,In_55);
xor U664 (N_664,In_2438,In_1888);
or U665 (N_665,In_400,In_567);
xor U666 (N_666,In_1870,In_1314);
nor U667 (N_667,In_2015,In_179);
or U668 (N_668,In_2224,In_1945);
xor U669 (N_669,In_925,In_1714);
or U670 (N_670,In_1074,In_1784);
nor U671 (N_671,In_1513,In_685);
xor U672 (N_672,In_1820,In_914);
nor U673 (N_673,In_541,In_1964);
xnor U674 (N_674,In_388,In_1634);
or U675 (N_675,In_1076,In_1402);
nand U676 (N_676,In_2320,In_273);
nor U677 (N_677,In_292,In_1762);
xnor U678 (N_678,In_232,In_553);
nor U679 (N_679,In_2120,In_2412);
or U680 (N_680,In_2178,In_1378);
and U681 (N_681,In_1835,In_691);
nand U682 (N_682,In_57,In_490);
or U683 (N_683,In_1181,In_1554);
and U684 (N_684,In_2314,In_1752);
nand U685 (N_685,In_1068,In_175);
xor U686 (N_686,In_978,In_163);
or U687 (N_687,In_1857,In_1241);
nor U688 (N_688,In_2328,In_927);
and U689 (N_689,In_1377,In_1177);
nand U690 (N_690,In_766,In_1975);
or U691 (N_691,In_1558,In_1120);
or U692 (N_692,In_199,In_489);
nand U693 (N_693,In_1300,In_1587);
nand U694 (N_694,In_1467,In_845);
nand U695 (N_695,In_414,In_615);
nand U696 (N_696,In_2111,In_589);
nor U697 (N_697,In_2395,In_1843);
nor U698 (N_698,In_1625,In_1323);
and U699 (N_699,In_1556,In_1840);
nand U700 (N_700,In_344,In_888);
nor U701 (N_701,In_222,In_2296);
nand U702 (N_702,In_990,In_940);
or U703 (N_703,In_849,In_438);
nor U704 (N_704,In_369,In_1984);
xnor U705 (N_705,In_1165,In_2213);
nand U706 (N_706,In_607,In_2403);
nor U707 (N_707,In_699,In_1941);
or U708 (N_708,In_2202,In_326);
nor U709 (N_709,In_2226,In_2069);
nand U710 (N_710,In_156,In_2290);
nand U711 (N_711,In_530,In_1774);
xnor U712 (N_712,In_1828,In_2409);
xnor U713 (N_713,In_1766,In_1173);
nand U714 (N_714,In_30,In_305);
or U715 (N_715,In_938,In_434);
nor U716 (N_716,In_1349,In_2119);
or U717 (N_717,In_1713,In_385);
xor U718 (N_718,In_1495,In_2300);
xnor U719 (N_719,In_463,In_2307);
xnor U720 (N_720,In_1392,In_330);
or U721 (N_721,In_1937,In_1650);
xor U722 (N_722,In_2191,In_1291);
xor U723 (N_723,In_707,In_2081);
or U724 (N_724,In_2180,In_2481);
or U725 (N_725,In_1492,In_2153);
xnor U726 (N_726,In_1129,In_1772);
and U727 (N_727,In_2073,In_634);
and U728 (N_728,In_1202,In_147);
nor U729 (N_729,In_2091,In_286);
nor U730 (N_730,In_1768,In_1089);
nand U731 (N_731,In_1311,In_2211);
nor U732 (N_732,In_1665,In_237);
nor U733 (N_733,In_864,In_1255);
nor U734 (N_734,In_52,In_2464);
or U735 (N_735,In_1235,In_902);
xor U736 (N_736,In_1262,In_98);
and U737 (N_737,In_2467,In_218);
nand U738 (N_738,In_1982,In_1175);
xnor U739 (N_739,In_1052,In_1897);
nand U740 (N_740,In_2347,In_1698);
or U741 (N_741,In_723,In_493);
or U742 (N_742,In_1164,In_1936);
nand U743 (N_743,In_2196,In_446);
nand U744 (N_744,In_269,In_573);
and U745 (N_745,In_1873,In_1006);
xnor U746 (N_746,In_2286,In_969);
nor U747 (N_747,In_1821,In_1951);
or U748 (N_748,In_566,In_2039);
or U749 (N_749,In_1250,In_1108);
nor U750 (N_750,In_774,In_2158);
nand U751 (N_751,In_720,In_905);
or U752 (N_752,In_127,In_939);
or U753 (N_753,In_2309,In_647);
and U754 (N_754,In_1735,In_48);
and U755 (N_755,In_2169,In_892);
xor U756 (N_756,In_663,In_1138);
nor U757 (N_757,In_1598,In_1508);
or U758 (N_758,In_1831,In_462);
nor U759 (N_759,In_1942,In_2253);
xor U760 (N_760,In_1037,In_2143);
or U761 (N_761,In_717,In_198);
nand U762 (N_762,In_1794,In_820);
xnor U763 (N_763,In_587,In_114);
xor U764 (N_764,In_2125,In_1935);
or U765 (N_765,In_962,In_837);
nor U766 (N_766,In_694,In_1689);
or U767 (N_767,In_714,In_2281);
nand U768 (N_768,In_1874,In_909);
or U769 (N_769,In_1077,In_2469);
and U770 (N_770,In_244,In_37);
nand U771 (N_771,In_2378,In_75);
nand U772 (N_772,In_868,In_391);
and U773 (N_773,In_39,In_1573);
xor U774 (N_774,In_882,In_2214);
nand U775 (N_775,In_454,In_2448);
or U776 (N_776,In_968,In_2370);
xnor U777 (N_777,In_2401,In_1266);
nand U778 (N_778,In_830,In_538);
xor U779 (N_779,In_308,In_736);
nor U780 (N_780,In_1017,In_2079);
or U781 (N_781,In_1109,In_1978);
nand U782 (N_782,In_22,In_1521);
and U783 (N_783,In_1438,In_995);
or U784 (N_784,In_877,In_1142);
or U785 (N_785,In_2275,In_2363);
xor U786 (N_786,In_620,In_2303);
nand U787 (N_787,In_1260,In_2425);
nand U788 (N_788,In_876,In_1388);
xor U789 (N_789,In_2053,In_728);
and U790 (N_790,In_2016,In_1750);
nor U791 (N_791,In_112,In_1364);
nand U792 (N_792,In_593,In_1824);
nand U793 (N_793,In_933,In_1497);
nand U794 (N_794,In_2384,In_121);
or U795 (N_795,In_692,In_78);
nand U796 (N_796,In_843,In_131);
xnor U797 (N_797,In_1152,In_1116);
xor U798 (N_798,In_2381,In_1699);
and U799 (N_799,In_894,In_2056);
or U800 (N_800,In_1960,In_713);
nand U801 (N_801,In_952,In_908);
and U802 (N_802,In_95,In_1198);
and U803 (N_803,In_1780,In_2327);
nor U804 (N_804,In_871,In_128);
nor U805 (N_805,In_597,In_1734);
nand U806 (N_806,In_523,In_2207);
and U807 (N_807,In_2238,In_5);
nand U808 (N_808,In_216,In_1777);
nand U809 (N_809,In_183,In_2097);
xnor U810 (N_810,In_2388,In_2084);
nor U811 (N_811,In_1422,In_170);
or U812 (N_812,In_491,In_652);
or U813 (N_813,In_508,In_285);
xor U814 (N_814,In_470,In_1137);
and U815 (N_815,In_468,In_61);
or U816 (N_816,In_682,In_1803);
and U817 (N_817,In_2028,In_1191);
nand U818 (N_818,In_1065,In_1088);
xor U819 (N_819,In_1372,In_124);
and U820 (N_820,In_2323,In_2205);
nand U821 (N_821,In_907,In_513);
xor U822 (N_822,In_1720,In_390);
xnor U823 (N_823,In_560,In_578);
nor U824 (N_824,In_2183,In_761);
nand U825 (N_825,In_1944,In_2246);
or U826 (N_826,In_536,In_191);
or U827 (N_827,In_1149,In_1039);
or U828 (N_828,In_525,In_1014);
nand U829 (N_829,In_1167,In_873);
nor U830 (N_830,In_2161,In_86);
and U831 (N_831,In_1756,In_988);
and U832 (N_832,In_120,In_1507);
xor U833 (N_833,In_957,In_2208);
xor U834 (N_834,In_356,In_2321);
nor U835 (N_835,In_2105,In_2195);
xor U836 (N_836,In_1135,In_2227);
nor U837 (N_837,In_233,In_1692);
xor U838 (N_838,In_2441,In_835);
or U839 (N_839,In_65,In_1278);
nor U840 (N_840,In_108,In_1196);
nand U841 (N_841,In_375,In_193);
nand U842 (N_842,In_2254,In_1357);
nor U843 (N_843,In_1434,In_1739);
nand U844 (N_844,In_1299,In_1988);
and U845 (N_845,In_1178,In_1871);
xor U846 (N_846,In_667,In_2366);
xor U847 (N_847,In_242,In_1499);
nor U848 (N_848,In_12,In_991);
and U849 (N_849,In_1427,In_1193);
nand U850 (N_850,In_2038,In_606);
and U851 (N_851,In_1426,In_801);
nor U852 (N_852,In_2032,In_950);
xor U853 (N_853,In_1622,In_1748);
or U854 (N_854,In_1757,In_2466);
nand U855 (N_855,In_746,In_41);
nand U856 (N_856,In_2450,In_1504);
and U857 (N_857,In_910,In_1974);
nor U858 (N_858,In_1745,In_1576);
xnor U859 (N_859,In_360,In_2115);
and U860 (N_860,In_819,In_1747);
nand U861 (N_861,In_2164,In_2162);
xor U862 (N_862,In_2128,In_1856);
or U863 (N_863,In_304,In_1965);
or U864 (N_864,In_831,In_1342);
nand U865 (N_865,In_799,In_1404);
nand U866 (N_866,In_1869,In_1502);
nand U867 (N_867,In_2332,In_1849);
or U868 (N_868,In_440,In_681);
nand U869 (N_869,In_246,In_2140);
xnor U870 (N_870,In_1928,In_1327);
nand U871 (N_871,In_1085,In_236);
and U872 (N_872,In_2187,In_1383);
and U873 (N_873,In_405,In_303);
nand U874 (N_874,In_1836,In_2405);
or U875 (N_875,In_457,In_99);
xor U876 (N_876,In_1867,In_1157);
nor U877 (N_877,In_1297,In_1715);
nand U878 (N_878,In_1123,In_2490);
nand U879 (N_879,In_1919,In_1396);
xor U880 (N_880,In_1115,In_2343);
xnor U881 (N_881,In_904,In_1976);
and U882 (N_882,In_1375,In_296);
or U883 (N_883,In_1400,In_257);
nand U884 (N_884,In_44,In_1069);
and U885 (N_885,In_2355,In_2497);
xor U886 (N_886,In_1590,In_1194);
and U887 (N_887,In_2398,In_1717);
and U888 (N_888,In_1560,In_951);
nand U889 (N_889,In_1072,In_1482);
and U890 (N_890,In_149,In_2261);
or U891 (N_891,In_527,In_171);
nor U892 (N_892,In_974,In_1263);
and U893 (N_893,In_1399,In_1898);
xnor U894 (N_894,In_778,In_2074);
nand U895 (N_895,In_207,In_1439);
xnor U896 (N_896,In_1295,In_221);
nor U897 (N_897,In_1145,In_1132);
and U898 (N_898,In_1980,In_2369);
or U899 (N_899,In_2000,In_1564);
nand U900 (N_900,In_705,In_213);
nor U901 (N_901,In_1234,In_1127);
and U902 (N_902,In_2492,In_1711);
nand U903 (N_903,In_43,In_1779);
nand U904 (N_904,In_901,In_1022);
and U905 (N_905,In_579,In_985);
nor U906 (N_906,In_2067,In_1754);
or U907 (N_907,In_35,In_1147);
and U908 (N_908,In_2455,In_1943);
and U909 (N_909,In_1996,In_2440);
nor U910 (N_910,In_1320,In_575);
and U911 (N_911,In_2042,In_208);
nor U912 (N_912,In_1918,In_2294);
and U913 (N_913,In_2060,In_1706);
or U914 (N_914,In_840,In_2052);
and U915 (N_915,In_1970,In_632);
nor U916 (N_916,In_6,In_584);
nand U917 (N_917,In_2365,In_481);
and U918 (N_918,In_125,In_1218);
or U919 (N_919,In_2200,In_444);
and U920 (N_920,In_2124,In_520);
nor U921 (N_921,In_1493,In_2297);
xnor U922 (N_922,In_2356,In_2095);
xor U923 (N_923,In_1162,In_2011);
nand U924 (N_924,In_2423,In_2199);
nand U925 (N_925,In_106,In_1731);
and U926 (N_926,In_1663,In_1962);
nand U927 (N_927,In_1707,In_1029);
nand U928 (N_928,In_2439,In_36);
nor U929 (N_929,In_2110,In_899);
and U930 (N_930,In_2035,In_2007);
and U931 (N_931,In_698,In_1324);
xor U932 (N_932,In_1286,In_1054);
and U933 (N_933,In_2437,In_2382);
and U934 (N_934,In_1016,In_1475);
and U935 (N_935,In_2377,In_1356);
nand U936 (N_936,In_975,In_376);
xor U937 (N_937,In_473,In_1450);
xor U938 (N_938,In_484,In_1691);
or U939 (N_939,In_1648,In_105);
and U940 (N_940,In_2411,In_58);
nand U941 (N_941,In_2421,In_979);
nand U942 (N_942,In_600,In_1837);
xnor U943 (N_943,In_1623,In_2239);
or U944 (N_944,In_526,In_1301);
nor U945 (N_945,In_547,In_1987);
nor U946 (N_946,In_814,In_783);
xnor U947 (N_947,In_522,In_2034);
nor U948 (N_948,In_757,In_2179);
or U949 (N_949,In_2354,In_1850);
and U950 (N_950,In_1742,In_239);
and U951 (N_951,In_467,In_1066);
and U952 (N_952,In_1656,In_1668);
nor U953 (N_953,In_1373,In_338);
and U954 (N_954,In_443,In_779);
nand U955 (N_955,In_1113,In_1555);
or U956 (N_956,In_1139,In_1956);
and U957 (N_957,In_1360,In_675);
nor U958 (N_958,In_895,In_2250);
and U959 (N_959,In_875,In_74);
nor U960 (N_960,In_2102,In_517);
nand U961 (N_961,In_531,In_2044);
nor U962 (N_962,In_1182,In_1023);
nor U963 (N_963,In_2133,In_1865);
nor U964 (N_964,In_341,In_563);
nand U965 (N_965,In_1679,In_2114);
nor U966 (N_966,In_1313,In_1842);
nor U967 (N_967,In_2156,In_1090);
and U968 (N_968,In_1395,In_1808);
nor U969 (N_969,In_1891,In_291);
and U970 (N_970,In_1834,In_1452);
or U971 (N_971,In_1394,In_2426);
xor U972 (N_972,In_1829,In_1860);
nor U973 (N_973,In_2396,In_2217);
nand U974 (N_974,In_2315,In_2248);
or U975 (N_975,In_1184,In_261);
nor U976 (N_976,In_1677,In_1251);
or U977 (N_977,In_948,In_1358);
nor U978 (N_978,In_1172,In_1310);
nor U979 (N_979,In_1350,In_1882);
or U980 (N_980,In_56,In_588);
xnor U981 (N_981,In_998,In_1094);
or U982 (N_982,In_815,In_1496);
nand U983 (N_983,In_1476,In_2078);
xor U984 (N_984,In_996,In_1605);
nand U985 (N_985,In_1002,In_512);
nand U986 (N_986,In_452,In_1612);
and U987 (N_987,In_1880,In_1726);
xor U988 (N_988,In_1197,In_1107);
or U989 (N_989,In_26,In_1666);
nor U990 (N_990,In_1032,In_833);
and U991 (N_991,In_2216,In_1619);
xnor U992 (N_992,In_759,In_1778);
nand U993 (N_993,In_965,In_1791);
xnor U994 (N_994,In_861,In_1651);
nand U995 (N_995,In_433,In_794);
nor U996 (N_996,In_659,In_133);
or U997 (N_997,In_1096,In_2223);
xor U998 (N_998,In_293,In_917);
or U999 (N_999,In_611,In_228);
nor U1000 (N_1000,In_729,In_2019);
nor U1001 (N_1001,In_210,In_1994);
nand U1002 (N_1002,In_1366,In_644);
nor U1003 (N_1003,In_53,In_2460);
nand U1004 (N_1004,In_1365,In_2190);
or U1005 (N_1005,In_555,In_238);
nor U1006 (N_1006,In_1520,In_1060);
or U1007 (N_1007,In_747,In_101);
nand U1008 (N_1008,In_2312,In_832);
xor U1009 (N_1009,In_372,In_3);
or U1010 (N_1010,In_782,In_2086);
nor U1011 (N_1011,In_1219,In_181);
nand U1012 (N_1012,In_592,In_339);
nor U1013 (N_1013,In_1213,In_1253);
xnor U1014 (N_1014,In_2357,In_2271);
or U1015 (N_1015,In_700,In_661);
or U1016 (N_1016,In_2041,In_92);
nand U1017 (N_1017,In_2472,In_1352);
xnor U1018 (N_1018,In_935,In_185);
nor U1019 (N_1019,In_189,In_870);
nand U1020 (N_1020,In_342,In_1886);
xnor U1021 (N_1021,In_1347,In_1995);
and U1022 (N_1022,In_2304,In_941);
nand U1023 (N_1023,In_865,In_2027);
xnor U1024 (N_1024,In_1776,In_604);
nand U1025 (N_1025,In_1655,In_1273);
xor U1026 (N_1026,In_1042,In_2088);
or U1027 (N_1027,In_1125,In_2171);
or U1028 (N_1028,In_2308,In_1710);
xnor U1029 (N_1029,In_595,In_1056);
nor U1030 (N_1030,In_2349,In_1887);
xor U1031 (N_1031,In_153,In_1112);
nand U1032 (N_1032,In_514,In_1952);
xnor U1033 (N_1033,In_932,In_485);
nor U1034 (N_1034,In_944,In_1967);
or U1035 (N_1035,In_903,In_970);
xnor U1036 (N_1036,In_769,In_1376);
nand U1037 (N_1037,In_403,In_234);
nor U1038 (N_1038,In_2458,In_501);
or U1039 (N_1039,In_749,In_511);
and U1040 (N_1040,In_416,In_2113);
or U1041 (N_1041,In_1649,In_1827);
and U1042 (N_1042,In_559,In_2033);
xor U1043 (N_1043,In_1485,In_804);
and U1044 (N_1044,In_678,In_610);
or U1045 (N_1045,In_1442,In_605);
nand U1046 (N_1046,In_2023,In_1306);
and U1047 (N_1047,In_1839,In_1738);
and U1048 (N_1048,In_1674,In_245);
or U1049 (N_1049,In_980,In_1641);
or U1050 (N_1050,In_1282,In_266);
and U1051 (N_1051,In_1620,In_703);
and U1052 (N_1052,In_10,In_2020);
nand U1053 (N_1053,In_21,In_1252);
nand U1054 (N_1054,In_2496,In_1773);
or U1055 (N_1055,In_231,In_616);
and U1056 (N_1056,In_2413,In_642);
and U1057 (N_1057,In_150,In_168);
nand U1058 (N_1058,In_656,In_1183);
xor U1059 (N_1059,In_1208,In_420);
nor U1060 (N_1060,In_960,In_1611);
or U1061 (N_1061,In_1397,In_1595);
nor U1062 (N_1062,In_1159,In_881);
xnor U1063 (N_1063,In_82,In_1614);
or U1064 (N_1064,In_1688,In_2380);
nor U1065 (N_1065,In_544,In_982);
and U1066 (N_1066,In_2372,In_194);
nand U1067 (N_1067,In_1205,In_976);
nor U1068 (N_1068,In_331,In_1401);
nor U1069 (N_1069,In_141,In_1920);
nand U1070 (N_1070,In_1126,In_1544);
and U1071 (N_1071,In_2219,In_2400);
or U1072 (N_1072,In_2317,In_2228);
nand U1073 (N_1073,In_670,In_677);
xor U1074 (N_1074,In_1437,In_562);
xor U1075 (N_1075,In_735,In_1639);
and U1076 (N_1076,In_2237,In_2006);
xnor U1077 (N_1077,In_697,In_744);
or U1078 (N_1078,In_1667,In_719);
and U1079 (N_1079,In_422,In_318);
or U1080 (N_1080,In_317,In_2376);
xnor U1081 (N_1081,In_250,In_913);
and U1082 (N_1082,In_461,In_2233);
nand U1083 (N_1083,In_1468,In_2435);
nor U1084 (N_1084,In_1712,In_2103);
xnor U1085 (N_1085,In_896,In_1274);
xor U1086 (N_1086,In_1380,In_1583);
xor U1087 (N_1087,In_2325,In_1406);
xor U1088 (N_1088,In_2072,In_70);
and U1089 (N_1089,In_2215,In_734);
and U1090 (N_1090,In_89,In_9);
or U1091 (N_1091,In_2486,In_1763);
nor U1092 (N_1092,In_1413,In_1953);
xnor U1093 (N_1093,In_1788,In_50);
or U1094 (N_1094,In_34,In_254);
or U1095 (N_1095,In_2022,In_1531);
nand U1096 (N_1096,In_1041,In_201);
or U1097 (N_1097,In_1854,In_643);
or U1098 (N_1098,In_2082,In_1804);
nor U1099 (N_1099,In_1480,In_986);
or U1100 (N_1100,In_1326,In_548);
xor U1101 (N_1101,In_1868,In_569);
xor U1102 (N_1102,In_1464,In_924);
nor U1103 (N_1103,In_768,In_2452);
or U1104 (N_1104,In_1767,In_1457);
and U1105 (N_1105,In_1296,In_627);
nand U1106 (N_1106,In_451,In_188);
nand U1107 (N_1107,In_1,In_1917);
nand U1108 (N_1108,In_1168,In_2313);
nor U1109 (N_1109,In_1675,In_1103);
xor U1110 (N_1110,In_1546,In_721);
nand U1111 (N_1111,In_551,In_1938);
and U1112 (N_1112,In_1192,In_2062);
nor U1113 (N_1113,In_1999,In_1812);
nor U1114 (N_1114,In_775,In_1637);
xnor U1115 (N_1115,In_742,In_2165);
nor U1116 (N_1116,In_829,In_1106);
nand U1117 (N_1117,In_1446,In_1237);
nor U1118 (N_1118,In_148,In_1800);
nand U1119 (N_1119,In_1505,In_1033);
or U1120 (N_1120,In_2344,In_1644);
nand U1121 (N_1121,In_1341,In_557);
nor U1122 (N_1122,In_1899,In_1532);
and U1123 (N_1123,In_1153,In_1169);
and U1124 (N_1124,In_879,In_1548);
xor U1125 (N_1125,In_1968,In_2065);
nor U1126 (N_1126,In_1385,In_1389);
or U1127 (N_1127,In_1013,In_500);
and U1128 (N_1128,In_842,In_1355);
or U1129 (N_1129,In_752,In_441);
or U1130 (N_1130,In_380,In_29);
nor U1131 (N_1131,In_1307,In_2362);
nor U1132 (N_1132,In_2106,In_2420);
and U1133 (N_1133,In_999,In_1817);
nand U1134 (N_1134,In_1565,In_860);
nor U1135 (N_1135,In_1185,In_301);
and U1136 (N_1136,In_465,In_455);
and U1137 (N_1137,In_922,In_1111);
nor U1138 (N_1138,In_1796,In_1592);
and U1139 (N_1139,In_773,In_853);
nor U1140 (N_1140,In_2194,In_1470);
and U1141 (N_1141,In_1529,In_1971);
nand U1142 (N_1142,In_435,In_1414);
nor U1143 (N_1143,In_1765,In_402);
xor U1144 (N_1144,In_1141,In_2093);
or U1145 (N_1145,In_2010,In_2482);
and U1146 (N_1146,In_1488,In_1838);
or U1147 (N_1147,In_381,In_824);
xnor U1148 (N_1148,In_1261,In_2383);
xnor U1149 (N_1149,In_977,In_2066);
or U1150 (N_1150,In_1334,In_622);
and U1151 (N_1151,In_315,In_1424);
nor U1152 (N_1152,In_1240,In_110);
or U1153 (N_1153,In_2494,In_915);
or U1154 (N_1154,In_2407,In_1471);
or U1155 (N_1155,In_983,In_60);
nor U1156 (N_1156,In_1673,In_1600);
or U1157 (N_1157,In_1500,In_2447);
and U1158 (N_1158,In_2350,In_2160);
nand U1159 (N_1159,In_487,In_2087);
and U1160 (N_1160,In_1846,In_1199);
xor U1161 (N_1161,In_1339,In_2272);
nand U1162 (N_1162,In_2,In_2263);
and U1163 (N_1163,In_1907,In_1057);
and U1164 (N_1164,In_1293,In_2026);
nand U1165 (N_1165,In_1382,In_374);
nor U1166 (N_1166,In_299,In_1025);
or U1167 (N_1167,In_505,In_867);
or U1168 (N_1168,In_2256,In_645);
nand U1169 (N_1169,In_1384,In_1660);
nor U1170 (N_1170,In_2168,In_1097);
and U1171 (N_1171,In_1061,In_429);
xnor U1172 (N_1172,In_1929,In_135);
nor U1173 (N_1173,In_1537,In_1431);
xor U1174 (N_1174,In_54,In_813);
or U1175 (N_1175,In_1894,In_197);
or U1176 (N_1176,In_883,In_1420);
xor U1177 (N_1177,In_1124,In_854);
nor U1178 (N_1178,In_859,In_1430);
nand U1179 (N_1179,In_2287,In_1034);
xor U1180 (N_1180,In_577,In_1254);
nor U1181 (N_1181,In_1279,In_1662);
and U1182 (N_1182,In_964,In_398);
nand U1183 (N_1183,In_91,In_1925);
or U1184 (N_1184,In_1119,In_352);
nand U1185 (N_1185,In_215,In_2379);
nor U1186 (N_1186,In_504,In_492);
xnor U1187 (N_1187,In_2186,In_1916);
and U1188 (N_1188,In_1151,In_2157);
nor U1189 (N_1189,In_1877,In_2045);
nand U1190 (N_1190,In_2491,In_806);
nand U1191 (N_1191,In_1332,In_2138);
nor U1192 (N_1192,In_2265,In_11);
and U1193 (N_1193,In_942,In_2005);
and U1194 (N_1194,In_785,In_1283);
nand U1195 (N_1195,In_1678,In_345);
and U1196 (N_1196,In_255,In_740);
or U1197 (N_1197,In_772,In_316);
and U1198 (N_1198,In_825,In_2159);
or U1199 (N_1199,In_1463,In_554);
nor U1200 (N_1200,In_280,In_1451);
nand U1201 (N_1201,In_2487,In_1543);
nand U1202 (N_1202,In_1412,In_690);
nand U1203 (N_1203,In_1645,In_2201);
and U1204 (N_1204,In_1881,In_277);
nand U1205 (N_1205,In_2348,In_521);
nor U1206 (N_1206,In_1729,In_1782);
nor U1207 (N_1207,In_1336,In_28);
xnor U1208 (N_1208,In_358,In_2371);
or U1209 (N_1209,In_788,In_706);
nor U1210 (N_1210,In_176,In_1539);
nor U1211 (N_1211,In_2076,In_1322);
and U1212 (N_1212,In_1436,In_2499);
or U1213 (N_1213,In_732,In_1719);
nand U1214 (N_1214,In_1991,In_1433);
and U1215 (N_1215,In_118,In_1481);
xor U1216 (N_1216,In_144,In_1233);
and U1217 (N_1217,In_449,In_1265);
nand U1218 (N_1218,In_1258,In_2457);
or U1219 (N_1219,In_2131,In_731);
nor U1220 (N_1220,In_1958,In_810);
xor U1221 (N_1221,In_2198,In_262);
nand U1222 (N_1222,In_1289,In_1478);
xnor U1223 (N_1223,In_1203,In_1593);
nor U1224 (N_1224,In_2051,In_169);
and U1225 (N_1225,In_1519,In_2118);
xor U1226 (N_1226,In_265,In_8);
nor U1227 (N_1227,In_2295,In_2446);
nor U1228 (N_1228,In_660,In_1716);
or U1229 (N_1229,In_1577,In_247);
nand U1230 (N_1230,In_1271,In_585);
and U1231 (N_1231,In_612,In_2444);
nor U1232 (N_1232,In_2136,In_1946);
and U1233 (N_1233,In_2122,In_1993);
nand U1234 (N_1234,In_2101,In_2037);
and U1235 (N_1235,In_2318,In_1909);
and U1236 (N_1236,In_844,In_1815);
xor U1237 (N_1237,In_205,In_1722);
nor U1238 (N_1238,In_1799,In_2036);
or U1239 (N_1239,In_268,In_2480);
xnor U1240 (N_1240,In_166,In_1428);
nand U1241 (N_1241,In_1092,In_2415);
or U1242 (N_1242,In_1207,In_495);
or U1243 (N_1243,In_2335,In_1680);
xnor U1244 (N_1244,In_427,In_2358);
nand U1245 (N_1245,In_2417,In_1517);
and U1246 (N_1246,In_2249,In_2279);
and U1247 (N_1247,In_253,In_811);
and U1248 (N_1248,In_1009,In_1490);
or U1249 (N_1249,In_63,In_1285);
and U1250 (N_1250,N_1205,N_437);
nor U1251 (N_1251,N_961,N_746);
nand U1252 (N_1252,N_9,N_979);
nor U1253 (N_1253,N_1130,N_419);
or U1254 (N_1254,N_233,N_1056);
nor U1255 (N_1255,N_433,N_498);
nand U1256 (N_1256,N_1210,N_813);
nand U1257 (N_1257,N_1088,N_1231);
xor U1258 (N_1258,N_1036,N_497);
or U1259 (N_1259,N_416,N_246);
nand U1260 (N_1260,N_271,N_1246);
and U1261 (N_1261,N_431,N_819);
xor U1262 (N_1262,N_1183,N_729);
and U1263 (N_1263,N_4,N_863);
nand U1264 (N_1264,N_412,N_275);
or U1265 (N_1265,N_581,N_1010);
and U1266 (N_1266,N_678,N_1204);
or U1267 (N_1267,N_1075,N_22);
nand U1268 (N_1268,N_1209,N_1012);
or U1269 (N_1269,N_35,N_90);
nor U1270 (N_1270,N_1192,N_993);
nor U1271 (N_1271,N_707,N_81);
nor U1272 (N_1272,N_260,N_761);
or U1273 (N_1273,N_231,N_239);
and U1274 (N_1274,N_633,N_719);
xnor U1275 (N_1275,N_135,N_641);
nor U1276 (N_1276,N_331,N_1069);
nand U1277 (N_1277,N_446,N_709);
or U1278 (N_1278,N_285,N_65);
xnor U1279 (N_1279,N_824,N_623);
xor U1280 (N_1280,N_1170,N_388);
nor U1281 (N_1281,N_1050,N_512);
nor U1282 (N_1282,N_775,N_831);
nand U1283 (N_1283,N_1175,N_31);
nand U1284 (N_1284,N_1113,N_1188);
nor U1285 (N_1285,N_844,N_413);
nand U1286 (N_1286,N_747,N_1054);
or U1287 (N_1287,N_537,N_434);
xor U1288 (N_1288,N_71,N_877);
or U1289 (N_1289,N_915,N_874);
or U1290 (N_1290,N_934,N_749);
or U1291 (N_1291,N_26,N_1234);
xor U1292 (N_1292,N_272,N_911);
and U1293 (N_1293,N_460,N_181);
or U1294 (N_1294,N_987,N_888);
or U1295 (N_1295,N_514,N_1092);
xnor U1296 (N_1296,N_1208,N_1080);
nand U1297 (N_1297,N_1212,N_525);
nor U1298 (N_1298,N_868,N_938);
xnor U1299 (N_1299,N_475,N_209);
nor U1300 (N_1300,N_311,N_38);
or U1301 (N_1301,N_882,N_715);
xor U1302 (N_1302,N_607,N_1112);
xnor U1303 (N_1303,N_16,N_745);
nand U1304 (N_1304,N_338,N_590);
or U1305 (N_1305,N_1,N_287);
nand U1306 (N_1306,N_1070,N_50);
or U1307 (N_1307,N_929,N_593);
nand U1308 (N_1308,N_935,N_658);
nor U1309 (N_1309,N_494,N_1040);
and U1310 (N_1310,N_300,N_20);
xor U1311 (N_1311,N_695,N_1177);
and U1312 (N_1312,N_278,N_118);
or U1313 (N_1313,N_774,N_472);
nand U1314 (N_1314,N_1206,N_1129);
nand U1315 (N_1315,N_1226,N_1245);
nor U1316 (N_1316,N_381,N_335);
or U1317 (N_1317,N_741,N_146);
or U1318 (N_1318,N_1082,N_1064);
and U1319 (N_1319,N_845,N_1158);
nor U1320 (N_1320,N_664,N_196);
nor U1321 (N_1321,N_722,N_559);
xnor U1322 (N_1322,N_1094,N_937);
or U1323 (N_1323,N_564,N_145);
nor U1324 (N_1324,N_718,N_941);
xor U1325 (N_1325,N_711,N_814);
xor U1326 (N_1326,N_679,N_931);
and U1327 (N_1327,N_1227,N_109);
and U1328 (N_1328,N_227,N_454);
and U1329 (N_1329,N_1216,N_313);
and U1330 (N_1330,N_265,N_171);
or U1331 (N_1331,N_716,N_691);
and U1332 (N_1332,N_792,N_1184);
nor U1333 (N_1333,N_49,N_925);
and U1334 (N_1334,N_574,N_465);
nor U1335 (N_1335,N_557,N_111);
or U1336 (N_1336,N_452,N_640);
or U1337 (N_1337,N_996,N_158);
xor U1338 (N_1338,N_1048,N_856);
xnor U1339 (N_1339,N_482,N_293);
nor U1340 (N_1340,N_500,N_87);
nor U1341 (N_1341,N_1148,N_83);
and U1342 (N_1342,N_45,N_624);
or U1343 (N_1343,N_767,N_126);
xnor U1344 (N_1344,N_1098,N_632);
nor U1345 (N_1345,N_392,N_1156);
nor U1346 (N_1346,N_933,N_781);
xor U1347 (N_1347,N_1190,N_427);
or U1348 (N_1348,N_1025,N_534);
and U1349 (N_1349,N_561,N_159);
nand U1350 (N_1350,N_849,N_462);
or U1351 (N_1351,N_1066,N_652);
nand U1352 (N_1352,N_714,N_765);
or U1353 (N_1353,N_974,N_86);
nor U1354 (N_1354,N_787,N_769);
nand U1355 (N_1355,N_1232,N_78);
nor U1356 (N_1356,N_613,N_597);
or U1357 (N_1357,N_550,N_1110);
or U1358 (N_1358,N_1244,N_881);
nor U1359 (N_1359,N_635,N_347);
nor U1360 (N_1360,N_994,N_217);
nand U1361 (N_1361,N_21,N_617);
nor U1362 (N_1362,N_897,N_1147);
xor U1363 (N_1363,N_1014,N_137);
xnor U1364 (N_1364,N_491,N_685);
nand U1365 (N_1365,N_316,N_755);
or U1366 (N_1366,N_591,N_1095);
and U1367 (N_1367,N_721,N_836);
or U1368 (N_1368,N_605,N_79);
and U1369 (N_1369,N_886,N_134);
xor U1370 (N_1370,N_1081,N_396);
and U1371 (N_1371,N_841,N_907);
nand U1372 (N_1372,N_639,N_602);
nor U1373 (N_1373,N_447,N_736);
or U1374 (N_1374,N_270,N_913);
xor U1375 (N_1375,N_1141,N_348);
xnor U1376 (N_1376,N_106,N_425);
nor U1377 (N_1377,N_1160,N_544);
xor U1378 (N_1378,N_560,N_124);
xor U1379 (N_1379,N_1108,N_307);
or U1380 (N_1380,N_893,N_870);
nor U1381 (N_1381,N_703,N_1006);
xor U1382 (N_1382,N_837,N_274);
nor U1383 (N_1383,N_1241,N_812);
and U1384 (N_1384,N_889,N_634);
xor U1385 (N_1385,N_162,N_546);
or U1386 (N_1386,N_663,N_555);
nand U1387 (N_1387,N_594,N_1127);
and U1388 (N_1388,N_1118,N_1109);
nor U1389 (N_1389,N_125,N_832);
xor U1390 (N_1390,N_478,N_536);
nor U1391 (N_1391,N_589,N_395);
nor U1392 (N_1392,N_1068,N_210);
or U1393 (N_1393,N_571,N_1124);
and U1394 (N_1394,N_399,N_170);
nor U1395 (N_1395,N_1011,N_1090);
nand U1396 (N_1396,N_1111,N_906);
xor U1397 (N_1397,N_122,N_1202);
nor U1398 (N_1398,N_430,N_511);
nand U1399 (N_1399,N_62,N_843);
nor U1400 (N_1400,N_379,N_1016);
xor U1401 (N_1401,N_253,N_687);
or U1402 (N_1402,N_840,N_1145);
and U1403 (N_1403,N_507,N_179);
or U1404 (N_1404,N_1091,N_1120);
or U1405 (N_1405,N_391,N_828);
xnor U1406 (N_1406,N_110,N_23);
nand U1407 (N_1407,N_809,N_905);
or U1408 (N_1408,N_1053,N_793);
nand U1409 (N_1409,N_1119,N_653);
or U1410 (N_1410,N_508,N_1235);
nor U1411 (N_1411,N_1165,N_1022);
or U1412 (N_1412,N_798,N_668);
and U1413 (N_1413,N_900,N_860);
nor U1414 (N_1414,N_1052,N_306);
and U1415 (N_1415,N_222,N_322);
xnor U1416 (N_1416,N_432,N_509);
and U1417 (N_1417,N_671,N_532);
and U1418 (N_1418,N_817,N_551);
or U1419 (N_1419,N_1243,N_1032);
nor U1420 (N_1420,N_378,N_64);
nand U1421 (N_1421,N_531,N_684);
nand U1422 (N_1422,N_450,N_515);
nand U1423 (N_1423,N_225,N_245);
xor U1424 (N_1424,N_586,N_93);
and U1425 (N_1425,N_139,N_55);
or U1426 (N_1426,N_1163,N_477);
nor U1427 (N_1427,N_58,N_85);
or U1428 (N_1428,N_651,N_1017);
nand U1429 (N_1429,N_839,N_788);
nor U1430 (N_1430,N_712,N_976);
nand U1431 (N_1431,N_655,N_1083);
and U1432 (N_1432,N_242,N_654);
nand U1433 (N_1433,N_1194,N_984);
nand U1434 (N_1434,N_582,N_220);
or U1435 (N_1435,N_308,N_1180);
or U1436 (N_1436,N_762,N_569);
xor U1437 (N_1437,N_1122,N_1023);
and U1438 (N_1438,N_228,N_318);
xnor U1439 (N_1439,N_943,N_1131);
xor U1440 (N_1440,N_1033,N_985);
xnor U1441 (N_1441,N_163,N_1001);
and U1442 (N_1442,N_1015,N_1055);
and U1443 (N_1443,N_10,N_401);
nor U1444 (N_1444,N_1085,N_838);
nor U1445 (N_1445,N_435,N_630);
and U1446 (N_1446,N_727,N_631);
and U1447 (N_1447,N_880,N_992);
or U1448 (N_1448,N_182,N_585);
xor U1449 (N_1449,N_302,N_506);
xnor U1450 (N_1450,N_528,N_1037);
xor U1451 (N_1451,N_160,N_377);
and U1452 (N_1452,N_1249,N_409);
xor U1453 (N_1453,N_1059,N_291);
nor U1454 (N_1454,N_1105,N_1142);
nor U1455 (N_1455,N_948,N_851);
or U1456 (N_1456,N_56,N_367);
nand U1457 (N_1457,N_169,N_2);
nor U1458 (N_1458,N_869,N_42);
nor U1459 (N_1459,N_1222,N_510);
nor U1460 (N_1460,N_572,N_407);
or U1461 (N_1461,N_833,N_1221);
nand U1462 (N_1462,N_1239,N_995);
and U1463 (N_1463,N_899,N_850);
or U1464 (N_1464,N_1116,N_305);
nor U1465 (N_1465,N_1060,N_336);
or U1466 (N_1466,N_892,N_226);
and U1467 (N_1467,N_1133,N_1007);
and U1468 (N_1468,N_315,N_70);
nand U1469 (N_1469,N_32,N_116);
nor U1470 (N_1470,N_1043,N_801);
and U1471 (N_1471,N_89,N_390);
xor U1472 (N_1472,N_1076,N_1162);
or U1473 (N_1473,N_0,N_1038);
or U1474 (N_1474,N_644,N_683);
nand U1475 (N_1475,N_88,N_424);
nor U1476 (N_1476,N_1115,N_292);
and U1477 (N_1477,N_807,N_80);
nor U1478 (N_1478,N_341,N_187);
xnor U1479 (N_1479,N_1106,N_219);
and U1480 (N_1480,N_690,N_871);
and U1481 (N_1481,N_603,N_1185);
and U1482 (N_1482,N_174,N_689);
nand U1483 (N_1483,N_1207,N_614);
xor U1484 (N_1484,N_626,N_75);
xor U1485 (N_1485,N_39,N_451);
or U1486 (N_1486,N_140,N_466);
xor U1487 (N_1487,N_143,N_173);
nor U1488 (N_1488,N_211,N_1174);
nand U1489 (N_1489,N_148,N_1041);
or U1490 (N_1490,N_54,N_611);
and U1491 (N_1491,N_578,N_327);
and U1492 (N_1492,N_945,N_445);
or U1493 (N_1493,N_763,N_958);
nor U1494 (N_1494,N_896,N_830);
and U1495 (N_1495,N_123,N_1186);
or U1496 (N_1496,N_916,N_1030);
xnor U1497 (N_1497,N_501,N_885);
nor U1498 (N_1498,N_520,N_625);
nor U1499 (N_1499,N_556,N_780);
and U1500 (N_1500,N_299,N_268);
or U1501 (N_1501,N_69,N_681);
or U1502 (N_1502,N_606,N_612);
and U1503 (N_1503,N_1000,N_29);
and U1504 (N_1504,N_883,N_1087);
and U1505 (N_1505,N_986,N_646);
xnor U1506 (N_1506,N_686,N_1215);
nor U1507 (N_1507,N_1020,N_519);
xor U1508 (N_1508,N_815,N_1067);
and U1509 (N_1509,N_1150,N_138);
and U1510 (N_1510,N_950,N_688);
nor U1511 (N_1511,N_471,N_288);
or U1512 (N_1512,N_261,N_195);
nor U1513 (N_1513,N_398,N_19);
nor U1514 (N_1514,N_11,N_154);
xor U1515 (N_1515,N_914,N_740);
xnor U1516 (N_1516,N_922,N_1155);
and U1517 (N_1517,N_576,N_149);
xnor U1518 (N_1518,N_280,N_522);
nor U1519 (N_1519,N_455,N_467);
nor U1520 (N_1520,N_577,N_329);
and U1521 (N_1521,N_332,N_980);
and U1522 (N_1522,N_304,N_732);
nand U1523 (N_1523,N_1074,N_172);
nor U1524 (N_1524,N_667,N_1144);
or U1525 (N_1525,N_737,N_872);
or U1526 (N_1526,N_1166,N_797);
or U1527 (N_1527,N_481,N_203);
nand U1528 (N_1528,N_526,N_354);
nand U1529 (N_1529,N_178,N_944);
xor U1530 (N_1530,N_901,N_734);
and U1531 (N_1531,N_155,N_1238);
nand U1532 (N_1532,N_67,N_1062);
xnor U1533 (N_1533,N_616,N_699);
nand U1534 (N_1534,N_960,N_405);
or U1535 (N_1535,N_121,N_129);
xor U1536 (N_1536,N_197,N_675);
and U1537 (N_1537,N_112,N_1140);
nor U1538 (N_1538,N_676,N_567);
xor U1539 (N_1539,N_865,N_759);
and U1540 (N_1540,N_926,N_1039);
xor U1541 (N_1541,N_829,N_1134);
and U1542 (N_1542,N_360,N_205);
xor U1543 (N_1543,N_1005,N_408);
nand U1544 (N_1544,N_175,N_453);
xor U1545 (N_1545,N_648,N_60);
nand U1546 (N_1546,N_1240,N_619);
or U1547 (N_1547,N_873,N_12);
xor U1548 (N_1548,N_818,N_344);
or U1549 (N_1549,N_750,N_72);
nor U1550 (N_1550,N_113,N_1019);
and U1551 (N_1551,N_212,N_133);
and U1552 (N_1552,N_965,N_61);
nor U1553 (N_1553,N_568,N_105);
xor U1554 (N_1554,N_1107,N_207);
xnor U1555 (N_1555,N_333,N_891);
nand U1556 (N_1556,N_864,N_1027);
xnor U1557 (N_1557,N_743,N_953);
or U1558 (N_1558,N_230,N_57);
and U1559 (N_1559,N_954,N_1125);
or U1560 (N_1560,N_662,N_1229);
or U1561 (N_1561,N_298,N_852);
nand U1562 (N_1562,N_682,N_200);
xor U1563 (N_1563,N_1248,N_723);
xor U1564 (N_1564,N_383,N_164);
and U1565 (N_1565,N_1179,N_166);
or U1566 (N_1566,N_132,N_202);
nand U1567 (N_1567,N_483,N_185);
xor U1568 (N_1568,N_25,N_100);
nand U1569 (N_1569,N_380,N_952);
or U1570 (N_1570,N_1169,N_1159);
xnor U1571 (N_1571,N_587,N_458);
and U1572 (N_1572,N_286,N_726);
xnor U1573 (N_1573,N_1008,N_368);
nor U1574 (N_1574,N_700,N_463);
xnor U1575 (N_1575,N_1230,N_468);
nand U1576 (N_1576,N_918,N_973);
or U1577 (N_1577,N_224,N_243);
or U1578 (N_1578,N_386,N_724);
nor U1579 (N_1579,N_328,N_521);
nand U1580 (N_1580,N_1164,N_442);
or U1581 (N_1581,N_672,N_1146);
and U1582 (N_1582,N_345,N_1072);
or U1583 (N_1583,N_1218,N_730);
and U1584 (N_1584,N_524,N_1220);
nand U1585 (N_1585,N_281,N_215);
nand U1586 (N_1586,N_191,N_107);
or U1587 (N_1587,N_1089,N_997);
nor U1588 (N_1588,N_258,N_73);
or U1589 (N_1589,N_1031,N_554);
xnor U1590 (N_1590,N_643,N_702);
nor U1591 (N_1591,N_40,N_825);
nor U1592 (N_1592,N_415,N_527);
and U1593 (N_1593,N_570,N_204);
and U1594 (N_1594,N_803,N_733);
and U1595 (N_1595,N_543,N_866);
nand U1596 (N_1596,N_991,N_82);
nor U1597 (N_1597,N_334,N_1104);
nand U1598 (N_1598,N_600,N_46);
nor U1599 (N_1599,N_811,N_1057);
nor U1600 (N_1600,N_320,N_249);
nand U1601 (N_1601,N_131,N_1084);
nand U1602 (N_1602,N_363,N_538);
nand U1603 (N_1603,N_800,N_441);
or U1604 (N_1604,N_642,N_939);
or U1605 (N_1605,N_842,N_284);
or U1606 (N_1606,N_779,N_439);
nand U1607 (N_1607,N_240,N_144);
or U1608 (N_1608,N_52,N_921);
xnor U1609 (N_1609,N_957,N_1101);
and U1610 (N_1610,N_198,N_247);
xnor U1611 (N_1611,N_720,N_1201);
xor U1612 (N_1612,N_479,N_95);
nor U1613 (N_1613,N_823,N_59);
nand U1614 (N_1614,N_638,N_353);
nor U1615 (N_1615,N_440,N_290);
or U1616 (N_1616,N_806,N_1247);
xnor U1617 (N_1617,N_400,N_43);
and U1618 (N_1618,N_33,N_221);
nor U1619 (N_1619,N_94,N_259);
nand U1620 (N_1620,N_41,N_382);
nor U1621 (N_1621,N_742,N_820);
nor U1622 (N_1622,N_627,N_562);
xor U1623 (N_1623,N_1195,N_5);
and U1624 (N_1624,N_764,N_622);
nand U1625 (N_1625,N_1182,N_340);
xnor U1626 (N_1626,N_37,N_63);
or U1627 (N_1627,N_708,N_988);
or U1628 (N_1628,N_474,N_92);
xnor U1629 (N_1629,N_604,N_325);
nor U1630 (N_1630,N_565,N_610);
nand U1631 (N_1631,N_887,N_476);
nand U1632 (N_1632,N_636,N_758);
nand U1633 (N_1633,N_620,N_76);
and U1634 (N_1634,N_1214,N_674);
nor U1635 (N_1635,N_417,N_1137);
or U1636 (N_1636,N_314,N_27);
xor U1637 (N_1637,N_397,N_1149);
nand U1638 (N_1638,N_1078,N_365);
nor U1639 (N_1639,N_637,N_91);
nor U1640 (N_1640,N_1047,N_495);
nand U1641 (N_1641,N_1193,N_1099);
xnor U1642 (N_1642,N_282,N_890);
xor U1643 (N_1643,N_753,N_1172);
xor U1644 (N_1644,N_867,N_264);
xnor U1645 (N_1645,N_924,N_251);
nand U1646 (N_1646,N_1224,N_673);
nor U1647 (N_1647,N_876,N_754);
and U1648 (N_1648,N_791,N_3);
xnor U1649 (N_1649,N_262,N_503);
nor U1650 (N_1650,N_1117,N_628);
and U1651 (N_1651,N_701,N_805);
nor U1652 (N_1652,N_99,N_910);
nor U1653 (N_1653,N_489,N_799);
nand U1654 (N_1654,N_821,N_372);
and U1655 (N_1655,N_218,N_180);
nor U1656 (N_1656,N_563,N_963);
xor U1657 (N_1657,N_490,N_6);
or U1658 (N_1658,N_17,N_932);
or U1659 (N_1659,N_15,N_553);
or U1660 (N_1660,N_1233,N_609);
and U1661 (N_1661,N_236,N_1073);
or U1662 (N_1662,N_912,N_539);
or U1663 (N_1663,N_919,N_1126);
and U1664 (N_1664,N_579,N_1034);
nor U1665 (N_1665,N_861,N_254);
or U1666 (N_1666,N_540,N_349);
or U1667 (N_1667,N_927,N_406);
nand U1668 (N_1668,N_238,N_199);
xor U1669 (N_1669,N_659,N_194);
nand U1670 (N_1670,N_456,N_1102);
nand U1671 (N_1671,N_165,N_942);
nand U1672 (N_1672,N_936,N_429);
nand U1673 (N_1673,N_168,N_967);
nand U1674 (N_1674,N_1029,N_959);
nor U1675 (N_1675,N_443,N_1061);
xor U1676 (N_1676,N_795,N_1139);
and U1677 (N_1677,N_650,N_428);
nand U1678 (N_1678,N_1065,N_1191);
nor U1679 (N_1679,N_518,N_731);
nor U1680 (N_1680,N_1079,N_898);
nor U1681 (N_1681,N_810,N_1153);
nand U1682 (N_1682,N_513,N_680);
xor U1683 (N_1683,N_255,N_1219);
nand U1684 (N_1684,N_136,N_999);
or U1685 (N_1685,N_1171,N_1096);
or U1686 (N_1686,N_422,N_1181);
and U1687 (N_1687,N_770,N_566);
nor U1688 (N_1688,N_1013,N_930);
or U1689 (N_1689,N_822,N_321);
nand U1690 (N_1690,N_789,N_234);
nand U1691 (N_1691,N_114,N_184);
and U1692 (N_1692,N_1028,N_414);
nand U1693 (N_1693,N_756,N_461);
and U1694 (N_1694,N_161,N_1154);
nor U1695 (N_1695,N_802,N_289);
nand U1696 (N_1696,N_189,N_738);
nand U1697 (N_1697,N_983,N_598);
nand U1698 (N_1698,N_710,N_237);
nand U1699 (N_1699,N_713,N_319);
or U1700 (N_1700,N_361,N_547);
or U1701 (N_1701,N_167,N_130);
and U1702 (N_1702,N_580,N_487);
or U1703 (N_1703,N_496,N_782);
nor U1704 (N_1704,N_1121,N_371);
and U1705 (N_1705,N_1103,N_962);
xnor U1706 (N_1706,N_804,N_657);
and U1707 (N_1707,N_188,N_357);
nor U1708 (N_1708,N_358,N_1093);
and U1709 (N_1709,N_1100,N_276);
nand U1710 (N_1710,N_909,N_588);
or U1711 (N_1711,N_1198,N_982);
nand U1712 (N_1712,N_469,N_410);
nor U1713 (N_1713,N_784,N_847);
nand U1714 (N_1714,N_317,N_192);
nand U1715 (N_1715,N_894,N_584);
nor U1716 (N_1716,N_459,N_421);
nor U1717 (N_1717,N_649,N_878);
xnor U1718 (N_1718,N_998,N_752);
nor U1719 (N_1719,N_7,N_596);
nor U1720 (N_1720,N_350,N_28);
nand U1721 (N_1721,N_951,N_1042);
xor U1722 (N_1722,N_1046,N_150);
xnor U1723 (N_1723,N_263,N_1004);
nand U1724 (N_1724,N_533,N_968);
and U1725 (N_1725,N_777,N_595);
xor U1726 (N_1726,N_794,N_356);
and U1727 (N_1727,N_404,N_504);
nand U1728 (N_1728,N_232,N_1045);
and U1729 (N_1729,N_369,N_485);
nand U1730 (N_1730,N_283,N_530);
xor U1731 (N_1731,N_103,N_492);
nor U1732 (N_1732,N_98,N_250);
and U1733 (N_1733,N_955,N_656);
nor U1734 (N_1734,N_1123,N_493);
xnor U1735 (N_1735,N_529,N_1196);
nand U1736 (N_1736,N_1143,N_426);
nor U1737 (N_1737,N_389,N_704);
xor U1738 (N_1738,N_665,N_1049);
and U1739 (N_1739,N_310,N_1237);
nor U1740 (N_1740,N_895,N_1003);
and U1741 (N_1741,N_208,N_48);
or U1742 (N_1742,N_785,N_875);
or U1743 (N_1743,N_975,N_343);
and U1744 (N_1744,N_206,N_342);
nand U1745 (N_1745,N_773,N_786);
xor U1746 (N_1746,N_201,N_879);
and U1747 (N_1747,N_1168,N_352);
xnor U1748 (N_1748,N_902,N_190);
nand U1749 (N_1749,N_1217,N_1018);
nor U1750 (N_1750,N_693,N_183);
nand U1751 (N_1751,N_705,N_294);
and U1752 (N_1752,N_1051,N_44);
or U1753 (N_1753,N_362,N_1021);
nor U1754 (N_1754,N_216,N_601);
nor U1755 (N_1755,N_488,N_694);
nor U1756 (N_1756,N_552,N_816);
xnor U1757 (N_1757,N_387,N_744);
or U1758 (N_1758,N_403,N_884);
nor U1759 (N_1759,N_666,N_373);
nand U1760 (N_1760,N_981,N_735);
nand U1761 (N_1761,N_855,N_296);
xor U1762 (N_1762,N_117,N_142);
nor U1763 (N_1763,N_923,N_351);
nand U1764 (N_1764,N_696,N_301);
or U1765 (N_1765,N_120,N_484);
xor U1766 (N_1766,N_670,N_647);
nand U1767 (N_1767,N_966,N_470);
nor U1768 (N_1768,N_835,N_1086);
and U1769 (N_1769,N_535,N_359);
or U1770 (N_1770,N_808,N_1176);
or U1771 (N_1771,N_502,N_309);
xnor U1772 (N_1772,N_68,N_51);
nand U1773 (N_1773,N_854,N_698);
xnor U1774 (N_1774,N_768,N_772);
nand U1775 (N_1775,N_677,N_928);
nor U1776 (N_1776,N_573,N_989);
nand U1777 (N_1777,N_252,N_725);
and U1778 (N_1778,N_757,N_346);
and U1779 (N_1779,N_1071,N_946);
nand U1780 (N_1780,N_516,N_949);
nand U1781 (N_1781,N_1026,N_1035);
or U1782 (N_1782,N_96,N_545);
or U1783 (N_1783,N_862,N_77);
nand U1784 (N_1784,N_47,N_248);
nor U1785 (N_1785,N_505,N_257);
and U1786 (N_1786,N_1161,N_53);
xnor U1787 (N_1787,N_541,N_826);
nand U1788 (N_1788,N_364,N_330);
xnor U1789 (N_1789,N_339,N_1157);
and U1790 (N_1790,N_549,N_751);
and U1791 (N_1791,N_473,N_1228);
nand U1792 (N_1792,N_420,N_947);
nor U1793 (N_1793,N_697,N_977);
nand U1794 (N_1794,N_629,N_393);
or U1795 (N_1795,N_1024,N_608);
and U1796 (N_1796,N_1097,N_1009);
nand U1797 (N_1797,N_599,N_1203);
and U1798 (N_1798,N_917,N_970);
and U1799 (N_1799,N_1002,N_1167);
and U1800 (N_1800,N_1044,N_337);
or U1801 (N_1801,N_853,N_1223);
or U1802 (N_1802,N_229,N_1189);
and U1803 (N_1803,N_127,N_858);
or U1804 (N_1804,N_706,N_14);
nand U1805 (N_1805,N_104,N_24);
nor U1806 (N_1806,N_1199,N_375);
or U1807 (N_1807,N_74,N_956);
and U1808 (N_1808,N_448,N_558);
or U1809 (N_1809,N_920,N_36);
nor U1810 (N_1810,N_223,N_517);
nand U1811 (N_1811,N_661,N_940);
xnor U1812 (N_1812,N_235,N_1178);
nand U1813 (N_1813,N_423,N_1211);
nand U1814 (N_1814,N_374,N_66);
nor U1815 (N_1815,N_1152,N_848);
nand U1816 (N_1816,N_277,N_990);
xnor U1817 (N_1817,N_244,N_575);
xor U1818 (N_1818,N_1173,N_592);
xnor U1819 (N_1819,N_748,N_269);
nor U1820 (N_1820,N_153,N_796);
or U1821 (N_1821,N_1213,N_846);
or U1822 (N_1822,N_760,N_266);
or U1823 (N_1823,N_1135,N_583);
and U1824 (N_1824,N_1058,N_1138);
nor U1825 (N_1825,N_464,N_1063);
nand U1826 (N_1826,N_1077,N_480);
xor U1827 (N_1827,N_34,N_438);
and U1828 (N_1828,N_30,N_692);
xor U1829 (N_1829,N_523,N_444);
nor U1830 (N_1830,N_1187,N_376);
nor U1831 (N_1831,N_621,N_267);
or U1832 (N_1832,N_141,N_618);
and U1833 (N_1833,N_18,N_8);
xnor U1834 (N_1834,N_324,N_418);
or U1835 (N_1835,N_256,N_128);
xor U1836 (N_1836,N_241,N_615);
nor U1837 (N_1837,N_834,N_1200);
nor U1838 (N_1838,N_303,N_1197);
xnor U1839 (N_1839,N_312,N_101);
or U1840 (N_1840,N_97,N_486);
nand U1841 (N_1841,N_156,N_152);
or U1842 (N_1842,N_1225,N_326);
and U1843 (N_1843,N_297,N_177);
xnor U1844 (N_1844,N_971,N_84);
or U1845 (N_1845,N_969,N_739);
nand U1846 (N_1846,N_119,N_1114);
nand U1847 (N_1847,N_370,N_385);
and U1848 (N_1848,N_776,N_778);
xnor U1849 (N_1849,N_157,N_193);
or U1850 (N_1850,N_394,N_904);
nand U1851 (N_1851,N_402,N_827);
nand U1852 (N_1852,N_783,N_908);
or U1853 (N_1853,N_355,N_186);
xor U1854 (N_1854,N_548,N_1128);
or U1855 (N_1855,N_151,N_790);
nor U1856 (N_1856,N_717,N_176);
nor U1857 (N_1857,N_1151,N_102);
nor U1858 (N_1858,N_384,N_669);
or U1859 (N_1859,N_857,N_728);
or U1860 (N_1860,N_147,N_13);
or U1861 (N_1861,N_903,N_323);
nor U1862 (N_1862,N_1136,N_859);
or U1863 (N_1863,N_295,N_771);
nand U1864 (N_1864,N_1132,N_449);
or U1865 (N_1865,N_964,N_978);
and U1866 (N_1866,N_1236,N_213);
and U1867 (N_1867,N_766,N_660);
xor U1868 (N_1868,N_366,N_273);
nand U1869 (N_1869,N_411,N_279);
or U1870 (N_1870,N_645,N_972);
xor U1871 (N_1871,N_542,N_115);
nand U1872 (N_1872,N_214,N_499);
xnor U1873 (N_1873,N_436,N_457);
or U1874 (N_1874,N_1242,N_108);
or U1875 (N_1875,N_242,N_1227);
nand U1876 (N_1876,N_1074,N_306);
xor U1877 (N_1877,N_788,N_895);
xnor U1878 (N_1878,N_18,N_1011);
and U1879 (N_1879,N_471,N_777);
nand U1880 (N_1880,N_876,N_756);
and U1881 (N_1881,N_1076,N_985);
nor U1882 (N_1882,N_1082,N_832);
or U1883 (N_1883,N_528,N_1043);
and U1884 (N_1884,N_1033,N_323);
nor U1885 (N_1885,N_652,N_422);
nand U1886 (N_1886,N_449,N_1159);
or U1887 (N_1887,N_597,N_675);
or U1888 (N_1888,N_936,N_676);
or U1889 (N_1889,N_1009,N_43);
nor U1890 (N_1890,N_377,N_1193);
or U1891 (N_1891,N_441,N_135);
or U1892 (N_1892,N_1181,N_377);
and U1893 (N_1893,N_66,N_144);
and U1894 (N_1894,N_975,N_695);
nand U1895 (N_1895,N_1017,N_336);
and U1896 (N_1896,N_685,N_451);
or U1897 (N_1897,N_1089,N_1235);
or U1898 (N_1898,N_750,N_993);
and U1899 (N_1899,N_708,N_390);
and U1900 (N_1900,N_991,N_45);
and U1901 (N_1901,N_1180,N_801);
nor U1902 (N_1902,N_304,N_750);
or U1903 (N_1903,N_245,N_423);
or U1904 (N_1904,N_960,N_807);
xnor U1905 (N_1905,N_224,N_593);
xor U1906 (N_1906,N_1114,N_212);
xnor U1907 (N_1907,N_1118,N_388);
xnor U1908 (N_1908,N_129,N_270);
and U1909 (N_1909,N_105,N_101);
nand U1910 (N_1910,N_204,N_1084);
xnor U1911 (N_1911,N_407,N_764);
and U1912 (N_1912,N_321,N_970);
nor U1913 (N_1913,N_1013,N_670);
nand U1914 (N_1914,N_247,N_741);
and U1915 (N_1915,N_518,N_820);
and U1916 (N_1916,N_193,N_1206);
xnor U1917 (N_1917,N_921,N_581);
and U1918 (N_1918,N_29,N_311);
nand U1919 (N_1919,N_206,N_148);
nor U1920 (N_1920,N_829,N_1008);
nor U1921 (N_1921,N_866,N_1181);
nor U1922 (N_1922,N_670,N_915);
or U1923 (N_1923,N_754,N_1027);
xor U1924 (N_1924,N_921,N_529);
nor U1925 (N_1925,N_158,N_933);
and U1926 (N_1926,N_1176,N_294);
nor U1927 (N_1927,N_866,N_699);
xnor U1928 (N_1928,N_797,N_981);
xnor U1929 (N_1929,N_130,N_79);
or U1930 (N_1930,N_1188,N_242);
xnor U1931 (N_1931,N_219,N_1012);
and U1932 (N_1932,N_478,N_307);
nor U1933 (N_1933,N_997,N_888);
or U1934 (N_1934,N_128,N_110);
nand U1935 (N_1935,N_911,N_705);
and U1936 (N_1936,N_936,N_148);
nor U1937 (N_1937,N_384,N_929);
nor U1938 (N_1938,N_1115,N_36);
xor U1939 (N_1939,N_369,N_623);
or U1940 (N_1940,N_1050,N_40);
xnor U1941 (N_1941,N_310,N_726);
and U1942 (N_1942,N_31,N_783);
nor U1943 (N_1943,N_534,N_1028);
nand U1944 (N_1944,N_1155,N_1237);
or U1945 (N_1945,N_696,N_1135);
nor U1946 (N_1946,N_1247,N_186);
xor U1947 (N_1947,N_1151,N_844);
or U1948 (N_1948,N_173,N_252);
nor U1949 (N_1949,N_538,N_964);
and U1950 (N_1950,N_365,N_960);
nor U1951 (N_1951,N_453,N_896);
or U1952 (N_1952,N_265,N_366);
nor U1953 (N_1953,N_1039,N_216);
and U1954 (N_1954,N_1013,N_1025);
and U1955 (N_1955,N_320,N_825);
nand U1956 (N_1956,N_49,N_333);
xor U1957 (N_1957,N_58,N_224);
nor U1958 (N_1958,N_543,N_1049);
nor U1959 (N_1959,N_812,N_329);
xnor U1960 (N_1960,N_753,N_93);
or U1961 (N_1961,N_831,N_910);
xor U1962 (N_1962,N_184,N_249);
and U1963 (N_1963,N_971,N_449);
nor U1964 (N_1964,N_596,N_199);
nor U1965 (N_1965,N_771,N_944);
xnor U1966 (N_1966,N_569,N_1209);
nand U1967 (N_1967,N_958,N_665);
and U1968 (N_1968,N_527,N_935);
or U1969 (N_1969,N_1212,N_1171);
nand U1970 (N_1970,N_43,N_75);
nor U1971 (N_1971,N_762,N_1134);
xnor U1972 (N_1972,N_202,N_885);
and U1973 (N_1973,N_557,N_361);
and U1974 (N_1974,N_611,N_1150);
xor U1975 (N_1975,N_499,N_1113);
xnor U1976 (N_1976,N_733,N_859);
xnor U1977 (N_1977,N_446,N_636);
nand U1978 (N_1978,N_822,N_435);
nand U1979 (N_1979,N_433,N_919);
or U1980 (N_1980,N_628,N_491);
nor U1981 (N_1981,N_1052,N_337);
nor U1982 (N_1982,N_627,N_358);
or U1983 (N_1983,N_1090,N_1064);
or U1984 (N_1984,N_314,N_1149);
and U1985 (N_1985,N_990,N_225);
and U1986 (N_1986,N_614,N_218);
or U1987 (N_1987,N_733,N_969);
nand U1988 (N_1988,N_43,N_48);
nand U1989 (N_1989,N_942,N_636);
nand U1990 (N_1990,N_202,N_412);
xnor U1991 (N_1991,N_1088,N_246);
nor U1992 (N_1992,N_831,N_933);
and U1993 (N_1993,N_91,N_1188);
xnor U1994 (N_1994,N_1222,N_702);
nor U1995 (N_1995,N_12,N_1192);
nor U1996 (N_1996,N_485,N_544);
or U1997 (N_1997,N_65,N_836);
and U1998 (N_1998,N_629,N_12);
nor U1999 (N_1999,N_991,N_585);
nand U2000 (N_2000,N_864,N_219);
xnor U2001 (N_2001,N_1118,N_162);
or U2002 (N_2002,N_1203,N_79);
and U2003 (N_2003,N_922,N_739);
or U2004 (N_2004,N_453,N_1114);
and U2005 (N_2005,N_509,N_434);
or U2006 (N_2006,N_1236,N_784);
or U2007 (N_2007,N_339,N_255);
xor U2008 (N_2008,N_1071,N_375);
xnor U2009 (N_2009,N_1159,N_758);
xor U2010 (N_2010,N_624,N_222);
or U2011 (N_2011,N_198,N_932);
nor U2012 (N_2012,N_879,N_825);
xor U2013 (N_2013,N_85,N_822);
and U2014 (N_2014,N_885,N_103);
nand U2015 (N_2015,N_921,N_206);
or U2016 (N_2016,N_1190,N_435);
nand U2017 (N_2017,N_251,N_307);
nor U2018 (N_2018,N_1023,N_930);
and U2019 (N_2019,N_618,N_1154);
nand U2020 (N_2020,N_741,N_784);
and U2021 (N_2021,N_663,N_291);
and U2022 (N_2022,N_96,N_40);
xnor U2023 (N_2023,N_843,N_1014);
and U2024 (N_2024,N_222,N_925);
nand U2025 (N_2025,N_721,N_398);
or U2026 (N_2026,N_915,N_900);
nor U2027 (N_2027,N_207,N_271);
and U2028 (N_2028,N_915,N_0);
or U2029 (N_2029,N_683,N_596);
or U2030 (N_2030,N_843,N_1055);
xor U2031 (N_2031,N_1247,N_1000);
and U2032 (N_2032,N_972,N_1198);
or U2033 (N_2033,N_1193,N_446);
nor U2034 (N_2034,N_1231,N_679);
and U2035 (N_2035,N_1110,N_396);
nor U2036 (N_2036,N_735,N_413);
xor U2037 (N_2037,N_862,N_361);
xor U2038 (N_2038,N_19,N_355);
or U2039 (N_2039,N_487,N_939);
nand U2040 (N_2040,N_124,N_1213);
xor U2041 (N_2041,N_245,N_374);
nor U2042 (N_2042,N_1138,N_151);
or U2043 (N_2043,N_399,N_193);
xnor U2044 (N_2044,N_1207,N_938);
or U2045 (N_2045,N_594,N_989);
xnor U2046 (N_2046,N_657,N_789);
nor U2047 (N_2047,N_786,N_570);
or U2048 (N_2048,N_46,N_676);
and U2049 (N_2049,N_441,N_490);
and U2050 (N_2050,N_316,N_299);
nand U2051 (N_2051,N_878,N_74);
and U2052 (N_2052,N_988,N_305);
nor U2053 (N_2053,N_898,N_1059);
nand U2054 (N_2054,N_79,N_119);
nand U2055 (N_2055,N_439,N_903);
and U2056 (N_2056,N_1011,N_733);
nand U2057 (N_2057,N_229,N_167);
or U2058 (N_2058,N_1212,N_202);
and U2059 (N_2059,N_951,N_0);
and U2060 (N_2060,N_153,N_123);
nor U2061 (N_2061,N_803,N_1081);
or U2062 (N_2062,N_1190,N_652);
or U2063 (N_2063,N_359,N_91);
xnor U2064 (N_2064,N_375,N_71);
xor U2065 (N_2065,N_720,N_1091);
nor U2066 (N_2066,N_436,N_870);
nor U2067 (N_2067,N_901,N_593);
and U2068 (N_2068,N_676,N_458);
and U2069 (N_2069,N_227,N_940);
and U2070 (N_2070,N_315,N_805);
and U2071 (N_2071,N_607,N_339);
nand U2072 (N_2072,N_1006,N_413);
or U2073 (N_2073,N_942,N_1199);
and U2074 (N_2074,N_756,N_783);
or U2075 (N_2075,N_317,N_1088);
or U2076 (N_2076,N_139,N_170);
nand U2077 (N_2077,N_622,N_647);
or U2078 (N_2078,N_642,N_801);
and U2079 (N_2079,N_326,N_579);
nor U2080 (N_2080,N_310,N_924);
xor U2081 (N_2081,N_1245,N_140);
xnor U2082 (N_2082,N_985,N_414);
nand U2083 (N_2083,N_822,N_748);
nor U2084 (N_2084,N_1228,N_895);
xnor U2085 (N_2085,N_1145,N_899);
xnor U2086 (N_2086,N_1115,N_703);
or U2087 (N_2087,N_227,N_210);
and U2088 (N_2088,N_87,N_1036);
nand U2089 (N_2089,N_920,N_654);
xnor U2090 (N_2090,N_350,N_121);
or U2091 (N_2091,N_1144,N_956);
xor U2092 (N_2092,N_85,N_875);
nor U2093 (N_2093,N_42,N_683);
and U2094 (N_2094,N_321,N_1159);
xnor U2095 (N_2095,N_552,N_36);
nand U2096 (N_2096,N_415,N_923);
and U2097 (N_2097,N_921,N_1163);
nand U2098 (N_2098,N_672,N_449);
or U2099 (N_2099,N_4,N_756);
and U2100 (N_2100,N_693,N_536);
xnor U2101 (N_2101,N_1225,N_632);
nor U2102 (N_2102,N_1095,N_1089);
nand U2103 (N_2103,N_706,N_138);
or U2104 (N_2104,N_967,N_402);
nand U2105 (N_2105,N_45,N_172);
xor U2106 (N_2106,N_1065,N_633);
nor U2107 (N_2107,N_837,N_1058);
and U2108 (N_2108,N_815,N_1182);
nand U2109 (N_2109,N_547,N_754);
xor U2110 (N_2110,N_408,N_657);
nor U2111 (N_2111,N_556,N_406);
nand U2112 (N_2112,N_291,N_806);
xnor U2113 (N_2113,N_1141,N_81);
and U2114 (N_2114,N_317,N_4);
or U2115 (N_2115,N_335,N_1085);
nor U2116 (N_2116,N_272,N_115);
nand U2117 (N_2117,N_735,N_374);
nor U2118 (N_2118,N_244,N_1149);
nand U2119 (N_2119,N_233,N_270);
nor U2120 (N_2120,N_684,N_1203);
nand U2121 (N_2121,N_154,N_590);
or U2122 (N_2122,N_32,N_917);
or U2123 (N_2123,N_671,N_121);
or U2124 (N_2124,N_1181,N_703);
xor U2125 (N_2125,N_869,N_484);
nor U2126 (N_2126,N_593,N_182);
or U2127 (N_2127,N_987,N_760);
nand U2128 (N_2128,N_889,N_739);
and U2129 (N_2129,N_1034,N_580);
and U2130 (N_2130,N_12,N_1012);
nor U2131 (N_2131,N_1007,N_1043);
nor U2132 (N_2132,N_38,N_453);
or U2133 (N_2133,N_784,N_229);
nor U2134 (N_2134,N_612,N_305);
xor U2135 (N_2135,N_9,N_618);
nand U2136 (N_2136,N_796,N_140);
nand U2137 (N_2137,N_319,N_736);
nor U2138 (N_2138,N_926,N_1104);
and U2139 (N_2139,N_340,N_918);
nor U2140 (N_2140,N_63,N_608);
nand U2141 (N_2141,N_28,N_447);
nand U2142 (N_2142,N_1116,N_104);
or U2143 (N_2143,N_504,N_778);
and U2144 (N_2144,N_1122,N_750);
or U2145 (N_2145,N_30,N_116);
nand U2146 (N_2146,N_1225,N_692);
xor U2147 (N_2147,N_160,N_1181);
and U2148 (N_2148,N_666,N_816);
xor U2149 (N_2149,N_101,N_1207);
and U2150 (N_2150,N_484,N_685);
nand U2151 (N_2151,N_541,N_1248);
nand U2152 (N_2152,N_385,N_470);
xor U2153 (N_2153,N_879,N_125);
nor U2154 (N_2154,N_1015,N_189);
or U2155 (N_2155,N_1021,N_1200);
or U2156 (N_2156,N_1214,N_963);
and U2157 (N_2157,N_441,N_867);
or U2158 (N_2158,N_1089,N_910);
xor U2159 (N_2159,N_231,N_982);
or U2160 (N_2160,N_1185,N_145);
nand U2161 (N_2161,N_558,N_260);
nand U2162 (N_2162,N_38,N_834);
xor U2163 (N_2163,N_1164,N_410);
or U2164 (N_2164,N_229,N_270);
xnor U2165 (N_2165,N_1170,N_311);
nor U2166 (N_2166,N_558,N_1041);
nand U2167 (N_2167,N_73,N_1156);
nor U2168 (N_2168,N_384,N_862);
or U2169 (N_2169,N_498,N_586);
xnor U2170 (N_2170,N_674,N_338);
nor U2171 (N_2171,N_923,N_1165);
xor U2172 (N_2172,N_193,N_221);
xor U2173 (N_2173,N_501,N_671);
xor U2174 (N_2174,N_956,N_669);
and U2175 (N_2175,N_1143,N_1011);
and U2176 (N_2176,N_737,N_616);
nand U2177 (N_2177,N_228,N_269);
and U2178 (N_2178,N_14,N_318);
nand U2179 (N_2179,N_1081,N_45);
and U2180 (N_2180,N_258,N_562);
nor U2181 (N_2181,N_184,N_1090);
xnor U2182 (N_2182,N_400,N_92);
xor U2183 (N_2183,N_334,N_1112);
xnor U2184 (N_2184,N_140,N_710);
xor U2185 (N_2185,N_88,N_696);
and U2186 (N_2186,N_1119,N_498);
nand U2187 (N_2187,N_1064,N_713);
nor U2188 (N_2188,N_206,N_503);
nand U2189 (N_2189,N_477,N_425);
xnor U2190 (N_2190,N_568,N_454);
nor U2191 (N_2191,N_438,N_1057);
xor U2192 (N_2192,N_251,N_207);
or U2193 (N_2193,N_190,N_1193);
nor U2194 (N_2194,N_1081,N_330);
nand U2195 (N_2195,N_442,N_418);
or U2196 (N_2196,N_773,N_646);
nor U2197 (N_2197,N_519,N_908);
nand U2198 (N_2198,N_716,N_1174);
nor U2199 (N_2199,N_749,N_593);
and U2200 (N_2200,N_154,N_951);
nand U2201 (N_2201,N_823,N_644);
xnor U2202 (N_2202,N_1110,N_963);
xnor U2203 (N_2203,N_84,N_621);
or U2204 (N_2204,N_444,N_684);
and U2205 (N_2205,N_666,N_311);
and U2206 (N_2206,N_372,N_335);
xnor U2207 (N_2207,N_123,N_856);
xor U2208 (N_2208,N_37,N_811);
xor U2209 (N_2209,N_1060,N_28);
or U2210 (N_2210,N_1065,N_95);
xnor U2211 (N_2211,N_490,N_819);
or U2212 (N_2212,N_1049,N_286);
nor U2213 (N_2213,N_273,N_1185);
or U2214 (N_2214,N_506,N_861);
nand U2215 (N_2215,N_747,N_204);
xor U2216 (N_2216,N_150,N_993);
or U2217 (N_2217,N_269,N_1248);
nor U2218 (N_2218,N_981,N_336);
and U2219 (N_2219,N_571,N_598);
and U2220 (N_2220,N_923,N_652);
xor U2221 (N_2221,N_119,N_884);
nor U2222 (N_2222,N_629,N_331);
nor U2223 (N_2223,N_1226,N_282);
nor U2224 (N_2224,N_1174,N_724);
nor U2225 (N_2225,N_933,N_845);
and U2226 (N_2226,N_226,N_659);
or U2227 (N_2227,N_51,N_6);
xor U2228 (N_2228,N_562,N_732);
and U2229 (N_2229,N_673,N_349);
nor U2230 (N_2230,N_765,N_571);
xor U2231 (N_2231,N_782,N_808);
xor U2232 (N_2232,N_1066,N_512);
xnor U2233 (N_2233,N_1082,N_768);
or U2234 (N_2234,N_335,N_202);
nand U2235 (N_2235,N_250,N_313);
or U2236 (N_2236,N_762,N_1074);
or U2237 (N_2237,N_432,N_270);
nand U2238 (N_2238,N_173,N_513);
and U2239 (N_2239,N_152,N_1161);
and U2240 (N_2240,N_1192,N_353);
nand U2241 (N_2241,N_843,N_1061);
nor U2242 (N_2242,N_1015,N_180);
xor U2243 (N_2243,N_1145,N_490);
and U2244 (N_2244,N_1033,N_905);
nor U2245 (N_2245,N_195,N_1006);
xnor U2246 (N_2246,N_214,N_271);
or U2247 (N_2247,N_343,N_852);
and U2248 (N_2248,N_467,N_402);
xor U2249 (N_2249,N_1235,N_824);
or U2250 (N_2250,N_364,N_475);
and U2251 (N_2251,N_896,N_25);
nor U2252 (N_2252,N_653,N_354);
and U2253 (N_2253,N_569,N_175);
nand U2254 (N_2254,N_1194,N_774);
xnor U2255 (N_2255,N_544,N_564);
xnor U2256 (N_2256,N_213,N_89);
or U2257 (N_2257,N_385,N_729);
nor U2258 (N_2258,N_524,N_645);
xor U2259 (N_2259,N_154,N_838);
xor U2260 (N_2260,N_46,N_283);
nor U2261 (N_2261,N_987,N_438);
xnor U2262 (N_2262,N_884,N_553);
xor U2263 (N_2263,N_1069,N_419);
xor U2264 (N_2264,N_1178,N_280);
or U2265 (N_2265,N_767,N_460);
or U2266 (N_2266,N_616,N_632);
and U2267 (N_2267,N_220,N_1059);
xor U2268 (N_2268,N_792,N_779);
nand U2269 (N_2269,N_420,N_975);
nand U2270 (N_2270,N_865,N_503);
nand U2271 (N_2271,N_325,N_248);
and U2272 (N_2272,N_1236,N_1034);
and U2273 (N_2273,N_916,N_718);
and U2274 (N_2274,N_314,N_602);
xor U2275 (N_2275,N_1102,N_367);
and U2276 (N_2276,N_751,N_263);
nand U2277 (N_2277,N_35,N_180);
or U2278 (N_2278,N_689,N_911);
or U2279 (N_2279,N_540,N_763);
or U2280 (N_2280,N_330,N_1118);
or U2281 (N_2281,N_873,N_814);
and U2282 (N_2282,N_630,N_487);
nand U2283 (N_2283,N_887,N_1199);
xnor U2284 (N_2284,N_18,N_764);
or U2285 (N_2285,N_699,N_969);
nor U2286 (N_2286,N_659,N_554);
nand U2287 (N_2287,N_97,N_707);
and U2288 (N_2288,N_490,N_65);
xnor U2289 (N_2289,N_960,N_631);
or U2290 (N_2290,N_840,N_1223);
and U2291 (N_2291,N_381,N_1059);
or U2292 (N_2292,N_596,N_733);
nor U2293 (N_2293,N_1082,N_385);
or U2294 (N_2294,N_404,N_970);
nand U2295 (N_2295,N_305,N_1194);
nor U2296 (N_2296,N_886,N_235);
nor U2297 (N_2297,N_110,N_961);
xor U2298 (N_2298,N_785,N_216);
nor U2299 (N_2299,N_809,N_640);
xor U2300 (N_2300,N_181,N_272);
nand U2301 (N_2301,N_995,N_763);
or U2302 (N_2302,N_1221,N_69);
xnor U2303 (N_2303,N_984,N_314);
nand U2304 (N_2304,N_97,N_1173);
and U2305 (N_2305,N_1245,N_299);
nor U2306 (N_2306,N_994,N_670);
nand U2307 (N_2307,N_723,N_684);
nand U2308 (N_2308,N_842,N_678);
xnor U2309 (N_2309,N_582,N_8);
xor U2310 (N_2310,N_1039,N_1238);
nand U2311 (N_2311,N_314,N_1029);
or U2312 (N_2312,N_1064,N_154);
nand U2313 (N_2313,N_977,N_615);
nand U2314 (N_2314,N_461,N_393);
nand U2315 (N_2315,N_869,N_47);
or U2316 (N_2316,N_780,N_273);
xnor U2317 (N_2317,N_113,N_602);
nor U2318 (N_2318,N_1091,N_590);
nor U2319 (N_2319,N_643,N_333);
or U2320 (N_2320,N_1136,N_1232);
xor U2321 (N_2321,N_682,N_68);
or U2322 (N_2322,N_370,N_62);
nor U2323 (N_2323,N_130,N_296);
or U2324 (N_2324,N_349,N_190);
nor U2325 (N_2325,N_98,N_356);
xnor U2326 (N_2326,N_903,N_790);
xnor U2327 (N_2327,N_762,N_294);
xnor U2328 (N_2328,N_1062,N_1003);
nand U2329 (N_2329,N_805,N_119);
and U2330 (N_2330,N_24,N_491);
and U2331 (N_2331,N_764,N_715);
nand U2332 (N_2332,N_733,N_1230);
nand U2333 (N_2333,N_627,N_855);
xor U2334 (N_2334,N_936,N_154);
nor U2335 (N_2335,N_173,N_1152);
xor U2336 (N_2336,N_1042,N_116);
and U2337 (N_2337,N_597,N_153);
and U2338 (N_2338,N_969,N_290);
nand U2339 (N_2339,N_1067,N_1069);
xor U2340 (N_2340,N_492,N_798);
xnor U2341 (N_2341,N_179,N_273);
or U2342 (N_2342,N_585,N_1132);
and U2343 (N_2343,N_726,N_83);
xor U2344 (N_2344,N_78,N_564);
or U2345 (N_2345,N_789,N_81);
or U2346 (N_2346,N_372,N_327);
nand U2347 (N_2347,N_1241,N_838);
or U2348 (N_2348,N_971,N_1127);
nand U2349 (N_2349,N_907,N_1098);
xnor U2350 (N_2350,N_777,N_830);
nor U2351 (N_2351,N_1247,N_1167);
or U2352 (N_2352,N_326,N_143);
nand U2353 (N_2353,N_215,N_147);
nand U2354 (N_2354,N_491,N_961);
xor U2355 (N_2355,N_398,N_319);
xnor U2356 (N_2356,N_1152,N_333);
nand U2357 (N_2357,N_986,N_76);
nor U2358 (N_2358,N_200,N_295);
or U2359 (N_2359,N_128,N_910);
xor U2360 (N_2360,N_188,N_826);
or U2361 (N_2361,N_439,N_706);
and U2362 (N_2362,N_284,N_1225);
xnor U2363 (N_2363,N_427,N_949);
and U2364 (N_2364,N_23,N_897);
nor U2365 (N_2365,N_26,N_655);
and U2366 (N_2366,N_1049,N_629);
and U2367 (N_2367,N_979,N_1198);
nand U2368 (N_2368,N_147,N_471);
nor U2369 (N_2369,N_746,N_1239);
xnor U2370 (N_2370,N_933,N_372);
and U2371 (N_2371,N_1131,N_231);
nor U2372 (N_2372,N_463,N_583);
nor U2373 (N_2373,N_888,N_1098);
or U2374 (N_2374,N_527,N_665);
xnor U2375 (N_2375,N_872,N_524);
and U2376 (N_2376,N_384,N_97);
or U2377 (N_2377,N_971,N_877);
xnor U2378 (N_2378,N_242,N_302);
nand U2379 (N_2379,N_151,N_394);
xor U2380 (N_2380,N_459,N_168);
nor U2381 (N_2381,N_1084,N_857);
xnor U2382 (N_2382,N_713,N_594);
nor U2383 (N_2383,N_277,N_644);
or U2384 (N_2384,N_255,N_138);
xnor U2385 (N_2385,N_685,N_768);
nor U2386 (N_2386,N_583,N_801);
or U2387 (N_2387,N_1,N_790);
and U2388 (N_2388,N_545,N_235);
and U2389 (N_2389,N_391,N_819);
xnor U2390 (N_2390,N_824,N_615);
and U2391 (N_2391,N_89,N_104);
and U2392 (N_2392,N_413,N_798);
xnor U2393 (N_2393,N_186,N_1035);
and U2394 (N_2394,N_119,N_812);
and U2395 (N_2395,N_404,N_561);
xor U2396 (N_2396,N_668,N_232);
xor U2397 (N_2397,N_953,N_733);
nor U2398 (N_2398,N_249,N_1085);
and U2399 (N_2399,N_155,N_949);
xnor U2400 (N_2400,N_1088,N_1141);
nand U2401 (N_2401,N_177,N_1225);
or U2402 (N_2402,N_239,N_47);
xnor U2403 (N_2403,N_78,N_729);
nand U2404 (N_2404,N_1064,N_523);
nand U2405 (N_2405,N_478,N_627);
or U2406 (N_2406,N_477,N_1122);
xor U2407 (N_2407,N_782,N_919);
or U2408 (N_2408,N_1103,N_1247);
and U2409 (N_2409,N_445,N_1042);
xnor U2410 (N_2410,N_289,N_1185);
nand U2411 (N_2411,N_1080,N_660);
nand U2412 (N_2412,N_1072,N_1078);
or U2413 (N_2413,N_24,N_224);
and U2414 (N_2414,N_195,N_1139);
nor U2415 (N_2415,N_469,N_552);
nor U2416 (N_2416,N_707,N_1159);
or U2417 (N_2417,N_169,N_1018);
or U2418 (N_2418,N_302,N_105);
nand U2419 (N_2419,N_141,N_282);
nor U2420 (N_2420,N_1207,N_662);
or U2421 (N_2421,N_431,N_703);
xor U2422 (N_2422,N_818,N_1094);
or U2423 (N_2423,N_684,N_736);
nand U2424 (N_2424,N_299,N_979);
xor U2425 (N_2425,N_699,N_316);
or U2426 (N_2426,N_1048,N_597);
or U2427 (N_2427,N_1117,N_1159);
and U2428 (N_2428,N_1003,N_1106);
nor U2429 (N_2429,N_1041,N_473);
nor U2430 (N_2430,N_470,N_1090);
xor U2431 (N_2431,N_113,N_748);
or U2432 (N_2432,N_1065,N_122);
nand U2433 (N_2433,N_267,N_1132);
xnor U2434 (N_2434,N_1008,N_474);
xnor U2435 (N_2435,N_996,N_929);
nand U2436 (N_2436,N_79,N_754);
or U2437 (N_2437,N_437,N_700);
nand U2438 (N_2438,N_512,N_468);
nand U2439 (N_2439,N_1137,N_736);
xnor U2440 (N_2440,N_938,N_1012);
or U2441 (N_2441,N_1222,N_96);
or U2442 (N_2442,N_848,N_703);
and U2443 (N_2443,N_41,N_29);
and U2444 (N_2444,N_353,N_535);
nand U2445 (N_2445,N_472,N_924);
nand U2446 (N_2446,N_560,N_1006);
nand U2447 (N_2447,N_480,N_1036);
nand U2448 (N_2448,N_44,N_839);
xor U2449 (N_2449,N_762,N_869);
nor U2450 (N_2450,N_1001,N_355);
and U2451 (N_2451,N_904,N_662);
and U2452 (N_2452,N_349,N_21);
and U2453 (N_2453,N_169,N_554);
xor U2454 (N_2454,N_1079,N_822);
or U2455 (N_2455,N_1058,N_872);
nor U2456 (N_2456,N_1016,N_780);
or U2457 (N_2457,N_838,N_1015);
xor U2458 (N_2458,N_595,N_1229);
and U2459 (N_2459,N_1029,N_1124);
or U2460 (N_2460,N_780,N_636);
or U2461 (N_2461,N_140,N_991);
xor U2462 (N_2462,N_233,N_886);
nand U2463 (N_2463,N_935,N_760);
or U2464 (N_2464,N_30,N_543);
nor U2465 (N_2465,N_115,N_184);
or U2466 (N_2466,N_468,N_1172);
and U2467 (N_2467,N_906,N_440);
xnor U2468 (N_2468,N_717,N_303);
nor U2469 (N_2469,N_1149,N_604);
or U2470 (N_2470,N_158,N_404);
xor U2471 (N_2471,N_988,N_322);
and U2472 (N_2472,N_1170,N_728);
and U2473 (N_2473,N_197,N_1139);
and U2474 (N_2474,N_46,N_1213);
and U2475 (N_2475,N_231,N_724);
or U2476 (N_2476,N_905,N_1216);
xor U2477 (N_2477,N_709,N_639);
xnor U2478 (N_2478,N_1175,N_1124);
xnor U2479 (N_2479,N_1245,N_678);
or U2480 (N_2480,N_584,N_252);
or U2481 (N_2481,N_948,N_59);
and U2482 (N_2482,N_629,N_93);
xnor U2483 (N_2483,N_21,N_641);
and U2484 (N_2484,N_617,N_521);
or U2485 (N_2485,N_615,N_514);
or U2486 (N_2486,N_258,N_240);
nor U2487 (N_2487,N_309,N_733);
nor U2488 (N_2488,N_1225,N_1056);
and U2489 (N_2489,N_110,N_1129);
xor U2490 (N_2490,N_179,N_634);
xor U2491 (N_2491,N_1139,N_706);
and U2492 (N_2492,N_292,N_779);
nand U2493 (N_2493,N_1169,N_785);
and U2494 (N_2494,N_625,N_602);
and U2495 (N_2495,N_362,N_976);
nand U2496 (N_2496,N_761,N_625);
nand U2497 (N_2497,N_292,N_133);
nor U2498 (N_2498,N_898,N_999);
or U2499 (N_2499,N_921,N_673);
nand U2500 (N_2500,N_1647,N_1791);
nor U2501 (N_2501,N_2180,N_1812);
nand U2502 (N_2502,N_1994,N_1585);
nor U2503 (N_2503,N_1792,N_1793);
or U2504 (N_2504,N_2073,N_1680);
xor U2505 (N_2505,N_2388,N_1623);
or U2506 (N_2506,N_1282,N_2197);
nor U2507 (N_2507,N_2306,N_2411);
or U2508 (N_2508,N_2480,N_1526);
and U2509 (N_2509,N_1936,N_2222);
nor U2510 (N_2510,N_1386,N_1930);
xor U2511 (N_2511,N_1993,N_1962);
and U2512 (N_2512,N_1693,N_1504);
nand U2513 (N_2513,N_2498,N_1360);
or U2514 (N_2514,N_1977,N_2391);
or U2515 (N_2515,N_2472,N_1322);
nand U2516 (N_2516,N_1580,N_1445);
or U2517 (N_2517,N_2419,N_1742);
nor U2518 (N_2518,N_2475,N_2333);
and U2519 (N_2519,N_2402,N_1508);
or U2520 (N_2520,N_1345,N_1902);
nor U2521 (N_2521,N_1704,N_1668);
or U2522 (N_2522,N_2154,N_2404);
xnor U2523 (N_2523,N_1667,N_1376);
or U2524 (N_2524,N_1932,N_1860);
nand U2525 (N_2525,N_1357,N_2387);
or U2526 (N_2526,N_1281,N_1428);
and U2527 (N_2527,N_1771,N_1632);
xnor U2528 (N_2528,N_1961,N_1903);
xor U2529 (N_2529,N_2208,N_2228);
xnor U2530 (N_2530,N_2492,N_2272);
nor U2531 (N_2531,N_1291,N_1723);
nand U2532 (N_2532,N_1631,N_1524);
nand U2533 (N_2533,N_1590,N_1583);
nand U2534 (N_2534,N_1456,N_2055);
nand U2535 (N_2535,N_2183,N_1879);
and U2536 (N_2536,N_2079,N_2085);
and U2537 (N_2537,N_2008,N_1724);
or U2538 (N_2538,N_1828,N_1819);
or U2539 (N_2539,N_2230,N_1890);
and U2540 (N_2540,N_2108,N_2372);
nand U2541 (N_2541,N_1467,N_2263);
nor U2542 (N_2542,N_2112,N_1595);
nor U2543 (N_2543,N_2194,N_1774);
nand U2544 (N_2544,N_2395,N_1379);
and U2545 (N_2545,N_1787,N_1306);
xnor U2546 (N_2546,N_2207,N_2407);
xnor U2547 (N_2547,N_2356,N_2458);
nor U2548 (N_2548,N_2470,N_1346);
and U2549 (N_2549,N_2167,N_1769);
or U2550 (N_2550,N_2165,N_1820);
or U2551 (N_2551,N_1556,N_1461);
nor U2552 (N_2552,N_2483,N_1751);
or U2553 (N_2553,N_2429,N_2384);
nor U2554 (N_2554,N_2091,N_2131);
xor U2555 (N_2555,N_1542,N_2126);
nor U2556 (N_2556,N_1454,N_2095);
and U2557 (N_2557,N_1988,N_1719);
nand U2558 (N_2558,N_1528,N_2269);
nor U2559 (N_2559,N_2314,N_2083);
and U2560 (N_2560,N_2030,N_1318);
nor U2561 (N_2561,N_1608,N_2493);
and U2562 (N_2562,N_1672,N_2216);
nand U2563 (N_2563,N_1489,N_2416);
and U2564 (N_2564,N_2206,N_2345);
and U2565 (N_2565,N_2441,N_1460);
nor U2566 (N_2566,N_2186,N_2293);
xor U2567 (N_2567,N_1914,N_2058);
nor U2568 (N_2568,N_2256,N_1601);
xor U2569 (N_2569,N_2425,N_1866);
xnor U2570 (N_2570,N_1929,N_1366);
nand U2571 (N_2571,N_2130,N_1412);
nor U2572 (N_2572,N_1344,N_1314);
and U2573 (N_2573,N_1644,N_1569);
nor U2574 (N_2574,N_1882,N_2427);
nand U2575 (N_2575,N_2336,N_2232);
xor U2576 (N_2576,N_1659,N_1339);
and U2577 (N_2577,N_1926,N_1829);
xor U2578 (N_2578,N_1992,N_2176);
or U2579 (N_2579,N_1759,N_1782);
and U2580 (N_2580,N_2305,N_2067);
xor U2581 (N_2581,N_2264,N_1614);
or U2582 (N_2582,N_1674,N_1514);
and U2583 (N_2583,N_1986,N_1676);
and U2584 (N_2584,N_1835,N_2065);
nor U2585 (N_2585,N_1266,N_1618);
or U2586 (N_2586,N_1352,N_1367);
xnor U2587 (N_2587,N_1840,N_1843);
xnor U2588 (N_2588,N_2036,N_1837);
xnor U2589 (N_2589,N_1698,N_1714);
nand U2590 (N_2590,N_2231,N_2442);
nand U2591 (N_2591,N_1854,N_2147);
xnor U2592 (N_2592,N_1520,N_1482);
or U2593 (N_2593,N_1781,N_1442);
or U2594 (N_2594,N_2409,N_1748);
and U2595 (N_2595,N_1857,N_2171);
nor U2596 (N_2596,N_1688,N_1588);
and U2597 (N_2597,N_2123,N_1721);
or U2598 (N_2598,N_1397,N_2412);
nor U2599 (N_2599,N_1368,N_2196);
and U2600 (N_2600,N_1576,N_1319);
and U2601 (N_2601,N_1378,N_2284);
xor U2602 (N_2602,N_2312,N_1985);
nor U2603 (N_2603,N_1878,N_2109);
nor U2604 (N_2604,N_1708,N_2227);
or U2605 (N_2605,N_2210,N_1931);
nand U2606 (N_2606,N_2444,N_2268);
and U2607 (N_2607,N_2087,N_1853);
nor U2608 (N_2608,N_2371,N_1349);
or U2609 (N_2609,N_1696,N_1701);
nor U2610 (N_2610,N_1395,N_2393);
nor U2611 (N_2611,N_1380,N_1348);
nor U2612 (N_2612,N_2029,N_2178);
or U2613 (N_2613,N_1746,N_2432);
nor U2614 (N_2614,N_1402,N_1800);
xnor U2615 (N_2615,N_1653,N_1868);
nor U2616 (N_2616,N_2344,N_2031);
and U2617 (N_2617,N_1754,N_1681);
nor U2618 (N_2618,N_1565,N_1256);
nand U2619 (N_2619,N_2054,N_1462);
or U2620 (N_2620,N_1921,N_1361);
nor U2621 (N_2621,N_2488,N_1705);
nor U2622 (N_2622,N_2436,N_1833);
nand U2623 (N_2623,N_1944,N_2358);
and U2624 (N_2624,N_2238,N_2459);
and U2625 (N_2625,N_1459,N_2111);
xor U2626 (N_2626,N_1656,N_1838);
xnor U2627 (N_2627,N_1293,N_1609);
xor U2628 (N_2628,N_2082,N_2364);
and U2629 (N_2629,N_1750,N_2383);
xor U2630 (N_2630,N_2330,N_1478);
or U2631 (N_2631,N_1852,N_1369);
nor U2632 (N_2632,N_2190,N_1422);
nor U2633 (N_2633,N_2369,N_1535);
and U2634 (N_2634,N_1738,N_2455);
nand U2635 (N_2635,N_2046,N_2377);
nand U2636 (N_2636,N_2150,N_1578);
nand U2637 (N_2637,N_1959,N_1259);
nand U2638 (N_2638,N_1303,N_1826);
nor U2639 (N_2639,N_2335,N_2355);
and U2640 (N_2640,N_1417,N_2061);
or U2641 (N_2641,N_1285,N_1373);
nor U2642 (N_2642,N_1548,N_1434);
nand U2643 (N_2643,N_1766,N_1315);
nand U2644 (N_2644,N_1734,N_1483);
nor U2645 (N_2645,N_2386,N_1323);
or U2646 (N_2646,N_1262,N_2137);
or U2647 (N_2647,N_2084,N_1779);
xor U2648 (N_2648,N_2205,N_2182);
nor U2649 (N_2649,N_1982,N_2350);
xnor U2650 (N_2650,N_1873,N_1939);
nand U2651 (N_2651,N_2203,N_1896);
and U2652 (N_2652,N_2234,N_1856);
or U2653 (N_2653,N_1399,N_2485);
nor U2654 (N_2654,N_2278,N_2053);
nor U2655 (N_2655,N_2001,N_2466);
nor U2656 (N_2656,N_2349,N_1343);
nand U2657 (N_2657,N_2149,N_2275);
or U2658 (N_2658,N_2144,N_2431);
xnor U2659 (N_2659,N_1855,N_2375);
xor U2660 (N_2660,N_1947,N_1481);
nor U2661 (N_2661,N_2174,N_1711);
and U2662 (N_2662,N_1935,N_1924);
nor U2663 (N_2663,N_2385,N_2357);
and U2664 (N_2664,N_1795,N_1621);
nor U2665 (N_2665,N_1385,N_1446);
or U2666 (N_2666,N_2202,N_2014);
xnor U2667 (N_2667,N_1519,N_1675);
and U2668 (N_2668,N_2456,N_1773);
and U2669 (N_2669,N_2328,N_1671);
xor U2670 (N_2670,N_1269,N_1485);
xor U2671 (N_2671,N_1752,N_1350);
or U2672 (N_2672,N_1332,N_1922);
xor U2673 (N_2673,N_2159,N_2401);
and U2674 (N_2674,N_1404,N_1471);
or U2675 (N_2675,N_1512,N_1786);
xor U2676 (N_2676,N_1398,N_1546);
and U2677 (N_2677,N_1299,N_1995);
or U2678 (N_2678,N_2099,N_1372);
xnor U2679 (N_2679,N_2155,N_1406);
nand U2680 (N_2680,N_2117,N_2451);
or U2681 (N_2681,N_1337,N_2307);
nor U2682 (N_2682,N_2047,N_1611);
nor U2683 (N_2683,N_1640,N_1919);
nand U2684 (N_2684,N_1717,N_2004);
nand U2685 (N_2685,N_1284,N_1770);
or U2686 (N_2686,N_2301,N_2226);
nand U2687 (N_2687,N_1999,N_1745);
and U2688 (N_2688,N_1276,N_2153);
nor U2689 (N_2689,N_1493,N_1405);
nor U2690 (N_2690,N_1606,N_1438);
or U2691 (N_2691,N_1682,N_2019);
nor U2692 (N_2692,N_2469,N_2347);
or U2693 (N_2693,N_2482,N_1305);
nor U2694 (N_2694,N_2465,N_1584);
xnor U2695 (N_2695,N_1265,N_2009);
or U2696 (N_2696,N_2170,N_1775);
xnor U2697 (N_2697,N_1341,N_2070);
nand U2698 (N_2698,N_1517,N_1286);
xnor U2699 (N_2699,N_2360,N_2016);
or U2700 (N_2700,N_2062,N_2020);
and U2701 (N_2701,N_2048,N_2160);
nand U2702 (N_2702,N_1713,N_2434);
nor U2703 (N_2703,N_1666,N_2288);
nor U2704 (N_2704,N_2022,N_2092);
nand U2705 (N_2705,N_2128,N_1987);
and U2706 (N_2706,N_1441,N_2448);
and U2707 (N_2707,N_1863,N_2236);
or U2708 (N_2708,N_1415,N_1927);
xor U2709 (N_2709,N_2365,N_1486);
or U2710 (N_2710,N_2033,N_1885);
nand U2711 (N_2711,N_1946,N_1297);
nand U2712 (N_2712,N_1541,N_1531);
and U2713 (N_2713,N_1788,N_2351);
nand U2714 (N_2714,N_2077,N_1340);
or U2715 (N_2715,N_1252,N_2088);
nand U2716 (N_2716,N_2408,N_1321);
nor U2717 (N_2717,N_1948,N_1908);
nand U2718 (N_2718,N_1883,N_1544);
and U2719 (N_2719,N_1938,N_2418);
xor U2720 (N_2720,N_2038,N_2152);
or U2721 (N_2721,N_1480,N_1311);
nand U2722 (N_2722,N_1661,N_2261);
nand U2723 (N_2723,N_1909,N_2239);
nor U2724 (N_2724,N_1765,N_2221);
nand U2725 (N_2725,N_1831,N_1957);
or U2726 (N_2726,N_2327,N_1448);
and U2727 (N_2727,N_1801,N_1420);
nor U2728 (N_2728,N_2390,N_1612);
nand U2729 (N_2729,N_2027,N_2303);
and U2730 (N_2730,N_1287,N_1848);
nand U2731 (N_2731,N_1970,N_1887);
or U2732 (N_2732,N_1639,N_2243);
and U2733 (N_2733,N_1298,N_1521);
or U2734 (N_2734,N_1642,N_1956);
nand U2735 (N_2735,N_2107,N_2346);
and U2736 (N_2736,N_2495,N_1384);
and U2737 (N_2737,N_1694,N_1657);
xnor U2738 (N_2738,N_1553,N_1491);
or U2739 (N_2739,N_1981,N_1525);
or U2740 (N_2740,N_1824,N_1960);
xor U2741 (N_2741,N_1566,N_2487);
nor U2742 (N_2742,N_2177,N_2248);
or U2743 (N_2743,N_1431,N_2340);
xor U2744 (N_2744,N_2281,N_2075);
nand U2745 (N_2745,N_1974,N_1501);
or U2746 (N_2746,N_2274,N_1679);
nand U2747 (N_2747,N_2074,N_1396);
and U2748 (N_2748,N_1744,N_1457);
and U2749 (N_2749,N_2296,N_2361);
nand U2750 (N_2750,N_2426,N_1300);
nand U2751 (N_2751,N_1643,N_1365);
nand U2752 (N_2752,N_1325,N_1400);
or U2753 (N_2753,N_1383,N_1997);
and U2754 (N_2754,N_1968,N_2025);
nor U2755 (N_2755,N_1953,N_2250);
nand U2756 (N_2756,N_1274,N_2140);
nand U2757 (N_2757,N_1329,N_1530);
and U2758 (N_2758,N_1725,N_1450);
or U2759 (N_2759,N_1624,N_1973);
or U2760 (N_2760,N_2026,N_1390);
or U2761 (N_2761,N_2331,N_2422);
nor U2762 (N_2762,N_1444,N_1880);
or U2763 (N_2763,N_1842,N_2367);
and U2764 (N_2764,N_1413,N_1859);
nor U2765 (N_2765,N_2343,N_2007);
and U2766 (N_2766,N_1338,N_2191);
nand U2767 (N_2767,N_2198,N_1407);
nor U2768 (N_2768,N_1333,N_1280);
and U2769 (N_2769,N_1971,N_2215);
nor U2770 (N_2770,N_2136,N_1753);
nand U2771 (N_2771,N_1794,N_2287);
and U2772 (N_2772,N_1277,N_1364);
or U2773 (N_2773,N_1638,N_1891);
and U2774 (N_2774,N_1394,N_1362);
or U2775 (N_2775,N_1296,N_1712);
or U2776 (N_2776,N_2072,N_1907);
xnor U2777 (N_2777,N_2181,N_1492);
xnor U2778 (N_2778,N_1858,N_2354);
and U2779 (N_2779,N_2114,N_2348);
and U2780 (N_2780,N_1976,N_2220);
and U2781 (N_2781,N_2242,N_1557);
and U2782 (N_2782,N_1628,N_1943);
nor U2783 (N_2783,N_1552,N_1586);
xor U2784 (N_2784,N_2490,N_2260);
xor U2785 (N_2785,N_1496,N_1756);
nand U2786 (N_2786,N_2024,N_1425);
nor U2787 (N_2787,N_1706,N_1509);
nand U2788 (N_2788,N_1302,N_1648);
nand U2789 (N_2789,N_2068,N_2496);
nor U2790 (N_2790,N_2291,N_1822);
or U2791 (N_2791,N_1503,N_1437);
and U2792 (N_2792,N_2478,N_2298);
xor U2793 (N_2793,N_2433,N_1761);
or U2794 (N_2794,N_2173,N_1844);
or U2795 (N_2795,N_1899,N_1874);
and U2796 (N_2796,N_2090,N_1414);
nor U2797 (N_2797,N_2414,N_1802);
and U2798 (N_2798,N_2018,N_1560);
nor U2799 (N_2799,N_2120,N_2449);
and U2800 (N_2800,N_2286,N_1602);
and U2801 (N_2801,N_1660,N_1790);
nand U2802 (N_2802,N_2132,N_2121);
nand U2803 (N_2803,N_1506,N_1727);
nand U2804 (N_2804,N_2104,N_1484);
nand U2805 (N_2805,N_2042,N_2253);
xor U2806 (N_2806,N_1370,N_2057);
nor U2807 (N_2807,N_1772,N_2420);
nand U2808 (N_2808,N_1374,N_1382);
nor U2809 (N_2809,N_2192,N_1529);
and U2810 (N_2810,N_1805,N_2209);
xor U2811 (N_2811,N_2035,N_2059);
nor U2812 (N_2812,N_1600,N_1898);
nor U2813 (N_2813,N_1558,N_2229);
nor U2814 (N_2814,N_1730,N_2211);
nand U2815 (N_2815,N_2311,N_2097);
nor U2816 (N_2816,N_1597,N_1388);
nor U2817 (N_2817,N_1587,N_2134);
xor U2818 (N_2818,N_1283,N_2435);
and U2819 (N_2819,N_1737,N_2225);
nand U2820 (N_2820,N_1598,N_2100);
nor U2821 (N_2821,N_2023,N_1726);
xnor U2822 (N_2822,N_1916,N_2040);
and U2823 (N_2823,N_2223,N_2280);
xor U2824 (N_2824,N_1591,N_1669);
or U2825 (N_2825,N_1409,N_2389);
xnor U2826 (N_2826,N_1377,N_1273);
nand U2827 (N_2827,N_2000,N_1250);
or U2828 (N_2828,N_1707,N_2060);
nand U2829 (N_2829,N_1685,N_1421);
or U2830 (N_2830,N_1267,N_1473);
and U2831 (N_2831,N_1917,N_1499);
or U2832 (N_2832,N_1545,N_1327);
nor U2833 (N_2833,N_2158,N_2244);
and U2834 (N_2834,N_1304,N_2235);
or U2835 (N_2835,N_2184,N_1447);
or U2836 (N_2836,N_1778,N_1443);
nand U2837 (N_2837,N_1523,N_1270);
and U2838 (N_2838,N_1351,N_1633);
xnor U2839 (N_2839,N_2201,N_1980);
or U2840 (N_2840,N_2285,N_1925);
nor U2841 (N_2841,N_1465,N_1923);
and U2842 (N_2842,N_2094,N_2486);
nor U2843 (N_2843,N_1476,N_2166);
xor U2844 (N_2844,N_2076,N_1662);
and U2845 (N_2845,N_1718,N_1964);
nand U2846 (N_2846,N_2370,N_1920);
nor U2847 (N_2847,N_1731,N_2473);
or U2848 (N_2848,N_1469,N_1371);
and U2849 (N_2849,N_1522,N_1911);
nor U2850 (N_2850,N_1949,N_1589);
xor U2851 (N_2851,N_1715,N_1255);
and U2852 (N_2852,N_1452,N_1593);
nand U2853 (N_2853,N_2044,N_2010);
and U2854 (N_2854,N_2450,N_1798);
nor U2855 (N_2855,N_1313,N_1451);
or U2856 (N_2856,N_2172,N_1354);
or U2857 (N_2857,N_2398,N_2359);
nand U2858 (N_2858,N_1955,N_2378);
xor U2859 (N_2859,N_2376,N_2116);
or U2860 (N_2860,N_2056,N_2113);
or U2861 (N_2861,N_2403,N_2168);
nand U2862 (N_2862,N_2457,N_1575);
nor U2863 (N_2863,N_2271,N_2329);
nand U2864 (N_2864,N_2279,N_1747);
and U2865 (N_2865,N_1969,N_1941);
nand U2866 (N_2866,N_1740,N_1776);
nand U2867 (N_2867,N_1881,N_2096);
xnor U2868 (N_2868,N_2479,N_1375);
nor U2869 (N_2869,N_2143,N_2169);
nand U2870 (N_2870,N_1419,N_2017);
nand U2871 (N_2871,N_1780,N_1564);
nor U2872 (N_2872,N_1335,N_2148);
xnor U2873 (N_2873,N_1651,N_1733);
and U2874 (N_2874,N_2462,N_1511);
xnor U2875 (N_2875,N_1806,N_1468);
nand U2876 (N_2876,N_1937,N_1257);
or U2877 (N_2877,N_1827,N_2445);
nor U2878 (N_2878,N_1472,N_1803);
xnor U2879 (N_2879,N_1841,N_1310);
xnor U2880 (N_2880,N_2266,N_1760);
nand U2881 (N_2881,N_1411,N_2497);
xnor U2882 (N_2882,N_2438,N_1905);
or U2883 (N_2883,N_1815,N_1387);
nand U2884 (N_2884,N_1626,N_1475);
nor U2885 (N_2885,N_1889,N_1784);
or U2886 (N_2886,N_1251,N_2300);
and U2887 (N_2887,N_2270,N_2352);
and U2888 (N_2888,N_1427,N_2247);
nand U2889 (N_2889,N_2124,N_1686);
nand U2890 (N_2890,N_1620,N_1573);
and U2891 (N_2891,N_2297,N_1763);
nand U2892 (N_2892,N_1757,N_2163);
nand U2893 (N_2893,N_2437,N_2302);
nand U2894 (N_2894,N_1984,N_2322);
or U2895 (N_2895,N_2325,N_2195);
or U2896 (N_2896,N_2443,N_2259);
or U2897 (N_2897,N_1488,N_1864);
nand U2898 (N_2898,N_1622,N_1507);
xor U2899 (N_2899,N_1670,N_1458);
or U2900 (N_2900,N_1515,N_1886);
and U2901 (N_2901,N_1996,N_2353);
nor U2902 (N_2902,N_1527,N_2454);
and U2903 (N_2903,N_2162,N_2460);
nand U2904 (N_2904,N_1646,N_2115);
and U2905 (N_2905,N_1991,N_2315);
and U2906 (N_2906,N_1677,N_1326);
xor U2907 (N_2907,N_2363,N_2321);
or U2908 (N_2908,N_2039,N_1453);
or U2909 (N_2909,N_1562,N_1804);
and U2910 (N_2910,N_1401,N_1555);
xnor U2911 (N_2911,N_1324,N_1967);
nand U2912 (N_2912,N_2283,N_1690);
or U2913 (N_2913,N_2362,N_1605);
and U2914 (N_2914,N_2368,N_2424);
or U2915 (N_2915,N_1876,N_1449);
and U2916 (N_2916,N_1290,N_2430);
xnor U2917 (N_2917,N_1913,N_2338);
or U2918 (N_2918,N_1741,N_1498);
xor U2919 (N_2919,N_2110,N_1664);
or U2920 (N_2920,N_1629,N_2101);
nand U2921 (N_2921,N_2323,N_1430);
or U2922 (N_2922,N_2006,N_1490);
or U2923 (N_2923,N_2041,N_1732);
and U2924 (N_2924,N_1710,N_1577);
and U2925 (N_2925,N_1764,N_1331);
or U2926 (N_2926,N_1554,N_1716);
nor U2927 (N_2927,N_1836,N_2316);
and U2928 (N_2928,N_2011,N_2217);
and U2929 (N_2929,N_2474,N_1634);
nor U2930 (N_2930,N_2118,N_2453);
nand U2931 (N_2931,N_1933,N_1574);
and U2932 (N_2932,N_1641,N_1813);
and U2933 (N_2933,N_1735,N_1821);
or U2934 (N_2934,N_1872,N_1570);
nand U2935 (N_2935,N_2468,N_1895);
nor U2936 (N_2936,N_2224,N_1301);
or U2937 (N_2937,N_2204,N_2063);
nand U2938 (N_2938,N_2146,N_2415);
nand U2939 (N_2939,N_2089,N_1432);
or U2940 (N_2940,N_1594,N_2374);
or U2941 (N_2941,N_2310,N_1998);
xor U2942 (N_2942,N_2200,N_1495);
or U2943 (N_2943,N_2440,N_1410);
nand U2944 (N_2944,N_1336,N_1513);
or U2945 (N_2945,N_1596,N_1619);
nand U2946 (N_2946,N_1940,N_1785);
nor U2947 (N_2947,N_1307,N_1615);
or U2948 (N_2948,N_1875,N_2255);
or U2949 (N_2949,N_1261,N_1839);
nor U2950 (N_2950,N_1539,N_1900);
or U2951 (N_2951,N_1470,N_1830);
xor U2952 (N_2952,N_1884,N_2381);
and U2953 (N_2953,N_2175,N_1423);
or U2954 (N_2954,N_1692,N_1550);
nor U2955 (N_2955,N_1983,N_2366);
nand U2956 (N_2956,N_2129,N_1536);
nand U2957 (N_2957,N_1264,N_1316);
or U2958 (N_2958,N_1865,N_1572);
or U2959 (N_2959,N_1292,N_1603);
and U2960 (N_2960,N_2463,N_2249);
xnor U2961 (N_2961,N_1559,N_1825);
nor U2962 (N_2962,N_1636,N_1356);
nor U2963 (N_2963,N_2277,N_2103);
xnor U2964 (N_2964,N_2382,N_1695);
nand U2965 (N_2965,N_2218,N_2294);
nor U2966 (N_2966,N_2299,N_1518);
or U2967 (N_2967,N_2105,N_1474);
nor U2968 (N_2968,N_1625,N_2187);
xor U2969 (N_2969,N_1654,N_1607);
nor U2970 (N_2970,N_2037,N_1497);
xor U2971 (N_2971,N_1807,N_1870);
or U2972 (N_2972,N_1652,N_2189);
nor U2973 (N_2973,N_2334,N_2342);
or U2974 (N_2974,N_2125,N_1464);
nand U2975 (N_2975,N_2021,N_1549);
and U2976 (N_2976,N_1347,N_2295);
nor U2977 (N_2977,N_2308,N_2254);
nand U2978 (N_2978,N_1418,N_1455);
and U2979 (N_2979,N_1709,N_1381);
nand U2980 (N_2980,N_1811,N_2258);
nor U2981 (N_2981,N_1436,N_2477);
nor U2982 (N_2982,N_1532,N_2484);
nand U2983 (N_2983,N_1845,N_1571);
and U2984 (N_2984,N_1818,N_2265);
and U2985 (N_2985,N_1439,N_1655);
nor U2986 (N_2986,N_2237,N_2417);
nor U2987 (N_2987,N_1579,N_1547);
or U2988 (N_2988,N_2257,N_1263);
nand U2989 (N_2989,N_1582,N_1278);
and U2990 (N_2990,N_1762,N_1505);
nor U2991 (N_2991,N_1699,N_2127);
nand U2992 (N_2992,N_2161,N_1816);
or U2993 (N_2993,N_1295,N_1834);
or U2994 (N_2994,N_1691,N_2034);
nand U2995 (N_2995,N_1915,N_1799);
nor U2996 (N_2996,N_1862,N_2142);
or U2997 (N_2997,N_1551,N_2476);
or U2998 (N_2998,N_1537,N_1888);
xnor U2999 (N_2999,N_1650,N_2141);
nor U3000 (N_3000,N_1894,N_2003);
nor U3001 (N_3001,N_2326,N_1275);
and U3002 (N_3002,N_2071,N_2396);
nand U3003 (N_3003,N_1975,N_2489);
xnor U3004 (N_3004,N_1649,N_1260);
and U3005 (N_3005,N_2423,N_1663);
or U3006 (N_3006,N_1288,N_1627);
or U3007 (N_3007,N_1989,N_1990);
xnor U3008 (N_3008,N_1877,N_1477);
xor U3009 (N_3009,N_1403,N_1810);
xor U3010 (N_3010,N_2421,N_1934);
nor U3011 (N_3011,N_1678,N_1392);
and U3012 (N_3012,N_2317,N_1645);
and U3013 (N_3013,N_1950,N_1966);
and U3014 (N_3014,N_1703,N_1893);
nand U3015 (N_3015,N_1683,N_1687);
or U3016 (N_3016,N_2012,N_1567);
and U3017 (N_3017,N_2282,N_1728);
nand U3018 (N_3018,N_1809,N_2133);
or U3019 (N_3019,N_1796,N_1722);
nand U3020 (N_3020,N_2313,N_1945);
and U3021 (N_3021,N_2332,N_2106);
nand U3022 (N_3022,N_1563,N_1466);
and U3023 (N_3023,N_1393,N_2319);
or U3024 (N_3024,N_1617,N_1429);
xnor U3025 (N_3025,N_2499,N_1391);
or U3026 (N_3026,N_2494,N_1906);
and U3027 (N_3027,N_2098,N_1673);
and U3028 (N_3028,N_1630,N_2273);
or U3029 (N_3029,N_2119,N_2394);
or U3030 (N_3030,N_1342,N_1253);
or U3031 (N_3031,N_1814,N_1808);
or U3032 (N_3032,N_2078,N_1684);
and U3033 (N_3033,N_1777,N_2481);
nand U3034 (N_3034,N_1353,N_1317);
nor U3035 (N_3035,N_2428,N_1637);
and U3036 (N_3036,N_1979,N_1308);
and U3037 (N_3037,N_1330,N_2439);
nand U3038 (N_3038,N_1942,N_2309);
xnor U3039 (N_3039,N_2043,N_1592);
nor U3040 (N_3040,N_1254,N_1869);
and U3041 (N_3041,N_2002,N_1736);
and U3042 (N_3042,N_2413,N_1416);
nor U3043 (N_3043,N_1268,N_2452);
and U3044 (N_3044,N_1823,N_2320);
nand U3045 (N_3045,N_2213,N_1952);
and U3046 (N_3046,N_1540,N_1904);
and U3047 (N_3047,N_1847,N_2064);
xor U3048 (N_3048,N_1892,N_2289);
nor U3049 (N_3049,N_1604,N_1568);
or U3050 (N_3050,N_1279,N_2185);
nand U3051 (N_3051,N_2135,N_2397);
and U3052 (N_3052,N_1861,N_2015);
and U3053 (N_3053,N_2373,N_1320);
nor U3054 (N_3054,N_2156,N_1897);
nand U3055 (N_3055,N_1487,N_1665);
or U3056 (N_3056,N_1312,N_1720);
nand U3057 (N_3057,N_1363,N_2267);
xor U3058 (N_3058,N_1702,N_2193);
nor U3059 (N_3059,N_1328,N_2049);
and U3060 (N_3060,N_2262,N_1258);
or U3061 (N_3061,N_1440,N_1758);
and U3062 (N_3062,N_2446,N_2122);
xor U3063 (N_3063,N_1817,N_1697);
xnor U3064 (N_3064,N_1768,N_1789);
or U3065 (N_3065,N_2179,N_2157);
and U3066 (N_3066,N_2052,N_2410);
xor U3067 (N_3067,N_2139,N_1435);
xor U3068 (N_3068,N_1972,N_2246);
and U3069 (N_3069,N_1951,N_2086);
nor U3070 (N_3070,N_1309,N_1850);
xor U3071 (N_3071,N_1534,N_2045);
nand U3072 (N_3072,N_1516,N_1846);
and U3073 (N_3073,N_2145,N_1928);
nand U3074 (N_3074,N_1610,N_2252);
xnor U3075 (N_3075,N_1494,N_2290);
nor U3076 (N_3076,N_2324,N_2051);
or U3077 (N_3077,N_2339,N_2405);
nand U3078 (N_3078,N_1359,N_1749);
nand U3079 (N_3079,N_1755,N_1867);
nand U3080 (N_3080,N_1797,N_1832);
nand U3081 (N_3081,N_2245,N_2251);
and U3082 (N_3082,N_1561,N_1901);
or U3083 (N_3083,N_1533,N_1294);
xor U3084 (N_3084,N_2406,N_1851);
nor U3085 (N_3085,N_1963,N_1739);
nor U3086 (N_3086,N_2304,N_1271);
and U3087 (N_3087,N_2212,N_1910);
or U3088 (N_3088,N_2400,N_2318);
nor U3089 (N_3089,N_2188,N_1463);
nand U3090 (N_3090,N_1743,N_2164);
xnor U3091 (N_3091,N_2028,N_2241);
and U3092 (N_3092,N_1978,N_1408);
xnor U3093 (N_3093,N_2341,N_1479);
nor U3094 (N_3094,N_1599,N_1289);
nand U3095 (N_3095,N_1389,N_1355);
and U3096 (N_3096,N_2069,N_1510);
xnor U3097 (N_3097,N_2467,N_2080);
and U3098 (N_3098,N_2471,N_2461);
or U3099 (N_3099,N_1581,N_1767);
xnor U3100 (N_3100,N_2102,N_1658);
nor U3101 (N_3101,N_2276,N_1729);
xnor U3102 (N_3102,N_1635,N_2447);
nand U3103 (N_3103,N_2050,N_1426);
nor U3104 (N_3104,N_1543,N_2392);
xnor U3105 (N_3105,N_1849,N_1700);
and U3106 (N_3106,N_1958,N_2138);
or U3107 (N_3107,N_1613,N_2491);
xor U3108 (N_3108,N_2214,N_1502);
or U3109 (N_3109,N_2240,N_2399);
and U3110 (N_3110,N_2292,N_2081);
or U3111 (N_3111,N_1358,N_1334);
nand U3112 (N_3112,N_1272,N_2464);
or U3113 (N_3113,N_1433,N_2013);
and U3114 (N_3114,N_1616,N_1965);
or U3115 (N_3115,N_2066,N_2151);
xor U3116 (N_3116,N_1500,N_2219);
nand U3117 (N_3117,N_2199,N_2379);
or U3118 (N_3118,N_1912,N_2337);
or U3119 (N_3119,N_1954,N_2380);
or U3120 (N_3120,N_1918,N_1871);
xnor U3121 (N_3121,N_1783,N_1424);
xnor U3122 (N_3122,N_2032,N_2005);
or U3123 (N_3123,N_2093,N_1689);
xor U3124 (N_3124,N_1538,N_2233);
nor U3125 (N_3125,N_2215,N_2211);
xor U3126 (N_3126,N_1414,N_1635);
or U3127 (N_3127,N_2428,N_1386);
xnor U3128 (N_3128,N_1969,N_1732);
and U3129 (N_3129,N_1847,N_1290);
nor U3130 (N_3130,N_1341,N_1679);
nand U3131 (N_3131,N_2453,N_2376);
or U3132 (N_3132,N_2275,N_1541);
xnor U3133 (N_3133,N_1514,N_1692);
nor U3134 (N_3134,N_1859,N_1520);
nor U3135 (N_3135,N_2138,N_2014);
nor U3136 (N_3136,N_2137,N_1294);
or U3137 (N_3137,N_1756,N_1976);
or U3138 (N_3138,N_2279,N_2000);
xnor U3139 (N_3139,N_1612,N_1359);
xnor U3140 (N_3140,N_2376,N_1632);
and U3141 (N_3141,N_2112,N_1335);
nand U3142 (N_3142,N_1930,N_2255);
and U3143 (N_3143,N_1375,N_1886);
or U3144 (N_3144,N_1976,N_1863);
nand U3145 (N_3145,N_1558,N_2220);
or U3146 (N_3146,N_1387,N_1852);
or U3147 (N_3147,N_1361,N_2437);
or U3148 (N_3148,N_1509,N_2336);
and U3149 (N_3149,N_1527,N_1865);
nand U3150 (N_3150,N_1711,N_1978);
nand U3151 (N_3151,N_2453,N_2367);
nor U3152 (N_3152,N_2372,N_1405);
nor U3153 (N_3153,N_2350,N_1254);
nand U3154 (N_3154,N_2001,N_1992);
or U3155 (N_3155,N_2107,N_2281);
xor U3156 (N_3156,N_1647,N_1883);
and U3157 (N_3157,N_1682,N_2351);
and U3158 (N_3158,N_1788,N_1949);
or U3159 (N_3159,N_1896,N_1500);
and U3160 (N_3160,N_2077,N_1573);
nand U3161 (N_3161,N_2054,N_2020);
nand U3162 (N_3162,N_2412,N_1349);
or U3163 (N_3163,N_1914,N_1684);
nor U3164 (N_3164,N_1654,N_1960);
and U3165 (N_3165,N_1390,N_1887);
or U3166 (N_3166,N_2415,N_1842);
or U3167 (N_3167,N_1319,N_2015);
nor U3168 (N_3168,N_1559,N_1481);
and U3169 (N_3169,N_1290,N_2490);
and U3170 (N_3170,N_2185,N_2146);
xor U3171 (N_3171,N_1329,N_2081);
or U3172 (N_3172,N_1252,N_2155);
nand U3173 (N_3173,N_2012,N_1704);
or U3174 (N_3174,N_2302,N_2157);
or U3175 (N_3175,N_1485,N_2003);
nand U3176 (N_3176,N_2051,N_2423);
and U3177 (N_3177,N_2206,N_2012);
and U3178 (N_3178,N_1660,N_2130);
xor U3179 (N_3179,N_1325,N_1963);
xnor U3180 (N_3180,N_2369,N_1807);
nand U3181 (N_3181,N_1556,N_2395);
and U3182 (N_3182,N_1812,N_1472);
xnor U3183 (N_3183,N_1806,N_1997);
or U3184 (N_3184,N_2376,N_1967);
xnor U3185 (N_3185,N_1494,N_2453);
or U3186 (N_3186,N_1379,N_2033);
xor U3187 (N_3187,N_1840,N_2313);
xnor U3188 (N_3188,N_2375,N_2012);
xor U3189 (N_3189,N_1562,N_1293);
nand U3190 (N_3190,N_2483,N_1592);
xnor U3191 (N_3191,N_1999,N_2068);
xor U3192 (N_3192,N_1378,N_1582);
nand U3193 (N_3193,N_1394,N_2176);
or U3194 (N_3194,N_1432,N_2078);
or U3195 (N_3195,N_1313,N_1261);
nand U3196 (N_3196,N_1411,N_2220);
and U3197 (N_3197,N_1587,N_2458);
and U3198 (N_3198,N_2126,N_1583);
or U3199 (N_3199,N_1836,N_1876);
nor U3200 (N_3200,N_2144,N_1376);
or U3201 (N_3201,N_2137,N_1970);
nand U3202 (N_3202,N_1643,N_1766);
and U3203 (N_3203,N_1749,N_1971);
nor U3204 (N_3204,N_2061,N_1654);
xnor U3205 (N_3205,N_1343,N_2281);
xnor U3206 (N_3206,N_2469,N_1590);
and U3207 (N_3207,N_2075,N_2307);
and U3208 (N_3208,N_1376,N_1857);
nor U3209 (N_3209,N_2318,N_1812);
nand U3210 (N_3210,N_1994,N_1993);
or U3211 (N_3211,N_1641,N_1882);
or U3212 (N_3212,N_1711,N_2347);
and U3213 (N_3213,N_1703,N_1686);
and U3214 (N_3214,N_1582,N_1752);
and U3215 (N_3215,N_2062,N_1714);
xor U3216 (N_3216,N_1361,N_2338);
and U3217 (N_3217,N_1421,N_2012);
xor U3218 (N_3218,N_2154,N_1746);
xnor U3219 (N_3219,N_1699,N_2049);
nor U3220 (N_3220,N_1277,N_2172);
nor U3221 (N_3221,N_1436,N_1301);
nor U3222 (N_3222,N_1598,N_1390);
and U3223 (N_3223,N_1940,N_2028);
nor U3224 (N_3224,N_1563,N_1281);
nor U3225 (N_3225,N_2104,N_2286);
or U3226 (N_3226,N_1574,N_2415);
nor U3227 (N_3227,N_1253,N_1839);
xnor U3228 (N_3228,N_2225,N_2065);
and U3229 (N_3229,N_1499,N_1760);
xnor U3230 (N_3230,N_1521,N_1420);
nor U3231 (N_3231,N_2066,N_2453);
nor U3232 (N_3232,N_1927,N_1571);
nor U3233 (N_3233,N_1564,N_2344);
nand U3234 (N_3234,N_2146,N_1420);
nor U3235 (N_3235,N_2397,N_1992);
and U3236 (N_3236,N_1959,N_2258);
nor U3237 (N_3237,N_1609,N_2148);
or U3238 (N_3238,N_1670,N_2105);
and U3239 (N_3239,N_2054,N_1514);
nor U3240 (N_3240,N_1770,N_1709);
xor U3241 (N_3241,N_2003,N_2089);
nand U3242 (N_3242,N_1351,N_1536);
xor U3243 (N_3243,N_1926,N_1334);
or U3244 (N_3244,N_1678,N_2315);
or U3245 (N_3245,N_2087,N_1640);
or U3246 (N_3246,N_2483,N_1632);
and U3247 (N_3247,N_2029,N_1953);
nand U3248 (N_3248,N_1599,N_2321);
or U3249 (N_3249,N_2139,N_2167);
or U3250 (N_3250,N_1401,N_1724);
or U3251 (N_3251,N_1349,N_2410);
nand U3252 (N_3252,N_1590,N_1316);
xnor U3253 (N_3253,N_2214,N_1333);
nor U3254 (N_3254,N_1276,N_2331);
nand U3255 (N_3255,N_2456,N_1319);
nor U3256 (N_3256,N_2280,N_1734);
xor U3257 (N_3257,N_1976,N_1616);
xor U3258 (N_3258,N_2066,N_1747);
nand U3259 (N_3259,N_2078,N_2069);
nor U3260 (N_3260,N_1555,N_2102);
nand U3261 (N_3261,N_1387,N_1684);
nor U3262 (N_3262,N_1587,N_1529);
xor U3263 (N_3263,N_1643,N_1882);
or U3264 (N_3264,N_1563,N_1300);
xnor U3265 (N_3265,N_2118,N_1601);
nand U3266 (N_3266,N_1424,N_1337);
or U3267 (N_3267,N_1466,N_1295);
nor U3268 (N_3268,N_1938,N_2491);
nor U3269 (N_3269,N_2034,N_2081);
nor U3270 (N_3270,N_2036,N_1863);
and U3271 (N_3271,N_1681,N_2041);
xor U3272 (N_3272,N_1949,N_2155);
and U3273 (N_3273,N_2108,N_2454);
and U3274 (N_3274,N_1694,N_1413);
nor U3275 (N_3275,N_1780,N_1343);
nor U3276 (N_3276,N_2374,N_1481);
and U3277 (N_3277,N_1806,N_2280);
nor U3278 (N_3278,N_1870,N_1862);
xnor U3279 (N_3279,N_2226,N_2362);
or U3280 (N_3280,N_1854,N_2146);
or U3281 (N_3281,N_1507,N_2396);
and U3282 (N_3282,N_2258,N_1325);
and U3283 (N_3283,N_2426,N_2274);
xor U3284 (N_3284,N_1825,N_1732);
nor U3285 (N_3285,N_2378,N_1457);
or U3286 (N_3286,N_1818,N_2361);
nor U3287 (N_3287,N_1489,N_1709);
xnor U3288 (N_3288,N_1282,N_2324);
xor U3289 (N_3289,N_2058,N_1343);
and U3290 (N_3290,N_1551,N_2439);
nor U3291 (N_3291,N_1794,N_2471);
or U3292 (N_3292,N_1601,N_1914);
nor U3293 (N_3293,N_1623,N_1842);
nor U3294 (N_3294,N_1705,N_1513);
nand U3295 (N_3295,N_2145,N_2334);
nor U3296 (N_3296,N_2264,N_1384);
nand U3297 (N_3297,N_2061,N_1944);
nand U3298 (N_3298,N_1668,N_1672);
xor U3299 (N_3299,N_2087,N_1961);
and U3300 (N_3300,N_1342,N_2140);
or U3301 (N_3301,N_1335,N_1268);
or U3302 (N_3302,N_1355,N_1754);
or U3303 (N_3303,N_1542,N_1629);
and U3304 (N_3304,N_1312,N_1964);
nor U3305 (N_3305,N_1394,N_1259);
xnor U3306 (N_3306,N_1626,N_1551);
xor U3307 (N_3307,N_2075,N_2152);
or U3308 (N_3308,N_1869,N_2004);
and U3309 (N_3309,N_2384,N_2368);
nor U3310 (N_3310,N_2163,N_1394);
xor U3311 (N_3311,N_2444,N_1690);
or U3312 (N_3312,N_2491,N_1888);
nor U3313 (N_3313,N_2184,N_1395);
or U3314 (N_3314,N_1892,N_1351);
nand U3315 (N_3315,N_2024,N_2040);
nor U3316 (N_3316,N_1475,N_1545);
nor U3317 (N_3317,N_2297,N_1407);
nand U3318 (N_3318,N_1301,N_2280);
nor U3319 (N_3319,N_1407,N_1706);
xor U3320 (N_3320,N_1673,N_2434);
or U3321 (N_3321,N_2437,N_1446);
and U3322 (N_3322,N_2423,N_1903);
and U3323 (N_3323,N_1956,N_1975);
and U3324 (N_3324,N_1318,N_1690);
and U3325 (N_3325,N_2346,N_1815);
or U3326 (N_3326,N_2394,N_2227);
and U3327 (N_3327,N_1742,N_2407);
and U3328 (N_3328,N_2162,N_2271);
and U3329 (N_3329,N_1437,N_2455);
nand U3330 (N_3330,N_2159,N_1657);
nand U3331 (N_3331,N_2384,N_2198);
nand U3332 (N_3332,N_1252,N_1744);
nor U3333 (N_3333,N_2362,N_1876);
xnor U3334 (N_3334,N_1473,N_2104);
and U3335 (N_3335,N_2008,N_2148);
and U3336 (N_3336,N_1850,N_1439);
or U3337 (N_3337,N_2434,N_2261);
or U3338 (N_3338,N_1509,N_1535);
or U3339 (N_3339,N_1489,N_1559);
nand U3340 (N_3340,N_2336,N_2227);
xnor U3341 (N_3341,N_1849,N_2067);
and U3342 (N_3342,N_1883,N_2457);
xor U3343 (N_3343,N_1563,N_1390);
nand U3344 (N_3344,N_2188,N_2486);
xnor U3345 (N_3345,N_2097,N_1896);
nand U3346 (N_3346,N_1869,N_1560);
or U3347 (N_3347,N_1787,N_2413);
nand U3348 (N_3348,N_1667,N_1636);
nor U3349 (N_3349,N_1824,N_1678);
nand U3350 (N_3350,N_2421,N_2216);
xnor U3351 (N_3351,N_1731,N_2448);
and U3352 (N_3352,N_1440,N_1415);
nor U3353 (N_3353,N_1294,N_2290);
nor U3354 (N_3354,N_1350,N_2407);
nand U3355 (N_3355,N_1606,N_1511);
nand U3356 (N_3356,N_1271,N_2029);
and U3357 (N_3357,N_2200,N_1357);
nor U3358 (N_3358,N_1501,N_1292);
nand U3359 (N_3359,N_2313,N_2041);
nand U3360 (N_3360,N_2368,N_1897);
nor U3361 (N_3361,N_1954,N_1554);
xnor U3362 (N_3362,N_1786,N_2199);
xor U3363 (N_3363,N_1662,N_1622);
or U3364 (N_3364,N_2321,N_2243);
or U3365 (N_3365,N_1388,N_1472);
nor U3366 (N_3366,N_2229,N_1872);
or U3367 (N_3367,N_1326,N_2004);
xnor U3368 (N_3368,N_1672,N_1379);
xnor U3369 (N_3369,N_1881,N_2047);
nor U3370 (N_3370,N_2367,N_1907);
xnor U3371 (N_3371,N_2049,N_2396);
nand U3372 (N_3372,N_1719,N_1880);
nor U3373 (N_3373,N_2261,N_1467);
or U3374 (N_3374,N_2222,N_1714);
or U3375 (N_3375,N_1506,N_2492);
nand U3376 (N_3376,N_1393,N_2267);
nor U3377 (N_3377,N_2144,N_2299);
nand U3378 (N_3378,N_2279,N_1640);
xnor U3379 (N_3379,N_1785,N_1604);
xor U3380 (N_3380,N_1596,N_1935);
nor U3381 (N_3381,N_1313,N_1814);
and U3382 (N_3382,N_1481,N_2222);
nor U3383 (N_3383,N_1808,N_1403);
nor U3384 (N_3384,N_2072,N_2408);
or U3385 (N_3385,N_2418,N_1611);
xnor U3386 (N_3386,N_1610,N_1401);
xnor U3387 (N_3387,N_1999,N_1547);
nand U3388 (N_3388,N_1922,N_1302);
nor U3389 (N_3389,N_1665,N_1306);
nor U3390 (N_3390,N_2210,N_1723);
and U3391 (N_3391,N_2036,N_1490);
or U3392 (N_3392,N_1637,N_1987);
nand U3393 (N_3393,N_1682,N_2072);
or U3394 (N_3394,N_1987,N_1363);
and U3395 (N_3395,N_1641,N_2394);
nand U3396 (N_3396,N_1643,N_1513);
or U3397 (N_3397,N_1514,N_1581);
and U3398 (N_3398,N_2062,N_1716);
or U3399 (N_3399,N_1617,N_2396);
and U3400 (N_3400,N_1689,N_2040);
nor U3401 (N_3401,N_1309,N_1590);
nor U3402 (N_3402,N_1257,N_1776);
or U3403 (N_3403,N_1480,N_2418);
nor U3404 (N_3404,N_2237,N_1435);
xnor U3405 (N_3405,N_2316,N_2127);
or U3406 (N_3406,N_2014,N_1482);
xnor U3407 (N_3407,N_2327,N_1854);
and U3408 (N_3408,N_1706,N_1383);
nor U3409 (N_3409,N_1580,N_1273);
nor U3410 (N_3410,N_1672,N_1411);
and U3411 (N_3411,N_1589,N_2085);
or U3412 (N_3412,N_1411,N_1912);
nand U3413 (N_3413,N_1525,N_1783);
nand U3414 (N_3414,N_1807,N_2180);
nor U3415 (N_3415,N_2347,N_2499);
nor U3416 (N_3416,N_2328,N_2057);
nor U3417 (N_3417,N_2428,N_2373);
nand U3418 (N_3418,N_2010,N_1276);
nor U3419 (N_3419,N_1409,N_2323);
nand U3420 (N_3420,N_1275,N_1331);
xnor U3421 (N_3421,N_1597,N_2450);
or U3422 (N_3422,N_1462,N_2003);
nor U3423 (N_3423,N_1998,N_2477);
or U3424 (N_3424,N_1593,N_1996);
nand U3425 (N_3425,N_1850,N_1721);
nor U3426 (N_3426,N_1647,N_2497);
or U3427 (N_3427,N_1440,N_1833);
nand U3428 (N_3428,N_2399,N_2076);
and U3429 (N_3429,N_1396,N_1962);
nor U3430 (N_3430,N_2457,N_1656);
nor U3431 (N_3431,N_2061,N_2317);
or U3432 (N_3432,N_1313,N_1654);
nor U3433 (N_3433,N_2377,N_1452);
xnor U3434 (N_3434,N_2416,N_1463);
xnor U3435 (N_3435,N_1735,N_2015);
xnor U3436 (N_3436,N_2242,N_1603);
nand U3437 (N_3437,N_2475,N_2415);
and U3438 (N_3438,N_1841,N_1843);
nor U3439 (N_3439,N_1410,N_2439);
xor U3440 (N_3440,N_2209,N_2013);
or U3441 (N_3441,N_1469,N_2201);
nor U3442 (N_3442,N_1855,N_2067);
nand U3443 (N_3443,N_1432,N_2157);
or U3444 (N_3444,N_1330,N_1971);
nand U3445 (N_3445,N_2336,N_2273);
nor U3446 (N_3446,N_2141,N_2486);
or U3447 (N_3447,N_2314,N_1344);
nor U3448 (N_3448,N_1834,N_1275);
or U3449 (N_3449,N_1822,N_1320);
xor U3450 (N_3450,N_1393,N_1481);
xnor U3451 (N_3451,N_1723,N_1466);
nor U3452 (N_3452,N_1688,N_1602);
nor U3453 (N_3453,N_1670,N_1260);
xnor U3454 (N_3454,N_2039,N_1416);
nand U3455 (N_3455,N_2326,N_2308);
or U3456 (N_3456,N_1372,N_2440);
xnor U3457 (N_3457,N_1846,N_1581);
nand U3458 (N_3458,N_1616,N_2226);
nand U3459 (N_3459,N_2312,N_1919);
or U3460 (N_3460,N_1376,N_2348);
nor U3461 (N_3461,N_1336,N_2075);
and U3462 (N_3462,N_1307,N_1624);
nand U3463 (N_3463,N_2149,N_1606);
xnor U3464 (N_3464,N_2179,N_1803);
xnor U3465 (N_3465,N_1635,N_1693);
and U3466 (N_3466,N_1928,N_1946);
nand U3467 (N_3467,N_1269,N_2081);
or U3468 (N_3468,N_1607,N_1930);
nor U3469 (N_3469,N_1384,N_1403);
nand U3470 (N_3470,N_2160,N_1344);
nor U3471 (N_3471,N_2289,N_1288);
nor U3472 (N_3472,N_2039,N_1974);
nor U3473 (N_3473,N_1683,N_2428);
xnor U3474 (N_3474,N_2148,N_1869);
nor U3475 (N_3475,N_1935,N_2085);
or U3476 (N_3476,N_1739,N_1795);
nand U3477 (N_3477,N_1523,N_1492);
and U3478 (N_3478,N_1857,N_1596);
nor U3479 (N_3479,N_1928,N_1514);
or U3480 (N_3480,N_1966,N_2438);
or U3481 (N_3481,N_1412,N_2495);
nand U3482 (N_3482,N_2447,N_2246);
nor U3483 (N_3483,N_2392,N_1994);
nand U3484 (N_3484,N_1715,N_2397);
and U3485 (N_3485,N_1425,N_2497);
and U3486 (N_3486,N_1419,N_2180);
or U3487 (N_3487,N_1714,N_1305);
xor U3488 (N_3488,N_2236,N_2019);
and U3489 (N_3489,N_1936,N_2114);
or U3490 (N_3490,N_2049,N_1980);
or U3491 (N_3491,N_2437,N_2227);
or U3492 (N_3492,N_1520,N_1568);
xor U3493 (N_3493,N_1250,N_1567);
and U3494 (N_3494,N_1288,N_2484);
nor U3495 (N_3495,N_2046,N_1708);
nand U3496 (N_3496,N_1809,N_1375);
xnor U3497 (N_3497,N_2167,N_2052);
or U3498 (N_3498,N_2424,N_2302);
or U3499 (N_3499,N_2335,N_1348);
and U3500 (N_3500,N_1394,N_1424);
nand U3501 (N_3501,N_2458,N_1684);
or U3502 (N_3502,N_1648,N_1524);
and U3503 (N_3503,N_1351,N_1565);
nand U3504 (N_3504,N_1452,N_1681);
and U3505 (N_3505,N_1634,N_1833);
and U3506 (N_3506,N_2210,N_2271);
nand U3507 (N_3507,N_1758,N_1640);
and U3508 (N_3508,N_1849,N_1526);
and U3509 (N_3509,N_1489,N_2153);
and U3510 (N_3510,N_2119,N_2231);
and U3511 (N_3511,N_1393,N_2411);
nor U3512 (N_3512,N_1588,N_1379);
nand U3513 (N_3513,N_1645,N_2164);
xnor U3514 (N_3514,N_1542,N_2077);
nor U3515 (N_3515,N_1390,N_2173);
or U3516 (N_3516,N_1831,N_1746);
xnor U3517 (N_3517,N_2048,N_2028);
nor U3518 (N_3518,N_1755,N_2237);
xnor U3519 (N_3519,N_1489,N_2085);
or U3520 (N_3520,N_1569,N_1799);
and U3521 (N_3521,N_2203,N_1989);
xnor U3522 (N_3522,N_1712,N_1502);
or U3523 (N_3523,N_2226,N_1641);
xnor U3524 (N_3524,N_2406,N_1385);
xor U3525 (N_3525,N_1278,N_1495);
nand U3526 (N_3526,N_1991,N_2387);
and U3527 (N_3527,N_2354,N_2108);
nor U3528 (N_3528,N_2417,N_2256);
nand U3529 (N_3529,N_2201,N_2048);
or U3530 (N_3530,N_1366,N_1763);
nand U3531 (N_3531,N_1889,N_2242);
nor U3532 (N_3532,N_1772,N_2325);
nor U3533 (N_3533,N_1609,N_2119);
or U3534 (N_3534,N_2179,N_2160);
or U3535 (N_3535,N_1553,N_1331);
or U3536 (N_3536,N_2320,N_2157);
nand U3537 (N_3537,N_2098,N_1401);
or U3538 (N_3538,N_1253,N_1281);
nor U3539 (N_3539,N_1543,N_2318);
xnor U3540 (N_3540,N_1457,N_1821);
or U3541 (N_3541,N_2115,N_1435);
nor U3542 (N_3542,N_2205,N_2001);
or U3543 (N_3543,N_2008,N_2103);
nor U3544 (N_3544,N_2212,N_1824);
nor U3545 (N_3545,N_2447,N_1556);
xor U3546 (N_3546,N_1295,N_1977);
and U3547 (N_3547,N_1850,N_1568);
or U3548 (N_3548,N_2041,N_1649);
xor U3549 (N_3549,N_2267,N_1847);
and U3550 (N_3550,N_1512,N_1641);
xnor U3551 (N_3551,N_1385,N_2007);
xnor U3552 (N_3552,N_1493,N_1835);
nand U3553 (N_3553,N_1359,N_2305);
or U3554 (N_3554,N_1357,N_1347);
xor U3555 (N_3555,N_1476,N_1696);
nor U3556 (N_3556,N_1533,N_1944);
or U3557 (N_3557,N_1441,N_2155);
or U3558 (N_3558,N_2074,N_2354);
nor U3559 (N_3559,N_2306,N_2415);
or U3560 (N_3560,N_2079,N_1370);
xor U3561 (N_3561,N_2494,N_2266);
and U3562 (N_3562,N_1639,N_1560);
nand U3563 (N_3563,N_1716,N_1704);
xnor U3564 (N_3564,N_2181,N_2250);
and U3565 (N_3565,N_1574,N_1517);
and U3566 (N_3566,N_2106,N_2284);
xnor U3567 (N_3567,N_1852,N_1292);
nor U3568 (N_3568,N_2191,N_1821);
or U3569 (N_3569,N_2288,N_2374);
nor U3570 (N_3570,N_1971,N_2461);
or U3571 (N_3571,N_1727,N_2191);
and U3572 (N_3572,N_2291,N_2145);
nand U3573 (N_3573,N_2104,N_2092);
nor U3574 (N_3574,N_1872,N_1919);
nand U3575 (N_3575,N_1343,N_1963);
and U3576 (N_3576,N_2233,N_1389);
xnor U3577 (N_3577,N_2248,N_1421);
nor U3578 (N_3578,N_1670,N_2059);
nand U3579 (N_3579,N_1440,N_2385);
and U3580 (N_3580,N_2062,N_1353);
and U3581 (N_3581,N_2406,N_1571);
or U3582 (N_3582,N_1813,N_2071);
nand U3583 (N_3583,N_2464,N_2236);
and U3584 (N_3584,N_2335,N_2315);
and U3585 (N_3585,N_2025,N_2150);
nor U3586 (N_3586,N_2391,N_1258);
nand U3587 (N_3587,N_2349,N_2449);
nor U3588 (N_3588,N_2414,N_1521);
nor U3589 (N_3589,N_2377,N_2247);
nor U3590 (N_3590,N_2078,N_2358);
and U3591 (N_3591,N_1817,N_2304);
nor U3592 (N_3592,N_2071,N_2293);
or U3593 (N_3593,N_1542,N_1562);
xnor U3594 (N_3594,N_1351,N_1259);
nor U3595 (N_3595,N_1274,N_2299);
and U3596 (N_3596,N_2348,N_2101);
or U3597 (N_3597,N_1420,N_1809);
or U3598 (N_3598,N_2109,N_2081);
nand U3599 (N_3599,N_1252,N_2399);
nand U3600 (N_3600,N_2298,N_1682);
and U3601 (N_3601,N_1951,N_1325);
xnor U3602 (N_3602,N_1517,N_1817);
nor U3603 (N_3603,N_2408,N_2211);
xnor U3604 (N_3604,N_2339,N_1410);
nand U3605 (N_3605,N_1752,N_1620);
nand U3606 (N_3606,N_2491,N_2249);
nor U3607 (N_3607,N_1434,N_1488);
or U3608 (N_3608,N_2243,N_1808);
xnor U3609 (N_3609,N_1639,N_2198);
and U3610 (N_3610,N_1760,N_2338);
nor U3611 (N_3611,N_2427,N_1840);
or U3612 (N_3612,N_1398,N_2366);
or U3613 (N_3613,N_1685,N_1292);
nand U3614 (N_3614,N_2142,N_1904);
nor U3615 (N_3615,N_2445,N_1460);
and U3616 (N_3616,N_2400,N_1868);
and U3617 (N_3617,N_1775,N_1441);
xnor U3618 (N_3618,N_1864,N_2097);
or U3619 (N_3619,N_1650,N_1922);
nand U3620 (N_3620,N_1488,N_1656);
nand U3621 (N_3621,N_1435,N_1645);
xnor U3622 (N_3622,N_2455,N_1549);
nand U3623 (N_3623,N_1334,N_2401);
xor U3624 (N_3624,N_1469,N_2364);
or U3625 (N_3625,N_1459,N_2469);
and U3626 (N_3626,N_1745,N_1962);
or U3627 (N_3627,N_1790,N_2317);
and U3628 (N_3628,N_2083,N_1826);
nand U3629 (N_3629,N_2239,N_1728);
nand U3630 (N_3630,N_1582,N_2424);
nand U3631 (N_3631,N_1949,N_2276);
or U3632 (N_3632,N_1878,N_2210);
and U3633 (N_3633,N_1580,N_2423);
nand U3634 (N_3634,N_1831,N_1333);
and U3635 (N_3635,N_1698,N_2138);
xor U3636 (N_3636,N_1717,N_2297);
or U3637 (N_3637,N_1901,N_1325);
nor U3638 (N_3638,N_1551,N_2191);
nand U3639 (N_3639,N_2194,N_2445);
xor U3640 (N_3640,N_2092,N_1267);
nor U3641 (N_3641,N_1383,N_1922);
nor U3642 (N_3642,N_1816,N_2450);
xnor U3643 (N_3643,N_1431,N_1410);
nor U3644 (N_3644,N_1340,N_1287);
nand U3645 (N_3645,N_1907,N_2083);
nand U3646 (N_3646,N_1990,N_1458);
nand U3647 (N_3647,N_1544,N_1558);
or U3648 (N_3648,N_1803,N_1875);
or U3649 (N_3649,N_2154,N_2304);
or U3650 (N_3650,N_1790,N_1405);
or U3651 (N_3651,N_1962,N_2046);
or U3652 (N_3652,N_1328,N_1873);
nand U3653 (N_3653,N_2376,N_1439);
nand U3654 (N_3654,N_1588,N_1613);
xor U3655 (N_3655,N_1561,N_1464);
nor U3656 (N_3656,N_1786,N_1768);
nor U3657 (N_3657,N_2286,N_2423);
xor U3658 (N_3658,N_1580,N_2480);
nand U3659 (N_3659,N_2310,N_2037);
and U3660 (N_3660,N_2469,N_2479);
and U3661 (N_3661,N_1382,N_2380);
or U3662 (N_3662,N_1791,N_2165);
nand U3663 (N_3663,N_2434,N_2478);
nor U3664 (N_3664,N_2447,N_1652);
xnor U3665 (N_3665,N_2298,N_1698);
nand U3666 (N_3666,N_2423,N_2025);
and U3667 (N_3667,N_1553,N_1679);
xor U3668 (N_3668,N_2122,N_1332);
nor U3669 (N_3669,N_2276,N_1510);
xnor U3670 (N_3670,N_1363,N_2464);
nor U3671 (N_3671,N_1912,N_1530);
nand U3672 (N_3672,N_1266,N_1444);
or U3673 (N_3673,N_1835,N_2222);
and U3674 (N_3674,N_1821,N_1898);
nand U3675 (N_3675,N_1331,N_1708);
or U3676 (N_3676,N_1621,N_1579);
or U3677 (N_3677,N_1419,N_1398);
nand U3678 (N_3678,N_1681,N_1981);
or U3679 (N_3679,N_2192,N_2197);
or U3680 (N_3680,N_1377,N_1999);
or U3681 (N_3681,N_1978,N_2421);
nor U3682 (N_3682,N_1555,N_2398);
nand U3683 (N_3683,N_1964,N_1648);
xor U3684 (N_3684,N_2468,N_2346);
and U3685 (N_3685,N_2124,N_1296);
nand U3686 (N_3686,N_2212,N_1327);
nand U3687 (N_3687,N_1794,N_2199);
xor U3688 (N_3688,N_1326,N_1449);
and U3689 (N_3689,N_2415,N_2119);
nor U3690 (N_3690,N_1795,N_1438);
nor U3691 (N_3691,N_1811,N_2054);
or U3692 (N_3692,N_1463,N_2414);
and U3693 (N_3693,N_2493,N_1885);
nor U3694 (N_3694,N_2378,N_1825);
nor U3695 (N_3695,N_2106,N_1823);
nor U3696 (N_3696,N_1335,N_1564);
or U3697 (N_3697,N_1908,N_1347);
or U3698 (N_3698,N_1981,N_1274);
nor U3699 (N_3699,N_1987,N_1341);
nand U3700 (N_3700,N_1754,N_1674);
and U3701 (N_3701,N_1636,N_2292);
nor U3702 (N_3702,N_2182,N_1584);
nand U3703 (N_3703,N_1606,N_1362);
or U3704 (N_3704,N_1424,N_1841);
or U3705 (N_3705,N_1938,N_1522);
nor U3706 (N_3706,N_2392,N_2258);
nand U3707 (N_3707,N_1466,N_1864);
nand U3708 (N_3708,N_2200,N_1891);
and U3709 (N_3709,N_2002,N_1926);
nand U3710 (N_3710,N_2167,N_1430);
xor U3711 (N_3711,N_2373,N_2143);
nand U3712 (N_3712,N_2195,N_1548);
nor U3713 (N_3713,N_2211,N_1591);
xnor U3714 (N_3714,N_1816,N_1962);
xnor U3715 (N_3715,N_2154,N_1838);
and U3716 (N_3716,N_1616,N_2375);
xor U3717 (N_3717,N_1599,N_2447);
xor U3718 (N_3718,N_1763,N_2397);
nand U3719 (N_3719,N_2128,N_1704);
and U3720 (N_3720,N_1329,N_1405);
xnor U3721 (N_3721,N_1631,N_1468);
nor U3722 (N_3722,N_1868,N_1667);
or U3723 (N_3723,N_1410,N_1587);
or U3724 (N_3724,N_1972,N_2421);
xnor U3725 (N_3725,N_1394,N_1666);
and U3726 (N_3726,N_1885,N_1362);
xor U3727 (N_3727,N_1732,N_1681);
or U3728 (N_3728,N_1449,N_1650);
nand U3729 (N_3729,N_1682,N_2444);
nand U3730 (N_3730,N_2438,N_2291);
xnor U3731 (N_3731,N_1984,N_2360);
nor U3732 (N_3732,N_1437,N_1930);
nand U3733 (N_3733,N_1533,N_1907);
or U3734 (N_3734,N_1913,N_1297);
or U3735 (N_3735,N_2265,N_1599);
or U3736 (N_3736,N_2149,N_2054);
nor U3737 (N_3737,N_2052,N_1579);
or U3738 (N_3738,N_1649,N_1546);
and U3739 (N_3739,N_1614,N_1348);
nor U3740 (N_3740,N_1939,N_2308);
nor U3741 (N_3741,N_1309,N_1643);
nand U3742 (N_3742,N_1915,N_2389);
nand U3743 (N_3743,N_1359,N_1317);
and U3744 (N_3744,N_1953,N_1966);
nor U3745 (N_3745,N_2041,N_1591);
or U3746 (N_3746,N_1929,N_2354);
or U3747 (N_3747,N_1675,N_1265);
or U3748 (N_3748,N_1926,N_2184);
xnor U3749 (N_3749,N_2384,N_1274);
or U3750 (N_3750,N_3749,N_3632);
and U3751 (N_3751,N_3148,N_3318);
xor U3752 (N_3752,N_3619,N_3435);
and U3753 (N_3753,N_3514,N_3053);
nand U3754 (N_3754,N_2870,N_2533);
nor U3755 (N_3755,N_3333,N_2628);
nand U3756 (N_3756,N_2599,N_3693);
and U3757 (N_3757,N_3169,N_2776);
xnor U3758 (N_3758,N_3717,N_2680);
xnor U3759 (N_3759,N_2681,N_2829);
xnor U3760 (N_3760,N_3118,N_3565);
xor U3761 (N_3761,N_3577,N_3414);
nand U3762 (N_3762,N_3358,N_2664);
nand U3763 (N_3763,N_3255,N_3573);
and U3764 (N_3764,N_3697,N_3413);
nand U3765 (N_3765,N_3334,N_3547);
nor U3766 (N_3766,N_2981,N_2661);
or U3767 (N_3767,N_3374,N_3379);
nor U3768 (N_3768,N_3308,N_3683);
nand U3769 (N_3769,N_2750,N_3437);
nand U3770 (N_3770,N_2757,N_2568);
or U3771 (N_3771,N_3409,N_3389);
or U3772 (N_3772,N_2943,N_3668);
or U3773 (N_3773,N_2954,N_3085);
or U3774 (N_3774,N_2920,N_3098);
or U3775 (N_3775,N_2843,N_2748);
nor U3776 (N_3776,N_3171,N_3504);
nor U3777 (N_3777,N_3337,N_2864);
and U3778 (N_3778,N_2835,N_2755);
nor U3779 (N_3779,N_2736,N_3377);
and U3780 (N_3780,N_2553,N_3044);
and U3781 (N_3781,N_2848,N_2907);
nor U3782 (N_3782,N_3142,N_2685);
or U3783 (N_3783,N_3160,N_2955);
nor U3784 (N_3784,N_3572,N_3328);
nand U3785 (N_3785,N_3278,N_2904);
xnor U3786 (N_3786,N_2917,N_2689);
xnor U3787 (N_3787,N_3679,N_2572);
nand U3788 (N_3788,N_3363,N_3542);
and U3789 (N_3789,N_3251,N_2519);
xor U3790 (N_3790,N_2631,N_3299);
or U3791 (N_3791,N_2559,N_3153);
or U3792 (N_3792,N_2765,N_3215);
or U3793 (N_3793,N_3271,N_2851);
and U3794 (N_3794,N_2965,N_2841);
and U3795 (N_3795,N_3604,N_3270);
and U3796 (N_3796,N_3631,N_3360);
xor U3797 (N_3797,N_3686,N_2566);
or U3798 (N_3798,N_2728,N_3638);
xnor U3799 (N_3799,N_3494,N_2550);
and U3800 (N_3800,N_3428,N_3112);
nor U3801 (N_3801,N_3320,N_2675);
or U3802 (N_3802,N_3716,N_3376);
nand U3803 (N_3803,N_2670,N_2871);
or U3804 (N_3804,N_2789,N_2510);
nand U3805 (N_3805,N_2961,N_3558);
nand U3806 (N_3806,N_2665,N_3102);
nor U3807 (N_3807,N_2772,N_3307);
nand U3808 (N_3808,N_3625,N_3141);
or U3809 (N_3809,N_2684,N_3402);
nor U3810 (N_3810,N_2731,N_2515);
nand U3811 (N_3811,N_3730,N_3212);
nor U3812 (N_3812,N_2593,N_2779);
nand U3813 (N_3813,N_3505,N_3474);
nor U3814 (N_3814,N_3605,N_2688);
xnor U3815 (N_3815,N_2601,N_3323);
xnor U3816 (N_3816,N_3512,N_2653);
nand U3817 (N_3817,N_2666,N_2902);
xnor U3818 (N_3818,N_2869,N_2898);
nand U3819 (N_3819,N_3701,N_3450);
and U3820 (N_3820,N_3626,N_2583);
nand U3821 (N_3821,N_3246,N_3436);
and U3822 (N_3822,N_2946,N_3346);
and U3823 (N_3823,N_3419,N_2791);
xnor U3824 (N_3824,N_2878,N_2874);
nor U3825 (N_3825,N_3310,N_2980);
nor U3826 (N_3826,N_2692,N_3609);
nor U3827 (N_3827,N_2913,N_3125);
nor U3828 (N_3828,N_2964,N_3264);
xor U3829 (N_3829,N_3082,N_2872);
or U3830 (N_3830,N_3628,N_3315);
or U3831 (N_3831,N_3015,N_3286);
and U3832 (N_3832,N_3535,N_3690);
nor U3833 (N_3833,N_3362,N_3088);
nor U3834 (N_3834,N_2865,N_3531);
nand U3835 (N_3835,N_3748,N_2635);
and U3836 (N_3836,N_2973,N_3059);
or U3837 (N_3837,N_3208,N_2773);
nand U3838 (N_3838,N_3029,N_2634);
nor U3839 (N_3839,N_3642,N_2682);
and U3840 (N_3840,N_2941,N_3403);
xor U3841 (N_3841,N_3637,N_3735);
nor U3842 (N_3842,N_2861,N_2794);
or U3843 (N_3843,N_3478,N_2839);
nand U3844 (N_3844,N_3273,N_2691);
xor U3845 (N_3845,N_2594,N_3449);
or U3846 (N_3846,N_3266,N_2517);
xor U3847 (N_3847,N_3438,N_3453);
and U3848 (N_3848,N_3464,N_2725);
nor U3849 (N_3849,N_3232,N_3695);
nand U3850 (N_3850,N_3150,N_2900);
nand U3851 (N_3851,N_2641,N_2614);
xnor U3852 (N_3852,N_2774,N_2737);
nand U3853 (N_3853,N_2727,N_3476);
nand U3854 (N_3854,N_3603,N_2534);
nand U3855 (N_3855,N_3726,N_3324);
and U3856 (N_3856,N_2958,N_3424);
or U3857 (N_3857,N_3116,N_2828);
xnor U3858 (N_3858,N_2970,N_3155);
or U3859 (N_3859,N_3483,N_3109);
nand U3860 (N_3860,N_2770,N_2969);
nor U3861 (N_3861,N_3131,N_3025);
nor U3862 (N_3862,N_3124,N_3120);
and U3863 (N_3863,N_2581,N_3222);
xor U3864 (N_3864,N_3496,N_2636);
or U3865 (N_3865,N_3624,N_2922);
xnor U3866 (N_3866,N_3032,N_3151);
and U3867 (N_3867,N_3064,N_2551);
or U3868 (N_3868,N_2524,N_3479);
xor U3869 (N_3869,N_3122,N_2518);
nand U3870 (N_3870,N_2527,N_3465);
and U3871 (N_3871,N_2811,N_2586);
xor U3872 (N_3872,N_3452,N_2645);
nand U3873 (N_3873,N_2542,N_2863);
nand U3874 (N_3874,N_2787,N_3700);
or U3875 (N_3875,N_2856,N_3050);
and U3876 (N_3876,N_2749,N_2901);
or U3877 (N_3877,N_3263,N_3640);
xnor U3878 (N_3878,N_3657,N_3062);
and U3879 (N_3879,N_3630,N_2632);
nor U3880 (N_3880,N_3612,N_3244);
and U3881 (N_3881,N_2968,N_3430);
nor U3882 (N_3882,N_2905,N_2962);
nor U3883 (N_3883,N_3396,N_3119);
or U3884 (N_3884,N_3093,N_2906);
or U3885 (N_3885,N_3506,N_3027);
or U3886 (N_3886,N_2944,N_3095);
and U3887 (N_3887,N_3063,N_3135);
and U3888 (N_3888,N_2712,N_3237);
or U3889 (N_3889,N_3649,N_2948);
or U3890 (N_3890,N_3007,N_3442);
and U3891 (N_3891,N_2529,N_3041);
xnor U3892 (N_3892,N_3530,N_3395);
nand U3893 (N_3893,N_3663,N_3676);
xor U3894 (N_3894,N_2590,N_2929);
nor U3895 (N_3895,N_2805,N_3168);
or U3896 (N_3896,N_3691,N_3257);
or U3897 (N_3897,N_3336,N_2535);
xnor U3898 (N_3898,N_2669,N_3427);
nor U3899 (N_3899,N_2503,N_2889);
and U3900 (N_3900,N_3046,N_3743);
and U3901 (N_3901,N_3342,N_2545);
and U3902 (N_3902,N_2934,N_3585);
nor U3903 (N_3903,N_3529,N_3117);
xor U3904 (N_3904,N_2756,N_3350);
nor U3905 (N_3905,N_2644,N_2814);
or U3906 (N_3906,N_3461,N_2927);
nand U3907 (N_3907,N_3728,N_3267);
nand U3908 (N_3908,N_3037,N_2933);
xnor U3909 (N_3909,N_3580,N_3186);
nor U3910 (N_3910,N_3513,N_2979);
and U3911 (N_3911,N_3378,N_3103);
xnor U3912 (N_3912,N_3740,N_2781);
xor U3913 (N_3913,N_3680,N_3129);
nand U3914 (N_3914,N_3429,N_3347);
nand U3915 (N_3915,N_2960,N_3134);
or U3916 (N_3916,N_3669,N_3367);
and U3917 (N_3917,N_3312,N_2588);
or U3918 (N_3918,N_3172,N_3627);
nor U3919 (N_3919,N_3383,N_2852);
and U3920 (N_3920,N_3105,N_3265);
nor U3921 (N_3921,N_3096,N_2595);
and U3922 (N_3922,N_3592,N_2626);
nand U3923 (N_3923,N_3611,N_2887);
or U3924 (N_3924,N_2678,N_2663);
or U3925 (N_3925,N_2709,N_3739);
xor U3926 (N_3926,N_2826,N_3445);
nor U3927 (N_3927,N_2598,N_2556);
nand U3928 (N_3928,N_2804,N_2806);
nand U3929 (N_3929,N_3720,N_3608);
and U3930 (N_3930,N_3011,N_3195);
or U3931 (N_3931,N_2652,N_3747);
xnor U3932 (N_3932,N_3227,N_3444);
and U3933 (N_3933,N_3144,N_3331);
and U3934 (N_3934,N_2989,N_3285);
or U3935 (N_3935,N_3517,N_3052);
and U3936 (N_3936,N_3238,N_3281);
and U3937 (N_3937,N_2506,N_2813);
nand U3938 (N_3938,N_3311,N_2825);
xnor U3939 (N_3939,N_3301,N_2771);
nand U3940 (N_3940,N_3731,N_3133);
nand U3941 (N_3941,N_2600,N_3723);
and U3942 (N_3942,N_2699,N_3524);
or U3943 (N_3943,N_3028,N_3736);
or U3944 (N_3944,N_2924,N_2734);
xnor U3945 (N_3945,N_3060,N_3578);
nor U3946 (N_3946,N_2650,N_3247);
xnor U3947 (N_3947,N_2660,N_3732);
nor U3948 (N_3948,N_2746,N_3317);
xor U3949 (N_3949,N_3713,N_2592);
nor U3950 (N_3950,N_3040,N_3470);
nand U3951 (N_3951,N_3656,N_2617);
or U3952 (N_3952,N_2679,N_2704);
xor U3953 (N_3953,N_3684,N_2584);
or U3954 (N_3954,N_3741,N_3510);
or U3955 (N_3955,N_3340,N_3399);
xnor U3956 (N_3956,N_3365,N_3545);
and U3957 (N_3957,N_2834,N_3493);
xnor U3958 (N_3958,N_3368,N_3551);
xor U3959 (N_3959,N_2821,N_3468);
nand U3960 (N_3960,N_3463,N_2705);
or U3961 (N_3961,N_2502,N_3228);
nand U3962 (N_3962,N_3454,N_3645);
nor U3963 (N_3963,N_3652,N_2655);
nand U3964 (N_3964,N_2802,N_3154);
or U3965 (N_3965,N_3552,N_3157);
xnor U3966 (N_3966,N_3045,N_3180);
nand U3967 (N_3967,N_2953,N_3137);
nor U3968 (N_3968,N_3282,N_2988);
nor U3969 (N_3969,N_3048,N_2701);
xor U3970 (N_3970,N_3138,N_2719);
nand U3971 (N_3971,N_3556,N_2571);
or U3972 (N_3972,N_3440,N_3650);
xnor U3973 (N_3973,N_2860,N_2511);
nand U3974 (N_3974,N_3502,N_2676);
xor U3975 (N_3975,N_3594,N_3108);
nor U3976 (N_3976,N_3372,N_3256);
nor U3977 (N_3977,N_3325,N_3644);
nor U3978 (N_3978,N_2622,N_3576);
and U3979 (N_3979,N_3224,N_3600);
xnor U3980 (N_3980,N_3375,N_3006);
or U3981 (N_3981,N_3036,N_3049);
nor U3982 (N_3982,N_3667,N_3192);
and U3983 (N_3983,N_3262,N_3618);
nand U3984 (N_3984,N_3021,N_3184);
nor U3985 (N_3985,N_3236,N_3393);
and U3986 (N_3986,N_3229,N_3745);
and U3987 (N_3987,N_3417,N_2591);
and U3988 (N_3988,N_3100,N_3167);
xor U3989 (N_3989,N_3182,N_3537);
or U3990 (N_3990,N_2623,N_2858);
xor U3991 (N_3991,N_2947,N_3269);
nor U3992 (N_3992,N_2763,N_3639);
nand U3993 (N_3993,N_2531,N_3658);
nor U3994 (N_3994,N_3054,N_3415);
nor U3995 (N_3995,N_2850,N_3487);
xor U3996 (N_3996,N_3010,N_2647);
nand U3997 (N_3997,N_3018,N_3410);
and U3998 (N_3998,N_3023,N_3712);
xnor U3999 (N_3999,N_2768,N_3614);
and U4000 (N_4000,N_2866,N_3164);
nand U4001 (N_4001,N_3326,N_3140);
nand U4002 (N_4002,N_2868,N_2708);
nor U4003 (N_4003,N_3560,N_3073);
nor U4004 (N_4004,N_2662,N_3290);
nand U4005 (N_4005,N_3406,N_3303);
nand U4006 (N_4006,N_3643,N_2937);
nor U4007 (N_4007,N_3139,N_2761);
xnor U4008 (N_4008,N_2996,N_3707);
xor U4009 (N_4009,N_3152,N_3615);
and U4010 (N_4010,N_2579,N_2615);
xnor U4011 (N_4011,N_3400,N_3293);
or U4012 (N_4012,N_3589,N_2743);
nand U4013 (N_4013,N_3200,N_3727);
and U4014 (N_4014,N_3484,N_2607);
and U4015 (N_4015,N_2546,N_3536);
or U4016 (N_4016,N_3356,N_3724);
nand U4017 (N_4017,N_3617,N_2677);
xnor U4018 (N_4018,N_2544,N_2564);
and U4019 (N_4019,N_2730,N_2891);
xor U4020 (N_4020,N_3515,N_2877);
nor U4021 (N_4021,N_2543,N_3574);
nand U4022 (N_4022,N_2683,N_2561);
or U4023 (N_4023,N_2882,N_3466);
and U4024 (N_4024,N_3191,N_2720);
nor U4025 (N_4025,N_2694,N_2831);
nand U4026 (N_4026,N_2792,N_3111);
or U4027 (N_4027,N_3194,N_2908);
nor U4028 (N_4028,N_3481,N_2508);
or U4029 (N_4029,N_3132,N_3128);
or U4030 (N_4030,N_2714,N_2798);
nor U4031 (N_4031,N_3366,N_2603);
xor U4032 (N_4032,N_2642,N_3621);
xor U4033 (N_4033,N_2610,N_2690);
xor U4034 (N_4034,N_2706,N_3653);
nand U4035 (N_4035,N_3391,N_3682);
and U4036 (N_4036,N_2778,N_3145);
xor U4037 (N_4037,N_3526,N_3404);
nand U4038 (N_4038,N_2523,N_2587);
or U4039 (N_4039,N_2646,N_3104);
nor U4040 (N_4040,N_2643,N_2633);
nor U4041 (N_4041,N_2926,N_3685);
nand U4042 (N_4042,N_2818,N_2513);
nand U4043 (N_4043,N_2975,N_2711);
or U4044 (N_4044,N_3534,N_3457);
and U4045 (N_4045,N_3380,N_3401);
nor U4046 (N_4046,N_2911,N_2606);
nand U4047 (N_4047,N_2555,N_3659);
nor U4048 (N_4048,N_3209,N_3675);
or U4049 (N_4049,N_3533,N_3586);
nor U4050 (N_4050,N_2541,N_2931);
nor U4051 (N_4051,N_3014,N_2925);
nor U4052 (N_4052,N_3361,N_2759);
xor U4053 (N_4053,N_3024,N_2500);
and U4054 (N_4054,N_3090,N_3408);
and U4055 (N_4055,N_3355,N_2986);
xnor U4056 (N_4056,N_3199,N_3569);
or U4057 (N_4057,N_2824,N_2695);
nand U4058 (N_4058,N_2621,N_3447);
and U4059 (N_4059,N_2796,N_2845);
and U4060 (N_4060,N_2914,N_3179);
xor U4061 (N_4061,N_2918,N_2942);
nor U4062 (N_4062,N_2638,N_3673);
nor U4063 (N_4063,N_3459,N_2659);
xnor U4064 (N_4064,N_2686,N_2580);
nor U4065 (N_4065,N_3189,N_3086);
or U4066 (N_4066,N_3706,N_3268);
or U4067 (N_4067,N_3170,N_3498);
or U4068 (N_4068,N_3008,N_2945);
nand U4069 (N_4069,N_2854,N_3012);
nor U4070 (N_4070,N_3418,N_2974);
xor U4071 (N_4071,N_2612,N_2838);
nor U4072 (N_4072,N_2935,N_3509);
nor U4073 (N_4073,N_3602,N_3338);
nor U4074 (N_4074,N_2745,N_3101);
xnor U4075 (N_4075,N_3259,N_3439);
or U4076 (N_4076,N_3662,N_3348);
or U4077 (N_4077,N_3711,N_2932);
xor U4078 (N_4078,N_3610,N_2987);
xor U4079 (N_4079,N_2896,N_3384);
nor U4080 (N_4080,N_3161,N_3300);
xor U4081 (N_4081,N_3177,N_3477);
or U4082 (N_4082,N_3382,N_3254);
xnor U4083 (N_4083,N_3471,N_3492);
or U4084 (N_4084,N_3291,N_3249);
and U4085 (N_4085,N_3051,N_3715);
and U4086 (N_4086,N_3013,N_2857);
xnor U4087 (N_4087,N_3280,N_2657);
and U4088 (N_4088,N_3423,N_3566);
nor U4089 (N_4089,N_3188,N_3357);
and U4090 (N_4090,N_3176,N_3213);
xor U4091 (N_4091,N_3149,N_3557);
nand U4092 (N_4092,N_3003,N_3369);
or U4093 (N_4093,N_2990,N_3329);
xnor U4094 (N_4094,N_3030,N_3646);
nor U4095 (N_4095,N_2827,N_3147);
or U4096 (N_4096,N_3276,N_2876);
nor U4097 (N_4097,N_3359,N_3033);
and U4098 (N_4098,N_2801,N_2867);
xnor U4099 (N_4099,N_2526,N_2880);
xnor U4100 (N_4100,N_3703,N_2732);
nand U4101 (N_4101,N_3397,N_3539);
or U4102 (N_4102,N_3486,N_3084);
nand U4103 (N_4103,N_3523,N_3070);
xnor U4104 (N_4104,N_2837,N_3113);
or U4105 (N_4105,N_2521,N_3330);
nor U4106 (N_4106,N_3622,N_2971);
or U4107 (N_4107,N_2717,N_2582);
and U4108 (N_4108,N_2799,N_2567);
xor U4109 (N_4109,N_3390,N_3567);
nand U4110 (N_4110,N_3692,N_3211);
nor U4111 (N_4111,N_2554,N_3596);
xnor U4112 (N_4112,N_3345,N_3252);
nor U4113 (N_4113,N_3681,N_3305);
or U4114 (N_4114,N_3598,N_3287);
nor U4115 (N_4115,N_3448,N_3056);
nand U4116 (N_4116,N_3538,N_2505);
nor U4117 (N_4117,N_3599,N_2873);
nand U4118 (N_4118,N_3629,N_3126);
and U4119 (N_4119,N_2884,N_3458);
nand U4120 (N_4120,N_3283,N_3674);
nand U4121 (N_4121,N_3110,N_3080);
xor U4122 (N_4122,N_2977,N_3425);
xnor U4123 (N_4123,N_2991,N_2853);
nor U4124 (N_4124,N_3373,N_3665);
or U4125 (N_4125,N_3107,N_2537);
nand U4126 (N_4126,N_2764,N_3055);
and U4127 (N_4127,N_2618,N_3127);
nor U4128 (N_4128,N_3197,N_3426);
xnor U4129 (N_4129,N_3441,N_2963);
nor U4130 (N_4130,N_3620,N_2895);
xor U4131 (N_4131,N_2672,N_3042);
nand U4132 (N_4132,N_3075,N_3201);
xnor U4133 (N_4133,N_2616,N_2549);
nand U4134 (N_4134,N_3322,N_2978);
xnor U4135 (N_4135,N_3016,N_2984);
xnor U4136 (N_4136,N_3087,N_2995);
xnor U4137 (N_4137,N_2573,N_3544);
xnor U4138 (N_4138,N_3193,N_3136);
xor U4139 (N_4139,N_3022,N_3722);
and U4140 (N_4140,N_3588,N_2909);
nand U4141 (N_4141,N_2687,N_2780);
xor U4142 (N_4142,N_2767,N_3729);
nor U4143 (N_4143,N_3704,N_3295);
nor U4144 (N_4144,N_3233,N_3555);
nor U4145 (N_4145,N_2993,N_3214);
xnor U4146 (N_4146,N_2921,N_3298);
or U4147 (N_4147,N_2693,N_2729);
nor U4148 (N_4148,N_2766,N_3187);
or U4149 (N_4149,N_2985,N_3163);
nand U4150 (N_4150,N_3527,N_3204);
nand U4151 (N_4151,N_2577,N_3623);
xor U4152 (N_4152,N_2639,N_3696);
xnor U4153 (N_4153,N_3079,N_3143);
nand U4154 (N_4154,N_2894,N_2910);
xnor U4155 (N_4155,N_2740,N_2957);
xor U4156 (N_4156,N_2696,N_2883);
nor U4157 (N_4157,N_3443,N_2951);
xor U4158 (N_4158,N_3220,N_2654);
xor U4159 (N_4159,N_3165,N_3198);
nor U4160 (N_4160,N_3114,N_3158);
or U4161 (N_4161,N_3516,N_2574);
nor U4162 (N_4162,N_2528,N_3549);
nor U4163 (N_4163,N_2795,N_3258);
xor U4164 (N_4164,N_2862,N_2578);
nand U4165 (N_4165,N_3035,N_2952);
xnor U4166 (N_4166,N_2552,N_3146);
nand U4167 (N_4167,N_3077,N_2507);
nor U4168 (N_4168,N_2859,N_2668);
nand U4169 (N_4169,N_2760,N_2849);
nor U4170 (N_4170,N_3061,N_3635);
xor U4171 (N_4171,N_3001,N_2999);
xnor U4172 (N_4172,N_3039,N_2620);
and U4173 (N_4173,N_3460,N_2629);
nand U4174 (N_4174,N_3313,N_2823);
or U4175 (N_4175,N_2967,N_3243);
nand U4176 (N_4176,N_2893,N_3304);
and U4177 (N_4177,N_3302,N_3433);
and U4178 (N_4178,N_2777,N_3210);
or U4179 (N_4179,N_2762,N_2548);
and U4180 (N_4180,N_2713,N_2716);
xnor U4181 (N_4181,N_2570,N_3467);
xor U4182 (N_4182,N_2881,N_3421);
xor U4183 (N_4183,N_3388,N_3456);
nor U4184 (N_4184,N_2721,N_3121);
xor U4185 (N_4185,N_3156,N_2788);
nor U4186 (N_4186,N_3687,N_2651);
xnor U4187 (N_4187,N_3570,N_2949);
xnor U4188 (N_4188,N_3123,N_3434);
nor U4189 (N_4189,N_3316,N_3593);
or U4190 (N_4190,N_2994,N_2723);
nand U4191 (N_4191,N_3094,N_3532);
or U4192 (N_4192,N_2936,N_3351);
or U4193 (N_4193,N_3491,N_3097);
and U4194 (N_4194,N_3541,N_2722);
and U4195 (N_4195,N_3175,N_2790);
xor U4196 (N_4196,N_3173,N_2930);
nand U4197 (N_4197,N_2919,N_3528);
or U4198 (N_4198,N_3591,N_3455);
nor U4199 (N_4199,N_2649,N_2613);
and U4200 (N_4200,N_2966,N_3431);
nand U4201 (N_4201,N_2624,N_3564);
nand U4202 (N_4202,N_2782,N_2674);
nand U4203 (N_4203,N_3568,N_3485);
nor U4204 (N_4204,N_2540,N_3522);
or U4205 (N_4205,N_3279,N_3344);
or U4206 (N_4206,N_3451,N_2899);
xor U4207 (N_4207,N_2539,N_3507);
and U4208 (N_4208,N_3065,N_3499);
nor U4209 (N_4209,N_3579,N_2605);
nand U4210 (N_4210,N_2959,N_3385);
and U4211 (N_4211,N_2855,N_3196);
nor U4212 (N_4212,N_3480,N_2892);
or U4213 (N_4213,N_3115,N_3130);
nor U4214 (N_4214,N_3420,N_3332);
xor U4215 (N_4215,N_2888,N_3718);
and U4216 (N_4216,N_3297,N_2915);
xnor U4217 (N_4217,N_3501,N_3206);
or U4218 (N_4218,N_3381,N_3031);
or U4219 (N_4219,N_2673,N_3248);
nor U4220 (N_4220,N_2885,N_3613);
nor U4221 (N_4221,N_2775,N_2800);
xnor U4222 (N_4222,N_3559,N_2563);
nand U4223 (N_4223,N_3482,N_2726);
or U4224 (N_4224,N_2569,N_3708);
or U4225 (N_4225,N_2836,N_3203);
or U4226 (N_4226,N_2982,N_3216);
nand U4227 (N_4227,N_3641,N_3250);
and U4228 (N_4228,N_3699,N_2602);
nand U4229 (N_4229,N_2803,N_3272);
xnor U4230 (N_4230,N_2997,N_3235);
nor U4231 (N_4231,N_3678,N_3540);
xnor U4232 (N_4232,N_3742,N_3289);
nor U4233 (N_4233,N_2753,N_3043);
nor U4234 (N_4234,N_3521,N_3242);
nand U4235 (N_4235,N_2976,N_3071);
or U4236 (N_4236,N_2512,N_3554);
nand U4237 (N_4237,N_2739,N_3074);
nor U4238 (N_4238,N_2560,N_2808);
and U4239 (N_4239,N_2733,N_3190);
nand U4240 (N_4240,N_2608,N_3660);
nand U4241 (N_4241,N_3392,N_3462);
and U4242 (N_4242,N_3553,N_3386);
xnor U4243 (N_4243,N_3546,N_3525);
xnor U4244 (N_4244,N_3671,N_3737);
nand U4245 (N_4245,N_3495,N_3387);
and U4246 (N_4246,N_3277,N_3089);
and U4247 (N_4247,N_3314,N_3019);
nor U4248 (N_4248,N_3672,N_3446);
xor U4249 (N_4249,N_3607,N_3581);
nand U4250 (N_4250,N_2585,N_3370);
xnor U4251 (N_4251,N_2785,N_2816);
xor U4252 (N_4252,N_2807,N_3664);
nand U4253 (N_4253,N_3511,N_3519);
nand U4254 (N_4254,N_3647,N_3719);
nor U4255 (N_4255,N_2627,N_3407);
nand U4256 (N_4256,N_3339,N_2671);
nor U4257 (N_4257,N_2702,N_2847);
nor U4258 (N_4258,N_2532,N_3092);
and U4259 (N_4259,N_3078,N_3047);
and U4260 (N_4260,N_3240,N_3321);
xor U4261 (N_4261,N_3705,N_3688);
xor U4262 (N_4262,N_3319,N_2886);
or U4263 (N_4263,N_3166,N_3159);
and U4264 (N_4264,N_2747,N_2897);
or U4265 (N_4265,N_3017,N_2504);
nor U4266 (N_4266,N_3239,N_2509);
and U4267 (N_4267,N_3026,N_2820);
nand U4268 (N_4268,N_3563,N_2596);
nor U4269 (N_4269,N_3744,N_3309);
and U4270 (N_4270,N_3274,N_3677);
xnor U4271 (N_4271,N_3654,N_3472);
nand U4272 (N_4272,N_3057,N_3327);
xnor U4273 (N_4273,N_3416,N_3202);
or U4274 (N_4274,N_2817,N_3174);
nand U4275 (N_4275,N_3231,N_3230);
or U4276 (N_4276,N_3666,N_3181);
xor U4277 (N_4277,N_3490,N_2783);
or U4278 (N_4278,N_2698,N_3606);
xnor U4279 (N_4279,N_3004,N_3497);
and U4280 (N_4280,N_2538,N_2648);
and U4281 (N_4281,N_3601,N_3571);
or U4282 (N_4282,N_2784,N_3587);
xnor U4283 (N_4283,N_2630,N_3091);
nand U4284 (N_4284,N_2939,N_3562);
nor U4285 (N_4285,N_3223,N_3306);
or U4286 (N_4286,N_2797,N_3595);
or U4287 (N_4287,N_3661,N_3002);
nand U4288 (N_4288,N_2833,N_3734);
nor U4289 (N_4289,N_2530,N_2516);
nor U4290 (N_4290,N_3343,N_2707);
or U4291 (N_4291,N_2903,N_3066);
nand U4292 (N_4292,N_2741,N_3000);
nand U4293 (N_4293,N_2536,N_3038);
and U4294 (N_4294,N_3207,N_3590);
and U4295 (N_4295,N_3636,N_2793);
and U4296 (N_4296,N_3543,N_2751);
nand U4297 (N_4297,N_2562,N_2557);
xor U4298 (N_4298,N_3584,N_2950);
nor U4299 (N_4299,N_3670,N_3398);
xor U4300 (N_4300,N_3072,N_2938);
nand U4301 (N_4301,N_3422,N_3725);
nor U4302 (N_4302,N_3352,N_2609);
and U4303 (N_4303,N_3005,N_2520);
nand U4304 (N_4304,N_3226,N_3698);
nand U4305 (N_4305,N_3341,N_2738);
or U4306 (N_4306,N_2565,N_2758);
or U4307 (N_4307,N_3694,N_2844);
xor U4308 (N_4308,N_3633,N_3710);
nor U4309 (N_4309,N_3475,N_3488);
xor U4310 (N_4310,N_3349,N_2710);
xor U4311 (N_4311,N_3294,N_2832);
and U4312 (N_4312,N_3575,N_3746);
nor U4313 (N_4313,N_3335,N_2744);
or U4314 (N_4314,N_3651,N_3245);
nand U4315 (N_4315,N_2667,N_3068);
nand U4316 (N_4316,N_3473,N_3500);
nand U4317 (N_4317,N_3067,N_3405);
or U4318 (N_4318,N_2875,N_2752);
and U4319 (N_4319,N_3353,N_3076);
xor U4320 (N_4320,N_3518,N_3234);
xor U4321 (N_4321,N_2625,N_2547);
and U4322 (N_4322,N_2700,N_2972);
nor U4323 (N_4323,N_3241,N_3394);
and U4324 (N_4324,N_3648,N_3260);
or U4325 (N_4325,N_3354,N_3205);
nand U4326 (N_4326,N_2916,N_3582);
and U4327 (N_4327,N_3020,N_2840);
nand U4328 (N_4328,N_3162,N_2589);
or U4329 (N_4329,N_2819,N_2998);
and U4330 (N_4330,N_3469,N_2597);
nand U4331 (N_4331,N_3738,N_3081);
and U4332 (N_4332,N_3709,N_3099);
xnor U4333 (N_4333,N_2619,N_3702);
nand U4334 (N_4334,N_3689,N_3503);
nor U4335 (N_4335,N_2810,N_2703);
and U4336 (N_4336,N_2501,N_2604);
xor U4337 (N_4337,N_2815,N_3550);
and U4338 (N_4338,N_2809,N_3219);
or U4339 (N_4339,N_2697,N_3371);
xor U4340 (N_4340,N_3284,N_3412);
and U4341 (N_4341,N_2992,N_2558);
or U4342 (N_4342,N_3432,N_3034);
xor U4343 (N_4343,N_2769,N_2718);
or U4344 (N_4344,N_3583,N_2812);
nor U4345 (N_4345,N_2525,N_3106);
nor U4346 (N_4346,N_3733,N_3225);
or U4347 (N_4347,N_2786,N_3069);
and U4348 (N_4348,N_3411,N_2983);
nor U4349 (N_4349,N_3261,N_3489);
nor U4350 (N_4350,N_3548,N_3292);
xnor U4351 (N_4351,N_3561,N_3178);
and U4352 (N_4352,N_2923,N_3183);
nor U4353 (N_4353,N_2611,N_2658);
and U4354 (N_4354,N_3275,N_3655);
and U4355 (N_4355,N_2640,N_3253);
xnor U4356 (N_4356,N_3520,N_2846);
xnor U4357 (N_4357,N_2656,N_3221);
nand U4358 (N_4358,N_2842,N_2715);
xnor U4359 (N_4359,N_3364,N_2879);
nand U4360 (N_4360,N_2940,N_2890);
nand U4361 (N_4361,N_3185,N_2754);
nor U4362 (N_4362,N_3296,N_3714);
nor U4363 (N_4363,N_3634,N_3508);
nor U4364 (N_4364,N_2724,N_2822);
xnor U4365 (N_4365,N_3288,N_3009);
and U4366 (N_4366,N_2576,N_3083);
xnor U4367 (N_4367,N_2912,N_2742);
nor U4368 (N_4368,N_2830,N_3058);
and U4369 (N_4369,N_2522,N_2637);
xor U4370 (N_4370,N_3721,N_3217);
nand U4371 (N_4371,N_3597,N_3218);
nand U4372 (N_4372,N_3616,N_2928);
xor U4373 (N_4373,N_2956,N_2514);
and U4374 (N_4374,N_2575,N_2735);
and U4375 (N_4375,N_3331,N_3424);
nand U4376 (N_4376,N_2780,N_3101);
and U4377 (N_4377,N_2829,N_2581);
and U4378 (N_4378,N_2898,N_2779);
nor U4379 (N_4379,N_3704,N_3293);
or U4380 (N_4380,N_2850,N_2710);
and U4381 (N_4381,N_3619,N_2726);
nand U4382 (N_4382,N_2810,N_3295);
nor U4383 (N_4383,N_3185,N_3418);
or U4384 (N_4384,N_3346,N_3186);
or U4385 (N_4385,N_2888,N_3490);
xnor U4386 (N_4386,N_3298,N_3740);
nor U4387 (N_4387,N_3018,N_2949);
nand U4388 (N_4388,N_3015,N_3113);
nand U4389 (N_4389,N_3209,N_2505);
nand U4390 (N_4390,N_3414,N_3167);
and U4391 (N_4391,N_2539,N_3095);
nor U4392 (N_4392,N_3731,N_3113);
nor U4393 (N_4393,N_2741,N_3215);
and U4394 (N_4394,N_3642,N_3667);
and U4395 (N_4395,N_3663,N_2532);
nand U4396 (N_4396,N_2910,N_2984);
nor U4397 (N_4397,N_2772,N_3093);
nand U4398 (N_4398,N_2651,N_3678);
nor U4399 (N_4399,N_3322,N_3587);
nand U4400 (N_4400,N_3269,N_2772);
and U4401 (N_4401,N_3743,N_2786);
nand U4402 (N_4402,N_2690,N_2877);
nand U4403 (N_4403,N_2767,N_3249);
nand U4404 (N_4404,N_2782,N_3499);
nor U4405 (N_4405,N_2790,N_3247);
nand U4406 (N_4406,N_2883,N_2991);
nor U4407 (N_4407,N_3515,N_3204);
or U4408 (N_4408,N_3512,N_3257);
xor U4409 (N_4409,N_2887,N_3679);
nand U4410 (N_4410,N_2907,N_2553);
and U4411 (N_4411,N_2650,N_3579);
nor U4412 (N_4412,N_3080,N_2648);
and U4413 (N_4413,N_2628,N_2964);
and U4414 (N_4414,N_2755,N_3042);
nand U4415 (N_4415,N_3082,N_3125);
nor U4416 (N_4416,N_3159,N_2634);
nor U4417 (N_4417,N_2750,N_2678);
xnor U4418 (N_4418,N_3718,N_2766);
nand U4419 (N_4419,N_2517,N_2999);
or U4420 (N_4420,N_3597,N_3095);
xor U4421 (N_4421,N_3094,N_2604);
nand U4422 (N_4422,N_3176,N_3215);
or U4423 (N_4423,N_3590,N_3130);
or U4424 (N_4424,N_2659,N_2932);
nor U4425 (N_4425,N_3365,N_3405);
nor U4426 (N_4426,N_3377,N_3411);
and U4427 (N_4427,N_2998,N_3525);
xor U4428 (N_4428,N_2504,N_2556);
nand U4429 (N_4429,N_3240,N_3281);
nand U4430 (N_4430,N_3376,N_3198);
nand U4431 (N_4431,N_2537,N_2630);
nand U4432 (N_4432,N_3643,N_3353);
nor U4433 (N_4433,N_2551,N_2894);
or U4434 (N_4434,N_2709,N_2752);
nor U4435 (N_4435,N_3734,N_3087);
nand U4436 (N_4436,N_2568,N_2878);
nand U4437 (N_4437,N_3185,N_2567);
xor U4438 (N_4438,N_2899,N_3506);
xor U4439 (N_4439,N_3115,N_3223);
and U4440 (N_4440,N_3337,N_2730);
nand U4441 (N_4441,N_2612,N_2642);
nand U4442 (N_4442,N_3484,N_3181);
nand U4443 (N_4443,N_3370,N_3162);
and U4444 (N_4444,N_3099,N_3104);
nand U4445 (N_4445,N_2535,N_3671);
nor U4446 (N_4446,N_2846,N_2789);
or U4447 (N_4447,N_3113,N_3301);
or U4448 (N_4448,N_3375,N_3626);
and U4449 (N_4449,N_3006,N_2631);
nand U4450 (N_4450,N_2638,N_3059);
and U4451 (N_4451,N_3300,N_2592);
nor U4452 (N_4452,N_3708,N_2721);
nand U4453 (N_4453,N_2607,N_3048);
or U4454 (N_4454,N_2661,N_2797);
nor U4455 (N_4455,N_2506,N_2509);
xor U4456 (N_4456,N_2688,N_3414);
or U4457 (N_4457,N_2982,N_3097);
or U4458 (N_4458,N_3241,N_3435);
xnor U4459 (N_4459,N_3080,N_2657);
and U4460 (N_4460,N_3425,N_3251);
and U4461 (N_4461,N_3190,N_3332);
xnor U4462 (N_4462,N_3347,N_3227);
and U4463 (N_4463,N_3337,N_3242);
xnor U4464 (N_4464,N_2755,N_2610);
and U4465 (N_4465,N_3324,N_3683);
xnor U4466 (N_4466,N_3527,N_2647);
xnor U4467 (N_4467,N_3390,N_2662);
nand U4468 (N_4468,N_2704,N_3308);
or U4469 (N_4469,N_3686,N_3106);
xnor U4470 (N_4470,N_3716,N_2815);
nor U4471 (N_4471,N_3269,N_3235);
and U4472 (N_4472,N_2990,N_2601);
or U4473 (N_4473,N_3246,N_3199);
nor U4474 (N_4474,N_2588,N_3494);
or U4475 (N_4475,N_3187,N_2779);
nand U4476 (N_4476,N_3069,N_2509);
or U4477 (N_4477,N_2836,N_3267);
nor U4478 (N_4478,N_3280,N_2606);
or U4479 (N_4479,N_2682,N_3224);
or U4480 (N_4480,N_3627,N_3340);
nand U4481 (N_4481,N_3220,N_3733);
nor U4482 (N_4482,N_3030,N_2612);
nand U4483 (N_4483,N_3160,N_3629);
nor U4484 (N_4484,N_3491,N_3559);
xor U4485 (N_4485,N_2960,N_2769);
xor U4486 (N_4486,N_2627,N_2802);
xnor U4487 (N_4487,N_3173,N_2726);
nand U4488 (N_4488,N_2536,N_3144);
xor U4489 (N_4489,N_3298,N_3184);
and U4490 (N_4490,N_3627,N_3112);
and U4491 (N_4491,N_2927,N_2806);
xnor U4492 (N_4492,N_2677,N_3393);
and U4493 (N_4493,N_2708,N_2914);
xor U4494 (N_4494,N_2955,N_3679);
xnor U4495 (N_4495,N_2724,N_3448);
xnor U4496 (N_4496,N_3491,N_3239);
xnor U4497 (N_4497,N_3142,N_2937);
xor U4498 (N_4498,N_3592,N_2512);
and U4499 (N_4499,N_3001,N_3312);
nand U4500 (N_4500,N_2821,N_3387);
and U4501 (N_4501,N_3419,N_3340);
nor U4502 (N_4502,N_2685,N_3542);
nor U4503 (N_4503,N_3529,N_2727);
and U4504 (N_4504,N_3618,N_3270);
or U4505 (N_4505,N_3399,N_2574);
and U4506 (N_4506,N_3663,N_3013);
or U4507 (N_4507,N_3389,N_3139);
xor U4508 (N_4508,N_3376,N_2853);
nand U4509 (N_4509,N_3003,N_3176);
xor U4510 (N_4510,N_2681,N_3223);
xor U4511 (N_4511,N_3006,N_3070);
xnor U4512 (N_4512,N_2819,N_2560);
and U4513 (N_4513,N_2848,N_3099);
nand U4514 (N_4514,N_2862,N_2706);
nand U4515 (N_4515,N_2705,N_3071);
nor U4516 (N_4516,N_2948,N_3663);
xnor U4517 (N_4517,N_3345,N_2734);
or U4518 (N_4518,N_3308,N_3144);
and U4519 (N_4519,N_3194,N_3119);
and U4520 (N_4520,N_2945,N_3678);
xnor U4521 (N_4521,N_3351,N_3164);
xnor U4522 (N_4522,N_2554,N_3137);
nand U4523 (N_4523,N_3257,N_3095);
nor U4524 (N_4524,N_2817,N_2867);
and U4525 (N_4525,N_3008,N_3174);
or U4526 (N_4526,N_3243,N_2847);
nor U4527 (N_4527,N_2800,N_2851);
xor U4528 (N_4528,N_3153,N_2933);
or U4529 (N_4529,N_3151,N_3449);
nor U4530 (N_4530,N_2797,N_2817);
nor U4531 (N_4531,N_2645,N_3489);
nand U4532 (N_4532,N_3085,N_2708);
nor U4533 (N_4533,N_3539,N_3291);
and U4534 (N_4534,N_3335,N_2737);
and U4535 (N_4535,N_3220,N_2660);
and U4536 (N_4536,N_2797,N_3244);
xnor U4537 (N_4537,N_3420,N_2762);
and U4538 (N_4538,N_2846,N_3557);
nor U4539 (N_4539,N_3022,N_3063);
xor U4540 (N_4540,N_2958,N_3320);
xor U4541 (N_4541,N_3198,N_2602);
nand U4542 (N_4542,N_2747,N_2877);
xor U4543 (N_4543,N_2865,N_3255);
xnor U4544 (N_4544,N_2619,N_2508);
or U4545 (N_4545,N_2899,N_3726);
or U4546 (N_4546,N_3243,N_2916);
nand U4547 (N_4547,N_2527,N_3304);
or U4548 (N_4548,N_3166,N_3685);
or U4549 (N_4549,N_3632,N_3009);
and U4550 (N_4550,N_3303,N_2512);
and U4551 (N_4551,N_3615,N_3624);
xnor U4552 (N_4552,N_2994,N_3298);
nor U4553 (N_4553,N_2904,N_2876);
and U4554 (N_4554,N_3110,N_3407);
xnor U4555 (N_4555,N_3341,N_2668);
xor U4556 (N_4556,N_2727,N_3457);
or U4557 (N_4557,N_2657,N_3164);
nand U4558 (N_4558,N_2607,N_3005);
or U4559 (N_4559,N_3180,N_3378);
nor U4560 (N_4560,N_2697,N_3294);
nand U4561 (N_4561,N_2846,N_2935);
nor U4562 (N_4562,N_2719,N_2988);
or U4563 (N_4563,N_3055,N_3000);
and U4564 (N_4564,N_2955,N_2534);
nor U4565 (N_4565,N_2743,N_2981);
or U4566 (N_4566,N_3380,N_3526);
or U4567 (N_4567,N_3537,N_3639);
xor U4568 (N_4568,N_3223,N_2678);
nand U4569 (N_4569,N_2712,N_3379);
or U4570 (N_4570,N_2898,N_3468);
nand U4571 (N_4571,N_2909,N_2878);
and U4572 (N_4572,N_2531,N_2606);
xnor U4573 (N_4573,N_3368,N_2837);
nor U4574 (N_4574,N_2799,N_3249);
nand U4575 (N_4575,N_3686,N_2590);
xor U4576 (N_4576,N_3460,N_3387);
nor U4577 (N_4577,N_2770,N_3257);
xor U4578 (N_4578,N_3341,N_3174);
nor U4579 (N_4579,N_2658,N_2866);
xnor U4580 (N_4580,N_3226,N_2890);
nor U4581 (N_4581,N_3439,N_3069);
nand U4582 (N_4582,N_3749,N_3098);
nor U4583 (N_4583,N_2528,N_3498);
nor U4584 (N_4584,N_3164,N_3204);
or U4585 (N_4585,N_2963,N_2601);
nor U4586 (N_4586,N_3554,N_3743);
nor U4587 (N_4587,N_3742,N_3044);
xor U4588 (N_4588,N_3319,N_3182);
xnor U4589 (N_4589,N_3480,N_3020);
nand U4590 (N_4590,N_3633,N_3602);
and U4591 (N_4591,N_3411,N_3160);
nor U4592 (N_4592,N_3059,N_3207);
nor U4593 (N_4593,N_2502,N_3306);
xor U4594 (N_4594,N_2658,N_3368);
xor U4595 (N_4595,N_3709,N_3295);
nor U4596 (N_4596,N_2731,N_2564);
and U4597 (N_4597,N_3602,N_2554);
nor U4598 (N_4598,N_2562,N_3658);
and U4599 (N_4599,N_3436,N_3104);
and U4600 (N_4600,N_2606,N_2724);
nand U4601 (N_4601,N_3470,N_2654);
xor U4602 (N_4602,N_3076,N_3702);
or U4603 (N_4603,N_2740,N_2575);
nand U4604 (N_4604,N_2690,N_3499);
or U4605 (N_4605,N_3312,N_2581);
xnor U4606 (N_4606,N_2950,N_2798);
nand U4607 (N_4607,N_3316,N_2845);
and U4608 (N_4608,N_2974,N_2907);
xnor U4609 (N_4609,N_3016,N_3209);
xor U4610 (N_4610,N_3425,N_2832);
and U4611 (N_4611,N_2882,N_3487);
nand U4612 (N_4612,N_2888,N_3088);
xnor U4613 (N_4613,N_3501,N_2528);
nand U4614 (N_4614,N_3733,N_3455);
or U4615 (N_4615,N_3687,N_2753);
xor U4616 (N_4616,N_3365,N_2929);
nor U4617 (N_4617,N_2598,N_2669);
xor U4618 (N_4618,N_2684,N_2798);
nor U4619 (N_4619,N_3008,N_3106);
nand U4620 (N_4620,N_2954,N_3325);
and U4621 (N_4621,N_3228,N_3378);
nand U4622 (N_4622,N_3124,N_3278);
or U4623 (N_4623,N_3685,N_2538);
or U4624 (N_4624,N_3431,N_3103);
nand U4625 (N_4625,N_2752,N_2926);
and U4626 (N_4626,N_3344,N_3609);
xor U4627 (N_4627,N_3542,N_3130);
xnor U4628 (N_4628,N_2612,N_3326);
nand U4629 (N_4629,N_2713,N_2894);
nand U4630 (N_4630,N_3293,N_3278);
or U4631 (N_4631,N_3402,N_3266);
or U4632 (N_4632,N_3352,N_3139);
nor U4633 (N_4633,N_2830,N_2703);
or U4634 (N_4634,N_3032,N_2866);
nor U4635 (N_4635,N_3279,N_3272);
or U4636 (N_4636,N_3266,N_2729);
nor U4637 (N_4637,N_3032,N_3180);
or U4638 (N_4638,N_2875,N_3152);
nor U4639 (N_4639,N_3545,N_2951);
and U4640 (N_4640,N_3139,N_2553);
xor U4641 (N_4641,N_3014,N_3379);
nand U4642 (N_4642,N_3049,N_3621);
nor U4643 (N_4643,N_3640,N_3490);
and U4644 (N_4644,N_2777,N_2853);
xnor U4645 (N_4645,N_3461,N_3578);
nand U4646 (N_4646,N_2987,N_3394);
nand U4647 (N_4647,N_2649,N_3495);
nor U4648 (N_4648,N_2887,N_3422);
nor U4649 (N_4649,N_2517,N_3732);
nor U4650 (N_4650,N_2632,N_3287);
xor U4651 (N_4651,N_2925,N_3115);
or U4652 (N_4652,N_3314,N_2917);
nor U4653 (N_4653,N_3432,N_3361);
nand U4654 (N_4654,N_3288,N_3229);
or U4655 (N_4655,N_3479,N_2910);
or U4656 (N_4656,N_3056,N_3664);
nor U4657 (N_4657,N_3600,N_3282);
nand U4658 (N_4658,N_3095,N_2545);
and U4659 (N_4659,N_2723,N_2656);
nand U4660 (N_4660,N_3005,N_3578);
and U4661 (N_4661,N_3056,N_3321);
nor U4662 (N_4662,N_3654,N_3389);
nor U4663 (N_4663,N_2768,N_3004);
and U4664 (N_4664,N_2573,N_2683);
nor U4665 (N_4665,N_3547,N_3646);
nand U4666 (N_4666,N_3577,N_2984);
or U4667 (N_4667,N_3349,N_3566);
nand U4668 (N_4668,N_3189,N_2824);
nor U4669 (N_4669,N_3388,N_3517);
or U4670 (N_4670,N_3656,N_2585);
nand U4671 (N_4671,N_3465,N_3138);
xnor U4672 (N_4672,N_3637,N_2996);
or U4673 (N_4673,N_3229,N_2767);
xor U4674 (N_4674,N_3413,N_2800);
xnor U4675 (N_4675,N_2505,N_3546);
xor U4676 (N_4676,N_2825,N_2563);
or U4677 (N_4677,N_3590,N_2975);
xnor U4678 (N_4678,N_2937,N_2743);
or U4679 (N_4679,N_3475,N_3111);
nand U4680 (N_4680,N_3184,N_3351);
xor U4681 (N_4681,N_3575,N_2749);
and U4682 (N_4682,N_3640,N_3511);
or U4683 (N_4683,N_3064,N_3089);
nor U4684 (N_4684,N_3682,N_2926);
or U4685 (N_4685,N_3412,N_3057);
and U4686 (N_4686,N_2502,N_3470);
or U4687 (N_4687,N_3297,N_3364);
xnor U4688 (N_4688,N_3646,N_3478);
xnor U4689 (N_4689,N_3000,N_2856);
nor U4690 (N_4690,N_2859,N_2657);
nand U4691 (N_4691,N_2911,N_3673);
nor U4692 (N_4692,N_2608,N_3455);
xor U4693 (N_4693,N_2821,N_3413);
nand U4694 (N_4694,N_3677,N_2951);
xor U4695 (N_4695,N_2959,N_2756);
nor U4696 (N_4696,N_2746,N_2525);
nor U4697 (N_4697,N_3678,N_3232);
nor U4698 (N_4698,N_3248,N_3014);
and U4699 (N_4699,N_3748,N_3273);
nor U4700 (N_4700,N_3410,N_3711);
or U4701 (N_4701,N_3386,N_2930);
or U4702 (N_4702,N_2600,N_3032);
or U4703 (N_4703,N_2948,N_3341);
nand U4704 (N_4704,N_3658,N_2662);
nand U4705 (N_4705,N_2725,N_2553);
xnor U4706 (N_4706,N_3495,N_3313);
and U4707 (N_4707,N_3217,N_2508);
and U4708 (N_4708,N_3346,N_2925);
nor U4709 (N_4709,N_3631,N_2971);
xor U4710 (N_4710,N_3390,N_3468);
nor U4711 (N_4711,N_2524,N_3009);
xor U4712 (N_4712,N_3244,N_3343);
and U4713 (N_4713,N_2659,N_2665);
or U4714 (N_4714,N_3126,N_3278);
and U4715 (N_4715,N_2851,N_2969);
nand U4716 (N_4716,N_3267,N_2694);
xnor U4717 (N_4717,N_2551,N_3524);
and U4718 (N_4718,N_3259,N_3334);
nand U4719 (N_4719,N_3329,N_3415);
or U4720 (N_4720,N_2515,N_3050);
xnor U4721 (N_4721,N_2815,N_3698);
nand U4722 (N_4722,N_3320,N_3695);
xor U4723 (N_4723,N_3298,N_3314);
nand U4724 (N_4724,N_3503,N_3349);
xnor U4725 (N_4725,N_2506,N_3562);
xnor U4726 (N_4726,N_3367,N_3417);
xor U4727 (N_4727,N_2584,N_3461);
and U4728 (N_4728,N_2749,N_3564);
nor U4729 (N_4729,N_2792,N_3269);
nor U4730 (N_4730,N_2673,N_3224);
nor U4731 (N_4731,N_2706,N_2913);
nand U4732 (N_4732,N_3173,N_3519);
nor U4733 (N_4733,N_2729,N_3218);
xnor U4734 (N_4734,N_2780,N_3262);
or U4735 (N_4735,N_2771,N_2615);
and U4736 (N_4736,N_3187,N_3524);
nor U4737 (N_4737,N_2618,N_3414);
and U4738 (N_4738,N_3086,N_3297);
nor U4739 (N_4739,N_3389,N_3719);
nor U4740 (N_4740,N_2933,N_3102);
and U4741 (N_4741,N_3302,N_3246);
nand U4742 (N_4742,N_2907,N_3114);
and U4743 (N_4743,N_3181,N_3365);
nor U4744 (N_4744,N_3655,N_2680);
xor U4745 (N_4745,N_3459,N_2945);
nand U4746 (N_4746,N_2992,N_3307);
nand U4747 (N_4747,N_2547,N_3214);
xor U4748 (N_4748,N_3555,N_3247);
and U4749 (N_4749,N_3319,N_3026);
and U4750 (N_4750,N_2771,N_3072);
nor U4751 (N_4751,N_2957,N_3649);
xnor U4752 (N_4752,N_2625,N_3294);
nand U4753 (N_4753,N_3666,N_3564);
nor U4754 (N_4754,N_2830,N_2739);
nand U4755 (N_4755,N_3728,N_3570);
nand U4756 (N_4756,N_3253,N_2622);
and U4757 (N_4757,N_3726,N_2728);
nand U4758 (N_4758,N_3192,N_3046);
and U4759 (N_4759,N_3157,N_3094);
xor U4760 (N_4760,N_3070,N_2917);
and U4761 (N_4761,N_2735,N_3529);
or U4762 (N_4762,N_3515,N_2769);
nor U4763 (N_4763,N_2785,N_2724);
and U4764 (N_4764,N_3109,N_2781);
xnor U4765 (N_4765,N_2506,N_2649);
xor U4766 (N_4766,N_2981,N_3639);
xnor U4767 (N_4767,N_2554,N_2639);
nand U4768 (N_4768,N_2788,N_2898);
and U4769 (N_4769,N_2994,N_3655);
nor U4770 (N_4770,N_2836,N_3070);
xor U4771 (N_4771,N_3002,N_3626);
or U4772 (N_4772,N_3478,N_2696);
and U4773 (N_4773,N_3239,N_3001);
xor U4774 (N_4774,N_2918,N_2611);
nor U4775 (N_4775,N_2971,N_3451);
nand U4776 (N_4776,N_2992,N_3259);
nor U4777 (N_4777,N_2504,N_3575);
xor U4778 (N_4778,N_3452,N_2543);
xor U4779 (N_4779,N_2513,N_3415);
and U4780 (N_4780,N_2653,N_2779);
nand U4781 (N_4781,N_3362,N_3032);
or U4782 (N_4782,N_3009,N_2825);
nor U4783 (N_4783,N_3740,N_2528);
or U4784 (N_4784,N_3335,N_3455);
nand U4785 (N_4785,N_2798,N_2886);
nor U4786 (N_4786,N_3184,N_2844);
xnor U4787 (N_4787,N_3215,N_2816);
and U4788 (N_4788,N_3236,N_3416);
and U4789 (N_4789,N_3085,N_3455);
or U4790 (N_4790,N_2924,N_3048);
and U4791 (N_4791,N_3190,N_3192);
nand U4792 (N_4792,N_3276,N_3677);
xnor U4793 (N_4793,N_2927,N_2956);
or U4794 (N_4794,N_3476,N_2774);
nor U4795 (N_4795,N_2717,N_3663);
or U4796 (N_4796,N_2731,N_2767);
xor U4797 (N_4797,N_3485,N_2823);
xor U4798 (N_4798,N_2928,N_3346);
nor U4799 (N_4799,N_3660,N_3670);
or U4800 (N_4800,N_3084,N_2723);
or U4801 (N_4801,N_2679,N_3459);
or U4802 (N_4802,N_3459,N_3170);
nor U4803 (N_4803,N_3051,N_3059);
xor U4804 (N_4804,N_3748,N_3656);
xor U4805 (N_4805,N_3149,N_2647);
nand U4806 (N_4806,N_3143,N_3029);
and U4807 (N_4807,N_2981,N_3235);
nor U4808 (N_4808,N_2767,N_3508);
nor U4809 (N_4809,N_3085,N_2761);
and U4810 (N_4810,N_2636,N_2967);
or U4811 (N_4811,N_3328,N_3069);
and U4812 (N_4812,N_2705,N_3504);
nand U4813 (N_4813,N_2904,N_3618);
xnor U4814 (N_4814,N_2671,N_3367);
xnor U4815 (N_4815,N_2588,N_3733);
and U4816 (N_4816,N_2946,N_3022);
nand U4817 (N_4817,N_2754,N_3433);
or U4818 (N_4818,N_3731,N_2999);
nand U4819 (N_4819,N_2764,N_3636);
xor U4820 (N_4820,N_3288,N_3467);
nor U4821 (N_4821,N_3165,N_3589);
nand U4822 (N_4822,N_2747,N_3007);
and U4823 (N_4823,N_2795,N_2966);
xnor U4824 (N_4824,N_3159,N_3617);
nor U4825 (N_4825,N_2506,N_2666);
nand U4826 (N_4826,N_3646,N_2805);
nand U4827 (N_4827,N_3213,N_3673);
nor U4828 (N_4828,N_2693,N_2960);
nand U4829 (N_4829,N_3538,N_3208);
nor U4830 (N_4830,N_3661,N_3546);
xor U4831 (N_4831,N_2961,N_3388);
and U4832 (N_4832,N_3185,N_3387);
nor U4833 (N_4833,N_3671,N_3586);
nor U4834 (N_4834,N_2739,N_3305);
nor U4835 (N_4835,N_3559,N_3537);
nor U4836 (N_4836,N_2991,N_2776);
nor U4837 (N_4837,N_2525,N_2998);
and U4838 (N_4838,N_3700,N_2616);
nand U4839 (N_4839,N_3274,N_2893);
or U4840 (N_4840,N_3199,N_3745);
nor U4841 (N_4841,N_2695,N_2526);
or U4842 (N_4842,N_2780,N_2760);
or U4843 (N_4843,N_3469,N_3298);
nand U4844 (N_4844,N_3001,N_3696);
nor U4845 (N_4845,N_3647,N_3383);
and U4846 (N_4846,N_3111,N_3305);
xor U4847 (N_4847,N_3412,N_2657);
and U4848 (N_4848,N_3350,N_3417);
and U4849 (N_4849,N_3478,N_3159);
or U4850 (N_4850,N_2653,N_2849);
nand U4851 (N_4851,N_3545,N_2678);
and U4852 (N_4852,N_2671,N_3626);
or U4853 (N_4853,N_3066,N_2852);
nand U4854 (N_4854,N_3147,N_2587);
nand U4855 (N_4855,N_3371,N_3667);
nand U4856 (N_4856,N_3214,N_3281);
xnor U4857 (N_4857,N_2727,N_2948);
and U4858 (N_4858,N_2986,N_3498);
xnor U4859 (N_4859,N_2747,N_2604);
nor U4860 (N_4860,N_3013,N_2780);
nor U4861 (N_4861,N_3658,N_2625);
and U4862 (N_4862,N_2588,N_3626);
nand U4863 (N_4863,N_2556,N_3235);
and U4864 (N_4864,N_2654,N_3598);
nor U4865 (N_4865,N_2834,N_3110);
and U4866 (N_4866,N_2836,N_3265);
or U4867 (N_4867,N_3268,N_2886);
nand U4868 (N_4868,N_3609,N_2786);
or U4869 (N_4869,N_3537,N_3027);
xor U4870 (N_4870,N_3744,N_2761);
xor U4871 (N_4871,N_2558,N_3148);
xnor U4872 (N_4872,N_3152,N_2534);
nor U4873 (N_4873,N_3213,N_2650);
and U4874 (N_4874,N_3048,N_3548);
nand U4875 (N_4875,N_3586,N_3415);
or U4876 (N_4876,N_2941,N_3414);
xnor U4877 (N_4877,N_2774,N_2521);
and U4878 (N_4878,N_3380,N_2764);
and U4879 (N_4879,N_3180,N_2809);
xnor U4880 (N_4880,N_3436,N_2896);
and U4881 (N_4881,N_3040,N_2952);
or U4882 (N_4882,N_3525,N_3251);
and U4883 (N_4883,N_3205,N_2914);
and U4884 (N_4884,N_3313,N_2860);
or U4885 (N_4885,N_3618,N_2918);
and U4886 (N_4886,N_2709,N_3641);
xor U4887 (N_4887,N_3320,N_2598);
and U4888 (N_4888,N_2824,N_2722);
nor U4889 (N_4889,N_3086,N_3409);
nor U4890 (N_4890,N_2763,N_2866);
nor U4891 (N_4891,N_3017,N_2507);
nand U4892 (N_4892,N_3720,N_2898);
xnor U4893 (N_4893,N_3059,N_3274);
and U4894 (N_4894,N_2993,N_3533);
nand U4895 (N_4895,N_3262,N_2549);
nor U4896 (N_4896,N_2896,N_3373);
xnor U4897 (N_4897,N_2780,N_3230);
nor U4898 (N_4898,N_2627,N_2928);
nor U4899 (N_4899,N_2963,N_3378);
xor U4900 (N_4900,N_3666,N_3405);
nand U4901 (N_4901,N_3601,N_2756);
xor U4902 (N_4902,N_3126,N_3228);
and U4903 (N_4903,N_3032,N_3375);
nand U4904 (N_4904,N_2986,N_2756);
nand U4905 (N_4905,N_3071,N_2878);
nor U4906 (N_4906,N_2838,N_3035);
nand U4907 (N_4907,N_2700,N_3373);
nand U4908 (N_4908,N_2797,N_3462);
or U4909 (N_4909,N_3572,N_2502);
and U4910 (N_4910,N_2770,N_2535);
or U4911 (N_4911,N_2640,N_3675);
or U4912 (N_4912,N_3304,N_3133);
or U4913 (N_4913,N_2576,N_3488);
and U4914 (N_4914,N_3588,N_2882);
xor U4915 (N_4915,N_2550,N_3724);
nor U4916 (N_4916,N_2667,N_3371);
nand U4917 (N_4917,N_3272,N_2877);
nor U4918 (N_4918,N_3004,N_2928);
xor U4919 (N_4919,N_3521,N_3491);
nand U4920 (N_4920,N_3257,N_2673);
nor U4921 (N_4921,N_3483,N_3132);
xnor U4922 (N_4922,N_2910,N_2500);
nand U4923 (N_4923,N_3569,N_3444);
nand U4924 (N_4924,N_2825,N_3280);
nand U4925 (N_4925,N_3433,N_3361);
xnor U4926 (N_4926,N_3368,N_3508);
nand U4927 (N_4927,N_2772,N_3336);
and U4928 (N_4928,N_2578,N_3351);
nor U4929 (N_4929,N_3162,N_3688);
xor U4930 (N_4930,N_3359,N_2577);
and U4931 (N_4931,N_2960,N_2614);
nor U4932 (N_4932,N_3081,N_2620);
xor U4933 (N_4933,N_3468,N_3244);
or U4934 (N_4934,N_3065,N_2693);
xnor U4935 (N_4935,N_2982,N_2845);
nand U4936 (N_4936,N_3535,N_3739);
or U4937 (N_4937,N_2616,N_3121);
nor U4938 (N_4938,N_2759,N_3491);
xor U4939 (N_4939,N_3126,N_3554);
nand U4940 (N_4940,N_2860,N_2561);
nor U4941 (N_4941,N_3194,N_2910);
or U4942 (N_4942,N_3715,N_3456);
nor U4943 (N_4943,N_3591,N_3560);
nand U4944 (N_4944,N_3337,N_3309);
or U4945 (N_4945,N_2580,N_2784);
nor U4946 (N_4946,N_2565,N_2918);
or U4947 (N_4947,N_3654,N_3201);
xnor U4948 (N_4948,N_3627,N_3306);
nor U4949 (N_4949,N_3130,N_3459);
xor U4950 (N_4950,N_2947,N_2506);
xor U4951 (N_4951,N_2578,N_2936);
and U4952 (N_4952,N_2913,N_3605);
and U4953 (N_4953,N_3339,N_2808);
and U4954 (N_4954,N_2674,N_3127);
nor U4955 (N_4955,N_2913,N_2815);
or U4956 (N_4956,N_3741,N_2685);
nand U4957 (N_4957,N_2538,N_2836);
nand U4958 (N_4958,N_3013,N_3011);
nand U4959 (N_4959,N_3659,N_2573);
and U4960 (N_4960,N_3325,N_3356);
and U4961 (N_4961,N_3472,N_2928);
nand U4962 (N_4962,N_3426,N_3730);
nor U4963 (N_4963,N_3063,N_2603);
or U4964 (N_4964,N_2830,N_3653);
xnor U4965 (N_4965,N_3514,N_3035);
xor U4966 (N_4966,N_3563,N_3464);
xnor U4967 (N_4967,N_3467,N_3454);
nor U4968 (N_4968,N_3062,N_3184);
nand U4969 (N_4969,N_2503,N_2975);
nor U4970 (N_4970,N_2868,N_2880);
nor U4971 (N_4971,N_3643,N_3015);
or U4972 (N_4972,N_3504,N_3229);
xnor U4973 (N_4973,N_3452,N_3713);
or U4974 (N_4974,N_2642,N_2768);
nor U4975 (N_4975,N_2600,N_3737);
nand U4976 (N_4976,N_2984,N_3506);
nand U4977 (N_4977,N_3290,N_2544);
or U4978 (N_4978,N_3259,N_3038);
nor U4979 (N_4979,N_3706,N_2885);
or U4980 (N_4980,N_3414,N_3679);
nor U4981 (N_4981,N_2987,N_3469);
and U4982 (N_4982,N_3551,N_3641);
and U4983 (N_4983,N_3551,N_3254);
nand U4984 (N_4984,N_3004,N_3396);
and U4985 (N_4985,N_2633,N_3065);
nor U4986 (N_4986,N_3168,N_3263);
xor U4987 (N_4987,N_2641,N_3563);
nand U4988 (N_4988,N_3156,N_3093);
nand U4989 (N_4989,N_3442,N_3289);
xor U4990 (N_4990,N_2843,N_3413);
xnor U4991 (N_4991,N_2760,N_2814);
nor U4992 (N_4992,N_2649,N_3742);
nand U4993 (N_4993,N_2838,N_2732);
nor U4994 (N_4994,N_3476,N_3314);
nor U4995 (N_4995,N_3518,N_2902);
or U4996 (N_4996,N_2777,N_2616);
xnor U4997 (N_4997,N_3315,N_2762);
nand U4998 (N_4998,N_3725,N_2826);
nand U4999 (N_4999,N_3485,N_3605);
or U5000 (N_5000,N_4700,N_3883);
xor U5001 (N_5001,N_4723,N_3768);
nor U5002 (N_5002,N_4861,N_4641);
and U5003 (N_5003,N_4749,N_4181);
nand U5004 (N_5004,N_4519,N_4414);
and U5005 (N_5005,N_4758,N_4193);
xnor U5006 (N_5006,N_3953,N_4960);
xor U5007 (N_5007,N_4243,N_4177);
or U5008 (N_5008,N_3755,N_4237);
xor U5009 (N_5009,N_4020,N_4744);
xnor U5010 (N_5010,N_4547,N_3978);
nor U5011 (N_5011,N_4435,N_4546);
nand U5012 (N_5012,N_4727,N_4620);
nand U5013 (N_5013,N_4596,N_4075);
and U5014 (N_5014,N_3945,N_3837);
and U5015 (N_5015,N_4799,N_3913);
nor U5016 (N_5016,N_4334,N_3879);
or U5017 (N_5017,N_4287,N_4567);
xor U5018 (N_5018,N_4092,N_3830);
or U5019 (N_5019,N_4695,N_3952);
nor U5020 (N_5020,N_3779,N_4467);
or U5021 (N_5021,N_4760,N_4374);
xor U5022 (N_5022,N_4431,N_4013);
and U5023 (N_5023,N_4011,N_4420);
or U5024 (N_5024,N_4750,N_4557);
xor U5025 (N_5025,N_4226,N_4327);
nand U5026 (N_5026,N_4080,N_4787);
nor U5027 (N_5027,N_3948,N_4742);
or U5028 (N_5028,N_4354,N_4136);
nor U5029 (N_5029,N_4003,N_4301);
nor U5030 (N_5030,N_3990,N_4077);
nand U5031 (N_5031,N_3886,N_4631);
nand U5032 (N_5032,N_4615,N_3991);
nor U5033 (N_5033,N_4937,N_4846);
or U5034 (N_5034,N_3910,N_4297);
xnor U5035 (N_5035,N_3798,N_4642);
and U5036 (N_5036,N_4432,N_4169);
and U5037 (N_5037,N_3759,N_4324);
and U5038 (N_5038,N_4681,N_4212);
and U5039 (N_5039,N_4685,N_4307);
and U5040 (N_5040,N_3822,N_4259);
and U5041 (N_5041,N_4189,N_4558);
xor U5042 (N_5042,N_4261,N_4663);
or U5043 (N_5043,N_3806,N_3944);
nor U5044 (N_5044,N_4292,N_4168);
nand U5045 (N_5045,N_4510,N_4361);
nand U5046 (N_5046,N_4221,N_4609);
xnor U5047 (N_5047,N_3930,N_3896);
xor U5048 (N_5048,N_4209,N_4483);
nand U5049 (N_5049,N_4920,N_3771);
or U5050 (N_5050,N_4199,N_4712);
xnor U5051 (N_5051,N_4233,N_4054);
xnor U5052 (N_5052,N_3914,N_3794);
and U5053 (N_5053,N_3773,N_4205);
xor U5054 (N_5054,N_4676,N_4931);
and U5055 (N_5055,N_4048,N_4577);
xor U5056 (N_5056,N_3926,N_4569);
nor U5057 (N_5057,N_4529,N_3942);
nor U5058 (N_5058,N_4608,N_4800);
and U5059 (N_5059,N_4564,N_4217);
xor U5060 (N_5060,N_4159,N_4272);
or U5061 (N_5061,N_3958,N_3792);
or U5062 (N_5062,N_3843,N_4900);
or U5063 (N_5063,N_4797,N_3826);
nand U5064 (N_5064,N_4521,N_4341);
nor U5065 (N_5065,N_3996,N_3937);
xor U5066 (N_5066,N_4008,N_4699);
and U5067 (N_5067,N_4893,N_4556);
nor U5068 (N_5068,N_4190,N_4965);
or U5069 (N_5069,N_4638,N_3970);
or U5070 (N_5070,N_4228,N_3935);
xor U5071 (N_5071,N_4767,N_4581);
nand U5072 (N_5072,N_4376,N_4686);
or U5073 (N_5073,N_4188,N_4145);
nor U5074 (N_5074,N_4491,N_4304);
xnor U5075 (N_5075,N_4339,N_3919);
and U5076 (N_5076,N_4829,N_4026);
and U5077 (N_5077,N_3957,N_4945);
or U5078 (N_5078,N_4299,N_4260);
nor U5079 (N_5079,N_4633,N_4213);
nand U5080 (N_5080,N_4129,N_4202);
nor U5081 (N_5081,N_4206,N_4288);
or U5082 (N_5082,N_4315,N_4618);
nand U5083 (N_5083,N_4834,N_4972);
nand U5084 (N_5084,N_4612,N_3797);
xnor U5085 (N_5085,N_4268,N_4939);
and U5086 (N_5086,N_4605,N_4105);
or U5087 (N_5087,N_3834,N_4671);
nand U5088 (N_5088,N_4009,N_4369);
nand U5089 (N_5089,N_4865,N_4667);
or U5090 (N_5090,N_4669,N_4479);
nor U5091 (N_5091,N_4300,N_4805);
and U5092 (N_5092,N_4746,N_4338);
and U5093 (N_5093,N_3868,N_3972);
nand U5094 (N_5094,N_4757,N_4047);
nor U5095 (N_5095,N_4678,N_3908);
nor U5096 (N_5096,N_4540,N_3998);
and U5097 (N_5097,N_4333,N_4824);
nor U5098 (N_5098,N_4842,N_3936);
xor U5099 (N_5099,N_4654,N_4860);
or U5100 (N_5100,N_4687,N_4684);
nand U5101 (N_5101,N_4910,N_4122);
or U5102 (N_5102,N_4215,N_4500);
nand U5103 (N_5103,N_4401,N_4889);
or U5104 (N_5104,N_3753,N_4879);
or U5105 (N_5105,N_4533,N_3808);
and U5106 (N_5106,N_4400,N_3802);
nand U5107 (N_5107,N_4033,N_4396);
nor U5108 (N_5108,N_4938,N_3891);
xnor U5109 (N_5109,N_4405,N_3774);
xor U5110 (N_5110,N_3988,N_3848);
nor U5111 (N_5111,N_4138,N_4722);
xor U5112 (N_5112,N_3880,N_4843);
and U5113 (N_5113,N_4406,N_4086);
nand U5114 (N_5114,N_4597,N_4155);
and U5115 (N_5115,N_4162,N_4492);
and U5116 (N_5116,N_4908,N_4358);
nor U5117 (N_5117,N_4314,N_3928);
and U5118 (N_5118,N_4065,N_4290);
nor U5119 (N_5119,N_4647,N_4562);
xnor U5120 (N_5120,N_4344,N_4457);
nand U5121 (N_5121,N_4715,N_3845);
xnor U5122 (N_5122,N_4921,N_4897);
nor U5123 (N_5123,N_4848,N_4850);
xnor U5124 (N_5124,N_4885,N_4192);
or U5125 (N_5125,N_4902,N_4508);
nand U5126 (N_5126,N_4929,N_3812);
and U5127 (N_5127,N_4303,N_4040);
or U5128 (N_5128,N_4954,N_4121);
or U5129 (N_5129,N_4518,N_3777);
and U5130 (N_5130,N_4216,N_4724);
nor U5131 (N_5131,N_4704,N_4777);
nor U5132 (N_5132,N_4208,N_4273);
xor U5133 (N_5133,N_4796,N_4068);
xor U5134 (N_5134,N_4941,N_4490);
nand U5135 (N_5135,N_4839,N_3923);
and U5136 (N_5136,N_4689,N_4183);
nand U5137 (N_5137,N_4201,N_4336);
or U5138 (N_5138,N_3756,N_4340);
and U5139 (N_5139,N_4610,N_3855);
or U5140 (N_5140,N_4607,N_3764);
nor U5141 (N_5141,N_3849,N_3751);
xor U5142 (N_5142,N_4565,N_4911);
xnor U5143 (N_5143,N_4450,N_3831);
nor U5144 (N_5144,N_4958,N_4982);
and U5145 (N_5145,N_3854,N_4692);
or U5146 (N_5146,N_4643,N_4347);
xor U5147 (N_5147,N_3968,N_4106);
or U5148 (N_5148,N_4688,N_4814);
nand U5149 (N_5149,N_4262,N_4674);
or U5150 (N_5150,N_3761,N_4868);
nand U5151 (N_5151,N_4094,N_4955);
xor U5152 (N_5152,N_3782,N_4079);
nand U5153 (N_5153,N_4587,N_4985);
nand U5154 (N_5154,N_3770,N_4321);
nand U5155 (N_5155,N_4127,N_3765);
and U5156 (N_5156,N_4161,N_4318);
and U5157 (N_5157,N_4291,N_4390);
and U5158 (N_5158,N_3795,N_4769);
or U5159 (N_5159,N_4974,N_3922);
or U5160 (N_5160,N_4646,N_4294);
and U5161 (N_5161,N_4725,N_4058);
nand U5162 (N_5162,N_4442,N_4527);
xnor U5163 (N_5163,N_4528,N_4320);
nand U5164 (N_5164,N_4433,N_3840);
or U5165 (N_5165,N_4143,N_4934);
nand U5166 (N_5166,N_4069,N_4813);
xor U5167 (N_5167,N_4660,N_4255);
or U5168 (N_5168,N_4496,N_4426);
or U5169 (N_5169,N_4025,N_4776);
or U5170 (N_5170,N_4514,N_3882);
nand U5171 (N_5171,N_4087,N_4096);
xnor U5172 (N_5172,N_4883,N_4266);
nor U5173 (N_5173,N_4439,N_4530);
and U5174 (N_5174,N_3790,N_3967);
nand U5175 (N_5175,N_4389,N_4708);
or U5176 (N_5176,N_4295,N_3989);
or U5177 (N_5177,N_4658,N_4670);
and U5178 (N_5178,N_4099,N_3841);
xor U5179 (N_5179,N_4651,N_4962);
and U5180 (N_5180,N_4055,N_4343);
and U5181 (N_5181,N_4480,N_3864);
nand U5182 (N_5182,N_4017,N_4733);
or U5183 (N_5183,N_4798,N_4554);
and U5184 (N_5184,N_4119,N_4981);
and U5185 (N_5185,N_4544,N_3899);
nand U5186 (N_5186,N_3807,N_4589);
and U5187 (N_5187,N_4229,N_4485);
xor U5188 (N_5188,N_4180,N_4182);
xor U5189 (N_5189,N_4640,N_4034);
nor U5190 (N_5190,N_4996,N_4498);
nor U5191 (N_5191,N_4046,N_4588);
or U5192 (N_5192,N_4909,N_3805);
and U5193 (N_5193,N_4768,N_4653);
and U5194 (N_5194,N_4319,N_4146);
nand U5195 (N_5195,N_4648,N_4482);
or U5196 (N_5196,N_4989,N_4819);
nand U5197 (N_5197,N_4041,N_4966);
xnor U5198 (N_5198,N_4027,N_4207);
and U5199 (N_5199,N_4575,N_4821);
xor U5200 (N_5200,N_4466,N_4306);
and U5201 (N_5201,N_4582,N_4252);
or U5202 (N_5202,N_3932,N_4736);
nor U5203 (N_5203,N_4896,N_4455);
xnor U5204 (N_5204,N_3762,N_4279);
and U5205 (N_5205,N_4083,N_4269);
nor U5206 (N_5206,N_4994,N_4050);
xnor U5207 (N_5207,N_3889,N_4826);
xor U5208 (N_5208,N_4352,N_3860);
xnor U5209 (N_5209,N_4384,N_4445);
nor U5210 (N_5210,N_4021,N_4731);
xnor U5211 (N_5211,N_4130,N_4331);
and U5212 (N_5212,N_4603,N_3897);
nor U5213 (N_5213,N_4032,N_3785);
xor U5214 (N_5214,N_4368,N_4976);
xor U5215 (N_5215,N_4894,N_4745);
and U5216 (N_5216,N_4249,N_4171);
and U5217 (N_5217,N_3817,N_4986);
xnor U5218 (N_5218,N_4015,N_4906);
nor U5219 (N_5219,N_4553,N_4147);
nor U5220 (N_5220,N_4815,N_4197);
nor U5221 (N_5221,N_3877,N_4363);
and U5222 (N_5222,N_4971,N_4253);
and U5223 (N_5223,N_4875,N_4112);
and U5224 (N_5224,N_4353,N_4617);
xor U5225 (N_5225,N_4023,N_4264);
xor U5226 (N_5226,N_3796,N_4936);
nand U5227 (N_5227,N_4018,N_3833);
nor U5228 (N_5228,N_4661,N_4379);
nor U5229 (N_5229,N_4473,N_3769);
nand U5230 (N_5230,N_4568,N_3815);
or U5231 (N_5231,N_4151,N_3832);
and U5232 (N_5232,N_4028,N_3917);
nor U5233 (N_5233,N_4545,N_3757);
and U5234 (N_5234,N_4827,N_3938);
xnor U5235 (N_5235,N_4748,N_3884);
and U5236 (N_5236,N_4576,N_4232);
xor U5237 (N_5237,N_4234,N_3955);
nand U5238 (N_5238,N_4841,N_4245);
or U5239 (N_5239,N_4186,N_4743);
nand U5240 (N_5240,N_4422,N_3778);
nand U5241 (N_5241,N_3867,N_3836);
or U5242 (N_5242,N_4195,N_4619);
or U5243 (N_5243,N_4901,N_4276);
nand U5244 (N_5244,N_4585,N_4828);
nand U5245 (N_5245,N_4090,N_4756);
nand U5246 (N_5246,N_4382,N_4502);
xnor U5247 (N_5247,N_4503,N_4351);
or U5248 (N_5248,N_4538,N_4851);
nor U5249 (N_5249,N_3997,N_4089);
nor U5250 (N_5250,N_4238,N_4728);
or U5251 (N_5251,N_4752,N_4256);
and U5252 (N_5252,N_4494,N_4730);
nand U5253 (N_5253,N_3862,N_3887);
and U5254 (N_5254,N_4056,N_3961);
xor U5255 (N_5255,N_4038,N_3859);
nor U5256 (N_5256,N_4359,N_4387);
nor U5257 (N_5257,N_4867,N_4397);
nand U5258 (N_5258,N_4782,N_4478);
xor U5259 (N_5259,N_4468,N_4580);
nor U5260 (N_5260,N_4584,N_4156);
or U5261 (N_5261,N_4785,N_4447);
and U5262 (N_5262,N_4677,N_4242);
nand U5263 (N_5263,N_4788,N_4286);
nor U5264 (N_5264,N_4223,N_4942);
and U5265 (N_5265,N_4998,N_4786);
or U5266 (N_5266,N_3939,N_4039);
and U5267 (N_5267,N_3844,N_3752);
nor U5268 (N_5268,N_4809,N_4991);
nand U5269 (N_5269,N_4928,N_4953);
and U5270 (N_5270,N_4634,N_4019);
or U5271 (N_5271,N_4114,N_3803);
or U5272 (N_5272,N_4191,N_4655);
nor U5273 (N_5273,N_3865,N_4762);
or U5274 (N_5274,N_4891,N_4184);
or U5275 (N_5275,N_4946,N_4082);
or U5276 (N_5276,N_4329,N_4871);
and U5277 (N_5277,N_4531,N_3881);
or U5278 (N_5278,N_4438,N_4471);
and U5279 (N_5279,N_4604,N_4870);
nor U5280 (N_5280,N_4664,N_4356);
and U5281 (N_5281,N_4738,N_4225);
and U5282 (N_5282,N_4332,N_4614);
nand U5283 (N_5283,N_4298,N_3827);
nor U5284 (N_5284,N_4622,N_4278);
nand U5285 (N_5285,N_3857,N_4905);
or U5286 (N_5286,N_4740,N_4408);
xor U5287 (N_5287,N_4649,N_4807);
nor U5288 (N_5288,N_4878,N_4853);
xnor U5289 (N_5289,N_4720,N_4916);
nor U5290 (N_5290,N_4579,N_3821);
nor U5291 (N_5291,N_4348,N_4719);
nand U5292 (N_5292,N_4394,N_4884);
or U5293 (N_5293,N_4006,N_3950);
nor U5294 (N_5294,N_3754,N_4410);
or U5295 (N_5295,N_4919,N_4505);
and U5296 (N_5296,N_4375,N_4029);
xor U5297 (N_5297,N_3946,N_4425);
nor U5298 (N_5298,N_4265,N_4682);
or U5299 (N_5299,N_3804,N_4091);
or U5300 (N_5300,N_4275,N_4949);
and U5301 (N_5301,N_4964,N_3973);
nand U5302 (N_5302,N_3979,N_4507);
and U5303 (N_5303,N_4950,N_3820);
xnor U5304 (N_5304,N_4062,N_4488);
xor U5305 (N_5305,N_3966,N_4293);
xnor U5306 (N_5306,N_4035,N_4759);
nor U5307 (N_5307,N_4084,N_4973);
or U5308 (N_5308,N_4385,N_3894);
xnor U5309 (N_5309,N_4227,N_4591);
xnor U5310 (N_5310,N_4751,N_4388);
nor U5311 (N_5311,N_4761,N_4574);
or U5312 (N_5312,N_4706,N_3963);
xnor U5313 (N_5313,N_4462,N_4637);
xnor U5314 (N_5314,N_4497,N_4449);
nand U5315 (N_5315,N_3793,N_4372);
nand U5316 (N_5316,N_3951,N_3981);
nor U5317 (N_5317,N_4045,N_4501);
and U5318 (N_5318,N_4990,N_3949);
or U5319 (N_5319,N_3892,N_4128);
and U5320 (N_5320,N_4702,N_4409);
nand U5321 (N_5321,N_4244,N_4924);
nand U5322 (N_5322,N_3801,N_4854);
or U5323 (N_5323,N_4078,N_3900);
or U5324 (N_5324,N_3788,N_4779);
nor U5325 (N_5325,N_4675,N_4811);
nand U5326 (N_5326,N_4428,N_3838);
or U5327 (N_5327,N_4052,N_3890);
or U5328 (N_5328,N_4940,N_4051);
xor U5329 (N_5329,N_4284,N_4943);
and U5330 (N_5330,N_4453,N_4739);
nor U5331 (N_5331,N_3964,N_4166);
nor U5332 (N_5332,N_4469,N_3915);
or U5333 (N_5333,N_4110,N_4543);
nand U5334 (N_5334,N_4624,N_4995);
or U5335 (N_5335,N_4666,N_4852);
nand U5336 (N_5336,N_4120,N_4683);
and U5337 (N_5337,N_4448,N_3818);
and U5338 (N_5338,N_4904,N_3789);
and U5339 (N_5339,N_4590,N_4322);
nor U5340 (N_5340,N_4463,N_4476);
xor U5341 (N_5341,N_4024,N_3791);
or U5342 (N_5342,N_3954,N_4402);
and U5343 (N_5343,N_4837,N_4072);
nor U5344 (N_5344,N_4081,N_4968);
or U5345 (N_5345,N_4713,N_4175);
and U5346 (N_5346,N_4862,N_3787);
and U5347 (N_5347,N_4693,N_4398);
or U5348 (N_5348,N_4464,N_4630);
and U5349 (N_5349,N_3906,N_4392);
and U5350 (N_5350,N_4210,N_3993);
xnor U5351 (N_5351,N_4817,N_4806);
nor U5352 (N_5352,N_4437,N_4561);
or U5353 (N_5353,N_4732,N_4419);
xor U5354 (N_5354,N_4176,N_4308);
or U5355 (N_5355,N_4116,N_4933);
nor U5356 (N_5356,N_4350,N_4481);
or U5357 (N_5357,N_4178,N_4309);
nand U5358 (N_5358,N_4551,N_4118);
nand U5359 (N_5359,N_4484,N_4204);
and U5360 (N_5360,N_4095,N_4423);
nand U5361 (N_5361,N_4915,N_3920);
nor U5362 (N_5362,N_3839,N_4446);
nand U5363 (N_5363,N_4113,N_4876);
nand U5364 (N_5364,N_4840,N_4066);
nand U5365 (N_5365,N_4317,N_4326);
and U5366 (N_5366,N_4167,N_4859);
and U5367 (N_5367,N_4133,N_4659);
and U5368 (N_5368,N_4951,N_4783);
xor U5369 (N_5369,N_3956,N_4067);
nor U5370 (N_5370,N_4330,N_4927);
and U5371 (N_5371,N_3987,N_4560);
and U5372 (N_5372,N_4523,N_4274);
xor U5373 (N_5373,N_4101,N_4516);
and U5374 (N_5374,N_4412,N_4137);
and U5375 (N_5375,N_3852,N_3901);
nor U5376 (N_5376,N_4271,N_4042);
nand U5377 (N_5377,N_3933,N_4887);
nor U5378 (N_5378,N_3858,N_4672);
nand U5379 (N_5379,N_4784,N_4458);
and U5380 (N_5380,N_4429,N_4367);
nor U5381 (N_5381,N_3965,N_4513);
and U5382 (N_5382,N_4917,N_3816);
xor U5383 (N_5383,N_4801,N_4775);
nand U5384 (N_5384,N_4855,N_3846);
nor U5385 (N_5385,N_4710,N_3861);
or U5386 (N_5386,N_3869,N_4311);
xor U5387 (N_5387,N_4912,N_4820);
nand U5388 (N_5388,N_4764,N_4282);
and U5389 (N_5389,N_3776,N_4694);
xor U5390 (N_5390,N_4992,N_3876);
nand U5391 (N_5391,N_4250,N_4595);
and U5392 (N_5392,N_4872,N_4360);
or U5393 (N_5393,N_4711,N_4214);
xor U5394 (N_5394,N_4125,N_3907);
nor U5395 (N_5395,N_4930,N_4858);
or U5396 (N_5396,N_3947,N_4888);
nand U5397 (N_5397,N_4198,N_4616);
or U5398 (N_5398,N_3904,N_4277);
nand U5399 (N_5399,N_4987,N_3941);
nor U5400 (N_5400,N_4157,N_3853);
or U5401 (N_5401,N_4635,N_4134);
or U5402 (N_5402,N_4370,N_4957);
nand U5403 (N_5403,N_4903,N_4316);
nand U5404 (N_5404,N_4697,N_4302);
and U5405 (N_5405,N_4218,N_4975);
and U5406 (N_5406,N_4434,N_4583);
xor U5407 (N_5407,N_4825,N_4549);
nor U5408 (N_5408,N_4060,N_4131);
nor U5409 (N_5409,N_4049,N_3969);
xor U5410 (N_5410,N_3888,N_4831);
and U5411 (N_5411,N_3905,N_3934);
or U5412 (N_5412,N_4451,N_4726);
xnor U5413 (N_5413,N_4816,N_4436);
or U5414 (N_5414,N_4044,N_3962);
or U5415 (N_5415,N_4014,N_4313);
nand U5416 (N_5416,N_4774,N_4312);
or U5417 (N_5417,N_3943,N_4541);
nor U5418 (N_5418,N_4611,N_3984);
xnor U5419 (N_5419,N_4153,N_4735);
nor U5420 (N_5420,N_3823,N_4224);
or U5421 (N_5421,N_4803,N_3772);
nand U5422 (N_5422,N_4572,N_4031);
and U5423 (N_5423,N_4076,N_4391);
and U5424 (N_5424,N_4657,N_4236);
xnor U5425 (N_5425,N_4160,N_4662);
xor U5426 (N_5426,N_4812,N_4737);
xor U5427 (N_5427,N_3863,N_4154);
nor U5428 (N_5428,N_4132,N_4717);
xnor U5429 (N_5429,N_3824,N_4534);
nor U5430 (N_5430,N_3775,N_4701);
or U5431 (N_5431,N_4863,N_3927);
or U5432 (N_5432,N_4328,N_4141);
nor U5433 (N_5433,N_4461,N_3992);
nand U5434 (N_5434,N_4836,N_4443);
nand U5435 (N_5435,N_3898,N_4323);
nor U5436 (N_5436,N_4810,N_3800);
nor U5437 (N_5437,N_4036,N_3763);
and U5438 (N_5438,N_4061,N_4555);
and U5439 (N_5439,N_4220,N_3811);
nand U5440 (N_5440,N_4140,N_4542);
and U5441 (N_5441,N_4085,N_4773);
xnor U5442 (N_5442,N_4606,N_4325);
and U5443 (N_5443,N_4838,N_4709);
nand U5444 (N_5444,N_4886,N_3960);
nor U5445 (N_5445,N_4763,N_4979);
and U5446 (N_5446,N_3916,N_4948);
nor U5447 (N_5447,N_4914,N_4165);
or U5448 (N_5448,N_4935,N_4866);
nor U5449 (N_5449,N_3983,N_4378);
xnor U5450 (N_5450,N_4802,N_4194);
or U5451 (N_5451,N_4980,N_4639);
nor U5452 (N_5452,N_4766,N_4499);
xor U5453 (N_5453,N_4487,N_4548);
xor U5454 (N_5454,N_4001,N_4117);
nor U5455 (N_5455,N_4627,N_4923);
or U5456 (N_5456,N_4922,N_4149);
nor U5457 (N_5457,N_4037,N_4063);
and U5458 (N_5458,N_4959,N_3766);
nor U5459 (N_5459,N_4296,N_4407);
nor U5460 (N_5460,N_4625,N_4559);
xnor U5461 (N_5461,N_3799,N_4179);
xnor U5462 (N_5462,N_4673,N_3866);
nand U5463 (N_5463,N_4399,N_3980);
nor U5464 (N_5464,N_4895,N_4222);
nand U5465 (N_5465,N_3760,N_3925);
nor U5466 (N_5466,N_4235,N_4517);
and U5467 (N_5467,N_3842,N_4822);
or U5468 (N_5468,N_4150,N_4102);
or U5469 (N_5469,N_4650,N_4602);
and U5470 (N_5470,N_4070,N_3829);
or U5471 (N_5471,N_4823,N_3871);
nand U5472 (N_5472,N_4833,N_3971);
and U5473 (N_5473,N_4281,N_4486);
or U5474 (N_5474,N_4219,N_4703);
nand U5475 (N_5475,N_4364,N_4778);
xnor U5476 (N_5476,N_3918,N_4474);
xor U5477 (N_5477,N_4537,N_3975);
xnor U5478 (N_5478,N_4636,N_4104);
or U5479 (N_5479,N_4386,N_4593);
or U5480 (N_5480,N_4107,N_3813);
nand U5481 (N_5481,N_4342,N_4355);
or U5482 (N_5482,N_4248,N_4377);
nor U5483 (N_5483,N_4148,N_4716);
xnor U5484 (N_5484,N_4470,N_4257);
xnor U5485 (N_5485,N_4093,N_3912);
xnor U5486 (N_5486,N_4515,N_3851);
nand U5487 (N_5487,N_4002,N_4495);
or U5488 (N_5488,N_3814,N_4246);
nor U5489 (N_5489,N_3825,N_4601);
xnor U5490 (N_5490,N_4566,N_4403);
or U5491 (N_5491,N_4251,N_3940);
and U5492 (N_5492,N_4522,N_4652);
xor U5493 (N_5493,N_4362,N_4240);
and U5494 (N_5494,N_4383,N_3873);
xnor U5495 (N_5495,N_4074,N_4097);
nand U5496 (N_5496,N_4795,N_3856);
and U5497 (N_5497,N_4644,N_4592);
nor U5498 (N_5498,N_4873,N_4600);
nand U5499 (N_5499,N_4539,N_3995);
nor U5500 (N_5500,N_4690,N_4881);
xnor U5501 (N_5501,N_4230,N_4967);
and U5502 (N_5502,N_4520,N_4707);
nand U5503 (N_5503,N_4411,N_4395);
nand U5504 (N_5504,N_4845,N_3819);
nand U5505 (N_5505,N_4441,N_4772);
nor U5506 (N_5506,N_4645,N_4830);
and U5507 (N_5507,N_4765,N_4944);
and U5508 (N_5508,N_4999,N_4754);
xnor U5509 (N_5509,N_4380,N_3982);
nand U5510 (N_5510,N_3874,N_3878);
and U5511 (N_5511,N_4440,N_3784);
nor U5512 (N_5512,N_4310,N_4890);
xor U5513 (N_5513,N_3985,N_4444);
nor U5514 (N_5514,N_4187,N_4005);
xor U5515 (N_5515,N_4741,N_4874);
xor U5516 (N_5516,N_3959,N_4144);
xor U5517 (N_5517,N_4978,N_4718);
xnor U5518 (N_5518,N_4012,N_4010);
xnor U5519 (N_5519,N_4196,N_3921);
xor U5520 (N_5520,N_4371,N_4416);
xnor U5521 (N_5521,N_3780,N_4808);
and U5522 (N_5522,N_4956,N_4705);
xnor U5523 (N_5523,N_4918,N_3902);
nand U5524 (N_5524,N_4135,N_3767);
or U5525 (N_5525,N_4164,N_3847);
nor U5526 (N_5526,N_4573,N_4793);
and U5527 (N_5527,N_4747,N_4780);
xnor U5528 (N_5528,N_4668,N_3986);
nand U5529 (N_5529,N_4349,N_3758);
xnor U5530 (N_5530,N_4626,N_4064);
or U5531 (N_5531,N_4115,N_4598);
and U5532 (N_5532,N_4932,N_3872);
nand U5533 (N_5533,N_4696,N_3977);
and U5534 (N_5534,N_4071,N_4365);
nor U5535 (N_5535,N_3875,N_4882);
or U5536 (N_5536,N_4714,N_4472);
nand U5537 (N_5537,N_4452,N_4926);
nand U5538 (N_5538,N_4109,N_4578);
xnor U5539 (N_5539,N_4000,N_4247);
xnor U5540 (N_5540,N_4270,N_3750);
nor U5541 (N_5541,N_3976,N_4913);
and U5542 (N_5542,N_4665,N_4781);
xor U5543 (N_5543,N_4997,N_4864);
nand U5544 (N_5544,N_4413,N_4509);
or U5545 (N_5545,N_4818,N_4124);
nor U5546 (N_5546,N_4427,N_4947);
nand U5547 (N_5547,N_3870,N_4952);
xor U5548 (N_5548,N_4856,N_4465);
or U5549 (N_5549,N_4475,N_4791);
and U5550 (N_5550,N_4289,N_4346);
and U5551 (N_5551,N_4454,N_4088);
xor U5552 (N_5552,N_4103,N_3885);
xor U5553 (N_5553,N_4849,N_4415);
xor U5554 (N_5554,N_4969,N_4899);
and U5555 (N_5555,N_4771,N_4170);
or U5556 (N_5556,N_4459,N_4877);
xor U5557 (N_5557,N_4804,N_4524);
nand U5558 (N_5558,N_4417,N_3895);
xor U5559 (N_5559,N_3994,N_4621);
and U5560 (N_5560,N_4173,N_4755);
nand U5561 (N_5561,N_4680,N_4239);
and U5562 (N_5562,N_3809,N_4504);
and U5563 (N_5563,N_3786,N_4489);
xnor U5564 (N_5564,N_4305,N_4381);
or U5565 (N_5565,N_3893,N_4963);
nand U5566 (N_5566,N_3999,N_4552);
and U5567 (N_5567,N_4172,N_4869);
xor U5568 (N_5568,N_4258,N_4357);
nand U5569 (N_5569,N_4016,N_4984);
nor U5570 (N_5570,N_4698,N_4835);
and U5571 (N_5571,N_4753,N_4656);
and U5572 (N_5572,N_4418,N_4231);
and U5573 (N_5573,N_4629,N_4424);
xor U5574 (N_5574,N_4030,N_3931);
or U5575 (N_5575,N_4880,N_4789);
and U5576 (N_5576,N_3850,N_4100);
xnor U5577 (N_5577,N_4421,N_4857);
or U5578 (N_5578,N_4512,N_4970);
nand U5579 (N_5579,N_4721,N_4337);
or U5580 (N_5580,N_4892,N_4285);
and U5581 (N_5581,N_4613,N_4570);
nor U5582 (N_5582,N_3911,N_4525);
and U5583 (N_5583,N_4594,N_4163);
xor U5584 (N_5584,N_4983,N_4563);
nand U5585 (N_5585,N_4053,N_4142);
and U5586 (N_5586,N_4263,N_4734);
and U5587 (N_5587,N_4022,N_4898);
nand U5588 (N_5588,N_4203,N_4628);
nand U5589 (N_5589,N_4847,N_4158);
nand U5590 (N_5590,N_3781,N_4691);
xnor U5591 (N_5591,N_4267,N_4057);
and U5592 (N_5592,N_4108,N_3924);
nand U5593 (N_5593,N_4550,N_4925);
xnor U5594 (N_5594,N_4977,N_3783);
and U5595 (N_5595,N_4794,N_4043);
nand U5596 (N_5596,N_3828,N_4460);
xor U5597 (N_5597,N_4832,N_4456);
nor U5598 (N_5598,N_4961,N_3974);
and U5599 (N_5599,N_4790,N_4373);
xor U5600 (N_5600,N_4430,N_4586);
nor U5601 (N_5601,N_4007,N_4200);
nand U5602 (N_5602,N_4174,N_4393);
or U5603 (N_5603,N_4770,N_3929);
xor U5604 (N_5604,N_3810,N_4335);
or U5605 (N_5605,N_4073,N_4477);
nor U5606 (N_5606,N_4679,N_4254);
or U5607 (N_5607,N_4185,N_4571);
nor U5608 (N_5608,N_4123,N_4988);
and U5609 (N_5609,N_4004,N_4366);
nor U5610 (N_5610,N_4098,N_4280);
or U5611 (N_5611,N_4844,N_4139);
or U5612 (N_5612,N_4493,N_4404);
xor U5613 (N_5613,N_3909,N_4907);
xnor U5614 (N_5614,N_4111,N_4283);
nand U5615 (N_5615,N_4535,N_3835);
and U5616 (N_5616,N_4511,N_4536);
and U5617 (N_5617,N_3903,N_4126);
nand U5618 (N_5618,N_4993,N_4599);
nand U5619 (N_5619,N_4532,N_4729);
nor U5620 (N_5620,N_4345,N_4506);
xor U5621 (N_5621,N_4526,N_4211);
nand U5622 (N_5622,N_4623,N_4241);
nor U5623 (N_5623,N_4152,N_4792);
xnor U5624 (N_5624,N_4059,N_4632);
xnor U5625 (N_5625,N_4675,N_4039);
and U5626 (N_5626,N_4296,N_4490);
nor U5627 (N_5627,N_4604,N_4296);
or U5628 (N_5628,N_4111,N_3908);
xor U5629 (N_5629,N_4090,N_4913);
or U5630 (N_5630,N_4814,N_4869);
nor U5631 (N_5631,N_4822,N_4705);
and U5632 (N_5632,N_3899,N_3954);
xnor U5633 (N_5633,N_4348,N_4652);
nor U5634 (N_5634,N_4227,N_4493);
or U5635 (N_5635,N_4306,N_4862);
and U5636 (N_5636,N_4736,N_4608);
and U5637 (N_5637,N_4864,N_4988);
xnor U5638 (N_5638,N_4046,N_3937);
and U5639 (N_5639,N_4434,N_4224);
nand U5640 (N_5640,N_4165,N_4760);
xnor U5641 (N_5641,N_4590,N_3961);
and U5642 (N_5642,N_4445,N_4312);
or U5643 (N_5643,N_4983,N_4604);
xor U5644 (N_5644,N_4692,N_4456);
xnor U5645 (N_5645,N_3753,N_4773);
xnor U5646 (N_5646,N_4717,N_4173);
nor U5647 (N_5647,N_4813,N_4145);
nand U5648 (N_5648,N_4144,N_4089);
or U5649 (N_5649,N_4137,N_4447);
nor U5650 (N_5650,N_4905,N_4132);
or U5651 (N_5651,N_4546,N_3936);
nor U5652 (N_5652,N_4682,N_4150);
nand U5653 (N_5653,N_4580,N_3924);
and U5654 (N_5654,N_4943,N_4898);
xnor U5655 (N_5655,N_4869,N_4730);
or U5656 (N_5656,N_3851,N_4581);
xor U5657 (N_5657,N_4401,N_3975);
and U5658 (N_5658,N_4700,N_4305);
xor U5659 (N_5659,N_4089,N_4383);
xor U5660 (N_5660,N_4652,N_4870);
and U5661 (N_5661,N_4687,N_4371);
or U5662 (N_5662,N_4097,N_4251);
or U5663 (N_5663,N_3957,N_4409);
and U5664 (N_5664,N_3858,N_4808);
nor U5665 (N_5665,N_4392,N_4863);
and U5666 (N_5666,N_3787,N_4043);
nand U5667 (N_5667,N_4094,N_3803);
nor U5668 (N_5668,N_4033,N_3845);
nor U5669 (N_5669,N_4581,N_3967);
and U5670 (N_5670,N_4355,N_4962);
nor U5671 (N_5671,N_4756,N_3843);
xnor U5672 (N_5672,N_3908,N_4027);
nor U5673 (N_5673,N_4262,N_3911);
xor U5674 (N_5674,N_4985,N_3930);
and U5675 (N_5675,N_4333,N_3903);
and U5676 (N_5676,N_3917,N_3952);
nor U5677 (N_5677,N_4433,N_4029);
nand U5678 (N_5678,N_4285,N_4510);
and U5679 (N_5679,N_4931,N_4014);
or U5680 (N_5680,N_4243,N_4880);
or U5681 (N_5681,N_4162,N_4541);
and U5682 (N_5682,N_4036,N_4056);
or U5683 (N_5683,N_4385,N_4163);
nand U5684 (N_5684,N_4721,N_4127);
and U5685 (N_5685,N_4222,N_4392);
xnor U5686 (N_5686,N_4825,N_4632);
nand U5687 (N_5687,N_4584,N_4547);
and U5688 (N_5688,N_3989,N_4073);
xnor U5689 (N_5689,N_4197,N_4335);
or U5690 (N_5690,N_4235,N_4736);
or U5691 (N_5691,N_4323,N_4095);
nor U5692 (N_5692,N_3775,N_4294);
xnor U5693 (N_5693,N_4564,N_4279);
nor U5694 (N_5694,N_4491,N_4245);
xor U5695 (N_5695,N_4988,N_4792);
nor U5696 (N_5696,N_4190,N_4569);
nand U5697 (N_5697,N_4588,N_4669);
nand U5698 (N_5698,N_4122,N_4288);
and U5699 (N_5699,N_4634,N_4034);
or U5700 (N_5700,N_4171,N_3829);
nor U5701 (N_5701,N_3957,N_3944);
nand U5702 (N_5702,N_4353,N_4525);
nor U5703 (N_5703,N_4474,N_4469);
nand U5704 (N_5704,N_4481,N_4142);
or U5705 (N_5705,N_4009,N_4724);
xor U5706 (N_5706,N_4738,N_4811);
nand U5707 (N_5707,N_4851,N_4917);
nand U5708 (N_5708,N_3948,N_4261);
nor U5709 (N_5709,N_4004,N_4377);
xor U5710 (N_5710,N_4585,N_4916);
xnor U5711 (N_5711,N_4959,N_4569);
nor U5712 (N_5712,N_4332,N_4879);
xnor U5713 (N_5713,N_4831,N_4944);
or U5714 (N_5714,N_4015,N_4804);
nor U5715 (N_5715,N_4875,N_4410);
or U5716 (N_5716,N_3923,N_4621);
xor U5717 (N_5717,N_4237,N_4360);
and U5718 (N_5718,N_4381,N_4253);
xnor U5719 (N_5719,N_4436,N_4790);
xnor U5720 (N_5720,N_3978,N_4010);
nand U5721 (N_5721,N_4567,N_3776);
and U5722 (N_5722,N_4566,N_4548);
nor U5723 (N_5723,N_3996,N_4722);
nor U5724 (N_5724,N_4581,N_4350);
xnor U5725 (N_5725,N_4191,N_4550);
nor U5726 (N_5726,N_4992,N_4151);
and U5727 (N_5727,N_4229,N_3972);
nand U5728 (N_5728,N_3851,N_4011);
nand U5729 (N_5729,N_4493,N_4503);
xor U5730 (N_5730,N_4819,N_3938);
nor U5731 (N_5731,N_3819,N_4293);
nor U5732 (N_5732,N_3971,N_3965);
and U5733 (N_5733,N_4409,N_4376);
nand U5734 (N_5734,N_4595,N_4599);
or U5735 (N_5735,N_4674,N_4535);
xnor U5736 (N_5736,N_4079,N_4184);
xor U5737 (N_5737,N_4423,N_3781);
and U5738 (N_5738,N_4581,N_4536);
nand U5739 (N_5739,N_4977,N_4253);
xnor U5740 (N_5740,N_4597,N_4959);
nor U5741 (N_5741,N_4807,N_4863);
xnor U5742 (N_5742,N_4262,N_4075);
nand U5743 (N_5743,N_4657,N_4243);
and U5744 (N_5744,N_4780,N_4937);
and U5745 (N_5745,N_3872,N_4145);
nor U5746 (N_5746,N_4108,N_4900);
xnor U5747 (N_5747,N_4370,N_4748);
nand U5748 (N_5748,N_3810,N_4191);
and U5749 (N_5749,N_4125,N_4686);
and U5750 (N_5750,N_4836,N_4784);
xor U5751 (N_5751,N_4499,N_3765);
nand U5752 (N_5752,N_3913,N_3770);
nor U5753 (N_5753,N_4225,N_4008);
xnor U5754 (N_5754,N_4487,N_4984);
xor U5755 (N_5755,N_4511,N_4488);
xor U5756 (N_5756,N_3997,N_4050);
and U5757 (N_5757,N_4093,N_4988);
xnor U5758 (N_5758,N_3799,N_4096);
and U5759 (N_5759,N_4996,N_4136);
and U5760 (N_5760,N_4289,N_4724);
nor U5761 (N_5761,N_4361,N_4419);
xor U5762 (N_5762,N_3876,N_3816);
xnor U5763 (N_5763,N_4118,N_4280);
xnor U5764 (N_5764,N_3923,N_4746);
and U5765 (N_5765,N_3991,N_4663);
or U5766 (N_5766,N_4287,N_4480);
or U5767 (N_5767,N_4096,N_4843);
nor U5768 (N_5768,N_3983,N_4412);
nor U5769 (N_5769,N_4386,N_3960);
xor U5770 (N_5770,N_4901,N_4031);
xnor U5771 (N_5771,N_4655,N_4764);
or U5772 (N_5772,N_4820,N_4218);
xnor U5773 (N_5773,N_4647,N_4683);
nand U5774 (N_5774,N_4091,N_4403);
xor U5775 (N_5775,N_4874,N_4270);
or U5776 (N_5776,N_4417,N_4817);
nor U5777 (N_5777,N_4499,N_4682);
nand U5778 (N_5778,N_4431,N_4537);
or U5779 (N_5779,N_4953,N_4215);
and U5780 (N_5780,N_4130,N_4968);
nor U5781 (N_5781,N_3907,N_4497);
xnor U5782 (N_5782,N_4664,N_4004);
xnor U5783 (N_5783,N_4772,N_3774);
or U5784 (N_5784,N_4504,N_4016);
nor U5785 (N_5785,N_4993,N_4696);
xnor U5786 (N_5786,N_4801,N_4371);
nor U5787 (N_5787,N_4164,N_4904);
nand U5788 (N_5788,N_4218,N_3801);
and U5789 (N_5789,N_4416,N_4264);
or U5790 (N_5790,N_4999,N_4955);
and U5791 (N_5791,N_3813,N_4745);
nand U5792 (N_5792,N_4165,N_4513);
xor U5793 (N_5793,N_4183,N_4336);
or U5794 (N_5794,N_4914,N_4436);
and U5795 (N_5795,N_4872,N_4919);
nand U5796 (N_5796,N_4825,N_3806);
or U5797 (N_5797,N_4890,N_4988);
nor U5798 (N_5798,N_4336,N_4602);
and U5799 (N_5799,N_3804,N_4024);
nand U5800 (N_5800,N_4471,N_4545);
or U5801 (N_5801,N_4926,N_4995);
or U5802 (N_5802,N_3775,N_3853);
nand U5803 (N_5803,N_3984,N_4005);
and U5804 (N_5804,N_3954,N_4028);
nand U5805 (N_5805,N_4485,N_4821);
xor U5806 (N_5806,N_4307,N_4004);
or U5807 (N_5807,N_4334,N_3922);
or U5808 (N_5808,N_4511,N_4799);
or U5809 (N_5809,N_3979,N_4501);
or U5810 (N_5810,N_4454,N_4749);
nor U5811 (N_5811,N_4329,N_3901);
or U5812 (N_5812,N_4496,N_4547);
nor U5813 (N_5813,N_4038,N_4159);
nand U5814 (N_5814,N_4718,N_4976);
nand U5815 (N_5815,N_4668,N_4311);
nand U5816 (N_5816,N_4049,N_4489);
or U5817 (N_5817,N_4060,N_4029);
and U5818 (N_5818,N_3773,N_4457);
or U5819 (N_5819,N_3905,N_3845);
nor U5820 (N_5820,N_4366,N_3937);
xor U5821 (N_5821,N_4568,N_4121);
nor U5822 (N_5822,N_4625,N_4196);
or U5823 (N_5823,N_3772,N_4559);
nor U5824 (N_5824,N_3783,N_4801);
xor U5825 (N_5825,N_3928,N_3849);
nor U5826 (N_5826,N_4639,N_4884);
or U5827 (N_5827,N_4061,N_4852);
xnor U5828 (N_5828,N_3794,N_3984);
xor U5829 (N_5829,N_3830,N_4718);
nand U5830 (N_5830,N_3803,N_4182);
nor U5831 (N_5831,N_4613,N_3757);
xor U5832 (N_5832,N_4153,N_4389);
xnor U5833 (N_5833,N_4047,N_4619);
xnor U5834 (N_5834,N_4159,N_3777);
xnor U5835 (N_5835,N_3781,N_4325);
xnor U5836 (N_5836,N_4027,N_4094);
nor U5837 (N_5837,N_4569,N_4382);
xor U5838 (N_5838,N_3900,N_3940);
nand U5839 (N_5839,N_4689,N_3930);
and U5840 (N_5840,N_3932,N_4661);
xor U5841 (N_5841,N_4865,N_4608);
nor U5842 (N_5842,N_3831,N_4242);
nor U5843 (N_5843,N_4667,N_4623);
or U5844 (N_5844,N_4570,N_4307);
nand U5845 (N_5845,N_4284,N_4730);
or U5846 (N_5846,N_4961,N_4716);
nor U5847 (N_5847,N_3901,N_4992);
nand U5848 (N_5848,N_4044,N_4388);
or U5849 (N_5849,N_4696,N_4235);
nand U5850 (N_5850,N_4114,N_4459);
nor U5851 (N_5851,N_4363,N_4737);
xnor U5852 (N_5852,N_4955,N_4695);
or U5853 (N_5853,N_4121,N_4214);
nand U5854 (N_5854,N_3950,N_3974);
or U5855 (N_5855,N_4200,N_4261);
nand U5856 (N_5856,N_4877,N_4045);
or U5857 (N_5857,N_4027,N_4244);
and U5858 (N_5858,N_4336,N_4865);
xor U5859 (N_5859,N_4456,N_3981);
nor U5860 (N_5860,N_4960,N_4711);
nand U5861 (N_5861,N_4343,N_4936);
or U5862 (N_5862,N_4740,N_4072);
nor U5863 (N_5863,N_4883,N_4275);
nand U5864 (N_5864,N_3907,N_4863);
nand U5865 (N_5865,N_4109,N_3852);
nor U5866 (N_5866,N_4649,N_3968);
and U5867 (N_5867,N_4246,N_3909);
nor U5868 (N_5868,N_4583,N_4560);
nor U5869 (N_5869,N_4915,N_4277);
and U5870 (N_5870,N_4946,N_4277);
xnor U5871 (N_5871,N_4457,N_4834);
or U5872 (N_5872,N_4331,N_4889);
or U5873 (N_5873,N_4366,N_4546);
or U5874 (N_5874,N_4626,N_3792);
nand U5875 (N_5875,N_3782,N_3893);
and U5876 (N_5876,N_4217,N_3976);
or U5877 (N_5877,N_4191,N_3936);
nand U5878 (N_5878,N_4122,N_4608);
and U5879 (N_5879,N_4202,N_4176);
or U5880 (N_5880,N_4224,N_4192);
nor U5881 (N_5881,N_4178,N_4218);
nand U5882 (N_5882,N_4982,N_4885);
nor U5883 (N_5883,N_3941,N_4197);
xor U5884 (N_5884,N_4797,N_3865);
nor U5885 (N_5885,N_4612,N_4702);
and U5886 (N_5886,N_4291,N_3840);
and U5887 (N_5887,N_3833,N_4425);
xnor U5888 (N_5888,N_4924,N_3952);
nor U5889 (N_5889,N_4783,N_4258);
xor U5890 (N_5890,N_4831,N_4528);
nand U5891 (N_5891,N_4065,N_4069);
nand U5892 (N_5892,N_4621,N_4054);
nor U5893 (N_5893,N_4388,N_4758);
xor U5894 (N_5894,N_4323,N_4017);
nand U5895 (N_5895,N_3904,N_4773);
nor U5896 (N_5896,N_4691,N_4965);
nor U5897 (N_5897,N_4923,N_4022);
and U5898 (N_5898,N_4843,N_4431);
nand U5899 (N_5899,N_3807,N_4163);
and U5900 (N_5900,N_4765,N_4630);
or U5901 (N_5901,N_4676,N_4589);
xor U5902 (N_5902,N_4419,N_4701);
xor U5903 (N_5903,N_3928,N_4967);
nor U5904 (N_5904,N_4337,N_4180);
xor U5905 (N_5905,N_3804,N_4667);
and U5906 (N_5906,N_3822,N_4754);
and U5907 (N_5907,N_4637,N_3929);
and U5908 (N_5908,N_4399,N_4890);
nor U5909 (N_5909,N_3825,N_4864);
or U5910 (N_5910,N_4879,N_4712);
xnor U5911 (N_5911,N_4795,N_3992);
and U5912 (N_5912,N_4838,N_4253);
xnor U5913 (N_5913,N_4384,N_4310);
and U5914 (N_5914,N_3935,N_4785);
and U5915 (N_5915,N_4795,N_4662);
nor U5916 (N_5916,N_4666,N_4458);
nand U5917 (N_5917,N_4956,N_4281);
or U5918 (N_5918,N_4493,N_4960);
nand U5919 (N_5919,N_4152,N_4360);
or U5920 (N_5920,N_4026,N_4999);
nor U5921 (N_5921,N_3873,N_4994);
nor U5922 (N_5922,N_4471,N_4190);
nor U5923 (N_5923,N_4148,N_3917);
or U5924 (N_5924,N_4783,N_3992);
or U5925 (N_5925,N_4800,N_4886);
or U5926 (N_5926,N_3827,N_4525);
or U5927 (N_5927,N_4403,N_3897);
and U5928 (N_5928,N_3836,N_4875);
nand U5929 (N_5929,N_4778,N_3894);
xnor U5930 (N_5930,N_4637,N_4325);
or U5931 (N_5931,N_4009,N_4483);
xnor U5932 (N_5932,N_4044,N_4462);
or U5933 (N_5933,N_4658,N_4822);
nand U5934 (N_5934,N_4601,N_4905);
nand U5935 (N_5935,N_4364,N_4860);
and U5936 (N_5936,N_4923,N_4065);
nand U5937 (N_5937,N_3875,N_3788);
xor U5938 (N_5938,N_4443,N_4951);
nor U5939 (N_5939,N_4404,N_3797);
or U5940 (N_5940,N_4462,N_4100);
or U5941 (N_5941,N_4280,N_4643);
nor U5942 (N_5942,N_4965,N_4943);
xnor U5943 (N_5943,N_4031,N_4695);
xor U5944 (N_5944,N_4863,N_4716);
nand U5945 (N_5945,N_3906,N_4327);
nor U5946 (N_5946,N_4354,N_4213);
and U5947 (N_5947,N_4216,N_4825);
and U5948 (N_5948,N_4861,N_4836);
and U5949 (N_5949,N_4797,N_3848);
nor U5950 (N_5950,N_4350,N_4125);
nor U5951 (N_5951,N_3875,N_4803);
nor U5952 (N_5952,N_4636,N_3976);
or U5953 (N_5953,N_3762,N_4271);
nor U5954 (N_5954,N_4395,N_4765);
or U5955 (N_5955,N_4354,N_4076);
xor U5956 (N_5956,N_4465,N_4418);
or U5957 (N_5957,N_4463,N_4612);
or U5958 (N_5958,N_4559,N_4214);
nand U5959 (N_5959,N_4214,N_4538);
or U5960 (N_5960,N_4260,N_3874);
or U5961 (N_5961,N_4555,N_4608);
or U5962 (N_5962,N_4362,N_4726);
or U5963 (N_5963,N_4849,N_4247);
nand U5964 (N_5964,N_4202,N_4883);
and U5965 (N_5965,N_4291,N_4294);
nand U5966 (N_5966,N_4391,N_4933);
nand U5967 (N_5967,N_4410,N_4245);
xnor U5968 (N_5968,N_4027,N_3963);
or U5969 (N_5969,N_3994,N_4754);
xnor U5970 (N_5970,N_4470,N_4950);
nor U5971 (N_5971,N_4713,N_3951);
xnor U5972 (N_5972,N_4522,N_4716);
and U5973 (N_5973,N_4442,N_4931);
or U5974 (N_5974,N_4246,N_4315);
nor U5975 (N_5975,N_4893,N_4855);
or U5976 (N_5976,N_3791,N_3820);
xnor U5977 (N_5977,N_3933,N_4826);
nor U5978 (N_5978,N_4304,N_4505);
and U5979 (N_5979,N_4099,N_4140);
or U5980 (N_5980,N_4218,N_3991);
nor U5981 (N_5981,N_3760,N_4008);
and U5982 (N_5982,N_4125,N_4254);
nand U5983 (N_5983,N_4954,N_3805);
nand U5984 (N_5984,N_4826,N_4691);
nand U5985 (N_5985,N_3990,N_4273);
and U5986 (N_5986,N_4148,N_3921);
nand U5987 (N_5987,N_4212,N_4252);
nand U5988 (N_5988,N_4560,N_3913);
nand U5989 (N_5989,N_4563,N_4994);
nand U5990 (N_5990,N_4500,N_4785);
xor U5991 (N_5991,N_4348,N_3968);
nor U5992 (N_5992,N_3798,N_4199);
nand U5993 (N_5993,N_4694,N_4570);
and U5994 (N_5994,N_4112,N_4230);
xor U5995 (N_5995,N_3954,N_4465);
or U5996 (N_5996,N_3863,N_3952);
and U5997 (N_5997,N_4412,N_4112);
nand U5998 (N_5998,N_4874,N_4947);
or U5999 (N_5999,N_4255,N_4879);
xor U6000 (N_6000,N_4745,N_4727);
and U6001 (N_6001,N_4654,N_3767);
and U6002 (N_6002,N_4366,N_4341);
and U6003 (N_6003,N_4418,N_4526);
xor U6004 (N_6004,N_3789,N_3766);
or U6005 (N_6005,N_3863,N_4999);
xnor U6006 (N_6006,N_4292,N_4122);
xor U6007 (N_6007,N_4515,N_4141);
or U6008 (N_6008,N_4056,N_3771);
and U6009 (N_6009,N_4376,N_4800);
and U6010 (N_6010,N_3964,N_4357);
nand U6011 (N_6011,N_4883,N_4436);
and U6012 (N_6012,N_3770,N_4153);
nor U6013 (N_6013,N_4908,N_4525);
xnor U6014 (N_6014,N_4713,N_4932);
nand U6015 (N_6015,N_4555,N_4912);
xnor U6016 (N_6016,N_3813,N_4488);
and U6017 (N_6017,N_4553,N_4935);
and U6018 (N_6018,N_4429,N_4323);
or U6019 (N_6019,N_4563,N_4269);
nor U6020 (N_6020,N_3806,N_4954);
and U6021 (N_6021,N_4884,N_3936);
nand U6022 (N_6022,N_4079,N_4246);
nand U6023 (N_6023,N_4943,N_4661);
xnor U6024 (N_6024,N_4204,N_3789);
nor U6025 (N_6025,N_4576,N_3911);
xor U6026 (N_6026,N_4541,N_3887);
nor U6027 (N_6027,N_4301,N_4962);
or U6028 (N_6028,N_4663,N_4919);
or U6029 (N_6029,N_4229,N_4510);
or U6030 (N_6030,N_4108,N_4825);
nor U6031 (N_6031,N_4722,N_3903);
nor U6032 (N_6032,N_4610,N_4611);
xnor U6033 (N_6033,N_4437,N_4259);
and U6034 (N_6034,N_4887,N_4101);
nor U6035 (N_6035,N_4445,N_3926);
nor U6036 (N_6036,N_4993,N_4509);
xnor U6037 (N_6037,N_4288,N_3800);
and U6038 (N_6038,N_4509,N_4308);
nand U6039 (N_6039,N_4470,N_3884);
or U6040 (N_6040,N_4852,N_3950);
or U6041 (N_6041,N_4721,N_4025);
xnor U6042 (N_6042,N_3874,N_4050);
nor U6043 (N_6043,N_4908,N_4064);
nand U6044 (N_6044,N_4868,N_4430);
or U6045 (N_6045,N_4318,N_4534);
nor U6046 (N_6046,N_4415,N_4599);
or U6047 (N_6047,N_4406,N_4490);
or U6048 (N_6048,N_4662,N_4211);
or U6049 (N_6049,N_4764,N_3816);
xnor U6050 (N_6050,N_4019,N_3799);
or U6051 (N_6051,N_3993,N_4480);
nor U6052 (N_6052,N_4005,N_3815);
xor U6053 (N_6053,N_4030,N_4275);
or U6054 (N_6054,N_4556,N_4511);
nand U6055 (N_6055,N_4721,N_4001);
or U6056 (N_6056,N_4073,N_4205);
nor U6057 (N_6057,N_3760,N_4628);
and U6058 (N_6058,N_4906,N_4957);
xnor U6059 (N_6059,N_4904,N_3864);
nor U6060 (N_6060,N_4523,N_4800);
nor U6061 (N_6061,N_4490,N_3786);
nand U6062 (N_6062,N_4671,N_4951);
and U6063 (N_6063,N_4536,N_4052);
nor U6064 (N_6064,N_4239,N_4901);
nand U6065 (N_6065,N_4352,N_3773);
xnor U6066 (N_6066,N_4842,N_4947);
nor U6067 (N_6067,N_4389,N_4508);
nand U6068 (N_6068,N_4996,N_4393);
and U6069 (N_6069,N_3983,N_4652);
or U6070 (N_6070,N_4110,N_4131);
or U6071 (N_6071,N_4118,N_4323);
or U6072 (N_6072,N_4590,N_4120);
or U6073 (N_6073,N_4210,N_4262);
xnor U6074 (N_6074,N_4930,N_4961);
or U6075 (N_6075,N_4300,N_4616);
xor U6076 (N_6076,N_4359,N_4640);
nor U6077 (N_6077,N_4381,N_4980);
nor U6078 (N_6078,N_4118,N_4318);
or U6079 (N_6079,N_3853,N_4772);
xnor U6080 (N_6080,N_4490,N_4440);
or U6081 (N_6081,N_4330,N_3883);
nor U6082 (N_6082,N_4130,N_4177);
or U6083 (N_6083,N_4766,N_4731);
nor U6084 (N_6084,N_4281,N_4398);
or U6085 (N_6085,N_4240,N_3940);
and U6086 (N_6086,N_4177,N_4545);
or U6087 (N_6087,N_3810,N_3828);
and U6088 (N_6088,N_4542,N_4361);
nor U6089 (N_6089,N_3783,N_4749);
and U6090 (N_6090,N_4366,N_3869);
xnor U6091 (N_6091,N_4905,N_4322);
or U6092 (N_6092,N_4927,N_3806);
nor U6093 (N_6093,N_4215,N_4609);
or U6094 (N_6094,N_4592,N_4873);
xor U6095 (N_6095,N_4066,N_3960);
or U6096 (N_6096,N_4411,N_4727);
xor U6097 (N_6097,N_4935,N_4537);
nor U6098 (N_6098,N_4419,N_4394);
nor U6099 (N_6099,N_4809,N_4228);
nor U6100 (N_6100,N_4483,N_4275);
nor U6101 (N_6101,N_4780,N_4029);
nand U6102 (N_6102,N_3777,N_4888);
nor U6103 (N_6103,N_4262,N_4224);
nand U6104 (N_6104,N_4604,N_3831);
nand U6105 (N_6105,N_4160,N_4625);
or U6106 (N_6106,N_4542,N_4607);
nor U6107 (N_6107,N_3974,N_3988);
or U6108 (N_6108,N_4670,N_4106);
nand U6109 (N_6109,N_4761,N_3818);
or U6110 (N_6110,N_4995,N_4463);
nor U6111 (N_6111,N_4675,N_3846);
xnor U6112 (N_6112,N_4552,N_4969);
or U6113 (N_6113,N_4395,N_4398);
xor U6114 (N_6114,N_4339,N_4344);
nor U6115 (N_6115,N_4408,N_4069);
and U6116 (N_6116,N_4036,N_4399);
xnor U6117 (N_6117,N_3931,N_3936);
xor U6118 (N_6118,N_4715,N_4854);
or U6119 (N_6119,N_4360,N_3765);
nand U6120 (N_6120,N_4029,N_4504);
nor U6121 (N_6121,N_4249,N_4273);
xor U6122 (N_6122,N_4876,N_3955);
nor U6123 (N_6123,N_4034,N_4388);
or U6124 (N_6124,N_3907,N_3815);
nor U6125 (N_6125,N_3801,N_4663);
or U6126 (N_6126,N_3790,N_4108);
nand U6127 (N_6127,N_3943,N_4495);
nand U6128 (N_6128,N_3840,N_4602);
nand U6129 (N_6129,N_4705,N_4773);
nor U6130 (N_6130,N_3988,N_4951);
nand U6131 (N_6131,N_4509,N_4603);
and U6132 (N_6132,N_4017,N_4078);
or U6133 (N_6133,N_4903,N_4536);
and U6134 (N_6134,N_4617,N_4277);
or U6135 (N_6135,N_3963,N_4496);
nor U6136 (N_6136,N_4662,N_4425);
or U6137 (N_6137,N_4546,N_4260);
and U6138 (N_6138,N_4456,N_4797);
xor U6139 (N_6139,N_4047,N_4974);
xnor U6140 (N_6140,N_4955,N_4143);
nand U6141 (N_6141,N_4521,N_4934);
and U6142 (N_6142,N_4476,N_3907);
and U6143 (N_6143,N_4790,N_3964);
and U6144 (N_6144,N_4222,N_4117);
nor U6145 (N_6145,N_4362,N_4289);
nand U6146 (N_6146,N_4597,N_4502);
and U6147 (N_6147,N_4898,N_4611);
nor U6148 (N_6148,N_3910,N_4667);
and U6149 (N_6149,N_4974,N_4980);
xor U6150 (N_6150,N_4757,N_4678);
nand U6151 (N_6151,N_3881,N_4276);
nor U6152 (N_6152,N_4607,N_3812);
or U6153 (N_6153,N_3945,N_4855);
nand U6154 (N_6154,N_4631,N_4077);
nor U6155 (N_6155,N_4480,N_3804);
or U6156 (N_6156,N_3828,N_4027);
and U6157 (N_6157,N_4007,N_3812);
xnor U6158 (N_6158,N_4496,N_4147);
and U6159 (N_6159,N_4645,N_4736);
xnor U6160 (N_6160,N_4698,N_4301);
or U6161 (N_6161,N_3877,N_4937);
and U6162 (N_6162,N_4237,N_4121);
or U6163 (N_6163,N_4274,N_4152);
or U6164 (N_6164,N_4461,N_4031);
xnor U6165 (N_6165,N_4487,N_3814);
xnor U6166 (N_6166,N_4540,N_4723);
or U6167 (N_6167,N_4901,N_3760);
and U6168 (N_6168,N_3985,N_4161);
xor U6169 (N_6169,N_4392,N_4265);
nand U6170 (N_6170,N_4076,N_4653);
or U6171 (N_6171,N_4882,N_4404);
nor U6172 (N_6172,N_4853,N_4176);
or U6173 (N_6173,N_3936,N_4389);
nor U6174 (N_6174,N_3940,N_4720);
and U6175 (N_6175,N_4636,N_4131);
xnor U6176 (N_6176,N_3763,N_4412);
xnor U6177 (N_6177,N_3981,N_4074);
or U6178 (N_6178,N_4611,N_4535);
or U6179 (N_6179,N_4955,N_4597);
xor U6180 (N_6180,N_4023,N_4111);
xor U6181 (N_6181,N_4463,N_4890);
nand U6182 (N_6182,N_4028,N_4017);
and U6183 (N_6183,N_4110,N_4072);
and U6184 (N_6184,N_4942,N_4181);
and U6185 (N_6185,N_4367,N_4503);
nor U6186 (N_6186,N_3950,N_4995);
xnor U6187 (N_6187,N_4344,N_4971);
nand U6188 (N_6188,N_4607,N_4716);
nor U6189 (N_6189,N_4019,N_4668);
nor U6190 (N_6190,N_3784,N_4103);
xor U6191 (N_6191,N_4306,N_4968);
xnor U6192 (N_6192,N_4979,N_4150);
and U6193 (N_6193,N_4427,N_3887);
or U6194 (N_6194,N_4566,N_4535);
and U6195 (N_6195,N_4704,N_4455);
and U6196 (N_6196,N_4162,N_4125);
and U6197 (N_6197,N_4400,N_4366);
and U6198 (N_6198,N_3902,N_4624);
or U6199 (N_6199,N_4131,N_3845);
nand U6200 (N_6200,N_4055,N_4996);
nand U6201 (N_6201,N_3930,N_4835);
nor U6202 (N_6202,N_4697,N_4456);
or U6203 (N_6203,N_4469,N_4985);
xnor U6204 (N_6204,N_4170,N_3829);
xnor U6205 (N_6205,N_4688,N_4690);
xor U6206 (N_6206,N_4393,N_4492);
and U6207 (N_6207,N_4643,N_4868);
nor U6208 (N_6208,N_4569,N_4135);
and U6209 (N_6209,N_4274,N_4671);
or U6210 (N_6210,N_4487,N_4164);
and U6211 (N_6211,N_3918,N_4943);
nor U6212 (N_6212,N_3922,N_3790);
or U6213 (N_6213,N_3862,N_3787);
nand U6214 (N_6214,N_4110,N_3809);
xor U6215 (N_6215,N_4880,N_4481);
nor U6216 (N_6216,N_4207,N_3954);
nand U6217 (N_6217,N_4438,N_4519);
or U6218 (N_6218,N_4349,N_4209);
xnor U6219 (N_6219,N_3992,N_4065);
xor U6220 (N_6220,N_4292,N_4543);
nand U6221 (N_6221,N_4966,N_4106);
xnor U6222 (N_6222,N_4315,N_4781);
xnor U6223 (N_6223,N_4252,N_3976);
or U6224 (N_6224,N_3788,N_4432);
xnor U6225 (N_6225,N_4388,N_3941);
nor U6226 (N_6226,N_4605,N_4343);
nor U6227 (N_6227,N_4223,N_3773);
or U6228 (N_6228,N_3929,N_4034);
and U6229 (N_6229,N_4237,N_4319);
xor U6230 (N_6230,N_4142,N_4507);
nor U6231 (N_6231,N_4972,N_4177);
or U6232 (N_6232,N_3969,N_4606);
nor U6233 (N_6233,N_3833,N_4424);
xnor U6234 (N_6234,N_4770,N_4321);
and U6235 (N_6235,N_3852,N_4925);
or U6236 (N_6236,N_4792,N_4347);
xnor U6237 (N_6237,N_4367,N_4744);
nor U6238 (N_6238,N_3826,N_4286);
and U6239 (N_6239,N_4425,N_3895);
nand U6240 (N_6240,N_4363,N_4423);
and U6241 (N_6241,N_4247,N_4619);
nor U6242 (N_6242,N_4658,N_4295);
nand U6243 (N_6243,N_3824,N_4954);
xor U6244 (N_6244,N_4320,N_4003);
xor U6245 (N_6245,N_3961,N_4819);
and U6246 (N_6246,N_4922,N_3927);
or U6247 (N_6247,N_4608,N_4619);
xnor U6248 (N_6248,N_4901,N_4030);
and U6249 (N_6249,N_4475,N_4911);
xnor U6250 (N_6250,N_5492,N_5682);
nor U6251 (N_6251,N_6103,N_5918);
nor U6252 (N_6252,N_5327,N_5425);
nand U6253 (N_6253,N_6139,N_5174);
and U6254 (N_6254,N_5664,N_5796);
or U6255 (N_6255,N_5116,N_5762);
nor U6256 (N_6256,N_5900,N_6047);
nand U6257 (N_6257,N_5381,N_6072);
and U6258 (N_6258,N_5952,N_6125);
and U6259 (N_6259,N_5244,N_5496);
nor U6260 (N_6260,N_5449,N_6163);
nor U6261 (N_6261,N_6017,N_5643);
nand U6262 (N_6262,N_5712,N_6028);
or U6263 (N_6263,N_6208,N_5936);
xor U6264 (N_6264,N_5033,N_6025);
nor U6265 (N_6265,N_5115,N_5316);
or U6266 (N_6266,N_6045,N_5532);
nor U6267 (N_6267,N_5774,N_5331);
nand U6268 (N_6268,N_5319,N_5976);
or U6269 (N_6269,N_6184,N_5265);
nand U6270 (N_6270,N_5259,N_5382);
or U6271 (N_6271,N_6115,N_5890);
nor U6272 (N_6272,N_5246,N_5704);
xnor U6273 (N_6273,N_5043,N_5340);
nor U6274 (N_6274,N_5117,N_5406);
and U6275 (N_6275,N_5751,N_5011);
and U6276 (N_6276,N_5547,N_5802);
nor U6277 (N_6277,N_5764,N_5019);
or U6278 (N_6278,N_6153,N_5880);
xor U6279 (N_6279,N_5094,N_5872);
nor U6280 (N_6280,N_5708,N_5882);
and U6281 (N_6281,N_5861,N_5143);
and U6282 (N_6282,N_6176,N_5077);
or U6283 (N_6283,N_5065,N_5909);
xor U6284 (N_6284,N_5201,N_5662);
or U6285 (N_6285,N_5630,N_5670);
or U6286 (N_6286,N_5658,N_5087);
nor U6287 (N_6287,N_5038,N_5864);
xor U6288 (N_6288,N_6190,N_5508);
or U6289 (N_6289,N_5167,N_5690);
or U6290 (N_6290,N_5758,N_5828);
nand U6291 (N_6291,N_5550,N_6071);
xnor U6292 (N_6292,N_5119,N_5454);
nand U6293 (N_6293,N_5266,N_6030);
and U6294 (N_6294,N_5911,N_5821);
xor U6295 (N_6295,N_5570,N_5130);
nand U6296 (N_6296,N_5634,N_5059);
xnor U6297 (N_6297,N_5018,N_5405);
and U6298 (N_6298,N_6170,N_5223);
or U6299 (N_6299,N_5079,N_6203);
or U6300 (N_6300,N_5848,N_5754);
and U6301 (N_6301,N_5495,N_5151);
and U6302 (N_6302,N_5233,N_5515);
xnor U6303 (N_6303,N_5363,N_6104);
or U6304 (N_6304,N_5009,N_5476);
nand U6305 (N_6305,N_5637,N_5017);
or U6306 (N_6306,N_5551,N_5456);
xor U6307 (N_6307,N_6085,N_5584);
xor U6308 (N_6308,N_6124,N_5855);
nor U6309 (N_6309,N_5687,N_5535);
nor U6310 (N_6310,N_6228,N_6201);
or U6311 (N_6311,N_5368,N_5204);
nor U6312 (N_6312,N_5322,N_5342);
and U6313 (N_6313,N_5410,N_5317);
and U6314 (N_6314,N_5049,N_5125);
nand U6315 (N_6315,N_5445,N_5501);
nor U6316 (N_6316,N_5280,N_5830);
and U6317 (N_6317,N_5301,N_5149);
nor U6318 (N_6318,N_6173,N_5845);
nor U6319 (N_6319,N_5040,N_5105);
nand U6320 (N_6320,N_5088,N_5507);
and U6321 (N_6321,N_6080,N_5652);
or U6322 (N_6322,N_6137,N_5219);
nor U6323 (N_6323,N_6038,N_5946);
nand U6324 (N_6324,N_5085,N_5228);
nor U6325 (N_6325,N_5984,N_5838);
nand U6326 (N_6326,N_5186,N_5112);
or U6327 (N_6327,N_5135,N_5992);
or U6328 (N_6328,N_5594,N_5734);
and U6329 (N_6329,N_5513,N_6185);
or U6330 (N_6330,N_5541,N_5055);
nor U6331 (N_6331,N_5620,N_5489);
nand U6332 (N_6332,N_5858,N_5494);
nand U6333 (N_6333,N_5983,N_5253);
nand U6334 (N_6334,N_5595,N_5249);
xnor U6335 (N_6335,N_6175,N_6008);
nor U6336 (N_6336,N_5942,N_5974);
or U6337 (N_6337,N_6181,N_5024);
nand U6338 (N_6338,N_5727,N_6174);
nand U6339 (N_6339,N_6101,N_6231);
xor U6340 (N_6340,N_6151,N_5225);
nand U6341 (N_6341,N_5856,N_5332);
or U6342 (N_6342,N_5181,N_5526);
nand U6343 (N_6343,N_5578,N_5711);
nand U6344 (N_6344,N_6059,N_5958);
nand U6345 (N_6345,N_6234,N_5299);
nor U6346 (N_6346,N_5698,N_6096);
xnor U6347 (N_6347,N_5592,N_5147);
xor U6348 (N_6348,N_5192,N_5298);
or U6349 (N_6349,N_5443,N_5433);
or U6350 (N_6350,N_6143,N_6225);
nor U6351 (N_6351,N_5282,N_5795);
nor U6352 (N_6352,N_5971,N_5837);
nor U6353 (N_6353,N_5060,N_6084);
xnor U6354 (N_6354,N_5925,N_5527);
nand U6355 (N_6355,N_5530,N_5409);
and U6356 (N_6356,N_5831,N_6034);
or U6357 (N_6357,N_5385,N_5020);
nor U6358 (N_6358,N_6044,N_6009);
xnor U6359 (N_6359,N_5173,N_5671);
and U6360 (N_6360,N_5525,N_6131);
and U6361 (N_6361,N_5258,N_5203);
xnor U6362 (N_6362,N_6140,N_6116);
xnor U6363 (N_6363,N_6235,N_5440);
nand U6364 (N_6364,N_5980,N_5270);
nand U6365 (N_6365,N_6001,N_5341);
nand U6366 (N_6366,N_5371,N_5310);
xnor U6367 (N_6367,N_6196,N_5654);
or U6368 (N_6368,N_5328,N_5345);
nor U6369 (N_6369,N_5887,N_6007);
nor U6370 (N_6370,N_5600,N_5252);
xor U6371 (N_6371,N_5091,N_5180);
nor U6372 (N_6372,N_5144,N_5164);
xor U6373 (N_6373,N_5553,N_5314);
xnor U6374 (N_6374,N_5365,N_5354);
or U6375 (N_6375,N_5063,N_5779);
or U6376 (N_6376,N_5997,N_5857);
and U6377 (N_6377,N_6110,N_5834);
nor U6378 (N_6378,N_5030,N_5048);
and U6379 (N_6379,N_5387,N_6249);
xnor U6380 (N_6380,N_6241,N_6068);
nand U6381 (N_6381,N_5086,N_5372);
nor U6382 (N_6382,N_6215,N_5081);
and U6383 (N_6383,N_5036,N_5102);
nand U6384 (N_6384,N_5874,N_5480);
and U6385 (N_6385,N_5408,N_5562);
and U6386 (N_6386,N_5563,N_6069);
xor U6387 (N_6387,N_6109,N_5719);
nand U6388 (N_6388,N_5614,N_6063);
and U6389 (N_6389,N_5694,N_5726);
and U6390 (N_6390,N_5128,N_5881);
and U6391 (N_6391,N_6018,N_5155);
xnor U6392 (N_6392,N_5208,N_5840);
nor U6393 (N_6393,N_5424,N_5082);
nor U6394 (N_6394,N_5669,N_5475);
xnor U6395 (N_6395,N_5278,N_6057);
nand U6396 (N_6396,N_5069,N_5871);
nand U6397 (N_6397,N_5300,N_5050);
nand U6398 (N_6398,N_6172,N_5302);
xor U6399 (N_6399,N_6200,N_6145);
or U6400 (N_6400,N_5574,N_5429);
nand U6401 (N_6401,N_5366,N_5137);
nand U6402 (N_6402,N_5885,N_6083);
and U6403 (N_6403,N_5545,N_5618);
xnor U6404 (N_6404,N_5879,N_5027);
xor U6405 (N_6405,N_5095,N_5817);
nand U6406 (N_6406,N_6219,N_5742);
xnor U6407 (N_6407,N_5703,N_5185);
xor U6408 (N_6408,N_5771,N_5292);
and U6409 (N_6409,N_5827,N_5623);
xor U6410 (N_6410,N_5142,N_5567);
xnor U6411 (N_6411,N_5188,N_6169);
and U6412 (N_6412,N_5474,N_6119);
or U6413 (N_6413,N_5775,N_5680);
nand U6414 (N_6414,N_5798,N_5770);
nor U6415 (N_6415,N_5394,N_5619);
nor U6416 (N_6416,N_5261,N_5622);
nand U6417 (N_6417,N_5296,N_5906);
nand U6418 (N_6418,N_5800,N_5807);
or U6419 (N_6419,N_5902,N_5511);
nand U6420 (N_6420,N_6081,N_5895);
or U6421 (N_6421,N_5737,N_5447);
and U6422 (N_6422,N_5362,N_5961);
and U6423 (N_6423,N_5931,N_5899);
nand U6424 (N_6424,N_5459,N_5355);
or U6425 (N_6425,N_5688,N_5254);
or U6426 (N_6426,N_6207,N_5833);
xor U6427 (N_6427,N_5490,N_5287);
xor U6428 (N_6428,N_5913,N_5210);
xnor U6429 (N_6429,N_6062,N_5989);
nor U6430 (N_6430,N_6093,N_5152);
and U6431 (N_6431,N_6221,N_5616);
xnor U6432 (N_6432,N_5315,N_5546);
and U6433 (N_6433,N_5604,N_5291);
xor U6434 (N_6434,N_5968,N_5179);
nand U6435 (N_6435,N_5632,N_5788);
xor U6436 (N_6436,N_6065,N_5401);
and U6437 (N_6437,N_5497,N_5755);
or U6438 (N_6438,N_5250,N_5555);
nand U6439 (N_6439,N_5528,N_6230);
and U6440 (N_6440,N_5006,N_5506);
nor U6441 (N_6441,N_5177,N_5548);
or U6442 (N_6442,N_5072,N_5538);
or U6443 (N_6443,N_5639,N_5446);
xor U6444 (N_6444,N_5139,N_5353);
and U6445 (N_6445,N_6024,N_5064);
and U6446 (N_6446,N_5740,N_5076);
or U6447 (N_6447,N_5303,N_5212);
nand U6448 (N_6448,N_6117,N_5450);
or U6449 (N_6449,N_5182,N_5403);
or U6450 (N_6450,N_5767,N_5191);
xnor U6451 (N_6451,N_6205,N_6199);
or U6452 (N_6452,N_6162,N_6011);
xor U6453 (N_6453,N_5383,N_6227);
and U6454 (N_6454,N_6014,N_5598);
nor U6455 (N_6455,N_5399,N_6058);
xor U6456 (N_6456,N_5170,N_5487);
xor U6457 (N_6457,N_6161,N_5517);
xnor U6458 (N_6458,N_5927,N_5759);
nor U6459 (N_6459,N_5686,N_5556);
or U6460 (N_6460,N_5376,N_5916);
and U6461 (N_6461,N_6089,N_5904);
xnor U6462 (N_6462,N_5901,N_5321);
and U6463 (N_6463,N_5364,N_5631);
and U6464 (N_6464,N_5972,N_5026);
and U6465 (N_6465,N_6029,N_5089);
xnor U6466 (N_6466,N_5812,N_6122);
nand U6467 (N_6467,N_6245,N_5001);
and U6468 (N_6468,N_6154,N_5732);
xor U6469 (N_6469,N_5947,N_5540);
nand U6470 (N_6470,N_5172,N_5935);
xnor U6471 (N_6471,N_5747,N_5836);
or U6472 (N_6472,N_5780,N_5733);
xnor U6473 (N_6473,N_5668,N_6005);
and U6474 (N_6474,N_5277,N_6088);
nor U6475 (N_6475,N_5999,N_5393);
or U6476 (N_6476,N_5470,N_5217);
nor U6477 (N_6477,N_5735,N_5978);
xnor U6478 (N_6478,N_6078,N_5558);
and U6479 (N_6479,N_5294,N_5176);
and U6480 (N_6480,N_6092,N_6033);
or U6481 (N_6481,N_5835,N_5973);
nand U6482 (N_6482,N_5295,N_5745);
xnor U6483 (N_6483,N_5851,N_5199);
xnor U6484 (N_6484,N_5564,N_5080);
nor U6485 (N_6485,N_5436,N_5552);
xnor U6486 (N_6486,N_5400,N_5998);
nand U6487 (N_6487,N_5245,N_5937);
and U6488 (N_6488,N_6127,N_5922);
xnor U6489 (N_6489,N_5760,N_5549);
nand U6490 (N_6490,N_5723,N_5260);
nand U6491 (N_6491,N_6134,N_5344);
nor U6492 (N_6492,N_6167,N_6098);
xnor U6493 (N_6493,N_6086,N_6168);
nor U6494 (N_6494,N_5533,N_5876);
xnor U6495 (N_6495,N_5412,N_5070);
nor U6496 (N_6496,N_5183,N_5361);
xor U6497 (N_6497,N_5166,N_5500);
or U6498 (N_6498,N_6158,N_5272);
and U6499 (N_6499,N_5090,N_5028);
xor U6500 (N_6500,N_5934,N_5569);
xor U6501 (N_6501,N_5285,N_5150);
nand U6502 (N_6502,N_5516,N_5964);
nand U6503 (N_6503,N_5386,N_6177);
xnor U6504 (N_6504,N_6111,N_5805);
or U6505 (N_6505,N_5903,N_5101);
nand U6506 (N_6506,N_5471,N_5785);
xor U6507 (N_6507,N_5843,N_5842);
or U6508 (N_6508,N_5438,N_6118);
nand U6509 (N_6509,N_5061,N_5455);
and U6510 (N_6510,N_6229,N_5263);
or U6511 (N_6511,N_6152,N_5502);
nor U6512 (N_6512,N_6186,N_5121);
nand U6513 (N_6513,N_5232,N_5162);
nor U6514 (N_6514,N_5012,N_6197);
or U6515 (N_6515,N_5777,N_5700);
xnor U6516 (N_6516,N_6052,N_5572);
nor U6517 (N_6517,N_5458,N_5666);
nand U6518 (N_6518,N_5790,N_5912);
xor U6519 (N_6519,N_5580,N_5271);
and U6520 (N_6520,N_6073,N_5693);
nand U6521 (N_6521,N_6036,N_5859);
and U6522 (N_6522,N_5384,N_5200);
nor U6523 (N_6523,N_6132,N_6076);
xor U6524 (N_6524,N_5052,N_5773);
or U6525 (N_6525,N_5655,N_5514);
nand U6526 (N_6526,N_5896,N_5350);
or U6527 (N_6527,N_6240,N_5753);
and U6528 (N_6528,N_6183,N_5276);
nand U6529 (N_6529,N_5957,N_5993);
nor U6530 (N_6530,N_6182,N_5606);
xor U6531 (N_6531,N_5356,N_5612);
and U6532 (N_6532,N_5377,N_5929);
or U6533 (N_6533,N_5312,N_5111);
or U6534 (N_6534,N_5073,N_5437);
nor U6535 (N_6535,N_5160,N_5389);
or U6536 (N_6536,N_5829,N_5242);
xnor U6537 (N_6537,N_5894,N_5194);
nor U6538 (N_6538,N_6238,N_6106);
or U6539 (N_6539,N_5818,N_6180);
nand U6540 (N_6540,N_5588,N_6070);
nand U6541 (N_6541,N_5923,N_6149);
or U6542 (N_6542,N_5846,N_5793);
nor U6543 (N_6543,N_5994,N_5256);
nand U6544 (N_6544,N_6136,N_5120);
xnor U6545 (N_6545,N_6043,N_5791);
xor U6546 (N_6546,N_5421,N_5118);
nand U6547 (N_6547,N_5815,N_5165);
or U6548 (N_6548,N_5205,N_5251);
nand U6549 (N_6549,N_5640,N_5692);
and U6550 (N_6550,N_5839,N_6141);
or U6551 (N_6551,N_5635,N_5097);
nand U6552 (N_6552,N_5472,N_6242);
xnor U6553 (N_6553,N_5482,N_5518);
nand U6554 (N_6554,N_5877,N_5907);
and U6555 (N_6555,N_5675,N_5596);
and U6556 (N_6556,N_5230,N_5949);
or U6557 (N_6557,N_5724,N_6067);
or U6558 (N_6558,N_5649,N_5531);
and U6559 (N_6559,N_5878,N_6102);
nor U6560 (N_6560,N_5921,N_5792);
nor U6561 (N_6561,N_6004,N_5672);
and U6562 (N_6562,N_5696,N_5781);
nor U6563 (N_6563,N_5352,N_5367);
nor U6564 (N_6564,N_5731,N_5710);
xor U6565 (N_6565,N_5196,N_6042);
nand U6566 (N_6566,N_5801,N_5042);
nand U6567 (N_6567,N_5676,N_5359);
and U6568 (N_6568,N_6056,N_5369);
nor U6569 (N_6569,N_5650,N_5163);
and U6570 (N_6570,N_6120,N_5797);
nor U6571 (N_6571,N_5722,N_5305);
nor U6572 (N_6572,N_5542,N_6015);
nor U6573 (N_6573,N_5597,N_5289);
or U6574 (N_6574,N_5811,N_6010);
and U6575 (N_6575,N_5267,N_5853);
nand U6576 (N_6576,N_5211,N_6246);
nand U6577 (N_6577,N_5068,N_5624);
xor U6578 (N_6578,N_5782,N_5602);
or U6579 (N_6579,N_5349,N_6051);
xnor U6580 (N_6580,N_5248,N_5813);
nand U6581 (N_6581,N_5615,N_5195);
nand U6582 (N_6582,N_6144,N_5083);
and U6583 (N_6583,N_5728,N_6178);
nand U6584 (N_6584,N_5794,N_5343);
nand U6585 (N_6585,N_5279,N_5307);
nand U6586 (N_6586,N_5736,N_5216);
xnor U6587 (N_6587,N_5746,N_5577);
and U6588 (N_6588,N_5391,N_5062);
and U6589 (N_6589,N_6129,N_5098);
nand U6590 (N_6590,N_6138,N_5110);
or U6591 (N_6591,N_5663,N_5706);
and U6592 (N_6592,N_5816,N_5697);
nand U6593 (N_6593,N_5713,N_5138);
nor U6594 (N_6594,N_5720,N_5948);
xnor U6595 (N_6595,N_5178,N_5132);
and U6596 (N_6596,N_5629,N_5730);
or U6597 (N_6597,N_5886,N_6217);
xor U6598 (N_6598,N_5933,N_5575);
or U6599 (N_6599,N_5648,N_5241);
nor U6600 (N_6600,N_5108,N_6090);
xor U6601 (N_6601,N_5107,N_5987);
and U6602 (N_6602,N_5411,N_6105);
nand U6603 (N_6603,N_5329,N_5021);
or U6604 (N_6604,N_5323,N_5257);
xor U6605 (N_6605,N_6160,N_5220);
nor U6606 (N_6606,N_6236,N_5491);
nand U6607 (N_6607,N_5415,N_5426);
xor U6608 (N_6608,N_5725,N_5557);
nand U6609 (N_6609,N_5114,N_6128);
nand U6610 (N_6610,N_5854,N_5863);
or U6611 (N_6611,N_5761,N_5678);
or U6612 (N_6612,N_5333,N_5778);
xnor U6613 (N_6613,N_5991,N_6216);
nor U6614 (N_6614,N_5847,N_6099);
nand U6615 (N_6615,N_5227,N_5419);
or U6616 (N_6616,N_5032,N_5351);
or U6617 (N_6617,N_5045,N_5529);
nor U6618 (N_6618,N_5825,N_5641);
and U6619 (N_6619,N_6218,N_5380);
nor U6620 (N_6620,N_5238,N_5716);
nand U6621 (N_6621,N_5892,N_6107);
and U6622 (N_6622,N_5136,N_5207);
or U6623 (N_6623,N_5875,N_5047);
xnor U6624 (N_6624,N_5397,N_5920);
nor U6625 (N_6625,N_5092,N_6050);
or U6626 (N_6626,N_5625,N_5520);
nand U6627 (N_6627,N_5283,N_5402);
xor U6628 (N_6628,N_5168,N_5681);
nand U6629 (N_6629,N_5420,N_5945);
and U6630 (N_6630,N_5414,N_5309);
and U6631 (N_6631,N_5591,N_6202);
and U6632 (N_6632,N_5585,N_5275);
xor U6633 (N_6633,N_5647,N_5699);
nor U6634 (N_6634,N_6039,N_6130);
xnor U6635 (N_6635,N_5274,N_5084);
or U6636 (N_6636,N_6082,N_5930);
and U6637 (N_6637,N_5659,N_5928);
nor U6638 (N_6638,N_5269,N_5589);
nand U6639 (N_6639,N_5129,N_6055);
and U6640 (N_6640,N_5483,N_5103);
and U6641 (N_6641,N_5417,N_5627);
xor U6642 (N_6642,N_5870,N_5560);
nand U6643 (N_6643,N_5691,N_5378);
nand U6644 (N_6644,N_5660,N_5473);
or U6645 (N_6645,N_6147,N_6209);
and U6646 (N_6646,N_5434,N_5910);
or U6647 (N_6647,N_5729,N_5236);
and U6648 (N_6648,N_5003,N_5963);
and U6649 (N_6649,N_5932,N_5441);
nor U6650 (N_6650,N_5867,N_5665);
nand U6651 (N_6651,N_6000,N_5981);
nand U6652 (N_6652,N_5008,N_5214);
nor U6653 (N_6653,N_5034,N_6233);
xor U6654 (N_6654,N_6123,N_5464);
xnor U6655 (N_6655,N_5237,N_5750);
nor U6656 (N_6656,N_5002,N_5536);
nor U6657 (N_6657,N_5783,N_5146);
or U6658 (N_6658,N_6243,N_5452);
or U6659 (N_6659,N_5919,N_5888);
xnor U6660 (N_6660,N_5617,N_5074);
nor U6661 (N_6661,N_6188,N_6021);
or U6662 (N_6662,N_5071,N_5486);
nor U6663 (N_6663,N_5453,N_5960);
and U6664 (N_6664,N_5803,N_5235);
or U6665 (N_6665,N_5939,N_6060);
nand U6666 (N_6666,N_6046,N_5705);
xnor U6667 (N_6667,N_6156,N_5581);
or U6668 (N_6668,N_5673,N_5738);
nand U6669 (N_6669,N_5375,N_5416);
nand U6670 (N_6670,N_5126,N_5926);
and U6671 (N_6671,N_5145,N_6198);
nand U6672 (N_6672,N_6019,N_5601);
and U6673 (N_6673,N_6210,N_6206);
nor U6674 (N_6674,N_5427,N_5171);
nand U6675 (N_6675,N_6006,N_6112);
xor U6676 (N_6676,N_5524,N_6239);
nand U6677 (N_6677,N_5335,N_5099);
nor U6678 (N_6678,N_5962,N_5626);
nor U6679 (N_6679,N_5784,N_5313);
and U6680 (N_6680,N_5039,N_5396);
nor U6681 (N_6681,N_5066,N_5175);
nand U6682 (N_6682,N_5852,N_6003);
and U6683 (N_6683,N_6022,N_5809);
nor U6684 (N_6684,N_5884,N_5897);
nor U6685 (N_6685,N_5757,N_5293);
and U6686 (N_6686,N_6204,N_6066);
and U6687 (N_6687,N_5789,N_5255);
and U6688 (N_6688,N_5224,N_5543);
xor U6689 (N_6689,N_5122,N_5599);
xor U6690 (N_6690,N_5005,N_5418);
and U6691 (N_6691,N_5124,N_5338);
and U6692 (N_6692,N_5306,N_5374);
nor U6693 (N_6693,N_5769,N_5579);
nand U6694 (N_6694,N_6027,N_5463);
xnor U6695 (N_6695,N_5810,N_5290);
nand U6696 (N_6696,N_6095,N_5457);
nand U6697 (N_6697,N_6074,N_5133);
and U6698 (N_6698,N_5264,N_6026);
nand U6699 (N_6699,N_6054,N_5869);
nand U6700 (N_6700,N_6037,N_6135);
xor U6701 (N_6701,N_5297,N_5586);
nor U6702 (N_6702,N_5683,N_5407);
and U6703 (N_6703,N_5046,N_5158);
and U6704 (N_6704,N_5814,N_5127);
nor U6705 (N_6705,N_5140,N_5106);
nand U6706 (N_6706,N_6053,N_5209);
nand U6707 (N_6707,N_5914,N_5908);
and U6708 (N_6708,N_5787,N_5539);
xnor U6709 (N_6709,N_5841,N_5218);
and U6710 (N_6710,N_5583,N_5898);
and U6711 (N_6711,N_5392,N_6226);
nor U6712 (N_6712,N_5741,N_5849);
xnor U6713 (N_6713,N_5054,N_5202);
or U6714 (N_6714,N_6126,N_5093);
or U6715 (N_6715,N_5187,N_5284);
nor U6716 (N_6716,N_6114,N_6150);
nor U6717 (N_6717,N_5941,N_5702);
or U6718 (N_6718,N_6087,N_5100);
nor U6719 (N_6719,N_6049,N_5982);
and U6720 (N_6720,N_5422,N_5056);
or U6721 (N_6721,N_5684,N_6214);
xnor U6722 (N_6722,N_5943,N_5893);
xor U6723 (N_6723,N_5123,N_5288);
nor U6724 (N_6724,N_5320,N_5304);
and U6725 (N_6725,N_5488,N_5721);
or U6726 (N_6726,N_6075,N_6023);
and U6727 (N_6727,N_5965,N_5559);
or U6728 (N_6728,N_5053,N_5905);
xnor U6729 (N_6729,N_5197,N_5823);
xor U6730 (N_6730,N_5953,N_5763);
and U6731 (N_6731,N_5339,N_5051);
and U6732 (N_6732,N_5281,N_5657);
and U6733 (N_6733,N_6002,N_5959);
nor U6734 (N_6734,N_5537,N_5695);
xor U6735 (N_6735,N_5431,N_6146);
and U6736 (N_6736,N_5234,N_5661);
xnor U6737 (N_6737,N_5766,N_5714);
xnor U6738 (N_6738,N_5607,N_5022);
or U6739 (N_6739,N_5370,N_5873);
xor U6740 (N_6740,N_5621,N_5915);
nor U6741 (N_6741,N_5995,N_6165);
nand U6742 (N_6742,N_5247,N_5357);
xor U6743 (N_6743,N_5576,N_5156);
or U6744 (N_6744,N_5786,N_6191);
nor U6745 (N_6745,N_5478,N_5967);
xnor U6746 (N_6746,N_5058,N_6244);
and U6747 (N_6747,N_5398,N_5970);
or U6748 (N_6748,N_5239,N_5715);
xor U6749 (N_6749,N_5776,N_5467);
xnor U6750 (N_6750,N_5819,N_5308);
nor U6751 (N_6751,N_5566,N_5031);
or U6752 (N_6752,N_5193,N_5677);
xnor U6753 (N_6753,N_5756,N_6020);
nor U6754 (N_6754,N_5709,N_5346);
nand U6755 (N_6755,N_5990,N_5035);
xor U6756 (N_6756,N_5609,N_5844);
nor U6757 (N_6757,N_6171,N_5969);
xnor U6758 (N_6758,N_5439,N_5744);
or U6759 (N_6759,N_5862,N_6213);
nand U6760 (N_6760,N_5868,N_5347);
xnor U6761 (N_6761,N_5651,N_5889);
and U6762 (N_6762,N_6061,N_5940);
nand U6763 (N_6763,N_5190,N_6016);
and U6764 (N_6764,N_6192,N_5373);
nor U6765 (N_6765,N_5498,N_6142);
or U6766 (N_6766,N_5286,N_5154);
nand U6767 (N_6767,N_5222,N_5324);
or U6768 (N_6768,N_5311,N_5044);
xnor U6769 (N_6769,N_5979,N_5950);
xor U6770 (N_6770,N_5161,N_6193);
nor U6771 (N_6771,N_5571,N_5603);
and U6772 (N_6772,N_5544,N_5718);
xnor U6773 (N_6773,N_5423,N_5004);
nor U6774 (N_6774,N_5485,N_5468);
xnor U6775 (N_6775,N_5273,N_5243);
nor U6776 (N_6776,N_5985,N_5390);
or U6777 (N_6777,N_5522,N_5226);
and U6778 (N_6778,N_5808,N_5206);
nor U6779 (N_6779,N_5534,N_6211);
or U6780 (N_6780,N_5826,N_5975);
xnor U6781 (N_6781,N_5772,N_5016);
and U6782 (N_6782,N_5334,N_5505);
or U6783 (N_6783,N_5554,N_5956);
xor U6784 (N_6784,N_5954,N_5689);
or U6785 (N_6785,N_5231,N_5109);
xor U6786 (N_6786,N_5013,N_5015);
nand U6787 (N_6787,N_5509,N_5850);
xor U6788 (N_6788,N_5213,N_6100);
nand U6789 (N_6789,N_5240,N_5938);
xor U6790 (N_6790,N_5318,N_5799);
and U6791 (N_6791,N_5413,N_5404);
or U6792 (N_6792,N_5451,N_5014);
nand U6793 (N_6793,N_6237,N_5573);
or U6794 (N_6794,N_6108,N_6187);
xor U6795 (N_6795,N_5866,N_5430);
nor U6796 (N_6796,N_5996,N_6157);
and U6797 (N_6797,N_5891,N_5337);
or U6798 (N_6798,N_5113,N_6220);
xnor U6799 (N_6799,N_5477,N_5484);
nor U6800 (N_6800,N_6064,N_5917);
or U6801 (N_6801,N_5804,N_6248);
or U6802 (N_6802,N_5986,N_5153);
nand U6803 (N_6803,N_5743,N_5628);
or U6804 (N_6804,N_5519,N_5348);
nand U6805 (N_6805,N_5096,N_5025);
xor U6806 (N_6806,N_6224,N_6032);
and U6807 (N_6807,N_5007,N_5966);
xnor U6808 (N_6808,N_6194,N_5636);
xnor U6809 (N_6809,N_5388,N_5752);
nor U6810 (N_6810,N_5717,N_6148);
nor U6811 (N_6811,N_5748,N_5221);
nor U6812 (N_6812,N_5325,N_5860);
xnor U6813 (N_6813,N_6094,N_5360);
nand U6814 (N_6814,N_6048,N_5448);
nand U6815 (N_6815,N_6212,N_5481);
nand U6816 (N_6816,N_6164,N_5590);
or U6817 (N_6817,N_5642,N_5512);
nand U6818 (N_6818,N_5262,N_5587);
nor U6819 (N_6819,N_5432,N_5646);
or U6820 (N_6820,N_5685,N_5593);
nor U6821 (N_6821,N_5510,N_6031);
nand U6822 (N_6822,N_5215,N_5565);
xnor U6823 (N_6823,N_5977,N_5067);
xnor U6824 (N_6824,N_5159,N_5674);
xor U6825 (N_6825,N_5608,N_5479);
nor U6826 (N_6826,N_5395,N_5820);
and U6827 (N_6827,N_5988,N_5057);
and U6828 (N_6828,N_5883,N_5739);
nand U6829 (N_6829,N_6159,N_5503);
xor U6830 (N_6830,N_5466,N_5148);
and U6831 (N_6831,N_6035,N_5131);
and U6832 (N_6832,N_5358,N_5610);
nor U6833 (N_6833,N_5667,N_5461);
and U6834 (N_6834,N_5078,N_5169);
and U6835 (N_6835,N_6121,N_5460);
nand U6836 (N_6836,N_6155,N_5336);
and U6837 (N_6837,N_5499,N_5465);
nand U6838 (N_6838,N_5444,N_5442);
and U6839 (N_6839,N_5023,N_6189);
nand U6840 (N_6840,N_6091,N_5822);
nor U6841 (N_6841,N_5944,N_5644);
and U6842 (N_6842,N_5000,N_5104);
nand U6843 (N_6843,N_6012,N_5582);
nand U6844 (N_6844,N_5633,N_5645);
or U6845 (N_6845,N_5189,N_5504);
nand U6846 (N_6846,N_6113,N_5010);
or U6847 (N_6847,N_5611,N_5824);
nand U6848 (N_6848,N_5832,N_5521);
and U6849 (N_6849,N_5605,N_5326);
nor U6850 (N_6850,N_5701,N_6179);
or U6851 (N_6851,N_5268,N_6013);
nand U6852 (N_6852,N_5924,N_6041);
nand U6853 (N_6853,N_5428,N_6077);
nor U6854 (N_6854,N_5653,N_6247);
or U6855 (N_6855,N_5379,N_5765);
or U6856 (N_6856,N_6223,N_6097);
or U6857 (N_6857,N_5037,N_5462);
xor U6858 (N_6858,N_5561,N_5435);
xor U6859 (N_6859,N_6166,N_5638);
xnor U6860 (N_6860,N_6133,N_5029);
xor U6861 (N_6861,N_5951,N_5749);
nor U6862 (N_6862,N_5141,N_5469);
nor U6863 (N_6863,N_5656,N_5041);
and U6864 (N_6864,N_5229,N_5955);
xnor U6865 (N_6865,N_5198,N_5330);
nand U6866 (N_6866,N_5707,N_5134);
nor U6867 (N_6867,N_5157,N_5523);
nor U6868 (N_6868,N_5865,N_6222);
and U6869 (N_6869,N_5613,N_5679);
and U6870 (N_6870,N_6079,N_6040);
xnor U6871 (N_6871,N_5075,N_5768);
or U6872 (N_6872,N_6232,N_5184);
nand U6873 (N_6873,N_6195,N_5568);
nand U6874 (N_6874,N_5493,N_5806);
nand U6875 (N_6875,N_5789,N_5612);
or U6876 (N_6876,N_6161,N_5676);
xor U6877 (N_6877,N_5148,N_5844);
nand U6878 (N_6878,N_5986,N_5778);
nor U6879 (N_6879,N_5687,N_6068);
nor U6880 (N_6880,N_6117,N_5779);
nand U6881 (N_6881,N_5213,N_5709);
xnor U6882 (N_6882,N_5666,N_5064);
or U6883 (N_6883,N_5136,N_5655);
or U6884 (N_6884,N_5881,N_5822);
or U6885 (N_6885,N_6040,N_5819);
nand U6886 (N_6886,N_5708,N_5860);
nand U6887 (N_6887,N_5535,N_5807);
nor U6888 (N_6888,N_5640,N_5957);
xor U6889 (N_6889,N_6101,N_6039);
or U6890 (N_6890,N_5790,N_5991);
or U6891 (N_6891,N_5977,N_5247);
and U6892 (N_6892,N_5335,N_6132);
nand U6893 (N_6893,N_5987,N_5622);
xnor U6894 (N_6894,N_5708,N_5346);
and U6895 (N_6895,N_5767,N_5218);
nand U6896 (N_6896,N_5453,N_5016);
xor U6897 (N_6897,N_5422,N_5232);
nand U6898 (N_6898,N_5086,N_5757);
or U6899 (N_6899,N_5371,N_5540);
nor U6900 (N_6900,N_5372,N_6183);
or U6901 (N_6901,N_5029,N_5949);
and U6902 (N_6902,N_5377,N_6067);
xor U6903 (N_6903,N_5676,N_5542);
nand U6904 (N_6904,N_6107,N_5621);
nor U6905 (N_6905,N_5987,N_5688);
and U6906 (N_6906,N_5341,N_5706);
nand U6907 (N_6907,N_5758,N_5257);
or U6908 (N_6908,N_5776,N_5308);
nor U6909 (N_6909,N_6005,N_5639);
and U6910 (N_6910,N_5849,N_6175);
nand U6911 (N_6911,N_6134,N_5629);
xor U6912 (N_6912,N_5822,N_5827);
or U6913 (N_6913,N_5888,N_5199);
and U6914 (N_6914,N_6037,N_6053);
xnor U6915 (N_6915,N_6074,N_5196);
xnor U6916 (N_6916,N_6043,N_5280);
nand U6917 (N_6917,N_5227,N_6002);
nor U6918 (N_6918,N_5492,N_5641);
nand U6919 (N_6919,N_6090,N_5165);
or U6920 (N_6920,N_5373,N_5343);
and U6921 (N_6921,N_5446,N_5889);
or U6922 (N_6922,N_5512,N_5755);
nand U6923 (N_6923,N_5639,N_6092);
nor U6924 (N_6924,N_5561,N_5405);
nor U6925 (N_6925,N_5838,N_5620);
nand U6926 (N_6926,N_5942,N_6037);
xnor U6927 (N_6927,N_5341,N_5132);
nor U6928 (N_6928,N_5192,N_5012);
xnor U6929 (N_6929,N_5009,N_5592);
and U6930 (N_6930,N_5762,N_6224);
or U6931 (N_6931,N_5541,N_5963);
nor U6932 (N_6932,N_5169,N_5489);
nand U6933 (N_6933,N_5982,N_5229);
xnor U6934 (N_6934,N_6173,N_5569);
nand U6935 (N_6935,N_5851,N_5592);
xnor U6936 (N_6936,N_5466,N_5585);
or U6937 (N_6937,N_5747,N_5310);
or U6938 (N_6938,N_6047,N_5390);
and U6939 (N_6939,N_5080,N_5408);
and U6940 (N_6940,N_5746,N_5076);
xor U6941 (N_6941,N_5370,N_5657);
or U6942 (N_6942,N_5063,N_5652);
xor U6943 (N_6943,N_6090,N_5444);
xor U6944 (N_6944,N_5381,N_5887);
or U6945 (N_6945,N_5302,N_5340);
nor U6946 (N_6946,N_6050,N_6120);
and U6947 (N_6947,N_6146,N_5342);
xnor U6948 (N_6948,N_5745,N_5820);
nor U6949 (N_6949,N_5262,N_5676);
xor U6950 (N_6950,N_5855,N_5461);
or U6951 (N_6951,N_5077,N_5022);
nand U6952 (N_6952,N_5199,N_6246);
nand U6953 (N_6953,N_5305,N_6169);
nor U6954 (N_6954,N_6208,N_5745);
and U6955 (N_6955,N_5011,N_5453);
and U6956 (N_6956,N_5256,N_6124);
or U6957 (N_6957,N_5064,N_5590);
and U6958 (N_6958,N_5513,N_5013);
nand U6959 (N_6959,N_5110,N_5055);
or U6960 (N_6960,N_5263,N_5480);
and U6961 (N_6961,N_5051,N_6186);
nand U6962 (N_6962,N_5929,N_5563);
nand U6963 (N_6963,N_5169,N_5249);
xnor U6964 (N_6964,N_5056,N_5662);
and U6965 (N_6965,N_5215,N_5639);
or U6966 (N_6966,N_5435,N_5838);
nand U6967 (N_6967,N_5468,N_5844);
xor U6968 (N_6968,N_5634,N_5621);
nand U6969 (N_6969,N_5353,N_5322);
nor U6970 (N_6970,N_5851,N_5055);
xor U6971 (N_6971,N_6061,N_5631);
xnor U6972 (N_6972,N_5673,N_5555);
nand U6973 (N_6973,N_5782,N_5506);
xnor U6974 (N_6974,N_6050,N_5558);
and U6975 (N_6975,N_5248,N_5276);
nand U6976 (N_6976,N_6070,N_6073);
and U6977 (N_6977,N_5517,N_5407);
nor U6978 (N_6978,N_6030,N_5246);
or U6979 (N_6979,N_6062,N_5592);
nand U6980 (N_6980,N_6210,N_5082);
and U6981 (N_6981,N_6196,N_5468);
nor U6982 (N_6982,N_5513,N_6171);
nor U6983 (N_6983,N_5094,N_5947);
or U6984 (N_6984,N_5392,N_5576);
nor U6985 (N_6985,N_5081,N_5249);
xnor U6986 (N_6986,N_5913,N_6184);
xor U6987 (N_6987,N_5402,N_5241);
xnor U6988 (N_6988,N_5039,N_5943);
and U6989 (N_6989,N_5425,N_5876);
nor U6990 (N_6990,N_6059,N_5146);
nor U6991 (N_6991,N_5815,N_5070);
nor U6992 (N_6992,N_5879,N_5754);
and U6993 (N_6993,N_5990,N_5067);
nand U6994 (N_6994,N_6167,N_5892);
nor U6995 (N_6995,N_6182,N_6246);
xnor U6996 (N_6996,N_5707,N_6014);
or U6997 (N_6997,N_5933,N_5295);
and U6998 (N_6998,N_5926,N_5817);
nand U6999 (N_6999,N_6056,N_5749);
nor U7000 (N_7000,N_6023,N_5158);
and U7001 (N_7001,N_5003,N_5394);
nor U7002 (N_7002,N_5076,N_5193);
and U7003 (N_7003,N_5186,N_5021);
and U7004 (N_7004,N_5505,N_5657);
or U7005 (N_7005,N_5023,N_5630);
nor U7006 (N_7006,N_5131,N_5784);
and U7007 (N_7007,N_5753,N_5709);
and U7008 (N_7008,N_5698,N_5933);
and U7009 (N_7009,N_6019,N_5215);
xor U7010 (N_7010,N_5195,N_5636);
and U7011 (N_7011,N_5188,N_5067);
and U7012 (N_7012,N_5719,N_5867);
nor U7013 (N_7013,N_5960,N_5533);
or U7014 (N_7014,N_5678,N_5566);
xnor U7015 (N_7015,N_5130,N_5328);
nor U7016 (N_7016,N_6232,N_5541);
nor U7017 (N_7017,N_5388,N_5741);
and U7018 (N_7018,N_5690,N_5445);
nand U7019 (N_7019,N_5531,N_5392);
xor U7020 (N_7020,N_5646,N_5157);
xnor U7021 (N_7021,N_6003,N_5068);
and U7022 (N_7022,N_5288,N_5902);
nand U7023 (N_7023,N_6163,N_5494);
nor U7024 (N_7024,N_5964,N_6135);
nor U7025 (N_7025,N_5778,N_6179);
nor U7026 (N_7026,N_5467,N_5128);
nor U7027 (N_7027,N_5339,N_5829);
or U7028 (N_7028,N_6200,N_5889);
nor U7029 (N_7029,N_6063,N_5196);
xor U7030 (N_7030,N_5287,N_5753);
nand U7031 (N_7031,N_5391,N_5022);
xor U7032 (N_7032,N_5098,N_5633);
and U7033 (N_7033,N_5755,N_6212);
and U7034 (N_7034,N_5363,N_6134);
and U7035 (N_7035,N_5697,N_5965);
nor U7036 (N_7036,N_5399,N_5701);
and U7037 (N_7037,N_5186,N_6033);
xor U7038 (N_7038,N_5240,N_5324);
xnor U7039 (N_7039,N_5842,N_6214);
nand U7040 (N_7040,N_5972,N_6130);
and U7041 (N_7041,N_5090,N_6041);
nand U7042 (N_7042,N_5652,N_5536);
nand U7043 (N_7043,N_5072,N_6048);
nor U7044 (N_7044,N_5794,N_5755);
nand U7045 (N_7045,N_5186,N_5680);
xnor U7046 (N_7046,N_5324,N_5867);
nor U7047 (N_7047,N_5951,N_5106);
or U7048 (N_7048,N_6094,N_5059);
xnor U7049 (N_7049,N_5846,N_5651);
or U7050 (N_7050,N_6118,N_5792);
nand U7051 (N_7051,N_5891,N_5406);
xor U7052 (N_7052,N_6187,N_5101);
nand U7053 (N_7053,N_6085,N_5720);
xor U7054 (N_7054,N_5433,N_5855);
xor U7055 (N_7055,N_5116,N_6143);
nor U7056 (N_7056,N_5315,N_5630);
nor U7057 (N_7057,N_5469,N_6188);
nand U7058 (N_7058,N_5680,N_5878);
xnor U7059 (N_7059,N_5629,N_5318);
or U7060 (N_7060,N_6160,N_5995);
nand U7061 (N_7061,N_6185,N_5844);
nand U7062 (N_7062,N_5320,N_5171);
or U7063 (N_7063,N_5724,N_5160);
and U7064 (N_7064,N_5627,N_5072);
nor U7065 (N_7065,N_5132,N_5726);
nand U7066 (N_7066,N_5992,N_5077);
xnor U7067 (N_7067,N_5390,N_5866);
and U7068 (N_7068,N_5341,N_5130);
or U7069 (N_7069,N_5340,N_5962);
xnor U7070 (N_7070,N_5680,N_5063);
and U7071 (N_7071,N_5384,N_5325);
nand U7072 (N_7072,N_6166,N_5675);
and U7073 (N_7073,N_5714,N_5291);
nand U7074 (N_7074,N_6239,N_5944);
or U7075 (N_7075,N_5145,N_5707);
xor U7076 (N_7076,N_5968,N_5884);
or U7077 (N_7077,N_5699,N_5792);
and U7078 (N_7078,N_6059,N_5503);
xnor U7079 (N_7079,N_5421,N_6190);
and U7080 (N_7080,N_6123,N_5059);
nor U7081 (N_7081,N_6231,N_5215);
xnor U7082 (N_7082,N_5433,N_5802);
or U7083 (N_7083,N_5293,N_5813);
nor U7084 (N_7084,N_5117,N_5988);
and U7085 (N_7085,N_6234,N_6175);
nor U7086 (N_7086,N_6236,N_5937);
and U7087 (N_7087,N_5852,N_5290);
or U7088 (N_7088,N_5443,N_6114);
or U7089 (N_7089,N_5818,N_5322);
or U7090 (N_7090,N_5079,N_6189);
nand U7091 (N_7091,N_5866,N_5611);
or U7092 (N_7092,N_5058,N_5417);
nand U7093 (N_7093,N_5815,N_5105);
or U7094 (N_7094,N_5956,N_5023);
xor U7095 (N_7095,N_6152,N_5680);
nor U7096 (N_7096,N_6061,N_5835);
or U7097 (N_7097,N_5947,N_5872);
nand U7098 (N_7098,N_6225,N_5037);
nor U7099 (N_7099,N_5555,N_5162);
nand U7100 (N_7100,N_6061,N_6112);
nand U7101 (N_7101,N_5788,N_5170);
and U7102 (N_7102,N_5430,N_6176);
nand U7103 (N_7103,N_6074,N_5658);
or U7104 (N_7104,N_5217,N_5777);
or U7105 (N_7105,N_5834,N_5935);
nor U7106 (N_7106,N_6220,N_6104);
and U7107 (N_7107,N_5208,N_5296);
nand U7108 (N_7108,N_5219,N_5509);
and U7109 (N_7109,N_5520,N_5079);
nand U7110 (N_7110,N_5181,N_5023);
xor U7111 (N_7111,N_5589,N_5248);
and U7112 (N_7112,N_6006,N_5797);
nor U7113 (N_7113,N_5682,N_6008);
nor U7114 (N_7114,N_5089,N_5525);
and U7115 (N_7115,N_6099,N_5258);
xnor U7116 (N_7116,N_5601,N_5254);
and U7117 (N_7117,N_5053,N_5412);
nand U7118 (N_7118,N_5091,N_5442);
xnor U7119 (N_7119,N_5208,N_6176);
xnor U7120 (N_7120,N_5504,N_6043);
nand U7121 (N_7121,N_5017,N_5467);
nand U7122 (N_7122,N_5331,N_5384);
or U7123 (N_7123,N_5458,N_6222);
or U7124 (N_7124,N_5482,N_5817);
nand U7125 (N_7125,N_5551,N_5574);
nand U7126 (N_7126,N_5995,N_6100);
or U7127 (N_7127,N_6204,N_5768);
and U7128 (N_7128,N_5488,N_5402);
xor U7129 (N_7129,N_5852,N_5663);
nand U7130 (N_7130,N_6212,N_5660);
or U7131 (N_7131,N_5291,N_6034);
nor U7132 (N_7132,N_5843,N_5939);
or U7133 (N_7133,N_5576,N_5435);
nand U7134 (N_7134,N_6132,N_5769);
xor U7135 (N_7135,N_5524,N_5770);
or U7136 (N_7136,N_5644,N_6052);
and U7137 (N_7137,N_5385,N_5781);
nand U7138 (N_7138,N_5789,N_5507);
nand U7139 (N_7139,N_5103,N_5636);
or U7140 (N_7140,N_5307,N_5705);
xnor U7141 (N_7141,N_5803,N_5370);
nand U7142 (N_7142,N_5659,N_5015);
nor U7143 (N_7143,N_6058,N_6040);
nor U7144 (N_7144,N_5295,N_5831);
and U7145 (N_7145,N_5089,N_5384);
nor U7146 (N_7146,N_6191,N_6095);
xor U7147 (N_7147,N_5038,N_5565);
nor U7148 (N_7148,N_6006,N_6053);
nor U7149 (N_7149,N_5678,N_5318);
or U7150 (N_7150,N_6038,N_6047);
or U7151 (N_7151,N_6107,N_6181);
or U7152 (N_7152,N_5324,N_5939);
and U7153 (N_7153,N_5387,N_5979);
xnor U7154 (N_7154,N_5533,N_5369);
and U7155 (N_7155,N_5764,N_6045);
and U7156 (N_7156,N_5011,N_6154);
nand U7157 (N_7157,N_5756,N_5229);
or U7158 (N_7158,N_5497,N_5230);
nor U7159 (N_7159,N_5011,N_5929);
and U7160 (N_7160,N_5384,N_6060);
xnor U7161 (N_7161,N_5692,N_5833);
nand U7162 (N_7162,N_5933,N_5009);
nand U7163 (N_7163,N_5135,N_5561);
xor U7164 (N_7164,N_5363,N_5775);
or U7165 (N_7165,N_5160,N_5005);
and U7166 (N_7166,N_5902,N_5441);
xor U7167 (N_7167,N_5688,N_5151);
nor U7168 (N_7168,N_5458,N_5362);
and U7169 (N_7169,N_5576,N_5750);
xor U7170 (N_7170,N_5012,N_5045);
and U7171 (N_7171,N_5815,N_6093);
xor U7172 (N_7172,N_5569,N_5498);
nand U7173 (N_7173,N_5294,N_5702);
and U7174 (N_7174,N_5637,N_5035);
nand U7175 (N_7175,N_5322,N_6108);
xor U7176 (N_7176,N_5941,N_5204);
nand U7177 (N_7177,N_5823,N_5487);
nor U7178 (N_7178,N_6149,N_5819);
nand U7179 (N_7179,N_6215,N_6076);
and U7180 (N_7180,N_5834,N_6180);
nand U7181 (N_7181,N_5598,N_5628);
xnor U7182 (N_7182,N_6134,N_6230);
nand U7183 (N_7183,N_5620,N_5125);
nand U7184 (N_7184,N_5978,N_5762);
nand U7185 (N_7185,N_5140,N_5842);
nor U7186 (N_7186,N_6046,N_5696);
and U7187 (N_7187,N_5544,N_5343);
nor U7188 (N_7188,N_6112,N_5706);
xor U7189 (N_7189,N_5636,N_5583);
xnor U7190 (N_7190,N_5022,N_5376);
nand U7191 (N_7191,N_5369,N_6193);
nor U7192 (N_7192,N_5561,N_6247);
xor U7193 (N_7193,N_5063,N_5210);
and U7194 (N_7194,N_5822,N_5887);
xnor U7195 (N_7195,N_5550,N_5927);
or U7196 (N_7196,N_6006,N_5775);
nand U7197 (N_7197,N_5686,N_5710);
nand U7198 (N_7198,N_5789,N_6152);
and U7199 (N_7199,N_5931,N_5770);
xor U7200 (N_7200,N_5838,N_5159);
and U7201 (N_7201,N_5267,N_5573);
and U7202 (N_7202,N_5659,N_5038);
or U7203 (N_7203,N_5053,N_5664);
nand U7204 (N_7204,N_5758,N_5658);
and U7205 (N_7205,N_5975,N_5969);
and U7206 (N_7206,N_5146,N_5070);
or U7207 (N_7207,N_6012,N_5648);
or U7208 (N_7208,N_5607,N_5506);
xor U7209 (N_7209,N_5028,N_5114);
xor U7210 (N_7210,N_5105,N_5643);
nor U7211 (N_7211,N_5155,N_6248);
or U7212 (N_7212,N_5205,N_5875);
nand U7213 (N_7213,N_5266,N_6032);
xor U7214 (N_7214,N_5668,N_5639);
xnor U7215 (N_7215,N_5544,N_5991);
xor U7216 (N_7216,N_5760,N_5660);
nand U7217 (N_7217,N_5276,N_6190);
nor U7218 (N_7218,N_6071,N_5655);
nor U7219 (N_7219,N_6153,N_5261);
xor U7220 (N_7220,N_5976,N_5922);
and U7221 (N_7221,N_6237,N_5834);
xnor U7222 (N_7222,N_6097,N_5256);
nand U7223 (N_7223,N_5599,N_5385);
xnor U7224 (N_7224,N_5846,N_5380);
xor U7225 (N_7225,N_5127,N_5895);
and U7226 (N_7226,N_5679,N_5990);
or U7227 (N_7227,N_5639,N_5255);
xor U7228 (N_7228,N_6100,N_5316);
or U7229 (N_7229,N_5972,N_5455);
nor U7230 (N_7230,N_5800,N_5380);
or U7231 (N_7231,N_6175,N_5930);
nor U7232 (N_7232,N_5574,N_5047);
xnor U7233 (N_7233,N_5014,N_5739);
and U7234 (N_7234,N_5535,N_5859);
nand U7235 (N_7235,N_5580,N_6035);
and U7236 (N_7236,N_5723,N_5655);
nand U7237 (N_7237,N_5277,N_6209);
and U7238 (N_7238,N_6047,N_5048);
nor U7239 (N_7239,N_5841,N_6179);
nor U7240 (N_7240,N_6098,N_5546);
nor U7241 (N_7241,N_5498,N_5666);
xor U7242 (N_7242,N_6209,N_6152);
nor U7243 (N_7243,N_6049,N_5445);
xnor U7244 (N_7244,N_5545,N_5465);
nand U7245 (N_7245,N_5496,N_5848);
nand U7246 (N_7246,N_5592,N_5207);
and U7247 (N_7247,N_5368,N_5190);
nor U7248 (N_7248,N_5169,N_5178);
and U7249 (N_7249,N_6220,N_5200);
xnor U7250 (N_7250,N_5322,N_5464);
nor U7251 (N_7251,N_6157,N_5276);
nand U7252 (N_7252,N_5858,N_6197);
or U7253 (N_7253,N_5630,N_5933);
xor U7254 (N_7254,N_5020,N_5286);
or U7255 (N_7255,N_5916,N_5802);
and U7256 (N_7256,N_5264,N_6102);
or U7257 (N_7257,N_5263,N_5959);
nor U7258 (N_7258,N_5024,N_5738);
nor U7259 (N_7259,N_5524,N_5487);
or U7260 (N_7260,N_5435,N_5183);
nand U7261 (N_7261,N_6123,N_5816);
or U7262 (N_7262,N_5961,N_5836);
nand U7263 (N_7263,N_5935,N_5652);
nand U7264 (N_7264,N_5918,N_5429);
nor U7265 (N_7265,N_5112,N_5114);
nor U7266 (N_7266,N_5677,N_5558);
nor U7267 (N_7267,N_6210,N_5132);
or U7268 (N_7268,N_6220,N_5948);
nor U7269 (N_7269,N_5619,N_5867);
nand U7270 (N_7270,N_5274,N_5710);
nand U7271 (N_7271,N_6012,N_6033);
nand U7272 (N_7272,N_5753,N_5202);
nor U7273 (N_7273,N_5457,N_5187);
nand U7274 (N_7274,N_5466,N_5035);
and U7275 (N_7275,N_5759,N_5792);
xnor U7276 (N_7276,N_6076,N_5166);
xor U7277 (N_7277,N_6193,N_5266);
xor U7278 (N_7278,N_5470,N_5462);
nand U7279 (N_7279,N_5981,N_5928);
xnor U7280 (N_7280,N_6199,N_5390);
and U7281 (N_7281,N_5430,N_5855);
nor U7282 (N_7282,N_5957,N_6013);
and U7283 (N_7283,N_5077,N_5839);
xnor U7284 (N_7284,N_5397,N_5391);
xor U7285 (N_7285,N_5961,N_6175);
and U7286 (N_7286,N_5642,N_5824);
nand U7287 (N_7287,N_5582,N_5489);
nor U7288 (N_7288,N_5747,N_5607);
xor U7289 (N_7289,N_5869,N_5582);
nand U7290 (N_7290,N_5798,N_6034);
xor U7291 (N_7291,N_5771,N_5146);
or U7292 (N_7292,N_5324,N_5937);
xnor U7293 (N_7293,N_5879,N_5994);
xnor U7294 (N_7294,N_5452,N_5492);
nor U7295 (N_7295,N_6080,N_5886);
or U7296 (N_7296,N_5697,N_5380);
nor U7297 (N_7297,N_6098,N_5048);
nor U7298 (N_7298,N_5733,N_5570);
xnor U7299 (N_7299,N_5398,N_5351);
or U7300 (N_7300,N_5152,N_5965);
nor U7301 (N_7301,N_5664,N_5345);
or U7302 (N_7302,N_5744,N_5784);
and U7303 (N_7303,N_5002,N_5181);
xor U7304 (N_7304,N_5534,N_5485);
xnor U7305 (N_7305,N_5720,N_5015);
nor U7306 (N_7306,N_5713,N_6028);
or U7307 (N_7307,N_5714,N_6055);
nand U7308 (N_7308,N_5010,N_5142);
nor U7309 (N_7309,N_5510,N_5700);
or U7310 (N_7310,N_5048,N_5961);
or U7311 (N_7311,N_5919,N_5537);
and U7312 (N_7312,N_5026,N_5925);
and U7313 (N_7313,N_6181,N_5095);
nor U7314 (N_7314,N_5646,N_6078);
and U7315 (N_7315,N_5227,N_5564);
or U7316 (N_7316,N_5630,N_5408);
and U7317 (N_7317,N_5760,N_6058);
nor U7318 (N_7318,N_6164,N_6144);
xnor U7319 (N_7319,N_5679,N_5111);
and U7320 (N_7320,N_5078,N_5262);
or U7321 (N_7321,N_5665,N_5275);
or U7322 (N_7322,N_6156,N_5107);
nand U7323 (N_7323,N_6151,N_5088);
or U7324 (N_7324,N_5740,N_5185);
nor U7325 (N_7325,N_5661,N_5915);
nand U7326 (N_7326,N_6037,N_5243);
nand U7327 (N_7327,N_5572,N_6110);
nand U7328 (N_7328,N_5747,N_5613);
nor U7329 (N_7329,N_5478,N_5551);
nand U7330 (N_7330,N_5813,N_6126);
and U7331 (N_7331,N_5329,N_5580);
nand U7332 (N_7332,N_5373,N_5401);
and U7333 (N_7333,N_5326,N_6007);
or U7334 (N_7334,N_5412,N_5720);
nor U7335 (N_7335,N_5963,N_5945);
xor U7336 (N_7336,N_5413,N_5218);
nand U7337 (N_7337,N_5298,N_5136);
and U7338 (N_7338,N_5948,N_5011);
and U7339 (N_7339,N_5432,N_5763);
or U7340 (N_7340,N_6032,N_6145);
and U7341 (N_7341,N_6020,N_6044);
or U7342 (N_7342,N_5643,N_6012);
nor U7343 (N_7343,N_5171,N_5215);
nor U7344 (N_7344,N_6059,N_5094);
nand U7345 (N_7345,N_5475,N_5181);
nand U7346 (N_7346,N_6140,N_5573);
xnor U7347 (N_7347,N_6080,N_6024);
nand U7348 (N_7348,N_5126,N_5322);
or U7349 (N_7349,N_5557,N_5678);
nor U7350 (N_7350,N_5888,N_5677);
xor U7351 (N_7351,N_5253,N_5563);
xnor U7352 (N_7352,N_6060,N_5707);
nand U7353 (N_7353,N_5502,N_5742);
and U7354 (N_7354,N_5372,N_5273);
and U7355 (N_7355,N_6151,N_5038);
or U7356 (N_7356,N_5545,N_5399);
and U7357 (N_7357,N_5034,N_5431);
xnor U7358 (N_7358,N_5313,N_5269);
xor U7359 (N_7359,N_6245,N_5021);
nor U7360 (N_7360,N_5229,N_5741);
xor U7361 (N_7361,N_6060,N_5144);
or U7362 (N_7362,N_6077,N_5845);
and U7363 (N_7363,N_5955,N_6096);
and U7364 (N_7364,N_5264,N_6191);
nand U7365 (N_7365,N_5207,N_5753);
xor U7366 (N_7366,N_5626,N_5248);
nor U7367 (N_7367,N_5621,N_5097);
nor U7368 (N_7368,N_5662,N_5152);
nor U7369 (N_7369,N_5676,N_5741);
and U7370 (N_7370,N_5737,N_5243);
and U7371 (N_7371,N_5713,N_5041);
nor U7372 (N_7372,N_5415,N_5443);
nor U7373 (N_7373,N_5158,N_6093);
or U7374 (N_7374,N_6032,N_5339);
and U7375 (N_7375,N_5708,N_5179);
nand U7376 (N_7376,N_5612,N_5721);
nor U7377 (N_7377,N_5058,N_5952);
or U7378 (N_7378,N_5870,N_5395);
xor U7379 (N_7379,N_6012,N_5272);
nor U7380 (N_7380,N_5810,N_5307);
nor U7381 (N_7381,N_5529,N_6062);
and U7382 (N_7382,N_5984,N_5768);
and U7383 (N_7383,N_5477,N_5245);
xnor U7384 (N_7384,N_5853,N_5989);
nor U7385 (N_7385,N_5841,N_5960);
xor U7386 (N_7386,N_5935,N_5150);
or U7387 (N_7387,N_5618,N_5283);
or U7388 (N_7388,N_5041,N_6051);
xor U7389 (N_7389,N_5442,N_5955);
nand U7390 (N_7390,N_5301,N_5947);
and U7391 (N_7391,N_5029,N_5625);
or U7392 (N_7392,N_5868,N_5155);
and U7393 (N_7393,N_5727,N_6132);
nor U7394 (N_7394,N_5560,N_5655);
or U7395 (N_7395,N_5311,N_5922);
and U7396 (N_7396,N_5463,N_5180);
and U7397 (N_7397,N_6123,N_5157);
xnor U7398 (N_7398,N_5063,N_6084);
or U7399 (N_7399,N_5650,N_5546);
and U7400 (N_7400,N_5069,N_5709);
nand U7401 (N_7401,N_5130,N_5864);
nor U7402 (N_7402,N_5792,N_6147);
or U7403 (N_7403,N_5906,N_5158);
xnor U7404 (N_7404,N_5198,N_5693);
nor U7405 (N_7405,N_6033,N_5171);
xor U7406 (N_7406,N_6245,N_5840);
nand U7407 (N_7407,N_5944,N_5555);
and U7408 (N_7408,N_5330,N_5897);
and U7409 (N_7409,N_5614,N_5488);
and U7410 (N_7410,N_6025,N_5372);
nor U7411 (N_7411,N_5565,N_5194);
nand U7412 (N_7412,N_5225,N_5238);
and U7413 (N_7413,N_5233,N_5743);
nand U7414 (N_7414,N_5080,N_6202);
and U7415 (N_7415,N_5036,N_5165);
nor U7416 (N_7416,N_5868,N_5024);
nor U7417 (N_7417,N_5414,N_5156);
or U7418 (N_7418,N_5542,N_5960);
xor U7419 (N_7419,N_5591,N_5005);
xor U7420 (N_7420,N_6062,N_5951);
nor U7421 (N_7421,N_5472,N_5241);
nand U7422 (N_7422,N_5729,N_6177);
and U7423 (N_7423,N_5798,N_5214);
nor U7424 (N_7424,N_5060,N_5435);
xor U7425 (N_7425,N_6168,N_5449);
nor U7426 (N_7426,N_5470,N_6097);
nand U7427 (N_7427,N_5619,N_5294);
or U7428 (N_7428,N_5208,N_5077);
or U7429 (N_7429,N_6206,N_6126);
nand U7430 (N_7430,N_5648,N_6237);
or U7431 (N_7431,N_6228,N_6246);
nor U7432 (N_7432,N_5552,N_5931);
or U7433 (N_7433,N_6025,N_5201);
and U7434 (N_7434,N_5813,N_5114);
nor U7435 (N_7435,N_5810,N_6213);
or U7436 (N_7436,N_5565,N_5643);
nand U7437 (N_7437,N_5631,N_5692);
or U7438 (N_7438,N_6211,N_5354);
and U7439 (N_7439,N_5408,N_6081);
nor U7440 (N_7440,N_5589,N_6238);
nor U7441 (N_7441,N_5377,N_6184);
or U7442 (N_7442,N_5378,N_5219);
and U7443 (N_7443,N_6030,N_5135);
or U7444 (N_7444,N_5123,N_5301);
nand U7445 (N_7445,N_5489,N_5452);
and U7446 (N_7446,N_6189,N_6038);
xor U7447 (N_7447,N_6207,N_5235);
nor U7448 (N_7448,N_5943,N_5346);
and U7449 (N_7449,N_5069,N_5661);
nand U7450 (N_7450,N_5933,N_6238);
nand U7451 (N_7451,N_5644,N_5443);
nand U7452 (N_7452,N_5508,N_5133);
nor U7453 (N_7453,N_5233,N_6052);
nor U7454 (N_7454,N_5034,N_6247);
xnor U7455 (N_7455,N_5770,N_5894);
or U7456 (N_7456,N_5763,N_6244);
and U7457 (N_7457,N_5231,N_5392);
and U7458 (N_7458,N_6195,N_6086);
or U7459 (N_7459,N_5830,N_5728);
xnor U7460 (N_7460,N_6192,N_5872);
or U7461 (N_7461,N_5435,N_5555);
and U7462 (N_7462,N_5966,N_5265);
nor U7463 (N_7463,N_5789,N_5782);
nand U7464 (N_7464,N_5304,N_5988);
xor U7465 (N_7465,N_5704,N_5583);
xor U7466 (N_7466,N_5928,N_5447);
nor U7467 (N_7467,N_5741,N_5278);
nor U7468 (N_7468,N_5985,N_5090);
nor U7469 (N_7469,N_5342,N_5581);
or U7470 (N_7470,N_5064,N_6237);
and U7471 (N_7471,N_5011,N_5185);
or U7472 (N_7472,N_5165,N_5223);
nor U7473 (N_7473,N_5651,N_5172);
and U7474 (N_7474,N_6135,N_6236);
nor U7475 (N_7475,N_6039,N_6225);
and U7476 (N_7476,N_5731,N_6166);
xnor U7477 (N_7477,N_6152,N_5519);
or U7478 (N_7478,N_5336,N_5904);
xor U7479 (N_7479,N_5247,N_5265);
nor U7480 (N_7480,N_5509,N_6068);
nand U7481 (N_7481,N_5374,N_5887);
nor U7482 (N_7482,N_5664,N_5554);
nor U7483 (N_7483,N_5404,N_5811);
and U7484 (N_7484,N_6237,N_5512);
or U7485 (N_7485,N_6116,N_5646);
nor U7486 (N_7486,N_5473,N_6106);
or U7487 (N_7487,N_5126,N_5365);
nor U7488 (N_7488,N_5908,N_5412);
or U7489 (N_7489,N_5391,N_6073);
or U7490 (N_7490,N_5596,N_5021);
or U7491 (N_7491,N_5335,N_5007);
or U7492 (N_7492,N_5590,N_5356);
xnor U7493 (N_7493,N_5636,N_5046);
or U7494 (N_7494,N_5346,N_6127);
or U7495 (N_7495,N_5693,N_6067);
and U7496 (N_7496,N_5452,N_5512);
nand U7497 (N_7497,N_6155,N_5915);
and U7498 (N_7498,N_5338,N_5941);
or U7499 (N_7499,N_5968,N_5663);
and U7500 (N_7500,N_6744,N_6548);
nor U7501 (N_7501,N_6718,N_7278);
xnor U7502 (N_7502,N_7304,N_6316);
xnor U7503 (N_7503,N_6863,N_7365);
and U7504 (N_7504,N_7313,N_6476);
and U7505 (N_7505,N_7458,N_6253);
nor U7506 (N_7506,N_7036,N_6262);
and U7507 (N_7507,N_7494,N_6934);
or U7508 (N_7508,N_6828,N_7455);
or U7509 (N_7509,N_6489,N_6766);
nor U7510 (N_7510,N_6662,N_6545);
and U7511 (N_7511,N_7100,N_7024);
nor U7512 (N_7512,N_6857,N_6319);
nand U7513 (N_7513,N_6963,N_6571);
and U7514 (N_7514,N_6357,N_6492);
xnor U7515 (N_7515,N_6944,N_7223);
xnor U7516 (N_7516,N_6398,N_6380);
nor U7517 (N_7517,N_7293,N_6425);
or U7518 (N_7518,N_6700,N_6608);
or U7519 (N_7519,N_6778,N_6692);
nor U7520 (N_7520,N_6855,N_6682);
nand U7521 (N_7521,N_6534,N_6366);
nand U7522 (N_7522,N_7316,N_7337);
or U7523 (N_7523,N_6802,N_7046);
xnor U7524 (N_7524,N_7208,N_6600);
or U7525 (N_7525,N_7355,N_7212);
or U7526 (N_7526,N_7136,N_7010);
nand U7527 (N_7527,N_6767,N_7126);
nand U7528 (N_7528,N_6730,N_7361);
nor U7529 (N_7529,N_6279,N_7194);
or U7530 (N_7530,N_6844,N_6404);
and U7531 (N_7531,N_7146,N_6549);
nand U7532 (N_7532,N_7075,N_6379);
or U7533 (N_7533,N_7470,N_6332);
and U7534 (N_7534,N_6735,N_6845);
or U7535 (N_7535,N_6593,N_6506);
nand U7536 (N_7536,N_7490,N_6475);
xor U7537 (N_7537,N_6756,N_7157);
nor U7538 (N_7538,N_6385,N_7368);
and U7539 (N_7539,N_6986,N_6340);
nor U7540 (N_7540,N_7182,N_6979);
or U7541 (N_7541,N_6301,N_6625);
xnor U7542 (N_7542,N_7250,N_6868);
xor U7543 (N_7543,N_7386,N_7043);
and U7544 (N_7544,N_6479,N_7122);
xor U7545 (N_7545,N_7413,N_6617);
nor U7546 (N_7546,N_7362,N_6813);
xnor U7547 (N_7547,N_7169,N_7346);
xor U7548 (N_7548,N_6999,N_6895);
nor U7549 (N_7549,N_7375,N_6620);
or U7550 (N_7550,N_6921,N_6418);
nor U7551 (N_7551,N_7161,N_6915);
or U7552 (N_7552,N_7281,N_6302);
nor U7553 (N_7553,N_6712,N_6790);
and U7554 (N_7554,N_7451,N_6837);
xnor U7555 (N_7555,N_7256,N_7391);
nor U7556 (N_7556,N_6515,N_7429);
or U7557 (N_7557,N_7061,N_6974);
or U7558 (N_7558,N_6629,N_6990);
xnor U7559 (N_7559,N_6360,N_6364);
xnor U7560 (N_7560,N_6602,N_7341);
or U7561 (N_7561,N_6519,N_7254);
xor U7562 (N_7562,N_7497,N_6776);
and U7563 (N_7563,N_6315,N_7094);
and U7564 (N_7564,N_7031,N_7128);
nor U7565 (N_7565,N_6912,N_6377);
nor U7566 (N_7566,N_7310,N_7311);
or U7567 (N_7567,N_6763,N_7242);
xnor U7568 (N_7568,N_6993,N_6502);
or U7569 (N_7569,N_6378,N_6856);
or U7570 (N_7570,N_6444,N_7183);
and U7571 (N_7571,N_7037,N_6458);
or U7572 (N_7572,N_7119,N_6526);
and U7573 (N_7573,N_6254,N_6498);
nand U7574 (N_7574,N_6334,N_6553);
xnor U7575 (N_7575,N_6890,N_7175);
or U7576 (N_7576,N_6699,N_7220);
and U7577 (N_7577,N_6591,N_7407);
and U7578 (N_7578,N_7132,N_6565);
nor U7579 (N_7579,N_6948,N_6356);
nand U7580 (N_7580,N_6395,N_7257);
nor U7581 (N_7581,N_6647,N_6293);
nor U7582 (N_7582,N_6995,N_7213);
and U7583 (N_7583,N_6327,N_6920);
nand U7584 (N_7584,N_6297,N_6815);
nor U7585 (N_7585,N_7308,N_6768);
nand U7586 (N_7586,N_6968,N_6977);
nor U7587 (N_7587,N_7403,N_6831);
xnor U7588 (N_7588,N_6349,N_6369);
nand U7589 (N_7589,N_6850,N_6611);
and U7590 (N_7590,N_6525,N_6323);
xnor U7591 (N_7591,N_7335,N_6757);
xnor U7592 (N_7592,N_6787,N_6630);
nand U7593 (N_7593,N_7356,N_6482);
nor U7594 (N_7594,N_6814,N_6717);
xor U7595 (N_7595,N_7457,N_7487);
or U7596 (N_7596,N_6582,N_6503);
nand U7597 (N_7597,N_6533,N_7493);
and U7598 (N_7598,N_6820,N_6905);
nor U7599 (N_7599,N_6447,N_7447);
nor U7600 (N_7600,N_6312,N_6307);
nor U7601 (N_7601,N_6347,N_7301);
nand U7602 (N_7602,N_7035,N_7013);
or U7603 (N_7603,N_6453,N_6930);
or U7604 (N_7604,N_7399,N_6528);
and U7605 (N_7605,N_6842,N_6936);
xor U7606 (N_7606,N_6732,N_6772);
or U7607 (N_7607,N_7460,N_7428);
nand U7608 (N_7608,N_7088,N_7081);
nor U7609 (N_7609,N_7070,N_7478);
xor U7610 (N_7610,N_7296,N_7397);
and U7611 (N_7611,N_6685,N_6803);
nor U7612 (N_7612,N_6733,N_7057);
or U7613 (N_7613,N_7319,N_7071);
and U7614 (N_7614,N_6881,N_7306);
or U7615 (N_7615,N_6740,N_6711);
nor U7616 (N_7616,N_7420,N_6439);
or U7617 (N_7617,N_6370,N_6816);
and U7618 (N_7618,N_6908,N_7229);
xnor U7619 (N_7619,N_6605,N_7097);
nor U7620 (N_7620,N_7402,N_7144);
xor U7621 (N_7621,N_6780,N_6691);
nor U7622 (N_7622,N_6885,N_7258);
and U7623 (N_7623,N_7450,N_6998);
and U7624 (N_7624,N_6367,N_7042);
and U7625 (N_7625,N_6913,N_7093);
or U7626 (N_7626,N_6409,N_6997);
or U7627 (N_7627,N_6461,N_6806);
nor U7628 (N_7628,N_7430,N_6636);
xnor U7629 (N_7629,N_6403,N_6989);
nand U7630 (N_7630,N_6562,N_7372);
and U7631 (N_7631,N_6296,N_6626);
and U7632 (N_7632,N_7090,N_6273);
xor U7633 (N_7633,N_6865,N_6697);
xor U7634 (N_7634,N_6960,N_7369);
nor U7635 (N_7635,N_6531,N_7444);
and U7636 (N_7636,N_6290,N_6640);
nand U7637 (N_7637,N_7202,N_6976);
xor U7638 (N_7638,N_6910,N_6781);
or U7639 (N_7639,N_6826,N_6959);
and U7640 (N_7640,N_6683,N_6318);
xor U7641 (N_7641,N_6670,N_6622);
nand U7642 (N_7642,N_7324,N_7082);
xnor U7643 (N_7643,N_6573,N_6566);
nor U7644 (N_7644,N_6961,N_6484);
nand U7645 (N_7645,N_7239,N_7154);
and U7646 (N_7646,N_6308,N_6259);
and U7647 (N_7647,N_6665,N_6333);
nor U7648 (N_7648,N_6901,N_7436);
and U7649 (N_7649,N_6753,N_7387);
or U7650 (N_7650,N_7411,N_6456);
or U7651 (N_7651,N_6300,N_6496);
xor U7652 (N_7652,N_7072,N_7464);
nor U7653 (N_7653,N_7181,N_7472);
nand U7654 (N_7654,N_7234,N_6788);
or U7655 (N_7655,N_6423,N_6615);
nand U7656 (N_7656,N_7153,N_6650);
and U7657 (N_7657,N_6338,N_6587);
xor U7658 (N_7658,N_7163,N_6657);
nand U7659 (N_7659,N_7376,N_6853);
xor U7660 (N_7660,N_6486,N_7338);
xor U7661 (N_7661,N_7095,N_6987);
nand U7662 (N_7662,N_7395,N_7323);
nor U7663 (N_7663,N_6554,N_6951);
nand U7664 (N_7664,N_6572,N_6906);
or U7665 (N_7665,N_6460,N_6433);
xor U7666 (N_7666,N_6282,N_6835);
xnor U7667 (N_7667,N_6914,N_7357);
nand U7668 (N_7668,N_6362,N_6745);
or U7669 (N_7669,N_7240,N_6497);
nor U7670 (N_7670,N_7244,N_6560);
xnor U7671 (N_7671,N_6755,N_6516);
or U7672 (N_7672,N_6263,N_6288);
or U7673 (N_7673,N_6372,N_7408);
and U7674 (N_7674,N_6544,N_6624);
xnor U7675 (N_7675,N_7063,N_6436);
nor U7676 (N_7676,N_6680,N_7080);
nand U7677 (N_7677,N_6775,N_7328);
nor U7678 (N_7678,N_7412,N_6435);
nand U7679 (N_7679,N_7066,N_6874);
and U7680 (N_7680,N_6564,N_7174);
nand U7681 (N_7681,N_7445,N_7262);
or U7682 (N_7682,N_7468,N_7047);
nand U7683 (N_7683,N_6722,N_6504);
and U7684 (N_7684,N_6546,N_6774);
and U7685 (N_7685,N_7235,N_6322);
or U7686 (N_7686,N_7120,N_6441);
and U7687 (N_7687,N_7400,N_6511);
nor U7688 (N_7688,N_7343,N_6406);
and U7689 (N_7689,N_7180,N_6298);
nand U7690 (N_7690,N_6883,N_6452);
nor U7691 (N_7691,N_6938,N_6801);
nor U7692 (N_7692,N_7367,N_7378);
and U7693 (N_7693,N_7315,N_6558);
and U7694 (N_7694,N_6747,N_7064);
nor U7695 (N_7695,N_7023,N_7152);
nand U7696 (N_7696,N_6884,N_6454);
or U7697 (N_7697,N_6373,N_7012);
nor U7698 (N_7698,N_7192,N_7265);
and U7699 (N_7699,N_7243,N_7252);
and U7700 (N_7700,N_6337,N_6759);
or U7701 (N_7701,N_7465,N_6306);
nand U7702 (N_7702,N_7204,N_7384);
and U7703 (N_7703,N_7251,N_6672);
and U7704 (N_7704,N_6720,N_6500);
xor U7705 (N_7705,N_6947,N_6879);
xor U7706 (N_7706,N_7442,N_6524);
and U7707 (N_7707,N_6607,N_7314);
nand U7708 (N_7708,N_6686,N_6785);
or U7709 (N_7709,N_7350,N_7205);
or U7710 (N_7710,N_7237,N_6595);
or U7711 (N_7711,N_6320,N_6443);
and U7712 (N_7712,N_7019,N_6494);
xor U7713 (N_7713,N_6400,N_6387);
xor U7714 (N_7714,N_7489,N_6677);
xnor U7715 (N_7715,N_6688,N_7419);
or U7716 (N_7716,N_7140,N_6576);
and U7717 (N_7717,N_7004,N_6950);
xnor U7718 (N_7718,N_6474,N_6668);
nor U7719 (N_7719,N_6632,N_7446);
nor U7720 (N_7720,N_7302,N_7438);
or U7721 (N_7721,N_6962,N_6749);
xor U7722 (N_7722,N_6501,N_6427);
or U7723 (N_7723,N_6705,N_6782);
and U7724 (N_7724,N_7422,N_6358);
and U7725 (N_7725,N_7137,N_7320);
xnor U7726 (N_7726,N_7459,N_6941);
nand U7727 (N_7727,N_7172,N_6750);
nor U7728 (N_7728,N_6840,N_6690);
or U7729 (N_7729,N_6764,N_6389);
nand U7730 (N_7730,N_6634,N_6597);
xnor U7731 (N_7731,N_6655,N_6876);
and U7732 (N_7732,N_6667,N_7317);
nand U7733 (N_7733,N_6746,N_6610);
and U7734 (N_7734,N_6361,N_6848);
nand U7735 (N_7735,N_7016,N_7077);
or U7736 (N_7736,N_7110,N_7309);
and U7737 (N_7737,N_6639,N_7474);
and U7738 (N_7738,N_7147,N_6946);
or U7739 (N_7739,N_7435,N_6555);
xnor U7740 (N_7740,N_6487,N_6585);
or U7741 (N_7741,N_6869,N_7363);
nor U7742 (N_7742,N_6825,N_7170);
and U7743 (N_7743,N_6859,N_7114);
or U7744 (N_7744,N_6911,N_6783);
xnor U7745 (N_7745,N_7032,N_7390);
nor U7746 (N_7746,N_7006,N_6994);
nand U7747 (N_7747,N_6949,N_6527);
xor U7748 (N_7748,N_7034,N_7273);
xor U7749 (N_7749,N_7233,N_6725);
and U7750 (N_7750,N_7449,N_6568);
nand U7751 (N_7751,N_6469,N_6383);
or U7752 (N_7752,N_7421,N_6687);
or U7753 (N_7753,N_7168,N_6898);
or U7754 (N_7754,N_6653,N_6638);
xnor U7755 (N_7755,N_7145,N_6265);
nand U7756 (N_7756,N_6886,N_6726);
xnor U7757 (N_7757,N_6939,N_6368);
xor U7758 (N_7758,N_7342,N_6547);
and U7759 (N_7759,N_6937,N_7210);
and U7760 (N_7760,N_7481,N_7427);
nand U7761 (N_7761,N_7186,N_6352);
and U7762 (N_7762,N_7156,N_6721);
xnor U7763 (N_7763,N_6541,N_6748);
or U7764 (N_7764,N_7065,N_6980);
or U7765 (N_7765,N_7050,N_7330);
or U7766 (N_7766,N_6738,N_7206);
and U7767 (N_7767,N_7188,N_7184);
or U7768 (N_7768,N_7260,N_6945);
and U7769 (N_7769,N_6613,N_6707);
nor U7770 (N_7770,N_6536,N_6335);
xor U7771 (N_7771,N_6678,N_7483);
or U7772 (N_7772,N_6286,N_7219);
nand U7773 (N_7773,N_6574,N_6399);
and U7774 (N_7774,N_7025,N_6715);
nand U7775 (N_7775,N_7373,N_7155);
or U7776 (N_7776,N_6978,N_6769);
nand U7777 (N_7777,N_6483,N_7045);
nor U7778 (N_7778,N_6648,N_6462);
and U7779 (N_7779,N_6810,N_6819);
xor U7780 (N_7780,N_7087,N_7415);
or U7781 (N_7781,N_7467,N_7414);
and U7782 (N_7782,N_7022,N_6751);
or U7783 (N_7783,N_7084,N_7086);
xor U7784 (N_7784,N_6255,N_6698);
and U7785 (N_7785,N_7134,N_7287);
nand U7786 (N_7786,N_6982,N_7284);
xor U7787 (N_7787,N_6275,N_6804);
xnor U7788 (N_7788,N_7117,N_7060);
nand U7789 (N_7789,N_6392,N_6909);
nand U7790 (N_7790,N_6927,N_6933);
or U7791 (N_7791,N_6342,N_6649);
nor U7792 (N_7792,N_6684,N_7021);
or U7793 (N_7793,N_7018,N_6713);
or U7794 (N_7794,N_6451,N_6644);
nor U7795 (N_7795,N_6538,N_6737);
xnor U7796 (N_7796,N_6919,N_6419);
nand U7797 (N_7797,N_6925,N_6867);
xnor U7798 (N_7798,N_6467,N_7111);
nor U7799 (N_7799,N_7300,N_7039);
nand U7800 (N_7800,N_6584,N_7392);
xnor U7801 (N_7801,N_7129,N_6345);
and U7802 (N_7802,N_7104,N_7150);
nor U7803 (N_7803,N_7339,N_6952);
xnor U7804 (N_7804,N_7448,N_6354);
xnor U7805 (N_7805,N_6614,N_6956);
nor U7806 (N_7806,N_6260,N_6429);
xor U7807 (N_7807,N_6971,N_6932);
nor U7808 (N_7808,N_7041,N_6343);
and U7809 (N_7809,N_6935,N_7165);
and U7810 (N_7810,N_6463,N_6818);
nand U7811 (N_7811,N_6900,N_6795);
or U7812 (N_7812,N_7048,N_6556);
nand U7813 (N_7813,N_6627,N_6955);
or U7814 (N_7814,N_6437,N_7198);
xor U7815 (N_7815,N_6535,N_7171);
xnor U7816 (N_7816,N_6264,N_7462);
and U7817 (N_7817,N_6359,N_7196);
xor U7818 (N_7818,N_7381,N_7345);
nor U7819 (N_7819,N_6637,N_6983);
nand U7820 (N_7820,N_7026,N_7014);
nor U7821 (N_7821,N_7000,N_6512);
and U7822 (N_7822,N_7276,N_6832);
or U7823 (N_7823,N_6917,N_6896);
nor U7824 (N_7824,N_6539,N_7406);
xor U7825 (N_7825,N_6659,N_7103);
and U7826 (N_7826,N_7005,N_7499);
nor U7827 (N_7827,N_6311,N_6807);
and U7828 (N_7828,N_6967,N_6922);
or U7829 (N_7829,N_7389,N_7469);
nand U7830 (N_7830,N_6739,N_6331);
xnor U7831 (N_7831,N_7167,N_6811);
xnor U7832 (N_7832,N_6660,N_7437);
xor U7833 (N_7833,N_6480,N_7141);
nand U7834 (N_7834,N_6827,N_7359);
and U7835 (N_7835,N_6251,N_6346);
nor U7836 (N_7836,N_6376,N_6916);
nor U7837 (N_7837,N_6645,N_6401);
xor U7838 (N_7838,N_7432,N_6621);
nor U7839 (N_7839,N_7133,N_6428);
and U7840 (N_7840,N_6996,N_7347);
or U7841 (N_7841,N_6523,N_6702);
nor U7842 (N_7842,N_7101,N_6542);
or U7843 (N_7843,N_6770,N_6988);
or U7844 (N_7844,N_7292,N_7106);
or U7845 (N_7845,N_7193,N_6877);
nand U7846 (N_7846,N_6731,N_6557);
nor U7847 (N_7847,N_7079,N_6864);
or U7848 (N_7848,N_6341,N_6822);
xnor U7849 (N_7849,N_6791,N_6674);
and U7850 (N_7850,N_7216,N_6870);
nor U7851 (N_7851,N_7227,N_7238);
and U7852 (N_7852,N_7340,N_7221);
and U7853 (N_7853,N_6953,N_6550);
xor U7854 (N_7854,N_7195,N_7318);
xor U7855 (N_7855,N_7479,N_7073);
xnor U7856 (N_7856,N_6817,N_7279);
nor U7857 (N_7857,N_6654,N_7360);
and U7858 (N_7858,N_7008,N_7271);
and U7859 (N_7859,N_7289,N_7108);
and U7860 (N_7860,N_7349,N_7211);
xor U7861 (N_7861,N_7272,N_7336);
nand U7862 (N_7862,N_7149,N_7326);
nand U7863 (N_7863,N_7148,N_6631);
xnor U7864 (N_7864,N_7374,N_7054);
xnor U7865 (N_7865,N_7473,N_7139);
nor U7866 (N_7866,N_7417,N_7040);
and U7867 (N_7867,N_6762,N_6330);
or U7868 (N_7868,N_6727,N_6348);
and U7869 (N_7869,N_7249,N_7476);
nor U7870 (N_7870,N_6796,N_7370);
or U7871 (N_7871,N_7076,N_7404);
nand U7872 (N_7872,N_6269,N_6723);
nor U7873 (N_7873,N_6284,N_6507);
xor U7874 (N_7874,N_7164,N_6570);
xor U7875 (N_7875,N_7201,N_6271);
nor U7876 (N_7876,N_6488,N_7297);
and U7877 (N_7877,N_7113,N_7398);
and U7878 (N_7878,N_6413,N_6289);
or U7879 (N_7879,N_6601,N_7142);
or U7880 (N_7880,N_7091,N_7380);
xnor U7881 (N_7881,N_6339,N_7344);
xnor U7882 (N_7882,N_7379,N_6405);
or U7883 (N_7883,N_6450,N_6847);
xnor U7884 (N_7884,N_6664,N_7290);
nand U7885 (N_7885,N_7052,N_6426);
nand U7886 (N_7886,N_7059,N_6256);
or U7887 (N_7887,N_7454,N_7354);
or U7888 (N_7888,N_6777,N_7015);
or U7889 (N_7889,N_6765,N_7049);
or U7890 (N_7890,N_6431,N_6798);
or U7891 (N_7891,N_6481,N_6442);
xor U7892 (N_7892,N_6800,N_6590);
or U7893 (N_7893,N_6887,N_6681);
nor U7894 (N_7894,N_6563,N_6371);
nor U7895 (N_7895,N_6924,N_7441);
or U7896 (N_7896,N_7083,N_7189);
xor U7897 (N_7897,N_6514,N_6841);
nor U7898 (N_7898,N_6477,N_7396);
nor U7899 (N_7899,N_7162,N_6799);
and U7900 (N_7900,N_7452,N_7173);
and U7901 (N_7901,N_6623,N_6305);
and U7902 (N_7902,N_7200,N_6420);
nand U7903 (N_7903,N_6742,N_6278);
xor U7904 (N_7904,N_6313,N_6943);
nand U7905 (N_7905,N_6789,N_7056);
nand U7906 (N_7906,N_6871,N_6412);
and U7907 (N_7907,N_7332,N_6981);
xor U7908 (N_7908,N_6635,N_7366);
xnor U7909 (N_7909,N_6729,N_6295);
and U7910 (N_7910,N_6382,N_6388);
or U7911 (N_7911,N_6455,N_6396);
or U7912 (N_7912,N_6336,N_6415);
or U7913 (N_7913,N_6679,N_7028);
nor U7914 (N_7914,N_6432,N_7069);
xor U7915 (N_7915,N_7443,N_6518);
xor U7916 (N_7916,N_6561,N_6880);
or U7917 (N_7917,N_7187,N_6440);
and U7918 (N_7918,N_6446,N_6438);
nand U7919 (N_7919,N_6324,N_7253);
xnor U7920 (N_7920,N_6430,N_6643);
nand U7921 (N_7921,N_7352,N_7245);
nand U7922 (N_7922,N_7485,N_6969);
nand U7923 (N_7923,N_7416,N_6491);
xnor U7924 (N_7924,N_7003,N_6706);
nor U7925 (N_7925,N_7107,N_6728);
nor U7926 (N_7926,N_6618,N_6860);
nor U7927 (N_7927,N_7247,N_6658);
and U7928 (N_7928,N_7383,N_7246);
or U7929 (N_7929,N_6779,N_7007);
or U7930 (N_7930,N_7423,N_7053);
and U7931 (N_7931,N_6812,N_7099);
or U7932 (N_7932,N_6652,N_6694);
nor U7933 (N_7933,N_6465,N_6902);
nand U7934 (N_7934,N_6459,N_6508);
nor U7935 (N_7935,N_7203,N_6709);
and U7936 (N_7936,N_6493,N_6408);
xnor U7937 (N_7937,N_7085,N_7275);
nor U7938 (N_7938,N_6966,N_6589);
nand U7939 (N_7939,N_7267,N_7394);
nor U7940 (N_7940,N_6421,N_6466);
and U7941 (N_7941,N_6390,N_6351);
or U7942 (N_7942,N_6708,N_6522);
nand U7943 (N_7943,N_7001,N_6588);
xnor U7944 (N_7944,N_6992,N_6809);
nand U7945 (N_7945,N_7176,N_6823);
or U7946 (N_7946,N_6517,N_6716);
nor U7947 (N_7947,N_6292,N_7334);
xor U7948 (N_7948,N_7312,N_7215);
nand U7949 (N_7949,N_7185,N_7484);
or U7950 (N_7950,N_6675,N_7480);
nor U7951 (N_7951,N_6250,N_7353);
or U7952 (N_7952,N_7295,N_6386);
xnor U7953 (N_7953,N_6397,N_6872);
or U7954 (N_7954,N_6411,N_6821);
or U7955 (N_7955,N_6457,N_6252);
or U7956 (N_7956,N_6701,N_6888);
and U7957 (N_7957,N_7030,N_6317);
nand U7958 (N_7958,N_7135,N_7322);
nor U7959 (N_7959,N_6651,N_6410);
nand U7960 (N_7960,N_7440,N_7274);
or U7961 (N_7961,N_6878,N_6374);
nand U7962 (N_7962,N_7331,N_7329);
and U7963 (N_7963,N_7498,N_6267);
or U7964 (N_7964,N_6580,N_6314);
nand U7965 (N_7965,N_6266,N_6957);
nor U7966 (N_7966,N_7348,N_6794);
or U7967 (N_7967,N_7388,N_6918);
xor U7968 (N_7968,N_6309,N_6505);
or U7969 (N_7969,N_6329,N_6473);
or U7970 (N_7970,N_6521,N_6891);
or U7971 (N_7971,N_6363,N_7291);
xnor U7972 (N_7972,N_7199,N_6666);
nor U7973 (N_7973,N_6468,N_7418);
nor U7974 (N_7974,N_6606,N_6592);
nor U7975 (N_7975,N_6628,N_6581);
nor U7976 (N_7976,N_6609,N_7011);
and U7977 (N_7977,N_7492,N_6833);
and U7978 (N_7978,N_6530,N_7303);
nand U7979 (N_7979,N_7058,N_6280);
and U7980 (N_7980,N_6579,N_6274);
nand U7981 (N_7981,N_6808,N_6646);
nand U7982 (N_7982,N_6355,N_6771);
nor U7983 (N_7983,N_6854,N_6540);
nand U7984 (N_7984,N_7471,N_6598);
xor U7985 (N_7985,N_6985,N_7305);
or U7986 (N_7986,N_6858,N_7495);
or U7987 (N_7987,N_6830,N_6495);
xnor U7988 (N_7988,N_7283,N_7109);
or U7989 (N_7989,N_6894,N_7261);
or U7990 (N_7990,N_6276,N_6543);
nand U7991 (N_7991,N_6422,N_6695);
xor U7992 (N_7992,N_7385,N_6394);
nor U7993 (N_7993,N_7197,N_6942);
and U7994 (N_7994,N_6743,N_6270);
xnor U7995 (N_7995,N_6866,N_6464);
nand U7996 (N_7996,N_6586,N_7377);
nor U7997 (N_7997,N_7424,N_7307);
nand U7998 (N_7998,N_7051,N_6510);
and U7999 (N_7999,N_6656,N_7434);
or U8000 (N_8000,N_7160,N_6299);
xnor U8001 (N_8001,N_6719,N_6291);
or U8002 (N_8002,N_6575,N_7190);
nor U8003 (N_8003,N_6703,N_7020);
nor U8004 (N_8004,N_7461,N_6984);
nand U8005 (N_8005,N_7092,N_7225);
nand U8006 (N_8006,N_7143,N_6633);
nor U8007 (N_8007,N_7089,N_6381);
nand U8008 (N_8008,N_7074,N_6603);
xor U8009 (N_8009,N_6285,N_6964);
and U8010 (N_8010,N_7207,N_6907);
nor U8011 (N_8011,N_7209,N_7105);
and U8012 (N_8012,N_7067,N_6724);
nor U8013 (N_8013,N_7294,N_7269);
xnor U8014 (N_8014,N_6773,N_7466);
nor U8015 (N_8015,N_7044,N_6824);
xnor U8016 (N_8016,N_7364,N_6294);
xnor U8017 (N_8017,N_6310,N_6402);
nor U8018 (N_8018,N_7486,N_7426);
xor U8019 (N_8019,N_6669,N_7496);
nor U8020 (N_8020,N_6829,N_7268);
or U8021 (N_8021,N_7112,N_7062);
nand U8022 (N_8022,N_7280,N_6472);
and U8023 (N_8023,N_6604,N_6897);
and U8024 (N_8024,N_7029,N_7425);
and U8025 (N_8025,N_6975,N_6792);
nand U8026 (N_8026,N_7038,N_7230);
nor U8027 (N_8027,N_6478,N_7488);
and U8028 (N_8028,N_6758,N_6375);
or U8029 (N_8029,N_6836,N_7179);
and U8030 (N_8030,N_7002,N_7439);
nand U8031 (N_8031,N_6325,N_6760);
and U8032 (N_8032,N_6414,N_6797);
nor U8033 (N_8033,N_6671,N_6529);
xnor U8034 (N_8034,N_7393,N_7096);
xor U8035 (N_8035,N_7264,N_6350);
nand U8036 (N_8036,N_6882,N_6834);
xnor U8037 (N_8037,N_6520,N_6714);
or U8038 (N_8038,N_6257,N_7123);
and U8039 (N_8039,N_6786,N_6904);
xor U8040 (N_8040,N_6752,N_6304);
nor U8041 (N_8041,N_6424,N_6596);
nor U8042 (N_8042,N_6272,N_6958);
nand U8043 (N_8043,N_7098,N_6619);
or U8044 (N_8044,N_7232,N_6599);
or U8045 (N_8045,N_7236,N_6594);
xnor U8046 (N_8046,N_6499,N_7325);
xnor U8047 (N_8047,N_6852,N_6929);
nand U8048 (N_8048,N_6710,N_6873);
nand U8049 (N_8049,N_7125,N_7078);
nor U8050 (N_8050,N_6485,N_6663);
nand U8051 (N_8051,N_7382,N_7228);
nor U8052 (N_8052,N_6326,N_7259);
nand U8053 (N_8053,N_6559,N_7151);
nor U8054 (N_8054,N_6928,N_6861);
and U8055 (N_8055,N_6893,N_6849);
or U8056 (N_8056,N_6509,N_6612);
or U8057 (N_8057,N_7138,N_7282);
or U8058 (N_8058,N_6391,N_7009);
or U8059 (N_8059,N_6490,N_7327);
and U8060 (N_8060,N_7286,N_7288);
and U8061 (N_8061,N_6328,N_6889);
nor U8062 (N_8062,N_6552,N_7017);
or U8063 (N_8063,N_6537,N_6676);
and U8064 (N_8064,N_6551,N_6344);
nor U8065 (N_8065,N_6761,N_6734);
xor U8066 (N_8066,N_7491,N_7255);
xor U8067 (N_8067,N_7102,N_6892);
nor U8068 (N_8068,N_6616,N_6843);
nor U8069 (N_8069,N_7116,N_7118);
and U8070 (N_8070,N_6353,N_6642);
xor U8071 (N_8071,N_7159,N_6384);
nor U8072 (N_8072,N_6641,N_6940);
and U8073 (N_8073,N_7027,N_7285);
or U8074 (N_8074,N_7158,N_7214);
xor U8075 (N_8075,N_6583,N_7298);
nor U8076 (N_8076,N_7410,N_6513);
nor U8077 (N_8077,N_6434,N_7263);
or U8078 (N_8078,N_6577,N_6416);
or U8079 (N_8079,N_7222,N_6970);
or U8080 (N_8080,N_6805,N_6417);
or U8081 (N_8081,N_6449,N_7321);
or U8082 (N_8082,N_6578,N_7241);
xor U8083 (N_8083,N_6923,N_7477);
nor U8084 (N_8084,N_7431,N_6567);
or U8085 (N_8085,N_7433,N_6281);
nor U8086 (N_8086,N_6471,N_7124);
and U8087 (N_8087,N_7456,N_6283);
nor U8088 (N_8088,N_6851,N_6972);
xnor U8089 (N_8089,N_7121,N_6965);
or U8090 (N_8090,N_7401,N_7405);
and U8091 (N_8091,N_7191,N_6470);
and U8092 (N_8092,N_6693,N_7218);
nand U8093 (N_8093,N_7226,N_7409);
nor U8094 (N_8094,N_6973,N_7453);
nand U8095 (N_8095,N_6277,N_7033);
and U8096 (N_8096,N_6393,N_6899);
or U8097 (N_8097,N_7358,N_6926);
nor U8098 (N_8098,N_7277,N_7217);
or U8099 (N_8099,N_6931,N_7130);
or U8100 (N_8100,N_6532,N_7475);
nor U8101 (N_8101,N_7270,N_6321);
nand U8102 (N_8102,N_7299,N_7127);
and U8103 (N_8103,N_7068,N_7482);
nor U8104 (N_8104,N_6696,N_7463);
xor U8105 (N_8105,N_6793,N_7248);
and U8106 (N_8106,N_6954,N_6862);
xor U8107 (N_8107,N_6689,N_6261);
and U8108 (N_8108,N_6287,N_6673);
or U8109 (N_8109,N_6704,N_7177);
xor U8110 (N_8110,N_7351,N_6569);
or U8111 (N_8111,N_7231,N_6736);
xor U8112 (N_8112,N_6784,N_6754);
nor U8113 (N_8113,N_6838,N_6903);
and U8114 (N_8114,N_6661,N_7178);
nor U8115 (N_8115,N_7115,N_6407);
and U8116 (N_8116,N_6365,N_7333);
and U8117 (N_8117,N_6846,N_7224);
nand U8118 (N_8118,N_6839,N_6991);
and U8119 (N_8119,N_7166,N_7055);
nand U8120 (N_8120,N_6303,N_7266);
nand U8121 (N_8121,N_6445,N_7131);
nor U8122 (N_8122,N_6268,N_6741);
and U8123 (N_8123,N_6875,N_6448);
nand U8124 (N_8124,N_7371,N_6258);
and U8125 (N_8125,N_7444,N_6956);
nor U8126 (N_8126,N_7450,N_6501);
xor U8127 (N_8127,N_7047,N_6252);
nand U8128 (N_8128,N_7101,N_6626);
nand U8129 (N_8129,N_7150,N_6640);
or U8130 (N_8130,N_7292,N_6475);
and U8131 (N_8131,N_7346,N_6697);
nand U8132 (N_8132,N_6891,N_7258);
xnor U8133 (N_8133,N_7479,N_6565);
or U8134 (N_8134,N_6509,N_6255);
xnor U8135 (N_8135,N_6684,N_7433);
or U8136 (N_8136,N_7340,N_7017);
nor U8137 (N_8137,N_6731,N_6644);
xnor U8138 (N_8138,N_6600,N_7127);
and U8139 (N_8139,N_7109,N_6358);
or U8140 (N_8140,N_6906,N_7466);
nand U8141 (N_8141,N_7266,N_7491);
or U8142 (N_8142,N_7393,N_7151);
or U8143 (N_8143,N_6536,N_6870);
or U8144 (N_8144,N_6623,N_6526);
nor U8145 (N_8145,N_6432,N_7047);
nand U8146 (N_8146,N_6530,N_7249);
nor U8147 (N_8147,N_6292,N_7015);
or U8148 (N_8148,N_6679,N_6403);
nand U8149 (N_8149,N_6826,N_7163);
and U8150 (N_8150,N_6505,N_7158);
nor U8151 (N_8151,N_6320,N_6768);
nand U8152 (N_8152,N_6970,N_6757);
xnor U8153 (N_8153,N_7384,N_6449);
nor U8154 (N_8154,N_7064,N_6512);
and U8155 (N_8155,N_6275,N_7016);
nor U8156 (N_8156,N_7054,N_7469);
or U8157 (N_8157,N_7253,N_7037);
nor U8158 (N_8158,N_6760,N_6592);
nor U8159 (N_8159,N_6632,N_6585);
nand U8160 (N_8160,N_7218,N_6993);
nor U8161 (N_8161,N_6305,N_7196);
xnor U8162 (N_8162,N_6824,N_7342);
and U8163 (N_8163,N_6889,N_6339);
nor U8164 (N_8164,N_6327,N_6677);
xor U8165 (N_8165,N_7117,N_7024);
and U8166 (N_8166,N_6552,N_6341);
nand U8167 (N_8167,N_6477,N_6926);
nand U8168 (N_8168,N_7473,N_7291);
or U8169 (N_8169,N_7026,N_7065);
nor U8170 (N_8170,N_6861,N_6732);
or U8171 (N_8171,N_6325,N_6330);
nand U8172 (N_8172,N_6429,N_6981);
and U8173 (N_8173,N_7056,N_6920);
and U8174 (N_8174,N_7475,N_7207);
or U8175 (N_8175,N_7014,N_7220);
nand U8176 (N_8176,N_6806,N_6695);
nand U8177 (N_8177,N_7498,N_6950);
nor U8178 (N_8178,N_6747,N_7399);
xnor U8179 (N_8179,N_7128,N_6903);
nor U8180 (N_8180,N_6721,N_7361);
and U8181 (N_8181,N_6873,N_7052);
and U8182 (N_8182,N_7252,N_7441);
nand U8183 (N_8183,N_6734,N_6359);
xor U8184 (N_8184,N_7276,N_6713);
xor U8185 (N_8185,N_7434,N_6377);
xor U8186 (N_8186,N_6360,N_6783);
nor U8187 (N_8187,N_6536,N_7132);
nand U8188 (N_8188,N_6856,N_7116);
xnor U8189 (N_8189,N_6359,N_7288);
nand U8190 (N_8190,N_6303,N_7378);
xnor U8191 (N_8191,N_6589,N_7433);
and U8192 (N_8192,N_7084,N_7077);
nor U8193 (N_8193,N_6418,N_6910);
or U8194 (N_8194,N_7402,N_6734);
nand U8195 (N_8195,N_6631,N_6833);
nor U8196 (N_8196,N_6726,N_6521);
or U8197 (N_8197,N_6594,N_7416);
and U8198 (N_8198,N_6304,N_7402);
or U8199 (N_8199,N_7238,N_7454);
nor U8200 (N_8200,N_6602,N_7286);
xnor U8201 (N_8201,N_6695,N_7302);
nor U8202 (N_8202,N_7030,N_6439);
or U8203 (N_8203,N_6622,N_6274);
and U8204 (N_8204,N_6872,N_6623);
nor U8205 (N_8205,N_6485,N_6633);
nand U8206 (N_8206,N_6807,N_7458);
nor U8207 (N_8207,N_7455,N_6414);
and U8208 (N_8208,N_7122,N_6908);
or U8209 (N_8209,N_7312,N_6285);
and U8210 (N_8210,N_6262,N_6775);
nand U8211 (N_8211,N_6770,N_7027);
or U8212 (N_8212,N_7087,N_6929);
nand U8213 (N_8213,N_6512,N_7054);
and U8214 (N_8214,N_6584,N_6560);
and U8215 (N_8215,N_7412,N_6844);
nor U8216 (N_8216,N_6602,N_7138);
nand U8217 (N_8217,N_6629,N_7478);
xor U8218 (N_8218,N_6477,N_6797);
and U8219 (N_8219,N_6466,N_7002);
xnor U8220 (N_8220,N_7423,N_6389);
nor U8221 (N_8221,N_7095,N_6782);
and U8222 (N_8222,N_6566,N_6558);
and U8223 (N_8223,N_7166,N_7390);
and U8224 (N_8224,N_6654,N_7095);
nand U8225 (N_8225,N_7484,N_6940);
nand U8226 (N_8226,N_6302,N_7172);
or U8227 (N_8227,N_6499,N_6692);
nand U8228 (N_8228,N_6756,N_6477);
or U8229 (N_8229,N_6843,N_7139);
xor U8230 (N_8230,N_6571,N_6393);
nor U8231 (N_8231,N_7301,N_7255);
and U8232 (N_8232,N_7203,N_6741);
or U8233 (N_8233,N_6429,N_7114);
xnor U8234 (N_8234,N_6251,N_6551);
nor U8235 (N_8235,N_7203,N_7150);
or U8236 (N_8236,N_7242,N_7126);
nor U8237 (N_8237,N_6424,N_7311);
nand U8238 (N_8238,N_6321,N_6344);
and U8239 (N_8239,N_6306,N_6811);
xor U8240 (N_8240,N_6600,N_6679);
and U8241 (N_8241,N_7290,N_6325);
nor U8242 (N_8242,N_7093,N_6733);
nor U8243 (N_8243,N_6516,N_6492);
or U8244 (N_8244,N_7176,N_6413);
nand U8245 (N_8245,N_7339,N_6720);
and U8246 (N_8246,N_6994,N_6708);
and U8247 (N_8247,N_6712,N_6507);
nand U8248 (N_8248,N_7020,N_6820);
or U8249 (N_8249,N_7173,N_6379);
nand U8250 (N_8250,N_6417,N_6952);
or U8251 (N_8251,N_7449,N_6284);
and U8252 (N_8252,N_7133,N_6466);
and U8253 (N_8253,N_7177,N_6857);
nor U8254 (N_8254,N_6975,N_7012);
and U8255 (N_8255,N_6862,N_7454);
xnor U8256 (N_8256,N_6332,N_6264);
nor U8257 (N_8257,N_7224,N_6314);
xor U8258 (N_8258,N_6910,N_7313);
xor U8259 (N_8259,N_7353,N_7289);
xnor U8260 (N_8260,N_6423,N_7320);
or U8261 (N_8261,N_7402,N_6499);
xor U8262 (N_8262,N_7371,N_6787);
nand U8263 (N_8263,N_7165,N_7369);
nand U8264 (N_8264,N_7041,N_7199);
nand U8265 (N_8265,N_6955,N_6759);
xor U8266 (N_8266,N_6645,N_7368);
nor U8267 (N_8267,N_7372,N_6525);
nor U8268 (N_8268,N_7036,N_6310);
xor U8269 (N_8269,N_6619,N_6427);
nor U8270 (N_8270,N_7171,N_6991);
or U8271 (N_8271,N_6805,N_7365);
xnor U8272 (N_8272,N_6678,N_7481);
nor U8273 (N_8273,N_6526,N_6857);
nand U8274 (N_8274,N_6780,N_7329);
and U8275 (N_8275,N_6421,N_7345);
or U8276 (N_8276,N_6394,N_7499);
nor U8277 (N_8277,N_6353,N_7387);
or U8278 (N_8278,N_6602,N_6861);
nand U8279 (N_8279,N_6439,N_7307);
or U8280 (N_8280,N_6589,N_6302);
or U8281 (N_8281,N_7453,N_6791);
nand U8282 (N_8282,N_6279,N_7279);
and U8283 (N_8283,N_7084,N_7059);
and U8284 (N_8284,N_6723,N_7070);
xnor U8285 (N_8285,N_6698,N_6711);
and U8286 (N_8286,N_7096,N_6508);
nor U8287 (N_8287,N_6855,N_7140);
or U8288 (N_8288,N_6699,N_6961);
xor U8289 (N_8289,N_7288,N_7295);
nand U8290 (N_8290,N_6887,N_6403);
nor U8291 (N_8291,N_7283,N_7360);
or U8292 (N_8292,N_6952,N_7351);
and U8293 (N_8293,N_6799,N_6276);
nor U8294 (N_8294,N_7422,N_7370);
xor U8295 (N_8295,N_6662,N_6735);
nor U8296 (N_8296,N_7488,N_6815);
nor U8297 (N_8297,N_6593,N_7415);
or U8298 (N_8298,N_6994,N_7190);
nand U8299 (N_8299,N_6875,N_6422);
and U8300 (N_8300,N_7426,N_7140);
nand U8301 (N_8301,N_6826,N_6517);
or U8302 (N_8302,N_6554,N_7405);
nand U8303 (N_8303,N_6470,N_6358);
or U8304 (N_8304,N_7223,N_6600);
xor U8305 (N_8305,N_6257,N_6553);
nor U8306 (N_8306,N_7097,N_7480);
nor U8307 (N_8307,N_7202,N_6927);
nand U8308 (N_8308,N_6965,N_7083);
and U8309 (N_8309,N_6338,N_6713);
or U8310 (N_8310,N_7414,N_7434);
or U8311 (N_8311,N_6878,N_7414);
xnor U8312 (N_8312,N_7248,N_6315);
xor U8313 (N_8313,N_7446,N_7385);
or U8314 (N_8314,N_6592,N_6972);
nand U8315 (N_8315,N_7098,N_6361);
nor U8316 (N_8316,N_7413,N_7231);
nand U8317 (N_8317,N_6617,N_6806);
xnor U8318 (N_8318,N_6394,N_6471);
or U8319 (N_8319,N_6977,N_6998);
nand U8320 (N_8320,N_6521,N_6802);
or U8321 (N_8321,N_6422,N_6388);
or U8322 (N_8322,N_6726,N_6719);
and U8323 (N_8323,N_7129,N_7239);
xor U8324 (N_8324,N_7326,N_7005);
and U8325 (N_8325,N_6495,N_7326);
xor U8326 (N_8326,N_7384,N_6915);
xnor U8327 (N_8327,N_6426,N_6799);
and U8328 (N_8328,N_7437,N_7327);
nor U8329 (N_8329,N_6985,N_6755);
and U8330 (N_8330,N_6858,N_7190);
and U8331 (N_8331,N_7368,N_7192);
xor U8332 (N_8332,N_6612,N_7359);
or U8333 (N_8333,N_7169,N_7409);
xnor U8334 (N_8334,N_6622,N_6872);
and U8335 (N_8335,N_7467,N_6968);
nor U8336 (N_8336,N_6395,N_7311);
nand U8337 (N_8337,N_6698,N_6628);
xor U8338 (N_8338,N_6661,N_7358);
nand U8339 (N_8339,N_6692,N_7253);
and U8340 (N_8340,N_7386,N_7288);
or U8341 (N_8341,N_7213,N_7458);
and U8342 (N_8342,N_7230,N_6593);
or U8343 (N_8343,N_7296,N_6709);
nand U8344 (N_8344,N_7123,N_6504);
nand U8345 (N_8345,N_6284,N_7315);
nand U8346 (N_8346,N_7329,N_6964);
and U8347 (N_8347,N_7092,N_6956);
xor U8348 (N_8348,N_6273,N_6382);
xor U8349 (N_8349,N_6420,N_6501);
nor U8350 (N_8350,N_6299,N_6810);
nor U8351 (N_8351,N_7198,N_6770);
nand U8352 (N_8352,N_6864,N_6677);
xor U8353 (N_8353,N_6365,N_6659);
nand U8354 (N_8354,N_7122,N_7476);
and U8355 (N_8355,N_6344,N_6695);
or U8356 (N_8356,N_7165,N_7393);
and U8357 (N_8357,N_6288,N_7339);
or U8358 (N_8358,N_6828,N_7124);
nand U8359 (N_8359,N_6565,N_6970);
nand U8360 (N_8360,N_7122,N_6467);
nor U8361 (N_8361,N_6993,N_7286);
or U8362 (N_8362,N_6444,N_7242);
xor U8363 (N_8363,N_7175,N_6787);
nor U8364 (N_8364,N_7371,N_6577);
nor U8365 (N_8365,N_6417,N_6988);
xor U8366 (N_8366,N_7412,N_6857);
xor U8367 (N_8367,N_7124,N_6725);
or U8368 (N_8368,N_6302,N_6425);
or U8369 (N_8369,N_6666,N_6505);
nor U8370 (N_8370,N_6762,N_7164);
or U8371 (N_8371,N_6983,N_6930);
or U8372 (N_8372,N_6699,N_7185);
nand U8373 (N_8373,N_6803,N_6260);
nand U8374 (N_8374,N_6466,N_6798);
nor U8375 (N_8375,N_6835,N_7277);
or U8376 (N_8376,N_7271,N_7173);
xnor U8377 (N_8377,N_6639,N_6473);
xor U8378 (N_8378,N_6902,N_6586);
nand U8379 (N_8379,N_6891,N_6512);
and U8380 (N_8380,N_6928,N_6339);
and U8381 (N_8381,N_7330,N_6613);
nor U8382 (N_8382,N_6471,N_6903);
or U8383 (N_8383,N_7282,N_6461);
or U8384 (N_8384,N_7274,N_6497);
xnor U8385 (N_8385,N_7071,N_6808);
nor U8386 (N_8386,N_6551,N_7103);
or U8387 (N_8387,N_7387,N_6674);
or U8388 (N_8388,N_7112,N_6472);
nand U8389 (N_8389,N_7314,N_7380);
and U8390 (N_8390,N_7118,N_7440);
and U8391 (N_8391,N_6528,N_7010);
and U8392 (N_8392,N_6850,N_6756);
nor U8393 (N_8393,N_6979,N_6964);
or U8394 (N_8394,N_6452,N_6716);
and U8395 (N_8395,N_6490,N_7197);
and U8396 (N_8396,N_6903,N_6610);
and U8397 (N_8397,N_7310,N_6645);
nor U8398 (N_8398,N_6978,N_6731);
and U8399 (N_8399,N_6617,N_6746);
or U8400 (N_8400,N_6323,N_7345);
nand U8401 (N_8401,N_6398,N_6659);
nand U8402 (N_8402,N_6528,N_6991);
nor U8403 (N_8403,N_7101,N_6822);
nand U8404 (N_8404,N_6291,N_6661);
or U8405 (N_8405,N_6785,N_7150);
nand U8406 (N_8406,N_6393,N_6671);
nand U8407 (N_8407,N_6531,N_7200);
nor U8408 (N_8408,N_7142,N_7270);
nor U8409 (N_8409,N_6884,N_6547);
nor U8410 (N_8410,N_7070,N_6975);
nor U8411 (N_8411,N_6440,N_6646);
xnor U8412 (N_8412,N_7481,N_6885);
nor U8413 (N_8413,N_7391,N_7334);
xor U8414 (N_8414,N_7378,N_7496);
or U8415 (N_8415,N_6740,N_6571);
and U8416 (N_8416,N_7338,N_7457);
nand U8417 (N_8417,N_6545,N_6352);
nand U8418 (N_8418,N_6831,N_6649);
or U8419 (N_8419,N_7465,N_7374);
nand U8420 (N_8420,N_7003,N_6946);
nor U8421 (N_8421,N_6835,N_6856);
nand U8422 (N_8422,N_6388,N_6843);
nor U8423 (N_8423,N_6468,N_7027);
nand U8424 (N_8424,N_6537,N_6486);
nand U8425 (N_8425,N_6552,N_6306);
xnor U8426 (N_8426,N_7008,N_6717);
nand U8427 (N_8427,N_7290,N_7405);
and U8428 (N_8428,N_6875,N_6885);
or U8429 (N_8429,N_6365,N_7100);
nand U8430 (N_8430,N_7173,N_6562);
nor U8431 (N_8431,N_7205,N_6616);
and U8432 (N_8432,N_6340,N_7032);
and U8433 (N_8433,N_6811,N_6652);
nor U8434 (N_8434,N_6457,N_6568);
nor U8435 (N_8435,N_6366,N_6921);
and U8436 (N_8436,N_6499,N_6704);
and U8437 (N_8437,N_7092,N_6439);
and U8438 (N_8438,N_7490,N_6292);
xnor U8439 (N_8439,N_6550,N_7260);
nor U8440 (N_8440,N_6809,N_7129);
xor U8441 (N_8441,N_6832,N_7195);
and U8442 (N_8442,N_6666,N_6821);
nor U8443 (N_8443,N_7123,N_7289);
or U8444 (N_8444,N_7188,N_7140);
or U8445 (N_8445,N_6851,N_7167);
xnor U8446 (N_8446,N_7479,N_7015);
nand U8447 (N_8447,N_6835,N_7160);
nand U8448 (N_8448,N_7120,N_7202);
nor U8449 (N_8449,N_7138,N_7370);
nand U8450 (N_8450,N_6692,N_6745);
nand U8451 (N_8451,N_6764,N_7361);
and U8452 (N_8452,N_6463,N_6524);
or U8453 (N_8453,N_6371,N_6331);
xor U8454 (N_8454,N_6755,N_6598);
or U8455 (N_8455,N_6426,N_6608);
nor U8456 (N_8456,N_6386,N_6708);
nand U8457 (N_8457,N_6338,N_7329);
nor U8458 (N_8458,N_6923,N_6393);
xnor U8459 (N_8459,N_6755,N_7309);
or U8460 (N_8460,N_6855,N_6329);
nor U8461 (N_8461,N_6456,N_7397);
nand U8462 (N_8462,N_7024,N_6611);
nor U8463 (N_8463,N_7259,N_7409);
nor U8464 (N_8464,N_6275,N_6927);
and U8465 (N_8465,N_6737,N_6835);
xnor U8466 (N_8466,N_7485,N_6667);
nor U8467 (N_8467,N_7473,N_6668);
xor U8468 (N_8468,N_6630,N_7264);
nand U8469 (N_8469,N_6680,N_6397);
nand U8470 (N_8470,N_7336,N_7318);
nand U8471 (N_8471,N_7419,N_7435);
or U8472 (N_8472,N_6667,N_6719);
xnor U8473 (N_8473,N_6269,N_7370);
or U8474 (N_8474,N_6546,N_6620);
and U8475 (N_8475,N_6829,N_6566);
xor U8476 (N_8476,N_7218,N_6794);
nand U8477 (N_8477,N_6837,N_6625);
xnor U8478 (N_8478,N_6594,N_6711);
nor U8479 (N_8479,N_6416,N_7008);
nand U8480 (N_8480,N_6464,N_6969);
or U8481 (N_8481,N_6431,N_6912);
nand U8482 (N_8482,N_6353,N_6653);
or U8483 (N_8483,N_6885,N_7360);
nor U8484 (N_8484,N_7370,N_6416);
and U8485 (N_8485,N_7252,N_7331);
and U8486 (N_8486,N_6250,N_6251);
nor U8487 (N_8487,N_6682,N_7051);
or U8488 (N_8488,N_6289,N_6342);
xor U8489 (N_8489,N_7344,N_7462);
or U8490 (N_8490,N_6290,N_7357);
xnor U8491 (N_8491,N_7448,N_6712);
xnor U8492 (N_8492,N_6266,N_7251);
and U8493 (N_8493,N_7029,N_6289);
nor U8494 (N_8494,N_6657,N_6601);
xor U8495 (N_8495,N_6948,N_7386);
or U8496 (N_8496,N_7122,N_6847);
or U8497 (N_8497,N_6512,N_7396);
or U8498 (N_8498,N_7021,N_6448);
nor U8499 (N_8499,N_7181,N_7309);
nand U8500 (N_8500,N_6751,N_6900);
xnor U8501 (N_8501,N_7176,N_6972);
and U8502 (N_8502,N_6398,N_7397);
nor U8503 (N_8503,N_6677,N_6529);
and U8504 (N_8504,N_7426,N_6378);
nor U8505 (N_8505,N_6643,N_6403);
nand U8506 (N_8506,N_7161,N_7377);
or U8507 (N_8507,N_6824,N_6788);
nor U8508 (N_8508,N_7238,N_7461);
nand U8509 (N_8509,N_6561,N_6536);
or U8510 (N_8510,N_6472,N_7418);
nand U8511 (N_8511,N_6629,N_7445);
or U8512 (N_8512,N_6756,N_7276);
or U8513 (N_8513,N_7400,N_6325);
nor U8514 (N_8514,N_6984,N_6842);
and U8515 (N_8515,N_6474,N_6343);
nor U8516 (N_8516,N_6731,N_7413);
or U8517 (N_8517,N_7416,N_6640);
nand U8518 (N_8518,N_7107,N_7029);
or U8519 (N_8519,N_7132,N_7052);
xnor U8520 (N_8520,N_7081,N_7261);
nor U8521 (N_8521,N_6370,N_6757);
nand U8522 (N_8522,N_6372,N_6841);
xor U8523 (N_8523,N_7077,N_6766);
and U8524 (N_8524,N_7064,N_6966);
or U8525 (N_8525,N_6527,N_6475);
nand U8526 (N_8526,N_7453,N_7073);
and U8527 (N_8527,N_7356,N_6500);
or U8528 (N_8528,N_7475,N_6952);
or U8529 (N_8529,N_6834,N_7046);
nor U8530 (N_8530,N_6793,N_6470);
nand U8531 (N_8531,N_6505,N_6947);
nor U8532 (N_8532,N_6284,N_6341);
and U8533 (N_8533,N_7389,N_7094);
nand U8534 (N_8534,N_6497,N_7128);
nand U8535 (N_8535,N_6742,N_6800);
and U8536 (N_8536,N_7086,N_7398);
or U8537 (N_8537,N_6542,N_6654);
and U8538 (N_8538,N_6381,N_6987);
or U8539 (N_8539,N_6707,N_7355);
or U8540 (N_8540,N_6477,N_6538);
nor U8541 (N_8541,N_7075,N_7395);
nor U8542 (N_8542,N_7132,N_6678);
nand U8543 (N_8543,N_6755,N_7146);
nand U8544 (N_8544,N_6537,N_6730);
nand U8545 (N_8545,N_7115,N_7053);
or U8546 (N_8546,N_6982,N_6560);
and U8547 (N_8547,N_6706,N_7172);
xnor U8548 (N_8548,N_7448,N_7181);
nor U8549 (N_8549,N_6807,N_7119);
nor U8550 (N_8550,N_6527,N_6664);
nand U8551 (N_8551,N_6625,N_7197);
xor U8552 (N_8552,N_7315,N_7492);
xnor U8553 (N_8553,N_6426,N_7422);
and U8554 (N_8554,N_6998,N_6695);
nor U8555 (N_8555,N_6756,N_7280);
nand U8556 (N_8556,N_7274,N_6584);
nand U8557 (N_8557,N_7018,N_7473);
nor U8558 (N_8558,N_6718,N_6304);
and U8559 (N_8559,N_6327,N_6337);
and U8560 (N_8560,N_6754,N_6587);
nor U8561 (N_8561,N_7053,N_6981);
xor U8562 (N_8562,N_6682,N_6681);
xnor U8563 (N_8563,N_6355,N_6947);
xnor U8564 (N_8564,N_6314,N_6960);
or U8565 (N_8565,N_6638,N_6881);
nor U8566 (N_8566,N_6830,N_6648);
and U8567 (N_8567,N_7163,N_6476);
nand U8568 (N_8568,N_6667,N_7097);
nor U8569 (N_8569,N_7049,N_6581);
nor U8570 (N_8570,N_7224,N_6598);
nor U8571 (N_8571,N_6588,N_6616);
xnor U8572 (N_8572,N_6330,N_7082);
xnor U8573 (N_8573,N_6473,N_6382);
nand U8574 (N_8574,N_6753,N_6649);
nor U8575 (N_8575,N_7359,N_6494);
and U8576 (N_8576,N_6589,N_6379);
nand U8577 (N_8577,N_7001,N_6982);
nand U8578 (N_8578,N_7349,N_6797);
nand U8579 (N_8579,N_6408,N_6327);
or U8580 (N_8580,N_7294,N_7221);
nand U8581 (N_8581,N_7390,N_6264);
xor U8582 (N_8582,N_6672,N_6534);
nand U8583 (N_8583,N_7210,N_6984);
nand U8584 (N_8584,N_7103,N_7454);
xnor U8585 (N_8585,N_6652,N_6855);
xnor U8586 (N_8586,N_6633,N_6574);
or U8587 (N_8587,N_7084,N_6506);
xor U8588 (N_8588,N_6713,N_7405);
and U8589 (N_8589,N_6518,N_7086);
and U8590 (N_8590,N_6289,N_7036);
xnor U8591 (N_8591,N_6476,N_6526);
nand U8592 (N_8592,N_6452,N_6714);
and U8593 (N_8593,N_6749,N_7081);
nand U8594 (N_8594,N_6661,N_7361);
xnor U8595 (N_8595,N_6989,N_7278);
nor U8596 (N_8596,N_6305,N_6386);
xor U8597 (N_8597,N_6515,N_7172);
nand U8598 (N_8598,N_6606,N_7270);
and U8599 (N_8599,N_6844,N_6343);
nand U8600 (N_8600,N_6703,N_6840);
and U8601 (N_8601,N_7307,N_7055);
nor U8602 (N_8602,N_7474,N_7494);
xnor U8603 (N_8603,N_6573,N_7487);
and U8604 (N_8604,N_6838,N_6497);
and U8605 (N_8605,N_7146,N_7323);
nand U8606 (N_8606,N_7294,N_6317);
and U8607 (N_8607,N_6873,N_6886);
nand U8608 (N_8608,N_6946,N_6593);
xor U8609 (N_8609,N_6381,N_7147);
xor U8610 (N_8610,N_6886,N_7050);
xnor U8611 (N_8611,N_7293,N_7066);
xor U8612 (N_8612,N_6938,N_6828);
xnor U8613 (N_8613,N_6728,N_7495);
and U8614 (N_8614,N_7451,N_6618);
xnor U8615 (N_8615,N_6488,N_7189);
nand U8616 (N_8616,N_6859,N_6436);
xor U8617 (N_8617,N_6835,N_6436);
nor U8618 (N_8618,N_7168,N_7057);
xor U8619 (N_8619,N_6960,N_7177);
nor U8620 (N_8620,N_6736,N_7146);
nand U8621 (N_8621,N_6647,N_6839);
or U8622 (N_8622,N_6482,N_7055);
or U8623 (N_8623,N_6968,N_7291);
and U8624 (N_8624,N_6855,N_6883);
or U8625 (N_8625,N_6573,N_6945);
nand U8626 (N_8626,N_7181,N_6730);
xor U8627 (N_8627,N_6858,N_6454);
nor U8628 (N_8628,N_6855,N_7319);
or U8629 (N_8629,N_6428,N_6371);
or U8630 (N_8630,N_6332,N_6929);
nor U8631 (N_8631,N_7110,N_6983);
nor U8632 (N_8632,N_7061,N_6313);
xor U8633 (N_8633,N_6891,N_7032);
and U8634 (N_8634,N_7274,N_7393);
nor U8635 (N_8635,N_7029,N_7229);
xnor U8636 (N_8636,N_7044,N_6595);
or U8637 (N_8637,N_6901,N_7482);
nand U8638 (N_8638,N_7019,N_7263);
xnor U8639 (N_8639,N_6629,N_6692);
nand U8640 (N_8640,N_7043,N_6614);
or U8641 (N_8641,N_7082,N_6593);
and U8642 (N_8642,N_6748,N_6780);
nand U8643 (N_8643,N_7042,N_6414);
and U8644 (N_8644,N_6604,N_6257);
and U8645 (N_8645,N_7378,N_6876);
xor U8646 (N_8646,N_7061,N_6546);
nor U8647 (N_8647,N_7023,N_6315);
nor U8648 (N_8648,N_6924,N_6630);
nand U8649 (N_8649,N_7143,N_6950);
nor U8650 (N_8650,N_7130,N_7434);
or U8651 (N_8651,N_7409,N_7037);
nor U8652 (N_8652,N_6551,N_7267);
nand U8653 (N_8653,N_6492,N_6728);
xnor U8654 (N_8654,N_7445,N_7404);
nand U8655 (N_8655,N_7098,N_6857);
and U8656 (N_8656,N_6303,N_7281);
nor U8657 (N_8657,N_6938,N_6285);
nand U8658 (N_8658,N_7258,N_6710);
or U8659 (N_8659,N_7460,N_6381);
xnor U8660 (N_8660,N_6934,N_7306);
xor U8661 (N_8661,N_6592,N_6340);
nand U8662 (N_8662,N_6548,N_6915);
or U8663 (N_8663,N_7379,N_6358);
nor U8664 (N_8664,N_6308,N_7285);
and U8665 (N_8665,N_7202,N_6645);
or U8666 (N_8666,N_6358,N_6989);
xnor U8667 (N_8667,N_7242,N_7320);
nand U8668 (N_8668,N_6914,N_7335);
nand U8669 (N_8669,N_6466,N_7351);
nand U8670 (N_8670,N_6623,N_6902);
nor U8671 (N_8671,N_6603,N_7090);
or U8672 (N_8672,N_6334,N_7462);
nor U8673 (N_8673,N_7469,N_7148);
or U8674 (N_8674,N_7369,N_7391);
or U8675 (N_8675,N_7116,N_6972);
and U8676 (N_8676,N_6973,N_7358);
and U8677 (N_8677,N_6253,N_6609);
xor U8678 (N_8678,N_7453,N_7117);
or U8679 (N_8679,N_7398,N_6344);
xor U8680 (N_8680,N_6404,N_7011);
and U8681 (N_8681,N_6921,N_7412);
or U8682 (N_8682,N_7378,N_6730);
nor U8683 (N_8683,N_7492,N_6730);
nand U8684 (N_8684,N_7053,N_7346);
or U8685 (N_8685,N_6438,N_6889);
nand U8686 (N_8686,N_6994,N_7394);
xnor U8687 (N_8687,N_6714,N_6367);
and U8688 (N_8688,N_6589,N_6999);
nand U8689 (N_8689,N_7179,N_6327);
nor U8690 (N_8690,N_7157,N_6945);
nor U8691 (N_8691,N_6494,N_6740);
or U8692 (N_8692,N_7196,N_6869);
or U8693 (N_8693,N_6327,N_7256);
or U8694 (N_8694,N_6965,N_6688);
and U8695 (N_8695,N_7228,N_6937);
nor U8696 (N_8696,N_6425,N_7067);
and U8697 (N_8697,N_6441,N_7015);
and U8698 (N_8698,N_6260,N_7218);
xnor U8699 (N_8699,N_7472,N_6726);
or U8700 (N_8700,N_7328,N_7256);
nand U8701 (N_8701,N_7227,N_6800);
or U8702 (N_8702,N_6394,N_6379);
or U8703 (N_8703,N_7205,N_7110);
xor U8704 (N_8704,N_7455,N_7048);
or U8705 (N_8705,N_7324,N_6792);
and U8706 (N_8706,N_6300,N_7312);
xor U8707 (N_8707,N_7352,N_7109);
nand U8708 (N_8708,N_6328,N_6368);
nor U8709 (N_8709,N_6307,N_6788);
nand U8710 (N_8710,N_6680,N_6774);
and U8711 (N_8711,N_6577,N_6824);
xnor U8712 (N_8712,N_7136,N_6906);
nor U8713 (N_8713,N_6893,N_7461);
nor U8714 (N_8714,N_6541,N_7057);
xnor U8715 (N_8715,N_7010,N_7054);
nor U8716 (N_8716,N_7435,N_6388);
nand U8717 (N_8717,N_6576,N_6432);
nor U8718 (N_8718,N_7071,N_6342);
xor U8719 (N_8719,N_7191,N_7016);
nor U8720 (N_8720,N_6368,N_6464);
nand U8721 (N_8721,N_7429,N_7267);
and U8722 (N_8722,N_7268,N_6957);
nor U8723 (N_8723,N_7082,N_7258);
xnor U8724 (N_8724,N_6512,N_7248);
and U8725 (N_8725,N_6848,N_7205);
or U8726 (N_8726,N_7434,N_7243);
xor U8727 (N_8727,N_6983,N_7008);
or U8728 (N_8728,N_6317,N_6726);
xor U8729 (N_8729,N_6963,N_6350);
xor U8730 (N_8730,N_6917,N_7360);
xor U8731 (N_8731,N_7424,N_7271);
xnor U8732 (N_8732,N_6689,N_7391);
nor U8733 (N_8733,N_6595,N_6381);
nor U8734 (N_8734,N_6505,N_6338);
nand U8735 (N_8735,N_7454,N_6576);
or U8736 (N_8736,N_6734,N_7235);
nor U8737 (N_8737,N_7214,N_6550);
xnor U8738 (N_8738,N_6650,N_7077);
and U8739 (N_8739,N_7362,N_6917);
nand U8740 (N_8740,N_7413,N_6268);
nand U8741 (N_8741,N_7003,N_7032);
xor U8742 (N_8742,N_7363,N_7269);
and U8743 (N_8743,N_6318,N_6751);
nand U8744 (N_8744,N_6981,N_7122);
nand U8745 (N_8745,N_7252,N_7081);
or U8746 (N_8746,N_6526,N_6830);
nor U8747 (N_8747,N_6917,N_6496);
or U8748 (N_8748,N_6617,N_7436);
nor U8749 (N_8749,N_6866,N_6573);
nand U8750 (N_8750,N_7891,N_7855);
nand U8751 (N_8751,N_8559,N_8451);
nand U8752 (N_8752,N_8716,N_7978);
nor U8753 (N_8753,N_8332,N_8733);
and U8754 (N_8754,N_7769,N_7544);
and U8755 (N_8755,N_8167,N_8527);
xnor U8756 (N_8756,N_7902,N_8729);
nor U8757 (N_8757,N_7812,N_8277);
or U8758 (N_8758,N_7672,N_8508);
and U8759 (N_8759,N_8554,N_8408);
xnor U8760 (N_8760,N_7934,N_8747);
nand U8761 (N_8761,N_7677,N_7922);
nand U8762 (N_8762,N_7614,N_8295);
or U8763 (N_8763,N_7543,N_8197);
xnor U8764 (N_8764,N_8123,N_8124);
or U8765 (N_8765,N_8454,N_8149);
or U8766 (N_8766,N_8352,N_8158);
or U8767 (N_8767,N_7625,N_8669);
and U8768 (N_8768,N_7719,N_8534);
or U8769 (N_8769,N_8067,N_7715);
xnor U8770 (N_8770,N_7987,N_7951);
nor U8771 (N_8771,N_8676,N_8170);
xnor U8772 (N_8772,N_7691,N_8009);
nand U8773 (N_8773,N_8431,N_8252);
or U8774 (N_8774,N_7565,N_7519);
or U8775 (N_8775,N_8380,N_7775);
nor U8776 (N_8776,N_7973,N_7985);
nand U8777 (N_8777,N_8414,N_7605);
or U8778 (N_8778,N_7774,N_7911);
nor U8779 (N_8779,N_7853,N_8594);
or U8780 (N_8780,N_8569,N_8028);
nor U8781 (N_8781,N_7604,N_8052);
and U8782 (N_8782,N_8563,N_8137);
nand U8783 (N_8783,N_8708,N_7959);
nor U8784 (N_8784,N_7773,N_7521);
and U8785 (N_8785,N_8440,N_8481);
nor U8786 (N_8786,N_8522,N_8572);
xnor U8787 (N_8787,N_7953,N_8697);
or U8788 (N_8788,N_7727,N_8281);
nand U8789 (N_8789,N_8696,N_7764);
xnor U8790 (N_8790,N_8429,N_8686);
xor U8791 (N_8791,N_8501,N_8063);
nand U8792 (N_8792,N_8417,N_8469);
nand U8793 (N_8793,N_7696,N_7548);
or U8794 (N_8794,N_8141,N_7776);
xnor U8795 (N_8795,N_8248,N_8358);
xor U8796 (N_8796,N_8085,N_8573);
xnor U8797 (N_8797,N_8433,N_8427);
xor U8798 (N_8798,N_8256,N_8404);
nor U8799 (N_8799,N_7708,N_7753);
and U8800 (N_8800,N_7811,N_7836);
or U8801 (N_8801,N_7539,N_8166);
xnor U8802 (N_8802,N_8341,N_8153);
nand U8803 (N_8803,N_8233,N_7659);
and U8804 (N_8804,N_8560,N_7700);
nor U8805 (N_8805,N_7921,N_8331);
xor U8806 (N_8806,N_7806,N_8025);
nand U8807 (N_8807,N_8577,N_8343);
xor U8808 (N_8808,N_7502,N_7829);
or U8809 (N_8809,N_7743,N_8714);
or U8810 (N_8810,N_8033,N_8693);
nand U8811 (N_8811,N_8611,N_8654);
nand U8812 (N_8812,N_8656,N_8583);
or U8813 (N_8813,N_8486,N_7901);
and U8814 (N_8814,N_8467,N_8407);
nor U8815 (N_8815,N_8627,N_8743);
xor U8816 (N_8816,N_7818,N_7622);
nand U8817 (N_8817,N_7856,N_8249);
nand U8818 (N_8818,N_8398,N_8212);
or U8819 (N_8819,N_8621,N_8095);
or U8820 (N_8820,N_7916,N_7630);
xor U8821 (N_8821,N_8000,N_8388);
and U8822 (N_8822,N_7796,N_8318);
xnor U8823 (N_8823,N_7827,N_7724);
or U8824 (N_8824,N_8078,N_8495);
nand U8825 (N_8825,N_8024,N_8293);
and U8826 (N_8826,N_7688,N_7522);
nor U8827 (N_8827,N_8551,N_8307);
xnor U8828 (N_8828,N_8425,N_7706);
xnor U8829 (N_8829,N_8634,N_8529);
or U8830 (N_8830,N_8374,N_8647);
or U8831 (N_8831,N_8242,N_8199);
xnor U8832 (N_8832,N_7643,N_7562);
nand U8833 (N_8833,N_8557,N_7616);
nor U8834 (N_8834,N_8313,N_7613);
or U8835 (N_8835,N_7640,N_7955);
or U8836 (N_8836,N_8315,N_8150);
nor U8837 (N_8837,N_7816,N_7506);
nand U8838 (N_8838,N_7866,N_8683);
nor U8839 (N_8839,N_7761,N_7908);
xor U8840 (N_8840,N_8644,N_8228);
and U8841 (N_8841,N_7992,N_7592);
and U8842 (N_8842,N_8173,N_8505);
xnor U8843 (N_8843,N_7892,N_7756);
and U8844 (N_8844,N_7500,N_7576);
and U8845 (N_8845,N_7567,N_8416);
nand U8846 (N_8846,N_8449,N_8533);
or U8847 (N_8847,N_8204,N_7697);
or U8848 (N_8848,N_7745,N_7781);
nand U8849 (N_8849,N_7684,N_7555);
and U8850 (N_8850,N_7644,N_7982);
and U8851 (N_8851,N_7792,N_7772);
or U8852 (N_8852,N_8734,N_7648);
nor U8853 (N_8853,N_8462,N_8579);
nor U8854 (N_8854,N_7633,N_7787);
or U8855 (N_8855,N_7854,N_7950);
nor U8856 (N_8856,N_8597,N_8118);
or U8857 (N_8857,N_7651,N_8463);
and U8858 (N_8858,N_7516,N_8311);
and U8859 (N_8859,N_8194,N_8283);
nand U8860 (N_8860,N_8446,N_8606);
nor U8861 (N_8861,N_7802,N_7600);
nor U8862 (N_8862,N_8324,N_8059);
xnor U8863 (N_8863,N_8221,N_8532);
nand U8864 (N_8864,N_7879,N_8452);
nor U8865 (N_8865,N_8112,N_8537);
and U8866 (N_8866,N_8596,N_8081);
and U8867 (N_8867,N_7733,N_7662);
or U8868 (N_8868,N_7569,N_8623);
nand U8869 (N_8869,N_7947,N_7874);
or U8870 (N_8870,N_8668,N_8581);
and U8871 (N_8871,N_7606,N_8222);
nor U8872 (N_8872,N_8397,N_8671);
and U8873 (N_8873,N_7841,N_8005);
nand U8874 (N_8874,N_8031,N_8284);
or U8875 (N_8875,N_8710,N_8163);
xnor U8876 (N_8876,N_7797,N_8631);
nand U8877 (N_8877,N_8565,N_7608);
nand U8878 (N_8878,N_8265,N_7877);
or U8879 (N_8879,N_7546,N_7586);
nor U8880 (N_8880,N_7615,N_7564);
and U8881 (N_8881,N_8741,N_8436);
and U8882 (N_8882,N_8615,N_8500);
xnor U8883 (N_8883,N_8737,N_8072);
xnor U8884 (N_8884,N_8518,N_8680);
nor U8885 (N_8885,N_8234,N_8480);
nor U8886 (N_8886,N_8069,N_7810);
nor U8887 (N_8887,N_7822,N_7735);
or U8888 (N_8888,N_7863,N_8202);
nor U8889 (N_8889,N_8323,N_8703);
and U8890 (N_8890,N_8539,N_7514);
and U8891 (N_8891,N_8147,N_8273);
nor U8892 (N_8892,N_7925,N_8278);
nor U8893 (N_8893,N_8238,N_7517);
xor U8894 (N_8894,N_8092,N_7634);
xnor U8895 (N_8895,N_8642,N_7558);
or U8896 (N_8896,N_8218,N_7656);
nand U8897 (N_8897,N_7794,N_7572);
nand U8898 (N_8898,N_8459,N_8291);
xnor U8899 (N_8899,N_7723,N_7886);
or U8900 (N_8900,N_8070,N_8400);
nor U8901 (N_8901,N_7831,N_8098);
nand U8902 (N_8902,N_8638,N_7748);
nand U8903 (N_8903,N_8333,N_8041);
and U8904 (N_8904,N_7965,N_8019);
nand U8905 (N_8905,N_8509,N_8636);
or U8906 (N_8906,N_8251,N_8205);
xnor U8907 (N_8907,N_8077,N_8213);
and U8908 (N_8908,N_8006,N_8447);
and U8909 (N_8909,N_8113,N_8259);
xnor U8910 (N_8910,N_8326,N_7559);
nor U8911 (N_8911,N_8571,N_7524);
or U8912 (N_8912,N_8330,N_8175);
and U8913 (N_8913,N_8237,N_8717);
and U8914 (N_8914,N_8575,N_8740);
nor U8915 (N_8915,N_8336,N_7563);
nand U8916 (N_8916,N_7515,N_8392);
xor U8917 (N_8917,N_7749,N_8356);
or U8918 (N_8918,N_7693,N_7807);
nor U8919 (N_8919,N_7638,N_8582);
nand U8920 (N_8920,N_8017,N_8187);
nand U8921 (N_8921,N_7872,N_7588);
nand U8922 (N_8922,N_8125,N_8513);
or U8923 (N_8923,N_8189,N_7971);
nor U8924 (N_8924,N_8567,N_7976);
nand U8925 (N_8925,N_8719,N_7612);
and U8926 (N_8926,N_8292,N_7858);
or U8927 (N_8927,N_8727,N_8007);
nor U8928 (N_8928,N_8306,N_8612);
nand U8929 (N_8929,N_8626,N_7601);
nand U8930 (N_8930,N_7805,N_8297);
nor U8931 (N_8931,N_8183,N_7652);
and U8932 (N_8932,N_8035,N_7547);
xor U8933 (N_8933,N_8337,N_8453);
xor U8934 (N_8934,N_8588,N_8060);
xnor U8935 (N_8935,N_7607,N_7714);
and U8936 (N_8936,N_8104,N_7939);
nor U8937 (N_8937,N_8203,N_8082);
nand U8938 (N_8938,N_7997,N_7636);
and U8939 (N_8939,N_7870,N_7956);
xor U8940 (N_8940,N_7979,N_8004);
xnor U8941 (N_8941,N_8715,N_8186);
and U8942 (N_8942,N_8381,N_8528);
xor U8943 (N_8943,N_8029,N_8748);
and U8944 (N_8944,N_8121,N_8196);
xnor U8945 (N_8945,N_7918,N_8541);
nand U8946 (N_8946,N_7848,N_8584);
nand U8947 (N_8947,N_8239,N_8725);
xnor U8948 (N_8948,N_7549,N_8286);
nor U8949 (N_8949,N_8516,N_8409);
or U8950 (N_8950,N_8523,N_8426);
xnor U8951 (N_8951,N_7669,N_7712);
and U8952 (N_8952,N_7532,N_8100);
xnor U8953 (N_8953,N_7860,N_7815);
and U8954 (N_8954,N_8240,N_8678);
xnor U8955 (N_8955,N_8110,N_7575);
nor U8956 (N_8956,N_8576,N_8386);
and U8957 (N_8957,N_7868,N_7778);
and U8958 (N_8958,N_7660,N_7977);
and U8959 (N_8959,N_8371,N_8483);
nand U8960 (N_8960,N_8488,N_7574);
nand U8961 (N_8961,N_8164,N_7611);
and U8962 (N_8962,N_8322,N_7758);
xor U8963 (N_8963,N_7535,N_8109);
and U8964 (N_8964,N_8329,N_7573);
nor U8965 (N_8965,N_8227,N_8701);
nand U8966 (N_8966,N_8672,N_8485);
and U8967 (N_8967,N_8266,N_7541);
nor U8968 (N_8968,N_8171,N_7690);
and U8969 (N_8969,N_7851,N_8650);
nor U8970 (N_8970,N_8319,N_7647);
nor U8971 (N_8971,N_8617,N_8271);
xnor U8972 (N_8972,N_7629,N_7751);
xnor U8973 (N_8973,N_8587,N_7603);
nand U8974 (N_8974,N_8340,N_8264);
xor U8975 (N_8975,N_7504,N_8015);
or U8976 (N_8976,N_8134,N_8514);
nand U8977 (N_8977,N_7523,N_8401);
and U8978 (N_8978,N_7779,N_7752);
xor U8979 (N_8979,N_8413,N_7533);
nand U8980 (N_8980,N_8062,N_8664);
nor U8981 (N_8981,N_8720,N_7801);
and U8982 (N_8982,N_8742,N_8154);
and U8983 (N_8983,N_8687,N_7846);
or U8984 (N_8984,N_8673,N_7942);
and U8985 (N_8985,N_8010,N_8298);
nand U8986 (N_8986,N_7940,N_8314);
and U8987 (N_8987,N_7917,N_7954);
nand U8988 (N_8988,N_7898,N_8721);
xnor U8989 (N_8989,N_8128,N_8335);
xnor U8990 (N_8990,N_7814,N_8032);
or U8991 (N_8991,N_7710,N_7895);
or U8992 (N_8992,N_8039,N_7963);
and U8993 (N_8993,N_8261,N_7845);
nand U8994 (N_8994,N_7980,N_8531);
xor U8995 (N_8995,N_7993,N_7763);
and U8996 (N_8996,N_7596,N_7676);
xnor U8997 (N_8997,N_8622,N_8290);
and U8998 (N_8998,N_8465,N_8544);
nor U8999 (N_8999,N_8043,N_7518);
nand U9000 (N_9000,N_8294,N_7771);
and U9001 (N_9001,N_8670,N_8040);
and U9002 (N_9002,N_8267,N_8609);
nand U9003 (N_9003,N_8198,N_7580);
xor U9004 (N_9004,N_7821,N_8061);
or U9005 (N_9005,N_7553,N_7933);
nand U9006 (N_9006,N_8373,N_8350);
xnor U9007 (N_9007,N_7692,N_7582);
xor U9008 (N_9008,N_8012,N_8225);
nand U9009 (N_9009,N_7840,N_7526);
xor U9010 (N_9010,N_7881,N_7850);
and U9011 (N_9011,N_8188,N_8589);
nand U9012 (N_9012,N_8393,N_8084);
or U9013 (N_9013,N_7678,N_7674);
nand U9014 (N_9014,N_8207,N_8677);
nand U9015 (N_9015,N_7508,N_8530);
nand U9016 (N_9016,N_7958,N_8605);
xor U9017 (N_9017,N_7791,N_8558);
and U9018 (N_9018,N_8482,N_7974);
nand U9019 (N_9019,N_8151,N_8176);
or U9020 (N_9020,N_8106,N_8599);
or U9021 (N_9021,N_8466,N_8030);
xnor U9022 (N_9022,N_8192,N_7928);
xor U9023 (N_9023,N_7875,N_8247);
xnor U9024 (N_9024,N_8450,N_8111);
xor U9025 (N_9025,N_7646,N_8200);
or U9026 (N_9026,N_7713,N_8232);
xor U9027 (N_9027,N_8155,N_8364);
nor U9028 (N_9028,N_8243,N_7903);
xor U9029 (N_9029,N_8246,N_8633);
nand U9030 (N_9030,N_8550,N_8214);
xor U9031 (N_9031,N_8684,N_8138);
nor U9032 (N_9032,N_8014,N_7534);
or U9033 (N_9033,N_8008,N_8377);
nor U9034 (N_9034,N_7949,N_7914);
xor U9035 (N_9035,N_7730,N_7687);
and U9036 (N_9036,N_8279,N_8328);
and U9037 (N_9037,N_8499,N_8280);
or U9038 (N_9038,N_7961,N_7788);
and U9039 (N_9039,N_8478,N_7780);
and U9040 (N_9040,N_7593,N_8665);
nand U9041 (N_9041,N_8068,N_7577);
xnor U9042 (N_9042,N_8658,N_8660);
nand U9043 (N_9043,N_8091,N_7755);
or U9044 (N_9044,N_7832,N_8735);
xnor U9045 (N_9045,N_7941,N_8075);
nor U9046 (N_9046,N_8722,N_8224);
xor U9047 (N_9047,N_8662,N_7990);
nor U9048 (N_9048,N_7888,N_8384);
xnor U9049 (N_9049,N_7599,N_7824);
nand U9050 (N_9050,N_7768,N_8476);
nor U9051 (N_9051,N_8058,N_7889);
nor U9052 (N_9052,N_8434,N_8287);
xnor U9053 (N_9053,N_8245,N_7740);
xnor U9054 (N_9054,N_8178,N_7790);
nor U9055 (N_9055,N_7587,N_8073);
or U9056 (N_9056,N_8339,N_7808);
and U9057 (N_9057,N_7915,N_8026);
nand U9058 (N_9058,N_8455,N_8094);
nor U9059 (N_9059,N_7671,N_8510);
or U9060 (N_9060,N_7762,N_8169);
and U9061 (N_9061,N_7847,N_7994);
or U9062 (N_9062,N_8056,N_8540);
and U9063 (N_9063,N_8274,N_8439);
and U9064 (N_9064,N_8553,N_8651);
nand U9065 (N_9065,N_8105,N_8027);
and U9066 (N_9066,N_8087,N_8564);
or U9067 (N_9067,N_7828,N_8076);
or U9068 (N_9068,N_8132,N_8182);
nand U9069 (N_9069,N_8270,N_8342);
or U9070 (N_9070,N_8399,N_8088);
nand U9071 (N_9071,N_8632,N_7938);
xnor U9072 (N_9072,N_8037,N_7972);
nor U9073 (N_9073,N_8115,N_8420);
nor U9074 (N_9074,N_7507,N_8497);
nor U9075 (N_9075,N_8174,N_8362);
nand U9076 (N_9076,N_7884,N_7864);
nor U9077 (N_9077,N_8231,N_8304);
nand U9078 (N_9078,N_8473,N_8548);
xnor U9079 (N_9079,N_8457,N_7770);
xnor U9080 (N_9080,N_7571,N_8679);
xnor U9081 (N_9081,N_7658,N_8526);
xor U9082 (N_9082,N_8161,N_7991);
or U9083 (N_9083,N_7667,N_8487);
xnor U9084 (N_9084,N_8236,N_7509);
or U9085 (N_9085,N_7741,N_8604);
nand U9086 (N_9086,N_7621,N_7531);
nand U9087 (N_9087,N_8625,N_7682);
and U9088 (N_9088,N_8148,N_8681);
xnor U9089 (N_9089,N_8699,N_7584);
nand U9090 (N_9090,N_8368,N_7641);
xnor U9091 (N_9091,N_8502,N_8593);
nand U9092 (N_9092,N_8591,N_8731);
nor U9093 (N_9093,N_7635,N_8360);
nor U9094 (N_9094,N_7725,N_7679);
xnor U9095 (N_9095,N_7746,N_8160);
and U9096 (N_9096,N_8327,N_8299);
nor U9097 (N_9097,N_7578,N_8445);
nor U9098 (N_9098,N_7817,N_7893);
and U9099 (N_9099,N_8272,N_8181);
nand U9100 (N_9100,N_8618,N_7750);
or U9101 (N_9101,N_8129,N_7654);
or U9102 (N_9102,N_8536,N_8269);
nor U9103 (N_9103,N_8394,N_8566);
xor U9104 (N_9104,N_8020,N_7556);
xnor U9105 (N_9105,N_7887,N_8241);
or U9106 (N_9106,N_8405,N_8641);
nor U9107 (N_9107,N_7861,N_8570);
nor U9108 (N_9108,N_8157,N_7919);
xnor U9109 (N_9109,N_8317,N_8285);
or U9110 (N_9110,N_7785,N_7989);
xnor U9111 (N_9111,N_7595,N_8744);
and U9112 (N_9112,N_7876,N_8613);
and U9113 (N_9113,N_8107,N_8038);
xor U9114 (N_9114,N_8300,N_8139);
xnor U9115 (N_9115,N_8220,N_7686);
nor U9116 (N_9116,N_8001,N_7830);
and U9117 (N_9117,N_7698,N_8490);
or U9118 (N_9118,N_7826,N_7589);
and U9119 (N_9119,N_8695,N_8345);
and U9120 (N_9120,N_7632,N_8011);
xnor U9121 (N_9121,N_7655,N_7561);
xor U9122 (N_9122,N_8496,N_7598);
xor U9123 (N_9123,N_8726,N_8143);
and U9124 (N_9124,N_8718,N_7804);
xor U9125 (N_9125,N_7800,N_7786);
or U9126 (N_9126,N_8739,N_8474);
nand U9127 (N_9127,N_8675,N_8250);
nand U9128 (N_9128,N_8504,N_7560);
nor U9129 (N_9129,N_8301,N_8296);
nor U9130 (N_9130,N_7890,N_8309);
nand U9131 (N_9131,N_7957,N_8355);
xor U9132 (N_9132,N_8666,N_8549);
nand U9133 (N_9133,N_8140,N_7783);
or U9134 (N_9134,N_7721,N_8461);
nand U9135 (N_9135,N_7967,N_7583);
and U9136 (N_9136,N_7711,N_8723);
nand U9137 (N_9137,N_7799,N_7964);
xor U9138 (N_9138,N_8630,N_8555);
and U9139 (N_9139,N_8177,N_7552);
and U9140 (N_9140,N_7623,N_7873);
xor U9141 (N_9141,N_7869,N_8136);
or U9142 (N_9142,N_8464,N_8172);
xnor U9143 (N_9143,N_7594,N_7747);
and U9144 (N_9144,N_7505,N_7906);
xor U9145 (N_9145,N_8066,N_7525);
xnor U9146 (N_9146,N_7536,N_7722);
and U9147 (N_9147,N_8353,N_8489);
and U9148 (N_9148,N_8580,N_7610);
xor U9149 (N_9149,N_8263,N_8209);
or U9150 (N_9150,N_7842,N_8262);
or U9151 (N_9151,N_7639,N_7728);
nor U9152 (N_9152,N_7789,N_7975);
xnor U9153 (N_9153,N_7726,N_8217);
and U9154 (N_9154,N_8344,N_8367);
nor U9155 (N_9155,N_8053,N_8180);
nand U9156 (N_9156,N_8506,N_7618);
or U9157 (N_9157,N_7766,N_8044);
and U9158 (N_9158,N_8620,N_8477);
nor U9159 (N_9159,N_7899,N_8437);
xor U9160 (N_9160,N_7694,N_8702);
or U9161 (N_9161,N_8403,N_7645);
nor U9162 (N_9162,N_8728,N_8391);
nand U9163 (N_9163,N_7701,N_7717);
xor U9164 (N_9164,N_7585,N_8211);
nand U9165 (N_9165,N_8458,N_7540);
nor U9166 (N_9166,N_8730,N_7983);
xnor U9167 (N_9167,N_8159,N_8711);
and U9168 (N_9168,N_8491,N_8479);
nand U9169 (N_9169,N_8685,N_8448);
nor U9170 (N_9170,N_8484,N_7910);
or U9171 (N_9171,N_8097,N_7670);
and U9172 (N_9172,N_8275,N_8302);
xor U9173 (N_9173,N_8648,N_8162);
nand U9174 (N_9174,N_8357,N_8258);
xnor U9175 (N_9175,N_7704,N_8472);
nand U9176 (N_9176,N_8691,N_7912);
nor U9177 (N_9177,N_8524,N_8661);
and U9178 (N_9178,N_8460,N_8131);
or U9179 (N_9179,N_7920,N_8372);
and U9180 (N_9180,N_8168,N_7952);
or U9181 (N_9181,N_8470,N_8430);
nor U9182 (N_9182,N_8276,N_8046);
or U9183 (N_9183,N_7936,N_7685);
nand U9184 (N_9184,N_8108,N_8190);
nand U9185 (N_9185,N_8216,N_8375);
and U9186 (N_9186,N_7720,N_7909);
and U9187 (N_9187,N_7649,N_8546);
or U9188 (N_9188,N_7627,N_7765);
and U9189 (N_9189,N_8542,N_8674);
xor U9190 (N_9190,N_8260,N_7865);
xnor U9191 (N_9191,N_7838,N_8325);
nand U9192 (N_9192,N_8152,N_8568);
and U9193 (N_9193,N_8303,N_7885);
and U9194 (N_9194,N_8607,N_8421);
nand U9195 (N_9195,N_7538,N_8629);
or U9196 (N_9196,N_8179,N_8036);
and U9197 (N_9197,N_8640,N_8378);
nor U9198 (N_9198,N_7568,N_8086);
xnor U9199 (N_9199,N_7716,N_8688);
xnor U9200 (N_9200,N_8709,N_8268);
or U9201 (N_9201,N_8419,N_8146);
nand U9202 (N_9202,N_8122,N_7849);
xor U9203 (N_9203,N_7737,N_7834);
xor U9204 (N_9204,N_8244,N_7839);
or U9205 (N_9205,N_8689,N_8657);
xnor U9206 (N_9206,N_7981,N_8119);
and U9207 (N_9207,N_7661,N_8387);
nand U9208 (N_9208,N_8590,N_8308);
and U9209 (N_9209,N_7637,N_7904);
xor U9210 (N_9210,N_8736,N_8601);
and U9211 (N_9211,N_7732,N_8493);
xnor U9212 (N_9212,N_8637,N_7597);
nor U9213 (N_9213,N_7935,N_7907);
and U9214 (N_9214,N_8423,N_8142);
nor U9215 (N_9215,N_7683,N_8643);
or U9216 (N_9216,N_7798,N_8208);
nor U9217 (N_9217,N_7510,N_7759);
xnor U9218 (N_9218,N_7527,N_8096);
or U9219 (N_9219,N_8114,N_8229);
nor U9220 (N_9220,N_8706,N_8468);
nand U9221 (N_9221,N_7859,N_8402);
xnor U9222 (N_9222,N_8471,N_8385);
or U9223 (N_9223,N_7566,N_8586);
nor U9224 (N_9224,N_8713,N_7996);
or U9225 (N_9225,N_8351,N_7545);
or U9226 (N_9226,N_8515,N_8707);
nor U9227 (N_9227,N_8120,N_8080);
nor U9228 (N_9228,N_8561,N_7742);
and U9229 (N_9229,N_8503,N_7988);
nand U9230 (N_9230,N_8406,N_7905);
and U9231 (N_9231,N_8545,N_8210);
nand U9232 (N_9232,N_7689,N_7664);
or U9233 (N_9233,N_8428,N_8363);
or U9234 (N_9234,N_8646,N_7998);
and U9235 (N_9235,N_8346,N_8395);
or U9236 (N_9236,N_7946,N_7550);
or U9237 (N_9237,N_7878,N_8021);
and U9238 (N_9238,N_8042,N_8156);
and U9239 (N_9239,N_8538,N_8547);
or U9240 (N_9240,N_8045,N_7666);
or U9241 (N_9241,N_8071,N_8127);
xnor U9242 (N_9242,N_8389,N_8525);
or U9243 (N_9243,N_8144,N_7937);
nor U9244 (N_9244,N_8635,N_8475);
or U9245 (N_9245,N_7926,N_7882);
or U9246 (N_9246,N_7777,N_8432);
and U9247 (N_9247,N_8418,N_7995);
xnor U9248 (N_9248,N_8610,N_8047);
and U9249 (N_9249,N_8282,N_8102);
and U9250 (N_9250,N_8376,N_8034);
or U9251 (N_9251,N_8507,N_8435);
xnor U9252 (N_9252,N_7628,N_7653);
nor U9253 (N_9253,N_7966,N_7813);
nand U9254 (N_9254,N_8690,N_7948);
or U9255 (N_9255,N_8145,N_8441);
nor U9256 (N_9256,N_8126,N_7668);
xnor U9257 (N_9257,N_7512,N_8226);
or U9258 (N_9258,N_8365,N_7913);
nand U9259 (N_9259,N_7537,N_7984);
nor U9260 (N_9260,N_8321,N_7729);
and U9261 (N_9261,N_8382,N_8379);
or U9262 (N_9262,N_8424,N_8746);
and U9263 (N_9263,N_8090,N_7579);
and U9264 (N_9264,N_8517,N_8598);
or U9265 (N_9265,N_7739,N_7871);
or U9266 (N_9266,N_8370,N_8492);
or U9267 (N_9267,N_8065,N_8608);
nor U9268 (N_9268,N_8732,N_8624);
or U9269 (N_9269,N_8659,N_8185);
xor U9270 (N_9270,N_8003,N_8602);
nand U9271 (N_9271,N_8018,N_8639);
nor U9272 (N_9272,N_7825,N_8512);
xor U9273 (N_9273,N_7520,N_7897);
xnor U9274 (N_9274,N_8055,N_8519);
nand U9275 (N_9275,N_8117,N_8556);
and U9276 (N_9276,N_8521,N_8002);
xor U9277 (N_9277,N_7923,N_7896);
xnor U9278 (N_9278,N_7960,N_8592);
or U9279 (N_9279,N_8700,N_8694);
nor U9280 (N_9280,N_8064,N_8682);
nand U9281 (N_9281,N_8438,N_8595);
nor U9282 (N_9282,N_8745,N_8585);
nor U9283 (N_9283,N_7757,N_8645);
xnor U9284 (N_9284,N_7820,N_8103);
xor U9285 (N_9285,N_7620,N_7570);
and U9286 (N_9286,N_8422,N_8444);
xor U9287 (N_9287,N_7894,N_8412);
and U9288 (N_9288,N_8184,N_7782);
and U9289 (N_9289,N_8655,N_8215);
nor U9290 (N_9290,N_7703,N_8079);
nand U9291 (N_9291,N_8411,N_8348);
or U9292 (N_9292,N_8235,N_8443);
and U9293 (N_9293,N_8649,N_7930);
or U9294 (N_9294,N_8410,N_8652);
nand U9295 (N_9295,N_8738,N_7675);
or U9296 (N_9296,N_8057,N_8206);
or U9297 (N_9297,N_7843,N_7803);
and U9298 (N_9298,N_7650,N_7734);
nor U9299 (N_9299,N_8049,N_7695);
nor U9300 (N_9300,N_8361,N_8135);
nand U9301 (N_9301,N_7986,N_8334);
nor U9302 (N_9302,N_7900,N_8383);
xnor U9303 (N_9303,N_7528,N_8316);
or U9304 (N_9304,N_8578,N_8089);
and U9305 (N_9305,N_8165,N_7927);
nor U9306 (N_9306,N_8498,N_8312);
or U9307 (N_9307,N_7680,N_7699);
and U9308 (N_9308,N_7793,N_7591);
nand U9309 (N_9309,N_8013,N_7970);
and U9310 (N_9310,N_8050,N_8305);
and U9311 (N_9311,N_7945,N_8442);
nor U9312 (N_9312,N_7809,N_8494);
nor U9313 (N_9313,N_7844,N_7823);
or U9314 (N_9314,N_7924,N_8619);
or U9315 (N_9315,N_8653,N_7932);
nand U9316 (N_9316,N_8191,N_7529);
xor U9317 (N_9317,N_7663,N_8320);
and U9318 (N_9318,N_7619,N_7511);
and U9319 (N_9319,N_8101,N_7857);
or U9320 (N_9320,N_8366,N_8705);
nor U9321 (N_9321,N_7880,N_8133);
nand U9322 (N_9322,N_7929,N_7681);
nor U9323 (N_9323,N_7657,N_7617);
xor U9324 (N_9324,N_8354,N_7883);
nand U9325 (N_9325,N_7968,N_8253);
nand U9326 (N_9326,N_8016,N_8562);
and U9327 (N_9327,N_8201,N_8223);
and U9328 (N_9328,N_7501,N_7931);
nand U9329 (N_9329,N_8347,N_7551);
and U9330 (N_9330,N_7731,N_7513);
or U9331 (N_9331,N_8099,N_8023);
or U9332 (N_9332,N_7702,N_8415);
or U9333 (N_9333,N_8288,N_8692);
nand U9334 (N_9334,N_8616,N_8116);
or U9335 (N_9335,N_8255,N_8054);
xnor U9336 (N_9336,N_7754,N_7705);
nor U9337 (N_9337,N_7784,N_8535);
xnor U9338 (N_9338,N_8195,N_7642);
and U9339 (N_9339,N_8359,N_7835);
and U9340 (N_9340,N_7795,N_8396);
nor U9341 (N_9341,N_7837,N_7709);
or U9342 (N_9342,N_7944,N_7624);
xnor U9343 (N_9343,N_8724,N_7581);
and U9344 (N_9344,N_7833,N_7962);
and U9345 (N_9345,N_8628,N_8219);
and U9346 (N_9346,N_7760,N_8193);
nor U9347 (N_9347,N_8022,N_8051);
or U9348 (N_9348,N_7718,N_7673);
nor U9349 (N_9349,N_8310,N_8704);
or U9350 (N_9350,N_7503,N_7542);
or U9351 (N_9351,N_8614,N_7736);
nand U9352 (N_9352,N_8130,N_8338);
and U9353 (N_9353,N_8230,N_8520);
xnor U9354 (N_9354,N_8289,N_7631);
and U9355 (N_9355,N_8712,N_8074);
nand U9356 (N_9356,N_8093,N_8552);
xor U9357 (N_9357,N_8667,N_7602);
and U9358 (N_9358,N_8369,N_8698);
nor U9359 (N_9359,N_8349,N_7852);
nor U9360 (N_9360,N_8749,N_8083);
and U9361 (N_9361,N_7969,N_8257);
and U9362 (N_9362,N_7590,N_7557);
xnor U9363 (N_9363,N_8600,N_7767);
nand U9364 (N_9364,N_8390,N_7530);
or U9365 (N_9365,N_8603,N_8663);
or U9366 (N_9366,N_7943,N_8574);
and U9367 (N_9367,N_7819,N_8254);
or U9368 (N_9368,N_7626,N_7744);
nand U9369 (N_9369,N_7609,N_8456);
and U9370 (N_9370,N_7999,N_7665);
xnor U9371 (N_9371,N_8048,N_8511);
xor U9372 (N_9372,N_7738,N_8543);
and U9373 (N_9373,N_7867,N_7707);
xor U9374 (N_9374,N_7862,N_7554);
nand U9375 (N_9375,N_8087,N_8312);
and U9376 (N_9376,N_8386,N_7836);
nor U9377 (N_9377,N_8278,N_8443);
or U9378 (N_9378,N_8194,N_7501);
and U9379 (N_9379,N_8654,N_7505);
or U9380 (N_9380,N_7515,N_7817);
xnor U9381 (N_9381,N_8280,N_8445);
or U9382 (N_9382,N_8309,N_8305);
and U9383 (N_9383,N_8323,N_7934);
nor U9384 (N_9384,N_7682,N_7637);
nand U9385 (N_9385,N_8088,N_8546);
and U9386 (N_9386,N_8554,N_7564);
xor U9387 (N_9387,N_8188,N_7977);
or U9388 (N_9388,N_8348,N_7517);
or U9389 (N_9389,N_7581,N_8549);
nor U9390 (N_9390,N_8117,N_8580);
nor U9391 (N_9391,N_7754,N_8694);
nor U9392 (N_9392,N_8273,N_8350);
nand U9393 (N_9393,N_8492,N_8305);
xor U9394 (N_9394,N_8746,N_8193);
xnor U9395 (N_9395,N_8512,N_8597);
or U9396 (N_9396,N_8520,N_8529);
or U9397 (N_9397,N_8495,N_7621);
nor U9398 (N_9398,N_7595,N_8419);
xor U9399 (N_9399,N_8594,N_8290);
nor U9400 (N_9400,N_7857,N_7989);
and U9401 (N_9401,N_7862,N_8246);
nand U9402 (N_9402,N_8327,N_8607);
nand U9403 (N_9403,N_8115,N_7862);
nand U9404 (N_9404,N_7921,N_8244);
xnor U9405 (N_9405,N_7730,N_7685);
nand U9406 (N_9406,N_8448,N_7591);
or U9407 (N_9407,N_7954,N_8344);
or U9408 (N_9408,N_8107,N_7535);
and U9409 (N_9409,N_7833,N_7879);
xnor U9410 (N_9410,N_8209,N_7943);
nand U9411 (N_9411,N_7704,N_8431);
or U9412 (N_9412,N_8597,N_8247);
nor U9413 (N_9413,N_8194,N_8609);
nor U9414 (N_9414,N_8703,N_7986);
and U9415 (N_9415,N_8150,N_8245);
and U9416 (N_9416,N_8564,N_8025);
nand U9417 (N_9417,N_7878,N_8329);
or U9418 (N_9418,N_8419,N_8258);
and U9419 (N_9419,N_8102,N_7978);
and U9420 (N_9420,N_8396,N_8169);
or U9421 (N_9421,N_8278,N_8635);
and U9422 (N_9422,N_8694,N_7968);
nor U9423 (N_9423,N_7552,N_7997);
nor U9424 (N_9424,N_8284,N_8381);
or U9425 (N_9425,N_7682,N_8030);
nand U9426 (N_9426,N_8174,N_8250);
nor U9427 (N_9427,N_7834,N_7687);
nand U9428 (N_9428,N_8267,N_8742);
nor U9429 (N_9429,N_8557,N_8058);
xnor U9430 (N_9430,N_8025,N_8395);
or U9431 (N_9431,N_8150,N_8273);
xnor U9432 (N_9432,N_8158,N_7925);
nand U9433 (N_9433,N_7776,N_7796);
nand U9434 (N_9434,N_8190,N_8737);
nor U9435 (N_9435,N_7544,N_8347);
xnor U9436 (N_9436,N_7695,N_8410);
nand U9437 (N_9437,N_8314,N_7607);
nand U9438 (N_9438,N_7795,N_7559);
or U9439 (N_9439,N_7781,N_7847);
or U9440 (N_9440,N_8551,N_8082);
nand U9441 (N_9441,N_7637,N_7784);
xnor U9442 (N_9442,N_8621,N_7896);
nand U9443 (N_9443,N_8586,N_8214);
xor U9444 (N_9444,N_7978,N_7619);
or U9445 (N_9445,N_7828,N_7607);
nand U9446 (N_9446,N_7534,N_8248);
xnor U9447 (N_9447,N_8438,N_8181);
xnor U9448 (N_9448,N_7920,N_8061);
and U9449 (N_9449,N_7794,N_8160);
xor U9450 (N_9450,N_8193,N_8298);
xor U9451 (N_9451,N_7869,N_8594);
nand U9452 (N_9452,N_8648,N_8275);
and U9453 (N_9453,N_7992,N_8749);
xor U9454 (N_9454,N_8625,N_8657);
xnor U9455 (N_9455,N_8137,N_8520);
nor U9456 (N_9456,N_8263,N_7614);
nor U9457 (N_9457,N_8548,N_8258);
and U9458 (N_9458,N_8276,N_8035);
xnor U9459 (N_9459,N_8043,N_7955);
or U9460 (N_9460,N_8370,N_7879);
xor U9461 (N_9461,N_8531,N_8391);
xnor U9462 (N_9462,N_8745,N_8352);
and U9463 (N_9463,N_7874,N_7784);
and U9464 (N_9464,N_7702,N_8124);
and U9465 (N_9465,N_7785,N_7570);
xor U9466 (N_9466,N_8573,N_8231);
or U9467 (N_9467,N_8512,N_8229);
or U9468 (N_9468,N_8236,N_8683);
or U9469 (N_9469,N_7839,N_8565);
nand U9470 (N_9470,N_7893,N_8124);
xor U9471 (N_9471,N_8555,N_8649);
and U9472 (N_9472,N_8202,N_7750);
and U9473 (N_9473,N_8333,N_8393);
and U9474 (N_9474,N_8293,N_8391);
nor U9475 (N_9475,N_8319,N_7664);
xnor U9476 (N_9476,N_8386,N_8519);
or U9477 (N_9477,N_8155,N_7758);
and U9478 (N_9478,N_8613,N_7622);
xnor U9479 (N_9479,N_7767,N_8042);
or U9480 (N_9480,N_8105,N_7757);
nor U9481 (N_9481,N_7827,N_7907);
nor U9482 (N_9482,N_7650,N_7747);
nor U9483 (N_9483,N_7538,N_8377);
nand U9484 (N_9484,N_8384,N_8647);
and U9485 (N_9485,N_8026,N_7702);
xor U9486 (N_9486,N_8054,N_7690);
or U9487 (N_9487,N_7911,N_8747);
nand U9488 (N_9488,N_8563,N_8597);
nand U9489 (N_9489,N_8016,N_7692);
xor U9490 (N_9490,N_8513,N_7825);
or U9491 (N_9491,N_8360,N_8542);
xor U9492 (N_9492,N_7876,N_8402);
xor U9493 (N_9493,N_8504,N_7918);
nand U9494 (N_9494,N_8150,N_8238);
nand U9495 (N_9495,N_7985,N_8507);
and U9496 (N_9496,N_8579,N_8615);
and U9497 (N_9497,N_7872,N_8545);
nor U9498 (N_9498,N_8589,N_8153);
nand U9499 (N_9499,N_8207,N_7835);
nand U9500 (N_9500,N_8663,N_7790);
and U9501 (N_9501,N_7771,N_7890);
xnor U9502 (N_9502,N_8549,N_8052);
nand U9503 (N_9503,N_8192,N_8283);
nand U9504 (N_9504,N_8436,N_7841);
or U9505 (N_9505,N_8333,N_7919);
or U9506 (N_9506,N_8561,N_7636);
nand U9507 (N_9507,N_8222,N_8687);
nor U9508 (N_9508,N_8478,N_7828);
or U9509 (N_9509,N_8305,N_8746);
or U9510 (N_9510,N_8010,N_8041);
or U9511 (N_9511,N_8475,N_8651);
and U9512 (N_9512,N_7511,N_7538);
nor U9513 (N_9513,N_7635,N_8712);
and U9514 (N_9514,N_7729,N_7688);
xnor U9515 (N_9515,N_8326,N_7671);
nand U9516 (N_9516,N_7892,N_8536);
nor U9517 (N_9517,N_8456,N_8025);
nor U9518 (N_9518,N_8073,N_8574);
nor U9519 (N_9519,N_8327,N_8700);
nor U9520 (N_9520,N_8311,N_8665);
nor U9521 (N_9521,N_8275,N_8337);
or U9522 (N_9522,N_7655,N_8697);
or U9523 (N_9523,N_8584,N_8477);
nor U9524 (N_9524,N_7535,N_7618);
nor U9525 (N_9525,N_7794,N_8226);
xor U9526 (N_9526,N_8742,N_7837);
nand U9527 (N_9527,N_8551,N_8141);
or U9528 (N_9528,N_7937,N_7543);
nor U9529 (N_9529,N_7682,N_8147);
nand U9530 (N_9530,N_8724,N_7794);
nand U9531 (N_9531,N_7741,N_8222);
xor U9532 (N_9532,N_8231,N_8195);
nand U9533 (N_9533,N_8139,N_8208);
nor U9534 (N_9534,N_7933,N_7543);
nand U9535 (N_9535,N_8307,N_7739);
nand U9536 (N_9536,N_7616,N_7669);
xnor U9537 (N_9537,N_8365,N_8060);
nand U9538 (N_9538,N_7524,N_8225);
nor U9539 (N_9539,N_8066,N_8370);
xnor U9540 (N_9540,N_7572,N_7639);
or U9541 (N_9541,N_7886,N_8644);
nand U9542 (N_9542,N_7805,N_7558);
nor U9543 (N_9543,N_8268,N_8021);
or U9544 (N_9544,N_7897,N_7671);
nand U9545 (N_9545,N_8040,N_7701);
nor U9546 (N_9546,N_7941,N_7549);
nand U9547 (N_9547,N_8223,N_8096);
xnor U9548 (N_9548,N_8673,N_8399);
xnor U9549 (N_9549,N_8367,N_7546);
nand U9550 (N_9550,N_7824,N_7901);
nor U9551 (N_9551,N_8579,N_8327);
and U9552 (N_9552,N_8730,N_8289);
and U9553 (N_9553,N_7684,N_8295);
or U9554 (N_9554,N_8392,N_7783);
or U9555 (N_9555,N_7612,N_7555);
xor U9556 (N_9556,N_7915,N_8004);
nor U9557 (N_9557,N_7660,N_7784);
xor U9558 (N_9558,N_7742,N_8021);
or U9559 (N_9559,N_8648,N_8084);
nor U9560 (N_9560,N_8057,N_8211);
nand U9561 (N_9561,N_7809,N_8728);
or U9562 (N_9562,N_8499,N_7781);
nand U9563 (N_9563,N_8455,N_7921);
nor U9564 (N_9564,N_7693,N_8227);
or U9565 (N_9565,N_8522,N_7518);
and U9566 (N_9566,N_8501,N_8096);
nand U9567 (N_9567,N_8546,N_7849);
nand U9568 (N_9568,N_8458,N_8210);
xor U9569 (N_9569,N_7865,N_8558);
xor U9570 (N_9570,N_8538,N_8438);
xnor U9571 (N_9571,N_8473,N_8149);
nand U9572 (N_9572,N_8601,N_8191);
xor U9573 (N_9573,N_7699,N_8355);
nand U9574 (N_9574,N_8560,N_8701);
or U9575 (N_9575,N_8022,N_8372);
nand U9576 (N_9576,N_8746,N_7733);
and U9577 (N_9577,N_7885,N_8505);
and U9578 (N_9578,N_7863,N_7657);
xnor U9579 (N_9579,N_7942,N_7597);
nand U9580 (N_9580,N_7934,N_7518);
nand U9581 (N_9581,N_8321,N_8136);
nor U9582 (N_9582,N_8240,N_8439);
xnor U9583 (N_9583,N_7658,N_8552);
nand U9584 (N_9584,N_7649,N_8307);
or U9585 (N_9585,N_8424,N_8160);
nor U9586 (N_9586,N_8460,N_8740);
or U9587 (N_9587,N_7909,N_8614);
or U9588 (N_9588,N_8384,N_8143);
and U9589 (N_9589,N_8286,N_8250);
nand U9590 (N_9590,N_8069,N_7930);
and U9591 (N_9591,N_8339,N_7768);
nand U9592 (N_9592,N_8475,N_7588);
nor U9593 (N_9593,N_8510,N_7819);
nor U9594 (N_9594,N_7857,N_7860);
and U9595 (N_9595,N_7577,N_7636);
nand U9596 (N_9596,N_8581,N_7619);
xnor U9597 (N_9597,N_8207,N_7838);
xor U9598 (N_9598,N_7979,N_7867);
xnor U9599 (N_9599,N_8618,N_7603);
xor U9600 (N_9600,N_8493,N_7706);
xnor U9601 (N_9601,N_8667,N_8740);
nand U9602 (N_9602,N_7970,N_8068);
nand U9603 (N_9603,N_8456,N_7988);
nor U9604 (N_9604,N_8651,N_8278);
or U9605 (N_9605,N_7734,N_8437);
or U9606 (N_9606,N_7998,N_8233);
and U9607 (N_9607,N_8029,N_7900);
nand U9608 (N_9608,N_7653,N_7519);
xor U9609 (N_9609,N_7862,N_8426);
nand U9610 (N_9610,N_7655,N_8507);
xnor U9611 (N_9611,N_7728,N_8708);
nor U9612 (N_9612,N_8162,N_7802);
and U9613 (N_9613,N_8408,N_7728);
and U9614 (N_9614,N_8151,N_8205);
and U9615 (N_9615,N_7828,N_8110);
and U9616 (N_9616,N_7804,N_8161);
nor U9617 (N_9617,N_7648,N_7554);
xnor U9618 (N_9618,N_8135,N_8314);
nor U9619 (N_9619,N_8338,N_7624);
xnor U9620 (N_9620,N_8293,N_8249);
xnor U9621 (N_9621,N_8635,N_7863);
or U9622 (N_9622,N_7865,N_8726);
and U9623 (N_9623,N_8464,N_8404);
nor U9624 (N_9624,N_8721,N_7811);
nand U9625 (N_9625,N_8378,N_7760);
nor U9626 (N_9626,N_8146,N_7677);
xor U9627 (N_9627,N_7717,N_8578);
xnor U9628 (N_9628,N_8399,N_7712);
or U9629 (N_9629,N_7765,N_8424);
and U9630 (N_9630,N_8291,N_7547);
nand U9631 (N_9631,N_8550,N_8019);
nor U9632 (N_9632,N_7864,N_8303);
nor U9633 (N_9633,N_8117,N_8095);
nor U9634 (N_9634,N_8042,N_8115);
nor U9635 (N_9635,N_7613,N_7502);
nand U9636 (N_9636,N_8363,N_8511);
and U9637 (N_9637,N_7721,N_8045);
nand U9638 (N_9638,N_7771,N_7554);
nor U9639 (N_9639,N_7580,N_7718);
or U9640 (N_9640,N_7943,N_7839);
or U9641 (N_9641,N_7712,N_7869);
nand U9642 (N_9642,N_8265,N_7878);
and U9643 (N_9643,N_7807,N_7682);
xnor U9644 (N_9644,N_7752,N_8690);
xor U9645 (N_9645,N_7727,N_8601);
or U9646 (N_9646,N_8696,N_8381);
nor U9647 (N_9647,N_8375,N_7823);
or U9648 (N_9648,N_8242,N_7760);
or U9649 (N_9649,N_8709,N_8546);
nand U9650 (N_9650,N_8329,N_7630);
or U9651 (N_9651,N_8091,N_7642);
xor U9652 (N_9652,N_7955,N_8276);
xor U9653 (N_9653,N_8259,N_8553);
nor U9654 (N_9654,N_8288,N_7903);
nand U9655 (N_9655,N_8368,N_7798);
nand U9656 (N_9656,N_8080,N_7756);
nor U9657 (N_9657,N_8376,N_7794);
or U9658 (N_9658,N_8132,N_8303);
nand U9659 (N_9659,N_7802,N_7797);
nand U9660 (N_9660,N_7601,N_8274);
nor U9661 (N_9661,N_7645,N_7615);
xor U9662 (N_9662,N_7622,N_8699);
nor U9663 (N_9663,N_7825,N_8245);
nand U9664 (N_9664,N_8497,N_7964);
or U9665 (N_9665,N_8539,N_8011);
xnor U9666 (N_9666,N_7637,N_7583);
or U9667 (N_9667,N_8695,N_8747);
nor U9668 (N_9668,N_7860,N_8558);
or U9669 (N_9669,N_7738,N_8436);
xor U9670 (N_9670,N_8634,N_8650);
nor U9671 (N_9671,N_7871,N_8181);
or U9672 (N_9672,N_8336,N_8062);
nor U9673 (N_9673,N_7912,N_8102);
and U9674 (N_9674,N_8441,N_8063);
nor U9675 (N_9675,N_8712,N_8473);
or U9676 (N_9676,N_8675,N_8305);
nor U9677 (N_9677,N_8410,N_8329);
or U9678 (N_9678,N_8481,N_7922);
and U9679 (N_9679,N_7506,N_7991);
xor U9680 (N_9680,N_8653,N_8281);
or U9681 (N_9681,N_8063,N_7502);
or U9682 (N_9682,N_8207,N_7907);
and U9683 (N_9683,N_7653,N_8378);
nor U9684 (N_9684,N_7771,N_7757);
nand U9685 (N_9685,N_7552,N_7500);
nand U9686 (N_9686,N_7606,N_7695);
and U9687 (N_9687,N_7836,N_7503);
nor U9688 (N_9688,N_7677,N_8640);
xor U9689 (N_9689,N_7833,N_8188);
nor U9690 (N_9690,N_8108,N_8347);
nor U9691 (N_9691,N_8212,N_7640);
xor U9692 (N_9692,N_7884,N_8191);
xnor U9693 (N_9693,N_8566,N_8675);
or U9694 (N_9694,N_7944,N_8612);
nor U9695 (N_9695,N_8648,N_8332);
xnor U9696 (N_9696,N_8142,N_7789);
and U9697 (N_9697,N_8193,N_7635);
and U9698 (N_9698,N_7910,N_7873);
nand U9699 (N_9699,N_7908,N_7766);
and U9700 (N_9700,N_8654,N_8027);
nand U9701 (N_9701,N_8057,N_8462);
nand U9702 (N_9702,N_8279,N_8076);
nand U9703 (N_9703,N_8195,N_7719);
nor U9704 (N_9704,N_7729,N_8127);
xnor U9705 (N_9705,N_7951,N_7571);
nand U9706 (N_9706,N_7921,N_8310);
nor U9707 (N_9707,N_8330,N_7655);
and U9708 (N_9708,N_8075,N_8693);
nor U9709 (N_9709,N_7615,N_8314);
nand U9710 (N_9710,N_7843,N_8074);
or U9711 (N_9711,N_8105,N_7890);
nand U9712 (N_9712,N_7697,N_8117);
and U9713 (N_9713,N_8179,N_7704);
nand U9714 (N_9714,N_8255,N_7580);
nand U9715 (N_9715,N_8670,N_7926);
or U9716 (N_9716,N_8166,N_8694);
or U9717 (N_9717,N_8240,N_8117);
nand U9718 (N_9718,N_8533,N_7974);
nor U9719 (N_9719,N_8376,N_7805);
or U9720 (N_9720,N_8433,N_8308);
nor U9721 (N_9721,N_8389,N_8114);
nor U9722 (N_9722,N_8619,N_8095);
nand U9723 (N_9723,N_7910,N_8128);
or U9724 (N_9724,N_8678,N_8049);
and U9725 (N_9725,N_8058,N_7947);
xnor U9726 (N_9726,N_8007,N_7620);
nor U9727 (N_9727,N_7882,N_8586);
and U9728 (N_9728,N_7985,N_7794);
nand U9729 (N_9729,N_8302,N_7869);
xor U9730 (N_9730,N_7816,N_8535);
and U9731 (N_9731,N_8501,N_7591);
xnor U9732 (N_9732,N_7962,N_7674);
or U9733 (N_9733,N_8405,N_7698);
xnor U9734 (N_9734,N_7596,N_8524);
nand U9735 (N_9735,N_7687,N_7639);
or U9736 (N_9736,N_7885,N_7763);
nor U9737 (N_9737,N_8658,N_8499);
nand U9738 (N_9738,N_7912,N_8564);
or U9739 (N_9739,N_8573,N_7536);
nand U9740 (N_9740,N_8721,N_8668);
nand U9741 (N_9741,N_7958,N_8072);
or U9742 (N_9742,N_8488,N_7542);
nor U9743 (N_9743,N_7782,N_7604);
or U9744 (N_9744,N_7535,N_8194);
xor U9745 (N_9745,N_8272,N_8006);
or U9746 (N_9746,N_7561,N_8313);
nand U9747 (N_9747,N_7745,N_8051);
and U9748 (N_9748,N_8400,N_8474);
nand U9749 (N_9749,N_7633,N_7524);
xnor U9750 (N_9750,N_7771,N_8094);
xnor U9751 (N_9751,N_7954,N_8093);
nor U9752 (N_9752,N_8155,N_8443);
nor U9753 (N_9753,N_7736,N_7654);
or U9754 (N_9754,N_7876,N_8390);
or U9755 (N_9755,N_8454,N_7568);
nor U9756 (N_9756,N_8311,N_8206);
nand U9757 (N_9757,N_8576,N_7947);
nor U9758 (N_9758,N_8342,N_7522);
nand U9759 (N_9759,N_7947,N_7820);
nor U9760 (N_9760,N_8594,N_8186);
and U9761 (N_9761,N_7692,N_7872);
nor U9762 (N_9762,N_7644,N_7927);
or U9763 (N_9763,N_8715,N_8104);
and U9764 (N_9764,N_8243,N_8233);
nor U9765 (N_9765,N_8058,N_8745);
nand U9766 (N_9766,N_8026,N_8138);
and U9767 (N_9767,N_8360,N_7847);
nor U9768 (N_9768,N_8226,N_7686);
and U9769 (N_9769,N_7543,N_8191);
xor U9770 (N_9770,N_7508,N_7920);
and U9771 (N_9771,N_7880,N_7780);
and U9772 (N_9772,N_8567,N_7931);
nand U9773 (N_9773,N_7926,N_7502);
xnor U9774 (N_9774,N_7941,N_7700);
nor U9775 (N_9775,N_7864,N_8307);
and U9776 (N_9776,N_8328,N_7510);
and U9777 (N_9777,N_8217,N_8436);
nand U9778 (N_9778,N_7858,N_8335);
nor U9779 (N_9779,N_7507,N_8368);
and U9780 (N_9780,N_7835,N_7552);
and U9781 (N_9781,N_8189,N_7822);
xor U9782 (N_9782,N_8255,N_7538);
xnor U9783 (N_9783,N_7638,N_8748);
nand U9784 (N_9784,N_8213,N_7548);
nor U9785 (N_9785,N_7783,N_8476);
nor U9786 (N_9786,N_7766,N_8744);
nor U9787 (N_9787,N_8325,N_7523);
nand U9788 (N_9788,N_7685,N_7588);
xor U9789 (N_9789,N_8533,N_8064);
nand U9790 (N_9790,N_8442,N_8520);
or U9791 (N_9791,N_8060,N_7982);
and U9792 (N_9792,N_8314,N_8631);
nand U9793 (N_9793,N_8185,N_7904);
nor U9794 (N_9794,N_7887,N_7510);
nor U9795 (N_9795,N_8262,N_7722);
or U9796 (N_9796,N_8443,N_8358);
xnor U9797 (N_9797,N_8124,N_7671);
and U9798 (N_9798,N_8283,N_8346);
or U9799 (N_9799,N_8734,N_8421);
nand U9800 (N_9800,N_8031,N_7775);
or U9801 (N_9801,N_7515,N_8131);
nand U9802 (N_9802,N_7600,N_8309);
and U9803 (N_9803,N_8318,N_8633);
or U9804 (N_9804,N_7514,N_8424);
xnor U9805 (N_9805,N_7533,N_7676);
and U9806 (N_9806,N_8730,N_8526);
and U9807 (N_9807,N_7715,N_7523);
nand U9808 (N_9808,N_8149,N_8211);
nor U9809 (N_9809,N_8369,N_7835);
nor U9810 (N_9810,N_8276,N_7538);
or U9811 (N_9811,N_8275,N_8258);
and U9812 (N_9812,N_7559,N_7802);
nor U9813 (N_9813,N_7959,N_8354);
xor U9814 (N_9814,N_7594,N_8506);
and U9815 (N_9815,N_8558,N_8049);
nand U9816 (N_9816,N_8063,N_8144);
nor U9817 (N_9817,N_8159,N_7855);
xnor U9818 (N_9818,N_8460,N_7938);
nand U9819 (N_9819,N_8304,N_8638);
nor U9820 (N_9820,N_8499,N_8278);
and U9821 (N_9821,N_7927,N_7998);
xnor U9822 (N_9822,N_8107,N_8611);
xor U9823 (N_9823,N_8582,N_8713);
nor U9824 (N_9824,N_7747,N_7933);
nor U9825 (N_9825,N_8545,N_7776);
or U9826 (N_9826,N_8654,N_7970);
nand U9827 (N_9827,N_7702,N_8688);
or U9828 (N_9828,N_7567,N_7837);
nand U9829 (N_9829,N_7865,N_7811);
nand U9830 (N_9830,N_7923,N_7792);
nand U9831 (N_9831,N_8738,N_8573);
xnor U9832 (N_9832,N_8298,N_8465);
nor U9833 (N_9833,N_8324,N_8486);
nor U9834 (N_9834,N_8014,N_8432);
nand U9835 (N_9835,N_8093,N_8486);
xor U9836 (N_9836,N_8183,N_8505);
or U9837 (N_9837,N_7828,N_7718);
or U9838 (N_9838,N_8212,N_8413);
or U9839 (N_9839,N_8069,N_8718);
nand U9840 (N_9840,N_8480,N_8521);
or U9841 (N_9841,N_8391,N_8676);
and U9842 (N_9842,N_8508,N_8293);
nor U9843 (N_9843,N_8448,N_8392);
and U9844 (N_9844,N_8319,N_8570);
and U9845 (N_9845,N_8529,N_7701);
or U9846 (N_9846,N_8095,N_7712);
nor U9847 (N_9847,N_8415,N_8181);
xor U9848 (N_9848,N_8066,N_7582);
or U9849 (N_9849,N_7552,N_8493);
nor U9850 (N_9850,N_8185,N_7529);
xor U9851 (N_9851,N_8508,N_8078);
nor U9852 (N_9852,N_8037,N_8557);
nand U9853 (N_9853,N_8166,N_7914);
nor U9854 (N_9854,N_7566,N_7552);
nand U9855 (N_9855,N_8305,N_8662);
or U9856 (N_9856,N_8687,N_7507);
nor U9857 (N_9857,N_8003,N_7949);
xor U9858 (N_9858,N_8541,N_8570);
and U9859 (N_9859,N_7738,N_7836);
xor U9860 (N_9860,N_8667,N_8053);
nor U9861 (N_9861,N_7520,N_7994);
nor U9862 (N_9862,N_8138,N_8400);
xnor U9863 (N_9863,N_8095,N_8177);
nand U9864 (N_9864,N_8313,N_8604);
or U9865 (N_9865,N_8193,N_7533);
or U9866 (N_9866,N_8558,N_7875);
or U9867 (N_9867,N_8478,N_7999);
and U9868 (N_9868,N_8580,N_8277);
or U9869 (N_9869,N_7531,N_8572);
nor U9870 (N_9870,N_7537,N_7642);
nor U9871 (N_9871,N_8067,N_7730);
or U9872 (N_9872,N_8533,N_7661);
xor U9873 (N_9873,N_8057,N_8490);
xor U9874 (N_9874,N_7593,N_8433);
xnor U9875 (N_9875,N_8621,N_8395);
nand U9876 (N_9876,N_8213,N_8639);
nand U9877 (N_9877,N_7671,N_8571);
nor U9878 (N_9878,N_8657,N_8323);
and U9879 (N_9879,N_8186,N_7710);
nand U9880 (N_9880,N_7844,N_7618);
or U9881 (N_9881,N_8053,N_8733);
nor U9882 (N_9882,N_8502,N_8066);
nor U9883 (N_9883,N_8471,N_8740);
xor U9884 (N_9884,N_8529,N_8099);
or U9885 (N_9885,N_8062,N_8016);
and U9886 (N_9886,N_7534,N_8602);
and U9887 (N_9887,N_7891,N_7925);
xor U9888 (N_9888,N_7810,N_8705);
nor U9889 (N_9889,N_8670,N_7843);
nor U9890 (N_9890,N_8593,N_8088);
nor U9891 (N_9891,N_7659,N_8534);
or U9892 (N_9892,N_7555,N_8561);
nand U9893 (N_9893,N_7720,N_7742);
xor U9894 (N_9894,N_8299,N_8216);
nor U9895 (N_9895,N_7547,N_8453);
and U9896 (N_9896,N_7979,N_8287);
nor U9897 (N_9897,N_7530,N_8038);
or U9898 (N_9898,N_7589,N_8359);
nand U9899 (N_9899,N_7957,N_8442);
nand U9900 (N_9900,N_8608,N_8286);
nand U9901 (N_9901,N_7801,N_7691);
xor U9902 (N_9902,N_7693,N_7555);
or U9903 (N_9903,N_8617,N_8544);
and U9904 (N_9904,N_8221,N_7658);
and U9905 (N_9905,N_7566,N_8471);
nand U9906 (N_9906,N_8489,N_7696);
and U9907 (N_9907,N_8392,N_8456);
and U9908 (N_9908,N_8504,N_8250);
nor U9909 (N_9909,N_7635,N_8715);
or U9910 (N_9910,N_8164,N_7672);
nor U9911 (N_9911,N_8263,N_7623);
and U9912 (N_9912,N_8128,N_7569);
or U9913 (N_9913,N_8398,N_7756);
nor U9914 (N_9914,N_8465,N_7898);
and U9915 (N_9915,N_8393,N_8167);
or U9916 (N_9916,N_8144,N_8315);
and U9917 (N_9917,N_8618,N_7760);
and U9918 (N_9918,N_8064,N_8528);
and U9919 (N_9919,N_8176,N_7745);
nor U9920 (N_9920,N_7813,N_7877);
or U9921 (N_9921,N_8001,N_7569);
and U9922 (N_9922,N_8484,N_8473);
xor U9923 (N_9923,N_8210,N_8075);
xor U9924 (N_9924,N_8587,N_7641);
xor U9925 (N_9925,N_8468,N_8463);
xor U9926 (N_9926,N_7600,N_8153);
nor U9927 (N_9927,N_7556,N_8320);
and U9928 (N_9928,N_7642,N_8277);
nor U9929 (N_9929,N_8569,N_8263);
or U9930 (N_9930,N_8163,N_7688);
nor U9931 (N_9931,N_8347,N_8486);
nor U9932 (N_9932,N_7827,N_8583);
xnor U9933 (N_9933,N_8229,N_8221);
and U9934 (N_9934,N_8202,N_8496);
nand U9935 (N_9935,N_7801,N_7525);
nand U9936 (N_9936,N_7757,N_8341);
nand U9937 (N_9937,N_8088,N_7987);
nand U9938 (N_9938,N_8289,N_8326);
xor U9939 (N_9939,N_7567,N_7931);
nand U9940 (N_9940,N_8166,N_7904);
nor U9941 (N_9941,N_8332,N_7702);
xnor U9942 (N_9942,N_8737,N_8516);
or U9943 (N_9943,N_7933,N_7762);
and U9944 (N_9944,N_7961,N_8468);
nor U9945 (N_9945,N_7901,N_8713);
and U9946 (N_9946,N_8108,N_7730);
nor U9947 (N_9947,N_7877,N_8193);
nor U9948 (N_9948,N_7910,N_8713);
xor U9949 (N_9949,N_7715,N_8617);
xor U9950 (N_9950,N_8651,N_7873);
and U9951 (N_9951,N_8374,N_8441);
and U9952 (N_9952,N_7743,N_7629);
xor U9953 (N_9953,N_8603,N_8149);
nand U9954 (N_9954,N_8117,N_8180);
or U9955 (N_9955,N_8426,N_8666);
and U9956 (N_9956,N_8569,N_8164);
and U9957 (N_9957,N_7823,N_7567);
nor U9958 (N_9958,N_8388,N_8002);
nand U9959 (N_9959,N_8068,N_7598);
and U9960 (N_9960,N_8714,N_8665);
or U9961 (N_9961,N_8416,N_7870);
nand U9962 (N_9962,N_8001,N_8596);
nand U9963 (N_9963,N_7644,N_8616);
xnor U9964 (N_9964,N_8024,N_8160);
or U9965 (N_9965,N_8499,N_7986);
xor U9966 (N_9966,N_8597,N_8595);
or U9967 (N_9967,N_7808,N_8563);
or U9968 (N_9968,N_7613,N_7631);
or U9969 (N_9969,N_7645,N_7702);
xor U9970 (N_9970,N_8063,N_8603);
nor U9971 (N_9971,N_8164,N_8696);
or U9972 (N_9972,N_8143,N_8747);
nand U9973 (N_9973,N_8029,N_8274);
and U9974 (N_9974,N_7710,N_7591);
nor U9975 (N_9975,N_8659,N_7540);
xor U9976 (N_9976,N_7870,N_8722);
nor U9977 (N_9977,N_8544,N_7501);
xnor U9978 (N_9978,N_7895,N_8400);
nand U9979 (N_9979,N_8176,N_8098);
xnor U9980 (N_9980,N_8563,N_8745);
nand U9981 (N_9981,N_8400,N_8608);
or U9982 (N_9982,N_8105,N_7940);
and U9983 (N_9983,N_7538,N_7804);
or U9984 (N_9984,N_8588,N_8105);
nand U9985 (N_9985,N_8671,N_7907);
nor U9986 (N_9986,N_8046,N_7668);
or U9987 (N_9987,N_8406,N_8683);
or U9988 (N_9988,N_7537,N_8536);
nor U9989 (N_9989,N_8283,N_7762);
nor U9990 (N_9990,N_8721,N_8288);
and U9991 (N_9991,N_8428,N_7991);
and U9992 (N_9992,N_8231,N_8641);
nor U9993 (N_9993,N_8043,N_8183);
nand U9994 (N_9994,N_8450,N_8085);
or U9995 (N_9995,N_8333,N_7971);
and U9996 (N_9996,N_7738,N_8643);
nand U9997 (N_9997,N_8469,N_7667);
nor U9998 (N_9998,N_7722,N_8027);
nor U9999 (N_9999,N_8461,N_7700);
nor U10000 (N_10000,N_9002,N_9594);
nand U10001 (N_10001,N_8983,N_9881);
and U10002 (N_10002,N_9300,N_9402);
or U10003 (N_10003,N_8905,N_9458);
and U10004 (N_10004,N_9800,N_8929);
nor U10005 (N_10005,N_9589,N_9155);
and U10006 (N_10006,N_8860,N_8907);
and U10007 (N_10007,N_9350,N_9896);
nor U10008 (N_10008,N_9719,N_9373);
and U10009 (N_10009,N_9378,N_9389);
or U10010 (N_10010,N_9428,N_9552);
nor U10011 (N_10011,N_9654,N_9999);
nor U10012 (N_10012,N_9283,N_9188);
nand U10013 (N_10013,N_8834,N_9854);
nor U10014 (N_10014,N_9651,N_9924);
xnor U10015 (N_10015,N_9519,N_9319);
and U10016 (N_10016,N_9391,N_9128);
nand U10017 (N_10017,N_9837,N_9045);
and U10018 (N_10018,N_9553,N_9108);
or U10019 (N_10019,N_9359,N_9811);
and U10020 (N_10020,N_9121,N_8821);
or U10021 (N_10021,N_9931,N_8855);
and U10022 (N_10022,N_9044,N_9993);
nand U10023 (N_10023,N_9194,N_9620);
and U10024 (N_10024,N_9830,N_9114);
and U10025 (N_10025,N_8925,N_9969);
nor U10026 (N_10026,N_9991,N_9029);
xor U10027 (N_10027,N_9132,N_9603);
nor U10028 (N_10028,N_8815,N_9047);
nand U10029 (N_10029,N_8963,N_9664);
or U10030 (N_10030,N_9082,N_8814);
nand U10031 (N_10031,N_9394,N_9454);
nor U10032 (N_10032,N_9213,N_9077);
xor U10033 (N_10033,N_9789,N_9827);
nor U10034 (N_10034,N_8948,N_9731);
nor U10035 (N_10035,N_8798,N_9890);
and U10036 (N_10036,N_9901,N_8951);
or U10037 (N_10037,N_9715,N_8763);
xnor U10038 (N_10038,N_8899,N_9900);
and U10039 (N_10039,N_9368,N_8940);
or U10040 (N_10040,N_9560,N_8790);
and U10041 (N_10041,N_9873,N_9413);
or U10042 (N_10042,N_9253,N_8956);
and U10043 (N_10043,N_8941,N_8943);
and U10044 (N_10044,N_9693,N_9533);
or U10045 (N_10045,N_8961,N_9727);
nor U10046 (N_10046,N_9066,N_9052);
or U10047 (N_10047,N_8906,N_9986);
and U10048 (N_10048,N_9950,N_9752);
nand U10049 (N_10049,N_9104,N_9946);
and U10050 (N_10050,N_9624,N_9298);
or U10051 (N_10051,N_9876,N_9617);
xnor U10052 (N_10052,N_9817,N_9371);
or U10053 (N_10053,N_9060,N_9465);
and U10054 (N_10054,N_8757,N_9706);
or U10055 (N_10055,N_9497,N_8893);
or U10056 (N_10056,N_9826,N_9843);
nand U10057 (N_10057,N_9702,N_9162);
nor U10058 (N_10058,N_9437,N_8867);
or U10059 (N_10059,N_9040,N_8954);
nand U10060 (N_10060,N_9922,N_8928);
xor U10061 (N_10061,N_9495,N_9857);
nor U10062 (N_10062,N_9917,N_9557);
and U10063 (N_10063,N_8969,N_9113);
and U10064 (N_10064,N_9705,N_9261);
nand U10065 (N_10065,N_9582,N_8824);
xnor U10066 (N_10066,N_9721,N_9425);
nand U10067 (N_10067,N_9059,N_9214);
and U10068 (N_10068,N_9849,N_9947);
xor U10069 (N_10069,N_8922,N_9509);
nor U10070 (N_10070,N_9980,N_9841);
or U10071 (N_10071,N_9531,N_9545);
and U10072 (N_10072,N_8979,N_9858);
xor U10073 (N_10073,N_9846,N_9814);
nor U10074 (N_10074,N_9302,N_9206);
and U10075 (N_10075,N_9701,N_9386);
and U10076 (N_10076,N_9272,N_9358);
and U10077 (N_10077,N_9680,N_9398);
xor U10078 (N_10078,N_9227,N_8785);
xnor U10079 (N_10079,N_9597,N_9536);
xor U10080 (N_10080,N_9645,N_9202);
xnor U10081 (N_10081,N_9856,N_9877);
nand U10082 (N_10082,N_8966,N_8764);
xor U10083 (N_10083,N_9469,N_9815);
xor U10084 (N_10084,N_9136,N_9898);
or U10085 (N_10085,N_9305,N_9430);
or U10086 (N_10086,N_9483,N_9403);
nand U10087 (N_10087,N_9152,N_9912);
or U10088 (N_10088,N_8885,N_9831);
nor U10089 (N_10089,N_9166,N_8780);
nor U10090 (N_10090,N_9260,N_9092);
or U10091 (N_10091,N_8851,N_9643);
nor U10092 (N_10092,N_8888,N_9862);
or U10093 (N_10093,N_9569,N_9310);
or U10094 (N_10094,N_9007,N_9279);
xnor U10095 (N_10095,N_9333,N_8946);
nor U10096 (N_10096,N_9161,N_9888);
and U10097 (N_10097,N_9178,N_9951);
or U10098 (N_10098,N_9665,N_9717);
and U10099 (N_10099,N_9418,N_9921);
xor U10100 (N_10100,N_9954,N_9904);
nand U10101 (N_10101,N_9764,N_8870);
and U10102 (N_10102,N_9175,N_9365);
nand U10103 (N_10103,N_9055,N_9666);
and U10104 (N_10104,N_9205,N_9758);
nand U10105 (N_10105,N_9526,N_9003);
nand U10106 (N_10106,N_9252,N_8794);
xnor U10107 (N_10107,N_8765,N_9457);
nor U10108 (N_10108,N_9655,N_8848);
nand U10109 (N_10109,N_9663,N_9297);
and U10110 (N_10110,N_9238,N_9196);
or U10111 (N_10111,N_9748,N_9006);
nor U10112 (N_10112,N_9215,N_9435);
xnor U10113 (N_10113,N_8988,N_9810);
nand U10114 (N_10114,N_8989,N_9875);
nand U10115 (N_10115,N_9791,N_9119);
xnor U10116 (N_10116,N_8758,N_8932);
and U10117 (N_10117,N_9125,N_8968);
nand U10118 (N_10118,N_9224,N_8923);
or U10119 (N_10119,N_9415,N_9266);
or U10120 (N_10120,N_9153,N_8783);
nor U10121 (N_10121,N_9571,N_9646);
xor U10122 (N_10122,N_9321,N_9192);
nand U10123 (N_10123,N_9289,N_8861);
nand U10124 (N_10124,N_9230,N_9525);
xor U10125 (N_10125,N_9769,N_9158);
nor U10126 (N_10126,N_9739,N_9895);
nand U10127 (N_10127,N_9661,N_9860);
nand U10128 (N_10128,N_9117,N_9584);
nor U10129 (N_10129,N_9548,N_8995);
and U10130 (N_10130,N_9541,N_9035);
or U10131 (N_10131,N_9464,N_9422);
nand U10132 (N_10132,N_9544,N_9523);
nand U10133 (N_10133,N_9303,N_9235);
and U10134 (N_10134,N_9245,N_8942);
xor U10135 (N_10135,N_9356,N_9145);
nand U10136 (N_10136,N_9973,N_9209);
nand U10137 (N_10137,N_8914,N_9514);
nand U10138 (N_10138,N_9507,N_8804);
or U10139 (N_10139,N_9601,N_8828);
and U10140 (N_10140,N_9894,N_9799);
or U10141 (N_10141,N_8816,N_9989);
nor U10142 (N_10142,N_9143,N_9122);
or U10143 (N_10143,N_8774,N_9907);
or U10144 (N_10144,N_8916,N_8823);
xnor U10145 (N_10145,N_8777,N_9200);
nand U10146 (N_10146,N_9746,N_8931);
nor U10147 (N_10147,N_9331,N_9743);
and U10148 (N_10148,N_8820,N_8875);
and U10149 (N_10149,N_9635,N_9713);
and U10150 (N_10150,N_9649,N_8844);
and U10151 (N_10151,N_9338,N_9820);
nand U10152 (N_10152,N_8853,N_9943);
xor U10153 (N_10153,N_9336,N_9351);
xor U10154 (N_10154,N_9053,N_9237);
nor U10155 (N_10155,N_9220,N_9349);
xor U10156 (N_10156,N_9091,N_9565);
and U10157 (N_10157,N_8874,N_9619);
nor U10158 (N_10158,N_9602,N_8864);
or U10159 (N_10159,N_9376,N_8975);
and U10160 (N_10160,N_9745,N_8866);
xnor U10161 (N_10161,N_9061,N_8789);
xnor U10162 (N_10162,N_9334,N_9543);
xnor U10163 (N_10163,N_8972,N_9700);
and U10164 (N_10164,N_9674,N_8793);
and U10165 (N_10165,N_9159,N_9808);
nand U10166 (N_10166,N_8967,N_9816);
nand U10167 (N_10167,N_9588,N_9149);
and U10168 (N_10168,N_8880,N_9886);
and U10169 (N_10169,N_9195,N_9870);
nand U10170 (N_10170,N_9294,N_9903);
and U10171 (N_10171,N_9505,N_9441);
and U10172 (N_10172,N_9797,N_9967);
xor U10173 (N_10173,N_9629,N_9712);
or U10174 (N_10174,N_9257,N_8809);
xnor U10175 (N_10175,N_8750,N_9424);
or U10176 (N_10176,N_9490,N_9018);
nand U10177 (N_10177,N_8799,N_9788);
nand U10178 (N_10178,N_8918,N_8825);
nor U10179 (N_10179,N_9242,N_9547);
and U10180 (N_10180,N_9173,N_9780);
nand U10181 (N_10181,N_9453,N_9879);
and U10182 (N_10182,N_9790,N_9236);
and U10183 (N_10183,N_9186,N_9889);
nor U10184 (N_10184,N_9934,N_9793);
or U10185 (N_10185,N_9513,N_9239);
nor U10186 (N_10186,N_9852,N_9442);
nand U10187 (N_10187,N_9126,N_9183);
or U10188 (N_10188,N_9050,N_9929);
and U10189 (N_10189,N_9062,N_9691);
xor U10190 (N_10190,N_9016,N_9987);
nor U10191 (N_10191,N_9738,N_9168);
nor U10192 (N_10192,N_9024,N_9784);
nand U10193 (N_10193,N_8840,N_9618);
xnor U10194 (N_10194,N_9539,N_9421);
and U10195 (N_10195,N_9440,N_9207);
and U10196 (N_10196,N_9234,N_9399);
and U10197 (N_10197,N_9580,N_9434);
xnor U10198 (N_10198,N_9414,N_9179);
and U10199 (N_10199,N_8753,N_9281);
nor U10200 (N_10200,N_9834,N_9498);
or U10201 (N_10201,N_8775,N_9823);
nor U10202 (N_10202,N_9286,N_9595);
or U10203 (N_10203,N_9313,N_9728);
nor U10204 (N_10204,N_9246,N_9976);
or U10205 (N_10205,N_9282,N_9076);
nor U10206 (N_10206,N_9600,N_9180);
or U10207 (N_10207,N_9240,N_9388);
nor U10208 (N_10208,N_9129,N_9070);
nand U10209 (N_10209,N_9165,N_9345);
xnor U10210 (N_10210,N_9148,N_9695);
and U10211 (N_10211,N_9170,N_9716);
xnor U10212 (N_10212,N_9804,N_9787);
nor U10213 (N_10213,N_9628,N_9561);
or U10214 (N_10214,N_9147,N_9019);
and U10215 (N_10215,N_9961,N_9754);
and U10216 (N_10216,N_9491,N_8886);
or U10217 (N_10217,N_8986,N_9120);
or U10218 (N_10218,N_8927,N_9426);
and U10219 (N_10219,N_9406,N_9277);
xor U10220 (N_10220,N_9593,N_9838);
or U10221 (N_10221,N_9008,N_9749);
nor U10222 (N_10222,N_9157,N_9959);
nor U10223 (N_10223,N_9938,N_9941);
and U10224 (N_10224,N_9981,N_9337);
and U10225 (N_10225,N_9258,N_9177);
or U10226 (N_10226,N_9032,N_9933);
xor U10227 (N_10227,N_9494,N_9952);
and U10228 (N_10228,N_9069,N_9433);
and U10229 (N_10229,N_8894,N_9099);
nor U10230 (N_10230,N_9819,N_8884);
or U10231 (N_10231,N_8822,N_9354);
nand U10232 (N_10232,N_9735,N_9673);
and U10233 (N_10233,N_9201,N_9757);
or U10234 (N_10234,N_9480,N_9208);
or U10235 (N_10235,N_9322,N_8772);
and U10236 (N_10236,N_8939,N_8872);
xnor U10237 (N_10237,N_9228,N_9219);
and U10238 (N_10238,N_9293,N_9276);
and U10239 (N_10239,N_9524,N_8795);
xnor U10240 (N_10240,N_9233,N_9792);
nor U10241 (N_10241,N_9855,N_9429);
nand U10242 (N_10242,N_8778,N_9822);
xnor U10243 (N_10243,N_9504,N_9079);
nand U10244 (N_10244,N_9871,N_9596);
nor U10245 (N_10245,N_9766,N_9486);
and U10246 (N_10246,N_9572,N_9585);
nand U10247 (N_10247,N_8751,N_9264);
nand U10248 (N_10248,N_8980,N_8827);
and U10249 (N_10249,N_9778,N_8993);
or U10250 (N_10250,N_9323,N_9777);
xor U10251 (N_10251,N_9291,N_8782);
xor U10252 (N_10252,N_8920,N_8887);
nand U10253 (N_10253,N_9982,N_9438);
or U10254 (N_10254,N_9068,N_9669);
or U10255 (N_10255,N_9184,N_9250);
or U10256 (N_10256,N_8971,N_9369);
and U10257 (N_10257,N_9927,N_9756);
and U10258 (N_10258,N_9703,N_8977);
xnor U10259 (N_10259,N_9073,N_9622);
nand U10260 (N_10260,N_9866,N_9920);
nand U10261 (N_10261,N_9482,N_9449);
and U10262 (N_10262,N_9867,N_9682);
and U10263 (N_10263,N_8761,N_8755);
nor U10264 (N_10264,N_9865,N_9915);
nand U10265 (N_10265,N_9225,N_9041);
and U10266 (N_10266,N_9171,N_9802);
xor U10267 (N_10267,N_9659,N_9658);
nand U10268 (N_10268,N_9839,N_9640);
xnor U10269 (N_10269,N_8960,N_9481);
xnor U10270 (N_10270,N_9880,N_9616);
and U10271 (N_10271,N_9353,N_9431);
nor U10272 (N_10272,N_9383,N_9592);
and U10273 (N_10273,N_8877,N_9384);
nor U10274 (N_10274,N_9299,N_9806);
xor U10275 (N_10275,N_9786,N_8973);
xor U10276 (N_10276,N_9998,N_9075);
nor U10277 (N_10277,N_9112,N_9939);
nand U10278 (N_10278,N_8806,N_9254);
and U10279 (N_10279,N_9835,N_8856);
or U10280 (N_10280,N_9146,N_9436);
and U10281 (N_10281,N_9231,N_9058);
and U10282 (N_10282,N_9681,N_9477);
or U10283 (N_10283,N_9330,N_9229);
nand U10284 (N_10284,N_9021,N_9393);
nor U10285 (N_10285,N_9106,N_9734);
nand U10286 (N_10286,N_9949,N_9983);
and U10287 (N_10287,N_9656,N_9443);
and U10288 (N_10288,N_9632,N_8953);
xnor U10289 (N_10289,N_9611,N_9471);
xnor U10290 (N_10290,N_9740,N_8926);
nand U10291 (N_10291,N_9244,N_9742);
and U10292 (N_10292,N_9015,N_9885);
or U10293 (N_10293,N_9218,N_9111);
or U10294 (N_10294,N_9753,N_9642);
nor U10295 (N_10295,N_9028,N_9517);
and U10296 (N_10296,N_9730,N_8846);
and U10297 (N_10297,N_8921,N_9566);
nand U10298 (N_10298,N_9647,N_9892);
xnor U10299 (N_10299,N_9361,N_8810);
and U10300 (N_10300,N_9172,N_9385);
xor U10301 (N_10301,N_9977,N_8903);
nor U10302 (N_10302,N_9785,N_9833);
or U10303 (N_10303,N_9247,N_9427);
nand U10304 (N_10304,N_9893,N_9290);
xor U10305 (N_10305,N_9312,N_9935);
xor U10306 (N_10306,N_9908,N_9670);
nand U10307 (N_10307,N_9573,N_9472);
nand U10308 (N_10308,N_9466,N_9897);
nand U10309 (N_10309,N_9086,N_8832);
nor U10310 (N_10310,N_9096,N_9380);
nand U10311 (N_10311,N_9304,N_9515);
nor U10312 (N_10312,N_8768,N_9049);
or U10313 (N_10313,N_8957,N_9853);
xnor U10314 (N_10314,N_9948,N_9563);
nand U10315 (N_10315,N_9473,N_8857);
or U10316 (N_10316,N_9057,N_8805);
nor U10317 (N_10317,N_9767,N_8917);
nor U10318 (N_10318,N_9134,N_9056);
or U10319 (N_10319,N_9733,N_9905);
nor U10320 (N_10320,N_9783,N_9295);
or U10321 (N_10321,N_9071,N_8817);
nor U10322 (N_10322,N_9474,N_8997);
and U10323 (N_10323,N_9970,N_9836);
and U10324 (N_10324,N_9088,N_9599);
or U10325 (N_10325,N_9328,N_9444);
nand U10326 (N_10326,N_8981,N_9499);
xor U10327 (N_10327,N_9031,N_9621);
nor U10328 (N_10328,N_9847,N_9825);
or U10329 (N_10329,N_9335,N_8770);
nor U10330 (N_10330,N_9615,N_9249);
or U10331 (N_10331,N_9420,N_8788);
or U10332 (N_10332,N_8762,N_9942);
and U10333 (N_10333,N_8800,N_8970);
and U10334 (N_10334,N_9211,N_9492);
nand U10335 (N_10335,N_8883,N_8933);
or U10336 (N_10336,N_9671,N_9906);
xor U10337 (N_10337,N_9005,N_9962);
xnor U10338 (N_10338,N_8792,N_9614);
and U10339 (N_10339,N_9567,N_9555);
or U10340 (N_10340,N_9559,N_8959);
nor U10341 (N_10341,N_9794,N_9568);
nor U10342 (N_10342,N_9704,N_8958);
xnor U10343 (N_10343,N_8919,N_9275);
xnor U10344 (N_10344,N_9583,N_9913);
xor U10345 (N_10345,N_9953,N_9193);
nor U10346 (N_10346,N_8991,N_9990);
nand U10347 (N_10347,N_9033,N_9714);
or U10348 (N_10348,N_9975,N_9039);
or U10349 (N_10349,N_9164,N_9578);
xnor U10350 (N_10350,N_9660,N_9127);
nor U10351 (N_10351,N_9637,N_8950);
nand U10352 (N_10352,N_8974,N_9190);
and U10353 (N_10353,N_9607,N_9925);
and U10354 (N_10354,N_9410,N_9707);
and U10355 (N_10355,N_9530,N_9102);
and U10356 (N_10356,N_9577,N_9496);
or U10357 (N_10357,N_9074,N_9613);
xor U10358 (N_10358,N_9226,N_9022);
xor U10359 (N_10359,N_8930,N_9636);
nand U10360 (N_10360,N_9914,N_9452);
xor U10361 (N_10361,N_8766,N_9736);
or U10362 (N_10362,N_9098,N_8879);
and U10363 (N_10363,N_9087,N_9737);
nand U10364 (N_10364,N_8852,N_8819);
and U10365 (N_10365,N_9185,N_9626);
and U10366 (N_10366,N_9285,N_9564);
and U10367 (N_10367,N_9280,N_9095);
xor U10368 (N_10368,N_9411,N_9850);
nor U10369 (N_10369,N_8826,N_9964);
or U10370 (N_10370,N_9212,N_9500);
xnor U10371 (N_10371,N_9639,N_8996);
nor U10372 (N_10372,N_9189,N_9634);
or U10373 (N_10373,N_9828,N_8900);
or U10374 (N_10374,N_9447,N_9324);
nand U10375 (N_10375,N_9824,N_9677);
or U10376 (N_10376,N_9037,N_9110);
nor U10377 (N_10377,N_8998,N_9397);
xnor U10378 (N_10378,N_9692,N_9940);
xor U10379 (N_10379,N_9030,N_8891);
nor U10380 (N_10380,N_9156,N_9124);
and U10381 (N_10381,N_9768,N_9803);
nor U10382 (N_10382,N_8831,N_9722);
nor U10383 (N_10383,N_9014,N_9775);
nor U10384 (N_10384,N_9273,N_9342);
nor U10385 (N_10385,N_9489,N_9537);
nor U10386 (N_10386,N_9902,N_8802);
nand U10387 (N_10387,N_9100,N_9538);
and U10388 (N_10388,N_8978,N_9529);
nor U10389 (N_10389,N_9510,N_9248);
xnor U10390 (N_10390,N_9267,N_9259);
or U10391 (N_10391,N_9417,N_8962);
and U10392 (N_10392,N_9137,N_9844);
nand U10393 (N_10393,N_8898,N_9375);
nand U10394 (N_10394,N_9360,N_8786);
nor U10395 (N_10395,N_9404,N_9340);
xor U10396 (N_10396,N_9478,N_9868);
and U10397 (N_10397,N_8811,N_9461);
nand U10398 (N_10398,N_9484,N_9899);
or U10399 (N_10399,N_9027,N_8773);
nor U10400 (N_10400,N_9861,N_8752);
and U10401 (N_10401,N_8797,N_9809);
or U10402 (N_10402,N_9678,N_8796);
nor U10403 (N_10403,N_9926,N_9093);
or U10404 (N_10404,N_9084,N_9199);
or U10405 (N_10405,N_9916,N_9762);
or U10406 (N_10406,N_8787,N_9796);
and U10407 (N_10407,N_9772,N_8901);
xnor U10408 (N_10408,N_9690,N_9832);
nor U10409 (N_10409,N_9366,N_9741);
nand U10410 (N_10410,N_9381,N_9936);
nor U10411 (N_10411,N_9503,N_9488);
nand U10412 (N_10412,N_9667,N_9653);
and U10413 (N_10413,N_9017,N_8803);
xor U10414 (N_10414,N_9487,N_8902);
or U10415 (N_10415,N_9840,N_9587);
nor U10416 (N_10416,N_9263,N_8873);
or U10417 (N_10417,N_9204,N_9141);
nor U10418 (N_10418,N_9910,N_9181);
and U10419 (N_10419,N_9988,N_9689);
nor U10420 (N_10420,N_8889,N_9374);
and U10421 (N_10421,N_9221,N_8838);
nor U10422 (N_10422,N_9115,N_9562);
or U10423 (N_10423,N_9818,N_9995);
nor U10424 (N_10424,N_9026,N_9996);
and U10425 (N_10425,N_9955,N_8836);
xnor U10426 (N_10426,N_9009,N_9506);
or U10427 (N_10427,N_9042,N_9025);
and U10428 (N_10428,N_9627,N_9699);
and U10429 (N_10429,N_9135,N_9944);
and U10430 (N_10430,N_8801,N_8912);
and U10431 (N_10431,N_9997,N_8813);
nor U10432 (N_10432,N_9222,N_9958);
nand U10433 (N_10433,N_8837,N_9608);
xor U10434 (N_10434,N_9038,N_9798);
and U10435 (N_10435,N_9329,N_9405);
nand U10436 (N_10436,N_9462,N_9390);
and U10437 (N_10437,N_9672,N_9937);
nor U10438 (N_10438,N_9644,N_9364);
nand U10439 (N_10439,N_8935,N_9012);
or U10440 (N_10440,N_8854,N_8830);
nand U10441 (N_10441,N_8987,N_9255);
nand U10442 (N_10442,N_9382,N_9064);
xnor U10443 (N_10443,N_9274,N_9151);
nand U10444 (N_10444,N_9774,N_9262);
nor U10445 (N_10445,N_9455,N_9210);
nor U10446 (N_10446,N_9232,N_9090);
xor U10447 (N_10447,N_9698,N_9325);
xnor U10448 (N_10448,N_9859,N_9470);
nand U10449 (N_10449,N_9341,N_9570);
and U10450 (N_10450,N_9043,N_9187);
nor U10451 (N_10451,N_9685,N_9918);
nand U10452 (N_10452,N_9103,N_8769);
xor U10453 (N_10453,N_9048,N_9668);
xnor U10454 (N_10454,N_9972,N_9864);
or U10455 (N_10455,N_9109,N_8760);
nor U10456 (N_10456,N_9154,N_8847);
nor U10457 (N_10457,N_9377,N_9508);
nand U10458 (N_10458,N_9747,N_9697);
xnor U10459 (N_10459,N_9779,N_9590);
nand U10460 (N_10460,N_9456,N_9432);
or U10461 (N_10461,N_9191,N_9367);
nor U10462 (N_10462,N_8829,N_9884);
nand U10463 (N_10463,N_9686,N_9054);
xor U10464 (N_10464,N_9416,N_9251);
nand U10465 (N_10465,N_9203,N_9930);
or U10466 (N_10466,N_8904,N_8849);
xnor U10467 (N_10467,N_9726,N_9270);
and U10468 (N_10468,N_9216,N_9795);
xnor U10469 (N_10469,N_8955,N_9306);
nor U10470 (N_10470,N_9805,N_9451);
nand U10471 (N_10471,N_8759,N_9842);
nand U10472 (N_10472,N_9650,N_9046);
xnor U10473 (N_10473,N_9710,N_9460);
nand U10474 (N_10474,N_9348,N_9966);
nor U10475 (N_10475,N_9140,N_9763);
or U10476 (N_10476,N_8839,N_8892);
nor U10477 (N_10477,N_8863,N_9314);
xnor U10478 (N_10478,N_9945,N_8909);
and U10479 (N_10479,N_9848,N_9409);
nand U10480 (N_10480,N_8833,N_9485);
xor U10481 (N_10481,N_8807,N_9339);
nand U10482 (N_10482,N_9511,N_9105);
or U10483 (N_10483,N_9150,N_8858);
nand U10484 (N_10484,N_8896,N_9287);
nor U10485 (N_10485,N_9542,N_8964);
and U10486 (N_10486,N_9586,N_9475);
nor U10487 (N_10487,N_9268,N_9520);
nor U10488 (N_10488,N_9528,N_9744);
nand U10489 (N_10489,N_9080,N_8982);
nor U10490 (N_10490,N_8882,N_9459);
nor U10491 (N_10491,N_8841,N_9807);
or U10492 (N_10492,N_9392,N_9610);
nand U10493 (N_10493,N_9065,N_8924);
and U10494 (N_10494,N_9708,N_9662);
and U10495 (N_10495,N_9308,N_9363);
nor U10496 (N_10496,N_9676,N_9501);
or U10497 (N_10497,N_9932,N_8945);
nand U10498 (N_10498,N_9067,N_8771);
xor U10499 (N_10499,N_9309,N_9732);
and U10500 (N_10500,N_8881,N_9874);
nand U10501 (N_10501,N_9476,N_9512);
nand U10502 (N_10502,N_9284,N_8999);
xor U10503 (N_10503,N_9133,N_9241);
or U10504 (N_10504,N_9243,N_9089);
nand U10505 (N_10505,N_8754,N_9423);
xnor U10506 (N_10506,N_9357,N_9493);
nor U10507 (N_10507,N_9863,N_9372);
nor U10508 (N_10508,N_9549,N_8812);
xnor U10509 (N_10509,N_9869,N_8869);
nand U10510 (N_10510,N_8842,N_9131);
xor U10511 (N_10511,N_9591,N_9142);
or U10512 (N_10512,N_9985,N_9540);
xnor U10513 (N_10513,N_9326,N_9004);
nor U10514 (N_10514,N_9138,N_9971);
and U10515 (N_10515,N_9821,N_9909);
or U10516 (N_10516,N_9311,N_9083);
or U10517 (N_10517,N_9521,N_9891);
or U10518 (N_10518,N_9527,N_9684);
and U10519 (N_10519,N_9729,N_9957);
xnor U10520 (N_10520,N_9094,N_9965);
xnor U10521 (N_10521,N_9174,N_9554);
and U10522 (N_10522,N_8808,N_8994);
and U10523 (N_10523,N_9288,N_9097);
xor U10524 (N_10524,N_8781,N_9446);
nor U10525 (N_10525,N_9269,N_9575);
nor U10526 (N_10526,N_9558,N_9343);
or U10527 (N_10527,N_9657,N_8936);
xnor U10528 (N_10528,N_9072,N_9307);
and U10529 (N_10529,N_9718,N_9332);
nand U10530 (N_10530,N_9387,N_8944);
and U10531 (N_10531,N_9760,N_9812);
or U10532 (N_10532,N_9407,N_9923);
xor U10533 (N_10533,N_9638,N_8776);
xnor U10534 (N_10534,N_9401,N_9773);
nor U10535 (N_10535,N_9606,N_9010);
nand U10536 (N_10536,N_9408,N_9502);
nand U10537 (N_10537,N_9036,N_9623);
nor U10538 (N_10538,N_9362,N_9063);
nand U10539 (N_10539,N_9759,N_8890);
or U10540 (N_10540,N_9412,N_8937);
nand U10541 (N_10541,N_9883,N_9468);
and U10542 (N_10542,N_9160,N_8862);
nand U10543 (N_10543,N_9450,N_9101);
xor U10544 (N_10544,N_8976,N_9751);
nand U10545 (N_10545,N_9327,N_9605);
xor U10546 (N_10546,N_9801,N_9872);
nand U10547 (N_10547,N_9984,N_9518);
xor U10548 (N_10548,N_9167,N_9724);
nor U10549 (N_10549,N_9217,N_9516);
and U10550 (N_10550,N_9223,N_9845);
and U10551 (N_10551,N_9318,N_9169);
xnor U10552 (N_10552,N_9765,N_8910);
nor U10553 (N_10553,N_9001,N_8908);
nor U10554 (N_10554,N_9439,N_9604);
nor U10555 (N_10555,N_9320,N_9301);
nand U10556 (N_10556,N_9000,N_9723);
xnor U10557 (N_10557,N_9887,N_9198);
nor U10558 (N_10558,N_9346,N_8915);
nand U10559 (N_10559,N_9770,N_9696);
or U10560 (N_10560,N_9919,N_9522);
and U10561 (N_10561,N_9535,N_8835);
or U10562 (N_10562,N_9396,N_9720);
xor U10563 (N_10563,N_8784,N_9347);
or U10564 (N_10564,N_8850,N_9344);
nand U10565 (N_10565,N_9020,N_9574);
nand U10566 (N_10566,N_9771,N_8949);
nand U10567 (N_10567,N_9448,N_9576);
and U10568 (N_10568,N_9315,N_9355);
nand U10569 (N_10569,N_9581,N_9598);
or U10570 (N_10570,N_8934,N_9445);
nand U10571 (N_10571,N_8878,N_8965);
xnor U10572 (N_10572,N_9782,N_9278);
nor U10573 (N_10573,N_9551,N_9316);
xnor U10574 (N_10574,N_9679,N_9878);
nand U10575 (N_10575,N_9761,N_9652);
nor U10576 (N_10576,N_9370,N_9265);
or U10577 (N_10577,N_8767,N_8938);
nor U10578 (N_10578,N_9963,N_9755);
nor U10579 (N_10579,N_9750,N_9694);
and U10580 (N_10580,N_9081,N_9400);
or U10581 (N_10581,N_9994,N_9296);
nor U10582 (N_10582,N_9683,N_8756);
xor U10583 (N_10583,N_8845,N_9725);
and U10584 (N_10584,N_8876,N_9534);
nand U10585 (N_10585,N_9118,N_9479);
and U10586 (N_10586,N_8897,N_8818);
nand U10587 (N_10587,N_9928,N_8865);
xor U10588 (N_10588,N_9011,N_9139);
or U10589 (N_10589,N_9271,N_9051);
and U10590 (N_10590,N_8985,N_9532);
nand U10591 (N_10591,N_9467,N_9630);
and U10592 (N_10592,N_8791,N_9463);
nand U10593 (N_10593,N_9813,N_9709);
and U10594 (N_10594,N_9144,N_8868);
nand U10595 (N_10595,N_9979,N_9612);
and U10596 (N_10596,N_9631,N_9123);
or U10597 (N_10597,N_9546,N_9882);
and U10598 (N_10598,N_8895,N_8952);
and U10599 (N_10599,N_9992,N_9956);
nand U10600 (N_10600,N_9163,N_9256);
xnor U10601 (N_10601,N_9085,N_8871);
xor U10602 (N_10602,N_9419,N_9352);
nand U10603 (N_10603,N_8947,N_9978);
nand U10604 (N_10604,N_9641,N_8990);
and U10605 (N_10605,N_9182,N_9675);
or U10606 (N_10606,N_9078,N_9851);
or U10607 (N_10607,N_9013,N_9550);
or U10608 (N_10608,N_9292,N_8859);
or U10609 (N_10609,N_9633,N_9556);
xor U10610 (N_10610,N_9625,N_9968);
nand U10611 (N_10611,N_9648,N_9687);
nor U10612 (N_10612,N_9911,N_9579);
xor U10613 (N_10613,N_8779,N_9023);
nor U10614 (N_10614,N_9379,N_9688);
nor U10615 (N_10615,N_8843,N_9609);
and U10616 (N_10616,N_8911,N_9395);
or U10617 (N_10617,N_9197,N_8984);
nor U10618 (N_10618,N_9974,N_9317);
nand U10619 (N_10619,N_9034,N_8913);
nand U10620 (N_10620,N_9107,N_9776);
or U10621 (N_10621,N_9960,N_9130);
and U10622 (N_10622,N_9829,N_8992);
nor U10623 (N_10623,N_9116,N_9711);
nor U10624 (N_10624,N_9781,N_9176);
nor U10625 (N_10625,N_8830,N_8946);
or U10626 (N_10626,N_8782,N_9805);
and U10627 (N_10627,N_8868,N_9514);
and U10628 (N_10628,N_9475,N_9035);
or U10629 (N_10629,N_9476,N_9087);
xor U10630 (N_10630,N_9424,N_8903);
and U10631 (N_10631,N_9277,N_9233);
nand U10632 (N_10632,N_9934,N_9672);
xor U10633 (N_10633,N_9513,N_9332);
xnor U10634 (N_10634,N_9006,N_9028);
xnor U10635 (N_10635,N_9585,N_8813);
or U10636 (N_10636,N_9948,N_8818);
nand U10637 (N_10637,N_8927,N_9773);
xor U10638 (N_10638,N_9220,N_9571);
nand U10639 (N_10639,N_9817,N_9355);
nor U10640 (N_10640,N_8944,N_8754);
xor U10641 (N_10641,N_8934,N_9366);
and U10642 (N_10642,N_9149,N_8825);
nand U10643 (N_10643,N_9188,N_9180);
xor U10644 (N_10644,N_9062,N_9585);
nand U10645 (N_10645,N_9408,N_9949);
nor U10646 (N_10646,N_9198,N_9363);
and U10647 (N_10647,N_9620,N_9464);
and U10648 (N_10648,N_9598,N_9053);
nor U10649 (N_10649,N_9211,N_9380);
nor U10650 (N_10650,N_8929,N_9267);
and U10651 (N_10651,N_8834,N_9907);
and U10652 (N_10652,N_9408,N_9414);
nor U10653 (N_10653,N_9754,N_9481);
or U10654 (N_10654,N_9401,N_9922);
nand U10655 (N_10655,N_9913,N_9288);
nor U10656 (N_10656,N_9119,N_9256);
or U10657 (N_10657,N_9461,N_8846);
xnor U10658 (N_10658,N_9558,N_9118);
xnor U10659 (N_10659,N_9443,N_9802);
nor U10660 (N_10660,N_8967,N_9979);
nor U10661 (N_10661,N_9313,N_9058);
xor U10662 (N_10662,N_9529,N_8838);
or U10663 (N_10663,N_9894,N_8979);
nor U10664 (N_10664,N_8865,N_8771);
or U10665 (N_10665,N_9725,N_9635);
xnor U10666 (N_10666,N_9037,N_9116);
xnor U10667 (N_10667,N_9119,N_9787);
nor U10668 (N_10668,N_9172,N_9553);
xor U10669 (N_10669,N_9395,N_9099);
nand U10670 (N_10670,N_9903,N_8810);
or U10671 (N_10671,N_9770,N_9328);
xor U10672 (N_10672,N_9306,N_9307);
nand U10673 (N_10673,N_8882,N_9433);
or U10674 (N_10674,N_9869,N_9710);
and U10675 (N_10675,N_9110,N_9835);
nand U10676 (N_10676,N_9431,N_9868);
nor U10677 (N_10677,N_9139,N_9779);
or U10678 (N_10678,N_9914,N_9673);
nor U10679 (N_10679,N_9874,N_9557);
xnor U10680 (N_10680,N_9994,N_9142);
or U10681 (N_10681,N_9897,N_9062);
nand U10682 (N_10682,N_9875,N_9542);
nand U10683 (N_10683,N_9495,N_9485);
or U10684 (N_10684,N_8856,N_9561);
and U10685 (N_10685,N_9013,N_9631);
and U10686 (N_10686,N_9101,N_9116);
or U10687 (N_10687,N_9091,N_8999);
nor U10688 (N_10688,N_8879,N_9369);
or U10689 (N_10689,N_9122,N_8925);
and U10690 (N_10690,N_9469,N_9108);
nor U10691 (N_10691,N_8904,N_9120);
xnor U10692 (N_10692,N_9303,N_8838);
and U10693 (N_10693,N_9611,N_9102);
or U10694 (N_10694,N_9327,N_9833);
xor U10695 (N_10695,N_9559,N_9806);
xnor U10696 (N_10696,N_8998,N_9302);
and U10697 (N_10697,N_9662,N_9034);
or U10698 (N_10698,N_9646,N_9296);
and U10699 (N_10699,N_9946,N_9154);
nor U10700 (N_10700,N_9192,N_8760);
or U10701 (N_10701,N_9528,N_9046);
or U10702 (N_10702,N_9476,N_9486);
nand U10703 (N_10703,N_8937,N_9206);
and U10704 (N_10704,N_9925,N_9017);
nand U10705 (N_10705,N_9813,N_9783);
and U10706 (N_10706,N_8821,N_8862);
or U10707 (N_10707,N_9354,N_9633);
xnor U10708 (N_10708,N_9536,N_9327);
and U10709 (N_10709,N_9984,N_9023);
nor U10710 (N_10710,N_8979,N_8845);
xnor U10711 (N_10711,N_9187,N_9748);
or U10712 (N_10712,N_9279,N_8784);
and U10713 (N_10713,N_8863,N_9434);
nand U10714 (N_10714,N_9560,N_9972);
or U10715 (N_10715,N_9785,N_9816);
nor U10716 (N_10716,N_9354,N_9231);
nor U10717 (N_10717,N_9503,N_9714);
xnor U10718 (N_10718,N_8920,N_8883);
nand U10719 (N_10719,N_8846,N_9303);
or U10720 (N_10720,N_9613,N_8882);
nor U10721 (N_10721,N_9973,N_8994);
or U10722 (N_10722,N_9060,N_8911);
or U10723 (N_10723,N_9571,N_9815);
xor U10724 (N_10724,N_9229,N_8997);
xnor U10725 (N_10725,N_9306,N_8866);
nor U10726 (N_10726,N_9943,N_8828);
and U10727 (N_10727,N_9186,N_9904);
and U10728 (N_10728,N_8971,N_8821);
or U10729 (N_10729,N_9990,N_9510);
nand U10730 (N_10730,N_9797,N_9831);
xnor U10731 (N_10731,N_9343,N_9566);
or U10732 (N_10732,N_9516,N_8884);
nand U10733 (N_10733,N_8844,N_9487);
xnor U10734 (N_10734,N_9233,N_9878);
xor U10735 (N_10735,N_9359,N_9910);
xnor U10736 (N_10736,N_9439,N_9939);
nand U10737 (N_10737,N_9787,N_9218);
or U10738 (N_10738,N_9451,N_9730);
and U10739 (N_10739,N_9616,N_8787);
xnor U10740 (N_10740,N_9888,N_9032);
nand U10741 (N_10741,N_9857,N_8848);
and U10742 (N_10742,N_8942,N_8824);
xor U10743 (N_10743,N_9891,N_9279);
xnor U10744 (N_10744,N_9754,N_9544);
nor U10745 (N_10745,N_9431,N_8914);
or U10746 (N_10746,N_9023,N_9870);
nand U10747 (N_10747,N_9767,N_9926);
and U10748 (N_10748,N_9956,N_8837);
or U10749 (N_10749,N_9580,N_8804);
nand U10750 (N_10750,N_8831,N_9219);
nand U10751 (N_10751,N_9621,N_9914);
xnor U10752 (N_10752,N_9955,N_8915);
xnor U10753 (N_10753,N_9569,N_9441);
or U10754 (N_10754,N_9223,N_9137);
nand U10755 (N_10755,N_9464,N_9835);
and U10756 (N_10756,N_9284,N_9180);
nand U10757 (N_10757,N_9504,N_9891);
and U10758 (N_10758,N_9106,N_9289);
xor U10759 (N_10759,N_9781,N_9066);
and U10760 (N_10760,N_9326,N_9654);
nor U10761 (N_10761,N_9412,N_9133);
xnor U10762 (N_10762,N_9888,N_9570);
nor U10763 (N_10763,N_8911,N_9444);
xor U10764 (N_10764,N_9314,N_9366);
or U10765 (N_10765,N_8769,N_9990);
and U10766 (N_10766,N_9697,N_8883);
or U10767 (N_10767,N_9986,N_9583);
xor U10768 (N_10768,N_9758,N_9216);
and U10769 (N_10769,N_9783,N_9867);
nor U10770 (N_10770,N_9021,N_9651);
nor U10771 (N_10771,N_9181,N_9199);
or U10772 (N_10772,N_9902,N_9654);
and U10773 (N_10773,N_9167,N_9424);
or U10774 (N_10774,N_9316,N_9890);
nor U10775 (N_10775,N_8904,N_9700);
nand U10776 (N_10776,N_9653,N_8870);
nand U10777 (N_10777,N_9691,N_9147);
nand U10778 (N_10778,N_9443,N_8942);
or U10779 (N_10779,N_9342,N_9796);
and U10780 (N_10780,N_9080,N_9832);
or U10781 (N_10781,N_9449,N_9335);
nand U10782 (N_10782,N_9891,N_8957);
and U10783 (N_10783,N_8953,N_9826);
xor U10784 (N_10784,N_9876,N_9542);
nor U10785 (N_10785,N_9915,N_9338);
nor U10786 (N_10786,N_9090,N_8846);
and U10787 (N_10787,N_9989,N_9276);
xnor U10788 (N_10788,N_9261,N_9085);
and U10789 (N_10789,N_9468,N_8988);
nor U10790 (N_10790,N_9430,N_9677);
xnor U10791 (N_10791,N_9399,N_9130);
nand U10792 (N_10792,N_8837,N_9420);
xnor U10793 (N_10793,N_9789,N_8940);
xor U10794 (N_10794,N_9022,N_8835);
nor U10795 (N_10795,N_9624,N_9524);
or U10796 (N_10796,N_8799,N_9845);
and U10797 (N_10797,N_9884,N_8999);
or U10798 (N_10798,N_9623,N_9189);
or U10799 (N_10799,N_8783,N_9841);
and U10800 (N_10800,N_9091,N_8991);
xnor U10801 (N_10801,N_9719,N_9912);
or U10802 (N_10802,N_9796,N_9886);
and U10803 (N_10803,N_9727,N_9094);
nand U10804 (N_10804,N_9538,N_9194);
xor U10805 (N_10805,N_9146,N_9127);
nand U10806 (N_10806,N_9825,N_9803);
nand U10807 (N_10807,N_9495,N_9062);
or U10808 (N_10808,N_9262,N_9218);
xor U10809 (N_10809,N_9878,N_9923);
xor U10810 (N_10810,N_9860,N_9157);
and U10811 (N_10811,N_9020,N_9669);
nand U10812 (N_10812,N_9825,N_9982);
xnor U10813 (N_10813,N_9291,N_9951);
or U10814 (N_10814,N_8967,N_9303);
nand U10815 (N_10815,N_9361,N_9247);
nand U10816 (N_10816,N_9709,N_9017);
and U10817 (N_10817,N_9382,N_9182);
xor U10818 (N_10818,N_9590,N_9876);
nor U10819 (N_10819,N_9634,N_8843);
nand U10820 (N_10820,N_9722,N_8891);
nor U10821 (N_10821,N_9975,N_9379);
nor U10822 (N_10822,N_8837,N_8999);
nand U10823 (N_10823,N_9359,N_9387);
or U10824 (N_10824,N_9271,N_9972);
and U10825 (N_10825,N_9251,N_8752);
and U10826 (N_10826,N_9391,N_9556);
nor U10827 (N_10827,N_9724,N_9976);
nor U10828 (N_10828,N_8789,N_9343);
and U10829 (N_10829,N_9736,N_9495);
or U10830 (N_10830,N_9762,N_9639);
nor U10831 (N_10831,N_9885,N_9835);
or U10832 (N_10832,N_9451,N_9942);
or U10833 (N_10833,N_9216,N_8796);
or U10834 (N_10834,N_9281,N_8949);
and U10835 (N_10835,N_9832,N_9610);
nor U10836 (N_10836,N_9962,N_9635);
nor U10837 (N_10837,N_9450,N_9926);
xor U10838 (N_10838,N_9653,N_9881);
nor U10839 (N_10839,N_9120,N_9652);
nand U10840 (N_10840,N_8764,N_9988);
or U10841 (N_10841,N_8759,N_9225);
and U10842 (N_10842,N_9516,N_9868);
and U10843 (N_10843,N_9751,N_9576);
and U10844 (N_10844,N_9247,N_9046);
nand U10845 (N_10845,N_9276,N_9688);
or U10846 (N_10846,N_9280,N_9001);
xnor U10847 (N_10847,N_9054,N_9259);
or U10848 (N_10848,N_9493,N_9896);
xor U10849 (N_10849,N_9292,N_9685);
xnor U10850 (N_10850,N_9876,N_8832);
or U10851 (N_10851,N_8801,N_8825);
nor U10852 (N_10852,N_8792,N_8934);
and U10853 (N_10853,N_9517,N_9689);
xor U10854 (N_10854,N_9227,N_8904);
or U10855 (N_10855,N_9897,N_9250);
or U10856 (N_10856,N_8990,N_9404);
and U10857 (N_10857,N_9748,N_9696);
nor U10858 (N_10858,N_9909,N_9409);
nand U10859 (N_10859,N_9434,N_9712);
xor U10860 (N_10860,N_9189,N_8936);
nand U10861 (N_10861,N_9811,N_9661);
xnor U10862 (N_10862,N_9259,N_9812);
xnor U10863 (N_10863,N_8817,N_9365);
nand U10864 (N_10864,N_9610,N_9200);
or U10865 (N_10865,N_9338,N_9406);
or U10866 (N_10866,N_9727,N_9297);
or U10867 (N_10867,N_9465,N_8809);
nor U10868 (N_10868,N_9871,N_9177);
and U10869 (N_10869,N_9567,N_9178);
xnor U10870 (N_10870,N_9034,N_9072);
or U10871 (N_10871,N_8830,N_9535);
nor U10872 (N_10872,N_9055,N_9588);
and U10873 (N_10873,N_9777,N_8780);
or U10874 (N_10874,N_8864,N_9208);
and U10875 (N_10875,N_9607,N_9719);
and U10876 (N_10876,N_9312,N_9990);
nand U10877 (N_10877,N_9866,N_9343);
xnor U10878 (N_10878,N_9282,N_9037);
nand U10879 (N_10879,N_9514,N_9044);
xnor U10880 (N_10880,N_9025,N_8804);
xnor U10881 (N_10881,N_9590,N_8973);
nand U10882 (N_10882,N_9312,N_9886);
xnor U10883 (N_10883,N_9805,N_9319);
nand U10884 (N_10884,N_9506,N_8835);
nand U10885 (N_10885,N_8795,N_9997);
or U10886 (N_10886,N_9325,N_9795);
or U10887 (N_10887,N_8856,N_9027);
or U10888 (N_10888,N_8839,N_9232);
xnor U10889 (N_10889,N_9565,N_9352);
nand U10890 (N_10890,N_9065,N_9011);
or U10891 (N_10891,N_8935,N_9233);
xor U10892 (N_10892,N_9937,N_9642);
xor U10893 (N_10893,N_9967,N_9289);
or U10894 (N_10894,N_9663,N_9158);
nand U10895 (N_10895,N_9235,N_9228);
nand U10896 (N_10896,N_9953,N_9995);
nand U10897 (N_10897,N_9142,N_9608);
nor U10898 (N_10898,N_9765,N_9729);
or U10899 (N_10899,N_8988,N_9973);
nor U10900 (N_10900,N_8772,N_8943);
xnor U10901 (N_10901,N_9574,N_9923);
and U10902 (N_10902,N_9489,N_9203);
nor U10903 (N_10903,N_9442,N_9737);
and U10904 (N_10904,N_9870,N_9531);
nand U10905 (N_10905,N_9828,N_9964);
xor U10906 (N_10906,N_9063,N_9664);
and U10907 (N_10907,N_9538,N_9537);
nor U10908 (N_10908,N_9160,N_9038);
nand U10909 (N_10909,N_9176,N_8805);
xor U10910 (N_10910,N_9113,N_9849);
nand U10911 (N_10911,N_9800,N_9994);
nand U10912 (N_10912,N_9919,N_9463);
xnor U10913 (N_10913,N_9784,N_9617);
xor U10914 (N_10914,N_9163,N_9637);
and U10915 (N_10915,N_8850,N_9572);
or U10916 (N_10916,N_9415,N_9628);
nand U10917 (N_10917,N_8875,N_9449);
nand U10918 (N_10918,N_9377,N_8837);
xnor U10919 (N_10919,N_8793,N_8778);
and U10920 (N_10920,N_9572,N_9740);
nand U10921 (N_10921,N_9955,N_9757);
nand U10922 (N_10922,N_9965,N_9004);
nor U10923 (N_10923,N_9945,N_8792);
xnor U10924 (N_10924,N_8784,N_9406);
nor U10925 (N_10925,N_9003,N_9272);
xnor U10926 (N_10926,N_9751,N_9044);
or U10927 (N_10927,N_8854,N_9727);
nor U10928 (N_10928,N_8751,N_8818);
nand U10929 (N_10929,N_9198,N_9048);
and U10930 (N_10930,N_8940,N_9982);
and U10931 (N_10931,N_9996,N_9053);
nand U10932 (N_10932,N_8999,N_9734);
nor U10933 (N_10933,N_9287,N_9683);
and U10934 (N_10934,N_9237,N_9446);
nor U10935 (N_10935,N_9849,N_9864);
nand U10936 (N_10936,N_9229,N_8840);
and U10937 (N_10937,N_8907,N_8769);
xnor U10938 (N_10938,N_9391,N_9415);
or U10939 (N_10939,N_9340,N_9983);
nor U10940 (N_10940,N_9137,N_9704);
and U10941 (N_10941,N_9295,N_9684);
nor U10942 (N_10942,N_8785,N_9224);
nand U10943 (N_10943,N_9924,N_8833);
nand U10944 (N_10944,N_8907,N_9321);
nand U10945 (N_10945,N_9733,N_9964);
nand U10946 (N_10946,N_8922,N_9031);
xnor U10947 (N_10947,N_8757,N_9155);
xnor U10948 (N_10948,N_9180,N_9224);
nor U10949 (N_10949,N_9380,N_9608);
xor U10950 (N_10950,N_8822,N_9506);
nor U10951 (N_10951,N_9001,N_9975);
and U10952 (N_10952,N_9874,N_9757);
and U10953 (N_10953,N_9447,N_9984);
nor U10954 (N_10954,N_8832,N_9426);
and U10955 (N_10955,N_9200,N_8799);
nor U10956 (N_10956,N_9988,N_9638);
nor U10957 (N_10957,N_9451,N_9950);
or U10958 (N_10958,N_8899,N_9846);
xor U10959 (N_10959,N_9207,N_9683);
or U10960 (N_10960,N_8930,N_9843);
xor U10961 (N_10961,N_9987,N_8802);
nor U10962 (N_10962,N_9666,N_9251);
nand U10963 (N_10963,N_9862,N_9246);
and U10964 (N_10964,N_9763,N_9047);
nor U10965 (N_10965,N_9761,N_9083);
xnor U10966 (N_10966,N_8837,N_8979);
xnor U10967 (N_10967,N_8861,N_9212);
xor U10968 (N_10968,N_8801,N_8881);
and U10969 (N_10969,N_9498,N_8943);
and U10970 (N_10970,N_8832,N_9556);
nand U10971 (N_10971,N_9822,N_8943);
nand U10972 (N_10972,N_9607,N_9250);
xnor U10973 (N_10973,N_9753,N_9182);
nand U10974 (N_10974,N_9626,N_9113);
nor U10975 (N_10975,N_9156,N_9945);
nand U10976 (N_10976,N_9228,N_9282);
xor U10977 (N_10977,N_9866,N_9884);
and U10978 (N_10978,N_9962,N_9793);
or U10979 (N_10979,N_9642,N_9587);
nor U10980 (N_10980,N_9789,N_9484);
nor U10981 (N_10981,N_9005,N_8855);
xnor U10982 (N_10982,N_9165,N_9748);
and U10983 (N_10983,N_9449,N_9371);
nand U10984 (N_10984,N_8897,N_9228);
xnor U10985 (N_10985,N_9940,N_9096);
or U10986 (N_10986,N_9028,N_9906);
or U10987 (N_10987,N_9404,N_9515);
nor U10988 (N_10988,N_8810,N_9754);
xnor U10989 (N_10989,N_9437,N_9815);
nor U10990 (N_10990,N_9528,N_9293);
and U10991 (N_10991,N_8959,N_9744);
or U10992 (N_10992,N_9162,N_8937);
and U10993 (N_10993,N_9061,N_9551);
or U10994 (N_10994,N_9766,N_9551);
nand U10995 (N_10995,N_9867,N_9551);
nor U10996 (N_10996,N_9600,N_9534);
or U10997 (N_10997,N_9270,N_9017);
nand U10998 (N_10998,N_9223,N_9814);
nor U10999 (N_10999,N_9496,N_9440);
and U11000 (N_11000,N_8823,N_8960);
or U11001 (N_11001,N_8902,N_9208);
nor U11002 (N_11002,N_9208,N_9040);
and U11003 (N_11003,N_8861,N_8817);
or U11004 (N_11004,N_8995,N_9626);
nor U11005 (N_11005,N_9406,N_9768);
or U11006 (N_11006,N_9038,N_9909);
or U11007 (N_11007,N_9963,N_9511);
nor U11008 (N_11008,N_9741,N_9445);
nor U11009 (N_11009,N_9656,N_8858);
nand U11010 (N_11010,N_9542,N_9736);
xor U11011 (N_11011,N_9733,N_9285);
nor U11012 (N_11012,N_9761,N_9794);
and U11013 (N_11013,N_9166,N_9874);
and U11014 (N_11014,N_9713,N_8858);
nor U11015 (N_11015,N_9421,N_9406);
xnor U11016 (N_11016,N_9217,N_9822);
nor U11017 (N_11017,N_9525,N_8820);
xor U11018 (N_11018,N_9643,N_9817);
and U11019 (N_11019,N_9850,N_9063);
or U11020 (N_11020,N_9289,N_9621);
nand U11021 (N_11021,N_9631,N_9171);
or U11022 (N_11022,N_9928,N_9717);
or U11023 (N_11023,N_9613,N_8778);
nor U11024 (N_11024,N_9810,N_9062);
or U11025 (N_11025,N_9164,N_9433);
nor U11026 (N_11026,N_9873,N_9270);
or U11027 (N_11027,N_8837,N_9521);
nand U11028 (N_11028,N_9625,N_8937);
xor U11029 (N_11029,N_9076,N_9701);
nor U11030 (N_11030,N_9484,N_9606);
nand U11031 (N_11031,N_9321,N_8909);
nand U11032 (N_11032,N_9412,N_9353);
nand U11033 (N_11033,N_9955,N_9903);
or U11034 (N_11034,N_9625,N_8829);
nor U11035 (N_11035,N_9529,N_9555);
xor U11036 (N_11036,N_9067,N_9723);
xor U11037 (N_11037,N_9778,N_9010);
nand U11038 (N_11038,N_9454,N_9190);
nand U11039 (N_11039,N_9594,N_9933);
xor U11040 (N_11040,N_9326,N_8764);
xor U11041 (N_11041,N_9999,N_9161);
or U11042 (N_11042,N_9730,N_9404);
nand U11043 (N_11043,N_9411,N_9629);
and U11044 (N_11044,N_8775,N_9095);
nand U11045 (N_11045,N_9573,N_9767);
or U11046 (N_11046,N_9116,N_9730);
nand U11047 (N_11047,N_9726,N_9858);
nand U11048 (N_11048,N_9852,N_8804);
nor U11049 (N_11049,N_9416,N_9828);
and U11050 (N_11050,N_9024,N_9028);
or U11051 (N_11051,N_9423,N_9828);
or U11052 (N_11052,N_9669,N_9705);
xor U11053 (N_11053,N_9389,N_9026);
nand U11054 (N_11054,N_9194,N_9897);
nor U11055 (N_11055,N_9697,N_9873);
nand U11056 (N_11056,N_8785,N_9044);
nor U11057 (N_11057,N_8893,N_9215);
or U11058 (N_11058,N_9650,N_9992);
nand U11059 (N_11059,N_9115,N_8889);
and U11060 (N_11060,N_9331,N_9815);
or U11061 (N_11061,N_9138,N_9794);
or U11062 (N_11062,N_8995,N_9926);
nand U11063 (N_11063,N_9390,N_8973);
nor U11064 (N_11064,N_9450,N_9629);
nor U11065 (N_11065,N_9167,N_9247);
nand U11066 (N_11066,N_9805,N_9019);
nand U11067 (N_11067,N_8821,N_9636);
and U11068 (N_11068,N_8919,N_9306);
or U11069 (N_11069,N_9907,N_9340);
nor U11070 (N_11070,N_9969,N_9147);
nand U11071 (N_11071,N_9365,N_9725);
or U11072 (N_11072,N_8932,N_9668);
or U11073 (N_11073,N_8914,N_9530);
nor U11074 (N_11074,N_8799,N_9275);
nand U11075 (N_11075,N_8839,N_8863);
and U11076 (N_11076,N_8963,N_9333);
and U11077 (N_11077,N_8872,N_9693);
and U11078 (N_11078,N_9622,N_9996);
xnor U11079 (N_11079,N_9761,N_9746);
or U11080 (N_11080,N_9123,N_8992);
xnor U11081 (N_11081,N_8817,N_9926);
and U11082 (N_11082,N_9167,N_9145);
nor U11083 (N_11083,N_9856,N_9396);
nor U11084 (N_11084,N_9123,N_9822);
nor U11085 (N_11085,N_9384,N_9973);
nor U11086 (N_11086,N_9945,N_8847);
and U11087 (N_11087,N_9355,N_9757);
and U11088 (N_11088,N_9475,N_9768);
xnor U11089 (N_11089,N_9463,N_9506);
and U11090 (N_11090,N_9252,N_9204);
nor U11091 (N_11091,N_9778,N_9707);
and U11092 (N_11092,N_9333,N_8888);
and U11093 (N_11093,N_9502,N_9476);
or U11094 (N_11094,N_9864,N_9256);
and U11095 (N_11095,N_9601,N_9738);
xnor U11096 (N_11096,N_9545,N_9420);
xor U11097 (N_11097,N_9558,N_9251);
and U11098 (N_11098,N_9805,N_9621);
and U11099 (N_11099,N_9391,N_9513);
and U11100 (N_11100,N_9713,N_9678);
and U11101 (N_11101,N_9454,N_9774);
nor U11102 (N_11102,N_9704,N_9762);
or U11103 (N_11103,N_9458,N_9328);
nand U11104 (N_11104,N_9550,N_9618);
xor U11105 (N_11105,N_9557,N_8843);
and U11106 (N_11106,N_9625,N_8938);
nor U11107 (N_11107,N_9437,N_9897);
and U11108 (N_11108,N_8893,N_8896);
and U11109 (N_11109,N_9438,N_9868);
nand U11110 (N_11110,N_9889,N_8928);
nor U11111 (N_11111,N_9237,N_9055);
nor U11112 (N_11112,N_9874,N_8787);
or U11113 (N_11113,N_9546,N_9718);
or U11114 (N_11114,N_8830,N_9127);
or U11115 (N_11115,N_9814,N_9295);
xor U11116 (N_11116,N_9505,N_8889);
and U11117 (N_11117,N_9337,N_9196);
or U11118 (N_11118,N_9818,N_9900);
and U11119 (N_11119,N_9882,N_8773);
nand U11120 (N_11120,N_9905,N_9092);
or U11121 (N_11121,N_8941,N_9683);
and U11122 (N_11122,N_9123,N_9455);
nor U11123 (N_11123,N_9999,N_9774);
xnor U11124 (N_11124,N_9660,N_9479);
and U11125 (N_11125,N_9999,N_9590);
nor U11126 (N_11126,N_8885,N_9970);
and U11127 (N_11127,N_9150,N_8750);
and U11128 (N_11128,N_9538,N_9261);
nor U11129 (N_11129,N_9698,N_9982);
xnor U11130 (N_11130,N_9783,N_9265);
nand U11131 (N_11131,N_9133,N_9126);
xnor U11132 (N_11132,N_9125,N_9933);
nor U11133 (N_11133,N_9357,N_8863);
xor U11134 (N_11134,N_9108,N_9447);
nand U11135 (N_11135,N_9575,N_9853);
nor U11136 (N_11136,N_9921,N_9121);
nand U11137 (N_11137,N_8818,N_8929);
nand U11138 (N_11138,N_9795,N_9159);
nand U11139 (N_11139,N_9407,N_8897);
or U11140 (N_11140,N_9019,N_9195);
or U11141 (N_11141,N_9484,N_9058);
nor U11142 (N_11142,N_9973,N_9520);
or U11143 (N_11143,N_9895,N_9405);
or U11144 (N_11144,N_9392,N_9580);
nor U11145 (N_11145,N_9576,N_9310);
xor U11146 (N_11146,N_9811,N_9757);
nand U11147 (N_11147,N_9922,N_9723);
or U11148 (N_11148,N_9403,N_9897);
or U11149 (N_11149,N_8969,N_9286);
nand U11150 (N_11150,N_9924,N_9544);
nand U11151 (N_11151,N_8835,N_9273);
nand U11152 (N_11152,N_9555,N_8840);
xnor U11153 (N_11153,N_9553,N_8896);
nand U11154 (N_11154,N_9270,N_9816);
and U11155 (N_11155,N_9892,N_9437);
nor U11156 (N_11156,N_9122,N_9499);
and U11157 (N_11157,N_9586,N_9193);
xor U11158 (N_11158,N_9552,N_8885);
and U11159 (N_11159,N_9774,N_9010);
and U11160 (N_11160,N_9370,N_9945);
xor U11161 (N_11161,N_9506,N_9921);
nor U11162 (N_11162,N_9808,N_9240);
nor U11163 (N_11163,N_9534,N_9539);
nand U11164 (N_11164,N_9267,N_9683);
or U11165 (N_11165,N_9448,N_9125);
xnor U11166 (N_11166,N_9928,N_9022);
nand U11167 (N_11167,N_8983,N_9248);
and U11168 (N_11168,N_9263,N_9763);
xnor U11169 (N_11169,N_9453,N_9893);
nor U11170 (N_11170,N_9184,N_9107);
and U11171 (N_11171,N_8897,N_9029);
nor U11172 (N_11172,N_9216,N_9960);
nor U11173 (N_11173,N_9201,N_9640);
xor U11174 (N_11174,N_9238,N_8967);
or U11175 (N_11175,N_9544,N_9307);
nor U11176 (N_11176,N_9578,N_9481);
and U11177 (N_11177,N_8947,N_9533);
or U11178 (N_11178,N_8969,N_9201);
nand U11179 (N_11179,N_8963,N_8769);
nor U11180 (N_11180,N_8921,N_8858);
xor U11181 (N_11181,N_8894,N_8815);
nand U11182 (N_11182,N_9596,N_9199);
and U11183 (N_11183,N_9547,N_9224);
and U11184 (N_11184,N_9876,N_9541);
and U11185 (N_11185,N_9089,N_9561);
nand U11186 (N_11186,N_9784,N_9439);
xnor U11187 (N_11187,N_9324,N_9008);
or U11188 (N_11188,N_9176,N_9966);
or U11189 (N_11189,N_8756,N_9537);
or U11190 (N_11190,N_9307,N_9477);
or U11191 (N_11191,N_9280,N_9075);
or U11192 (N_11192,N_9141,N_9657);
nor U11193 (N_11193,N_9826,N_9968);
nand U11194 (N_11194,N_8882,N_9004);
nand U11195 (N_11195,N_9181,N_9775);
xnor U11196 (N_11196,N_9561,N_9623);
and U11197 (N_11197,N_9680,N_9592);
nand U11198 (N_11198,N_9565,N_9831);
and U11199 (N_11199,N_9672,N_9230);
nor U11200 (N_11200,N_8826,N_9409);
or U11201 (N_11201,N_9218,N_8834);
nor U11202 (N_11202,N_8905,N_9808);
xor U11203 (N_11203,N_9597,N_9771);
xor U11204 (N_11204,N_8799,N_9626);
or U11205 (N_11205,N_8994,N_9126);
xor U11206 (N_11206,N_8774,N_9960);
xnor U11207 (N_11207,N_9190,N_9881);
and U11208 (N_11208,N_9955,N_9861);
and U11209 (N_11209,N_9371,N_9931);
nand U11210 (N_11210,N_9326,N_8936);
nand U11211 (N_11211,N_9954,N_8919);
or U11212 (N_11212,N_8802,N_9633);
xor U11213 (N_11213,N_8818,N_9536);
xnor U11214 (N_11214,N_9916,N_9661);
and U11215 (N_11215,N_9667,N_8977);
xor U11216 (N_11216,N_9813,N_9203);
nor U11217 (N_11217,N_9283,N_9128);
nand U11218 (N_11218,N_9883,N_9377);
or U11219 (N_11219,N_9917,N_9987);
nand U11220 (N_11220,N_9040,N_9430);
and U11221 (N_11221,N_9065,N_8917);
nor U11222 (N_11222,N_8949,N_9249);
xor U11223 (N_11223,N_9773,N_9510);
nand U11224 (N_11224,N_8977,N_9040);
nor U11225 (N_11225,N_8866,N_9043);
nor U11226 (N_11226,N_8972,N_9504);
and U11227 (N_11227,N_9281,N_9435);
nor U11228 (N_11228,N_9031,N_9442);
xnor U11229 (N_11229,N_9078,N_8760);
nor U11230 (N_11230,N_9207,N_9049);
nor U11231 (N_11231,N_8850,N_8947);
and U11232 (N_11232,N_9819,N_9961);
nor U11233 (N_11233,N_9361,N_8897);
nand U11234 (N_11234,N_9874,N_9666);
nor U11235 (N_11235,N_9602,N_9091);
nor U11236 (N_11236,N_9282,N_8806);
nand U11237 (N_11237,N_8806,N_9938);
and U11238 (N_11238,N_9600,N_9369);
nand U11239 (N_11239,N_9354,N_9278);
xnor U11240 (N_11240,N_9435,N_9613);
nor U11241 (N_11241,N_9895,N_9939);
or U11242 (N_11242,N_9559,N_9316);
and U11243 (N_11243,N_9679,N_9827);
and U11244 (N_11244,N_8983,N_8934);
or U11245 (N_11245,N_9380,N_9373);
and U11246 (N_11246,N_9413,N_9468);
and U11247 (N_11247,N_8893,N_9749);
and U11248 (N_11248,N_8920,N_8937);
and U11249 (N_11249,N_9553,N_9589);
xnor U11250 (N_11250,N_11152,N_10852);
and U11251 (N_11251,N_10166,N_11046);
nand U11252 (N_11252,N_10666,N_11148);
nor U11253 (N_11253,N_10264,N_10815);
and U11254 (N_11254,N_10114,N_10562);
nand U11255 (N_11255,N_10393,N_10828);
nor U11256 (N_11256,N_10418,N_11033);
or U11257 (N_11257,N_11070,N_10153);
nand U11258 (N_11258,N_10410,N_10040);
nand U11259 (N_11259,N_10122,N_10246);
nor U11260 (N_11260,N_11117,N_10078);
and U11261 (N_11261,N_10136,N_10521);
nor U11262 (N_11262,N_10889,N_10262);
or U11263 (N_11263,N_10454,N_10368);
xnor U11264 (N_11264,N_10660,N_10607);
xnor U11265 (N_11265,N_10425,N_10629);
nand U11266 (N_11266,N_10737,N_11111);
and U11267 (N_11267,N_10713,N_11059);
xor U11268 (N_11268,N_10198,N_10579);
nor U11269 (N_11269,N_11249,N_10907);
or U11270 (N_11270,N_11150,N_10447);
nand U11271 (N_11271,N_11040,N_10070);
xor U11272 (N_11272,N_11206,N_10398);
nand U11273 (N_11273,N_10000,N_10935);
or U11274 (N_11274,N_10848,N_10577);
nand U11275 (N_11275,N_10505,N_10496);
xnor U11276 (N_11276,N_10213,N_10271);
and U11277 (N_11277,N_11030,N_10309);
or U11278 (N_11278,N_10769,N_10144);
nand U11279 (N_11279,N_11051,N_10443);
xor U11280 (N_11280,N_10734,N_10911);
nor U11281 (N_11281,N_10707,N_11042);
xor U11282 (N_11282,N_10442,N_10975);
xnor U11283 (N_11283,N_10301,N_10155);
nand U11284 (N_11284,N_10093,N_10902);
or U11285 (N_11285,N_10958,N_10016);
nor U11286 (N_11286,N_10929,N_10132);
or U11287 (N_11287,N_11204,N_10874);
nor U11288 (N_11288,N_10576,N_11143);
and U11289 (N_11289,N_10850,N_11242);
xor U11290 (N_11290,N_10635,N_10998);
nor U11291 (N_11291,N_10719,N_11065);
xor U11292 (N_11292,N_10300,N_10677);
and U11293 (N_11293,N_10840,N_10401);
xnor U11294 (N_11294,N_10777,N_10940);
or U11295 (N_11295,N_11175,N_10408);
xnor U11296 (N_11296,N_11011,N_10849);
xnor U11297 (N_11297,N_10817,N_10133);
nor U11298 (N_11298,N_10383,N_10971);
and U11299 (N_11299,N_10129,N_10077);
or U11300 (N_11300,N_11220,N_10483);
and U11301 (N_11301,N_11158,N_10714);
and U11302 (N_11302,N_10786,N_10740);
xnor U11303 (N_11303,N_11137,N_11079);
nor U11304 (N_11304,N_10021,N_10382);
or U11305 (N_11305,N_10482,N_10915);
or U11306 (N_11306,N_10285,N_10330);
xor U11307 (N_11307,N_11008,N_11125);
nand U11308 (N_11308,N_10580,N_11201);
or U11309 (N_11309,N_10705,N_11044);
xor U11310 (N_11310,N_10112,N_10227);
nor U11311 (N_11311,N_10993,N_10168);
nor U11312 (N_11312,N_10015,N_10668);
or U11313 (N_11313,N_11060,N_10731);
nor U11314 (N_11314,N_10844,N_10258);
and U11315 (N_11315,N_10823,N_10716);
nor U11316 (N_11316,N_10363,N_10331);
or U11317 (N_11317,N_10634,N_10047);
xnor U11318 (N_11318,N_10266,N_11248);
xnor U11319 (N_11319,N_10180,N_11225);
or U11320 (N_11320,N_10515,N_10609);
or U11321 (N_11321,N_10488,N_10433);
or U11322 (N_11322,N_11166,N_10775);
and U11323 (N_11323,N_10657,N_10320);
or U11324 (N_11324,N_11050,N_11126);
xnor U11325 (N_11325,N_10241,N_10517);
xor U11326 (N_11326,N_10806,N_11012);
and U11327 (N_11327,N_11029,N_10696);
or U11328 (N_11328,N_10291,N_10995);
nand U11329 (N_11329,N_10834,N_10934);
and U11330 (N_11330,N_10767,N_10930);
or U11331 (N_11331,N_10319,N_10581);
or U11332 (N_11332,N_11239,N_10328);
nor U11333 (N_11333,N_10321,N_11192);
nand U11334 (N_11334,N_10768,N_10123);
xnor U11335 (N_11335,N_10392,N_11077);
and U11336 (N_11336,N_10141,N_10456);
nand U11337 (N_11337,N_10450,N_10394);
or U11338 (N_11338,N_10094,N_10989);
or U11339 (N_11339,N_10352,N_10182);
xor U11340 (N_11340,N_10207,N_10630);
nor U11341 (N_11341,N_10882,N_10599);
xnor U11342 (N_11342,N_10477,N_10898);
or U11343 (N_11343,N_10596,N_10396);
or U11344 (N_11344,N_10072,N_10640);
nor U11345 (N_11345,N_10350,N_11082);
or U11346 (N_11346,N_10551,N_10440);
nand U11347 (N_11347,N_10279,N_10073);
or U11348 (N_11348,N_10897,N_10825);
nor U11349 (N_11349,N_11089,N_11247);
nor U11350 (N_11350,N_10499,N_11216);
nand U11351 (N_11351,N_10561,N_10067);
and U11352 (N_11352,N_10507,N_10652);
xor U11353 (N_11353,N_11130,N_10868);
nor U11354 (N_11354,N_10520,N_10348);
nand U11355 (N_11355,N_10709,N_10049);
nor U11356 (N_11356,N_10495,N_10306);
or U11357 (N_11357,N_10895,N_11056);
nor U11358 (N_11358,N_10186,N_10616);
and U11359 (N_11359,N_10171,N_10472);
nand U11360 (N_11360,N_10608,N_10762);
nand U11361 (N_11361,N_10994,N_10687);
nand U11362 (N_11362,N_10504,N_10980);
nor U11363 (N_11363,N_10999,N_10455);
xnor U11364 (N_11364,N_10727,N_10358);
nand U11365 (N_11365,N_10741,N_10905);
nand U11366 (N_11366,N_10923,N_10283);
or U11367 (N_11367,N_10604,N_10754);
nand U11368 (N_11368,N_10458,N_11103);
and U11369 (N_11369,N_10359,N_10005);
or U11370 (N_11370,N_10624,N_10978);
or U11371 (N_11371,N_10872,N_10548);
nor U11372 (N_11372,N_10397,N_10778);
nor U11373 (N_11373,N_11146,N_11240);
or U11374 (N_11374,N_10222,N_11107);
nor U11375 (N_11375,N_10941,N_11189);
and U11376 (N_11376,N_11018,N_10221);
nor U11377 (N_11377,N_10289,N_10829);
nand U11378 (N_11378,N_10298,N_10617);
or U11379 (N_11379,N_10263,N_10431);
or U11380 (N_11380,N_11246,N_10802);
xor U11381 (N_11381,N_10625,N_10231);
and U11382 (N_11382,N_10406,N_10374);
nor U11383 (N_11383,N_10583,N_10063);
and U11384 (N_11384,N_10386,N_10726);
xnor U11385 (N_11385,N_11109,N_10412);
or U11386 (N_11386,N_10295,N_10402);
nand U11387 (N_11387,N_10312,N_11156);
nand U11388 (N_11388,N_10772,N_10343);
or U11389 (N_11389,N_11088,N_10535);
nor U11390 (N_11390,N_11217,N_10908);
nand U11391 (N_11391,N_10627,N_10225);
or U11392 (N_11392,N_11177,N_10025);
xnor U11393 (N_11393,N_10034,N_10066);
nand U11394 (N_11394,N_10332,N_10195);
nor U11395 (N_11395,N_11154,N_10335);
nor U11396 (N_11396,N_10918,N_10739);
or U11397 (N_11397,N_10459,N_11147);
and U11398 (N_11398,N_10228,N_10883);
nand U11399 (N_11399,N_10826,N_10269);
xor U11400 (N_11400,N_10595,N_10038);
or U11401 (N_11401,N_11232,N_10623);
xor U11402 (N_11402,N_10602,N_10145);
xor U11403 (N_11403,N_10710,N_10818);
nand U11404 (N_11404,N_11049,N_11184);
xnor U11405 (N_11405,N_10774,N_11035);
xnor U11406 (N_11406,N_10513,N_11032);
nor U11407 (N_11407,N_10871,N_11087);
nor U11408 (N_11408,N_10367,N_11006);
nand U11409 (N_11409,N_10165,N_10765);
and U11410 (N_11410,N_10916,N_10187);
xor U11411 (N_11411,N_10653,N_10003);
and U11412 (N_11412,N_10196,N_11074);
and U11413 (N_11413,N_10749,N_10858);
xnor U11414 (N_11414,N_11183,N_10791);
and U11415 (N_11415,N_11119,N_10528);
or U11416 (N_11416,N_11134,N_11023);
and U11417 (N_11417,N_10120,N_10906);
and U11418 (N_11418,N_11172,N_11243);
xor U11419 (N_11419,N_10091,N_11066);
and U11420 (N_11420,N_10208,N_11025);
and U11421 (N_11421,N_11027,N_10371);
xor U11422 (N_11422,N_10944,N_10805);
or U11423 (N_11423,N_10886,N_10031);
nor U11424 (N_11424,N_10534,N_10681);
xnor U11425 (N_11425,N_11004,N_10065);
and U11426 (N_11426,N_10743,N_10830);
xor U11427 (N_11427,N_11017,N_10820);
and U11428 (N_11428,N_10365,N_11054);
xor U11429 (N_11429,N_10574,N_10983);
nor U11430 (N_11430,N_10282,N_10113);
nand U11431 (N_11431,N_10856,N_10245);
or U11432 (N_11432,N_10920,N_10092);
or U11433 (N_11433,N_10685,N_10914);
nor U11434 (N_11434,N_10899,N_10554);
or U11435 (N_11435,N_10135,N_10011);
or U11436 (N_11436,N_10215,N_10096);
xnor U11437 (N_11437,N_10981,N_10233);
or U11438 (N_11438,N_11132,N_10502);
nor U11439 (N_11439,N_10189,N_10267);
xnor U11440 (N_11440,N_10509,N_10277);
or U11441 (N_11441,N_10827,N_11028);
nor U11442 (N_11442,N_10248,N_10865);
nand U11443 (N_11443,N_10061,N_11120);
nor U11444 (N_11444,N_10703,N_10351);
and U11445 (N_11445,N_10493,N_10342);
nand U11446 (N_11446,N_10952,N_10140);
and U11447 (N_11447,N_11036,N_10308);
nand U11448 (N_11448,N_10471,N_11064);
nor U11449 (N_11449,N_11047,N_10861);
and U11450 (N_11450,N_10302,N_10002);
nor U11451 (N_11451,N_11139,N_10892);
and U11452 (N_11452,N_10972,N_10316);
nand U11453 (N_11453,N_11149,N_10591);
nor U11454 (N_11454,N_10966,N_11212);
xor U11455 (N_11455,N_10413,N_10256);
and U11456 (N_11456,N_11171,N_10014);
nor U11457 (N_11457,N_10953,N_11092);
nor U11458 (N_11458,N_10621,N_10671);
nand U11459 (N_11459,N_10232,N_10950);
nor U11460 (N_11460,N_10807,N_10299);
and U11461 (N_11461,N_10119,N_10212);
xor U11462 (N_11462,N_10226,N_10795);
and U11463 (N_11463,N_10148,N_10322);
nor U11464 (N_11464,N_10730,N_10023);
xnor U11465 (N_11465,N_10990,N_11179);
xor U11466 (N_11466,N_10587,N_10121);
or U11467 (N_11467,N_10880,N_11245);
nor U11468 (N_11468,N_10116,N_10891);
xnor U11469 (N_11469,N_10400,N_10525);
nor U11470 (N_11470,N_10833,N_10109);
nor U11471 (N_11471,N_10613,N_10467);
nand U11472 (N_11472,N_10259,N_10388);
nor U11473 (N_11473,N_11019,N_10679);
nor U11474 (N_11474,N_10542,N_10427);
or U11475 (N_11475,N_10252,N_10188);
and U11476 (N_11476,N_10690,N_10434);
nor U11477 (N_11477,N_10028,N_10030);
and U11478 (N_11478,N_10887,N_10516);
nand U11479 (N_11479,N_11221,N_10361);
xnor U11480 (N_11480,N_10736,N_10503);
nand U11481 (N_11481,N_10404,N_11101);
nand U11482 (N_11482,N_10029,N_10179);
or U11483 (N_11483,N_11191,N_11007);
and U11484 (N_11484,N_10466,N_10824);
or U11485 (N_11485,N_10530,N_10700);
or U11486 (N_11486,N_11169,N_11112);
and U11487 (N_11487,N_10430,N_10662);
nand U11488 (N_11488,N_10378,N_10728);
and U11489 (N_11489,N_10451,N_11159);
xor U11490 (N_11490,N_10890,N_10519);
or U11491 (N_11491,N_10288,N_10474);
and U11492 (N_11492,N_10606,N_10103);
or U11493 (N_11493,N_10732,N_10346);
xnor U11494 (N_11494,N_10162,N_10573);
xor U11495 (N_11495,N_10315,N_10610);
nand U11496 (N_11496,N_10879,N_10480);
nand U11497 (N_11497,N_10968,N_10976);
nand U11498 (N_11498,N_10645,N_11157);
xor U11499 (N_11499,N_10748,N_10088);
nor U11500 (N_11500,N_10711,N_10755);
xor U11501 (N_11501,N_10810,N_10062);
or U11502 (N_11502,N_11118,N_10564);
xnor U11503 (N_11503,N_10747,N_10462);
nor U11504 (N_11504,N_10366,N_10476);
or U11505 (N_11505,N_11133,N_11224);
and U11506 (N_11506,N_10997,N_10760);
xor U11507 (N_11507,N_10018,N_10684);
or U11508 (N_11508,N_10831,N_10694);
nor U11509 (N_11509,N_10536,N_10074);
xnor U11510 (N_11510,N_11005,N_10903);
or U11511 (N_11511,N_10647,N_10203);
nor U11512 (N_11512,N_10860,N_10142);
or U11513 (N_11513,N_10855,N_10704);
or U11514 (N_11514,N_10523,N_10039);
nand U11515 (N_11515,N_11009,N_10571);
and U11516 (N_11516,N_11227,N_10919);
or U11517 (N_11517,N_10446,N_11197);
or U11518 (N_11518,N_10105,N_11188);
nor U11519 (N_11519,N_10384,N_10152);
nand U11520 (N_11520,N_10185,N_10261);
and U11521 (N_11521,N_10723,N_10866);
nor U11522 (N_11522,N_10742,N_10565);
and U11523 (N_11523,N_10927,N_10364);
xnor U11524 (N_11524,N_11003,N_10275);
or U11525 (N_11525,N_10293,N_11160);
xnor U11526 (N_11526,N_10052,N_11039);
xnor U11527 (N_11527,N_10033,N_10104);
or U11528 (N_11528,N_10798,N_10082);
and U11529 (N_11529,N_10893,N_10835);
or U11530 (N_11530,N_10559,N_10071);
nand U11531 (N_11531,N_10991,N_10644);
nand U11532 (N_11532,N_10421,N_10812);
nor U11533 (N_11533,N_10804,N_10598);
xor U11534 (N_11534,N_10729,N_10485);
xor U11535 (N_11535,N_10572,N_10310);
or U11536 (N_11536,N_10799,N_10510);
nor U11537 (N_11537,N_10324,N_10721);
and U11538 (N_11538,N_11213,N_10201);
xnor U11539 (N_11539,N_10008,N_11096);
and U11540 (N_11540,N_10379,N_10566);
and U11541 (N_11541,N_11161,N_10611);
or U11542 (N_11542,N_10593,N_10284);
and U11543 (N_11543,N_10193,N_10238);
nor U11544 (N_11544,N_11108,N_10797);
nand U11545 (N_11545,N_11097,N_10819);
and U11546 (N_11546,N_10184,N_10390);
nor U11547 (N_11547,N_10060,N_11145);
nand U11548 (N_11548,N_10270,N_10753);
or U11549 (N_11549,N_10733,N_10963);
and U11550 (N_11550,N_10912,N_11153);
or U11551 (N_11551,N_10955,N_10842);
or U11552 (N_11552,N_10313,N_10712);
or U11553 (N_11553,N_10537,N_10646);
and U11554 (N_11554,N_11095,N_10042);
nand U11555 (N_11555,N_10009,N_10389);
xnor U11556 (N_11556,N_10682,N_10514);
nand U11557 (N_11557,N_11078,N_10859);
or U11558 (N_11558,N_10095,N_10377);
nand U11559 (N_11559,N_10800,N_10854);
or U11560 (N_11560,N_10917,N_11142);
nand U11561 (N_11561,N_10338,N_10385);
nor U11562 (N_11562,N_10896,N_10235);
nand U11563 (N_11563,N_10154,N_10048);
nand U11564 (N_11564,N_10290,N_10924);
nor U11565 (N_11565,N_10839,N_11098);
nor U11566 (N_11566,N_10957,N_10575);
or U11567 (N_11567,N_10169,N_11045);
nand U11568 (N_11568,N_10676,N_10656);
xor U11569 (N_11569,N_10424,N_10437);
nand U11570 (N_11570,N_10090,N_11053);
xnor U11571 (N_11571,N_10027,N_10294);
nor U11572 (N_11572,N_10612,N_10803);
nor U11573 (N_11573,N_11084,N_10761);
nor U11574 (N_11574,N_10234,N_10813);
xnor U11575 (N_11575,N_10395,N_10636);
xnor U11576 (N_11576,N_11002,N_10010);
and U11577 (N_11577,N_10544,N_10639);
nor U11578 (N_11578,N_10560,N_11072);
nand U11579 (N_11579,N_10438,N_10680);
or U11580 (N_11580,N_10670,N_10128);
and U11581 (N_11581,N_10307,N_10329);
or U11582 (N_11582,N_11076,N_10718);
or U11583 (N_11583,N_10555,N_10278);
or U11584 (N_11584,N_10550,N_10100);
xnor U11585 (N_11585,N_10445,N_10349);
nor U11586 (N_11586,N_10181,N_10419);
and U11587 (N_11587,N_10875,N_10304);
xor U11588 (N_11588,N_10257,N_10691);
nor U11589 (N_11589,N_11106,N_11235);
nand U11590 (N_11590,N_11193,N_10921);
or U11591 (N_11591,N_10672,N_10191);
xnor U11592 (N_11592,N_10925,N_10006);
or U11593 (N_11593,N_10337,N_10947);
xnor U11594 (N_11594,N_10594,N_11124);
and U11595 (N_11595,N_10904,N_10693);
nor U11596 (N_11596,N_10372,N_11187);
nor U11597 (N_11597,N_10417,N_10318);
and U11598 (N_11598,N_10603,N_10655);
nor U11599 (N_11599,N_11200,N_10878);
xor U11600 (N_11600,N_10273,N_10541);
and U11601 (N_11601,N_10585,N_10578);
nand U11602 (N_11602,N_11163,N_10001);
nand U11603 (N_11603,N_10230,N_10864);
xor U11604 (N_11604,N_11020,N_10420);
nand U11605 (N_11605,N_10176,N_10847);
xnor U11606 (N_11606,N_11016,N_10036);
and U11607 (N_11607,N_10744,N_11211);
and U11608 (N_11608,N_10757,N_10763);
or U11609 (N_11609,N_10926,N_11144);
and U11610 (N_11610,N_11001,N_10956);
xor U11611 (N_11611,N_10965,N_10522);
xnor U11612 (N_11612,N_10058,N_10853);
nand U11613 (N_11613,N_10317,N_10706);
nand U11614 (N_11614,N_10881,N_11122);
and U11615 (N_11615,N_10081,N_10843);
nor U11616 (N_11616,N_10177,N_10464);
or U11617 (N_11617,N_10945,N_10083);
nor U11618 (N_11618,N_10174,N_11127);
nand U11619 (N_11619,N_11218,N_10012);
nor U11620 (N_11620,N_10461,N_10518);
nand U11621 (N_11621,N_10143,N_10910);
nand U11622 (N_11622,N_10097,N_10111);
nor U11623 (N_11623,N_10862,N_10751);
or U11624 (N_11624,N_10068,N_10650);
nor U11625 (N_11625,N_11062,N_10970);
nand U11626 (N_11626,N_10490,N_10592);
and U11627 (N_11627,N_10987,N_10452);
nand U11628 (N_11628,N_10151,N_10876);
xnor U11629 (N_11629,N_10399,N_10381);
or U11630 (N_11630,N_10932,N_10689);
or U11631 (N_11631,N_10867,N_11010);
xnor U11632 (N_11632,N_10563,N_10552);
nand U11633 (N_11633,N_10167,N_11207);
and U11634 (N_11634,N_10558,N_10199);
xor U11635 (N_11635,N_10590,N_11234);
and U11636 (N_11636,N_10415,N_10722);
nand U11637 (N_11637,N_10954,N_10501);
and U11638 (N_11638,N_11090,N_10409);
or U11639 (N_11639,N_10979,N_10131);
or U11640 (N_11640,N_10615,N_10701);
or U11641 (N_11641,N_10928,N_10759);
nand U11642 (N_11642,N_11026,N_11052);
and U11643 (N_11643,N_10909,N_10255);
or U11644 (N_11644,N_10407,N_10922);
or U11645 (N_11645,N_10345,N_10137);
and U11646 (N_11646,N_11091,N_10391);
nand U11647 (N_11647,N_10297,N_10715);
and U11648 (N_11648,N_10210,N_11174);
and U11649 (N_11649,N_10673,N_10202);
nor U11650 (N_11650,N_10139,N_10387);
nand U11651 (N_11651,N_10216,N_10223);
or U11652 (N_11652,N_10512,N_10138);
xor U11653 (N_11653,N_10484,N_10832);
nand U11654 (N_11654,N_11136,N_10106);
nor U11655 (N_11655,N_10046,N_11190);
nand U11656 (N_11656,N_10977,N_10347);
nor U11657 (N_11657,N_11013,N_10355);
nor U11658 (N_11658,N_10549,N_10984);
or U11659 (N_11659,N_10089,N_10822);
and U11660 (N_11660,N_10962,N_10695);
xnor U11661 (N_11661,N_11182,N_10821);
and U11662 (N_11662,N_10781,N_10600);
nor U11663 (N_11663,N_11055,N_10236);
xor U11664 (N_11664,N_10055,N_10683);
xnor U11665 (N_11665,N_10531,N_10738);
nand U11666 (N_11666,N_10626,N_10790);
nand U11667 (N_11667,N_10200,N_11233);
xor U11668 (N_11668,N_10344,N_10533);
nor U11669 (N_11669,N_11000,N_10857);
nand U11670 (N_11670,N_10532,N_10057);
or U11671 (N_11671,N_10086,N_10175);
and U11672 (N_11672,N_11181,N_11205);
or U11673 (N_11673,N_10816,N_10362);
xor U11674 (N_11674,N_10087,N_10481);
nand U11675 (N_11675,N_11194,N_10524);
or U11676 (N_11676,N_10931,N_11170);
and U11677 (N_11677,N_10638,N_10661);
nor U11678 (N_11678,N_10117,N_10149);
xnor U11679 (N_11679,N_10435,N_11229);
or U11680 (N_11680,N_10107,N_10453);
and U11681 (N_11681,N_10240,N_10678);
nor U11682 (N_11682,N_10894,N_11244);
and U11683 (N_11683,N_10973,N_10292);
xor U11684 (N_11684,N_10588,N_11100);
nor U11685 (N_11685,N_11099,N_10527);
or U11686 (N_11686,N_10782,N_11178);
and U11687 (N_11687,N_11203,N_10569);
nor U11688 (N_11688,N_10281,N_10101);
nor U11689 (N_11689,N_10156,N_10674);
or U11690 (N_11690,N_10220,N_11105);
and U11691 (N_11691,N_10641,N_11024);
and U11692 (N_11692,N_10584,N_10885);
xnor U11693 (N_11693,N_10080,N_10218);
and U11694 (N_11694,N_10664,N_10500);
nand U11695 (N_11695,N_11162,N_10163);
nor U11696 (N_11696,N_11165,N_10796);
xnor U11697 (N_11697,N_10102,N_10597);
nor U11698 (N_11698,N_11073,N_11061);
and U11699 (N_11699,N_11031,N_10076);
xor U11700 (N_11700,N_10568,N_11080);
xnor U11701 (N_11701,N_10913,N_10247);
xnor U11702 (N_11702,N_11114,N_10369);
nor U11703 (N_11703,N_10988,N_10750);
and U11704 (N_11704,N_10115,N_10637);
and U11705 (N_11705,N_10614,N_10967);
xnor U11706 (N_11706,N_10992,N_10339);
and U11707 (N_11707,N_10020,N_10814);
nor U11708 (N_11708,N_11135,N_10004);
xnor U11709 (N_11709,N_10444,N_10631);
xor U11710 (N_11710,N_10974,N_11083);
and U11711 (N_11711,N_10205,N_10134);
nor U11712 (N_11712,N_10422,N_10720);
nand U11713 (N_11713,N_10801,N_11021);
nand U11714 (N_11714,N_10041,N_11164);
xnor U11715 (N_11715,N_10697,N_11071);
nand U11716 (N_11716,N_10869,N_10229);
xor U11717 (N_11717,N_10570,N_10209);
and U11718 (N_11718,N_10305,N_11173);
nand U11719 (N_11719,N_11104,N_10669);
or U11720 (N_11720,N_10771,N_11129);
xor U11721 (N_11721,N_11214,N_10756);
nand U11722 (N_11722,N_11043,N_10013);
xnor U11723 (N_11723,N_10037,N_11186);
and U11724 (N_11724,N_11196,N_10888);
xnor U11725 (N_11725,N_10628,N_10237);
and U11726 (N_11726,N_10448,N_10665);
and U11727 (N_11727,N_10836,N_10900);
and U11728 (N_11728,N_10160,N_11176);
or U11729 (N_11729,N_10242,N_10054);
and U11730 (N_11730,N_10649,N_10035);
nand U11731 (N_11731,N_10632,N_10863);
nor U11732 (N_11732,N_10045,N_11075);
xnor U11733 (N_11733,N_10959,N_10556);
xnor U11734 (N_11734,N_10428,N_10375);
and U11735 (N_11735,N_10125,N_10582);
xnor U11736 (N_11736,N_10758,N_10260);
xnor U11737 (N_11737,N_11102,N_11022);
nand U11738 (N_11738,N_11048,N_10708);
nand U11739 (N_11739,N_11069,N_10633);
xor U11740 (N_11740,N_10296,N_10019);
nand U11741 (N_11741,N_11210,N_11241);
and U11742 (N_11742,N_10426,N_10026);
or U11743 (N_11743,N_10688,N_11168);
xnor U11744 (N_11744,N_10079,N_10780);
nand U11745 (N_11745,N_10274,N_11113);
and U11746 (N_11746,N_10118,N_10024);
or U11747 (N_11747,N_10075,N_10648);
nand U11748 (N_11748,N_10197,N_10779);
or U11749 (N_11749,N_10960,N_10475);
xor U11750 (N_11750,N_10792,N_10845);
and U11751 (N_11751,N_10124,N_10334);
xor U11752 (N_11752,N_10050,N_10376);
xnor U11753 (N_11753,N_10746,N_10098);
xor U11754 (N_11754,N_10964,N_10340);
and U11755 (N_11755,N_10311,N_11121);
or U11756 (N_11756,N_10949,N_11086);
or U11757 (N_11757,N_11081,N_10099);
and U11758 (N_11758,N_10468,N_10414);
and U11759 (N_11759,N_10370,N_11219);
nor U11760 (N_11760,N_10794,N_10439);
xor U11761 (N_11761,N_10314,N_10353);
xor U11762 (N_11762,N_10251,N_10686);
xor U11763 (N_11763,N_10429,N_10276);
nand U11764 (N_11764,N_10333,N_11208);
nand U11765 (N_11765,N_10360,N_11068);
nand U11766 (N_11766,N_10272,N_10056);
nand U11767 (N_11767,N_10059,N_11038);
xor U11768 (N_11768,N_10996,N_11094);
nor U11769 (N_11769,N_10619,N_10405);
and U11770 (N_11770,N_10497,N_11202);
and U11771 (N_11771,N_10735,N_10498);
nand U11772 (N_11772,N_10489,N_10543);
nor U11773 (N_11773,N_10546,N_11058);
xnor U11774 (N_11774,N_10547,N_10667);
nand U11775 (N_11775,N_10942,N_10506);
nor U11776 (N_11776,N_10933,N_10557);
or U11777 (N_11777,N_11140,N_11155);
nand U11778 (N_11778,N_11151,N_10752);
or U11779 (N_11779,N_11014,N_11215);
and U11780 (N_11780,N_11238,N_10253);
nand U11781 (N_11781,N_10449,N_10146);
xnor U11782 (N_11782,N_11195,N_11128);
or U11783 (N_11783,N_10206,N_10717);
nand U11784 (N_11784,N_10161,N_10357);
or U11785 (N_11785,N_10511,N_10130);
xor U11786 (N_11786,N_10873,N_10250);
nand U11787 (N_11787,N_10380,N_10841);
nor U11788 (N_11788,N_10441,N_10007);
nor U11789 (N_11789,N_10494,N_10937);
xor U11790 (N_11790,N_10287,N_10659);
or U11791 (N_11791,N_10110,N_10173);
nand U11792 (N_11792,N_11199,N_10939);
or U11793 (N_11793,N_10190,N_10784);
xnor U11794 (N_11794,N_10423,N_10526);
or U11795 (N_11795,N_10508,N_10725);
xor U11796 (N_11796,N_10044,N_10159);
nand U11797 (N_11797,N_10985,N_10809);
and U11798 (N_11798,N_10032,N_10479);
or U11799 (N_11799,N_10457,N_10326);
or U11800 (N_11800,N_11115,N_10538);
xnor U11801 (N_11801,N_10053,N_10356);
nor U11802 (N_11802,N_11110,N_10465);
nand U11803 (N_11803,N_10460,N_10268);
and U11804 (N_11804,N_10051,N_10663);
nand U11805 (N_11805,N_10192,N_10325);
or U11806 (N_11806,N_10788,N_10303);
and U11807 (N_11807,N_11167,N_10172);
or U11808 (N_11808,N_10463,N_10127);
nor U11809 (N_11809,N_10787,N_10214);
nand U11810 (N_11810,N_10157,N_10354);
and U11811 (N_11811,N_10764,N_10766);
nor U11812 (N_11812,N_11041,N_10492);
nor U11813 (N_11813,N_10487,N_10219);
or U11814 (N_11814,N_10884,N_10618);
and U11815 (N_11815,N_10589,N_11180);
nor U11816 (N_11816,N_10545,N_11037);
and U11817 (N_11817,N_10491,N_10938);
nor U11818 (N_11818,N_11034,N_10478);
xor U11819 (N_11819,N_10783,N_11230);
xnor U11820 (N_11820,N_10808,N_10951);
or U11821 (N_11821,N_10211,N_11116);
and U11822 (N_11822,N_11063,N_10473);
and U11823 (N_11823,N_10108,N_10651);
or U11824 (N_11824,N_10776,N_11093);
xor U11825 (N_11825,N_10323,N_11226);
nand U11826 (N_11826,N_10789,N_10553);
xor U11827 (N_11827,N_10702,N_10017);
and U11828 (N_11828,N_10064,N_10901);
nor U11829 (N_11829,N_10770,N_10982);
and U11830 (N_11830,N_10341,N_10403);
xor U11831 (N_11831,N_10658,N_10851);
nand U11832 (N_11832,N_10986,N_10943);
xnor U11833 (N_11833,N_10336,N_10043);
nand U11834 (N_11834,N_10254,N_11015);
nor U11835 (N_11835,N_10126,N_10373);
nand U11836 (N_11836,N_11209,N_10793);
or U11837 (N_11837,N_10773,N_10158);
xor U11838 (N_11838,N_10265,N_10280);
nor U11839 (N_11839,N_11223,N_10969);
xnor U11840 (N_11840,N_10601,N_10470);
nand U11841 (N_11841,N_11067,N_11236);
xor U11842 (N_11842,N_10948,N_10436);
and U11843 (N_11843,N_10084,N_10692);
nor U11844 (N_11844,N_10085,N_10877);
or U11845 (N_11845,N_10654,N_10217);
or U11846 (N_11846,N_10069,N_10838);
nand U11847 (N_11847,N_10224,N_10785);
or U11848 (N_11848,N_10243,N_10170);
or U11849 (N_11849,N_11185,N_10622);
nand U11850 (N_11850,N_10164,N_11231);
or U11851 (N_11851,N_10620,N_11123);
xor U11852 (N_11852,N_10567,N_10432);
or U11853 (N_11853,N_10249,N_10416);
and U11854 (N_11854,N_10469,N_10605);
xor U11855 (N_11855,N_10642,N_11228);
nor U11856 (N_11856,N_10327,N_11237);
and U11857 (N_11857,N_11131,N_11141);
nand U11858 (N_11858,N_10239,N_11222);
nand U11859 (N_11859,N_10150,N_10846);
nor U11860 (N_11860,N_10486,N_10147);
nand U11861 (N_11861,N_10540,N_10698);
nand U11862 (N_11862,N_10811,N_10022);
and U11863 (N_11863,N_10643,N_10675);
nand U11864 (N_11864,N_11057,N_10586);
and U11865 (N_11865,N_10961,N_10539);
and U11866 (N_11866,N_10178,N_10411);
nand U11867 (N_11867,N_10244,N_10529);
xnor U11868 (N_11868,N_10936,N_11198);
nor U11869 (N_11869,N_10204,N_10946);
and U11870 (N_11870,N_10194,N_11085);
nand U11871 (N_11871,N_10870,N_10286);
or U11872 (N_11872,N_10699,N_11138);
nor U11873 (N_11873,N_10837,N_10183);
and U11874 (N_11874,N_10745,N_10724);
and U11875 (N_11875,N_10851,N_10646);
xor U11876 (N_11876,N_10455,N_10789);
nand U11877 (N_11877,N_11051,N_10114);
or U11878 (N_11878,N_10596,N_10529);
xnor U11879 (N_11879,N_10264,N_10947);
or U11880 (N_11880,N_10681,N_10353);
nor U11881 (N_11881,N_10971,N_10970);
nand U11882 (N_11882,N_10935,N_10185);
xor U11883 (N_11883,N_10016,N_10725);
xor U11884 (N_11884,N_10708,N_10132);
nor U11885 (N_11885,N_11086,N_11204);
xor U11886 (N_11886,N_10608,N_10429);
nand U11887 (N_11887,N_10413,N_10128);
xor U11888 (N_11888,N_10249,N_11073);
nor U11889 (N_11889,N_10618,N_10319);
nand U11890 (N_11890,N_10502,N_10137);
or U11891 (N_11891,N_10431,N_11055);
xor U11892 (N_11892,N_11228,N_10583);
xnor U11893 (N_11893,N_10940,N_10387);
nand U11894 (N_11894,N_10223,N_11161);
xnor U11895 (N_11895,N_10530,N_10659);
xor U11896 (N_11896,N_10370,N_10558);
nand U11897 (N_11897,N_10094,N_10939);
or U11898 (N_11898,N_10994,N_10321);
and U11899 (N_11899,N_10736,N_10883);
xnor U11900 (N_11900,N_10936,N_10601);
xnor U11901 (N_11901,N_11013,N_10126);
xnor U11902 (N_11902,N_10110,N_10776);
or U11903 (N_11903,N_10162,N_11029);
nand U11904 (N_11904,N_11094,N_11039);
xnor U11905 (N_11905,N_10793,N_10753);
or U11906 (N_11906,N_10445,N_11094);
and U11907 (N_11907,N_10820,N_10546);
or U11908 (N_11908,N_10062,N_11009);
nand U11909 (N_11909,N_10195,N_10842);
xor U11910 (N_11910,N_10835,N_10352);
xnor U11911 (N_11911,N_10848,N_10793);
nor U11912 (N_11912,N_10738,N_10733);
and U11913 (N_11913,N_10221,N_10130);
xnor U11914 (N_11914,N_11076,N_10808);
xnor U11915 (N_11915,N_10730,N_10318);
xor U11916 (N_11916,N_10475,N_11246);
or U11917 (N_11917,N_10573,N_10712);
and U11918 (N_11918,N_10841,N_10785);
or U11919 (N_11919,N_10586,N_11210);
nand U11920 (N_11920,N_10601,N_10820);
or U11921 (N_11921,N_11236,N_10670);
and U11922 (N_11922,N_10769,N_11032);
and U11923 (N_11923,N_11090,N_10038);
nor U11924 (N_11924,N_10316,N_10238);
or U11925 (N_11925,N_10544,N_10992);
nand U11926 (N_11926,N_10834,N_10459);
nand U11927 (N_11927,N_10358,N_10099);
nand U11928 (N_11928,N_10066,N_10731);
xnor U11929 (N_11929,N_10223,N_10267);
and U11930 (N_11930,N_11203,N_11097);
or U11931 (N_11931,N_11029,N_10015);
nor U11932 (N_11932,N_11188,N_11178);
xor U11933 (N_11933,N_10534,N_10407);
and U11934 (N_11934,N_10130,N_11031);
nand U11935 (N_11935,N_10276,N_10650);
xor U11936 (N_11936,N_10820,N_10413);
xor U11937 (N_11937,N_11132,N_10459);
or U11938 (N_11938,N_10842,N_10573);
or U11939 (N_11939,N_10263,N_10071);
nand U11940 (N_11940,N_10147,N_11007);
or U11941 (N_11941,N_10756,N_10067);
or U11942 (N_11942,N_10162,N_10933);
xnor U11943 (N_11943,N_10847,N_10407);
nor U11944 (N_11944,N_11201,N_10779);
and U11945 (N_11945,N_10120,N_10451);
nor U11946 (N_11946,N_10565,N_10105);
and U11947 (N_11947,N_10692,N_10017);
or U11948 (N_11948,N_10393,N_10201);
xnor U11949 (N_11949,N_11068,N_10501);
nand U11950 (N_11950,N_10247,N_10970);
xnor U11951 (N_11951,N_10516,N_10475);
and U11952 (N_11952,N_10225,N_10016);
nand U11953 (N_11953,N_11249,N_10785);
and U11954 (N_11954,N_10427,N_10259);
xor U11955 (N_11955,N_10169,N_10035);
or U11956 (N_11956,N_10982,N_10282);
nand U11957 (N_11957,N_10772,N_10229);
and U11958 (N_11958,N_10357,N_10363);
and U11959 (N_11959,N_10988,N_10554);
and U11960 (N_11960,N_11048,N_10163);
nand U11961 (N_11961,N_10629,N_10985);
or U11962 (N_11962,N_11139,N_10472);
and U11963 (N_11963,N_10124,N_10584);
nand U11964 (N_11964,N_10005,N_10591);
and U11965 (N_11965,N_10523,N_11001);
or U11966 (N_11966,N_10866,N_11049);
and U11967 (N_11967,N_10215,N_10347);
nand U11968 (N_11968,N_10398,N_10123);
nor U11969 (N_11969,N_10221,N_10669);
or U11970 (N_11970,N_10979,N_10517);
nor U11971 (N_11971,N_10110,N_11093);
and U11972 (N_11972,N_10928,N_11076);
xnor U11973 (N_11973,N_10816,N_10777);
nor U11974 (N_11974,N_10280,N_11114);
and U11975 (N_11975,N_11183,N_10256);
and U11976 (N_11976,N_10870,N_10744);
xor U11977 (N_11977,N_10438,N_11169);
and U11978 (N_11978,N_10520,N_11107);
xor U11979 (N_11979,N_10392,N_10354);
xnor U11980 (N_11980,N_10889,N_10292);
or U11981 (N_11981,N_10291,N_10200);
xnor U11982 (N_11982,N_10181,N_11062);
and U11983 (N_11983,N_11000,N_11033);
xor U11984 (N_11984,N_10593,N_10092);
and U11985 (N_11985,N_10209,N_10538);
and U11986 (N_11986,N_10418,N_10495);
and U11987 (N_11987,N_10204,N_10481);
and U11988 (N_11988,N_10182,N_10556);
and U11989 (N_11989,N_11120,N_11016);
or U11990 (N_11990,N_11024,N_10525);
and U11991 (N_11991,N_10792,N_10920);
xnor U11992 (N_11992,N_11185,N_10251);
nand U11993 (N_11993,N_10483,N_10145);
nor U11994 (N_11994,N_10876,N_10663);
xor U11995 (N_11995,N_10223,N_10055);
nor U11996 (N_11996,N_10715,N_10622);
xor U11997 (N_11997,N_10655,N_10501);
or U11998 (N_11998,N_10914,N_10898);
xnor U11999 (N_11999,N_10533,N_10651);
and U12000 (N_12000,N_10123,N_10786);
xor U12001 (N_12001,N_10116,N_11131);
or U12002 (N_12002,N_10417,N_10733);
and U12003 (N_12003,N_10179,N_10417);
or U12004 (N_12004,N_10574,N_10467);
nand U12005 (N_12005,N_10797,N_10146);
and U12006 (N_12006,N_11069,N_10149);
nor U12007 (N_12007,N_10220,N_10452);
nor U12008 (N_12008,N_10085,N_10977);
and U12009 (N_12009,N_10604,N_11119);
nor U12010 (N_12010,N_11192,N_10356);
nor U12011 (N_12011,N_11003,N_10978);
nor U12012 (N_12012,N_10278,N_10399);
xor U12013 (N_12013,N_10327,N_10390);
or U12014 (N_12014,N_10305,N_11171);
xor U12015 (N_12015,N_10141,N_11045);
nand U12016 (N_12016,N_10679,N_10970);
and U12017 (N_12017,N_11007,N_10963);
nor U12018 (N_12018,N_10441,N_10785);
xor U12019 (N_12019,N_10405,N_10323);
xor U12020 (N_12020,N_11150,N_10765);
or U12021 (N_12021,N_10497,N_10040);
and U12022 (N_12022,N_10532,N_10446);
xnor U12023 (N_12023,N_10789,N_10954);
xor U12024 (N_12024,N_10922,N_10130);
and U12025 (N_12025,N_10054,N_10999);
and U12026 (N_12026,N_11175,N_10900);
xnor U12027 (N_12027,N_10479,N_10936);
or U12028 (N_12028,N_10303,N_10973);
nor U12029 (N_12029,N_10572,N_10412);
nand U12030 (N_12030,N_10186,N_10266);
or U12031 (N_12031,N_10243,N_10773);
xor U12032 (N_12032,N_11052,N_10169);
or U12033 (N_12033,N_10115,N_10138);
nand U12034 (N_12034,N_10726,N_10156);
nand U12035 (N_12035,N_10516,N_10784);
nand U12036 (N_12036,N_11089,N_10209);
nor U12037 (N_12037,N_10574,N_10583);
xor U12038 (N_12038,N_10997,N_10543);
or U12039 (N_12039,N_10537,N_11231);
nor U12040 (N_12040,N_11193,N_10822);
and U12041 (N_12041,N_11141,N_11193);
nor U12042 (N_12042,N_10827,N_11243);
and U12043 (N_12043,N_10048,N_10464);
nor U12044 (N_12044,N_10664,N_11166);
xnor U12045 (N_12045,N_10866,N_11248);
or U12046 (N_12046,N_10925,N_11063);
or U12047 (N_12047,N_10731,N_10269);
nand U12048 (N_12048,N_10723,N_11203);
nand U12049 (N_12049,N_10927,N_10053);
or U12050 (N_12050,N_10270,N_10910);
or U12051 (N_12051,N_10233,N_10074);
nor U12052 (N_12052,N_10715,N_10204);
nor U12053 (N_12053,N_10043,N_10657);
xor U12054 (N_12054,N_10612,N_10547);
nand U12055 (N_12055,N_10863,N_10560);
nor U12056 (N_12056,N_10912,N_10328);
nand U12057 (N_12057,N_10182,N_10818);
and U12058 (N_12058,N_11007,N_10266);
or U12059 (N_12059,N_10340,N_10630);
and U12060 (N_12060,N_10807,N_10562);
xnor U12061 (N_12061,N_11246,N_10034);
xnor U12062 (N_12062,N_10230,N_10038);
nor U12063 (N_12063,N_10770,N_10565);
and U12064 (N_12064,N_10582,N_10791);
or U12065 (N_12065,N_10818,N_11201);
xnor U12066 (N_12066,N_10831,N_10555);
nor U12067 (N_12067,N_11093,N_10387);
and U12068 (N_12068,N_10185,N_10537);
nand U12069 (N_12069,N_10394,N_10576);
nor U12070 (N_12070,N_10979,N_11043);
and U12071 (N_12071,N_10539,N_11208);
or U12072 (N_12072,N_11178,N_10387);
xor U12073 (N_12073,N_10019,N_10666);
and U12074 (N_12074,N_11110,N_11036);
or U12075 (N_12075,N_10776,N_10903);
or U12076 (N_12076,N_10257,N_10342);
nor U12077 (N_12077,N_10424,N_10363);
nand U12078 (N_12078,N_10557,N_11007);
xnor U12079 (N_12079,N_10176,N_10457);
nor U12080 (N_12080,N_10114,N_10678);
and U12081 (N_12081,N_10765,N_10615);
nor U12082 (N_12082,N_10186,N_10327);
nor U12083 (N_12083,N_10528,N_10332);
or U12084 (N_12084,N_10429,N_10029);
nor U12085 (N_12085,N_11232,N_11100);
nor U12086 (N_12086,N_10859,N_11153);
or U12087 (N_12087,N_10533,N_10963);
xnor U12088 (N_12088,N_10577,N_10556);
nor U12089 (N_12089,N_10454,N_10853);
xnor U12090 (N_12090,N_10103,N_10310);
and U12091 (N_12091,N_10141,N_10056);
nor U12092 (N_12092,N_11207,N_10417);
and U12093 (N_12093,N_10496,N_10117);
and U12094 (N_12094,N_10341,N_10266);
and U12095 (N_12095,N_10610,N_11183);
nand U12096 (N_12096,N_11231,N_10669);
and U12097 (N_12097,N_10755,N_10321);
and U12098 (N_12098,N_10673,N_10418);
xnor U12099 (N_12099,N_11214,N_10804);
or U12100 (N_12100,N_10801,N_10574);
xor U12101 (N_12101,N_11243,N_11210);
nor U12102 (N_12102,N_11100,N_10652);
nand U12103 (N_12103,N_11110,N_10813);
or U12104 (N_12104,N_10974,N_10852);
nand U12105 (N_12105,N_10703,N_11036);
or U12106 (N_12106,N_10598,N_10044);
nand U12107 (N_12107,N_10616,N_11016);
and U12108 (N_12108,N_10447,N_10460);
nand U12109 (N_12109,N_10287,N_10825);
and U12110 (N_12110,N_10703,N_10259);
and U12111 (N_12111,N_11118,N_10977);
or U12112 (N_12112,N_10765,N_10292);
or U12113 (N_12113,N_10171,N_10205);
and U12114 (N_12114,N_10503,N_10835);
nor U12115 (N_12115,N_11139,N_10370);
nand U12116 (N_12116,N_11100,N_10973);
xnor U12117 (N_12117,N_10664,N_10038);
and U12118 (N_12118,N_10774,N_10183);
xor U12119 (N_12119,N_10669,N_10521);
nand U12120 (N_12120,N_11095,N_10587);
and U12121 (N_12121,N_10371,N_11068);
and U12122 (N_12122,N_10682,N_10524);
or U12123 (N_12123,N_10037,N_10514);
nor U12124 (N_12124,N_10492,N_10975);
nor U12125 (N_12125,N_10473,N_10355);
xor U12126 (N_12126,N_11030,N_10023);
and U12127 (N_12127,N_10014,N_10298);
xor U12128 (N_12128,N_10446,N_11048);
nor U12129 (N_12129,N_10604,N_10114);
and U12130 (N_12130,N_10829,N_10394);
nand U12131 (N_12131,N_10784,N_10633);
xnor U12132 (N_12132,N_10061,N_10094);
and U12133 (N_12133,N_10261,N_10819);
or U12134 (N_12134,N_10311,N_10635);
nand U12135 (N_12135,N_10952,N_10303);
and U12136 (N_12136,N_10523,N_10689);
and U12137 (N_12137,N_10461,N_10049);
and U12138 (N_12138,N_10119,N_11240);
xor U12139 (N_12139,N_10741,N_10878);
xor U12140 (N_12140,N_10023,N_10696);
nor U12141 (N_12141,N_11100,N_10387);
nor U12142 (N_12142,N_10050,N_10915);
nand U12143 (N_12143,N_10478,N_10528);
nor U12144 (N_12144,N_11148,N_10020);
nand U12145 (N_12145,N_10910,N_10367);
and U12146 (N_12146,N_10515,N_10116);
nand U12147 (N_12147,N_10342,N_10694);
xnor U12148 (N_12148,N_11171,N_10556);
or U12149 (N_12149,N_10716,N_10149);
and U12150 (N_12150,N_10113,N_10216);
and U12151 (N_12151,N_10430,N_10875);
xor U12152 (N_12152,N_10218,N_10607);
xor U12153 (N_12153,N_10852,N_10217);
nand U12154 (N_12154,N_11217,N_10376);
nor U12155 (N_12155,N_10686,N_10581);
nand U12156 (N_12156,N_10256,N_10358);
xor U12157 (N_12157,N_10510,N_10683);
xnor U12158 (N_12158,N_11103,N_10386);
nand U12159 (N_12159,N_10275,N_10191);
xor U12160 (N_12160,N_10140,N_10760);
nand U12161 (N_12161,N_11063,N_11009);
nor U12162 (N_12162,N_11055,N_10817);
nand U12163 (N_12163,N_10742,N_10627);
and U12164 (N_12164,N_10306,N_10529);
or U12165 (N_12165,N_11096,N_10961);
and U12166 (N_12166,N_10188,N_10161);
xnor U12167 (N_12167,N_10110,N_10067);
and U12168 (N_12168,N_10923,N_10185);
xor U12169 (N_12169,N_11150,N_11146);
nor U12170 (N_12170,N_10604,N_10680);
nand U12171 (N_12171,N_11160,N_11236);
nand U12172 (N_12172,N_11183,N_10553);
xnor U12173 (N_12173,N_10799,N_11041);
xnor U12174 (N_12174,N_10829,N_10561);
or U12175 (N_12175,N_10922,N_11068);
and U12176 (N_12176,N_10637,N_10292);
and U12177 (N_12177,N_10687,N_10217);
nor U12178 (N_12178,N_10214,N_10945);
xnor U12179 (N_12179,N_10912,N_10916);
xnor U12180 (N_12180,N_11089,N_10020);
nor U12181 (N_12181,N_10218,N_10676);
or U12182 (N_12182,N_10314,N_10026);
nor U12183 (N_12183,N_10887,N_11244);
nand U12184 (N_12184,N_10450,N_10643);
and U12185 (N_12185,N_11161,N_10641);
and U12186 (N_12186,N_10425,N_10027);
nor U12187 (N_12187,N_10253,N_10648);
xor U12188 (N_12188,N_10383,N_11040);
xnor U12189 (N_12189,N_10609,N_10912);
nand U12190 (N_12190,N_10299,N_10942);
nand U12191 (N_12191,N_10023,N_10857);
xnor U12192 (N_12192,N_10001,N_11142);
nor U12193 (N_12193,N_10447,N_10200);
xor U12194 (N_12194,N_10166,N_10104);
nand U12195 (N_12195,N_10544,N_11249);
or U12196 (N_12196,N_10541,N_11206);
xnor U12197 (N_12197,N_10087,N_11137);
xnor U12198 (N_12198,N_10137,N_10556);
nor U12199 (N_12199,N_10583,N_10416);
nand U12200 (N_12200,N_11155,N_10748);
or U12201 (N_12201,N_10358,N_10540);
xnor U12202 (N_12202,N_10504,N_10738);
nand U12203 (N_12203,N_10933,N_10034);
and U12204 (N_12204,N_10981,N_11048);
or U12205 (N_12205,N_10753,N_11243);
or U12206 (N_12206,N_10180,N_10269);
nor U12207 (N_12207,N_11090,N_10425);
xor U12208 (N_12208,N_10401,N_10600);
nand U12209 (N_12209,N_10237,N_10903);
and U12210 (N_12210,N_11244,N_10004);
xnor U12211 (N_12211,N_10997,N_11185);
and U12212 (N_12212,N_10290,N_11172);
and U12213 (N_12213,N_10661,N_11211);
xor U12214 (N_12214,N_10361,N_10399);
and U12215 (N_12215,N_10566,N_11049);
xor U12216 (N_12216,N_10931,N_10605);
or U12217 (N_12217,N_11086,N_10890);
nor U12218 (N_12218,N_10974,N_10584);
or U12219 (N_12219,N_10123,N_10883);
or U12220 (N_12220,N_10925,N_10578);
and U12221 (N_12221,N_10882,N_10331);
nor U12222 (N_12222,N_10147,N_10904);
nor U12223 (N_12223,N_11163,N_10258);
and U12224 (N_12224,N_10614,N_10462);
nor U12225 (N_12225,N_10745,N_10091);
or U12226 (N_12226,N_10088,N_10349);
xor U12227 (N_12227,N_11147,N_11058);
and U12228 (N_12228,N_11222,N_10251);
nand U12229 (N_12229,N_10508,N_11198);
nor U12230 (N_12230,N_10435,N_11136);
xnor U12231 (N_12231,N_10071,N_11130);
nor U12232 (N_12232,N_10907,N_10207);
nor U12233 (N_12233,N_10412,N_10207);
nand U12234 (N_12234,N_10815,N_10679);
xor U12235 (N_12235,N_11103,N_11241);
nand U12236 (N_12236,N_10654,N_10922);
nor U12237 (N_12237,N_10938,N_11110);
nand U12238 (N_12238,N_10101,N_10171);
nand U12239 (N_12239,N_10477,N_10551);
nor U12240 (N_12240,N_10224,N_10372);
nor U12241 (N_12241,N_11043,N_10160);
or U12242 (N_12242,N_10719,N_11038);
nor U12243 (N_12243,N_10651,N_10256);
or U12244 (N_12244,N_10988,N_10953);
nor U12245 (N_12245,N_10013,N_11000);
xor U12246 (N_12246,N_10083,N_10640);
or U12247 (N_12247,N_11233,N_10226);
nand U12248 (N_12248,N_11112,N_10209);
and U12249 (N_12249,N_10761,N_10769);
and U12250 (N_12250,N_10552,N_10695);
xor U12251 (N_12251,N_11202,N_10595);
nand U12252 (N_12252,N_10671,N_10205);
or U12253 (N_12253,N_10654,N_10297);
nor U12254 (N_12254,N_10839,N_10678);
nand U12255 (N_12255,N_10555,N_10265);
and U12256 (N_12256,N_10884,N_10631);
or U12257 (N_12257,N_10549,N_10992);
or U12258 (N_12258,N_11103,N_10118);
xor U12259 (N_12259,N_10726,N_10231);
nand U12260 (N_12260,N_10264,N_10701);
and U12261 (N_12261,N_10416,N_10872);
nor U12262 (N_12262,N_10050,N_10192);
or U12263 (N_12263,N_10853,N_10932);
xor U12264 (N_12264,N_11183,N_10134);
nor U12265 (N_12265,N_10164,N_10996);
or U12266 (N_12266,N_10138,N_10068);
nor U12267 (N_12267,N_10244,N_10525);
nand U12268 (N_12268,N_10226,N_10517);
or U12269 (N_12269,N_10266,N_11150);
nand U12270 (N_12270,N_10184,N_10779);
nor U12271 (N_12271,N_10832,N_10814);
and U12272 (N_12272,N_10668,N_10253);
or U12273 (N_12273,N_11226,N_10830);
xor U12274 (N_12274,N_10882,N_10714);
or U12275 (N_12275,N_10951,N_11125);
xor U12276 (N_12276,N_10496,N_10869);
nand U12277 (N_12277,N_10849,N_10634);
or U12278 (N_12278,N_10863,N_10377);
nor U12279 (N_12279,N_10248,N_11062);
nor U12280 (N_12280,N_10215,N_10500);
xor U12281 (N_12281,N_10619,N_10758);
and U12282 (N_12282,N_10629,N_10110);
nand U12283 (N_12283,N_10455,N_10171);
nor U12284 (N_12284,N_10846,N_10558);
nand U12285 (N_12285,N_10511,N_10030);
nand U12286 (N_12286,N_10546,N_10405);
nand U12287 (N_12287,N_10791,N_10620);
nand U12288 (N_12288,N_11049,N_10225);
nand U12289 (N_12289,N_11017,N_11079);
and U12290 (N_12290,N_10988,N_10324);
and U12291 (N_12291,N_10443,N_10561);
xor U12292 (N_12292,N_10010,N_10472);
nand U12293 (N_12293,N_11088,N_10622);
and U12294 (N_12294,N_10293,N_11208);
nand U12295 (N_12295,N_10689,N_10723);
nand U12296 (N_12296,N_10179,N_10864);
nand U12297 (N_12297,N_11054,N_10925);
or U12298 (N_12298,N_10755,N_10295);
xnor U12299 (N_12299,N_10076,N_10315);
nor U12300 (N_12300,N_10495,N_10206);
and U12301 (N_12301,N_10612,N_10646);
or U12302 (N_12302,N_11081,N_10353);
or U12303 (N_12303,N_10112,N_10888);
nand U12304 (N_12304,N_10117,N_10293);
nor U12305 (N_12305,N_10589,N_10559);
nor U12306 (N_12306,N_10077,N_10239);
xnor U12307 (N_12307,N_10789,N_10897);
nor U12308 (N_12308,N_10785,N_10769);
nor U12309 (N_12309,N_10757,N_10845);
nand U12310 (N_12310,N_10794,N_10945);
and U12311 (N_12311,N_10951,N_10892);
nand U12312 (N_12312,N_10875,N_10649);
and U12313 (N_12313,N_11082,N_10955);
or U12314 (N_12314,N_10027,N_10498);
nor U12315 (N_12315,N_10962,N_10100);
xnor U12316 (N_12316,N_10097,N_11101);
nand U12317 (N_12317,N_10298,N_10282);
xor U12318 (N_12318,N_10235,N_11134);
or U12319 (N_12319,N_10001,N_10390);
or U12320 (N_12320,N_11032,N_11229);
or U12321 (N_12321,N_10242,N_10259);
and U12322 (N_12322,N_10842,N_10211);
nand U12323 (N_12323,N_10239,N_10296);
xor U12324 (N_12324,N_10772,N_10456);
nand U12325 (N_12325,N_10495,N_10393);
xnor U12326 (N_12326,N_10577,N_11043);
nor U12327 (N_12327,N_10837,N_10121);
nand U12328 (N_12328,N_11094,N_11050);
nand U12329 (N_12329,N_10018,N_10042);
nand U12330 (N_12330,N_10922,N_10053);
or U12331 (N_12331,N_11188,N_10364);
nor U12332 (N_12332,N_10847,N_11007);
xnor U12333 (N_12333,N_11071,N_10783);
or U12334 (N_12334,N_10224,N_10820);
nand U12335 (N_12335,N_10282,N_10621);
nor U12336 (N_12336,N_11010,N_10358);
xor U12337 (N_12337,N_10858,N_10812);
nand U12338 (N_12338,N_11181,N_11090);
nand U12339 (N_12339,N_10828,N_11025);
xor U12340 (N_12340,N_10861,N_10661);
xnor U12341 (N_12341,N_10015,N_11143);
xor U12342 (N_12342,N_11027,N_11074);
xor U12343 (N_12343,N_10165,N_10637);
and U12344 (N_12344,N_10690,N_10817);
nand U12345 (N_12345,N_10803,N_10851);
xnor U12346 (N_12346,N_10214,N_11056);
xnor U12347 (N_12347,N_10257,N_10007);
nor U12348 (N_12348,N_10223,N_10413);
nand U12349 (N_12349,N_10653,N_11185);
or U12350 (N_12350,N_10184,N_10918);
xnor U12351 (N_12351,N_10762,N_10760);
nand U12352 (N_12352,N_11187,N_10985);
nor U12353 (N_12353,N_10981,N_10685);
or U12354 (N_12354,N_11157,N_10312);
nor U12355 (N_12355,N_10845,N_10402);
nor U12356 (N_12356,N_10474,N_11210);
nor U12357 (N_12357,N_10106,N_10926);
or U12358 (N_12358,N_11024,N_10255);
nor U12359 (N_12359,N_11087,N_10260);
nand U12360 (N_12360,N_10506,N_10617);
nor U12361 (N_12361,N_10915,N_10805);
nor U12362 (N_12362,N_10193,N_10568);
and U12363 (N_12363,N_10899,N_10949);
nor U12364 (N_12364,N_10736,N_10281);
nand U12365 (N_12365,N_10280,N_10023);
nor U12366 (N_12366,N_10854,N_11163);
xnor U12367 (N_12367,N_10756,N_10491);
xor U12368 (N_12368,N_10749,N_10084);
and U12369 (N_12369,N_11122,N_10565);
or U12370 (N_12370,N_10821,N_10541);
xnor U12371 (N_12371,N_10450,N_10932);
and U12372 (N_12372,N_10811,N_11109);
nor U12373 (N_12373,N_10736,N_10630);
and U12374 (N_12374,N_10291,N_10138);
and U12375 (N_12375,N_11045,N_11035);
nor U12376 (N_12376,N_10861,N_11181);
nor U12377 (N_12377,N_10376,N_10969);
or U12378 (N_12378,N_11199,N_11213);
xnor U12379 (N_12379,N_10628,N_10148);
or U12380 (N_12380,N_10233,N_10801);
or U12381 (N_12381,N_11170,N_10694);
nor U12382 (N_12382,N_11164,N_10097);
nor U12383 (N_12383,N_11101,N_10303);
xnor U12384 (N_12384,N_10325,N_11184);
and U12385 (N_12385,N_11127,N_10674);
nor U12386 (N_12386,N_10337,N_10193);
and U12387 (N_12387,N_10322,N_10390);
nor U12388 (N_12388,N_11057,N_10366);
nor U12389 (N_12389,N_10474,N_11103);
nand U12390 (N_12390,N_10788,N_10229);
or U12391 (N_12391,N_10699,N_11191);
xor U12392 (N_12392,N_10897,N_10250);
nand U12393 (N_12393,N_10133,N_10033);
and U12394 (N_12394,N_10609,N_10844);
or U12395 (N_12395,N_10666,N_10313);
nand U12396 (N_12396,N_11112,N_10335);
nor U12397 (N_12397,N_11029,N_10764);
and U12398 (N_12398,N_11249,N_10235);
nand U12399 (N_12399,N_10399,N_11061);
nand U12400 (N_12400,N_11049,N_10368);
nand U12401 (N_12401,N_10288,N_10984);
nor U12402 (N_12402,N_11187,N_10686);
or U12403 (N_12403,N_10107,N_10641);
or U12404 (N_12404,N_11036,N_10980);
or U12405 (N_12405,N_10281,N_10221);
or U12406 (N_12406,N_11137,N_10939);
or U12407 (N_12407,N_10872,N_10550);
nor U12408 (N_12408,N_11209,N_11060);
nor U12409 (N_12409,N_10592,N_10306);
xnor U12410 (N_12410,N_10921,N_10656);
nand U12411 (N_12411,N_10098,N_10969);
and U12412 (N_12412,N_10549,N_10763);
xor U12413 (N_12413,N_10133,N_10167);
or U12414 (N_12414,N_10667,N_10906);
nor U12415 (N_12415,N_10238,N_10888);
nor U12416 (N_12416,N_10745,N_10973);
or U12417 (N_12417,N_10203,N_10949);
and U12418 (N_12418,N_10313,N_10578);
or U12419 (N_12419,N_10849,N_10772);
nor U12420 (N_12420,N_10014,N_10986);
xor U12421 (N_12421,N_10303,N_10435);
nor U12422 (N_12422,N_10240,N_10298);
nand U12423 (N_12423,N_10384,N_10514);
xnor U12424 (N_12424,N_11018,N_10994);
xor U12425 (N_12425,N_11135,N_10660);
or U12426 (N_12426,N_10638,N_10241);
or U12427 (N_12427,N_11178,N_10720);
and U12428 (N_12428,N_10740,N_10209);
and U12429 (N_12429,N_10644,N_10656);
and U12430 (N_12430,N_10273,N_10298);
xor U12431 (N_12431,N_10611,N_10155);
or U12432 (N_12432,N_10651,N_10207);
xnor U12433 (N_12433,N_10022,N_11016);
nor U12434 (N_12434,N_10484,N_10595);
nand U12435 (N_12435,N_10273,N_10486);
and U12436 (N_12436,N_10157,N_10331);
or U12437 (N_12437,N_11176,N_10479);
or U12438 (N_12438,N_11131,N_10541);
and U12439 (N_12439,N_10320,N_10282);
and U12440 (N_12440,N_10099,N_10874);
xor U12441 (N_12441,N_10579,N_10732);
nor U12442 (N_12442,N_10967,N_10308);
nor U12443 (N_12443,N_10077,N_10812);
or U12444 (N_12444,N_10282,N_11205);
nand U12445 (N_12445,N_10391,N_11007);
nor U12446 (N_12446,N_11019,N_11104);
nand U12447 (N_12447,N_11146,N_10474);
and U12448 (N_12448,N_10733,N_10266);
or U12449 (N_12449,N_11021,N_10803);
or U12450 (N_12450,N_10014,N_10820);
xnor U12451 (N_12451,N_10430,N_10447);
nor U12452 (N_12452,N_10729,N_10769);
nor U12453 (N_12453,N_10880,N_10976);
xor U12454 (N_12454,N_10651,N_10045);
xnor U12455 (N_12455,N_11059,N_10363);
xnor U12456 (N_12456,N_10454,N_11053);
or U12457 (N_12457,N_11131,N_10471);
nand U12458 (N_12458,N_10746,N_11096);
nand U12459 (N_12459,N_10779,N_10384);
or U12460 (N_12460,N_10246,N_10406);
nor U12461 (N_12461,N_10834,N_10021);
nor U12462 (N_12462,N_10161,N_10865);
nand U12463 (N_12463,N_10408,N_10602);
or U12464 (N_12464,N_10902,N_11231);
or U12465 (N_12465,N_10273,N_10636);
xnor U12466 (N_12466,N_10295,N_10118);
or U12467 (N_12467,N_10092,N_10381);
xnor U12468 (N_12468,N_10575,N_10846);
and U12469 (N_12469,N_10234,N_10161);
and U12470 (N_12470,N_10816,N_10262);
and U12471 (N_12471,N_10648,N_10714);
nand U12472 (N_12472,N_10133,N_11115);
xor U12473 (N_12473,N_10016,N_10939);
and U12474 (N_12474,N_10920,N_10070);
or U12475 (N_12475,N_10304,N_10419);
xor U12476 (N_12476,N_10779,N_10359);
xor U12477 (N_12477,N_10189,N_10665);
and U12478 (N_12478,N_10495,N_10198);
xnor U12479 (N_12479,N_10082,N_10135);
and U12480 (N_12480,N_10688,N_10230);
or U12481 (N_12481,N_10894,N_10587);
nand U12482 (N_12482,N_10554,N_10671);
or U12483 (N_12483,N_11146,N_11173);
nand U12484 (N_12484,N_11215,N_11105);
nor U12485 (N_12485,N_11230,N_10811);
nor U12486 (N_12486,N_10679,N_10972);
or U12487 (N_12487,N_10922,N_10854);
xor U12488 (N_12488,N_10295,N_10285);
xor U12489 (N_12489,N_10763,N_10806);
nor U12490 (N_12490,N_10685,N_10662);
or U12491 (N_12491,N_10346,N_10309);
nand U12492 (N_12492,N_10299,N_10663);
nor U12493 (N_12493,N_10528,N_10997);
nand U12494 (N_12494,N_10308,N_10896);
nand U12495 (N_12495,N_10250,N_11226);
and U12496 (N_12496,N_10169,N_11240);
nand U12497 (N_12497,N_10827,N_11042);
nor U12498 (N_12498,N_10927,N_10471);
or U12499 (N_12499,N_10420,N_10493);
nand U12500 (N_12500,N_11969,N_11493);
xor U12501 (N_12501,N_12196,N_11714);
or U12502 (N_12502,N_11368,N_12369);
or U12503 (N_12503,N_12136,N_11763);
nand U12504 (N_12504,N_11473,N_12471);
and U12505 (N_12505,N_11488,N_11390);
nor U12506 (N_12506,N_12025,N_12068);
xnor U12507 (N_12507,N_12328,N_12029);
nor U12508 (N_12508,N_11287,N_11960);
or U12509 (N_12509,N_12122,N_11898);
and U12510 (N_12510,N_11722,N_12318);
xor U12511 (N_12511,N_12284,N_11756);
xnor U12512 (N_12512,N_11550,N_11948);
xnor U12513 (N_12513,N_11329,N_12483);
xor U12514 (N_12514,N_11583,N_12329);
xnor U12515 (N_12515,N_12453,N_11262);
and U12516 (N_12516,N_12071,N_11569);
nor U12517 (N_12517,N_12141,N_11646);
nor U12518 (N_12518,N_12049,N_11676);
and U12519 (N_12519,N_11618,N_11444);
xnor U12520 (N_12520,N_11528,N_11386);
or U12521 (N_12521,N_11438,N_11917);
nand U12522 (N_12522,N_11650,N_12433);
and U12523 (N_12523,N_11812,N_12211);
and U12524 (N_12524,N_11467,N_12004);
or U12525 (N_12525,N_12451,N_12175);
nand U12526 (N_12526,N_11779,N_12380);
xor U12527 (N_12527,N_11310,N_12394);
nand U12528 (N_12528,N_11652,N_11522);
nand U12529 (N_12529,N_12073,N_11540);
xnor U12530 (N_12530,N_11864,N_11346);
nand U12531 (N_12531,N_11733,N_11869);
nor U12532 (N_12532,N_12174,N_11786);
and U12533 (N_12533,N_12045,N_11562);
or U12534 (N_12534,N_11956,N_11985);
or U12535 (N_12535,N_12359,N_11399);
nand U12536 (N_12536,N_11952,N_11635);
nor U12537 (N_12537,N_12110,N_12276);
nor U12538 (N_12538,N_11315,N_11318);
nand U12539 (N_12539,N_12269,N_12186);
xor U12540 (N_12540,N_12367,N_12240);
or U12541 (N_12541,N_11633,N_12140);
or U12542 (N_12542,N_11566,N_12476);
xor U12543 (N_12543,N_12147,N_11776);
and U12544 (N_12544,N_11749,N_11766);
and U12545 (N_12545,N_11311,N_11589);
nand U12546 (N_12546,N_12443,N_12387);
nor U12547 (N_12547,N_11447,N_11451);
nand U12548 (N_12548,N_11526,N_11545);
nand U12549 (N_12549,N_11920,N_11790);
nand U12550 (N_12550,N_12111,N_12492);
xnor U12551 (N_12551,N_12388,N_12270);
nor U12552 (N_12552,N_12094,N_11362);
or U12553 (N_12553,N_12378,N_11515);
nand U12554 (N_12554,N_12324,N_12044);
and U12555 (N_12555,N_11289,N_11813);
or U12556 (N_12556,N_12330,N_11699);
xnor U12557 (N_12557,N_11608,N_11865);
xor U12558 (N_12558,N_11416,N_12121);
xnor U12559 (N_12559,N_11638,N_11874);
and U12560 (N_12560,N_12470,N_12295);
nor U12561 (N_12561,N_11902,N_12233);
or U12562 (N_12562,N_11290,N_12048);
nand U12563 (N_12563,N_11335,N_12265);
and U12564 (N_12564,N_11365,N_11951);
nand U12565 (N_12565,N_12146,N_11272);
nand U12566 (N_12566,N_12345,N_12159);
xnor U12567 (N_12567,N_11372,N_11876);
nor U12568 (N_12568,N_12181,N_11989);
and U12569 (N_12569,N_12493,N_12484);
xnor U12570 (N_12570,N_11990,N_11421);
xor U12571 (N_12571,N_11619,N_11701);
or U12572 (N_12572,N_12206,N_11840);
and U12573 (N_12573,N_11600,N_11556);
nor U12574 (N_12574,N_11634,N_11928);
or U12575 (N_12575,N_11643,N_12237);
and U12576 (N_12576,N_12158,N_11552);
nor U12577 (N_12577,N_11387,N_11542);
and U12578 (N_12578,N_11516,N_11453);
xnor U12579 (N_12579,N_11975,N_12148);
and U12580 (N_12580,N_11624,N_11342);
xnor U12581 (N_12581,N_12098,N_12489);
or U12582 (N_12582,N_12225,N_11477);
nand U12583 (N_12583,N_11724,N_12127);
or U12584 (N_12584,N_12400,N_11403);
xnor U12585 (N_12585,N_11737,N_11498);
nand U12586 (N_12586,N_12007,N_11674);
nand U12587 (N_12587,N_11564,N_12368);
nand U12588 (N_12588,N_12301,N_12249);
nor U12589 (N_12589,N_12477,N_11879);
xnor U12590 (N_12590,N_12473,N_11767);
or U12591 (N_12591,N_12198,N_12143);
and U12592 (N_12592,N_12227,N_11464);
nand U12593 (N_12593,N_12074,N_11509);
nand U12594 (N_12594,N_11506,N_11578);
nand U12595 (N_12595,N_12303,N_11844);
or U12596 (N_12596,N_11980,N_11715);
and U12597 (N_12597,N_12251,N_11941);
nor U12598 (N_12598,N_12238,N_11487);
nor U12599 (N_12599,N_12307,N_11405);
nor U12600 (N_12600,N_12219,N_11751);
or U12601 (N_12601,N_11910,N_11470);
and U12602 (N_12602,N_12188,N_11883);
or U12603 (N_12603,N_12364,N_12397);
and U12604 (N_12604,N_12455,N_11866);
nor U12605 (N_12605,N_12106,N_11423);
nand U12606 (N_12606,N_12480,N_12138);
nand U12607 (N_12607,N_12457,N_11859);
xnor U12608 (N_12608,N_11503,N_12180);
or U12609 (N_12609,N_11300,N_11384);
and U12610 (N_12610,N_11553,N_12218);
nand U12611 (N_12611,N_12228,N_11870);
nor U12612 (N_12612,N_12360,N_11445);
xnor U12613 (N_12613,N_11663,N_12323);
nand U12614 (N_12614,N_11871,N_11338);
and U12615 (N_12615,N_11430,N_11449);
and U12616 (N_12616,N_12195,N_12282);
xor U12617 (N_12617,N_12467,N_11424);
or U12618 (N_12618,N_11986,N_11432);
or U12619 (N_12619,N_12461,N_11884);
xnor U12620 (N_12620,N_12463,N_12450);
and U12621 (N_12621,N_12145,N_12267);
xnor U12622 (N_12622,N_12039,N_11582);
and U12623 (N_12623,N_11484,N_11662);
or U12624 (N_12624,N_11773,N_11687);
or U12625 (N_12625,N_12032,N_11966);
and U12626 (N_12626,N_11426,N_11429);
nand U12627 (N_12627,N_12379,N_12280);
and U12628 (N_12628,N_11856,N_11350);
or U12629 (N_12629,N_11734,N_11595);
nand U12630 (N_12630,N_11826,N_12221);
nand U12631 (N_12631,N_12056,N_12396);
nor U12632 (N_12632,N_12348,N_11567);
xor U12633 (N_12633,N_12452,N_11532);
xnor U12634 (N_12634,N_11323,N_11795);
and U12635 (N_12635,N_12449,N_11913);
and U12636 (N_12636,N_11725,N_11260);
or U12637 (N_12637,N_11909,N_11292);
and U12638 (N_12638,N_11997,N_11847);
and U12639 (N_12639,N_11769,N_11958);
nand U12640 (N_12640,N_11831,N_12352);
or U12641 (N_12641,N_12028,N_11721);
or U12642 (N_12642,N_11620,N_11630);
and U12643 (N_12643,N_11857,N_11736);
and U12644 (N_12644,N_11609,N_11692);
and U12645 (N_12645,N_12254,N_11875);
or U12646 (N_12646,N_12070,N_12320);
nand U12647 (N_12647,N_11584,N_11546);
nand U12648 (N_12648,N_12339,N_11801);
or U12649 (N_12649,N_12478,N_11726);
xnor U12650 (N_12650,N_12179,N_11732);
xor U12651 (N_12651,N_11750,N_12137);
nand U12652 (N_12652,N_12021,N_11418);
or U12653 (N_12653,N_12084,N_11984);
nor U12654 (N_12654,N_11436,N_12172);
nand U12655 (N_12655,N_12445,N_12187);
and U12656 (N_12656,N_12031,N_11837);
nor U12657 (N_12657,N_11848,N_11929);
and U12658 (N_12658,N_11500,N_12075);
and U12659 (N_12659,N_11998,N_11382);
xnor U12660 (N_12660,N_12101,N_11427);
nand U12661 (N_12661,N_11574,N_11458);
or U12662 (N_12662,N_11658,N_11435);
nor U12663 (N_12663,N_11393,N_11881);
xor U12664 (N_12664,N_11781,N_11838);
nor U12665 (N_12665,N_11480,N_12335);
and U12666 (N_12666,N_12439,N_12042);
or U12667 (N_12667,N_11330,N_11842);
xor U12668 (N_12668,N_11557,N_12223);
or U12669 (N_12669,N_12413,N_11759);
and U12670 (N_12670,N_12234,N_12142);
and U12671 (N_12671,N_11852,N_11700);
and U12672 (N_12672,N_11681,N_11568);
and U12673 (N_12673,N_11683,N_11544);
xnor U12674 (N_12674,N_11784,N_12003);
xor U12675 (N_12675,N_11299,N_12432);
and U12676 (N_12676,N_11959,N_11413);
nor U12677 (N_12677,N_12277,N_11370);
nor U12678 (N_12678,N_12023,N_12459);
xor U12679 (N_12679,N_11369,N_11392);
nand U12680 (N_12680,N_12382,N_11268);
xor U12681 (N_12681,N_11706,N_11450);
nand U12682 (N_12682,N_11926,N_12057);
and U12683 (N_12683,N_11601,N_12222);
or U12684 (N_12684,N_11476,N_11351);
and U12685 (N_12685,N_12216,N_12311);
or U12686 (N_12686,N_12060,N_11353);
and U12687 (N_12687,N_11697,N_11925);
xor U12688 (N_12688,N_12469,N_11291);
or U12689 (N_12689,N_11944,N_12168);
and U12690 (N_12690,N_12430,N_11481);
and U12691 (N_12691,N_11478,N_12244);
or U12692 (N_12692,N_11520,N_12210);
nor U12693 (N_12693,N_12185,N_11823);
and U12694 (N_12694,N_11381,N_12093);
nand U12695 (N_12695,N_11366,N_11294);
or U12696 (N_12696,N_11474,N_12481);
xor U12697 (N_12697,N_11905,N_12299);
nand U12698 (N_12698,N_12114,N_12474);
nand U12699 (N_12699,N_11337,N_11862);
and U12700 (N_12700,N_11694,N_11617);
xnor U12701 (N_12701,N_11901,N_12064);
and U12702 (N_12702,N_11753,N_12434);
nand U12703 (N_12703,N_11996,N_12108);
nand U12704 (N_12704,N_12373,N_11462);
xnor U12705 (N_12705,N_11672,N_11973);
and U12706 (N_12706,N_11252,N_12333);
nor U12707 (N_12707,N_11334,N_11810);
nand U12708 (N_12708,N_11938,N_11296);
and U12709 (N_12709,N_12343,N_11271);
xor U12710 (N_12710,N_12479,N_11570);
nand U12711 (N_12711,N_11954,N_12340);
nor U12712 (N_12712,N_12212,N_11629);
and U12713 (N_12713,N_12207,N_11460);
nor U12714 (N_12714,N_11541,N_12266);
and U12715 (N_12715,N_11911,N_11757);
or U12716 (N_12716,N_12043,N_12016);
and U12717 (N_12717,N_11796,N_12118);
nor U12718 (N_12718,N_11730,N_11896);
or U12719 (N_12719,N_12447,N_11855);
xor U12720 (N_12720,N_11765,N_12006);
and U12721 (N_12721,N_11961,N_11906);
and U12722 (N_12722,N_12128,N_11853);
xor U12723 (N_12723,N_11915,N_11306);
or U12724 (N_12724,N_11356,N_12072);
nor U12725 (N_12725,N_11828,N_12317);
and U12726 (N_12726,N_12164,N_11454);
xor U12727 (N_12727,N_11554,N_12253);
xor U12728 (N_12728,N_12058,N_11811);
xnor U12729 (N_12729,N_11265,N_11317);
or U12730 (N_12730,N_12066,N_12202);
nand U12731 (N_12731,N_11547,N_11711);
or U12732 (N_12732,N_11965,N_12321);
and U12733 (N_12733,N_11641,N_11907);
nor U12734 (N_12734,N_11950,N_12184);
xnor U12735 (N_12735,N_12341,N_11835);
nor U12736 (N_12736,N_11704,N_11277);
or U12737 (N_12737,N_12290,N_11836);
and U12738 (N_12738,N_11892,N_11282);
xnor U12739 (N_12739,N_12120,N_11972);
or U12740 (N_12740,N_12349,N_11508);
and U12741 (N_12741,N_12259,N_12063);
or U12742 (N_12742,N_12465,N_11596);
xnor U12743 (N_12743,N_11616,N_11485);
and U12744 (N_12744,N_11533,N_12182);
nand U12745 (N_12745,N_12416,N_12117);
nand U12746 (N_12746,N_12095,N_12363);
and U12747 (N_12747,N_11534,N_11364);
and U12748 (N_12748,N_11309,N_12342);
nand U12749 (N_12749,N_12208,N_11657);
and U12750 (N_12750,N_11953,N_12395);
or U12751 (N_12751,N_11684,N_11739);
nor U12752 (N_12752,N_11285,N_11380);
or U12753 (N_12753,N_12308,N_11555);
nand U12754 (N_12754,N_12313,N_11845);
nor U12755 (N_12755,N_11459,N_11933);
xnor U12756 (N_12756,N_11814,N_12440);
and U12757 (N_12757,N_11347,N_12437);
nor U12758 (N_12758,N_12428,N_11758);
xnor U12759 (N_12759,N_11780,N_12034);
nand U12760 (N_12760,N_12454,N_12337);
xor U12761 (N_12761,N_11431,N_11888);
nand U12762 (N_12762,N_11978,N_11628);
nor U12763 (N_12763,N_11916,N_11723);
or U12764 (N_12764,N_12012,N_12157);
nand U12765 (N_12765,N_11280,N_12173);
xor U12766 (N_12766,N_11686,N_11955);
nand U12767 (N_12767,N_11349,N_12386);
or U12768 (N_12768,N_11819,N_12242);
nor U12769 (N_12769,N_11573,N_12486);
xor U12770 (N_12770,N_11551,N_11841);
or U12771 (N_12771,N_12002,N_12319);
nand U12772 (N_12772,N_11752,N_12005);
or U12773 (N_12773,N_11827,N_11499);
or U12774 (N_12774,N_11472,N_12370);
nand U12775 (N_12775,N_11331,N_11830);
nor U12776 (N_12776,N_11278,N_12377);
or U12777 (N_12777,N_12361,N_12085);
or U12778 (N_12778,N_11713,N_11873);
nor U12779 (N_12779,N_11832,N_11670);
nor U12780 (N_12780,N_11250,N_12241);
or U12781 (N_12781,N_12485,N_11468);
nand U12782 (N_12782,N_11525,N_12354);
nor U12783 (N_12783,N_11994,N_11668);
and U12784 (N_12784,N_12306,N_12126);
nor U12785 (N_12785,N_12422,N_12166);
or U12786 (N_12786,N_12178,N_12403);
nand U12787 (N_12787,N_12252,N_12061);
xnor U12788 (N_12788,N_12331,N_12000);
and U12789 (N_12789,N_11303,N_12183);
nor U12790 (N_12790,N_11495,N_11486);
nand U12791 (N_12791,N_11389,N_11304);
nand U12792 (N_12792,N_11466,N_11995);
nand U12793 (N_12793,N_12035,N_11712);
nand U12794 (N_12794,N_11602,N_11669);
xor U12795 (N_12795,N_12078,N_12418);
and U12796 (N_12796,N_11361,N_12410);
nor U12797 (N_12797,N_11576,N_11266);
nand U12798 (N_12798,N_12059,N_11678);
nor U12799 (N_12799,N_12488,N_11344);
nand U12800 (N_12800,N_12327,N_12213);
xor U12801 (N_12801,N_12129,N_11425);
xor U12802 (N_12802,N_11549,N_11673);
and U12803 (N_12803,N_12134,N_11388);
nand U12804 (N_12804,N_12033,N_11257);
nand U12805 (N_12805,N_11964,N_12024);
and U12806 (N_12806,N_11510,N_12281);
or U12807 (N_12807,N_12390,N_11849);
xor U12808 (N_12808,N_11607,N_11446);
and U12809 (N_12809,N_12165,N_12351);
nor U12810 (N_12810,N_12498,N_11377);
and U12811 (N_12811,N_12090,N_11579);
nor U12812 (N_12812,N_11647,N_12041);
xor U12813 (N_12813,N_11420,N_11705);
xnor U12814 (N_12814,N_11404,N_11439);
xnor U12815 (N_12815,N_12419,N_11882);
nand U12816 (N_12816,N_12217,N_12472);
nand U12817 (N_12817,N_11688,N_12197);
or U12818 (N_12818,N_11908,N_12018);
or U12819 (N_12819,N_12248,N_12374);
nand U12820 (N_12820,N_12417,N_12116);
and U12821 (N_12821,N_12232,N_12286);
xnor U12822 (N_12822,N_11611,N_11340);
nor U12823 (N_12823,N_11422,N_11333);
or U12824 (N_12824,N_12325,N_12274);
or U12825 (N_12825,N_11585,N_11690);
nand U12826 (N_12826,N_11817,N_11411);
nand U12827 (N_12827,N_11798,N_12398);
xnor U12828 (N_12828,N_11656,N_12322);
nand U12829 (N_12829,N_12412,N_11359);
nand U12830 (N_12830,N_11850,N_11443);
nand U12831 (N_12831,N_12069,N_11258);
and U12832 (N_12832,N_11639,N_11398);
or U12833 (N_12833,N_12229,N_11613);
and U12834 (N_12834,N_11626,N_11651);
xor U12835 (N_12835,N_12466,N_12287);
or U12836 (N_12836,N_11854,N_12442);
nand U12837 (N_12837,N_11637,N_11809);
nand U12838 (N_12838,N_12139,N_12104);
and U12839 (N_12839,N_11320,N_11703);
xor U12840 (N_12840,N_11592,N_12214);
nand U12841 (N_12841,N_12392,N_12393);
or U12842 (N_12842,N_12102,N_11735);
xnor U12843 (N_12843,N_12105,N_11441);
and U12844 (N_12844,N_11923,N_11527);
nor U12845 (N_12845,N_11519,N_11327);
nand U12846 (N_12846,N_11783,N_12047);
xor U12847 (N_12847,N_11867,N_11858);
and U12848 (N_12848,N_12149,N_11878);
nand U12849 (N_12849,N_12298,N_12201);
nand U12850 (N_12850,N_11976,N_11537);
or U12851 (N_12851,N_12456,N_12278);
xor U12852 (N_12852,N_12191,N_11702);
nor U12853 (N_12853,N_12366,N_11934);
nand U12854 (N_12854,N_12247,N_12203);
and U12855 (N_12855,N_12239,N_12406);
and U12856 (N_12856,N_11689,N_11625);
and U12857 (N_12857,N_12355,N_11479);
xor U12858 (N_12858,N_11475,N_12020);
or U12859 (N_12859,N_12081,N_12441);
or U12860 (N_12860,N_11904,N_11580);
and U12861 (N_12861,N_11374,N_11482);
or U12862 (N_12862,N_12153,N_11627);
nand U12863 (N_12863,N_11744,N_12160);
nor U12864 (N_12864,N_12076,N_12080);
or U12865 (N_12865,N_11259,N_12487);
and U12866 (N_12866,N_12170,N_11371);
and U12867 (N_12867,N_11710,N_12399);
nand U12868 (N_12868,N_12176,N_11437);
xor U12869 (N_12869,N_11483,N_11789);
and U12870 (N_12870,N_11314,N_12425);
and U12871 (N_12871,N_12190,N_11718);
nand U12872 (N_12872,N_11820,N_12017);
nand U12873 (N_12873,N_11598,N_11968);
xnor U12874 (N_12874,N_11833,N_12346);
xnor U12875 (N_12875,N_11452,N_11900);
or U12876 (N_12876,N_11383,N_12344);
nor U12877 (N_12877,N_12096,N_12491);
and U12878 (N_12878,N_12409,N_11312);
nand U12879 (N_12879,N_12230,N_11360);
nor U12880 (N_12880,N_11709,N_11937);
or U12881 (N_12881,N_12262,N_11772);
xnor U12882 (N_12882,N_11825,N_12427);
nor U12883 (N_12883,N_11660,N_11815);
nand U12884 (N_12884,N_11988,N_12332);
xor U12885 (N_12885,N_11469,N_11269);
nor U12886 (N_12886,N_11792,N_12243);
or U12887 (N_12887,N_12167,N_11893);
xor U12888 (N_12888,N_11373,N_12050);
nand U12889 (N_12889,N_11914,N_11587);
and U12890 (N_12890,N_12291,N_12376);
nand U12891 (N_12891,N_12192,N_12091);
nor U12892 (N_12892,N_11255,N_12271);
or U12893 (N_12893,N_11513,N_11979);
xor U12894 (N_12894,N_12067,N_11782);
or U12895 (N_12895,N_11942,N_11787);
and U12896 (N_12896,N_11463,N_11332);
or U12897 (N_12897,N_11407,N_11685);
and U12898 (N_12898,N_11778,N_11693);
or U12899 (N_12899,N_12040,N_11572);
and U12900 (N_12900,N_11729,N_12338);
or U12901 (N_12901,N_11805,N_12365);
nor U12902 (N_12902,N_12304,N_12036);
nand U12903 (N_12903,N_12458,N_11894);
xnor U12904 (N_12904,N_11395,N_11256);
or U12905 (N_12905,N_11974,N_11491);
nor U12906 (N_12906,N_11461,N_11631);
or U12907 (N_12907,N_12082,N_11829);
and U12908 (N_12908,N_11590,N_11341);
or U12909 (N_12909,N_11409,N_12079);
nand U12910 (N_12910,N_12089,N_12296);
xor U12911 (N_12911,N_11575,N_11497);
xor U12912 (N_12912,N_11940,N_11741);
and U12913 (N_12913,N_11943,N_11274);
xnor U12914 (N_12914,N_12499,N_11912);
or U12915 (N_12915,N_11529,N_11804);
or U12916 (N_12916,N_11276,N_11970);
nand U12917 (N_12917,N_11921,N_11936);
nor U12918 (N_12918,N_12152,N_11748);
and U12919 (N_12919,N_11496,N_11514);
and U12920 (N_12920,N_11622,N_11675);
and U12921 (N_12921,N_11927,N_11428);
xor U12922 (N_12922,N_12279,N_12334);
nand U12923 (N_12923,N_12300,N_11696);
and U12924 (N_12924,N_12046,N_11419);
and U12925 (N_12925,N_12011,N_11251);
nand U12926 (N_12926,N_11536,N_11263);
nand U12927 (N_12927,N_12275,N_12426);
xor U12928 (N_12928,N_11889,N_11728);
or U12929 (N_12929,N_12130,N_11999);
nor U12930 (N_12930,N_11623,N_12171);
nand U12931 (N_12931,N_11808,N_11872);
nor U12932 (N_12932,N_11535,N_12215);
or U12933 (N_12933,N_12150,N_11680);
xor U12934 (N_12934,N_11414,N_11716);
and U12935 (N_12935,N_11947,N_11963);
nand U12936 (N_12936,N_11376,N_11307);
or U12937 (N_12937,N_11324,N_12235);
xnor U12938 (N_12938,N_11679,N_11621);
nand U12939 (N_12939,N_11806,N_11665);
nor U12940 (N_12940,N_11731,N_11559);
nand U12941 (N_12941,N_12008,N_12054);
nor U12942 (N_12942,N_11412,N_12169);
and U12943 (N_12943,N_12177,N_12131);
and U12944 (N_12944,N_11935,N_11456);
or U12945 (N_12945,N_12475,N_11586);
and U12946 (N_12946,N_11408,N_11642);
nor U12947 (N_12947,N_11385,N_11614);
nor U12948 (N_12948,N_12283,N_11885);
nor U12949 (N_12949,N_12404,N_11899);
nor U12950 (N_12950,N_11415,N_11501);
xor U12951 (N_12951,N_11987,N_12133);
nand U12952 (N_12952,N_11301,N_12372);
or U12953 (N_12953,N_11313,N_12420);
nand U12954 (N_12954,N_11818,N_11530);
or U12955 (N_12955,N_11571,N_11261);
or U12956 (N_12956,N_12415,N_11636);
and U12957 (N_12957,N_12030,N_12163);
xor U12958 (N_12958,N_12256,N_12144);
xnor U12959 (N_12959,N_11771,N_12087);
xnor U12960 (N_12960,N_12448,N_11877);
nor U12961 (N_12961,N_11270,N_11747);
nand U12962 (N_12962,N_12263,N_11339);
or U12963 (N_12963,N_11967,N_11945);
xor U12964 (N_12964,N_11667,N_11682);
xor U12965 (N_12965,N_11824,N_11745);
nand U12966 (N_12966,N_11367,N_12051);
or U12967 (N_12967,N_11983,N_11396);
and U12968 (N_12968,N_12257,N_12293);
and U12969 (N_12969,N_12384,N_11794);
xnor U12970 (N_12970,N_11918,N_11939);
nor U12971 (N_12971,N_11887,N_12305);
nor U12972 (N_12972,N_12401,N_11655);
nor U12973 (N_12973,N_12383,N_12009);
nor U12974 (N_12974,N_12112,N_11594);
or U12975 (N_12975,N_11707,N_11253);
or U12976 (N_12976,N_12408,N_12316);
and U12977 (N_12977,N_11465,N_12220);
xnor U12978 (N_12978,N_11560,N_11777);
xnor U12979 (N_12979,N_11659,N_12250);
and U12980 (N_12980,N_11354,N_11717);
and U12981 (N_12981,N_12189,N_12115);
xnor U12982 (N_12982,N_12272,N_11846);
nand U12983 (N_12983,N_11326,N_11316);
nand U12984 (N_12984,N_12381,N_11695);
nand U12985 (N_12985,N_11774,N_11494);
or U12986 (N_12986,N_11754,N_12444);
xnor U12987 (N_12987,N_11577,N_11603);
or U12988 (N_12988,N_12151,N_11558);
nor U12989 (N_12989,N_12022,N_11932);
xnor U12990 (N_12990,N_11691,N_12260);
xnor U12991 (N_12991,N_12391,N_11793);
or U12992 (N_12992,N_11281,N_12107);
or U12993 (N_12993,N_11588,N_12109);
and U12994 (N_12994,N_12038,N_11378);
xnor U12995 (N_12995,N_12015,N_12446);
nor U12996 (N_12996,N_11302,N_12464);
and U12997 (N_12997,N_12100,N_11406);
and U12998 (N_12998,N_12088,N_12424);
or U12999 (N_12999,N_12052,N_11283);
xor U13000 (N_13000,N_11720,N_12314);
or U13001 (N_13001,N_12209,N_11922);
nor U13002 (N_13002,N_12224,N_12288);
or U13003 (N_13003,N_11348,N_11962);
or U13004 (N_13004,N_11448,N_11518);
or U13005 (N_13005,N_12001,N_12496);
nand U13006 (N_13006,N_11517,N_12124);
xor U13007 (N_13007,N_11295,N_11512);
xnor U13008 (N_13008,N_12482,N_11839);
and U13009 (N_13009,N_11604,N_11298);
nand U13010 (N_13010,N_11785,N_11543);
and U13011 (N_13011,N_11890,N_11742);
nor U13012 (N_13012,N_11632,N_12460);
or U13013 (N_13013,N_11606,N_11861);
and U13014 (N_13014,N_12161,N_11645);
or U13015 (N_13015,N_11661,N_11505);
nor U13016 (N_13016,N_12435,N_12255);
nand U13017 (N_13017,N_11357,N_11433);
nor U13018 (N_13018,N_11993,N_12103);
or U13019 (N_13019,N_11816,N_11971);
or U13020 (N_13020,N_12326,N_11834);
nand U13021 (N_13021,N_11597,N_12097);
nor U13022 (N_13022,N_12155,N_12062);
and U13023 (N_13023,N_11581,N_11982);
xor U13024 (N_13024,N_11760,N_12292);
nor U13025 (N_13025,N_11727,N_12205);
xor U13026 (N_13026,N_11325,N_11363);
or U13027 (N_13027,N_12385,N_11489);
nand U13028 (N_13028,N_12309,N_11615);
and U13029 (N_13029,N_11402,N_11664);
or U13030 (N_13030,N_11797,N_12375);
nor U13031 (N_13031,N_11400,N_12421);
or U13032 (N_13032,N_11610,N_11770);
nand U13033 (N_13033,N_11799,N_12350);
xor U13034 (N_13034,N_12357,N_11511);
nand U13035 (N_13035,N_11293,N_11440);
or U13036 (N_13036,N_11949,N_12086);
and U13037 (N_13037,N_11738,N_12123);
nor U13038 (N_13038,N_12053,N_11561);
or U13039 (N_13039,N_11254,N_11957);
nor U13040 (N_13040,N_11565,N_11719);
nand U13041 (N_13041,N_12289,N_12193);
or U13042 (N_13042,N_11538,N_11746);
or U13043 (N_13043,N_12246,N_12132);
nand U13044 (N_13044,N_11868,N_11843);
or U13045 (N_13045,N_12065,N_11308);
nor U13046 (N_13046,N_12113,N_11328);
xor U13047 (N_13047,N_11394,N_12010);
nand U13048 (N_13048,N_12099,N_12199);
nor U13049 (N_13049,N_12294,N_12347);
nor U13050 (N_13050,N_11507,N_12494);
nor U13051 (N_13051,N_11455,N_11708);
nand U13052 (N_13052,N_11851,N_11397);
nand U13053 (N_13053,N_11644,N_11802);
nor U13054 (N_13054,N_11352,N_11946);
nand U13055 (N_13055,N_12495,N_11288);
or U13056 (N_13056,N_12037,N_12302);
xor U13057 (N_13057,N_11442,N_11321);
or U13058 (N_13058,N_12297,N_12402);
nand U13059 (N_13059,N_11273,N_11355);
nor U13060 (N_13060,N_11490,N_11930);
or U13061 (N_13061,N_12200,N_12356);
xor U13062 (N_13062,N_12055,N_11599);
and U13063 (N_13063,N_11391,N_11343);
xor U13064 (N_13064,N_11895,N_12414);
and U13065 (N_13065,N_11593,N_11764);
xnor U13066 (N_13066,N_11903,N_11375);
and U13067 (N_13067,N_11807,N_12162);
and U13068 (N_13068,N_11991,N_12371);
or U13069 (N_13069,N_11531,N_11800);
or U13070 (N_13070,N_12154,N_11504);
nand U13071 (N_13071,N_12429,N_11981);
nand U13072 (N_13072,N_11345,N_11605);
xnor U13073 (N_13073,N_11755,N_12497);
or U13074 (N_13074,N_12125,N_11322);
nor U13075 (N_13075,N_11791,N_11860);
or U13076 (N_13076,N_11305,N_12407);
xnor U13077 (N_13077,N_11275,N_12405);
nand U13078 (N_13078,N_11539,N_11563);
xor U13079 (N_13079,N_11880,N_12261);
or U13080 (N_13080,N_11471,N_11417);
or U13081 (N_13081,N_11548,N_12135);
nor U13082 (N_13082,N_11743,N_12336);
xnor U13083 (N_13083,N_12353,N_11677);
and U13084 (N_13084,N_11502,N_12204);
nand U13085 (N_13085,N_11264,N_11379);
or U13086 (N_13086,N_11336,N_11492);
nand U13087 (N_13087,N_11649,N_12156);
xnor U13088 (N_13088,N_11931,N_11358);
or U13089 (N_13089,N_11822,N_11524);
and U13090 (N_13090,N_12119,N_11897);
nor U13091 (N_13091,N_12014,N_11740);
nand U13092 (N_13092,N_11919,N_12285);
nand U13093 (N_13093,N_11788,N_12027);
xnor U13094 (N_13094,N_11319,N_11863);
and U13095 (N_13095,N_11401,N_11410);
xor U13096 (N_13096,N_12315,N_11648);
nand U13097 (N_13097,N_12438,N_12194);
xnor U13098 (N_13098,N_11803,N_12423);
nand U13099 (N_13099,N_11671,N_11698);
nor U13100 (N_13100,N_11654,N_11591);
nor U13101 (N_13101,N_11775,N_11977);
xor U13102 (N_13102,N_12490,N_11821);
nor U13103 (N_13103,N_11434,N_12273);
or U13104 (N_13104,N_11286,N_12431);
nand U13105 (N_13105,N_11653,N_12436);
nand U13106 (N_13106,N_12083,N_11297);
xnor U13107 (N_13107,N_11924,N_12226);
and U13108 (N_13108,N_12268,N_11457);
nand U13109 (N_13109,N_12312,N_12026);
nor U13110 (N_13110,N_12468,N_12358);
or U13111 (N_13111,N_12013,N_11279);
xnor U13112 (N_13112,N_12019,N_12462);
nor U13113 (N_13113,N_11284,N_12310);
or U13114 (N_13114,N_11666,N_12077);
or U13115 (N_13115,N_11521,N_12236);
nand U13116 (N_13116,N_12092,N_11768);
xnor U13117 (N_13117,N_11612,N_12264);
nand U13118 (N_13118,N_12245,N_12411);
xor U13119 (N_13119,N_12389,N_12258);
and U13120 (N_13120,N_11523,N_11640);
and U13121 (N_13121,N_12362,N_11992);
nor U13122 (N_13122,N_11891,N_11762);
nor U13123 (N_13123,N_11886,N_11761);
xor U13124 (N_13124,N_12231,N_11267);
and U13125 (N_13125,N_11574,N_12110);
xnor U13126 (N_13126,N_12105,N_11303);
nand U13127 (N_13127,N_12212,N_11495);
and U13128 (N_13128,N_12159,N_12458);
and U13129 (N_13129,N_11773,N_11277);
and U13130 (N_13130,N_12461,N_11543);
or U13131 (N_13131,N_12153,N_11353);
nor U13132 (N_13132,N_11280,N_12367);
or U13133 (N_13133,N_12115,N_12478);
or U13134 (N_13134,N_11673,N_12083);
and U13135 (N_13135,N_12479,N_11551);
and U13136 (N_13136,N_11320,N_11429);
and U13137 (N_13137,N_11692,N_11649);
and U13138 (N_13138,N_11279,N_12461);
nand U13139 (N_13139,N_12096,N_12095);
nand U13140 (N_13140,N_12247,N_11980);
nor U13141 (N_13141,N_11688,N_12352);
nand U13142 (N_13142,N_11430,N_11556);
and U13143 (N_13143,N_11879,N_11903);
nor U13144 (N_13144,N_12150,N_11504);
nand U13145 (N_13145,N_11583,N_11713);
xnor U13146 (N_13146,N_11560,N_12176);
and U13147 (N_13147,N_12206,N_11865);
nand U13148 (N_13148,N_11798,N_12268);
nand U13149 (N_13149,N_12479,N_12431);
or U13150 (N_13150,N_11664,N_11602);
nand U13151 (N_13151,N_11361,N_11476);
xnor U13152 (N_13152,N_12252,N_11324);
nor U13153 (N_13153,N_11723,N_12390);
nor U13154 (N_13154,N_12199,N_12450);
nand U13155 (N_13155,N_12086,N_12459);
nor U13156 (N_13156,N_11959,N_12020);
or U13157 (N_13157,N_12354,N_12464);
and U13158 (N_13158,N_11531,N_11692);
or U13159 (N_13159,N_12479,N_11469);
xnor U13160 (N_13160,N_11333,N_11357);
nor U13161 (N_13161,N_11735,N_11638);
nand U13162 (N_13162,N_12371,N_12162);
nor U13163 (N_13163,N_11731,N_11669);
or U13164 (N_13164,N_11978,N_12471);
xor U13165 (N_13165,N_11920,N_11983);
or U13166 (N_13166,N_11407,N_11490);
nand U13167 (N_13167,N_11913,N_12398);
nand U13168 (N_13168,N_12203,N_12367);
nand U13169 (N_13169,N_11693,N_12366);
nand U13170 (N_13170,N_11421,N_11899);
or U13171 (N_13171,N_11789,N_11446);
nor U13172 (N_13172,N_11776,N_12427);
nor U13173 (N_13173,N_11923,N_11679);
xnor U13174 (N_13174,N_11362,N_12368);
xor U13175 (N_13175,N_11527,N_11570);
and U13176 (N_13176,N_11673,N_11461);
nor U13177 (N_13177,N_11983,N_11930);
nor U13178 (N_13178,N_12031,N_12460);
xnor U13179 (N_13179,N_11847,N_12062);
nor U13180 (N_13180,N_11569,N_11290);
nand U13181 (N_13181,N_11463,N_12107);
or U13182 (N_13182,N_12228,N_12250);
nand U13183 (N_13183,N_11959,N_12076);
nor U13184 (N_13184,N_11624,N_12375);
nand U13185 (N_13185,N_11538,N_11590);
nand U13186 (N_13186,N_12134,N_11595);
and U13187 (N_13187,N_12273,N_12345);
nand U13188 (N_13188,N_11263,N_11419);
or U13189 (N_13189,N_12214,N_11279);
and U13190 (N_13190,N_11623,N_11923);
nor U13191 (N_13191,N_11599,N_11938);
and U13192 (N_13192,N_11564,N_11294);
or U13193 (N_13193,N_11325,N_11339);
nand U13194 (N_13194,N_11343,N_11974);
nand U13195 (N_13195,N_11418,N_11646);
and U13196 (N_13196,N_12112,N_11675);
xor U13197 (N_13197,N_11626,N_11945);
nand U13198 (N_13198,N_11934,N_11976);
or U13199 (N_13199,N_12148,N_11937);
nor U13200 (N_13200,N_12491,N_12445);
xor U13201 (N_13201,N_11757,N_12245);
nor U13202 (N_13202,N_11598,N_12090);
or U13203 (N_13203,N_12252,N_11514);
xnor U13204 (N_13204,N_12160,N_12382);
and U13205 (N_13205,N_12302,N_11840);
nor U13206 (N_13206,N_11801,N_11607);
nor U13207 (N_13207,N_12214,N_12251);
nor U13208 (N_13208,N_11570,N_11705);
and U13209 (N_13209,N_11738,N_11541);
nand U13210 (N_13210,N_12297,N_11661);
nor U13211 (N_13211,N_11935,N_11266);
and U13212 (N_13212,N_11904,N_11449);
or U13213 (N_13213,N_11254,N_12436);
nor U13214 (N_13214,N_11812,N_11649);
or U13215 (N_13215,N_11281,N_12089);
and U13216 (N_13216,N_12313,N_11386);
nor U13217 (N_13217,N_12052,N_12390);
xor U13218 (N_13218,N_11316,N_11441);
or U13219 (N_13219,N_11334,N_11840);
xor U13220 (N_13220,N_11981,N_11772);
xnor U13221 (N_13221,N_11977,N_11815);
xnor U13222 (N_13222,N_11941,N_11841);
or U13223 (N_13223,N_11738,N_12153);
and U13224 (N_13224,N_11270,N_11401);
nor U13225 (N_13225,N_12250,N_12075);
xor U13226 (N_13226,N_12294,N_11741);
and U13227 (N_13227,N_11293,N_11951);
nor U13228 (N_13228,N_11719,N_11805);
nor U13229 (N_13229,N_12163,N_11358);
and U13230 (N_13230,N_11640,N_11686);
nand U13231 (N_13231,N_12248,N_11604);
nor U13232 (N_13232,N_11964,N_12232);
or U13233 (N_13233,N_11848,N_12132);
nor U13234 (N_13234,N_11621,N_11720);
and U13235 (N_13235,N_11697,N_11819);
and U13236 (N_13236,N_11705,N_12129);
and U13237 (N_13237,N_11733,N_11865);
xor U13238 (N_13238,N_12036,N_11453);
or U13239 (N_13239,N_11780,N_12184);
nand U13240 (N_13240,N_11903,N_12124);
nor U13241 (N_13241,N_12476,N_11670);
or U13242 (N_13242,N_12151,N_11396);
and U13243 (N_13243,N_11587,N_12119);
and U13244 (N_13244,N_11767,N_12201);
or U13245 (N_13245,N_11568,N_11998);
and U13246 (N_13246,N_12117,N_12087);
or U13247 (N_13247,N_11852,N_11516);
and U13248 (N_13248,N_11676,N_11398);
and U13249 (N_13249,N_11524,N_11981);
nor U13250 (N_13250,N_12342,N_11424);
xor U13251 (N_13251,N_12028,N_11670);
nand U13252 (N_13252,N_11490,N_12305);
nor U13253 (N_13253,N_12495,N_11434);
or U13254 (N_13254,N_11586,N_11548);
nor U13255 (N_13255,N_11298,N_12357);
nand U13256 (N_13256,N_12336,N_12384);
nand U13257 (N_13257,N_12086,N_11470);
nand U13258 (N_13258,N_11631,N_12491);
nor U13259 (N_13259,N_11667,N_11540);
xor U13260 (N_13260,N_11364,N_11527);
and U13261 (N_13261,N_12180,N_12259);
or U13262 (N_13262,N_11898,N_11439);
nor U13263 (N_13263,N_11686,N_11550);
xnor U13264 (N_13264,N_12037,N_12028);
nand U13265 (N_13265,N_11311,N_11420);
nor U13266 (N_13266,N_12072,N_11630);
xor U13267 (N_13267,N_12404,N_11266);
and U13268 (N_13268,N_11803,N_11662);
nor U13269 (N_13269,N_11729,N_12322);
or U13270 (N_13270,N_11322,N_12318);
or U13271 (N_13271,N_11989,N_11503);
nor U13272 (N_13272,N_11848,N_11618);
or U13273 (N_13273,N_12064,N_11596);
xnor U13274 (N_13274,N_12215,N_11851);
nand U13275 (N_13275,N_12288,N_12011);
or U13276 (N_13276,N_12419,N_11659);
or U13277 (N_13277,N_11991,N_11851);
xnor U13278 (N_13278,N_12474,N_12489);
xnor U13279 (N_13279,N_11567,N_12150);
xor U13280 (N_13280,N_12023,N_11673);
nor U13281 (N_13281,N_12444,N_11808);
and U13282 (N_13282,N_11494,N_12497);
xor U13283 (N_13283,N_12473,N_11827);
xor U13284 (N_13284,N_12166,N_12026);
or U13285 (N_13285,N_11706,N_11836);
nor U13286 (N_13286,N_11917,N_11313);
nand U13287 (N_13287,N_11768,N_11285);
nand U13288 (N_13288,N_11952,N_11302);
or U13289 (N_13289,N_12326,N_11283);
and U13290 (N_13290,N_11881,N_12233);
nand U13291 (N_13291,N_11375,N_12254);
or U13292 (N_13292,N_11538,N_11321);
and U13293 (N_13293,N_12329,N_11565);
or U13294 (N_13294,N_12061,N_11815);
nand U13295 (N_13295,N_11649,N_12255);
or U13296 (N_13296,N_11473,N_11462);
nor U13297 (N_13297,N_11934,N_12201);
and U13298 (N_13298,N_11668,N_12255);
nand U13299 (N_13299,N_11648,N_11971);
nand U13300 (N_13300,N_12208,N_11465);
and U13301 (N_13301,N_12312,N_11775);
and U13302 (N_13302,N_11353,N_11480);
xor U13303 (N_13303,N_11508,N_11741);
nand U13304 (N_13304,N_11817,N_11324);
and U13305 (N_13305,N_11511,N_11263);
and U13306 (N_13306,N_11793,N_12312);
or U13307 (N_13307,N_11375,N_11368);
nor U13308 (N_13308,N_12180,N_11327);
and U13309 (N_13309,N_12191,N_12395);
or U13310 (N_13310,N_11806,N_12042);
nand U13311 (N_13311,N_11593,N_12042);
nor U13312 (N_13312,N_11903,N_11951);
xnor U13313 (N_13313,N_11292,N_11588);
nor U13314 (N_13314,N_12327,N_12047);
or U13315 (N_13315,N_11325,N_12223);
and U13316 (N_13316,N_12202,N_11450);
or U13317 (N_13317,N_12278,N_11314);
nand U13318 (N_13318,N_11435,N_11251);
or U13319 (N_13319,N_11714,N_11689);
and U13320 (N_13320,N_11486,N_12311);
nor U13321 (N_13321,N_11956,N_11396);
or U13322 (N_13322,N_12384,N_11532);
nor U13323 (N_13323,N_11965,N_11444);
and U13324 (N_13324,N_11691,N_12202);
and U13325 (N_13325,N_11506,N_11809);
and U13326 (N_13326,N_11804,N_12429);
and U13327 (N_13327,N_11813,N_12112);
or U13328 (N_13328,N_11425,N_11548);
nor U13329 (N_13329,N_11871,N_12341);
and U13330 (N_13330,N_11476,N_11747);
and U13331 (N_13331,N_11524,N_11451);
nand U13332 (N_13332,N_11381,N_11805);
nor U13333 (N_13333,N_11912,N_11928);
xor U13334 (N_13334,N_11546,N_11266);
and U13335 (N_13335,N_11591,N_12186);
nor U13336 (N_13336,N_12430,N_11813);
nor U13337 (N_13337,N_12004,N_11541);
nor U13338 (N_13338,N_12155,N_12348);
nor U13339 (N_13339,N_12219,N_11988);
nor U13340 (N_13340,N_12425,N_11438);
xnor U13341 (N_13341,N_11713,N_11900);
or U13342 (N_13342,N_11778,N_11583);
nor U13343 (N_13343,N_12139,N_11374);
nand U13344 (N_13344,N_11535,N_11714);
and U13345 (N_13345,N_11714,N_11458);
xor U13346 (N_13346,N_12235,N_11405);
nand U13347 (N_13347,N_11252,N_12169);
nand U13348 (N_13348,N_12166,N_12259);
or U13349 (N_13349,N_11513,N_11250);
xnor U13350 (N_13350,N_12418,N_11908);
xor U13351 (N_13351,N_11671,N_11821);
nand U13352 (N_13352,N_11437,N_11818);
or U13353 (N_13353,N_11282,N_11908);
or U13354 (N_13354,N_11288,N_11893);
xnor U13355 (N_13355,N_12068,N_12169);
nand U13356 (N_13356,N_11573,N_11895);
or U13357 (N_13357,N_11822,N_11692);
nand U13358 (N_13358,N_12400,N_11793);
nor U13359 (N_13359,N_11831,N_11834);
or U13360 (N_13360,N_11594,N_11837);
and U13361 (N_13361,N_11719,N_12061);
xor U13362 (N_13362,N_11943,N_11876);
and U13363 (N_13363,N_12151,N_11560);
nor U13364 (N_13364,N_12413,N_12442);
xnor U13365 (N_13365,N_11406,N_11579);
nor U13366 (N_13366,N_12142,N_12225);
nor U13367 (N_13367,N_11301,N_12468);
nand U13368 (N_13368,N_12321,N_11649);
nor U13369 (N_13369,N_12270,N_11536);
nor U13370 (N_13370,N_11784,N_11663);
or U13371 (N_13371,N_11906,N_12199);
nand U13372 (N_13372,N_11488,N_11391);
nand U13373 (N_13373,N_11999,N_11586);
nand U13374 (N_13374,N_11850,N_11779);
nand U13375 (N_13375,N_11783,N_12323);
nand U13376 (N_13376,N_11547,N_12179);
xor U13377 (N_13377,N_12249,N_12033);
or U13378 (N_13378,N_11959,N_11345);
nor U13379 (N_13379,N_11297,N_11756);
nand U13380 (N_13380,N_11517,N_11752);
and U13381 (N_13381,N_11713,N_11683);
or U13382 (N_13382,N_11678,N_12084);
xnor U13383 (N_13383,N_11534,N_11716);
xnor U13384 (N_13384,N_11269,N_11724);
or U13385 (N_13385,N_11898,N_11479);
xor U13386 (N_13386,N_11792,N_12075);
and U13387 (N_13387,N_11668,N_11504);
xor U13388 (N_13388,N_11686,N_11608);
xnor U13389 (N_13389,N_11917,N_11578);
or U13390 (N_13390,N_12149,N_11477);
xnor U13391 (N_13391,N_12091,N_12306);
xnor U13392 (N_13392,N_12006,N_11647);
nand U13393 (N_13393,N_12346,N_11544);
nand U13394 (N_13394,N_12166,N_12497);
nor U13395 (N_13395,N_11265,N_12308);
and U13396 (N_13396,N_11901,N_11764);
nor U13397 (N_13397,N_12120,N_12250);
or U13398 (N_13398,N_11540,N_11947);
nand U13399 (N_13399,N_11984,N_12218);
nand U13400 (N_13400,N_12201,N_11683);
or U13401 (N_13401,N_12415,N_12325);
or U13402 (N_13402,N_12147,N_11573);
and U13403 (N_13403,N_11322,N_11506);
nand U13404 (N_13404,N_12069,N_11322);
nor U13405 (N_13405,N_12189,N_12025);
or U13406 (N_13406,N_12083,N_11388);
nor U13407 (N_13407,N_11709,N_11583);
xnor U13408 (N_13408,N_11251,N_11802);
xnor U13409 (N_13409,N_12405,N_12109);
xnor U13410 (N_13410,N_12242,N_12290);
xor U13411 (N_13411,N_12190,N_12231);
nor U13412 (N_13412,N_11350,N_11488);
or U13413 (N_13413,N_12365,N_12366);
nor U13414 (N_13414,N_11341,N_11880);
nand U13415 (N_13415,N_12327,N_11819);
nor U13416 (N_13416,N_11310,N_12380);
nor U13417 (N_13417,N_11361,N_11684);
and U13418 (N_13418,N_11931,N_11578);
or U13419 (N_13419,N_11921,N_12206);
and U13420 (N_13420,N_11789,N_11401);
xor U13421 (N_13421,N_11386,N_11403);
or U13422 (N_13422,N_12143,N_11323);
nor U13423 (N_13423,N_12395,N_12024);
and U13424 (N_13424,N_11656,N_11556);
or U13425 (N_13425,N_12015,N_11803);
nor U13426 (N_13426,N_11451,N_11540);
or U13427 (N_13427,N_12029,N_11528);
and U13428 (N_13428,N_12306,N_11434);
and U13429 (N_13429,N_11740,N_11766);
or U13430 (N_13430,N_12048,N_11258);
or U13431 (N_13431,N_11526,N_12188);
nor U13432 (N_13432,N_11633,N_11527);
nand U13433 (N_13433,N_12085,N_11564);
xor U13434 (N_13434,N_12245,N_11461);
xor U13435 (N_13435,N_11391,N_11799);
or U13436 (N_13436,N_12270,N_12414);
or U13437 (N_13437,N_11441,N_12469);
or U13438 (N_13438,N_11789,N_11570);
xor U13439 (N_13439,N_12411,N_11555);
nor U13440 (N_13440,N_11561,N_11383);
xor U13441 (N_13441,N_12404,N_12093);
and U13442 (N_13442,N_12389,N_12168);
xor U13443 (N_13443,N_12089,N_11635);
or U13444 (N_13444,N_11665,N_12023);
xor U13445 (N_13445,N_12451,N_11721);
nand U13446 (N_13446,N_11323,N_11879);
nand U13447 (N_13447,N_11679,N_12070);
xor U13448 (N_13448,N_12072,N_11980);
nor U13449 (N_13449,N_11399,N_12050);
and U13450 (N_13450,N_12466,N_11882);
nor U13451 (N_13451,N_11694,N_11389);
or U13452 (N_13452,N_12099,N_12396);
or U13453 (N_13453,N_11523,N_11614);
nor U13454 (N_13454,N_12167,N_12239);
xor U13455 (N_13455,N_12281,N_12307);
nor U13456 (N_13456,N_12141,N_11686);
or U13457 (N_13457,N_11293,N_11969);
or U13458 (N_13458,N_11621,N_11852);
nor U13459 (N_13459,N_11666,N_11518);
or U13460 (N_13460,N_11714,N_11823);
nand U13461 (N_13461,N_11754,N_11631);
or U13462 (N_13462,N_11683,N_11808);
and U13463 (N_13463,N_11383,N_11388);
nor U13464 (N_13464,N_12286,N_12321);
or U13465 (N_13465,N_11734,N_11351);
nand U13466 (N_13466,N_11620,N_11887);
xor U13467 (N_13467,N_11834,N_11815);
or U13468 (N_13468,N_11252,N_11892);
xor U13469 (N_13469,N_11860,N_11525);
nor U13470 (N_13470,N_12377,N_11591);
or U13471 (N_13471,N_12259,N_11902);
xor U13472 (N_13472,N_11268,N_12306);
nand U13473 (N_13473,N_11970,N_11907);
and U13474 (N_13474,N_12301,N_12142);
nor U13475 (N_13475,N_11465,N_11811);
nand U13476 (N_13476,N_11965,N_11632);
xor U13477 (N_13477,N_11543,N_11908);
and U13478 (N_13478,N_11944,N_12352);
or U13479 (N_13479,N_11847,N_11820);
xnor U13480 (N_13480,N_11836,N_11812);
xor U13481 (N_13481,N_11804,N_12492);
and U13482 (N_13482,N_11489,N_12433);
nor U13483 (N_13483,N_11753,N_11657);
xnor U13484 (N_13484,N_11727,N_11607);
xor U13485 (N_13485,N_12320,N_12020);
nor U13486 (N_13486,N_11577,N_12003);
nand U13487 (N_13487,N_12056,N_12408);
or U13488 (N_13488,N_11586,N_11803);
xnor U13489 (N_13489,N_11601,N_11901);
nand U13490 (N_13490,N_11910,N_11946);
nand U13491 (N_13491,N_12227,N_11554);
and U13492 (N_13492,N_11786,N_11861);
and U13493 (N_13493,N_12293,N_11964);
nor U13494 (N_13494,N_11928,N_11382);
or U13495 (N_13495,N_12240,N_11633);
nand U13496 (N_13496,N_11960,N_12136);
nor U13497 (N_13497,N_12213,N_11314);
and U13498 (N_13498,N_11499,N_12492);
nand U13499 (N_13499,N_12380,N_11669);
or U13500 (N_13500,N_11575,N_11931);
and U13501 (N_13501,N_12252,N_11431);
nand U13502 (N_13502,N_11381,N_12499);
xor U13503 (N_13503,N_11589,N_11393);
nor U13504 (N_13504,N_11287,N_12241);
or U13505 (N_13505,N_11271,N_12041);
xor U13506 (N_13506,N_11539,N_11287);
and U13507 (N_13507,N_11413,N_11648);
and U13508 (N_13508,N_11862,N_11826);
and U13509 (N_13509,N_12352,N_12046);
or U13510 (N_13510,N_11746,N_12098);
and U13511 (N_13511,N_11914,N_11719);
or U13512 (N_13512,N_11339,N_12264);
nor U13513 (N_13513,N_12438,N_12381);
xor U13514 (N_13514,N_11827,N_12470);
xnor U13515 (N_13515,N_11359,N_11372);
nor U13516 (N_13516,N_12253,N_11764);
or U13517 (N_13517,N_12285,N_11908);
and U13518 (N_13518,N_11274,N_12314);
and U13519 (N_13519,N_12359,N_11320);
xnor U13520 (N_13520,N_11716,N_11950);
or U13521 (N_13521,N_12066,N_12184);
or U13522 (N_13522,N_12046,N_11842);
xor U13523 (N_13523,N_11940,N_12025);
or U13524 (N_13524,N_12331,N_11913);
nand U13525 (N_13525,N_11447,N_12232);
nor U13526 (N_13526,N_11413,N_11780);
nand U13527 (N_13527,N_12309,N_11717);
and U13528 (N_13528,N_12395,N_12456);
nor U13529 (N_13529,N_11616,N_11804);
or U13530 (N_13530,N_12407,N_12225);
xnor U13531 (N_13531,N_11790,N_11880);
and U13532 (N_13532,N_11422,N_11366);
or U13533 (N_13533,N_11904,N_12356);
and U13534 (N_13534,N_12184,N_12490);
and U13535 (N_13535,N_11409,N_12404);
and U13536 (N_13536,N_11777,N_12478);
xnor U13537 (N_13537,N_12274,N_12173);
xnor U13538 (N_13538,N_11990,N_11646);
xnor U13539 (N_13539,N_11908,N_12109);
or U13540 (N_13540,N_11953,N_11345);
nand U13541 (N_13541,N_11326,N_11604);
nand U13542 (N_13542,N_11985,N_12037);
nor U13543 (N_13543,N_11378,N_11828);
nor U13544 (N_13544,N_12234,N_12145);
xor U13545 (N_13545,N_12267,N_11649);
and U13546 (N_13546,N_11701,N_11580);
nor U13547 (N_13547,N_12136,N_12150);
xor U13548 (N_13548,N_12166,N_11918);
or U13549 (N_13549,N_11399,N_11526);
nor U13550 (N_13550,N_12353,N_11740);
nor U13551 (N_13551,N_11340,N_11437);
xor U13552 (N_13552,N_12399,N_12471);
or U13553 (N_13553,N_11377,N_12338);
xnor U13554 (N_13554,N_12234,N_11703);
nor U13555 (N_13555,N_11253,N_11703);
xnor U13556 (N_13556,N_12119,N_12392);
or U13557 (N_13557,N_12251,N_11887);
nand U13558 (N_13558,N_11671,N_11599);
nor U13559 (N_13559,N_11454,N_11419);
and U13560 (N_13560,N_11255,N_12082);
xnor U13561 (N_13561,N_12449,N_12081);
and U13562 (N_13562,N_12384,N_12394);
nand U13563 (N_13563,N_11865,N_11875);
xor U13564 (N_13564,N_11674,N_12080);
or U13565 (N_13565,N_12125,N_11408);
and U13566 (N_13566,N_11468,N_11344);
or U13567 (N_13567,N_12003,N_12212);
nand U13568 (N_13568,N_11727,N_11916);
nor U13569 (N_13569,N_11278,N_12174);
nor U13570 (N_13570,N_11443,N_11448);
or U13571 (N_13571,N_11607,N_11377);
xnor U13572 (N_13572,N_12062,N_11369);
or U13573 (N_13573,N_11534,N_12258);
and U13574 (N_13574,N_11300,N_11392);
or U13575 (N_13575,N_11425,N_11707);
or U13576 (N_13576,N_11878,N_12384);
xnor U13577 (N_13577,N_12082,N_12425);
nor U13578 (N_13578,N_12469,N_11462);
nand U13579 (N_13579,N_11690,N_11805);
nor U13580 (N_13580,N_12469,N_12492);
or U13581 (N_13581,N_11603,N_11713);
xnor U13582 (N_13582,N_11291,N_11453);
nand U13583 (N_13583,N_12095,N_12162);
xor U13584 (N_13584,N_11396,N_11282);
and U13585 (N_13585,N_12317,N_12031);
xnor U13586 (N_13586,N_11687,N_12377);
or U13587 (N_13587,N_11822,N_12314);
or U13588 (N_13588,N_11394,N_11837);
nand U13589 (N_13589,N_11599,N_11547);
xor U13590 (N_13590,N_11745,N_11961);
or U13591 (N_13591,N_12140,N_12240);
nor U13592 (N_13592,N_11906,N_11476);
xnor U13593 (N_13593,N_12041,N_12127);
nand U13594 (N_13594,N_12228,N_12302);
or U13595 (N_13595,N_11704,N_12005);
and U13596 (N_13596,N_12016,N_12285);
xnor U13597 (N_13597,N_12356,N_11957);
xnor U13598 (N_13598,N_11371,N_12021);
nor U13599 (N_13599,N_11954,N_11441);
nor U13600 (N_13600,N_11397,N_11834);
and U13601 (N_13601,N_12434,N_11601);
xor U13602 (N_13602,N_11584,N_11310);
or U13603 (N_13603,N_11839,N_11573);
nor U13604 (N_13604,N_11760,N_11553);
and U13605 (N_13605,N_12341,N_12429);
nor U13606 (N_13606,N_12268,N_12289);
and U13607 (N_13607,N_11346,N_12354);
and U13608 (N_13608,N_11872,N_11654);
and U13609 (N_13609,N_12018,N_11959);
nand U13610 (N_13610,N_11527,N_11615);
xor U13611 (N_13611,N_11712,N_12131);
xnor U13612 (N_13612,N_11337,N_11801);
nand U13613 (N_13613,N_12463,N_11988);
xor U13614 (N_13614,N_11479,N_11827);
or U13615 (N_13615,N_11410,N_11373);
or U13616 (N_13616,N_11722,N_12471);
and U13617 (N_13617,N_11575,N_11607);
xnor U13618 (N_13618,N_12230,N_11962);
xor U13619 (N_13619,N_11697,N_11295);
or U13620 (N_13620,N_11659,N_11293);
or U13621 (N_13621,N_12248,N_12113);
xnor U13622 (N_13622,N_11497,N_11787);
and U13623 (N_13623,N_12305,N_11802);
nand U13624 (N_13624,N_11319,N_12017);
or U13625 (N_13625,N_11892,N_11806);
nand U13626 (N_13626,N_11735,N_11394);
nand U13627 (N_13627,N_12348,N_12231);
nand U13628 (N_13628,N_11536,N_11951);
nand U13629 (N_13629,N_11439,N_11742);
nand U13630 (N_13630,N_11801,N_11826);
and U13631 (N_13631,N_11857,N_12232);
xnor U13632 (N_13632,N_11272,N_12282);
xor U13633 (N_13633,N_11552,N_11285);
or U13634 (N_13634,N_11380,N_11530);
nor U13635 (N_13635,N_12196,N_11511);
nand U13636 (N_13636,N_11399,N_12208);
xor U13637 (N_13637,N_12304,N_12415);
nand U13638 (N_13638,N_11356,N_11824);
or U13639 (N_13639,N_11973,N_12481);
and U13640 (N_13640,N_12413,N_12052);
nand U13641 (N_13641,N_12488,N_11581);
or U13642 (N_13642,N_11282,N_12116);
xnor U13643 (N_13643,N_11266,N_11957);
and U13644 (N_13644,N_11512,N_11706);
nand U13645 (N_13645,N_11281,N_11563);
and U13646 (N_13646,N_11782,N_12194);
or U13647 (N_13647,N_11864,N_11678);
nand U13648 (N_13648,N_11336,N_12454);
xor U13649 (N_13649,N_12025,N_12020);
xnor U13650 (N_13650,N_11449,N_12022);
nand U13651 (N_13651,N_12153,N_11944);
nor U13652 (N_13652,N_12199,N_11664);
and U13653 (N_13653,N_11553,N_12013);
xnor U13654 (N_13654,N_11473,N_11648);
nor U13655 (N_13655,N_11976,N_12458);
xor U13656 (N_13656,N_11512,N_12208);
nor U13657 (N_13657,N_11619,N_12219);
and U13658 (N_13658,N_11930,N_11255);
or U13659 (N_13659,N_11798,N_12442);
and U13660 (N_13660,N_12381,N_12057);
and U13661 (N_13661,N_11880,N_12280);
xor U13662 (N_13662,N_11805,N_12124);
xnor U13663 (N_13663,N_11722,N_11488);
nor U13664 (N_13664,N_11398,N_11319);
or U13665 (N_13665,N_12468,N_11809);
nor U13666 (N_13666,N_12479,N_11861);
or U13667 (N_13667,N_12126,N_11628);
nor U13668 (N_13668,N_11798,N_11771);
and U13669 (N_13669,N_12049,N_11574);
nor U13670 (N_13670,N_11397,N_12000);
or U13671 (N_13671,N_11576,N_12089);
or U13672 (N_13672,N_12136,N_12204);
xor U13673 (N_13673,N_12100,N_11573);
xnor U13674 (N_13674,N_12443,N_11406);
nor U13675 (N_13675,N_12348,N_11529);
nand U13676 (N_13676,N_12009,N_11403);
xor U13677 (N_13677,N_11636,N_12098);
xor U13678 (N_13678,N_11850,N_12255);
nor U13679 (N_13679,N_12425,N_12078);
nor U13680 (N_13680,N_11460,N_11639);
nor U13681 (N_13681,N_11954,N_11462);
or U13682 (N_13682,N_11631,N_11902);
or U13683 (N_13683,N_11994,N_12203);
xor U13684 (N_13684,N_11638,N_11818);
xor U13685 (N_13685,N_12464,N_11313);
xor U13686 (N_13686,N_11628,N_12417);
nand U13687 (N_13687,N_11428,N_12145);
or U13688 (N_13688,N_11596,N_11673);
and U13689 (N_13689,N_12046,N_12139);
or U13690 (N_13690,N_11318,N_11714);
nor U13691 (N_13691,N_11990,N_11257);
xor U13692 (N_13692,N_12251,N_11903);
nor U13693 (N_13693,N_11299,N_11731);
xnor U13694 (N_13694,N_12426,N_12283);
xor U13695 (N_13695,N_11923,N_12190);
or U13696 (N_13696,N_11281,N_12254);
nor U13697 (N_13697,N_11500,N_11878);
and U13698 (N_13698,N_11539,N_11837);
or U13699 (N_13699,N_11819,N_12071);
or U13700 (N_13700,N_12333,N_12208);
or U13701 (N_13701,N_11331,N_11777);
nor U13702 (N_13702,N_12011,N_12000);
or U13703 (N_13703,N_11871,N_12386);
nand U13704 (N_13704,N_11940,N_11903);
xnor U13705 (N_13705,N_12112,N_11406);
nor U13706 (N_13706,N_11897,N_11625);
and U13707 (N_13707,N_11296,N_12306);
and U13708 (N_13708,N_12204,N_11659);
nand U13709 (N_13709,N_11462,N_11347);
xor U13710 (N_13710,N_11359,N_11856);
and U13711 (N_13711,N_11918,N_12310);
nor U13712 (N_13712,N_12468,N_11434);
or U13713 (N_13713,N_11612,N_11316);
nor U13714 (N_13714,N_12385,N_11355);
nor U13715 (N_13715,N_11385,N_11973);
or U13716 (N_13716,N_12032,N_12140);
nor U13717 (N_13717,N_11965,N_11764);
xnor U13718 (N_13718,N_11645,N_11777);
nor U13719 (N_13719,N_11517,N_12431);
or U13720 (N_13720,N_12282,N_11969);
xor U13721 (N_13721,N_12477,N_12252);
xnor U13722 (N_13722,N_11876,N_11839);
nor U13723 (N_13723,N_12432,N_12098);
nand U13724 (N_13724,N_12433,N_11362);
or U13725 (N_13725,N_11323,N_11913);
xnor U13726 (N_13726,N_11654,N_11339);
xor U13727 (N_13727,N_12278,N_12336);
or U13728 (N_13728,N_11602,N_12151);
xnor U13729 (N_13729,N_11875,N_11357);
xor U13730 (N_13730,N_11522,N_12303);
or U13731 (N_13731,N_11297,N_11435);
xnor U13732 (N_13732,N_12441,N_12336);
nand U13733 (N_13733,N_11669,N_11685);
xor U13734 (N_13734,N_12405,N_11780);
nor U13735 (N_13735,N_12314,N_12352);
xnor U13736 (N_13736,N_12454,N_11926);
xor U13737 (N_13737,N_11971,N_11542);
nand U13738 (N_13738,N_12271,N_12032);
nand U13739 (N_13739,N_11510,N_12415);
nand U13740 (N_13740,N_11599,N_12149);
nand U13741 (N_13741,N_11779,N_11491);
or U13742 (N_13742,N_12440,N_12188);
and U13743 (N_13743,N_11269,N_11848);
nand U13744 (N_13744,N_11436,N_11679);
nor U13745 (N_13745,N_12287,N_11552);
and U13746 (N_13746,N_12237,N_11514);
and U13747 (N_13747,N_11641,N_11301);
nor U13748 (N_13748,N_12412,N_11942);
nor U13749 (N_13749,N_12288,N_11357);
nor U13750 (N_13750,N_13276,N_12528);
xnor U13751 (N_13751,N_13252,N_13027);
nor U13752 (N_13752,N_13315,N_13083);
xor U13753 (N_13753,N_12606,N_13453);
xor U13754 (N_13754,N_13685,N_13556);
and U13755 (N_13755,N_13074,N_13652);
xnor U13756 (N_13756,N_13360,N_13618);
or U13757 (N_13757,N_13466,N_13290);
nor U13758 (N_13758,N_12775,N_12684);
or U13759 (N_13759,N_13526,N_13624);
or U13760 (N_13760,N_13585,N_13563);
and U13761 (N_13761,N_12961,N_13342);
xor U13762 (N_13762,N_13527,N_13375);
or U13763 (N_13763,N_12573,N_12830);
and U13764 (N_13764,N_13484,N_13345);
nor U13765 (N_13765,N_13031,N_13233);
nor U13766 (N_13766,N_13603,N_13254);
and U13767 (N_13767,N_13644,N_12512);
and U13768 (N_13768,N_13749,N_12691);
or U13769 (N_13769,N_13374,N_12980);
and U13770 (N_13770,N_13009,N_12847);
or U13771 (N_13771,N_13082,N_13543);
nand U13772 (N_13772,N_12553,N_12751);
and U13773 (N_13773,N_13152,N_13525);
and U13774 (N_13774,N_13545,N_12653);
xor U13775 (N_13775,N_12987,N_12682);
or U13776 (N_13776,N_12798,N_13056);
nor U13777 (N_13777,N_12953,N_13447);
xor U13778 (N_13778,N_13000,N_13279);
and U13779 (N_13779,N_13717,N_13210);
xor U13780 (N_13780,N_13109,N_12610);
nor U13781 (N_13781,N_13413,N_13474);
xor U13782 (N_13782,N_13550,N_12647);
and U13783 (N_13783,N_12758,N_12716);
or U13784 (N_13784,N_12575,N_12501);
or U13785 (N_13785,N_13528,N_13204);
xor U13786 (N_13786,N_13215,N_13492);
or U13787 (N_13787,N_13132,N_13005);
xnor U13788 (N_13788,N_12959,N_12895);
nand U13789 (N_13789,N_13054,N_12664);
nor U13790 (N_13790,N_12570,N_13533);
nand U13791 (N_13791,N_12784,N_12527);
nand U13792 (N_13792,N_13145,N_13437);
nor U13793 (N_13793,N_12760,N_13193);
nor U13794 (N_13794,N_13679,N_13277);
xor U13795 (N_13795,N_13274,N_13505);
nand U13796 (N_13796,N_13720,N_13119);
nand U13797 (N_13797,N_13240,N_13257);
or U13798 (N_13798,N_13302,N_13676);
and U13799 (N_13799,N_12652,N_13183);
or U13800 (N_13800,N_12717,N_13017);
nor U13801 (N_13801,N_13021,N_13001);
and U13802 (N_13802,N_12718,N_13120);
or U13803 (N_13803,N_13591,N_12555);
nor U13804 (N_13804,N_13680,N_13620);
xnor U13805 (N_13805,N_13245,N_12627);
and U13806 (N_13806,N_12529,N_12695);
nor U13807 (N_13807,N_12825,N_13593);
xor U13808 (N_13808,N_12506,N_13369);
nand U13809 (N_13809,N_13485,N_13206);
nand U13810 (N_13810,N_12694,N_12663);
or U13811 (N_13811,N_12869,N_13643);
xnor U13812 (N_13812,N_12983,N_13673);
and U13813 (N_13813,N_12856,N_13426);
nor U13814 (N_13814,N_12886,N_13586);
nand U13815 (N_13815,N_12672,N_12614);
nor U13816 (N_13816,N_12697,N_13371);
nor U13817 (N_13817,N_13534,N_12851);
and U13818 (N_13818,N_13154,N_12912);
or U13819 (N_13819,N_13363,N_13216);
nor U13820 (N_13820,N_12777,N_12797);
xor U13821 (N_13821,N_12612,N_13306);
or U13822 (N_13822,N_13364,N_12981);
xnor U13823 (N_13823,N_12843,N_12752);
and U13824 (N_13824,N_12540,N_13509);
nor U13825 (N_13825,N_13303,N_12918);
or U13826 (N_13826,N_13539,N_12715);
or U13827 (N_13827,N_13079,N_13139);
nand U13828 (N_13828,N_13106,N_12988);
and U13829 (N_13829,N_12617,N_13366);
nor U13830 (N_13830,N_13071,N_13128);
xnor U13831 (N_13831,N_13708,N_13450);
or U13832 (N_13832,N_13649,N_13181);
xor U13833 (N_13833,N_13259,N_13008);
xor U13834 (N_13834,N_13331,N_13713);
or U13835 (N_13835,N_13659,N_12638);
xor U13836 (N_13836,N_13177,N_13036);
and U13837 (N_13837,N_13260,N_13495);
or U13838 (N_13838,N_12850,N_13481);
or U13839 (N_13839,N_12542,N_13100);
nand U13840 (N_13840,N_12676,N_13712);
nor U13841 (N_13841,N_13326,N_12552);
nor U13842 (N_13842,N_13115,N_13358);
or U13843 (N_13843,N_13340,N_12789);
nand U13844 (N_13844,N_13404,N_12738);
nand U13845 (N_13845,N_13599,N_13162);
or U13846 (N_13846,N_12649,N_13740);
nand U13847 (N_13847,N_13157,N_13710);
and U13848 (N_13848,N_13304,N_13349);
nor U13849 (N_13849,N_13656,N_12748);
or U13850 (N_13850,N_13235,N_13415);
nor U13851 (N_13851,N_12754,N_13043);
nor U13852 (N_13852,N_13703,N_12931);
or U13853 (N_13853,N_12696,N_12668);
xor U13854 (N_13854,N_13239,N_13727);
and U13855 (N_13855,N_12920,N_13590);
or U13856 (N_13856,N_13488,N_13144);
nand U13857 (N_13857,N_13695,N_12761);
xor U13858 (N_13858,N_12853,N_12858);
nor U13859 (N_13859,N_13524,N_13108);
or U13860 (N_13860,N_13573,N_13531);
and U13861 (N_13861,N_13739,N_13126);
xnor U13862 (N_13862,N_12947,N_12703);
and U13863 (N_13863,N_13323,N_13367);
and U13864 (N_13864,N_13217,N_12729);
nor U13865 (N_13865,N_12873,N_13060);
and U13866 (N_13866,N_13295,N_13732);
and U13867 (N_13867,N_12689,N_12782);
xnor U13868 (N_13868,N_12844,N_13702);
nand U13869 (N_13869,N_13305,N_12616);
and U13870 (N_13870,N_12826,N_13052);
and U13871 (N_13871,N_13149,N_12897);
xnor U13872 (N_13872,N_12513,N_13230);
and U13873 (N_13873,N_12533,N_12769);
or U13874 (N_13874,N_13464,N_13307);
nor U13875 (N_13875,N_13212,N_13407);
nand U13876 (N_13876,N_12724,N_13151);
or U13877 (N_13877,N_12572,N_13111);
or U13878 (N_13878,N_13704,N_13609);
nor U13879 (N_13879,N_12997,N_12966);
nand U13880 (N_13880,N_13461,N_13122);
nor U13881 (N_13881,N_12957,N_13434);
or U13882 (N_13882,N_13642,N_13388);
nor U13883 (N_13883,N_13357,N_13559);
or U13884 (N_13884,N_12887,N_12785);
xnor U13885 (N_13885,N_12547,N_12597);
xnor U13886 (N_13886,N_13365,N_13153);
or U13887 (N_13887,N_13209,N_13133);
xor U13888 (N_13888,N_13146,N_12609);
or U13889 (N_13889,N_13537,N_12965);
nor U13890 (N_13890,N_13150,N_12720);
xor U13891 (N_13891,N_13467,N_13019);
or U13892 (N_13892,N_12815,N_13168);
nand U13893 (N_13893,N_12776,N_12984);
nor U13894 (N_13894,N_12690,N_13701);
xnor U13895 (N_13895,N_13012,N_13377);
or U13896 (N_13896,N_13722,N_13350);
nand U13897 (N_13897,N_13471,N_13243);
xnor U13898 (N_13898,N_12817,N_13334);
or U13899 (N_13899,N_13707,N_13417);
xor U13900 (N_13900,N_13613,N_13747);
or U13901 (N_13901,N_12680,N_12973);
nor U13902 (N_13902,N_13298,N_12801);
xor U13903 (N_13903,N_13013,N_13156);
nor U13904 (N_13904,N_13200,N_12732);
nor U13905 (N_13905,N_12945,N_13744);
nand U13906 (N_13906,N_13194,N_12600);
and U13907 (N_13907,N_12635,N_13422);
xnor U13908 (N_13908,N_12639,N_13011);
or U13909 (N_13909,N_12835,N_12943);
nand U13910 (N_13910,N_12814,N_12833);
and U13911 (N_13911,N_12834,N_13692);
nand U13912 (N_13912,N_13458,N_12950);
nor U13913 (N_13913,N_12505,N_12865);
xor U13914 (N_13914,N_12637,N_12656);
nand U13915 (N_13915,N_13397,N_13072);
or U13916 (N_13916,N_12687,N_13552);
xnor U13917 (N_13917,N_12927,N_12753);
or U13918 (N_13918,N_13654,N_12962);
and U13919 (N_13919,N_13454,N_13657);
nand U13920 (N_13920,N_13287,N_12942);
nor U13921 (N_13921,N_13034,N_13638);
or U13922 (N_13922,N_13045,N_13625);
and U13923 (N_13923,N_13414,N_13251);
nand U13924 (N_13924,N_12793,N_13028);
or U13925 (N_13925,N_13630,N_13443);
nor U13926 (N_13926,N_13570,N_13487);
nor U13927 (N_13927,N_13494,N_13136);
nor U13928 (N_13928,N_12795,N_12561);
xnor U13929 (N_13929,N_13411,N_12813);
nor U13930 (N_13930,N_12708,N_13222);
nor U13931 (N_13931,N_13420,N_13476);
nand U13932 (N_13932,N_13691,N_13285);
xnor U13933 (N_13933,N_13372,N_13339);
and U13934 (N_13934,N_13095,N_12538);
or U13935 (N_13935,N_12891,N_13379);
and U13936 (N_13936,N_13113,N_13463);
and U13937 (N_13937,N_12909,N_13399);
nor U13938 (N_13938,N_12678,N_12580);
nand U13939 (N_13939,N_13275,N_12642);
nand U13940 (N_13940,N_12667,N_12818);
nor U13941 (N_13941,N_12526,N_13147);
nor U13942 (N_13942,N_13538,N_13288);
nand U13943 (N_13943,N_12620,N_13405);
or U13944 (N_13944,N_13265,N_13737);
xnor U13945 (N_13945,N_12866,N_12952);
nand U13946 (N_13946,N_13196,N_12846);
nor U13947 (N_13947,N_12946,N_13557);
or U13948 (N_13948,N_12764,N_12872);
nor U13949 (N_13949,N_13195,N_12935);
nand U13950 (N_13950,N_13301,N_13098);
and U13951 (N_13951,N_12750,N_12601);
nand U13952 (N_13952,N_12670,N_13174);
or U13953 (N_13953,N_12730,N_12675);
nor U13954 (N_13954,N_12829,N_13078);
and U13955 (N_13955,N_13075,N_13632);
or U13956 (N_13956,N_12624,N_12790);
nand U13957 (N_13957,N_12936,N_13601);
or U13958 (N_13958,N_13688,N_12976);
nand U13959 (N_13959,N_13007,N_13448);
nand U13960 (N_13960,N_13127,N_13352);
or U13961 (N_13961,N_13743,N_13410);
nand U13962 (N_13962,N_13587,N_12646);
nor U13963 (N_13963,N_13328,N_13716);
xnor U13964 (N_13964,N_13635,N_13532);
xnor U13965 (N_13965,N_12618,N_13103);
and U13966 (N_13966,N_13333,N_13121);
or U13967 (N_13967,N_12737,N_12692);
or U13968 (N_13968,N_13393,N_13706);
xnor U13969 (N_13969,N_12594,N_13547);
nor U13970 (N_13970,N_12802,N_13663);
or U13971 (N_13971,N_12607,N_13714);
nand U13972 (N_13972,N_13715,N_12993);
xnor U13973 (N_13973,N_13626,N_13497);
xnor U13974 (N_13974,N_12622,N_13387);
xnor U13975 (N_13975,N_13185,N_12581);
nand U13976 (N_13976,N_13610,N_12991);
nor U13977 (N_13977,N_12955,N_12990);
xnor U13978 (N_13978,N_12517,N_13672);
nor U13979 (N_13979,N_13180,N_13023);
xnor U13980 (N_13980,N_13343,N_13700);
nand U13981 (N_13981,N_13611,N_12960);
xnor U13982 (N_13982,N_13456,N_13155);
nor U13983 (N_13983,N_12577,N_12565);
or U13984 (N_13984,N_13359,N_13311);
xnor U13985 (N_13985,N_13172,N_12688);
nor U13986 (N_13986,N_13655,N_12679);
or U13987 (N_13987,N_13517,N_12660);
xnor U13988 (N_13988,N_13175,N_13406);
xnor U13989 (N_13989,N_12623,N_12892);
and U13990 (N_13990,N_13207,N_13548);
or U13991 (N_13991,N_13661,N_13064);
or U13992 (N_13992,N_13272,N_12636);
and U13993 (N_13993,N_13480,N_13390);
and U13994 (N_13994,N_13341,N_13619);
and U13995 (N_13995,N_13068,N_12712);
or U13996 (N_13996,N_13616,N_12763);
nor U13997 (N_13997,N_12655,N_13465);
nand U13998 (N_13998,N_12550,N_12762);
xor U13999 (N_13999,N_12500,N_12852);
nor U14000 (N_14000,N_12605,N_12954);
xnor U14001 (N_14001,N_13634,N_12992);
or U14002 (N_14002,N_13094,N_13629);
and U14003 (N_14003,N_12848,N_13338);
nand U14004 (N_14004,N_13211,N_12574);
xnor U14005 (N_14005,N_13478,N_13502);
nand U14006 (N_14006,N_12779,N_13313);
nor U14007 (N_14007,N_13425,N_12583);
nor U14008 (N_14008,N_13696,N_13114);
nand U14009 (N_14009,N_13429,N_13493);
nand U14010 (N_14010,N_13091,N_13244);
and U14011 (N_14011,N_12564,N_13640);
nor U14012 (N_14012,N_13577,N_13510);
or U14013 (N_14013,N_13419,N_13728);
and U14014 (N_14014,N_13489,N_12863);
nor U14015 (N_14015,N_12736,N_12832);
xor U14016 (N_14016,N_13729,N_12502);
or U14017 (N_14017,N_13442,N_12578);
nor U14018 (N_14018,N_13682,N_13598);
and U14019 (N_14019,N_13173,N_13070);
or U14020 (N_14020,N_13435,N_13310);
nor U14021 (N_14021,N_12780,N_13227);
or U14022 (N_14022,N_13504,N_13131);
or U14023 (N_14023,N_13512,N_13617);
and U14024 (N_14024,N_13581,N_13580);
or U14025 (N_14025,N_12840,N_13316);
and U14026 (N_14026,N_12940,N_13329);
or U14027 (N_14027,N_12928,N_13674);
or U14028 (N_14028,N_13482,N_13612);
and U14029 (N_14029,N_12969,N_13058);
nor U14030 (N_14030,N_13745,N_13440);
xnor U14031 (N_14031,N_12799,N_13469);
or U14032 (N_14032,N_13241,N_12903);
or U14033 (N_14033,N_12948,N_12939);
xnor U14034 (N_14034,N_13123,N_12906);
nand U14035 (N_14035,N_12537,N_12849);
or U14036 (N_14036,N_13541,N_13347);
xnor U14037 (N_14037,N_12979,N_12591);
nor U14038 (N_14038,N_13730,N_12711);
xnor U14039 (N_14039,N_13032,N_13069);
nand U14040 (N_14040,N_13086,N_13294);
and U14041 (N_14041,N_13242,N_13726);
nor U14042 (N_14042,N_12820,N_12706);
xor U14043 (N_14043,N_13403,N_12956);
xnor U14044 (N_14044,N_12563,N_13675);
and U14045 (N_14045,N_13263,N_13699);
nor U14046 (N_14046,N_12598,N_12571);
or U14047 (N_14047,N_13530,N_13565);
nand U14048 (N_14048,N_13041,N_12919);
or U14049 (N_14049,N_13582,N_13600);
nor U14050 (N_14050,N_13690,N_13567);
and U14051 (N_14051,N_12968,N_12800);
and U14052 (N_14052,N_13346,N_13391);
nand U14053 (N_14053,N_13073,N_13639);
or U14054 (N_14054,N_12504,N_13723);
and U14055 (N_14055,N_13020,N_13579);
nand U14056 (N_14056,N_12838,N_13686);
nor U14057 (N_14057,N_12566,N_13725);
or U14058 (N_14058,N_12809,N_13451);
nand U14059 (N_14059,N_12593,N_13327);
and U14060 (N_14060,N_13110,N_13499);
and U14061 (N_14061,N_13293,N_13319);
nand U14062 (N_14062,N_13540,N_13256);
or U14063 (N_14063,N_12876,N_13101);
and U14064 (N_14064,N_12592,N_12805);
and U14065 (N_14065,N_12929,N_13602);
and U14066 (N_14066,N_13394,N_12702);
nand U14067 (N_14067,N_13025,N_13090);
and U14068 (N_14068,N_13189,N_13055);
or U14069 (N_14069,N_13627,N_12974);
and U14070 (N_14070,N_12628,N_12518);
nand U14071 (N_14071,N_13116,N_13169);
nand U14072 (N_14072,N_13164,N_12546);
and U14073 (N_14073,N_13398,N_13412);
or U14074 (N_14074,N_13318,N_12648);
and U14075 (N_14075,N_12665,N_12788);
nand U14076 (N_14076,N_12824,N_13046);
xor U14077 (N_14077,N_12770,N_13588);
nand U14078 (N_14078,N_13436,N_13247);
or U14079 (N_14079,N_13536,N_13158);
xnor U14080 (N_14080,N_13496,N_12878);
or U14081 (N_14081,N_13125,N_13409);
nand U14082 (N_14082,N_12604,N_12905);
xor U14083 (N_14083,N_13067,N_13741);
xnor U14084 (N_14084,N_12860,N_13087);
or U14085 (N_14085,N_12917,N_13026);
xor U14086 (N_14086,N_13354,N_12644);
xnor U14087 (N_14087,N_12633,N_12921);
nand U14088 (N_14088,N_12657,N_12569);
or U14089 (N_14089,N_12567,N_12854);
nor U14090 (N_14090,N_12722,N_13472);
nor U14091 (N_14091,N_12837,N_12701);
nor U14092 (N_14092,N_13568,N_13278);
or U14093 (N_14093,N_13187,N_13376);
nand U14094 (N_14094,N_12756,N_12808);
xnor U14095 (N_14095,N_12559,N_13322);
and U14096 (N_14096,N_13184,N_13416);
nand U14097 (N_14097,N_13002,N_13596);
nand U14098 (N_14098,N_12870,N_13330);
and U14099 (N_14099,N_13284,N_13667);
nor U14100 (N_14100,N_13137,N_12731);
and U14101 (N_14101,N_13253,N_12902);
and U14102 (N_14102,N_13214,N_12503);
or U14103 (N_14103,N_12996,N_12907);
and U14104 (N_14104,N_12705,N_12508);
nor U14105 (N_14105,N_13736,N_12686);
nand U14106 (N_14106,N_12661,N_13006);
nor U14107 (N_14107,N_12629,N_13400);
xnor U14108 (N_14108,N_12796,N_13283);
nor U14109 (N_14109,N_12515,N_12733);
and U14110 (N_14110,N_13192,N_12579);
nor U14111 (N_14111,N_13604,N_12507);
nand U14112 (N_14112,N_12611,N_13261);
xnor U14113 (N_14113,N_13291,N_12932);
nor U14114 (N_14114,N_12710,N_13300);
or U14115 (N_14115,N_13368,N_12619);
nand U14116 (N_14116,N_12524,N_12888);
xnor U14117 (N_14117,N_13191,N_12771);
nor U14118 (N_14118,N_12930,N_13324);
nand U14119 (N_14119,N_13062,N_13024);
and U14120 (N_14120,N_12707,N_12908);
nor U14121 (N_14121,N_12978,N_13402);
nand U14122 (N_14122,N_13418,N_12728);
or U14123 (N_14123,N_13566,N_12744);
xor U14124 (N_14124,N_12934,N_13135);
nor U14125 (N_14125,N_13621,N_12551);
and U14126 (N_14126,N_13520,N_13096);
nor U14127 (N_14127,N_13592,N_13197);
nor U14128 (N_14128,N_13560,N_13445);
nor U14129 (N_14129,N_12742,N_13653);
or U14130 (N_14130,N_13199,N_13507);
nor U14131 (N_14131,N_12781,N_12868);
or U14132 (N_14132,N_13018,N_13554);
or U14133 (N_14133,N_12713,N_13015);
xnor U14134 (N_14134,N_12643,N_13353);
nor U14135 (N_14135,N_12613,N_12774);
xnor U14136 (N_14136,N_12584,N_12971);
nor U14137 (N_14137,N_13694,N_13104);
nand U14138 (N_14138,N_13039,N_13076);
nor U14139 (N_14139,N_13546,N_13665);
xnor U14140 (N_14140,N_13569,N_12944);
and U14141 (N_14141,N_13424,N_13268);
or U14142 (N_14142,N_12759,N_12549);
or U14143 (N_14143,N_12659,N_12650);
nor U14144 (N_14144,N_13143,N_13501);
xor U14145 (N_14145,N_13198,N_12519);
nor U14146 (N_14146,N_13490,N_13430);
or U14147 (N_14147,N_13503,N_12726);
or U14148 (N_14148,N_12864,N_13236);
and U14149 (N_14149,N_13053,N_13178);
nor U14150 (N_14150,N_13061,N_13683);
xor U14151 (N_14151,N_13452,N_13176);
and U14152 (N_14152,N_12882,N_13641);
nor U14153 (N_14153,N_13317,N_13049);
nand U14154 (N_14154,N_13385,N_12958);
nand U14155 (N_14155,N_13583,N_12937);
xnor U14156 (N_14156,N_13022,N_13595);
or U14157 (N_14157,N_13511,N_12915);
nand U14158 (N_14158,N_13670,N_12794);
nand U14159 (N_14159,N_13479,N_13035);
or U14160 (N_14160,N_12674,N_13112);
nor U14161 (N_14161,N_13721,N_12821);
xor U14162 (N_14162,N_13271,N_13491);
or U14163 (N_14163,N_13718,N_13332);
or U14164 (N_14164,N_12884,N_13124);
and U14165 (N_14165,N_12894,N_13042);
or U14166 (N_14166,N_12862,N_13171);
or U14167 (N_14167,N_12735,N_13529);
nor U14168 (N_14168,N_13614,N_13561);
and U14169 (N_14169,N_13220,N_12545);
nand U14170 (N_14170,N_13608,N_12630);
xnor U14171 (N_14171,N_12587,N_12977);
nand U14172 (N_14172,N_12641,N_13255);
xnor U14173 (N_14173,N_12839,N_13188);
nor U14174 (N_14174,N_13645,N_12914);
and U14175 (N_14175,N_12924,N_13202);
or U14176 (N_14176,N_12881,N_13562);
or U14177 (N_14177,N_12938,N_12651);
and U14178 (N_14178,N_13084,N_13709);
nor U14179 (N_14179,N_12812,N_12831);
nand U14180 (N_14180,N_12985,N_13201);
nand U14181 (N_14181,N_13089,N_13698);
or U14182 (N_14182,N_12998,N_12893);
and U14183 (N_14183,N_13282,N_13386);
nand U14184 (N_14184,N_13389,N_12975);
nand U14185 (N_14185,N_12880,N_12514);
and U14186 (N_14186,N_13408,N_13669);
xor U14187 (N_14187,N_13003,N_12995);
nor U14188 (N_14188,N_13299,N_13232);
or U14189 (N_14189,N_13597,N_12807);
and U14190 (N_14190,N_13014,N_13733);
nor U14191 (N_14191,N_12709,N_13134);
nand U14192 (N_14192,N_13179,N_12539);
nand U14193 (N_14193,N_13637,N_13381);
xnor U14194 (N_14194,N_12585,N_12811);
or U14195 (N_14195,N_12520,N_12874);
and U14196 (N_14196,N_13382,N_13362);
xor U14197 (N_14197,N_13130,N_12755);
nand U14198 (N_14198,N_13622,N_13658);
and U14199 (N_14199,N_13099,N_13498);
nand U14200 (N_14200,N_13351,N_12766);
nor U14201 (N_14201,N_13457,N_13088);
nand U14202 (N_14202,N_13544,N_12621);
nand U14203 (N_14203,N_12899,N_12548);
nor U14204 (N_14204,N_13396,N_12857);
nor U14205 (N_14205,N_13395,N_13057);
nor U14206 (N_14206,N_13519,N_12693);
nor U14207 (N_14207,N_13508,N_13384);
nor U14208 (N_14208,N_13065,N_12877);
or U14209 (N_14209,N_13711,N_12964);
nor U14210 (N_14210,N_13421,N_13671);
or U14211 (N_14211,N_13477,N_12525);
nand U14212 (N_14212,N_13459,N_13219);
and U14213 (N_14213,N_12989,N_13129);
or U14214 (N_14214,N_13446,N_13205);
nand U14215 (N_14215,N_13746,N_12522);
nand U14216 (N_14216,N_13428,N_13273);
xnor U14217 (N_14217,N_12836,N_12783);
xor U14218 (N_14218,N_12615,N_12589);
nor U14219 (N_14219,N_13373,N_13607);
nor U14220 (N_14220,N_13037,N_12855);
or U14221 (N_14221,N_13506,N_12677);
nor U14222 (N_14222,N_13281,N_12602);
or U14223 (N_14223,N_13218,N_12509);
and U14224 (N_14224,N_12671,N_13589);
or U14225 (N_14225,N_12595,N_13292);
nor U14226 (N_14226,N_12757,N_13697);
nor U14227 (N_14227,N_13444,N_13684);
nand U14228 (N_14228,N_12510,N_12925);
nor U14229 (N_14229,N_13648,N_13050);
and U14230 (N_14230,N_13325,N_13578);
xor U14231 (N_14231,N_12822,N_12669);
or U14232 (N_14232,N_13564,N_13475);
and U14233 (N_14233,N_12772,N_13160);
xnor U14234 (N_14234,N_13664,N_12913);
or U14235 (N_14235,N_13433,N_13269);
nand U14236 (N_14236,N_12586,N_13383);
nand U14237 (N_14237,N_13280,N_13555);
nand U14238 (N_14238,N_12590,N_12645);
nor U14239 (N_14239,N_13170,N_13576);
nand U14240 (N_14240,N_13237,N_13165);
and U14241 (N_14241,N_13182,N_13225);
nor U14242 (N_14242,N_13030,N_13650);
nor U14243 (N_14243,N_12734,N_13264);
and U14244 (N_14244,N_13572,N_12666);
and U14245 (N_14245,N_12972,N_12768);
and U14246 (N_14246,N_12654,N_13047);
or U14247 (N_14247,N_13623,N_12883);
and U14248 (N_14248,N_12640,N_13378);
nand U14249 (N_14249,N_13748,N_13224);
nor U14250 (N_14250,N_12951,N_13594);
xnor U14251 (N_14251,N_13522,N_13735);
nor U14252 (N_14252,N_13553,N_13483);
nand U14253 (N_14253,N_13551,N_13724);
nor U14254 (N_14254,N_12900,N_12923);
xor U14255 (N_14255,N_12773,N_12632);
nand U14256 (N_14256,N_13033,N_12626);
nand U14257 (N_14257,N_13348,N_13297);
nand U14258 (N_14258,N_13266,N_13431);
nand U14259 (N_14259,N_13606,N_13734);
and U14260 (N_14260,N_12749,N_13051);
or U14261 (N_14261,N_12719,N_13571);
xor U14262 (N_14262,N_12994,N_12896);
and U14263 (N_14263,N_13460,N_12739);
and U14264 (N_14264,N_12791,N_13267);
nand U14265 (N_14265,N_13647,N_12740);
or U14266 (N_14266,N_13141,N_12556);
or U14267 (N_14267,N_13059,N_12700);
xor U14268 (N_14268,N_12534,N_12532);
and U14269 (N_14269,N_12608,N_13248);
nor U14270 (N_14270,N_13668,N_13321);
nand U14271 (N_14271,N_13468,N_12767);
xor U14272 (N_14272,N_12588,N_13662);
nand U14273 (N_14273,N_12658,N_13077);
nand U14274 (N_14274,N_13010,N_13558);
nor U14275 (N_14275,N_13549,N_12554);
xor U14276 (N_14276,N_12949,N_12911);
nor U14277 (N_14277,N_13223,N_13605);
xor U14278 (N_14278,N_12898,N_13441);
xor U14279 (N_14279,N_13270,N_13004);
nand U14280 (N_14280,N_12704,N_13308);
nor U14281 (N_14281,N_13314,N_13633);
or U14282 (N_14282,N_12599,N_12625);
nand U14283 (N_14283,N_13226,N_12541);
nor U14284 (N_14284,N_13651,N_13677);
nand U14285 (N_14285,N_12819,N_13167);
nor U14286 (N_14286,N_13048,N_13742);
or U14287 (N_14287,N_13660,N_13118);
xnor U14288 (N_14288,N_12516,N_13337);
nor U14289 (N_14289,N_12875,N_13515);
or U14290 (N_14290,N_13221,N_13231);
or U14291 (N_14291,N_13615,N_12926);
nor U14292 (N_14292,N_13102,N_12727);
nor U14293 (N_14293,N_12871,N_12699);
xnor U14294 (N_14294,N_13462,N_13190);
xor U14295 (N_14295,N_13470,N_12634);
nand U14296 (N_14296,N_13380,N_13636);
xor U14297 (N_14297,N_12582,N_12859);
and U14298 (N_14298,N_13423,N_13449);
nand U14299 (N_14299,N_13705,N_12890);
xnor U14300 (N_14300,N_13455,N_13105);
xor U14301 (N_14301,N_13085,N_13666);
or U14302 (N_14302,N_13246,N_13081);
xor U14303 (N_14303,N_13262,N_13523);
nand U14304 (N_14304,N_13542,N_12568);
xor U14305 (N_14305,N_12681,N_13029);
nor U14306 (N_14306,N_12714,N_13092);
xnor U14307 (N_14307,N_12673,N_13584);
xor U14308 (N_14308,N_12963,N_13681);
or U14309 (N_14309,N_13689,N_13238);
xnor U14310 (N_14310,N_13335,N_12841);
or U14311 (N_14311,N_12861,N_13370);
nor U14312 (N_14312,N_12787,N_13392);
xor U14313 (N_14313,N_12721,N_13646);
or U14314 (N_14314,N_12816,N_12596);
xor U14315 (N_14315,N_13258,N_13486);
xnor U14316 (N_14316,N_13229,N_13355);
or U14317 (N_14317,N_12778,N_12982);
or U14318 (N_14318,N_13438,N_13163);
xnor U14319 (N_14319,N_13516,N_13063);
nor U14320 (N_14320,N_12662,N_12531);
nor U14321 (N_14321,N_12885,N_12879);
xor U14322 (N_14322,N_13514,N_12922);
nor U14323 (N_14323,N_12970,N_13521);
or U14324 (N_14324,N_13628,N_13312);
and U14325 (N_14325,N_13535,N_13289);
or U14326 (N_14326,N_12746,N_13693);
nand U14327 (N_14327,N_12560,N_12999);
nand U14328 (N_14328,N_12901,N_12723);
xnor U14329 (N_14329,N_13093,N_12530);
nand U14330 (N_14330,N_13148,N_12576);
nand U14331 (N_14331,N_13401,N_13117);
nand U14332 (N_14332,N_13142,N_13687);
nand U14333 (N_14333,N_12867,N_12803);
nand U14334 (N_14334,N_12828,N_12535);
nor U14335 (N_14335,N_13320,N_12792);
nor U14336 (N_14336,N_13080,N_12823);
nor U14337 (N_14337,N_12562,N_12941);
xnor U14338 (N_14338,N_12933,N_13203);
xor U14339 (N_14339,N_13719,N_12967);
nor U14340 (N_14340,N_13286,N_12845);
or U14341 (N_14341,N_13678,N_13336);
xor U14342 (N_14342,N_12986,N_13097);
or U14343 (N_14343,N_12827,N_12557);
xnor U14344 (N_14344,N_12543,N_12889);
and U14345 (N_14345,N_12725,N_13575);
and U14346 (N_14346,N_12521,N_13361);
and U14347 (N_14347,N_13296,N_13427);
xnor U14348 (N_14348,N_12631,N_12743);
xnor U14349 (N_14349,N_12741,N_13166);
nand U14350 (N_14350,N_13140,N_13574);
or U14351 (N_14351,N_12698,N_12523);
nor U14352 (N_14352,N_12842,N_12544);
nand U14353 (N_14353,N_12904,N_13044);
or U14354 (N_14354,N_13161,N_12511);
and U14355 (N_14355,N_13228,N_13731);
nor U14356 (N_14356,N_13016,N_13213);
and U14357 (N_14357,N_12765,N_12810);
or U14358 (N_14358,N_13208,N_13249);
xor U14359 (N_14359,N_13040,N_12910);
nand U14360 (N_14360,N_12536,N_13250);
and U14361 (N_14361,N_13344,N_13473);
nor U14362 (N_14362,N_13738,N_12745);
or U14363 (N_14363,N_12747,N_13518);
or U14364 (N_14364,N_12786,N_12806);
or U14365 (N_14365,N_13234,N_12603);
nand U14366 (N_14366,N_13500,N_13138);
xor U14367 (N_14367,N_13159,N_13186);
xor U14368 (N_14368,N_12916,N_12685);
and U14369 (N_14369,N_12683,N_12804);
xnor U14370 (N_14370,N_13432,N_13066);
xor U14371 (N_14371,N_13107,N_13038);
xnor U14372 (N_14372,N_13513,N_13309);
nor U14373 (N_14373,N_13439,N_13631);
xor U14374 (N_14374,N_12558,N_13356);
nand U14375 (N_14375,N_13355,N_13649);
nor U14376 (N_14376,N_13037,N_13328);
xor U14377 (N_14377,N_12502,N_12636);
nor U14378 (N_14378,N_13102,N_12865);
nor U14379 (N_14379,N_13009,N_13640);
or U14380 (N_14380,N_12873,N_13217);
and U14381 (N_14381,N_12941,N_12543);
and U14382 (N_14382,N_13334,N_12907);
nand U14383 (N_14383,N_13271,N_12871);
and U14384 (N_14384,N_12852,N_12958);
nor U14385 (N_14385,N_12649,N_12719);
nand U14386 (N_14386,N_12996,N_13206);
nor U14387 (N_14387,N_13149,N_12855);
or U14388 (N_14388,N_12976,N_13395);
xor U14389 (N_14389,N_13601,N_13315);
or U14390 (N_14390,N_13315,N_12813);
and U14391 (N_14391,N_13490,N_13606);
nand U14392 (N_14392,N_13694,N_13642);
or U14393 (N_14393,N_13284,N_13496);
nand U14394 (N_14394,N_12681,N_12968);
and U14395 (N_14395,N_13547,N_13532);
xor U14396 (N_14396,N_12853,N_12547);
nand U14397 (N_14397,N_12981,N_12631);
nand U14398 (N_14398,N_13416,N_13038);
and U14399 (N_14399,N_13175,N_12905);
and U14400 (N_14400,N_12522,N_13617);
xor U14401 (N_14401,N_13399,N_13543);
or U14402 (N_14402,N_12752,N_13556);
or U14403 (N_14403,N_13295,N_12669);
nor U14404 (N_14404,N_12957,N_13275);
or U14405 (N_14405,N_13462,N_13454);
or U14406 (N_14406,N_12653,N_13299);
nand U14407 (N_14407,N_12936,N_13522);
xnor U14408 (N_14408,N_13601,N_13101);
nand U14409 (N_14409,N_12723,N_12642);
or U14410 (N_14410,N_12753,N_13109);
and U14411 (N_14411,N_12907,N_13298);
xor U14412 (N_14412,N_12869,N_13728);
or U14413 (N_14413,N_13006,N_13337);
nand U14414 (N_14414,N_13395,N_12736);
xor U14415 (N_14415,N_13521,N_13192);
or U14416 (N_14416,N_13583,N_13381);
xor U14417 (N_14417,N_13709,N_12557);
and U14418 (N_14418,N_12924,N_13590);
xnor U14419 (N_14419,N_13071,N_12633);
or U14420 (N_14420,N_13398,N_12546);
or U14421 (N_14421,N_13415,N_12507);
xnor U14422 (N_14422,N_12679,N_12728);
xnor U14423 (N_14423,N_12891,N_12527);
and U14424 (N_14424,N_13320,N_13451);
and U14425 (N_14425,N_12708,N_12709);
nand U14426 (N_14426,N_13512,N_13454);
or U14427 (N_14427,N_13580,N_13119);
nand U14428 (N_14428,N_13260,N_12725);
xnor U14429 (N_14429,N_13383,N_12744);
xnor U14430 (N_14430,N_13050,N_12510);
nand U14431 (N_14431,N_13509,N_13746);
nor U14432 (N_14432,N_12565,N_13473);
xor U14433 (N_14433,N_12564,N_12710);
xor U14434 (N_14434,N_13709,N_13517);
xnor U14435 (N_14435,N_12533,N_12644);
nor U14436 (N_14436,N_12782,N_13640);
nand U14437 (N_14437,N_13338,N_13146);
or U14438 (N_14438,N_13505,N_13039);
and U14439 (N_14439,N_12595,N_12935);
or U14440 (N_14440,N_13206,N_12744);
xnor U14441 (N_14441,N_12957,N_12920);
nand U14442 (N_14442,N_12924,N_12538);
xnor U14443 (N_14443,N_12669,N_13580);
or U14444 (N_14444,N_12841,N_12881);
and U14445 (N_14445,N_12556,N_13172);
or U14446 (N_14446,N_13708,N_13409);
nand U14447 (N_14447,N_12979,N_12576);
or U14448 (N_14448,N_13538,N_13343);
nand U14449 (N_14449,N_13561,N_13518);
xnor U14450 (N_14450,N_12600,N_12967);
xnor U14451 (N_14451,N_12579,N_12567);
xnor U14452 (N_14452,N_13003,N_13269);
nand U14453 (N_14453,N_13268,N_13149);
xor U14454 (N_14454,N_13440,N_12589);
or U14455 (N_14455,N_13679,N_13151);
nand U14456 (N_14456,N_13107,N_13415);
or U14457 (N_14457,N_12884,N_12571);
or U14458 (N_14458,N_13583,N_13434);
nand U14459 (N_14459,N_13704,N_12827);
or U14460 (N_14460,N_13475,N_13129);
and U14461 (N_14461,N_13141,N_12885);
xnor U14462 (N_14462,N_13242,N_12932);
or U14463 (N_14463,N_13547,N_13209);
nand U14464 (N_14464,N_13549,N_13135);
nor U14465 (N_14465,N_12711,N_12889);
nor U14466 (N_14466,N_13688,N_13032);
or U14467 (N_14467,N_13729,N_12739);
and U14468 (N_14468,N_12868,N_13711);
nand U14469 (N_14469,N_13742,N_13039);
and U14470 (N_14470,N_13037,N_13630);
xnor U14471 (N_14471,N_13020,N_13701);
xor U14472 (N_14472,N_13509,N_12880);
xnor U14473 (N_14473,N_13026,N_12989);
or U14474 (N_14474,N_13133,N_13135);
nor U14475 (N_14475,N_13546,N_13323);
nor U14476 (N_14476,N_13282,N_12891);
nand U14477 (N_14477,N_12928,N_13727);
xnor U14478 (N_14478,N_12781,N_12656);
nand U14479 (N_14479,N_13153,N_12584);
nand U14480 (N_14480,N_12745,N_13309);
or U14481 (N_14481,N_12838,N_12562);
xnor U14482 (N_14482,N_12502,N_13173);
nor U14483 (N_14483,N_13002,N_12869);
nor U14484 (N_14484,N_12784,N_13357);
nor U14485 (N_14485,N_13641,N_13638);
xnor U14486 (N_14486,N_13636,N_13669);
nand U14487 (N_14487,N_13290,N_13355);
or U14488 (N_14488,N_13525,N_13107);
and U14489 (N_14489,N_12981,N_13570);
nand U14490 (N_14490,N_13635,N_12951);
nand U14491 (N_14491,N_13079,N_13292);
and U14492 (N_14492,N_13565,N_13055);
and U14493 (N_14493,N_13641,N_13191);
nor U14494 (N_14494,N_12910,N_12729);
nand U14495 (N_14495,N_12528,N_13183);
and U14496 (N_14496,N_13631,N_12502);
xor U14497 (N_14497,N_13694,N_13641);
and U14498 (N_14498,N_12649,N_13293);
nor U14499 (N_14499,N_12941,N_12958);
nor U14500 (N_14500,N_13422,N_13076);
and U14501 (N_14501,N_12810,N_12507);
nor U14502 (N_14502,N_13594,N_12810);
xnor U14503 (N_14503,N_12610,N_12864);
nand U14504 (N_14504,N_12647,N_13146);
or U14505 (N_14505,N_13453,N_13282);
nor U14506 (N_14506,N_13190,N_13235);
or U14507 (N_14507,N_13649,N_13648);
or U14508 (N_14508,N_13162,N_13571);
nand U14509 (N_14509,N_13461,N_12834);
or U14510 (N_14510,N_13749,N_12550);
or U14511 (N_14511,N_13367,N_13577);
xnor U14512 (N_14512,N_13682,N_12803);
and U14513 (N_14513,N_13101,N_12602);
nand U14514 (N_14514,N_13713,N_12622);
and U14515 (N_14515,N_13609,N_13327);
and U14516 (N_14516,N_13583,N_12742);
nor U14517 (N_14517,N_13006,N_13296);
xnor U14518 (N_14518,N_13196,N_12712);
nand U14519 (N_14519,N_12983,N_12612);
or U14520 (N_14520,N_12978,N_13452);
or U14521 (N_14521,N_12565,N_13663);
xnor U14522 (N_14522,N_12606,N_13376);
xnor U14523 (N_14523,N_12906,N_13164);
nor U14524 (N_14524,N_13425,N_13095);
nand U14525 (N_14525,N_12587,N_12876);
and U14526 (N_14526,N_13183,N_12849);
or U14527 (N_14527,N_13101,N_12606);
or U14528 (N_14528,N_12787,N_12748);
nand U14529 (N_14529,N_13502,N_12904);
and U14530 (N_14530,N_13156,N_13383);
nor U14531 (N_14531,N_13742,N_12623);
xor U14532 (N_14532,N_13408,N_12657);
xnor U14533 (N_14533,N_12751,N_13649);
xnor U14534 (N_14534,N_13732,N_12586);
nand U14535 (N_14535,N_13748,N_13403);
nand U14536 (N_14536,N_13395,N_13047);
nor U14537 (N_14537,N_13690,N_12615);
nor U14538 (N_14538,N_12791,N_13039);
nand U14539 (N_14539,N_13039,N_13341);
or U14540 (N_14540,N_13030,N_13131);
xnor U14541 (N_14541,N_13255,N_12846);
nand U14542 (N_14542,N_13000,N_13365);
xnor U14543 (N_14543,N_13575,N_13141);
nor U14544 (N_14544,N_12964,N_13472);
and U14545 (N_14545,N_12895,N_13516);
xnor U14546 (N_14546,N_13388,N_13308);
xor U14547 (N_14547,N_13032,N_13744);
or U14548 (N_14548,N_12663,N_13105);
nand U14549 (N_14549,N_13698,N_12900);
nand U14550 (N_14550,N_12877,N_12895);
xnor U14551 (N_14551,N_13537,N_13029);
nor U14552 (N_14552,N_13532,N_13066);
and U14553 (N_14553,N_12829,N_13018);
xnor U14554 (N_14554,N_12635,N_12638);
nand U14555 (N_14555,N_13046,N_13370);
and U14556 (N_14556,N_13160,N_12900);
xnor U14557 (N_14557,N_13449,N_13097);
xnor U14558 (N_14558,N_13459,N_12734);
nor U14559 (N_14559,N_13175,N_13623);
nand U14560 (N_14560,N_12542,N_12841);
nor U14561 (N_14561,N_12552,N_12955);
xnor U14562 (N_14562,N_13004,N_12973);
and U14563 (N_14563,N_12780,N_13178);
nand U14564 (N_14564,N_13002,N_12663);
xnor U14565 (N_14565,N_13634,N_12812);
or U14566 (N_14566,N_12505,N_13103);
nand U14567 (N_14567,N_13602,N_13376);
and U14568 (N_14568,N_13550,N_13627);
nor U14569 (N_14569,N_13479,N_13455);
and U14570 (N_14570,N_13090,N_13203);
nand U14571 (N_14571,N_12847,N_13603);
nand U14572 (N_14572,N_13108,N_13026);
xnor U14573 (N_14573,N_12809,N_13448);
and U14574 (N_14574,N_13250,N_12994);
and U14575 (N_14575,N_12597,N_12635);
and U14576 (N_14576,N_12967,N_12946);
or U14577 (N_14577,N_13596,N_12849);
nor U14578 (N_14578,N_13670,N_12687);
or U14579 (N_14579,N_13717,N_13452);
and U14580 (N_14580,N_12809,N_13367);
nand U14581 (N_14581,N_12859,N_13382);
nand U14582 (N_14582,N_13174,N_12598);
xnor U14583 (N_14583,N_12700,N_12979);
nor U14584 (N_14584,N_12728,N_13225);
nand U14585 (N_14585,N_13464,N_13132);
nand U14586 (N_14586,N_13509,N_12914);
and U14587 (N_14587,N_13535,N_12797);
xor U14588 (N_14588,N_13036,N_13524);
nand U14589 (N_14589,N_12568,N_13285);
nor U14590 (N_14590,N_13599,N_13613);
nor U14591 (N_14591,N_12597,N_13342);
and U14592 (N_14592,N_13138,N_13651);
xor U14593 (N_14593,N_12778,N_13716);
nor U14594 (N_14594,N_13263,N_13142);
or U14595 (N_14595,N_13424,N_12776);
nand U14596 (N_14596,N_13379,N_13362);
nor U14597 (N_14597,N_13728,N_12937);
or U14598 (N_14598,N_12526,N_12512);
nand U14599 (N_14599,N_12859,N_13630);
or U14600 (N_14600,N_12604,N_12573);
nor U14601 (N_14601,N_12552,N_13290);
and U14602 (N_14602,N_12517,N_12832);
and U14603 (N_14603,N_13484,N_13559);
and U14604 (N_14604,N_13663,N_13013);
or U14605 (N_14605,N_12852,N_13276);
or U14606 (N_14606,N_12574,N_13177);
or U14607 (N_14607,N_13412,N_12829);
and U14608 (N_14608,N_13206,N_13432);
and U14609 (N_14609,N_13096,N_12510);
nor U14610 (N_14610,N_13409,N_12580);
nand U14611 (N_14611,N_12550,N_12530);
nand U14612 (N_14612,N_13257,N_13524);
and U14613 (N_14613,N_12990,N_13241);
or U14614 (N_14614,N_12945,N_13207);
or U14615 (N_14615,N_13723,N_13123);
or U14616 (N_14616,N_12673,N_13389);
and U14617 (N_14617,N_13542,N_12659);
nand U14618 (N_14618,N_12932,N_12761);
nand U14619 (N_14619,N_13646,N_13484);
nand U14620 (N_14620,N_13455,N_12984);
xnor U14621 (N_14621,N_12939,N_12652);
xnor U14622 (N_14622,N_13191,N_12992);
xnor U14623 (N_14623,N_13669,N_13154);
or U14624 (N_14624,N_13312,N_13290);
nor U14625 (N_14625,N_13136,N_13595);
xor U14626 (N_14626,N_13572,N_12675);
xnor U14627 (N_14627,N_12711,N_13483);
and U14628 (N_14628,N_13491,N_13333);
xnor U14629 (N_14629,N_13685,N_13338);
or U14630 (N_14630,N_13478,N_12506);
nor U14631 (N_14631,N_13729,N_12709);
or U14632 (N_14632,N_13569,N_13510);
and U14633 (N_14633,N_12671,N_13473);
nand U14634 (N_14634,N_12927,N_13046);
or U14635 (N_14635,N_12813,N_13389);
nor U14636 (N_14636,N_12515,N_13159);
nand U14637 (N_14637,N_13231,N_12716);
or U14638 (N_14638,N_13633,N_13526);
xor U14639 (N_14639,N_13225,N_13713);
nor U14640 (N_14640,N_12583,N_13654);
nand U14641 (N_14641,N_13671,N_13709);
nand U14642 (N_14642,N_13552,N_13186);
xnor U14643 (N_14643,N_12774,N_12877);
nand U14644 (N_14644,N_13134,N_12531);
and U14645 (N_14645,N_13361,N_12552);
nor U14646 (N_14646,N_13012,N_13655);
or U14647 (N_14647,N_13701,N_13081);
nand U14648 (N_14648,N_13478,N_12604);
or U14649 (N_14649,N_12960,N_13177);
nor U14650 (N_14650,N_13593,N_13375);
nor U14651 (N_14651,N_12923,N_12606);
nor U14652 (N_14652,N_12782,N_12800);
nand U14653 (N_14653,N_12830,N_13566);
xnor U14654 (N_14654,N_12905,N_13162);
nand U14655 (N_14655,N_13049,N_12741);
and U14656 (N_14656,N_12554,N_13741);
or U14657 (N_14657,N_13737,N_13694);
or U14658 (N_14658,N_12810,N_13632);
nand U14659 (N_14659,N_12556,N_13112);
and U14660 (N_14660,N_13626,N_13464);
and U14661 (N_14661,N_13369,N_13109);
xor U14662 (N_14662,N_13063,N_13738);
and U14663 (N_14663,N_12975,N_13509);
nor U14664 (N_14664,N_13578,N_13188);
nand U14665 (N_14665,N_12990,N_13537);
or U14666 (N_14666,N_12887,N_12916);
or U14667 (N_14667,N_12726,N_13645);
nand U14668 (N_14668,N_13062,N_13536);
xnor U14669 (N_14669,N_13469,N_12824);
nand U14670 (N_14670,N_12828,N_12779);
or U14671 (N_14671,N_13258,N_13444);
nor U14672 (N_14672,N_12900,N_13019);
xor U14673 (N_14673,N_12840,N_12515);
or U14674 (N_14674,N_12531,N_13428);
and U14675 (N_14675,N_13650,N_12654);
nor U14676 (N_14676,N_13511,N_13708);
nand U14677 (N_14677,N_12807,N_13590);
and U14678 (N_14678,N_13364,N_13318);
xor U14679 (N_14679,N_13462,N_13667);
nor U14680 (N_14680,N_12661,N_13714);
nand U14681 (N_14681,N_12893,N_12612);
xor U14682 (N_14682,N_13616,N_13390);
nand U14683 (N_14683,N_12610,N_12513);
nor U14684 (N_14684,N_13686,N_13513);
nand U14685 (N_14685,N_13181,N_12868);
nor U14686 (N_14686,N_13208,N_13020);
nand U14687 (N_14687,N_12666,N_13258);
nand U14688 (N_14688,N_13372,N_12974);
nor U14689 (N_14689,N_13661,N_13574);
nand U14690 (N_14690,N_13237,N_12685);
nand U14691 (N_14691,N_12738,N_13530);
nor U14692 (N_14692,N_12673,N_13116);
and U14693 (N_14693,N_13418,N_13170);
or U14694 (N_14694,N_13733,N_12749);
xor U14695 (N_14695,N_13742,N_12719);
xnor U14696 (N_14696,N_13172,N_12684);
or U14697 (N_14697,N_12575,N_12750);
nor U14698 (N_14698,N_12749,N_13498);
nor U14699 (N_14699,N_13270,N_13366);
xor U14700 (N_14700,N_13046,N_13201);
or U14701 (N_14701,N_13590,N_13460);
or U14702 (N_14702,N_12832,N_13191);
nand U14703 (N_14703,N_13529,N_12550);
xor U14704 (N_14704,N_13555,N_12619);
xnor U14705 (N_14705,N_13268,N_12625);
nor U14706 (N_14706,N_12788,N_13241);
and U14707 (N_14707,N_13469,N_13096);
xnor U14708 (N_14708,N_13389,N_12932);
and U14709 (N_14709,N_13637,N_13546);
nor U14710 (N_14710,N_13005,N_12574);
and U14711 (N_14711,N_13498,N_13278);
and U14712 (N_14712,N_12933,N_12733);
xor U14713 (N_14713,N_12650,N_13458);
nor U14714 (N_14714,N_13536,N_13331);
and U14715 (N_14715,N_13283,N_12955);
and U14716 (N_14716,N_13645,N_13173);
and U14717 (N_14717,N_13229,N_13147);
and U14718 (N_14718,N_13572,N_13614);
or U14719 (N_14719,N_13298,N_12953);
xor U14720 (N_14720,N_12521,N_12957);
xor U14721 (N_14721,N_12995,N_13469);
xor U14722 (N_14722,N_13683,N_13528);
nor U14723 (N_14723,N_12514,N_12903);
nand U14724 (N_14724,N_13738,N_13544);
and U14725 (N_14725,N_12640,N_13066);
or U14726 (N_14726,N_13675,N_13378);
nor U14727 (N_14727,N_13602,N_13328);
or U14728 (N_14728,N_12854,N_12747);
and U14729 (N_14729,N_13006,N_13379);
and U14730 (N_14730,N_12689,N_12667);
xor U14731 (N_14731,N_13511,N_13154);
or U14732 (N_14732,N_13678,N_13716);
nand U14733 (N_14733,N_13141,N_13675);
and U14734 (N_14734,N_12775,N_12966);
and U14735 (N_14735,N_13086,N_12523);
nor U14736 (N_14736,N_12814,N_12816);
nor U14737 (N_14737,N_12626,N_12905);
nor U14738 (N_14738,N_13688,N_13484);
nand U14739 (N_14739,N_12512,N_13275);
xnor U14740 (N_14740,N_12613,N_13270);
nand U14741 (N_14741,N_12929,N_13286);
or U14742 (N_14742,N_12823,N_12523);
xor U14743 (N_14743,N_12717,N_12810);
nand U14744 (N_14744,N_13513,N_12784);
or U14745 (N_14745,N_13244,N_13595);
and U14746 (N_14746,N_13496,N_12726);
xor U14747 (N_14747,N_13271,N_12709);
or U14748 (N_14748,N_13640,N_13688);
nor U14749 (N_14749,N_13507,N_12577);
xor U14750 (N_14750,N_13000,N_13712);
nand U14751 (N_14751,N_13241,N_13466);
or U14752 (N_14752,N_13552,N_12807);
or U14753 (N_14753,N_12562,N_12836);
nand U14754 (N_14754,N_13252,N_13601);
nand U14755 (N_14755,N_12798,N_12611);
nand U14756 (N_14756,N_13526,N_13006);
nand U14757 (N_14757,N_13394,N_13585);
or U14758 (N_14758,N_13532,N_12832);
nand U14759 (N_14759,N_12826,N_12593);
xnor U14760 (N_14760,N_12544,N_13542);
and U14761 (N_14761,N_12951,N_12743);
xor U14762 (N_14762,N_12977,N_13019);
nor U14763 (N_14763,N_13739,N_13622);
nand U14764 (N_14764,N_13144,N_12969);
xor U14765 (N_14765,N_12552,N_13098);
nand U14766 (N_14766,N_13044,N_13517);
nor U14767 (N_14767,N_13706,N_13679);
xor U14768 (N_14768,N_13090,N_13559);
and U14769 (N_14769,N_13125,N_13547);
nand U14770 (N_14770,N_13072,N_12891);
and U14771 (N_14771,N_13628,N_13040);
or U14772 (N_14772,N_12789,N_13269);
or U14773 (N_14773,N_12911,N_12552);
or U14774 (N_14774,N_13641,N_12791);
or U14775 (N_14775,N_13608,N_12570);
nor U14776 (N_14776,N_12584,N_12710);
nand U14777 (N_14777,N_12806,N_12742);
and U14778 (N_14778,N_12880,N_13471);
xor U14779 (N_14779,N_13313,N_13252);
xnor U14780 (N_14780,N_13672,N_12612);
or U14781 (N_14781,N_13155,N_13393);
and U14782 (N_14782,N_13277,N_12818);
or U14783 (N_14783,N_12617,N_12705);
xor U14784 (N_14784,N_13305,N_12683);
or U14785 (N_14785,N_12969,N_13556);
xnor U14786 (N_14786,N_13744,N_13109);
and U14787 (N_14787,N_12940,N_12904);
and U14788 (N_14788,N_13085,N_12884);
nor U14789 (N_14789,N_13170,N_13696);
nand U14790 (N_14790,N_13549,N_13344);
and U14791 (N_14791,N_13111,N_12923);
xor U14792 (N_14792,N_12945,N_12518);
or U14793 (N_14793,N_12908,N_13220);
nand U14794 (N_14794,N_13706,N_13217);
xnor U14795 (N_14795,N_13668,N_12830);
or U14796 (N_14796,N_13659,N_12581);
nand U14797 (N_14797,N_12526,N_13522);
and U14798 (N_14798,N_13104,N_12673);
nor U14799 (N_14799,N_12682,N_13708);
nor U14800 (N_14800,N_13281,N_12644);
nand U14801 (N_14801,N_12813,N_13690);
nand U14802 (N_14802,N_13492,N_13048);
nor U14803 (N_14803,N_13262,N_13346);
or U14804 (N_14804,N_12562,N_13117);
and U14805 (N_14805,N_12812,N_13138);
xor U14806 (N_14806,N_12839,N_13456);
and U14807 (N_14807,N_13160,N_13580);
nand U14808 (N_14808,N_13411,N_13328);
xnor U14809 (N_14809,N_13333,N_13311);
nand U14810 (N_14810,N_13583,N_13276);
xnor U14811 (N_14811,N_13456,N_13242);
and U14812 (N_14812,N_12777,N_12971);
or U14813 (N_14813,N_12752,N_12788);
xnor U14814 (N_14814,N_13028,N_12615);
nor U14815 (N_14815,N_13150,N_13449);
and U14816 (N_14816,N_13569,N_12852);
and U14817 (N_14817,N_12500,N_13636);
and U14818 (N_14818,N_13235,N_12969);
xnor U14819 (N_14819,N_13296,N_12657);
and U14820 (N_14820,N_12554,N_13221);
nor U14821 (N_14821,N_12972,N_13172);
nor U14822 (N_14822,N_12786,N_13724);
nand U14823 (N_14823,N_13154,N_13465);
xor U14824 (N_14824,N_13266,N_13462);
or U14825 (N_14825,N_13376,N_12774);
xor U14826 (N_14826,N_12508,N_12933);
or U14827 (N_14827,N_12610,N_13325);
nand U14828 (N_14828,N_12680,N_13289);
nand U14829 (N_14829,N_13676,N_13170);
or U14830 (N_14830,N_12789,N_12764);
xor U14831 (N_14831,N_13126,N_12752);
xor U14832 (N_14832,N_12548,N_13055);
nand U14833 (N_14833,N_13723,N_12554);
nor U14834 (N_14834,N_13661,N_12625);
or U14835 (N_14835,N_12514,N_12921);
nand U14836 (N_14836,N_13297,N_12846);
nor U14837 (N_14837,N_13061,N_13604);
and U14838 (N_14838,N_13317,N_13188);
or U14839 (N_14839,N_13709,N_12588);
nor U14840 (N_14840,N_12848,N_12664);
or U14841 (N_14841,N_13729,N_12973);
nor U14842 (N_14842,N_13240,N_13061);
nand U14843 (N_14843,N_13281,N_12787);
and U14844 (N_14844,N_12821,N_13579);
xnor U14845 (N_14845,N_12575,N_12698);
and U14846 (N_14846,N_13379,N_12861);
or U14847 (N_14847,N_13411,N_13585);
or U14848 (N_14848,N_13590,N_13276);
or U14849 (N_14849,N_12565,N_12843);
nand U14850 (N_14850,N_13648,N_12617);
and U14851 (N_14851,N_12809,N_13439);
and U14852 (N_14852,N_13339,N_12568);
and U14853 (N_14853,N_12553,N_12999);
and U14854 (N_14854,N_13688,N_13197);
nand U14855 (N_14855,N_13541,N_12749);
or U14856 (N_14856,N_13455,N_12739);
xnor U14857 (N_14857,N_13350,N_13563);
xnor U14858 (N_14858,N_13386,N_12782);
or U14859 (N_14859,N_12649,N_13221);
nand U14860 (N_14860,N_13224,N_13273);
and U14861 (N_14861,N_13140,N_12983);
and U14862 (N_14862,N_13442,N_12661);
nand U14863 (N_14863,N_13020,N_12652);
and U14864 (N_14864,N_13179,N_12831);
nor U14865 (N_14865,N_13642,N_12936);
nor U14866 (N_14866,N_12985,N_13492);
nand U14867 (N_14867,N_12757,N_13379);
and U14868 (N_14868,N_13311,N_13633);
nor U14869 (N_14869,N_12779,N_13538);
or U14870 (N_14870,N_12838,N_13353);
nand U14871 (N_14871,N_13408,N_13045);
nor U14872 (N_14872,N_13166,N_13572);
nor U14873 (N_14873,N_13304,N_13455);
and U14874 (N_14874,N_13234,N_12511);
nor U14875 (N_14875,N_13486,N_12866);
nor U14876 (N_14876,N_13008,N_13733);
nor U14877 (N_14877,N_12771,N_12587);
nand U14878 (N_14878,N_13487,N_13536);
nor U14879 (N_14879,N_13642,N_12982);
xor U14880 (N_14880,N_13624,N_13182);
xnor U14881 (N_14881,N_12512,N_12879);
nand U14882 (N_14882,N_13101,N_13333);
xor U14883 (N_14883,N_13585,N_13113);
or U14884 (N_14884,N_12530,N_13705);
and U14885 (N_14885,N_13546,N_13630);
xnor U14886 (N_14886,N_13530,N_12975);
nor U14887 (N_14887,N_12962,N_12700);
or U14888 (N_14888,N_13283,N_13342);
nand U14889 (N_14889,N_13051,N_12928);
nand U14890 (N_14890,N_13625,N_13440);
and U14891 (N_14891,N_12880,N_12554);
nand U14892 (N_14892,N_13315,N_13307);
xnor U14893 (N_14893,N_13642,N_12952);
nand U14894 (N_14894,N_12964,N_13203);
nand U14895 (N_14895,N_12963,N_13094);
nor U14896 (N_14896,N_13372,N_13267);
nand U14897 (N_14897,N_13187,N_13532);
or U14898 (N_14898,N_13665,N_12529);
and U14899 (N_14899,N_13035,N_13056);
xor U14900 (N_14900,N_13250,N_12775);
or U14901 (N_14901,N_12518,N_12869);
or U14902 (N_14902,N_12600,N_12930);
nor U14903 (N_14903,N_12895,N_12562);
and U14904 (N_14904,N_13455,N_12817);
nor U14905 (N_14905,N_12820,N_12617);
nor U14906 (N_14906,N_13079,N_13648);
xnor U14907 (N_14907,N_12600,N_13575);
and U14908 (N_14908,N_13426,N_13547);
xnor U14909 (N_14909,N_12966,N_12540);
and U14910 (N_14910,N_13123,N_12984);
nor U14911 (N_14911,N_12996,N_13439);
or U14912 (N_14912,N_13264,N_13602);
xnor U14913 (N_14913,N_12983,N_13320);
xor U14914 (N_14914,N_13182,N_12888);
nor U14915 (N_14915,N_13176,N_13231);
nand U14916 (N_14916,N_12532,N_13042);
xnor U14917 (N_14917,N_13563,N_12691);
xor U14918 (N_14918,N_12527,N_12602);
nand U14919 (N_14919,N_13247,N_12890);
and U14920 (N_14920,N_12548,N_13710);
and U14921 (N_14921,N_13234,N_13067);
xnor U14922 (N_14922,N_13560,N_13093);
xor U14923 (N_14923,N_12907,N_13363);
nor U14924 (N_14924,N_13398,N_12624);
xnor U14925 (N_14925,N_12629,N_13188);
or U14926 (N_14926,N_13539,N_13074);
nand U14927 (N_14927,N_13621,N_13313);
nor U14928 (N_14928,N_13427,N_12566);
nor U14929 (N_14929,N_13227,N_12909);
or U14930 (N_14930,N_13231,N_13354);
or U14931 (N_14931,N_12646,N_13500);
nand U14932 (N_14932,N_12608,N_12791);
nand U14933 (N_14933,N_12967,N_12658);
nor U14934 (N_14934,N_13680,N_12736);
or U14935 (N_14935,N_13004,N_13539);
or U14936 (N_14936,N_13460,N_12601);
or U14937 (N_14937,N_13652,N_12721);
or U14938 (N_14938,N_13415,N_13568);
and U14939 (N_14939,N_12956,N_13482);
xor U14940 (N_14940,N_13586,N_12632);
xor U14941 (N_14941,N_13188,N_13026);
and U14942 (N_14942,N_12676,N_12805);
and U14943 (N_14943,N_13696,N_13673);
xnor U14944 (N_14944,N_13462,N_13518);
nand U14945 (N_14945,N_13589,N_13087);
xnor U14946 (N_14946,N_13695,N_12555);
and U14947 (N_14947,N_13350,N_13476);
and U14948 (N_14948,N_13693,N_12852);
nor U14949 (N_14949,N_13617,N_13047);
or U14950 (N_14950,N_12740,N_13660);
xnor U14951 (N_14951,N_13261,N_13395);
nor U14952 (N_14952,N_13503,N_13574);
xnor U14953 (N_14953,N_13451,N_13492);
and U14954 (N_14954,N_13138,N_13597);
and U14955 (N_14955,N_13316,N_13030);
nand U14956 (N_14956,N_13106,N_12655);
or U14957 (N_14957,N_13556,N_13580);
or U14958 (N_14958,N_13200,N_12554);
and U14959 (N_14959,N_13065,N_13698);
nand U14960 (N_14960,N_12507,N_13398);
nor U14961 (N_14961,N_13665,N_12894);
and U14962 (N_14962,N_13236,N_13262);
nand U14963 (N_14963,N_13350,N_12987);
nand U14964 (N_14964,N_13507,N_13737);
xnor U14965 (N_14965,N_12653,N_13130);
nor U14966 (N_14966,N_13180,N_12887);
nand U14967 (N_14967,N_12651,N_13378);
and U14968 (N_14968,N_12972,N_12944);
xnor U14969 (N_14969,N_13341,N_13623);
nor U14970 (N_14970,N_13504,N_13665);
nor U14971 (N_14971,N_13307,N_13052);
or U14972 (N_14972,N_13135,N_13625);
or U14973 (N_14973,N_13593,N_12630);
or U14974 (N_14974,N_13140,N_13085);
or U14975 (N_14975,N_12550,N_13622);
nor U14976 (N_14976,N_13202,N_12873);
nand U14977 (N_14977,N_13523,N_13492);
nand U14978 (N_14978,N_13128,N_12652);
xor U14979 (N_14979,N_12588,N_13644);
and U14980 (N_14980,N_13313,N_12569);
nor U14981 (N_14981,N_13040,N_13467);
xor U14982 (N_14982,N_12679,N_12818);
nor U14983 (N_14983,N_13558,N_12561);
xnor U14984 (N_14984,N_12993,N_12732);
xor U14985 (N_14985,N_12652,N_13465);
and U14986 (N_14986,N_12967,N_12709);
nor U14987 (N_14987,N_13044,N_13413);
or U14988 (N_14988,N_13412,N_13717);
nor U14989 (N_14989,N_13588,N_13561);
and U14990 (N_14990,N_13710,N_13006);
and U14991 (N_14991,N_13520,N_12655);
nand U14992 (N_14992,N_12835,N_13136);
nand U14993 (N_14993,N_13537,N_13371);
nor U14994 (N_14994,N_13449,N_13154);
nor U14995 (N_14995,N_12605,N_12898);
nor U14996 (N_14996,N_12908,N_13274);
nand U14997 (N_14997,N_13713,N_12792);
nor U14998 (N_14998,N_12637,N_13611);
nor U14999 (N_14999,N_12841,N_13408);
xnor U15000 (N_15000,N_14919,N_14303);
or U15001 (N_15001,N_14687,N_14893);
or U15002 (N_15002,N_14573,N_14180);
nand U15003 (N_15003,N_14488,N_14165);
nor U15004 (N_15004,N_14663,N_14970);
and U15005 (N_15005,N_14873,N_14444);
or U15006 (N_15006,N_13768,N_14759);
nand U15007 (N_15007,N_14083,N_13853);
nor U15008 (N_15008,N_13979,N_13924);
or U15009 (N_15009,N_13995,N_14302);
and U15010 (N_15010,N_14194,N_14055);
xnor U15011 (N_15011,N_14361,N_14560);
nand U15012 (N_15012,N_14753,N_13892);
nand U15013 (N_15013,N_14876,N_13858);
or U15014 (N_15014,N_14046,N_14182);
and U15015 (N_15015,N_14716,N_13815);
and U15016 (N_15016,N_14157,N_14696);
xor U15017 (N_15017,N_13758,N_14599);
nand U15018 (N_15018,N_14930,N_13947);
nand U15019 (N_15019,N_14621,N_14153);
nor U15020 (N_15020,N_14534,N_14646);
xnor U15021 (N_15021,N_14918,N_13911);
nor U15022 (N_15022,N_14172,N_14031);
nor U15023 (N_15023,N_14975,N_13854);
nor U15024 (N_15024,N_14027,N_14672);
nor U15025 (N_15025,N_14339,N_13915);
or U15026 (N_15026,N_14337,N_14983);
and U15027 (N_15027,N_14911,N_14944);
xnor U15028 (N_15028,N_14197,N_14866);
xnor U15029 (N_15029,N_14790,N_14283);
xnor U15030 (N_15030,N_14788,N_14967);
xnor U15031 (N_15031,N_13786,N_14722);
xnor U15032 (N_15032,N_14270,N_14076);
xnor U15033 (N_15033,N_14735,N_14120);
nand U15034 (N_15034,N_14200,N_14282);
and U15035 (N_15035,N_14360,N_14224);
and U15036 (N_15036,N_14441,N_13863);
or U15037 (N_15037,N_14176,N_14518);
nor U15038 (N_15038,N_14563,N_14665);
and U15039 (N_15039,N_13798,N_13752);
and U15040 (N_15040,N_14269,N_14587);
xor U15041 (N_15041,N_14700,N_14523);
nand U15042 (N_15042,N_14150,N_13826);
xnor U15043 (N_15043,N_14832,N_14223);
and U15044 (N_15044,N_13937,N_14388);
xor U15045 (N_15045,N_14782,N_13806);
nand U15046 (N_15046,N_14236,N_13883);
nor U15047 (N_15047,N_14245,N_14152);
xor U15048 (N_15048,N_14792,N_14884);
nor U15049 (N_15049,N_14324,N_14660);
or U15050 (N_15050,N_13955,N_13970);
xnor U15051 (N_15051,N_13959,N_14809);
nor U15052 (N_15052,N_14814,N_14325);
xnor U15053 (N_15053,N_14341,N_14418);
or U15054 (N_15054,N_14010,N_14793);
or U15055 (N_15055,N_13941,N_14542);
and U15056 (N_15056,N_14928,N_14969);
xnor U15057 (N_15057,N_14304,N_14246);
or U15058 (N_15058,N_14773,N_13803);
xor U15059 (N_15059,N_14903,N_14477);
and U15060 (N_15060,N_14037,N_14216);
xor U15061 (N_15061,N_14936,N_14439);
xnor U15062 (N_15062,N_14065,N_14220);
xnor U15063 (N_15063,N_14358,N_14190);
or U15064 (N_15064,N_13813,N_14327);
or U15065 (N_15065,N_14988,N_14247);
nand U15066 (N_15066,N_14066,N_14907);
nand U15067 (N_15067,N_14993,N_14353);
and U15068 (N_15068,N_14750,N_14338);
and U15069 (N_15069,N_14511,N_14841);
nand U15070 (N_15070,N_14104,N_14167);
xnor U15071 (N_15071,N_14752,N_14734);
nor U15072 (N_15072,N_13865,N_13781);
nand U15073 (N_15073,N_14422,N_14342);
and U15074 (N_15074,N_14865,N_14105);
nor U15075 (N_15075,N_13868,N_14350);
nor U15076 (N_15076,N_14267,N_14968);
nor U15077 (N_15077,N_13958,N_14533);
xor U15078 (N_15078,N_14382,N_13994);
nand U15079 (N_15079,N_14473,N_13816);
nand U15080 (N_15080,N_13932,N_14710);
nor U15081 (N_15081,N_13841,N_14319);
nand U15082 (N_15082,N_13871,N_14440);
and U15083 (N_15083,N_14498,N_14854);
or U15084 (N_15084,N_14667,N_14503);
xnor U15085 (N_15085,N_14931,N_13774);
xnor U15086 (N_15086,N_14600,N_14254);
and U15087 (N_15087,N_14427,N_14080);
xnor U15088 (N_15088,N_14374,N_14438);
and U15089 (N_15089,N_14965,N_14668);
nor U15090 (N_15090,N_14308,N_14170);
or U15091 (N_15091,N_14138,N_13862);
xor U15092 (N_15092,N_14310,N_13800);
and U15093 (N_15093,N_13876,N_13890);
nand U15094 (N_15094,N_14399,N_14862);
nor U15095 (N_15095,N_14015,N_14326);
or U15096 (N_15096,N_14766,N_14530);
or U15097 (N_15097,N_13930,N_14289);
or U15098 (N_15098,N_14562,N_14078);
nor U15099 (N_15099,N_14297,N_14195);
or U15100 (N_15100,N_14491,N_14758);
nor U15101 (N_15101,N_14333,N_13791);
xor U15102 (N_15102,N_13807,N_14492);
xnor U15103 (N_15103,N_14974,N_14677);
nand U15104 (N_15104,N_13866,N_14739);
nand U15105 (N_15105,N_13808,N_14964);
nor U15106 (N_15106,N_14740,N_14410);
and U15107 (N_15107,N_13809,N_13850);
nor U15108 (N_15108,N_13952,N_13936);
nand U15109 (N_15109,N_14725,N_14014);
or U15110 (N_15110,N_14284,N_14049);
or U15111 (N_15111,N_14217,N_14939);
xor U15112 (N_15112,N_14203,N_14679);
and U15113 (N_15113,N_14485,N_14933);
and U15114 (N_15114,N_14372,N_13997);
xnor U15115 (N_15115,N_14652,N_14743);
and U15116 (N_15116,N_14068,N_14156);
nor U15117 (N_15117,N_13913,N_14777);
or U15118 (N_15118,N_14070,N_14584);
or U15119 (N_15119,N_14095,N_14100);
and U15120 (N_15120,N_14432,N_14532);
xor U15121 (N_15121,N_13895,N_14858);
xor U15122 (N_15122,N_14566,N_14047);
xnor U15123 (N_15123,N_14997,N_13904);
nand U15124 (N_15124,N_14359,N_13940);
nand U15125 (N_15125,N_14513,N_14411);
and U15126 (N_15126,N_14020,N_13977);
or U15127 (N_15127,N_14586,N_14092);
nand U15128 (N_15128,N_14248,N_14481);
nand U15129 (N_15129,N_14051,N_14611);
and U15130 (N_15130,N_14775,N_14574);
xor U15131 (N_15131,N_14746,N_14959);
nor U15132 (N_15132,N_14458,N_14373);
nand U15133 (N_15133,N_14464,N_14545);
and U15134 (N_15134,N_14762,N_14768);
xor U15135 (N_15135,N_14772,N_14553);
nor U15136 (N_15136,N_14756,N_14657);
nor U15137 (N_15137,N_13756,N_14312);
or U15138 (N_15138,N_14541,N_14886);
and U15139 (N_15139,N_14711,N_14629);
nor U15140 (N_15140,N_14384,N_14986);
nand U15141 (N_15141,N_14575,N_14380);
xnor U15142 (N_15142,N_14769,N_14749);
xnor U15143 (N_15143,N_13795,N_14883);
nand U15144 (N_15144,N_14653,N_14589);
nor U15145 (N_15145,N_13967,N_14641);
xor U15146 (N_15146,N_13948,N_14268);
and U15147 (N_15147,N_14213,N_14824);
xor U15148 (N_15148,N_14540,N_13822);
nand U15149 (N_15149,N_14158,N_14954);
nand U15150 (N_15150,N_14287,N_14826);
nor U15151 (N_15151,N_14771,N_14340);
or U15152 (N_15152,N_14362,N_13766);
or U15153 (N_15153,N_14510,N_14898);
or U15154 (N_15154,N_13907,N_14443);
or U15155 (N_15155,N_14785,N_14659);
and U15156 (N_15156,N_14184,N_14872);
or U15157 (N_15157,N_14789,N_14416);
nor U15158 (N_15158,N_14980,N_14596);
and U15159 (N_15159,N_13834,N_14757);
nor U15160 (N_15160,N_14597,N_14045);
or U15161 (N_15161,N_14215,N_14622);
and U15162 (N_15162,N_14979,N_14798);
xor U15163 (N_15163,N_13828,N_14693);
nor U15164 (N_15164,N_14730,N_13975);
nand U15165 (N_15165,N_14181,N_13893);
nand U15166 (N_15166,N_14487,N_14094);
or U15167 (N_15167,N_13987,N_14895);
or U15168 (N_15168,N_14126,N_13945);
nand U15169 (N_15169,N_14155,N_14009);
nand U15170 (N_15170,N_14494,N_14001);
and U15171 (N_15171,N_14407,N_14786);
nor U15172 (N_15172,N_14177,N_13917);
nor U15173 (N_15173,N_14259,N_14484);
nand U15174 (N_15174,N_14842,N_14332);
xor U15175 (N_15175,N_13825,N_14670);
and U15176 (N_15176,N_14859,N_13833);
and U15177 (N_15177,N_14817,N_14040);
xor U15178 (N_15178,N_13981,N_14064);
nand U15179 (N_15179,N_14313,N_14995);
or U15180 (N_15180,N_14957,N_14160);
and U15181 (N_15181,N_14744,N_13962);
nor U15182 (N_15182,N_14527,N_13903);
or U15183 (N_15183,N_14069,N_14921);
xnor U15184 (N_15184,N_14174,N_14524);
xnor U15185 (N_15185,N_14415,N_13933);
or U15186 (N_15186,N_14520,N_13976);
xnor U15187 (N_15187,N_14420,N_14594);
nand U15188 (N_15188,N_14937,N_14209);
nor U15189 (N_15189,N_14956,N_14683);
nor U15190 (N_15190,N_14007,N_14910);
and U15191 (N_15191,N_14550,N_14808);
xnor U15192 (N_15192,N_14378,N_14026);
or U15193 (N_15193,N_13971,N_13881);
and U15194 (N_15194,N_14222,N_14508);
and U15195 (N_15195,N_14229,N_13830);
nand U15196 (N_15196,N_13753,N_14807);
nand U15197 (N_15197,N_13773,N_14901);
nand U15198 (N_15198,N_14868,N_14273);
nand U15199 (N_15199,N_14475,N_14426);
or U15200 (N_15200,N_14990,N_14042);
nor U15201 (N_15201,N_14776,N_14462);
and U15202 (N_15202,N_14626,N_14602);
or U15203 (N_15203,N_13931,N_13760);
and U15204 (N_15204,N_14189,N_14011);
xor U15205 (N_15205,N_14419,N_14264);
nor U15206 (N_15206,N_14827,N_14914);
and U15207 (N_15207,N_14093,N_14457);
and U15208 (N_15208,N_14391,N_14175);
and U15209 (N_15209,N_14173,N_14201);
and U15210 (N_15210,N_14024,N_14115);
nand U15211 (N_15211,N_13943,N_13999);
or U15212 (N_15212,N_13942,N_14537);
nand U15213 (N_15213,N_14429,N_14811);
or U15214 (N_15214,N_14552,N_14783);
and U15215 (N_15215,N_14650,N_14465);
xor U15216 (N_15216,N_14234,N_14806);
and U15217 (N_15217,N_14228,N_14831);
nor U15218 (N_15218,N_13950,N_14179);
or U15219 (N_15219,N_14818,N_14674);
nor U15220 (N_15220,N_14241,N_14163);
xnor U15221 (N_15221,N_13873,N_14075);
xor U15222 (N_15222,N_14522,N_14941);
nor U15223 (N_15223,N_13867,N_14436);
or U15224 (N_15224,N_14315,N_13843);
or U15225 (N_15225,N_13934,N_14847);
nor U15226 (N_15226,N_13764,N_13842);
nand U15227 (N_15227,N_13778,N_13794);
or U15228 (N_15228,N_14676,N_14816);
nor U15229 (N_15229,N_14583,N_14991);
and U15230 (N_15230,N_14855,N_13784);
nor U15231 (N_15231,N_14005,N_14616);
xnor U15232 (N_15232,N_14635,N_14277);
or U15233 (N_15233,N_14747,N_13805);
nor U15234 (N_15234,N_14149,N_14891);
nor U15235 (N_15235,N_14061,N_14161);
or U15236 (N_15236,N_14030,N_14137);
nand U15237 (N_15237,N_14850,N_14888);
nor U15238 (N_15238,N_14673,N_14110);
xor U15239 (N_15239,N_14395,N_14091);
nor U15240 (N_15240,N_14951,N_14021);
nor U15241 (N_15241,N_14403,N_14043);
nor U15242 (N_15242,N_14882,N_14715);
xnor U15243 (N_15243,N_14344,N_14774);
and U15244 (N_15244,N_14396,N_14293);
or U15245 (N_15245,N_13921,N_14848);
xor U15246 (N_15246,N_14205,N_13991);
xor U15247 (N_15247,N_14751,N_14637);
nand U15248 (N_15248,N_14721,N_14474);
and U15249 (N_15249,N_14880,N_13851);
xor U15250 (N_15250,N_14028,N_13993);
and U15251 (N_15251,N_14431,N_13920);
or U15252 (N_15252,N_14881,N_13819);
nor U15253 (N_15253,N_13989,N_14169);
and U15254 (N_15254,N_14056,N_13922);
and U15255 (N_15255,N_14219,N_14546);
nor U15256 (N_15256,N_14675,N_14377);
xnor U15257 (N_15257,N_14837,N_14764);
or U15258 (N_15258,N_14334,N_14192);
and U15259 (N_15259,N_14301,N_13780);
and U15260 (N_15260,N_14390,N_14828);
or U15261 (N_15261,N_14942,N_14112);
xnor U15262 (N_15262,N_14425,N_14250);
and U15263 (N_15263,N_13923,N_14606);
nand U15264 (N_15264,N_14002,N_14478);
and U15265 (N_15265,N_14517,N_13886);
xor U15266 (N_15266,N_14035,N_14823);
or U15267 (N_15267,N_13817,N_14820);
or U15268 (N_15268,N_14370,N_14736);
nand U15269 (N_15269,N_14551,N_14143);
nor U15270 (N_15270,N_14453,N_14086);
nand U15271 (N_15271,N_13787,N_14193);
nor U15272 (N_15272,N_13877,N_14879);
nand U15273 (N_15273,N_13887,N_14840);
or U15274 (N_15274,N_13832,N_14320);
xnor U15275 (N_15275,N_14952,N_14707);
nand U15276 (N_15276,N_14932,N_14732);
nor U15277 (N_15277,N_14973,N_14405);
or U15278 (N_15278,N_14631,N_14927);
xor U15279 (N_15279,N_14019,N_14681);
nand U15280 (N_15280,N_14796,N_13884);
and U15281 (N_15281,N_14733,N_14651);
nand U15282 (N_15282,N_14398,N_14349);
and U15283 (N_15283,N_13779,N_14875);
xor U15284 (N_15284,N_14829,N_14121);
and U15285 (N_15285,N_14452,N_14394);
nand U15286 (N_15286,N_14463,N_14794);
xnor U15287 (N_15287,N_14408,N_13935);
or U15288 (N_15288,N_14502,N_13972);
xnor U15289 (N_15289,N_13852,N_14328);
nor U15290 (N_15290,N_14648,N_13944);
nand U15291 (N_15291,N_14098,N_13896);
nand U15292 (N_15292,N_14843,N_14012);
xor U15293 (N_15293,N_14500,N_14274);
or U15294 (N_15294,N_14692,N_13759);
and U15295 (N_15295,N_14509,N_14953);
nand U15296 (N_15296,N_14628,N_14255);
or U15297 (N_15297,N_14085,N_14008);
xor U15298 (N_15298,N_14423,N_14833);
nor U15299 (N_15299,N_14188,N_14935);
nand U15300 (N_15300,N_14421,N_14591);
nor U15301 (N_15301,N_14572,N_14168);
nand U15302 (N_15302,N_13831,N_14581);
nor U15303 (N_15303,N_14800,N_14140);
or U15304 (N_15304,N_14669,N_14978);
nand U15305 (N_15305,N_14963,N_14977);
nor U15306 (N_15306,N_14543,N_14428);
and U15307 (N_15307,N_14922,N_14625);
and U15308 (N_15308,N_14052,N_13870);
nand U15309 (N_15309,N_13909,N_14501);
nand U15310 (N_15310,N_14642,N_14242);
or U15311 (N_15311,N_14240,N_13790);
nor U15312 (N_15312,N_14556,N_14263);
xor U15313 (N_15313,N_14210,N_14356);
nand U15314 (N_15314,N_14731,N_14369);
or U15315 (N_15315,N_14719,N_14206);
and U15316 (N_15316,N_14900,N_14630);
nand U15317 (N_15317,N_14036,N_14761);
nor U15318 (N_15318,N_14430,N_14839);
or U15319 (N_15319,N_14044,N_14728);
and U15320 (N_15320,N_14982,N_14726);
nand U15321 (N_15321,N_14489,N_13783);
xor U15322 (N_15322,N_13998,N_14393);
or U15323 (N_15323,N_13772,N_14643);
or U15324 (N_15324,N_14280,N_14934);
nor U15325 (N_15325,N_14013,N_14185);
nor U15326 (N_15326,N_14299,N_14887);
xor U15327 (N_15327,N_14835,N_14318);
nor U15328 (N_15328,N_14519,N_14878);
nor U15329 (N_15329,N_13754,N_14039);
nand U15330 (N_15330,N_14476,N_14097);
nor U15331 (N_15331,N_14703,N_14166);
xor U15332 (N_15332,N_13906,N_13776);
or U15333 (N_15333,N_13844,N_13793);
and U15334 (N_15334,N_13878,N_14468);
nor U15335 (N_15335,N_13872,N_14226);
or U15336 (N_15336,N_14614,N_14557);
nor U15337 (N_15337,N_14874,N_14142);
nand U15338 (N_15338,N_14528,N_14196);
and U15339 (N_15339,N_14135,N_14763);
or U15340 (N_15340,N_14955,N_14208);
or U15341 (N_15341,N_14576,N_14985);
and U15342 (N_15342,N_13782,N_14992);
and U15343 (N_15343,N_14819,N_14507);
nand U15344 (N_15344,N_13902,N_14691);
or U15345 (N_15345,N_14400,N_14999);
and U15346 (N_15346,N_14128,N_14971);
and U15347 (N_15347,N_14605,N_14564);
nand U15348 (N_15348,N_14547,N_14445);
nand U15349 (N_15349,N_14544,N_13848);
nor U15350 (N_15350,N_14003,N_14081);
xnor U15351 (N_15351,N_14860,N_14760);
or U15352 (N_15352,N_14561,N_14480);
and U15353 (N_15353,N_14905,N_13847);
xnor U15354 (N_15354,N_14699,N_14376);
and U15355 (N_15355,N_14368,N_14727);
xnor U15356 (N_15356,N_14632,N_14434);
xor U15357 (N_15357,N_14336,N_14885);
nand U15358 (N_15358,N_13812,N_14579);
and U15359 (N_15359,N_14946,N_14278);
or U15360 (N_15360,N_14469,N_14330);
xnor U15361 (N_15361,N_14912,N_14697);
or U15362 (N_15362,N_13855,N_14615);
xor U15363 (N_15363,N_14825,N_14577);
nor U15364 (N_15364,N_14450,N_14059);
xor U15365 (N_15365,N_14067,N_13891);
nand U15366 (N_15366,N_14702,N_14588);
nor U15367 (N_15367,N_14689,N_14034);
and U15368 (N_15368,N_14805,N_14183);
xor U15369 (N_15369,N_14943,N_14144);
nand U15370 (N_15370,N_14821,N_14290);
and U15371 (N_15371,N_13810,N_14791);
xnor U15372 (N_15372,N_13767,N_13889);
xor U15373 (N_15373,N_14146,N_14371);
or U15374 (N_15374,N_13785,N_14765);
or U15375 (N_15375,N_14448,N_14386);
and U15376 (N_15376,N_14096,N_14926);
or U15377 (N_15377,N_13755,N_14506);
nand U15378 (N_15378,N_14984,N_14131);
or U15379 (N_15379,N_13980,N_14025);
nor U15380 (N_15380,N_14253,N_14671);
nor U15381 (N_15381,N_14364,N_14662);
or U15382 (N_15382,N_14109,N_14238);
or U15383 (N_15383,N_13927,N_14352);
nor U15384 (N_15384,N_14249,N_14383);
nand U15385 (N_15385,N_14317,N_13879);
or U15386 (N_15386,N_14038,N_14365);
nor U15387 (N_15387,N_13880,N_14565);
or U15388 (N_15388,N_14295,N_14237);
nand U15389 (N_15389,N_14244,N_14869);
nand U15390 (N_15390,N_14033,N_14276);
nand U15391 (N_15391,N_14770,N_14938);
nand U15392 (N_15392,N_13956,N_14559);
xnor U15393 (N_15393,N_14851,N_14111);
or U15394 (N_15394,N_14617,N_14863);
nor U15395 (N_15395,N_14685,N_14191);
or U15396 (N_15396,N_14472,N_14998);
and U15397 (N_15397,N_14389,N_13859);
or U15398 (N_15398,N_14275,N_14114);
and U15399 (N_15399,N_13861,N_14134);
or U15400 (N_15400,N_14207,N_14571);
xnor U15401 (N_15401,N_14531,N_14417);
nand U15402 (N_15402,N_14694,N_14505);
or U15403 (N_15403,N_13961,N_14397);
or U15404 (N_15404,N_13856,N_14235);
nand U15405 (N_15405,N_14610,N_14392);
xnor U15406 (N_15406,N_13954,N_14698);
or U15407 (N_15407,N_14845,N_14723);
nor U15408 (N_15408,N_14218,N_14767);
or U15409 (N_15409,N_14256,N_14154);
xor U15410 (N_15410,N_14950,N_14345);
nor U15411 (N_15411,N_14619,N_14424);
or U15412 (N_15412,N_14032,N_13761);
xor U15413 (N_15413,N_14057,N_14225);
xor U15414 (N_15414,N_14082,N_14958);
or U15415 (N_15415,N_14016,N_14381);
nor U15416 (N_15416,N_14446,N_14291);
or U15417 (N_15417,N_14567,N_14962);
nor U15418 (N_15418,N_14198,N_14529);
or U15419 (N_15419,N_14655,N_14754);
nor U15420 (N_15420,N_14199,N_13824);
and U15421 (N_15421,N_14456,N_14890);
nor U15422 (N_15422,N_14343,N_14041);
xnor U15423 (N_15423,N_14871,N_14633);
nand U15424 (N_15424,N_14569,N_14412);
nor U15425 (N_15425,N_14585,N_14311);
xor U15426 (N_15426,N_14535,N_14089);
xor U15427 (N_15427,N_14961,N_14601);
or U15428 (N_15428,N_14106,N_14678);
xor U15429 (N_15429,N_13839,N_14145);
xor U15430 (N_15430,N_14300,N_14164);
xor U15431 (N_15431,N_14706,N_14316);
and U15432 (N_15432,N_14062,N_14558);
nand U15433 (N_15433,N_14894,N_13835);
nand U15434 (N_15434,N_14271,N_13928);
xor U15435 (N_15435,N_14515,N_14258);
or U15436 (N_15436,N_13983,N_14306);
or U15437 (N_15437,N_14401,N_14211);
nor U15438 (N_15438,N_14366,N_14251);
or U15439 (N_15439,N_14495,N_14022);
and U15440 (N_15440,N_14296,N_13978);
xnor U15441 (N_15441,N_14261,N_14549);
or U15442 (N_15442,N_13910,N_14202);
nand U15443 (N_15443,N_14636,N_14108);
and U15444 (N_15444,N_14603,N_14402);
xor U15445 (N_15445,N_14741,N_14779);
xnor U15446 (N_15446,N_13919,N_14604);
nor U15447 (N_15447,N_14947,N_13882);
xnor U15448 (N_15448,N_14525,N_14063);
nor U15449 (N_15449,N_14634,N_13804);
or U15450 (N_15450,N_14000,N_14496);
or U15451 (N_15451,N_14795,N_13899);
xor U15452 (N_15452,N_14802,N_13951);
or U15453 (N_15453,N_13914,N_14504);
nand U15454 (N_15454,N_14088,N_14889);
nand U15455 (N_15455,N_14355,N_14654);
nand U15456 (N_15456,N_13762,N_14084);
or U15457 (N_15457,N_13926,N_13765);
or U15458 (N_15458,N_14272,N_14781);
nor U15459 (N_15459,N_14688,N_14467);
and U15460 (N_15460,N_14351,N_14486);
nor U15461 (N_15461,N_13957,N_14708);
and U15462 (N_15462,N_14923,N_14624);
or U15463 (N_15463,N_14784,N_14347);
nand U15464 (N_15464,N_14618,N_14288);
xor U15465 (N_15465,N_13823,N_14292);
nand U15466 (N_15466,N_13946,N_14053);
xnor U15467 (N_15467,N_13849,N_14680);
or U15468 (N_15468,N_14666,N_14892);
xor U15469 (N_15469,N_14058,N_14623);
or U15470 (N_15470,N_14686,N_14231);
xnor U15471 (N_15471,N_14279,N_14592);
nand U15472 (N_15472,N_13771,N_14018);
and U15473 (N_15473,N_13864,N_14813);
or U15474 (N_15474,N_14107,N_14227);
xor U15475 (N_15475,N_14864,N_14897);
or U15476 (N_15476,N_14171,N_14870);
nand U15477 (N_15477,N_14593,N_14664);
or U15478 (N_15478,N_14849,N_13964);
or U15479 (N_15479,N_14929,N_14704);
nor U15480 (N_15480,N_14357,N_14204);
and U15481 (N_15481,N_13905,N_13960);
nor U15482 (N_15482,N_14090,N_14981);
xor U15483 (N_15483,N_13949,N_13845);
or U15484 (N_15484,N_14125,N_14645);
nor U15485 (N_15485,N_14101,N_14470);
and U15486 (N_15486,N_13929,N_14479);
xnor U15487 (N_15487,N_14915,N_14598);
xor U15488 (N_15488,N_14987,N_14538);
nor U15489 (N_15489,N_14582,N_14127);
nor U15490 (N_15490,N_14714,N_14379);
xor U15491 (N_15491,N_14178,N_14133);
nand U15492 (N_15492,N_13965,N_14239);
nand U15493 (N_15493,N_14830,N_13770);
nor U15494 (N_15494,N_14004,N_14077);
nor U15495 (N_15495,N_14252,N_14804);
and U15496 (N_15496,N_13818,N_14354);
nor U15497 (N_15497,N_14904,N_14834);
xnor U15498 (N_15498,N_14314,N_14815);
xnor U15499 (N_15499,N_13763,N_13811);
nor U15500 (N_15500,N_14755,N_14130);
xor U15501 (N_15501,N_14265,N_14442);
and U15502 (N_15502,N_14713,N_14989);
nor U15503 (N_15503,N_14822,N_14006);
or U15504 (N_15504,N_13837,N_13938);
nand U15505 (N_15505,N_14404,N_14136);
nand U15506 (N_15506,N_14590,N_14490);
or U15507 (N_15507,N_14724,N_14335);
xor U15508 (N_15508,N_14972,N_14409);
nor U15509 (N_15509,N_14709,N_14305);
nand U15510 (N_15510,N_14132,N_14701);
xor U15511 (N_15511,N_14079,N_14966);
or U15512 (N_15512,N_13984,N_14899);
xor U15513 (N_15513,N_14612,N_14838);
xor U15514 (N_15514,N_14148,N_13829);
and U15515 (N_15515,N_14151,N_14712);
nand U15516 (N_15516,N_14738,N_13869);
nand U15517 (N_15517,N_14578,N_14029);
xor U15518 (N_15518,N_13969,N_14413);
or U15519 (N_15519,N_14960,N_14499);
nor U15520 (N_15520,N_13796,N_14745);
nand U15521 (N_15521,N_13894,N_14129);
or U15522 (N_15522,N_14639,N_14186);
or U15523 (N_15523,N_14017,N_14187);
or U15524 (N_15524,N_14690,N_14742);
and U15525 (N_15525,N_14638,N_14620);
xnor U15526 (N_15526,N_14945,N_13966);
nor U15527 (N_15527,N_14920,N_14117);
and U15528 (N_15528,N_14801,N_14925);
nor U15529 (N_15529,N_14799,N_14387);
or U15530 (N_15530,N_14141,N_14122);
nor U15531 (N_15531,N_14048,N_13992);
nand U15532 (N_15532,N_13990,N_13982);
xor U15533 (N_15533,N_14414,N_14516);
nor U15534 (N_15534,N_13838,N_14159);
xor U15535 (N_15535,N_14656,N_14023);
nand U15536 (N_15536,N_14260,N_14346);
nand U15537 (N_15537,N_13918,N_14536);
nand U15538 (N_15538,N_14072,N_13901);
and U15539 (N_15539,N_13789,N_14406);
and U15540 (N_15540,N_13827,N_14321);
or U15541 (N_15541,N_14644,N_14717);
xor U15542 (N_15542,N_14294,N_14459);
or U15543 (N_15543,N_14695,N_14323);
nand U15544 (N_15544,N_13857,N_13985);
and U15545 (N_15545,N_14113,N_14329);
and U15546 (N_15546,N_14435,N_14471);
and U15547 (N_15547,N_14307,N_14778);
nor U15548 (N_15548,N_14949,N_14118);
nand U15549 (N_15549,N_14810,N_13757);
and U15550 (N_15550,N_13860,N_14385);
and U15551 (N_15551,N_14257,N_14857);
and U15552 (N_15552,N_14521,N_13769);
nand U15553 (N_15553,N_14483,N_14896);
xor U15554 (N_15554,N_14526,N_14787);
or U15555 (N_15555,N_14924,N_13797);
and U15556 (N_15556,N_13751,N_14482);
nand U15557 (N_15557,N_14948,N_13912);
xor U15558 (N_15558,N_14568,N_14071);
nor U15559 (N_15559,N_14322,N_13788);
nand U15560 (N_15560,N_14996,N_14803);
or U15561 (N_15561,N_14367,N_14627);
or U15562 (N_15562,N_14454,N_14917);
or U15563 (N_15563,N_13925,N_14497);
and U15564 (N_15564,N_13750,N_13820);
xor U15565 (N_15565,N_14461,N_14050);
nor U15566 (N_15566,N_14433,N_14856);
and U15567 (N_15567,N_14909,N_14437);
xnor U15568 (N_15568,N_14451,N_14607);
and U15569 (N_15569,N_14060,N_14608);
nor U15570 (N_15570,N_13840,N_13939);
or U15571 (N_15571,N_14580,N_14554);
and U15572 (N_15572,N_13996,N_14514);
and U15573 (N_15573,N_13821,N_14214);
and U15574 (N_15574,N_14262,N_14281);
nand U15575 (N_15575,N_14449,N_13874);
xnor U15576 (N_15576,N_14073,N_13973);
nand U15577 (N_15577,N_13777,N_14363);
xor U15578 (N_15578,N_14298,N_14555);
nand U15579 (N_15579,N_14729,N_14913);
xor U15580 (N_15580,N_14877,N_14139);
or U15581 (N_15581,N_14102,N_13836);
or U15582 (N_15582,N_14908,N_13888);
xor U15583 (N_15583,N_13885,N_14852);
xnor U15584 (N_15584,N_14493,N_14867);
xor U15585 (N_15585,N_13953,N_13968);
nand U15586 (N_15586,N_14812,N_14647);
xnor U15587 (N_15587,N_14902,N_13963);
nand U15588 (N_15588,N_14844,N_14548);
xnor U15589 (N_15589,N_14976,N_13974);
xnor U15590 (N_15590,N_14613,N_14661);
xnor U15591 (N_15591,N_14348,N_13916);
or U15592 (N_15592,N_14116,N_13900);
xnor U15593 (N_15593,N_13986,N_14658);
xnor U15594 (N_15594,N_14853,N_14162);
or U15595 (N_15595,N_14230,N_14595);
or U15596 (N_15596,N_13801,N_14705);
or U15597 (N_15597,N_14286,N_13799);
nand U15598 (N_15598,N_14266,N_14221);
or U15599 (N_15599,N_13802,N_14861);
nand U15600 (N_15600,N_14054,N_14649);
xor U15601 (N_15601,N_14570,N_13814);
xor U15602 (N_15602,N_14718,N_14748);
xor U15603 (N_15603,N_13792,N_14124);
nor U15604 (N_15604,N_14940,N_14684);
nand U15605 (N_15605,N_14147,N_14460);
xnor U15606 (N_15606,N_14285,N_14375);
nand U15607 (N_15607,N_13898,N_14609);
nor U15608 (N_15608,N_14780,N_14309);
or U15609 (N_15609,N_14103,N_13897);
nor U15610 (N_15610,N_13846,N_14119);
and U15611 (N_15611,N_13875,N_14466);
and U15612 (N_15612,N_14906,N_14243);
xnor U15613 (N_15613,N_14640,N_13775);
and U15614 (N_15614,N_14682,N_13988);
and U15615 (N_15615,N_14212,N_14512);
nand U15616 (N_15616,N_14331,N_14994);
nand U15617 (N_15617,N_14539,N_14123);
and U15618 (N_15618,N_14233,N_14099);
xor U15619 (N_15619,N_14232,N_14846);
nor U15620 (N_15620,N_14737,N_14836);
xnor U15621 (N_15621,N_14074,N_14087);
and U15622 (N_15622,N_14916,N_14720);
nor U15623 (N_15623,N_14797,N_13908);
or U15624 (N_15624,N_14455,N_14447);
nand U15625 (N_15625,N_14476,N_14191);
nand U15626 (N_15626,N_14962,N_14138);
nand U15627 (N_15627,N_14102,N_14097);
or U15628 (N_15628,N_14341,N_14631);
and U15629 (N_15629,N_14136,N_14002);
or U15630 (N_15630,N_13846,N_14755);
xor U15631 (N_15631,N_14685,N_14892);
nand U15632 (N_15632,N_14141,N_14805);
or U15633 (N_15633,N_14826,N_14092);
nor U15634 (N_15634,N_13961,N_14075);
nand U15635 (N_15635,N_13862,N_14260);
nor U15636 (N_15636,N_13850,N_14796);
nor U15637 (N_15637,N_14338,N_14749);
nor U15638 (N_15638,N_14222,N_14533);
nand U15639 (N_15639,N_13760,N_14324);
xor U15640 (N_15640,N_14721,N_14197);
nand U15641 (N_15641,N_14740,N_13917);
xnor U15642 (N_15642,N_14924,N_13957);
nor U15643 (N_15643,N_13785,N_14456);
and U15644 (N_15644,N_13900,N_13835);
nor U15645 (N_15645,N_14283,N_14758);
or U15646 (N_15646,N_14509,N_14379);
nor U15647 (N_15647,N_13760,N_14232);
nor U15648 (N_15648,N_14637,N_14974);
or U15649 (N_15649,N_14048,N_14424);
nor U15650 (N_15650,N_14158,N_14459);
xor U15651 (N_15651,N_14385,N_14693);
or U15652 (N_15652,N_14180,N_14453);
nand U15653 (N_15653,N_14728,N_13884);
xnor U15654 (N_15654,N_14251,N_13977);
or U15655 (N_15655,N_14632,N_14014);
nand U15656 (N_15656,N_13824,N_14573);
and U15657 (N_15657,N_14935,N_14418);
nand U15658 (N_15658,N_14619,N_14538);
nand U15659 (N_15659,N_14826,N_14533);
nand U15660 (N_15660,N_14279,N_14071);
or U15661 (N_15661,N_13856,N_14657);
nand U15662 (N_15662,N_14455,N_13801);
and U15663 (N_15663,N_13791,N_14133);
nor U15664 (N_15664,N_14572,N_14713);
nand U15665 (N_15665,N_14555,N_14362);
nor U15666 (N_15666,N_14215,N_14898);
or U15667 (N_15667,N_13893,N_13922);
and U15668 (N_15668,N_14332,N_14878);
nand U15669 (N_15669,N_14888,N_13912);
xor U15670 (N_15670,N_14343,N_14085);
xnor U15671 (N_15671,N_13864,N_13790);
and U15672 (N_15672,N_14339,N_14666);
or U15673 (N_15673,N_13860,N_14093);
xnor U15674 (N_15674,N_14914,N_14394);
nand U15675 (N_15675,N_14873,N_14870);
and U15676 (N_15676,N_14921,N_14007);
nor U15677 (N_15677,N_14316,N_14772);
or U15678 (N_15678,N_14326,N_14888);
nor U15679 (N_15679,N_14858,N_13978);
nand U15680 (N_15680,N_13920,N_13752);
and U15681 (N_15681,N_14274,N_13979);
nor U15682 (N_15682,N_13888,N_14090);
and U15683 (N_15683,N_14056,N_14670);
and U15684 (N_15684,N_14952,N_14488);
and U15685 (N_15685,N_14865,N_13962);
nor U15686 (N_15686,N_14158,N_14982);
nand U15687 (N_15687,N_14648,N_13953);
or U15688 (N_15688,N_14490,N_14156);
and U15689 (N_15689,N_14891,N_14474);
nand U15690 (N_15690,N_14342,N_13957);
and U15691 (N_15691,N_14803,N_14942);
nand U15692 (N_15692,N_14386,N_13980);
and U15693 (N_15693,N_14884,N_13894);
or U15694 (N_15694,N_14912,N_14062);
nand U15695 (N_15695,N_14753,N_14181);
and U15696 (N_15696,N_14209,N_14250);
nand U15697 (N_15697,N_14003,N_14858);
nand U15698 (N_15698,N_13774,N_13777);
nor U15699 (N_15699,N_13781,N_14363);
nor U15700 (N_15700,N_14363,N_13788);
nor U15701 (N_15701,N_14641,N_13883);
and U15702 (N_15702,N_14432,N_14875);
and U15703 (N_15703,N_13898,N_14445);
and U15704 (N_15704,N_14818,N_14080);
nor U15705 (N_15705,N_14522,N_14432);
and U15706 (N_15706,N_13918,N_14767);
xor U15707 (N_15707,N_14488,N_13935);
xor U15708 (N_15708,N_14974,N_14115);
and U15709 (N_15709,N_14310,N_13937);
and U15710 (N_15710,N_14526,N_14850);
nor U15711 (N_15711,N_14407,N_14094);
xor U15712 (N_15712,N_14942,N_13775);
or U15713 (N_15713,N_14365,N_14345);
or U15714 (N_15714,N_14627,N_14156);
nor U15715 (N_15715,N_14055,N_14927);
nor U15716 (N_15716,N_13869,N_14518);
or U15717 (N_15717,N_14672,N_14679);
nand U15718 (N_15718,N_14455,N_14637);
nor U15719 (N_15719,N_14337,N_14104);
xor U15720 (N_15720,N_14817,N_14182);
xnor U15721 (N_15721,N_14870,N_14578);
or U15722 (N_15722,N_14013,N_14573);
and U15723 (N_15723,N_14326,N_13934);
nand U15724 (N_15724,N_14073,N_14179);
or U15725 (N_15725,N_14729,N_14659);
nor U15726 (N_15726,N_14425,N_13853);
or U15727 (N_15727,N_14818,N_13985);
and U15728 (N_15728,N_14636,N_14671);
and U15729 (N_15729,N_13798,N_14640);
nand U15730 (N_15730,N_14302,N_14993);
nand U15731 (N_15731,N_13790,N_14150);
or U15732 (N_15732,N_13757,N_14431);
nand U15733 (N_15733,N_14667,N_14387);
nor U15734 (N_15734,N_14124,N_14881);
nand U15735 (N_15735,N_14232,N_14549);
xnor U15736 (N_15736,N_14050,N_14296);
nor U15737 (N_15737,N_14115,N_13955);
or U15738 (N_15738,N_14981,N_14385);
nor U15739 (N_15739,N_14378,N_14959);
nor U15740 (N_15740,N_13841,N_14560);
or U15741 (N_15741,N_14309,N_14592);
nor U15742 (N_15742,N_14262,N_14428);
or U15743 (N_15743,N_14794,N_13849);
nand U15744 (N_15744,N_13919,N_14464);
and U15745 (N_15745,N_14926,N_14288);
or U15746 (N_15746,N_14345,N_14861);
xnor U15747 (N_15747,N_14224,N_14039);
or U15748 (N_15748,N_14008,N_14391);
or U15749 (N_15749,N_14139,N_14769);
nand U15750 (N_15750,N_14100,N_14669);
nand U15751 (N_15751,N_13828,N_14744);
xnor U15752 (N_15752,N_13937,N_14781);
and U15753 (N_15753,N_14962,N_14383);
and U15754 (N_15754,N_14087,N_14940);
and U15755 (N_15755,N_14045,N_13882);
nand U15756 (N_15756,N_14016,N_14416);
or U15757 (N_15757,N_13911,N_14679);
or U15758 (N_15758,N_14476,N_13863);
and U15759 (N_15759,N_13860,N_14801);
or U15760 (N_15760,N_14664,N_14553);
or U15761 (N_15761,N_14380,N_14825);
and U15762 (N_15762,N_14515,N_14519);
xor U15763 (N_15763,N_14067,N_14925);
or U15764 (N_15764,N_14848,N_14533);
nor U15765 (N_15765,N_14737,N_13831);
or U15766 (N_15766,N_13827,N_14915);
xnor U15767 (N_15767,N_14140,N_14497);
nand U15768 (N_15768,N_14773,N_14953);
nor U15769 (N_15769,N_14537,N_14861);
xnor U15770 (N_15770,N_13897,N_14371);
or U15771 (N_15771,N_14044,N_14525);
nor U15772 (N_15772,N_14541,N_14325);
nor U15773 (N_15773,N_14148,N_13965);
nand U15774 (N_15774,N_14780,N_14332);
and U15775 (N_15775,N_14301,N_14924);
or U15776 (N_15776,N_14930,N_14248);
and U15777 (N_15777,N_14195,N_14134);
nand U15778 (N_15778,N_13865,N_13878);
xor U15779 (N_15779,N_13883,N_13855);
and U15780 (N_15780,N_13821,N_14578);
xnor U15781 (N_15781,N_14797,N_14731);
or U15782 (N_15782,N_13869,N_13876);
or U15783 (N_15783,N_14494,N_14086);
xor U15784 (N_15784,N_14064,N_14826);
xor U15785 (N_15785,N_14535,N_13906);
xnor U15786 (N_15786,N_13988,N_14867);
nand U15787 (N_15787,N_13946,N_14382);
xor U15788 (N_15788,N_14778,N_14446);
nand U15789 (N_15789,N_14287,N_14032);
or U15790 (N_15790,N_13887,N_14889);
nor U15791 (N_15791,N_14814,N_14954);
xor U15792 (N_15792,N_14088,N_14671);
nor U15793 (N_15793,N_14529,N_14009);
nor U15794 (N_15794,N_14236,N_14258);
nor U15795 (N_15795,N_14654,N_14012);
xor U15796 (N_15796,N_13933,N_14402);
nor U15797 (N_15797,N_14819,N_14535);
nor U15798 (N_15798,N_14795,N_14251);
and U15799 (N_15799,N_14137,N_14284);
xor U15800 (N_15800,N_14480,N_14812);
nand U15801 (N_15801,N_13893,N_14994);
or U15802 (N_15802,N_14725,N_14391);
or U15803 (N_15803,N_14921,N_14408);
nor U15804 (N_15804,N_14874,N_14435);
xor U15805 (N_15805,N_14224,N_14716);
nor U15806 (N_15806,N_13805,N_14944);
nand U15807 (N_15807,N_14991,N_14154);
nand U15808 (N_15808,N_13918,N_14046);
xor U15809 (N_15809,N_13820,N_14410);
nor U15810 (N_15810,N_14957,N_14600);
nand U15811 (N_15811,N_14753,N_14370);
nor U15812 (N_15812,N_14708,N_14523);
xor U15813 (N_15813,N_14029,N_14181);
and U15814 (N_15814,N_14297,N_14012);
nand U15815 (N_15815,N_13809,N_14282);
nand U15816 (N_15816,N_13874,N_14996);
xor U15817 (N_15817,N_13815,N_14951);
and U15818 (N_15818,N_13828,N_14899);
nor U15819 (N_15819,N_14779,N_14213);
or U15820 (N_15820,N_13771,N_14271);
and U15821 (N_15821,N_14258,N_13752);
nand U15822 (N_15822,N_13950,N_13853);
nor U15823 (N_15823,N_14331,N_14323);
or U15824 (N_15824,N_14176,N_14099);
or U15825 (N_15825,N_14116,N_14724);
nor U15826 (N_15826,N_13887,N_14298);
or U15827 (N_15827,N_14282,N_14956);
nor U15828 (N_15828,N_14056,N_14148);
or U15829 (N_15829,N_14619,N_14593);
xnor U15830 (N_15830,N_14490,N_14811);
nand U15831 (N_15831,N_14525,N_13810);
xnor U15832 (N_15832,N_14667,N_14289);
and U15833 (N_15833,N_13777,N_14784);
or U15834 (N_15834,N_14479,N_14847);
nand U15835 (N_15835,N_14147,N_14520);
nor U15836 (N_15836,N_14496,N_13949);
nand U15837 (N_15837,N_14087,N_14228);
or U15838 (N_15838,N_14013,N_14652);
or U15839 (N_15839,N_13996,N_14932);
xor U15840 (N_15840,N_14968,N_13864);
nor U15841 (N_15841,N_13977,N_14205);
or U15842 (N_15842,N_13975,N_14221);
xor U15843 (N_15843,N_14597,N_14220);
nor U15844 (N_15844,N_14914,N_14177);
and U15845 (N_15845,N_14696,N_14115);
or U15846 (N_15846,N_14334,N_14997);
xnor U15847 (N_15847,N_13786,N_14395);
nand U15848 (N_15848,N_14920,N_14362);
and U15849 (N_15849,N_14963,N_14525);
and U15850 (N_15850,N_13878,N_14385);
nor U15851 (N_15851,N_13993,N_14061);
nor U15852 (N_15852,N_14746,N_14400);
and U15853 (N_15853,N_14962,N_14351);
nand U15854 (N_15854,N_14779,N_13844);
nor U15855 (N_15855,N_14960,N_14529);
or U15856 (N_15856,N_14592,N_14798);
or U15857 (N_15857,N_13987,N_13958);
nand U15858 (N_15858,N_14126,N_14922);
and U15859 (N_15859,N_14151,N_14266);
nand U15860 (N_15860,N_14416,N_14292);
xnor U15861 (N_15861,N_14947,N_13769);
and U15862 (N_15862,N_14967,N_14479);
nand U15863 (N_15863,N_13764,N_14191);
nand U15864 (N_15864,N_14740,N_14144);
xor U15865 (N_15865,N_13847,N_14036);
nor U15866 (N_15866,N_13829,N_13814);
or U15867 (N_15867,N_14442,N_14957);
or U15868 (N_15868,N_14518,N_14102);
xor U15869 (N_15869,N_13878,N_13965);
nor U15870 (N_15870,N_14218,N_13896);
nor U15871 (N_15871,N_14905,N_14544);
nor U15872 (N_15872,N_14511,N_13803);
and U15873 (N_15873,N_14003,N_14381);
and U15874 (N_15874,N_13764,N_14285);
or U15875 (N_15875,N_14657,N_14289);
nor U15876 (N_15876,N_14016,N_14619);
nor U15877 (N_15877,N_14003,N_14295);
nand U15878 (N_15878,N_14070,N_14167);
nand U15879 (N_15879,N_14135,N_14994);
nand U15880 (N_15880,N_14004,N_13894);
or U15881 (N_15881,N_14238,N_14215);
and U15882 (N_15882,N_14704,N_14061);
nand U15883 (N_15883,N_14850,N_14780);
nor U15884 (N_15884,N_14401,N_13982);
xor U15885 (N_15885,N_13810,N_14935);
nor U15886 (N_15886,N_14328,N_14853);
xnor U15887 (N_15887,N_14805,N_14572);
or U15888 (N_15888,N_14101,N_14317);
xor U15889 (N_15889,N_13951,N_13977);
nor U15890 (N_15890,N_13974,N_14071);
or U15891 (N_15891,N_14587,N_14973);
nor U15892 (N_15892,N_14311,N_14853);
or U15893 (N_15893,N_13876,N_14118);
and U15894 (N_15894,N_14723,N_14186);
and U15895 (N_15895,N_14301,N_14220);
xnor U15896 (N_15896,N_14291,N_14723);
and U15897 (N_15897,N_14771,N_14063);
nand U15898 (N_15898,N_13871,N_14800);
nand U15899 (N_15899,N_14344,N_13959);
nor U15900 (N_15900,N_14983,N_14616);
xor U15901 (N_15901,N_14423,N_14651);
xnor U15902 (N_15902,N_14670,N_14730);
and U15903 (N_15903,N_14920,N_14307);
nand U15904 (N_15904,N_14815,N_14919);
nor U15905 (N_15905,N_14415,N_14623);
nand U15906 (N_15906,N_14873,N_14537);
or U15907 (N_15907,N_14157,N_13879);
nor U15908 (N_15908,N_14476,N_14859);
and U15909 (N_15909,N_14658,N_14272);
nand U15910 (N_15910,N_14579,N_14751);
and U15911 (N_15911,N_14647,N_14255);
or U15912 (N_15912,N_14705,N_14140);
nand U15913 (N_15913,N_14100,N_14143);
nand U15914 (N_15914,N_14169,N_14102);
nand U15915 (N_15915,N_14059,N_14645);
nand U15916 (N_15916,N_14741,N_14272);
nor U15917 (N_15917,N_14516,N_14989);
or U15918 (N_15918,N_14185,N_14915);
or U15919 (N_15919,N_14468,N_14287);
or U15920 (N_15920,N_14563,N_14546);
nor U15921 (N_15921,N_14553,N_14240);
nor U15922 (N_15922,N_14555,N_13767);
or U15923 (N_15923,N_14369,N_14831);
nand U15924 (N_15924,N_13815,N_14471);
nand U15925 (N_15925,N_14274,N_14630);
nor U15926 (N_15926,N_14751,N_14505);
nand U15927 (N_15927,N_14796,N_14675);
nand U15928 (N_15928,N_14726,N_14868);
and U15929 (N_15929,N_14972,N_14356);
nand U15930 (N_15930,N_14195,N_14013);
xor U15931 (N_15931,N_13834,N_14478);
and U15932 (N_15932,N_14077,N_14369);
xor U15933 (N_15933,N_13857,N_14490);
xor U15934 (N_15934,N_14157,N_14496);
nor U15935 (N_15935,N_14460,N_14638);
nor U15936 (N_15936,N_14248,N_14927);
nand U15937 (N_15937,N_14169,N_13840);
or U15938 (N_15938,N_14064,N_14119);
xor U15939 (N_15939,N_13893,N_14764);
and U15940 (N_15940,N_13928,N_14541);
or U15941 (N_15941,N_13884,N_13779);
or U15942 (N_15942,N_14600,N_14061);
and U15943 (N_15943,N_14410,N_14701);
xor U15944 (N_15944,N_14515,N_13829);
nor U15945 (N_15945,N_14353,N_14183);
nor U15946 (N_15946,N_14259,N_14271);
and U15947 (N_15947,N_13845,N_14975);
and U15948 (N_15948,N_13859,N_14236);
nand U15949 (N_15949,N_14210,N_13849);
xnor U15950 (N_15950,N_14638,N_14502);
nand U15951 (N_15951,N_13938,N_14434);
xor U15952 (N_15952,N_14653,N_13756);
nand U15953 (N_15953,N_14760,N_14844);
nand U15954 (N_15954,N_14482,N_14132);
or U15955 (N_15955,N_14544,N_14575);
nand U15956 (N_15956,N_13829,N_14350);
nand U15957 (N_15957,N_13938,N_14315);
nor U15958 (N_15958,N_13894,N_13848);
nor U15959 (N_15959,N_14914,N_14951);
nand U15960 (N_15960,N_14993,N_14125);
nor U15961 (N_15961,N_14256,N_14320);
nand U15962 (N_15962,N_14961,N_14006);
nand U15963 (N_15963,N_14106,N_14099);
nand U15964 (N_15964,N_14590,N_13864);
and U15965 (N_15965,N_14839,N_13793);
nand U15966 (N_15966,N_14795,N_14021);
or U15967 (N_15967,N_13883,N_14408);
or U15968 (N_15968,N_14069,N_14378);
nor U15969 (N_15969,N_14046,N_14258);
nor U15970 (N_15970,N_14878,N_13890);
and U15971 (N_15971,N_13966,N_14999);
xnor U15972 (N_15972,N_14420,N_13851);
xor U15973 (N_15973,N_14517,N_14186);
nand U15974 (N_15974,N_14774,N_13968);
nor U15975 (N_15975,N_14655,N_14967);
nor U15976 (N_15976,N_14476,N_13967);
and U15977 (N_15977,N_13890,N_14792);
xor U15978 (N_15978,N_13859,N_14286);
xnor U15979 (N_15979,N_14753,N_14565);
or U15980 (N_15980,N_14581,N_14673);
xnor U15981 (N_15981,N_14310,N_14629);
or U15982 (N_15982,N_14097,N_13970);
nor U15983 (N_15983,N_13775,N_14165);
nand U15984 (N_15984,N_14929,N_14542);
and U15985 (N_15985,N_14742,N_14353);
nand U15986 (N_15986,N_14590,N_14340);
or U15987 (N_15987,N_14670,N_13837);
xor U15988 (N_15988,N_14593,N_14147);
or U15989 (N_15989,N_13857,N_14608);
nand U15990 (N_15990,N_14467,N_14001);
and U15991 (N_15991,N_14914,N_13952);
xnor U15992 (N_15992,N_14258,N_14078);
or U15993 (N_15993,N_14869,N_14900);
xor U15994 (N_15994,N_14420,N_14150);
and U15995 (N_15995,N_13944,N_14606);
nor U15996 (N_15996,N_14635,N_13958);
or U15997 (N_15997,N_13805,N_13890);
xnor U15998 (N_15998,N_14866,N_14442);
or U15999 (N_15999,N_14525,N_14410);
nand U16000 (N_16000,N_14194,N_14970);
and U16001 (N_16001,N_13879,N_14760);
or U16002 (N_16002,N_13765,N_14769);
or U16003 (N_16003,N_14927,N_14264);
xnor U16004 (N_16004,N_13982,N_14999);
nor U16005 (N_16005,N_14312,N_14299);
nand U16006 (N_16006,N_14068,N_14764);
or U16007 (N_16007,N_14707,N_14377);
nor U16008 (N_16008,N_13793,N_14879);
xor U16009 (N_16009,N_14263,N_14521);
nor U16010 (N_16010,N_14231,N_14532);
nand U16011 (N_16011,N_14649,N_14051);
or U16012 (N_16012,N_14690,N_14514);
nor U16013 (N_16013,N_14395,N_14962);
and U16014 (N_16014,N_14986,N_14373);
nand U16015 (N_16015,N_13866,N_14191);
xor U16016 (N_16016,N_13983,N_13868);
or U16017 (N_16017,N_14034,N_14739);
nand U16018 (N_16018,N_14126,N_13929);
xnor U16019 (N_16019,N_14894,N_14859);
nor U16020 (N_16020,N_14850,N_14670);
nand U16021 (N_16021,N_14421,N_13787);
xnor U16022 (N_16022,N_13999,N_13875);
xor U16023 (N_16023,N_14227,N_13866);
nor U16024 (N_16024,N_14180,N_13917);
or U16025 (N_16025,N_13948,N_14788);
or U16026 (N_16026,N_13779,N_14327);
nand U16027 (N_16027,N_13938,N_13790);
or U16028 (N_16028,N_14943,N_13770);
or U16029 (N_16029,N_14628,N_14443);
xnor U16030 (N_16030,N_14196,N_13907);
xor U16031 (N_16031,N_14952,N_14361);
or U16032 (N_16032,N_14102,N_14249);
nand U16033 (N_16033,N_14793,N_14820);
or U16034 (N_16034,N_14510,N_14798);
xor U16035 (N_16035,N_14271,N_14784);
nor U16036 (N_16036,N_14559,N_13837);
xnor U16037 (N_16037,N_14234,N_13976);
or U16038 (N_16038,N_13864,N_14301);
and U16039 (N_16039,N_14057,N_13906);
or U16040 (N_16040,N_13966,N_14952);
and U16041 (N_16041,N_14923,N_14407);
xnor U16042 (N_16042,N_14072,N_14057);
xor U16043 (N_16043,N_14271,N_14102);
or U16044 (N_16044,N_14370,N_14053);
or U16045 (N_16045,N_13981,N_13799);
nand U16046 (N_16046,N_14024,N_14263);
nand U16047 (N_16047,N_14097,N_13854);
or U16048 (N_16048,N_14627,N_14058);
or U16049 (N_16049,N_14444,N_14253);
and U16050 (N_16050,N_14755,N_14545);
nand U16051 (N_16051,N_14754,N_14962);
nor U16052 (N_16052,N_14372,N_14076);
and U16053 (N_16053,N_14301,N_14618);
xnor U16054 (N_16054,N_14945,N_13957);
nand U16055 (N_16055,N_13976,N_14118);
nor U16056 (N_16056,N_13783,N_14129);
xnor U16057 (N_16057,N_13874,N_14457);
and U16058 (N_16058,N_14240,N_13796);
xor U16059 (N_16059,N_14850,N_13857);
or U16060 (N_16060,N_14423,N_14910);
and U16061 (N_16061,N_14692,N_14675);
or U16062 (N_16062,N_14936,N_13837);
xor U16063 (N_16063,N_14776,N_14082);
nand U16064 (N_16064,N_14301,N_14842);
nor U16065 (N_16065,N_14027,N_14962);
and U16066 (N_16066,N_13887,N_14943);
or U16067 (N_16067,N_13876,N_14143);
and U16068 (N_16068,N_14086,N_13987);
and U16069 (N_16069,N_14068,N_14345);
xnor U16070 (N_16070,N_14086,N_13787);
nand U16071 (N_16071,N_14600,N_13772);
nand U16072 (N_16072,N_13904,N_14480);
and U16073 (N_16073,N_14545,N_14930);
or U16074 (N_16074,N_13895,N_14679);
nor U16075 (N_16075,N_13869,N_14210);
and U16076 (N_16076,N_14930,N_14849);
and U16077 (N_16077,N_14814,N_14333);
nor U16078 (N_16078,N_13805,N_14919);
and U16079 (N_16079,N_14573,N_14768);
nor U16080 (N_16080,N_13782,N_14166);
and U16081 (N_16081,N_14767,N_13932);
nor U16082 (N_16082,N_14054,N_14379);
nor U16083 (N_16083,N_13793,N_14053);
and U16084 (N_16084,N_14039,N_14816);
nand U16085 (N_16085,N_14614,N_14008);
xor U16086 (N_16086,N_13999,N_14633);
nand U16087 (N_16087,N_14827,N_14832);
or U16088 (N_16088,N_13781,N_14319);
or U16089 (N_16089,N_14117,N_14609);
xor U16090 (N_16090,N_14077,N_14501);
xor U16091 (N_16091,N_13779,N_13826);
or U16092 (N_16092,N_13750,N_14830);
or U16093 (N_16093,N_14739,N_14348);
or U16094 (N_16094,N_14643,N_14522);
nand U16095 (N_16095,N_14057,N_13820);
nor U16096 (N_16096,N_14333,N_13832);
and U16097 (N_16097,N_13876,N_14147);
xnor U16098 (N_16098,N_14480,N_14909);
or U16099 (N_16099,N_14889,N_14616);
or U16100 (N_16100,N_14303,N_13997);
nand U16101 (N_16101,N_14622,N_14882);
xor U16102 (N_16102,N_14640,N_14511);
nor U16103 (N_16103,N_13784,N_13759);
and U16104 (N_16104,N_14862,N_14306);
nor U16105 (N_16105,N_14602,N_14724);
xnor U16106 (N_16106,N_14446,N_13819);
xor U16107 (N_16107,N_14162,N_14110);
nand U16108 (N_16108,N_13942,N_14422);
nand U16109 (N_16109,N_14870,N_14585);
and U16110 (N_16110,N_14170,N_13886);
or U16111 (N_16111,N_14604,N_14157);
nand U16112 (N_16112,N_13962,N_14601);
and U16113 (N_16113,N_14348,N_14626);
nor U16114 (N_16114,N_14060,N_14702);
xnor U16115 (N_16115,N_14245,N_14392);
nor U16116 (N_16116,N_14732,N_14697);
or U16117 (N_16117,N_14471,N_13985);
xnor U16118 (N_16118,N_14387,N_14440);
nand U16119 (N_16119,N_14960,N_14591);
xor U16120 (N_16120,N_13759,N_13913);
or U16121 (N_16121,N_14215,N_14875);
nor U16122 (N_16122,N_14234,N_14656);
nand U16123 (N_16123,N_14684,N_14686);
nand U16124 (N_16124,N_14970,N_14471);
or U16125 (N_16125,N_13797,N_14317);
or U16126 (N_16126,N_13844,N_14888);
xor U16127 (N_16127,N_13826,N_14897);
or U16128 (N_16128,N_14463,N_14567);
nor U16129 (N_16129,N_14387,N_13841);
nor U16130 (N_16130,N_14835,N_13927);
nor U16131 (N_16131,N_14615,N_14304);
and U16132 (N_16132,N_14637,N_14800);
and U16133 (N_16133,N_14976,N_14569);
or U16134 (N_16134,N_14411,N_13814);
nor U16135 (N_16135,N_14929,N_13946);
and U16136 (N_16136,N_14144,N_14252);
and U16137 (N_16137,N_14490,N_13786);
or U16138 (N_16138,N_14133,N_14461);
or U16139 (N_16139,N_13750,N_14349);
nor U16140 (N_16140,N_14726,N_14417);
nand U16141 (N_16141,N_13810,N_14634);
xnor U16142 (N_16142,N_14248,N_13802);
nand U16143 (N_16143,N_13930,N_14029);
nor U16144 (N_16144,N_13934,N_14057);
or U16145 (N_16145,N_14384,N_14645);
and U16146 (N_16146,N_14991,N_14597);
xor U16147 (N_16147,N_14259,N_13810);
and U16148 (N_16148,N_14483,N_14599);
xnor U16149 (N_16149,N_14774,N_13872);
xnor U16150 (N_16150,N_14684,N_14958);
or U16151 (N_16151,N_14586,N_14117);
nand U16152 (N_16152,N_14945,N_14183);
xnor U16153 (N_16153,N_14683,N_13934);
xnor U16154 (N_16154,N_13852,N_14333);
or U16155 (N_16155,N_13873,N_14629);
and U16156 (N_16156,N_13897,N_14101);
xnor U16157 (N_16157,N_14330,N_14397);
nor U16158 (N_16158,N_14768,N_14236);
and U16159 (N_16159,N_14370,N_14311);
xnor U16160 (N_16160,N_13817,N_14536);
or U16161 (N_16161,N_14432,N_14840);
or U16162 (N_16162,N_13788,N_14647);
or U16163 (N_16163,N_14994,N_14897);
nand U16164 (N_16164,N_14436,N_14592);
nand U16165 (N_16165,N_14545,N_13849);
and U16166 (N_16166,N_14344,N_14319);
nor U16167 (N_16167,N_14634,N_14672);
xnor U16168 (N_16168,N_13942,N_14368);
xor U16169 (N_16169,N_13955,N_14016);
nor U16170 (N_16170,N_14700,N_14408);
or U16171 (N_16171,N_14966,N_14235);
and U16172 (N_16172,N_14913,N_14993);
nor U16173 (N_16173,N_14225,N_14466);
and U16174 (N_16174,N_14790,N_14245);
nand U16175 (N_16175,N_14848,N_14470);
or U16176 (N_16176,N_14693,N_14094);
xor U16177 (N_16177,N_14766,N_14807);
nand U16178 (N_16178,N_14024,N_14719);
nand U16179 (N_16179,N_14882,N_14210);
nand U16180 (N_16180,N_14628,N_14281);
and U16181 (N_16181,N_13812,N_14447);
xnor U16182 (N_16182,N_14556,N_14761);
nor U16183 (N_16183,N_14465,N_14894);
and U16184 (N_16184,N_13827,N_14785);
nand U16185 (N_16185,N_14269,N_13825);
xnor U16186 (N_16186,N_14489,N_13788);
xor U16187 (N_16187,N_14518,N_14362);
xor U16188 (N_16188,N_14229,N_14706);
or U16189 (N_16189,N_14958,N_13772);
nand U16190 (N_16190,N_14350,N_13770);
xnor U16191 (N_16191,N_14180,N_14758);
and U16192 (N_16192,N_14884,N_14789);
nor U16193 (N_16193,N_14131,N_14917);
nand U16194 (N_16194,N_14898,N_13861);
or U16195 (N_16195,N_14061,N_14343);
xor U16196 (N_16196,N_14648,N_14786);
and U16197 (N_16197,N_14228,N_14584);
and U16198 (N_16198,N_14386,N_14808);
nor U16199 (N_16199,N_14407,N_14994);
xor U16200 (N_16200,N_14668,N_14907);
xnor U16201 (N_16201,N_13922,N_14707);
nand U16202 (N_16202,N_13776,N_14235);
and U16203 (N_16203,N_13831,N_14715);
xor U16204 (N_16204,N_13818,N_14796);
and U16205 (N_16205,N_14789,N_14188);
xnor U16206 (N_16206,N_14496,N_14330);
and U16207 (N_16207,N_14060,N_14927);
or U16208 (N_16208,N_13752,N_13842);
nor U16209 (N_16209,N_14444,N_14140);
or U16210 (N_16210,N_14336,N_13956);
xnor U16211 (N_16211,N_14983,N_14152);
and U16212 (N_16212,N_14611,N_14155);
or U16213 (N_16213,N_14752,N_14530);
and U16214 (N_16214,N_14102,N_14772);
xor U16215 (N_16215,N_13904,N_14502);
or U16216 (N_16216,N_14027,N_14002);
and U16217 (N_16217,N_14943,N_14461);
nor U16218 (N_16218,N_14073,N_13991);
nor U16219 (N_16219,N_14361,N_14960);
nor U16220 (N_16220,N_14490,N_14192);
and U16221 (N_16221,N_14210,N_14693);
nand U16222 (N_16222,N_14873,N_14138);
or U16223 (N_16223,N_14183,N_13763);
and U16224 (N_16224,N_14386,N_13762);
or U16225 (N_16225,N_14518,N_14360);
xor U16226 (N_16226,N_13869,N_14575);
nand U16227 (N_16227,N_14721,N_14103);
nand U16228 (N_16228,N_13981,N_14411);
nor U16229 (N_16229,N_14193,N_14264);
or U16230 (N_16230,N_14244,N_13970);
or U16231 (N_16231,N_14489,N_14531);
nand U16232 (N_16232,N_14847,N_14840);
and U16233 (N_16233,N_13845,N_13846);
xnor U16234 (N_16234,N_13964,N_14103);
and U16235 (N_16235,N_14276,N_14458);
nor U16236 (N_16236,N_13800,N_14275);
xnor U16237 (N_16237,N_13926,N_14108);
nand U16238 (N_16238,N_14046,N_14142);
and U16239 (N_16239,N_13754,N_14403);
nand U16240 (N_16240,N_14322,N_14015);
and U16241 (N_16241,N_14757,N_13755);
nand U16242 (N_16242,N_14321,N_14800);
nand U16243 (N_16243,N_13824,N_14168);
and U16244 (N_16244,N_14759,N_14143);
nor U16245 (N_16245,N_14597,N_13843);
or U16246 (N_16246,N_13868,N_14041);
and U16247 (N_16247,N_13833,N_14298);
and U16248 (N_16248,N_13802,N_14453);
nand U16249 (N_16249,N_14625,N_14015);
xnor U16250 (N_16250,N_15130,N_15970);
nand U16251 (N_16251,N_15938,N_15770);
nand U16252 (N_16252,N_15926,N_15417);
nor U16253 (N_16253,N_15112,N_15351);
and U16254 (N_16254,N_16083,N_15355);
nand U16255 (N_16255,N_15369,N_15301);
and U16256 (N_16256,N_15051,N_15203);
or U16257 (N_16257,N_15454,N_15491);
nor U16258 (N_16258,N_16210,N_15471);
nand U16259 (N_16259,N_15577,N_15319);
xor U16260 (N_16260,N_15478,N_15264);
nor U16261 (N_16261,N_15704,N_15699);
or U16262 (N_16262,N_15661,N_15107);
or U16263 (N_16263,N_15860,N_16229);
xnor U16264 (N_16264,N_15855,N_16107);
nand U16265 (N_16265,N_15487,N_16040);
nand U16266 (N_16266,N_15888,N_16235);
nor U16267 (N_16267,N_15912,N_15984);
xor U16268 (N_16268,N_15324,N_16221);
and U16269 (N_16269,N_15019,N_15354);
and U16270 (N_16270,N_15286,N_15435);
xor U16271 (N_16271,N_15509,N_15200);
or U16272 (N_16272,N_15928,N_15557);
xor U16273 (N_16273,N_15348,N_16049);
nand U16274 (N_16274,N_15421,N_15458);
nand U16275 (N_16275,N_16120,N_15309);
and U16276 (N_16276,N_16013,N_15931);
nand U16277 (N_16277,N_15409,N_15574);
nand U16278 (N_16278,N_16226,N_16145);
or U16279 (N_16279,N_15238,N_15433);
nand U16280 (N_16280,N_16177,N_15016);
and U16281 (N_16281,N_16023,N_15958);
nor U16282 (N_16282,N_15767,N_15386);
nand U16283 (N_16283,N_16183,N_15973);
and U16284 (N_16284,N_15066,N_15990);
nand U16285 (N_16285,N_15793,N_15282);
and U16286 (N_16286,N_15545,N_15546);
nand U16287 (N_16287,N_15356,N_15617);
or U16288 (N_16288,N_16154,N_16127);
or U16289 (N_16289,N_15105,N_15539);
nor U16290 (N_16290,N_16108,N_15028);
and U16291 (N_16291,N_15822,N_15812);
nand U16292 (N_16292,N_16129,N_15100);
or U16293 (N_16293,N_15663,N_15749);
and U16294 (N_16294,N_15675,N_15117);
and U16295 (N_16295,N_16042,N_15394);
or U16296 (N_16296,N_15082,N_16173);
xnor U16297 (N_16297,N_15195,N_15963);
and U16298 (N_16298,N_15125,N_15366);
xnor U16299 (N_16299,N_15978,N_15263);
and U16300 (N_16300,N_15731,N_15897);
and U16301 (N_16301,N_15833,N_15845);
and U16302 (N_16302,N_15173,N_15153);
and U16303 (N_16303,N_15053,N_16112);
xor U16304 (N_16304,N_16068,N_15152);
nor U16305 (N_16305,N_15279,N_15490);
and U16306 (N_16306,N_15875,N_15087);
nor U16307 (N_16307,N_15229,N_15951);
nor U16308 (N_16308,N_16078,N_15843);
xnor U16309 (N_16309,N_15725,N_15123);
nor U16310 (N_16310,N_15469,N_15939);
or U16311 (N_16311,N_15806,N_15294);
and U16312 (N_16312,N_15538,N_15601);
and U16313 (N_16313,N_15726,N_15586);
nor U16314 (N_16314,N_15135,N_15077);
or U16315 (N_16315,N_15465,N_15742);
and U16316 (N_16316,N_15643,N_16220);
xor U16317 (N_16317,N_15404,N_15936);
and U16318 (N_16318,N_16224,N_15657);
nor U16319 (N_16319,N_16181,N_15995);
nor U16320 (N_16320,N_16062,N_15341);
or U16321 (N_16321,N_16111,N_15187);
xnor U16322 (N_16322,N_15484,N_15694);
or U16323 (N_16323,N_16237,N_15473);
and U16324 (N_16324,N_15868,N_16004);
xnor U16325 (N_16325,N_15623,N_15411);
xor U16326 (N_16326,N_15737,N_16222);
and U16327 (N_16327,N_16170,N_15405);
or U16328 (N_16328,N_15240,N_15798);
nor U16329 (N_16329,N_15083,N_15442);
nand U16330 (N_16330,N_15246,N_16072);
or U16331 (N_16331,N_15878,N_16217);
nor U16332 (N_16332,N_15204,N_15450);
nor U16333 (N_16333,N_15278,N_15089);
xnor U16334 (N_16334,N_15296,N_15647);
nand U16335 (N_16335,N_15390,N_15228);
nand U16336 (N_16336,N_15470,N_15714);
xnor U16337 (N_16337,N_15242,N_15856);
nor U16338 (N_16338,N_15965,N_15250);
and U16339 (N_16339,N_15558,N_15804);
nor U16340 (N_16340,N_15646,N_15413);
nor U16341 (N_16341,N_15498,N_16071);
nand U16342 (N_16342,N_15660,N_16060);
xor U16343 (N_16343,N_16169,N_15190);
nand U16344 (N_16344,N_16219,N_15924);
nor U16345 (N_16345,N_15476,N_15841);
xor U16346 (N_16346,N_15058,N_15998);
nor U16347 (N_16347,N_15175,N_15245);
nor U16348 (N_16348,N_16162,N_15779);
or U16349 (N_16349,N_16191,N_15482);
or U16350 (N_16350,N_15099,N_15680);
or U16351 (N_16351,N_15813,N_15085);
or U16352 (N_16352,N_15340,N_16234);
and U16353 (N_16353,N_15270,N_16212);
or U16354 (N_16354,N_15684,N_15604);
or U16355 (N_16355,N_15292,N_16048);
nor U16356 (N_16356,N_15441,N_15853);
or U16357 (N_16357,N_15588,N_15093);
xor U16358 (N_16358,N_15371,N_15464);
nand U16359 (N_16359,N_16018,N_15969);
nand U16360 (N_16360,N_15560,N_15671);
nor U16361 (N_16361,N_15015,N_15313);
xor U16362 (N_16362,N_15687,N_16115);
nand U16363 (N_16363,N_15307,N_15126);
xor U16364 (N_16364,N_15649,N_16090);
or U16365 (N_16365,N_15258,N_15955);
nand U16366 (N_16366,N_16184,N_16079);
nor U16367 (N_16367,N_15373,N_15511);
and U16368 (N_16368,N_15254,N_15257);
xor U16369 (N_16369,N_15773,N_15420);
nand U16370 (N_16370,N_15920,N_15035);
nand U16371 (N_16371,N_15846,N_15344);
nor U16372 (N_16372,N_16092,N_15243);
and U16373 (N_16373,N_15662,N_15947);
xor U16374 (N_16374,N_15724,N_15885);
nand U16375 (N_16375,N_16139,N_15131);
and U16376 (N_16376,N_16053,N_15437);
nand U16377 (N_16377,N_15440,N_15041);
and U16378 (N_16378,N_15320,N_15987);
nand U16379 (N_16379,N_15052,N_15055);
nand U16380 (N_16380,N_15345,N_15104);
or U16381 (N_16381,N_15328,N_15139);
nand U16382 (N_16382,N_16244,N_16093);
nand U16383 (N_16383,N_15388,N_15350);
nand U16384 (N_16384,N_15580,N_15284);
and U16385 (N_16385,N_15311,N_16179);
xor U16386 (N_16386,N_16006,N_15525);
nor U16387 (N_16387,N_15039,N_15766);
nor U16388 (N_16388,N_15962,N_15732);
xor U16389 (N_16389,N_15907,N_16246);
or U16390 (N_16390,N_15098,N_15029);
xnor U16391 (N_16391,N_16082,N_15431);
xor U16392 (N_16392,N_15740,N_15480);
and U16393 (N_16393,N_15882,N_15327);
and U16394 (N_16394,N_15786,N_15976);
and U16395 (N_16395,N_15049,N_15864);
nor U16396 (N_16396,N_15909,N_15971);
or U16397 (N_16397,N_16094,N_15475);
and U16398 (N_16398,N_15408,N_15391);
nand U16399 (N_16399,N_16011,N_15669);
or U16400 (N_16400,N_15208,N_15664);
nand U16401 (N_16401,N_15196,N_15628);
xnor U16402 (N_16402,N_15738,N_15997);
and U16403 (N_16403,N_16105,N_15225);
or U16404 (N_16404,N_15956,N_15518);
xor U16405 (N_16405,N_16225,N_15559);
nand U16406 (N_16406,N_16102,N_15206);
nand U16407 (N_16407,N_15893,N_15268);
xor U16408 (N_16408,N_15552,N_16178);
nand U16409 (N_16409,N_15038,N_15202);
nand U16410 (N_16410,N_15718,N_16084);
nor U16411 (N_16411,N_16003,N_16027);
nor U16412 (N_16412,N_15692,N_15572);
nor U16413 (N_16413,N_15721,N_15727);
or U16414 (N_16414,N_15137,N_15387);
xor U16415 (N_16415,N_15067,N_15095);
and U16416 (N_16416,N_15269,N_15199);
nand U16417 (N_16417,N_15748,N_15462);
nand U16418 (N_16418,N_15784,N_15445);
or U16419 (N_16419,N_15312,N_15753);
and U16420 (N_16420,N_15744,N_16052);
xnor U16421 (N_16421,N_15873,N_15554);
nor U16422 (N_16422,N_15362,N_15803);
nand U16423 (N_16423,N_16054,N_15815);
and U16424 (N_16424,N_15068,N_15638);
xor U16425 (N_16425,N_15050,N_15443);
and U16426 (N_16426,N_15565,N_15548);
nor U16427 (N_16427,N_15707,N_15180);
nand U16428 (N_16428,N_16138,N_15094);
or U16429 (N_16429,N_15674,N_15523);
and U16430 (N_16430,N_16058,N_15876);
and U16431 (N_16431,N_15788,N_15211);
nand U16432 (N_16432,N_15004,N_15221);
nor U16433 (N_16433,N_16020,N_15508);
xnor U16434 (N_16434,N_15233,N_16242);
xnor U16435 (N_16435,N_15020,N_15210);
nor U16436 (N_16436,N_15375,N_16156);
or U16437 (N_16437,N_15556,N_15380);
and U16438 (N_16438,N_15310,N_15046);
nor U16439 (N_16439,N_16016,N_15468);
nor U16440 (N_16440,N_15519,N_15616);
and U16441 (N_16441,N_16041,N_15585);
and U16442 (N_16442,N_15755,N_15715);
or U16443 (N_16443,N_15459,N_15584);
or U16444 (N_16444,N_15639,N_15814);
or U16445 (N_16445,N_15506,N_15184);
nand U16446 (N_16446,N_15881,N_15600);
nand U16447 (N_16447,N_16119,N_15834);
nor U16448 (N_16448,N_15591,N_15280);
xnor U16449 (N_16449,N_16085,N_15863);
nand U16450 (N_16450,N_15308,N_16168);
or U16451 (N_16451,N_15503,N_15502);
and U16452 (N_16452,N_15781,N_15810);
and U16453 (N_16453,N_15492,N_15101);
or U16454 (N_16454,N_15836,N_15866);
xnor U16455 (N_16455,N_16194,N_15166);
and U16456 (N_16456,N_16061,N_15119);
and U16457 (N_16457,N_15181,N_15385);
and U16458 (N_16458,N_16035,N_15381);
or U16459 (N_16459,N_15446,N_15842);
xor U16460 (N_16460,N_16007,N_15378);
nor U16461 (N_16461,N_16103,N_15595);
nor U16462 (N_16462,N_15553,N_15857);
nor U16463 (N_16463,N_16158,N_16073);
or U16464 (N_16464,N_15261,N_15384);
and U16465 (N_16465,N_15921,N_15274);
nand U16466 (N_16466,N_15343,N_15383);
nand U16467 (N_16467,N_16233,N_15696);
xnor U16468 (N_16468,N_15031,N_15143);
nand U16469 (N_16469,N_16200,N_15256);
and U16470 (N_16470,N_15630,N_15967);
and U16471 (N_16471,N_15422,N_15949);
xnor U16472 (N_16472,N_15006,N_16151);
nand U16473 (N_16473,N_15013,N_15392);
xnor U16474 (N_16474,N_15259,N_15412);
nor U16475 (N_16475,N_15132,N_15494);
or U16476 (N_16476,N_16069,N_15379);
nor U16477 (N_16477,N_15772,N_15064);
and U16478 (N_16478,N_15960,N_15870);
or U16479 (N_16479,N_15654,N_16187);
nand U16480 (N_16480,N_15697,N_15722);
nand U16481 (N_16481,N_15197,N_15914);
and U16482 (N_16482,N_15075,N_15711);
nor U16483 (N_16483,N_15406,N_15449);
and U16484 (N_16484,N_15787,N_16017);
or U16485 (N_16485,N_16051,N_15612);
xor U16486 (N_16486,N_15795,N_15592);
and U16487 (N_16487,N_15542,N_16193);
and U16488 (N_16488,N_15040,N_15042);
nor U16489 (N_16489,N_15136,N_15402);
nand U16490 (N_16490,N_15235,N_15410);
and U16491 (N_16491,N_15564,N_15666);
and U16492 (N_16492,N_15763,N_15683);
and U16493 (N_16493,N_15000,N_15453);
or U16494 (N_16494,N_15879,N_15705);
and U16495 (N_16495,N_15377,N_15934);
nor U16496 (N_16496,N_15782,N_15801);
xor U16497 (N_16497,N_15957,N_15447);
nor U16498 (N_16498,N_15505,N_15636);
or U16499 (N_16499,N_15522,N_16230);
nor U16500 (N_16500,N_15644,N_15218);
or U16501 (N_16501,N_16218,N_15824);
and U16502 (N_16502,N_15608,N_15809);
or U16503 (N_16503,N_16149,N_15906);
nor U16504 (N_16504,N_15589,N_15232);
xnor U16505 (N_16505,N_15959,N_15890);
nor U16506 (N_16506,N_15562,N_15544);
and U16507 (N_16507,N_16022,N_16086);
or U16508 (N_16508,N_15178,N_15528);
nor U16509 (N_16509,N_15339,N_15305);
nand U16510 (N_16510,N_15950,N_16148);
or U16511 (N_16511,N_16046,N_16021);
nor U16512 (N_16512,N_15037,N_15819);
xor U16513 (N_16513,N_15504,N_16172);
xor U16514 (N_16514,N_16063,N_15656);
xor U16515 (N_16515,N_15302,N_15436);
or U16516 (N_16516,N_15485,N_15764);
nor U16517 (N_16517,N_15156,N_15551);
or U16518 (N_16518,N_15874,N_15342);
xor U16519 (N_16519,N_15164,N_16197);
nor U16520 (N_16520,N_15014,N_15393);
xor U16521 (N_16521,N_15635,N_15414);
and U16522 (N_16522,N_15376,N_15260);
nor U16523 (N_16523,N_15317,N_16088);
nor U16524 (N_16524,N_15102,N_15062);
nor U16525 (N_16525,N_15529,N_15789);
nor U16526 (N_16526,N_15072,N_15444);
nor U16527 (N_16527,N_15847,N_16249);
and U16528 (N_16528,N_15266,N_15226);
nand U16529 (N_16529,N_15059,N_15398);
nand U16530 (N_16530,N_15188,N_15273);
xor U16531 (N_16531,N_15536,N_15625);
or U16532 (N_16532,N_15061,N_16089);
nor U16533 (N_16533,N_15964,N_15207);
or U16534 (N_16534,N_16030,N_16248);
nor U16535 (N_16535,N_15018,N_15905);
nor U16536 (N_16536,N_16232,N_15849);
nor U16537 (N_16537,N_16070,N_15360);
nand U16538 (N_16538,N_15079,N_16064);
or U16539 (N_16539,N_15658,N_16029);
and U16540 (N_16540,N_16125,N_15255);
nand U16541 (N_16541,N_15710,N_15757);
nor U16542 (N_16542,N_15179,N_15512);
nor U16543 (N_16543,N_15507,N_16207);
and U16544 (N_16544,N_16171,N_15673);
nand U16545 (N_16545,N_15216,N_15561);
or U16546 (N_16546,N_15768,N_16015);
or U16547 (N_16547,N_16157,N_16198);
nand U16548 (N_16548,N_15330,N_15872);
or U16549 (N_16549,N_15220,N_15155);
nor U16550 (N_16550,N_15891,N_16160);
and U16551 (N_16551,N_15792,N_15916);
or U16552 (N_16552,N_15747,N_16159);
nor U16553 (N_16553,N_16012,N_15982);
and U16554 (N_16554,N_15915,N_15579);
and U16555 (N_16555,N_15937,N_15713);
or U16556 (N_16556,N_16142,N_15986);
and U16557 (N_16557,N_15267,N_15057);
xnor U16558 (N_16558,N_15641,N_15651);
nor U16559 (N_16559,N_16247,N_15415);
nand U16560 (N_16560,N_15746,N_15637);
or U16561 (N_16561,N_16096,N_16009);
xor U16562 (N_16562,N_15852,N_15823);
nand U16563 (N_16563,N_15448,N_15160);
and U16564 (N_16564,N_15821,N_15850);
nor U16565 (N_16565,N_15290,N_15213);
and U16566 (N_16566,N_15115,N_15429);
xnor U16567 (N_16567,N_15403,N_15432);
and U16568 (N_16568,N_16039,N_15794);
or U16569 (N_16569,N_15128,N_15659);
or U16570 (N_16570,N_15515,N_15993);
xor U16571 (N_16571,N_15854,N_16155);
nor U16572 (N_16572,N_15337,N_15602);
xnor U16573 (N_16573,N_15975,N_15182);
nor U16574 (N_16574,N_15165,N_15146);
or U16575 (N_16575,N_16121,N_16065);
xnor U16576 (N_16576,N_16190,N_15114);
and U16577 (N_16577,N_15543,N_15516);
xnor U16578 (N_16578,N_15698,N_15321);
and U16579 (N_16579,N_15493,N_15474);
nand U16580 (N_16580,N_15865,N_15289);
and U16581 (N_16581,N_15596,N_15839);
nor U16582 (N_16582,N_15291,N_15904);
nor U16583 (N_16583,N_15036,N_15489);
xor U16584 (N_16584,N_15730,N_15681);
xor U16585 (N_16585,N_15010,N_15609);
or U16586 (N_16586,N_15729,N_15158);
or U16587 (N_16587,N_15761,N_15800);
nand U16588 (N_16588,N_15288,N_15838);
xor U16589 (N_16589,N_16240,N_16206);
xnor U16590 (N_16590,N_16005,N_16123);
nand U16591 (N_16591,N_15008,N_15370);
or U16592 (N_16592,N_16141,N_15954);
xnor U16593 (N_16593,N_15108,N_16067);
nor U16594 (N_16594,N_15887,N_16223);
and U16595 (N_16595,N_15778,N_16161);
nor U16596 (N_16596,N_15594,N_15048);
and U16597 (N_16597,N_16081,N_16147);
nand U16598 (N_16598,N_15347,N_15106);
nand U16599 (N_16599,N_15032,N_15120);
nor U16600 (N_16600,N_15816,N_15603);
or U16601 (N_16601,N_15901,N_15626);
nor U16602 (N_16602,N_15428,N_15080);
nand U16603 (N_16603,N_15599,N_15790);
and U16604 (N_16604,N_15510,N_15201);
xor U16605 (N_16605,N_15023,N_15996);
and U16606 (N_16606,N_16126,N_16214);
xor U16607 (N_16607,N_15946,N_15071);
and U16608 (N_16608,N_16166,N_15030);
and U16609 (N_16609,N_15940,N_15776);
and U16610 (N_16610,N_16034,N_15497);
nand U16611 (N_16611,N_15111,N_15176);
nor U16612 (N_16612,N_15265,N_15249);
xor U16613 (N_16613,N_15500,N_16095);
nand U16614 (N_16614,N_15452,N_16231);
or U16615 (N_16615,N_16001,N_15871);
nor U16616 (N_16616,N_16010,N_15483);
or U16617 (N_16617,N_15917,N_16080);
nand U16618 (N_16618,N_15122,N_15769);
or U16619 (N_16619,N_15808,N_15648);
xor U16620 (N_16620,N_15933,N_15253);
xnor U16621 (N_16621,N_15520,N_15336);
or U16622 (N_16622,N_15169,N_15192);
nor U16623 (N_16623,N_15531,N_15247);
nor U16624 (N_16624,N_15894,N_16047);
nand U16625 (N_16625,N_15419,N_15331);
xor U16626 (N_16626,N_15695,N_15418);
and U16627 (N_16627,N_15365,N_15820);
nand U16628 (N_16628,N_15241,N_15363);
xnor U16629 (N_16629,N_15081,N_16074);
or U16630 (N_16630,N_15495,N_15183);
xor U16631 (N_16631,N_15719,N_16146);
and U16632 (N_16632,N_15368,N_15709);
and U16633 (N_16633,N_15091,N_15239);
and U16634 (N_16634,N_15981,N_16199);
xor U16635 (N_16635,N_15172,N_15252);
nor U16636 (N_16636,N_15582,N_15943);
or U16637 (N_16637,N_15622,N_15895);
xor U16638 (N_16638,N_15389,N_15227);
nor U16639 (N_16639,N_15382,N_15598);
nor U16640 (N_16640,N_15802,N_15831);
nand U16641 (N_16641,N_15688,N_15298);
xnor U16642 (N_16642,N_15499,N_15027);
and U16643 (N_16643,N_15848,N_16195);
and U16644 (N_16644,N_15161,N_15645);
nor U16645 (N_16645,N_15323,N_15640);
xor U16646 (N_16646,N_15631,N_16024);
nor U16647 (N_16647,N_16209,N_15547);
and U16648 (N_16648,N_15248,N_16205);
xnor U16649 (N_16649,N_15113,N_15002);
nor U16650 (N_16650,N_15952,N_16110);
nor U16651 (N_16651,N_15234,N_15655);
nor U16652 (N_16652,N_15889,N_15706);
nand U16653 (N_16653,N_15138,N_15733);
and U16654 (N_16654,N_15244,N_15700);
or U16655 (N_16655,N_15886,N_16100);
nor U16656 (N_16656,N_15026,N_15999);
or U16657 (N_16657,N_15177,N_15065);
or U16658 (N_16658,N_15096,N_15899);
nand U16659 (N_16659,N_15762,N_15851);
and U16660 (N_16660,N_15652,N_15124);
nand U16661 (N_16661,N_15614,N_16144);
xor U16662 (N_16662,N_15877,N_16038);
xnor U16663 (N_16663,N_15892,N_15828);
nand U16664 (N_16664,N_15679,N_15619);
nor U16665 (N_16665,N_15283,N_15457);
xnor U16666 (N_16666,N_15667,N_15224);
nand U16667 (N_16667,N_16130,N_15653);
nand U16668 (N_16668,N_15205,N_15222);
and U16669 (N_16669,N_15460,N_15488);
and U16670 (N_16670,N_15859,N_15230);
nor U16671 (N_16671,N_15620,N_15672);
nor U16672 (N_16672,N_16185,N_15514);
nand U16673 (N_16673,N_15948,N_15678);
nand U16674 (N_16674,N_15980,N_15352);
xnor U16675 (N_16675,N_15883,N_15144);
or U16676 (N_16676,N_15171,N_15918);
nand U16677 (N_16677,N_15424,N_15191);
nand U16678 (N_16678,N_15593,N_15012);
nand U16679 (N_16679,N_15743,N_15606);
or U16680 (N_16680,N_16241,N_15805);
and U16681 (N_16681,N_15129,N_16031);
nor U16682 (N_16682,N_15771,N_15723);
and U16683 (N_16683,N_15011,N_15400);
nand U16684 (N_16684,N_15701,N_15994);
and U16685 (N_16685,N_15407,N_15929);
nand U16686 (N_16686,N_15069,N_15303);
or U16687 (N_16687,N_15676,N_16036);
xor U16688 (N_16688,N_15359,N_15295);
nand U16689 (N_16689,N_15486,N_15092);
or U16690 (N_16690,N_15425,N_15736);
nand U16691 (N_16691,N_15276,N_16128);
and U16692 (N_16692,N_16227,N_15903);
nor U16693 (N_16693,N_15159,N_15045);
and U16694 (N_16694,N_15541,N_15991);
nor U16695 (N_16695,N_15133,N_15416);
and U16696 (N_16696,N_15968,N_16117);
or U16697 (N_16697,N_15333,N_15597);
xor U16698 (N_16698,N_15118,N_15090);
xor U16699 (N_16699,N_15237,N_15335);
xor U16700 (N_16700,N_16164,N_15116);
nand U16701 (N_16701,N_15044,N_15739);
nor U16702 (N_16702,N_15880,N_15322);
nor U16703 (N_16703,N_16182,N_15756);
nand U16704 (N_16704,N_15009,N_15334);
nand U16705 (N_16705,N_16118,N_16087);
and U16706 (N_16706,N_15170,N_15043);
nand U16707 (N_16707,N_16124,N_15306);
nor U16708 (N_16708,N_16152,N_15481);
nor U16709 (N_16709,N_15670,N_15862);
xnor U16710 (N_16710,N_16056,N_15219);
nor U16711 (N_16711,N_15945,N_16203);
xor U16712 (N_16712,N_15293,N_15605);
nor U16713 (N_16713,N_15932,N_15022);
nand U16714 (N_16714,N_15780,N_15472);
nor U16715 (N_16715,N_15157,N_15463);
nor U16716 (N_16716,N_16211,N_15613);
or U16717 (N_16717,N_15451,N_15977);
nand U16718 (N_16718,N_15985,N_15154);
or U16719 (N_16719,N_15086,N_15765);
or U16720 (N_16720,N_15989,N_15992);
nand U16721 (N_16721,N_15162,N_16033);
and U16722 (N_16722,N_16026,N_16189);
or U16723 (N_16723,N_15353,N_16192);
nor U16724 (N_16724,N_15209,N_16143);
xnor U16725 (N_16725,N_15642,N_15140);
nor U16726 (N_16726,N_15021,N_15563);
nor U16727 (N_16727,N_15858,N_15686);
and U16728 (N_16728,N_15285,N_15149);
and U16729 (N_16729,N_16043,N_15919);
nand U16730 (N_16730,N_15097,N_15534);
or U16731 (N_16731,N_15752,N_15186);
and U16732 (N_16732,N_16032,N_16114);
and U16733 (N_16733,N_15634,N_16097);
xor U16734 (N_16734,N_15007,N_15003);
nand U16735 (N_16735,N_15632,N_15466);
xnor U16736 (N_16736,N_15627,N_15925);
and U16737 (N_16737,N_15844,N_15607);
or U16738 (N_16738,N_15913,N_15867);
and U16739 (N_16739,N_16055,N_15109);
nand U16740 (N_16740,N_15685,N_15194);
nor U16741 (N_16741,N_16037,N_15785);
xnor U16742 (N_16742,N_15817,N_15720);
nand U16743 (N_16743,N_15650,N_15902);
nor U16744 (N_16744,N_15575,N_15791);
xnor U16745 (N_16745,N_15702,N_15717);
nor U16746 (N_16746,N_15615,N_16188);
nor U16747 (N_16747,N_15076,N_15103);
nor U16748 (N_16748,N_15329,N_15167);
nor U16749 (N_16749,N_15953,N_16059);
and U16750 (N_16750,N_15665,N_15633);
or U16751 (N_16751,N_16140,N_15760);
nor U16752 (N_16752,N_16201,N_16213);
or U16753 (N_16753,N_15775,N_15110);
nand U16754 (N_16754,N_15961,N_16109);
nor U16755 (N_16755,N_15741,N_15825);
or U16756 (N_16756,N_15287,N_15299);
nand U16757 (N_16757,N_15533,N_15972);
nand U16758 (N_16758,N_15134,N_15555);
or U16759 (N_16759,N_15297,N_16000);
and U16760 (N_16760,N_16153,N_15734);
nor U16761 (N_16761,N_15078,N_15426);
nor U16762 (N_16762,N_15826,N_15535);
xnor U16763 (N_16763,N_15818,N_15532);
and U16764 (N_16764,N_15621,N_15576);
nor U16765 (N_16765,N_15214,N_15691);
xor U16766 (N_16766,N_15477,N_15829);
or U16767 (N_16767,N_16075,N_16101);
nand U16768 (N_16768,N_15189,N_15682);
or U16769 (N_16769,N_16025,N_16202);
nor U16770 (N_16770,N_16134,N_16098);
or U16771 (N_16771,N_15521,N_16204);
nor U16772 (N_16772,N_15467,N_15537);
nand U16773 (N_16773,N_15272,N_15750);
nor U16774 (N_16774,N_15185,N_15927);
and U16775 (N_16775,N_15212,N_15088);
nor U16776 (N_16776,N_15900,N_15395);
nand U16777 (N_16777,N_15735,N_16106);
nor U16778 (N_16778,N_15524,N_15569);
and U16779 (N_16779,N_15799,N_15930);
xnor U16780 (N_16780,N_15501,N_15054);
and U16781 (N_16781,N_15271,N_15783);
nor U16782 (N_16782,N_15060,N_15567);
and U16783 (N_16783,N_15223,N_15438);
xor U16784 (N_16784,N_16163,N_15423);
xor U16785 (N_16785,N_15550,N_16028);
nor U16786 (N_16786,N_15456,N_15151);
nand U16787 (N_16787,N_15145,N_16165);
xnor U16788 (N_16788,N_16180,N_15427);
nor U16789 (N_16789,N_15193,N_16045);
nor U16790 (N_16790,N_15708,N_15896);
or U16791 (N_16791,N_15455,N_16131);
xor U16792 (N_16792,N_15908,N_15861);
xor U16793 (N_16793,N_15361,N_16243);
nand U16794 (N_16794,N_16167,N_15215);
or U16795 (N_16795,N_15578,N_16076);
or U16796 (N_16796,N_15966,N_15728);
nor U16797 (N_16797,N_16135,N_15358);
and U16798 (N_16798,N_15005,N_15988);
nand U16799 (N_16799,N_15326,N_15084);
nand U16800 (N_16800,N_15677,N_15759);
nor U16801 (N_16801,N_15745,N_16150);
xor U16802 (N_16802,N_15884,N_15811);
nor U16803 (N_16803,N_15587,N_15832);
and U16804 (N_16804,N_15461,N_15367);
nor U16805 (N_16805,N_15332,N_15835);
nor U16806 (N_16806,N_15526,N_15690);
nor U16807 (N_16807,N_15479,N_16133);
or U16808 (N_16808,N_15517,N_15399);
and U16809 (N_16809,N_15325,N_15570);
nor U16810 (N_16810,N_15121,N_16044);
or U16811 (N_16811,N_15150,N_15869);
xor U16812 (N_16812,N_15513,N_15439);
nor U16813 (N_16813,N_15610,N_15063);
xor U16814 (N_16814,N_15668,N_15025);
nand U16815 (N_16815,N_16186,N_15074);
nor U16816 (N_16816,N_15496,N_16002);
nor U16817 (N_16817,N_16077,N_16196);
xnor U16818 (N_16818,N_15979,N_16238);
or U16819 (N_16819,N_15236,N_16136);
xnor U16820 (N_16820,N_15774,N_15174);
or U16821 (N_16821,N_15944,N_15198);
xnor U16822 (N_16822,N_15941,N_16215);
nor U16823 (N_16823,N_15549,N_15372);
xnor U16824 (N_16824,N_16050,N_15797);
nor U16825 (N_16825,N_15316,N_15911);
and U16826 (N_16826,N_15716,N_15047);
nor U16827 (N_16827,N_15275,N_15540);
and U16828 (N_16828,N_16132,N_15147);
or U16829 (N_16829,N_16122,N_15689);
nand U16830 (N_16830,N_16176,N_15070);
nand U16831 (N_16831,N_15073,N_16057);
nor U16832 (N_16832,N_15168,N_15796);
or U16833 (N_16833,N_15530,N_15300);
nor U16834 (N_16834,N_16066,N_16175);
and U16835 (N_16835,N_15141,N_15568);
nor U16836 (N_16836,N_15571,N_15898);
xor U16837 (N_16837,N_15566,N_15357);
nor U16838 (N_16838,N_15807,N_15338);
nand U16839 (N_16839,N_15364,N_15581);
nor U16840 (N_16840,N_15922,N_16216);
and U16841 (N_16841,N_15983,N_15611);
xnor U16842 (N_16842,N_15056,N_15349);
or U16843 (N_16843,N_16104,N_15974);
and U16844 (N_16844,N_15231,N_15374);
and U16845 (N_16845,N_16245,N_15837);
xnor U16846 (N_16846,N_15346,N_15527);
and U16847 (N_16847,N_15573,N_15430);
xor U16848 (N_16848,N_16239,N_16091);
nand U16849 (N_16849,N_15318,N_15830);
or U16850 (N_16850,N_15148,N_15923);
nor U16851 (N_16851,N_15693,N_15034);
or U16852 (N_16852,N_15401,N_16174);
and U16853 (N_16853,N_15017,N_15751);
nand U16854 (N_16854,N_15262,N_15142);
nand U16855 (N_16855,N_15583,N_16019);
xor U16856 (N_16856,N_15001,N_16236);
and U16857 (N_16857,N_15314,N_15910);
and U16858 (N_16858,N_15127,N_16008);
or U16859 (N_16859,N_16113,N_15758);
nand U16860 (N_16860,N_15217,N_15618);
xor U16861 (N_16861,N_16014,N_16116);
xor U16862 (N_16862,N_15163,N_15629);
or U16863 (N_16863,N_15754,N_15033);
or U16864 (N_16864,N_15434,N_15840);
or U16865 (N_16865,N_15277,N_15827);
xnor U16866 (N_16866,N_15251,N_15942);
xnor U16867 (N_16867,N_16137,N_15590);
xor U16868 (N_16868,N_15712,N_15315);
nand U16869 (N_16869,N_16208,N_15396);
or U16870 (N_16870,N_15624,N_15281);
and U16871 (N_16871,N_16099,N_15703);
and U16872 (N_16872,N_16228,N_15777);
xor U16873 (N_16873,N_15024,N_15397);
and U16874 (N_16874,N_15935,N_15304);
nor U16875 (N_16875,N_15062,N_15458);
nand U16876 (N_16876,N_15299,N_16175);
xnor U16877 (N_16877,N_15464,N_15406);
xnor U16878 (N_16878,N_16193,N_16099);
nor U16879 (N_16879,N_16097,N_16001);
xor U16880 (N_16880,N_15064,N_15366);
nor U16881 (N_16881,N_15969,N_15865);
xor U16882 (N_16882,N_15312,N_15923);
and U16883 (N_16883,N_15171,N_15187);
and U16884 (N_16884,N_15284,N_15633);
and U16885 (N_16885,N_15929,N_15544);
nand U16886 (N_16886,N_16074,N_15295);
nand U16887 (N_16887,N_16125,N_15732);
nor U16888 (N_16888,N_15474,N_16096);
nand U16889 (N_16889,N_16228,N_15742);
nand U16890 (N_16890,N_16205,N_15381);
xor U16891 (N_16891,N_15015,N_15242);
xnor U16892 (N_16892,N_15740,N_15782);
xnor U16893 (N_16893,N_15146,N_15241);
or U16894 (N_16894,N_16176,N_15646);
nor U16895 (N_16895,N_16116,N_15471);
nor U16896 (N_16896,N_15642,N_15428);
and U16897 (N_16897,N_16079,N_15683);
nor U16898 (N_16898,N_15896,N_15147);
and U16899 (N_16899,N_15676,N_15197);
nor U16900 (N_16900,N_15102,N_15247);
nand U16901 (N_16901,N_15112,N_16177);
nor U16902 (N_16902,N_15647,N_15712);
xor U16903 (N_16903,N_16080,N_15057);
nor U16904 (N_16904,N_15083,N_15898);
nand U16905 (N_16905,N_15418,N_16010);
nor U16906 (N_16906,N_15417,N_15665);
nor U16907 (N_16907,N_15310,N_16097);
and U16908 (N_16908,N_15408,N_15452);
nor U16909 (N_16909,N_16192,N_15993);
and U16910 (N_16910,N_15133,N_15362);
and U16911 (N_16911,N_15334,N_16223);
nand U16912 (N_16912,N_16190,N_15920);
and U16913 (N_16913,N_15451,N_15928);
or U16914 (N_16914,N_15060,N_15169);
nand U16915 (N_16915,N_16039,N_15032);
or U16916 (N_16916,N_16038,N_15105);
and U16917 (N_16917,N_15800,N_15333);
and U16918 (N_16918,N_15752,N_15757);
and U16919 (N_16919,N_15941,N_15222);
xnor U16920 (N_16920,N_15109,N_16108);
nor U16921 (N_16921,N_15241,N_15036);
xor U16922 (N_16922,N_15294,N_15513);
and U16923 (N_16923,N_15153,N_16211);
or U16924 (N_16924,N_15911,N_15409);
or U16925 (N_16925,N_16197,N_15019);
and U16926 (N_16926,N_16058,N_15887);
nand U16927 (N_16927,N_15943,N_15450);
xor U16928 (N_16928,N_15790,N_15332);
or U16929 (N_16929,N_15900,N_15328);
or U16930 (N_16930,N_15136,N_15683);
nor U16931 (N_16931,N_16171,N_15325);
nand U16932 (N_16932,N_15712,N_15555);
or U16933 (N_16933,N_15852,N_15184);
and U16934 (N_16934,N_15028,N_15499);
xnor U16935 (N_16935,N_15733,N_15309);
and U16936 (N_16936,N_15685,N_16148);
nand U16937 (N_16937,N_15877,N_15476);
and U16938 (N_16938,N_15175,N_15299);
nor U16939 (N_16939,N_16113,N_15407);
xnor U16940 (N_16940,N_16040,N_15598);
and U16941 (N_16941,N_15573,N_15553);
nand U16942 (N_16942,N_15671,N_15165);
xor U16943 (N_16943,N_15412,N_16000);
or U16944 (N_16944,N_15172,N_15771);
nor U16945 (N_16945,N_16148,N_15158);
nor U16946 (N_16946,N_15077,N_16201);
or U16947 (N_16947,N_15840,N_16080);
and U16948 (N_16948,N_16024,N_15812);
nand U16949 (N_16949,N_15745,N_16077);
nor U16950 (N_16950,N_15824,N_15786);
nor U16951 (N_16951,N_15412,N_15258);
or U16952 (N_16952,N_15703,N_15792);
xor U16953 (N_16953,N_15569,N_15827);
nor U16954 (N_16954,N_15845,N_15797);
and U16955 (N_16955,N_16236,N_16229);
and U16956 (N_16956,N_15142,N_15322);
nor U16957 (N_16957,N_15746,N_15669);
nand U16958 (N_16958,N_15742,N_16047);
xnor U16959 (N_16959,N_15691,N_15080);
or U16960 (N_16960,N_15411,N_16097);
xnor U16961 (N_16961,N_15639,N_16185);
and U16962 (N_16962,N_15207,N_16204);
and U16963 (N_16963,N_15213,N_15693);
nand U16964 (N_16964,N_15852,N_15605);
nor U16965 (N_16965,N_15982,N_16185);
xnor U16966 (N_16966,N_16191,N_16208);
nand U16967 (N_16967,N_15002,N_15464);
nand U16968 (N_16968,N_15195,N_15135);
nor U16969 (N_16969,N_15634,N_15128);
nor U16970 (N_16970,N_15314,N_15567);
nand U16971 (N_16971,N_15245,N_15584);
nor U16972 (N_16972,N_15277,N_15234);
xor U16973 (N_16973,N_15692,N_15368);
and U16974 (N_16974,N_15881,N_15628);
nor U16975 (N_16975,N_15030,N_15828);
or U16976 (N_16976,N_15429,N_15982);
or U16977 (N_16977,N_15567,N_15742);
nand U16978 (N_16978,N_15666,N_15955);
and U16979 (N_16979,N_15873,N_15597);
and U16980 (N_16980,N_16015,N_15629);
nand U16981 (N_16981,N_15690,N_15661);
nor U16982 (N_16982,N_16132,N_15314);
nor U16983 (N_16983,N_15365,N_16241);
or U16984 (N_16984,N_16053,N_15740);
xor U16985 (N_16985,N_15482,N_16037);
xor U16986 (N_16986,N_15565,N_15972);
xor U16987 (N_16987,N_15154,N_15780);
nand U16988 (N_16988,N_15106,N_15512);
nor U16989 (N_16989,N_15860,N_15910);
and U16990 (N_16990,N_15287,N_15915);
or U16991 (N_16991,N_16141,N_15343);
nand U16992 (N_16992,N_16048,N_15695);
or U16993 (N_16993,N_16103,N_16095);
and U16994 (N_16994,N_16080,N_16143);
or U16995 (N_16995,N_15730,N_15142);
and U16996 (N_16996,N_15037,N_15959);
and U16997 (N_16997,N_15503,N_15960);
nor U16998 (N_16998,N_15959,N_15520);
nor U16999 (N_16999,N_16227,N_15373);
nand U17000 (N_17000,N_15996,N_15151);
nand U17001 (N_17001,N_15634,N_15905);
nand U17002 (N_17002,N_16121,N_16023);
nand U17003 (N_17003,N_16125,N_15480);
nor U17004 (N_17004,N_15982,N_15498);
xnor U17005 (N_17005,N_15336,N_15813);
and U17006 (N_17006,N_15589,N_16043);
nand U17007 (N_17007,N_15384,N_15486);
nor U17008 (N_17008,N_15610,N_15555);
xor U17009 (N_17009,N_15428,N_15462);
and U17010 (N_17010,N_16099,N_16022);
or U17011 (N_17011,N_15450,N_15840);
or U17012 (N_17012,N_15236,N_16119);
xor U17013 (N_17013,N_16117,N_16219);
nor U17014 (N_17014,N_15736,N_16206);
xnor U17015 (N_17015,N_15248,N_15903);
nand U17016 (N_17016,N_15497,N_15347);
and U17017 (N_17017,N_15192,N_16213);
nor U17018 (N_17018,N_15123,N_15483);
or U17019 (N_17019,N_15489,N_15384);
nor U17020 (N_17020,N_15554,N_15575);
and U17021 (N_17021,N_16187,N_15090);
or U17022 (N_17022,N_15927,N_15003);
xnor U17023 (N_17023,N_16013,N_16098);
or U17024 (N_17024,N_16114,N_15669);
nand U17025 (N_17025,N_15005,N_15221);
or U17026 (N_17026,N_15848,N_16070);
xnor U17027 (N_17027,N_15279,N_15028);
xor U17028 (N_17028,N_16208,N_15635);
xnor U17029 (N_17029,N_15913,N_15835);
nor U17030 (N_17030,N_15809,N_15922);
and U17031 (N_17031,N_15335,N_15530);
nor U17032 (N_17032,N_15891,N_15761);
nor U17033 (N_17033,N_15397,N_15207);
nand U17034 (N_17034,N_15139,N_15678);
xnor U17035 (N_17035,N_15082,N_15081);
xnor U17036 (N_17036,N_15469,N_15561);
xnor U17037 (N_17037,N_15575,N_15060);
nor U17038 (N_17038,N_15008,N_15913);
xnor U17039 (N_17039,N_15813,N_16079);
nand U17040 (N_17040,N_15805,N_15943);
nor U17041 (N_17041,N_15162,N_15311);
and U17042 (N_17042,N_15690,N_15089);
xnor U17043 (N_17043,N_16225,N_15615);
xor U17044 (N_17044,N_15250,N_15772);
nor U17045 (N_17045,N_15989,N_15482);
and U17046 (N_17046,N_15939,N_16075);
or U17047 (N_17047,N_15583,N_15060);
xor U17048 (N_17048,N_15249,N_15078);
or U17049 (N_17049,N_16223,N_15091);
and U17050 (N_17050,N_15324,N_16222);
or U17051 (N_17051,N_15181,N_15054);
nor U17052 (N_17052,N_15204,N_16192);
or U17053 (N_17053,N_15463,N_16218);
and U17054 (N_17054,N_16202,N_16091);
and U17055 (N_17055,N_16092,N_15207);
xor U17056 (N_17056,N_15726,N_15434);
nor U17057 (N_17057,N_15866,N_15100);
nor U17058 (N_17058,N_15251,N_16068);
and U17059 (N_17059,N_15078,N_15912);
nor U17060 (N_17060,N_15448,N_16152);
nor U17061 (N_17061,N_15738,N_15365);
nand U17062 (N_17062,N_16229,N_15111);
nand U17063 (N_17063,N_15864,N_15996);
and U17064 (N_17064,N_15327,N_16165);
nor U17065 (N_17065,N_15755,N_15159);
xor U17066 (N_17066,N_15360,N_15824);
xnor U17067 (N_17067,N_15304,N_15875);
nor U17068 (N_17068,N_15062,N_15630);
and U17069 (N_17069,N_15224,N_15750);
xor U17070 (N_17070,N_15639,N_15905);
nand U17071 (N_17071,N_15857,N_15870);
or U17072 (N_17072,N_15561,N_15640);
or U17073 (N_17073,N_15388,N_16038);
xor U17074 (N_17074,N_16224,N_15147);
or U17075 (N_17075,N_16142,N_15623);
and U17076 (N_17076,N_15099,N_15524);
nor U17077 (N_17077,N_15236,N_15714);
xnor U17078 (N_17078,N_15018,N_15687);
xnor U17079 (N_17079,N_15947,N_15577);
nor U17080 (N_17080,N_15376,N_15314);
nor U17081 (N_17081,N_16009,N_15760);
xor U17082 (N_17082,N_15538,N_16223);
nor U17083 (N_17083,N_15102,N_15622);
and U17084 (N_17084,N_15318,N_15585);
xnor U17085 (N_17085,N_15174,N_16170);
and U17086 (N_17086,N_16095,N_16006);
and U17087 (N_17087,N_15915,N_15615);
nor U17088 (N_17088,N_15213,N_15668);
nor U17089 (N_17089,N_15468,N_15286);
xor U17090 (N_17090,N_16057,N_15339);
or U17091 (N_17091,N_15602,N_16170);
nor U17092 (N_17092,N_15386,N_15128);
xnor U17093 (N_17093,N_15881,N_15197);
nand U17094 (N_17094,N_15037,N_15767);
nor U17095 (N_17095,N_15154,N_15471);
xor U17096 (N_17096,N_15961,N_16062);
or U17097 (N_17097,N_15487,N_16002);
nand U17098 (N_17098,N_15278,N_15583);
or U17099 (N_17099,N_15754,N_15056);
or U17100 (N_17100,N_15987,N_16153);
and U17101 (N_17101,N_15068,N_16062);
nand U17102 (N_17102,N_15190,N_15512);
xor U17103 (N_17103,N_15390,N_15596);
and U17104 (N_17104,N_16096,N_15273);
nand U17105 (N_17105,N_15747,N_15390);
nor U17106 (N_17106,N_15799,N_15104);
xor U17107 (N_17107,N_15587,N_15305);
and U17108 (N_17108,N_15423,N_15878);
and U17109 (N_17109,N_15943,N_15716);
nand U17110 (N_17110,N_15608,N_15177);
nor U17111 (N_17111,N_15935,N_15432);
xor U17112 (N_17112,N_15002,N_15786);
nand U17113 (N_17113,N_15216,N_15388);
xor U17114 (N_17114,N_15539,N_16179);
xnor U17115 (N_17115,N_16089,N_15942);
xnor U17116 (N_17116,N_15332,N_15704);
nor U17117 (N_17117,N_15269,N_15171);
nor U17118 (N_17118,N_15440,N_15905);
xor U17119 (N_17119,N_16073,N_15753);
xnor U17120 (N_17120,N_15951,N_15805);
nor U17121 (N_17121,N_15694,N_15855);
xnor U17122 (N_17122,N_15652,N_15921);
or U17123 (N_17123,N_16167,N_15236);
or U17124 (N_17124,N_15977,N_16127);
nor U17125 (N_17125,N_15447,N_15664);
nor U17126 (N_17126,N_15940,N_15478);
xnor U17127 (N_17127,N_15162,N_15010);
nand U17128 (N_17128,N_15230,N_15475);
or U17129 (N_17129,N_15041,N_15018);
xor U17130 (N_17130,N_15078,N_15647);
or U17131 (N_17131,N_15411,N_15033);
nand U17132 (N_17132,N_15718,N_15162);
nor U17133 (N_17133,N_15893,N_15480);
or U17134 (N_17134,N_15409,N_15870);
or U17135 (N_17135,N_16167,N_15675);
nand U17136 (N_17136,N_15724,N_15518);
or U17137 (N_17137,N_15592,N_15374);
xor U17138 (N_17138,N_15519,N_15132);
and U17139 (N_17139,N_15479,N_15144);
or U17140 (N_17140,N_15103,N_15665);
xor U17141 (N_17141,N_15718,N_16225);
nor U17142 (N_17142,N_15836,N_15787);
nand U17143 (N_17143,N_15089,N_15220);
nor U17144 (N_17144,N_15346,N_16208);
nor U17145 (N_17145,N_15702,N_15549);
nand U17146 (N_17146,N_15587,N_15704);
and U17147 (N_17147,N_16145,N_15394);
xnor U17148 (N_17148,N_15592,N_15006);
and U17149 (N_17149,N_15609,N_15229);
nor U17150 (N_17150,N_15691,N_15796);
nand U17151 (N_17151,N_16240,N_16045);
nand U17152 (N_17152,N_15087,N_15794);
or U17153 (N_17153,N_15495,N_15172);
and U17154 (N_17154,N_15011,N_15631);
nand U17155 (N_17155,N_16093,N_16044);
nor U17156 (N_17156,N_15075,N_15135);
nor U17157 (N_17157,N_15548,N_15292);
or U17158 (N_17158,N_15536,N_16055);
or U17159 (N_17159,N_15655,N_15866);
nand U17160 (N_17160,N_15195,N_15369);
nor U17161 (N_17161,N_15120,N_15857);
or U17162 (N_17162,N_15384,N_15217);
or U17163 (N_17163,N_15599,N_15151);
or U17164 (N_17164,N_16193,N_15922);
and U17165 (N_17165,N_15882,N_15403);
xnor U17166 (N_17166,N_15317,N_15344);
or U17167 (N_17167,N_15575,N_16119);
nand U17168 (N_17168,N_16035,N_15191);
xor U17169 (N_17169,N_15453,N_15544);
nand U17170 (N_17170,N_15658,N_15968);
or U17171 (N_17171,N_16057,N_15958);
nor U17172 (N_17172,N_16227,N_15000);
nor U17173 (N_17173,N_15188,N_15732);
or U17174 (N_17174,N_16222,N_15225);
nand U17175 (N_17175,N_15720,N_15178);
and U17176 (N_17176,N_15399,N_15487);
or U17177 (N_17177,N_15025,N_15171);
and U17178 (N_17178,N_15553,N_16005);
or U17179 (N_17179,N_16154,N_15064);
nor U17180 (N_17180,N_16107,N_15735);
and U17181 (N_17181,N_15666,N_15333);
and U17182 (N_17182,N_16038,N_15316);
and U17183 (N_17183,N_15557,N_15044);
or U17184 (N_17184,N_15971,N_16086);
nand U17185 (N_17185,N_15715,N_15438);
or U17186 (N_17186,N_15380,N_15966);
nor U17187 (N_17187,N_16158,N_15718);
and U17188 (N_17188,N_16212,N_15405);
and U17189 (N_17189,N_16156,N_15295);
xnor U17190 (N_17190,N_16162,N_16186);
nor U17191 (N_17191,N_15142,N_15988);
and U17192 (N_17192,N_15587,N_15237);
nand U17193 (N_17193,N_15883,N_15456);
nand U17194 (N_17194,N_15087,N_15123);
nor U17195 (N_17195,N_16233,N_15484);
nor U17196 (N_17196,N_15307,N_15259);
xor U17197 (N_17197,N_15425,N_15189);
nor U17198 (N_17198,N_15555,N_15058);
nor U17199 (N_17199,N_15511,N_15910);
or U17200 (N_17200,N_16191,N_15102);
xnor U17201 (N_17201,N_15267,N_15141);
xor U17202 (N_17202,N_15904,N_16216);
or U17203 (N_17203,N_15960,N_15560);
nand U17204 (N_17204,N_15296,N_15273);
or U17205 (N_17205,N_15178,N_16022);
or U17206 (N_17206,N_15373,N_15740);
xnor U17207 (N_17207,N_15116,N_15995);
or U17208 (N_17208,N_15068,N_15947);
xnor U17209 (N_17209,N_15706,N_15805);
nand U17210 (N_17210,N_16061,N_16133);
nand U17211 (N_17211,N_16124,N_15393);
nor U17212 (N_17212,N_16244,N_15678);
and U17213 (N_17213,N_15791,N_15668);
and U17214 (N_17214,N_16224,N_15378);
nand U17215 (N_17215,N_15644,N_15852);
and U17216 (N_17216,N_16170,N_15138);
and U17217 (N_17217,N_15485,N_16071);
or U17218 (N_17218,N_15666,N_15422);
or U17219 (N_17219,N_16019,N_15242);
or U17220 (N_17220,N_15821,N_16109);
or U17221 (N_17221,N_15343,N_15717);
and U17222 (N_17222,N_15150,N_16042);
nand U17223 (N_17223,N_15852,N_15429);
xor U17224 (N_17224,N_15821,N_16039);
xnor U17225 (N_17225,N_15220,N_15946);
nor U17226 (N_17226,N_16064,N_15348);
nor U17227 (N_17227,N_15499,N_15463);
and U17228 (N_17228,N_15132,N_16201);
nor U17229 (N_17229,N_15677,N_15214);
nor U17230 (N_17230,N_15133,N_15545);
xor U17231 (N_17231,N_15569,N_15795);
nand U17232 (N_17232,N_15218,N_15391);
or U17233 (N_17233,N_15996,N_15157);
and U17234 (N_17234,N_15510,N_15972);
or U17235 (N_17235,N_16142,N_15959);
xor U17236 (N_17236,N_15963,N_16027);
xnor U17237 (N_17237,N_15711,N_15528);
and U17238 (N_17238,N_16082,N_15839);
nand U17239 (N_17239,N_15765,N_15408);
and U17240 (N_17240,N_15656,N_15704);
or U17241 (N_17241,N_15283,N_16197);
nor U17242 (N_17242,N_15608,N_15385);
nor U17243 (N_17243,N_16019,N_15876);
nand U17244 (N_17244,N_15445,N_15563);
nor U17245 (N_17245,N_16055,N_15898);
or U17246 (N_17246,N_15574,N_15107);
nand U17247 (N_17247,N_15566,N_15157);
nor U17248 (N_17248,N_15733,N_16101);
nor U17249 (N_17249,N_16030,N_15493);
and U17250 (N_17250,N_15185,N_15650);
nor U17251 (N_17251,N_16136,N_15363);
and U17252 (N_17252,N_15859,N_15056);
nor U17253 (N_17253,N_15168,N_16212);
nand U17254 (N_17254,N_15597,N_15639);
xor U17255 (N_17255,N_15682,N_16171);
xnor U17256 (N_17256,N_16049,N_16159);
nand U17257 (N_17257,N_15492,N_15118);
nor U17258 (N_17258,N_16205,N_15823);
nand U17259 (N_17259,N_15623,N_15237);
xor U17260 (N_17260,N_15431,N_15796);
nor U17261 (N_17261,N_16143,N_15989);
and U17262 (N_17262,N_15043,N_15361);
xor U17263 (N_17263,N_15496,N_15335);
nand U17264 (N_17264,N_15199,N_15778);
or U17265 (N_17265,N_15327,N_16120);
nand U17266 (N_17266,N_15543,N_15945);
nor U17267 (N_17267,N_15163,N_15607);
xnor U17268 (N_17268,N_16047,N_15321);
nand U17269 (N_17269,N_15468,N_15512);
xnor U17270 (N_17270,N_15697,N_16146);
xor U17271 (N_17271,N_16007,N_15177);
and U17272 (N_17272,N_15947,N_15478);
nor U17273 (N_17273,N_15477,N_16049);
and U17274 (N_17274,N_15120,N_16115);
nor U17275 (N_17275,N_15600,N_15510);
and U17276 (N_17276,N_15321,N_15879);
nor U17277 (N_17277,N_15758,N_15278);
and U17278 (N_17278,N_15404,N_15366);
xnor U17279 (N_17279,N_15998,N_15508);
and U17280 (N_17280,N_15669,N_15367);
xor U17281 (N_17281,N_15381,N_16232);
or U17282 (N_17282,N_15881,N_15243);
nor U17283 (N_17283,N_16147,N_15370);
xor U17284 (N_17284,N_15366,N_15855);
or U17285 (N_17285,N_15079,N_15308);
or U17286 (N_17286,N_15696,N_15144);
nand U17287 (N_17287,N_15868,N_15583);
nand U17288 (N_17288,N_15945,N_16055);
nor U17289 (N_17289,N_15299,N_16128);
and U17290 (N_17290,N_15070,N_15283);
xnor U17291 (N_17291,N_15760,N_15884);
nor U17292 (N_17292,N_15678,N_15441);
xnor U17293 (N_17293,N_15622,N_15159);
or U17294 (N_17294,N_16033,N_16208);
or U17295 (N_17295,N_15473,N_15064);
xor U17296 (N_17296,N_15126,N_15530);
or U17297 (N_17297,N_16001,N_15636);
nor U17298 (N_17298,N_15279,N_15175);
nor U17299 (N_17299,N_15168,N_15227);
and U17300 (N_17300,N_15975,N_15788);
and U17301 (N_17301,N_16117,N_15037);
and U17302 (N_17302,N_15364,N_16034);
nor U17303 (N_17303,N_15101,N_15586);
nand U17304 (N_17304,N_15801,N_15878);
nor U17305 (N_17305,N_15174,N_15679);
and U17306 (N_17306,N_15928,N_15063);
nand U17307 (N_17307,N_15543,N_15322);
nor U17308 (N_17308,N_16172,N_15693);
or U17309 (N_17309,N_15472,N_15704);
nand U17310 (N_17310,N_15966,N_15598);
nor U17311 (N_17311,N_15611,N_15264);
nor U17312 (N_17312,N_15618,N_15429);
xor U17313 (N_17313,N_15590,N_15862);
nand U17314 (N_17314,N_15677,N_15384);
nor U17315 (N_17315,N_15617,N_15370);
nand U17316 (N_17316,N_15933,N_15068);
xor U17317 (N_17317,N_15616,N_15230);
nor U17318 (N_17318,N_15088,N_15856);
or U17319 (N_17319,N_16154,N_15881);
xor U17320 (N_17320,N_15140,N_15024);
nor U17321 (N_17321,N_15082,N_15721);
and U17322 (N_17322,N_15724,N_15035);
nand U17323 (N_17323,N_16162,N_15533);
nor U17324 (N_17324,N_15928,N_15136);
and U17325 (N_17325,N_15830,N_15047);
nor U17326 (N_17326,N_15525,N_15083);
nor U17327 (N_17327,N_15103,N_16198);
nand U17328 (N_17328,N_15383,N_15157);
or U17329 (N_17329,N_15355,N_15223);
or U17330 (N_17330,N_15526,N_15168);
and U17331 (N_17331,N_15972,N_15091);
nor U17332 (N_17332,N_16114,N_15286);
xor U17333 (N_17333,N_15137,N_15011);
nand U17334 (N_17334,N_15461,N_15420);
xor U17335 (N_17335,N_15066,N_16073);
or U17336 (N_17336,N_15845,N_15893);
and U17337 (N_17337,N_15218,N_15925);
nor U17338 (N_17338,N_15192,N_15812);
nand U17339 (N_17339,N_15451,N_15070);
xor U17340 (N_17340,N_15645,N_15928);
or U17341 (N_17341,N_15176,N_15871);
and U17342 (N_17342,N_15535,N_16237);
nand U17343 (N_17343,N_15715,N_15958);
nor U17344 (N_17344,N_15280,N_15426);
and U17345 (N_17345,N_16232,N_15571);
nor U17346 (N_17346,N_15158,N_15035);
nor U17347 (N_17347,N_15672,N_15150);
nand U17348 (N_17348,N_15424,N_15147);
and U17349 (N_17349,N_15848,N_16063);
or U17350 (N_17350,N_15695,N_15337);
or U17351 (N_17351,N_16004,N_16100);
nor U17352 (N_17352,N_15689,N_16099);
xor U17353 (N_17353,N_15535,N_16027);
or U17354 (N_17354,N_15928,N_15139);
and U17355 (N_17355,N_15178,N_15752);
nor U17356 (N_17356,N_15824,N_15873);
nand U17357 (N_17357,N_15088,N_16073);
xor U17358 (N_17358,N_15078,N_16206);
or U17359 (N_17359,N_15524,N_15674);
nand U17360 (N_17360,N_15380,N_15351);
and U17361 (N_17361,N_15182,N_15910);
nor U17362 (N_17362,N_15434,N_16192);
nor U17363 (N_17363,N_15825,N_15756);
nand U17364 (N_17364,N_15370,N_15421);
xnor U17365 (N_17365,N_16184,N_16131);
or U17366 (N_17366,N_15267,N_16248);
xnor U17367 (N_17367,N_15380,N_16096);
and U17368 (N_17368,N_15729,N_15745);
nand U17369 (N_17369,N_16177,N_15923);
and U17370 (N_17370,N_15743,N_15496);
nand U17371 (N_17371,N_15433,N_15875);
and U17372 (N_17372,N_15101,N_15408);
and U17373 (N_17373,N_15803,N_15594);
xor U17374 (N_17374,N_15758,N_15732);
nand U17375 (N_17375,N_16114,N_15240);
or U17376 (N_17376,N_15583,N_15688);
nand U17377 (N_17377,N_16211,N_15160);
xor U17378 (N_17378,N_15652,N_15605);
and U17379 (N_17379,N_16127,N_15354);
nand U17380 (N_17380,N_16161,N_15433);
or U17381 (N_17381,N_16134,N_15980);
or U17382 (N_17382,N_15539,N_15533);
or U17383 (N_17383,N_15169,N_15607);
nand U17384 (N_17384,N_16189,N_15989);
or U17385 (N_17385,N_16025,N_15218);
xnor U17386 (N_17386,N_15154,N_15284);
nor U17387 (N_17387,N_15234,N_15667);
xor U17388 (N_17388,N_15066,N_16127);
nand U17389 (N_17389,N_15757,N_15690);
nor U17390 (N_17390,N_15787,N_15463);
xnor U17391 (N_17391,N_15911,N_15220);
xnor U17392 (N_17392,N_15090,N_15031);
nand U17393 (N_17393,N_16233,N_15902);
or U17394 (N_17394,N_15519,N_15007);
and U17395 (N_17395,N_15387,N_15109);
or U17396 (N_17396,N_15443,N_15041);
xnor U17397 (N_17397,N_15723,N_15986);
and U17398 (N_17398,N_15637,N_15817);
xor U17399 (N_17399,N_15687,N_15813);
xnor U17400 (N_17400,N_15143,N_15631);
nor U17401 (N_17401,N_15614,N_15687);
or U17402 (N_17402,N_16151,N_15350);
xnor U17403 (N_17403,N_16051,N_15073);
and U17404 (N_17404,N_16122,N_15181);
nor U17405 (N_17405,N_15149,N_15170);
or U17406 (N_17406,N_16177,N_15267);
or U17407 (N_17407,N_15205,N_15308);
nor U17408 (N_17408,N_15731,N_15502);
xor U17409 (N_17409,N_15325,N_16214);
nor U17410 (N_17410,N_16223,N_15677);
nand U17411 (N_17411,N_15145,N_15245);
nand U17412 (N_17412,N_15436,N_15140);
nor U17413 (N_17413,N_16044,N_15874);
or U17414 (N_17414,N_15160,N_15322);
nor U17415 (N_17415,N_16240,N_15255);
and U17416 (N_17416,N_15630,N_16178);
xor U17417 (N_17417,N_15959,N_16015);
or U17418 (N_17418,N_15009,N_16149);
or U17419 (N_17419,N_15942,N_16009);
xnor U17420 (N_17420,N_15136,N_15531);
and U17421 (N_17421,N_15299,N_16003);
nand U17422 (N_17422,N_15563,N_15108);
or U17423 (N_17423,N_15693,N_15595);
xnor U17424 (N_17424,N_15724,N_16028);
nand U17425 (N_17425,N_15301,N_15880);
or U17426 (N_17426,N_15132,N_16174);
nor U17427 (N_17427,N_15716,N_15726);
nand U17428 (N_17428,N_15373,N_15731);
and U17429 (N_17429,N_15456,N_16019);
nor U17430 (N_17430,N_15286,N_15909);
and U17431 (N_17431,N_15796,N_15962);
xor U17432 (N_17432,N_15460,N_15790);
nor U17433 (N_17433,N_15148,N_15977);
xor U17434 (N_17434,N_16160,N_15717);
nor U17435 (N_17435,N_16194,N_15285);
and U17436 (N_17436,N_15022,N_15045);
nand U17437 (N_17437,N_16108,N_15618);
xor U17438 (N_17438,N_15345,N_15932);
xnor U17439 (N_17439,N_15155,N_16023);
nor U17440 (N_17440,N_15666,N_15730);
xor U17441 (N_17441,N_15528,N_15820);
or U17442 (N_17442,N_15174,N_15978);
nand U17443 (N_17443,N_16135,N_15404);
nand U17444 (N_17444,N_16138,N_15505);
xor U17445 (N_17445,N_15720,N_16193);
and U17446 (N_17446,N_15155,N_15261);
nand U17447 (N_17447,N_15312,N_15332);
nand U17448 (N_17448,N_15402,N_15500);
nor U17449 (N_17449,N_15601,N_15977);
xor U17450 (N_17450,N_16028,N_15093);
and U17451 (N_17451,N_15814,N_15626);
nor U17452 (N_17452,N_15256,N_15873);
nand U17453 (N_17453,N_15305,N_15717);
nor U17454 (N_17454,N_15334,N_15210);
nand U17455 (N_17455,N_15678,N_15583);
and U17456 (N_17456,N_16155,N_15245);
xnor U17457 (N_17457,N_15911,N_15525);
nand U17458 (N_17458,N_16170,N_15792);
and U17459 (N_17459,N_15517,N_15084);
xnor U17460 (N_17460,N_15345,N_16213);
or U17461 (N_17461,N_15854,N_15141);
xor U17462 (N_17462,N_15301,N_15975);
nand U17463 (N_17463,N_15720,N_15813);
xor U17464 (N_17464,N_15466,N_16241);
nor U17465 (N_17465,N_15524,N_15826);
xor U17466 (N_17466,N_15851,N_15376);
nand U17467 (N_17467,N_15221,N_15329);
nand U17468 (N_17468,N_15942,N_15203);
and U17469 (N_17469,N_15686,N_15824);
and U17470 (N_17470,N_16217,N_15425);
xor U17471 (N_17471,N_15015,N_15486);
nor U17472 (N_17472,N_16219,N_16087);
and U17473 (N_17473,N_15510,N_15572);
nor U17474 (N_17474,N_15317,N_15436);
and U17475 (N_17475,N_15668,N_16049);
xnor U17476 (N_17476,N_15456,N_15304);
and U17477 (N_17477,N_15824,N_16043);
and U17478 (N_17478,N_15486,N_15812);
nor U17479 (N_17479,N_15879,N_15615);
nor U17480 (N_17480,N_15868,N_15627);
xnor U17481 (N_17481,N_15270,N_15407);
xnor U17482 (N_17482,N_15659,N_15295);
or U17483 (N_17483,N_15494,N_15256);
and U17484 (N_17484,N_15291,N_15635);
nand U17485 (N_17485,N_15138,N_15643);
and U17486 (N_17486,N_15043,N_15974);
and U17487 (N_17487,N_15477,N_15649);
xor U17488 (N_17488,N_16107,N_15101);
xnor U17489 (N_17489,N_15953,N_15843);
xor U17490 (N_17490,N_15934,N_15201);
or U17491 (N_17491,N_15066,N_15346);
xor U17492 (N_17492,N_15161,N_15023);
nor U17493 (N_17493,N_15468,N_15199);
xor U17494 (N_17494,N_16060,N_15145);
nand U17495 (N_17495,N_16238,N_16234);
and U17496 (N_17496,N_15350,N_15879);
or U17497 (N_17497,N_15029,N_15094);
and U17498 (N_17498,N_15415,N_16029);
and U17499 (N_17499,N_15549,N_15404);
xnor U17500 (N_17500,N_16500,N_16336);
and U17501 (N_17501,N_16860,N_17162);
xor U17502 (N_17502,N_16813,N_17237);
nand U17503 (N_17503,N_17338,N_17381);
nand U17504 (N_17504,N_16676,N_16326);
nand U17505 (N_17505,N_16856,N_16266);
xnor U17506 (N_17506,N_17481,N_16779);
nand U17507 (N_17507,N_17291,N_16818);
or U17508 (N_17508,N_16750,N_17475);
nand U17509 (N_17509,N_16299,N_16358);
and U17510 (N_17510,N_16380,N_16342);
and U17511 (N_17511,N_16279,N_16317);
or U17512 (N_17512,N_17358,N_17002);
nand U17513 (N_17513,N_17473,N_16257);
and U17514 (N_17514,N_17422,N_17198);
or U17515 (N_17515,N_16740,N_16271);
nor U17516 (N_17516,N_16654,N_17290);
xnor U17517 (N_17517,N_16822,N_16385);
nand U17518 (N_17518,N_16868,N_16967);
and U17519 (N_17519,N_17455,N_16406);
nand U17520 (N_17520,N_16826,N_17335);
nand U17521 (N_17521,N_16564,N_17313);
or U17522 (N_17522,N_17200,N_16887);
or U17523 (N_17523,N_16855,N_17468);
nand U17524 (N_17524,N_17416,N_17280);
xnor U17525 (N_17525,N_17462,N_16330);
xnor U17526 (N_17526,N_16400,N_16424);
nor U17527 (N_17527,N_17193,N_17220);
nor U17528 (N_17528,N_16394,N_16786);
nand U17529 (N_17529,N_17009,N_16384);
nand U17530 (N_17530,N_16973,N_17165);
and U17531 (N_17531,N_16490,N_16663);
nor U17532 (N_17532,N_16834,N_16777);
nand U17533 (N_17533,N_16691,N_16339);
or U17534 (N_17534,N_16681,N_16802);
nor U17535 (N_17535,N_16450,N_16690);
nor U17536 (N_17536,N_16426,N_16914);
nand U17537 (N_17537,N_16594,N_16667);
or U17538 (N_17538,N_17407,N_16316);
and U17539 (N_17539,N_16412,N_16994);
xor U17540 (N_17540,N_16805,N_16431);
nand U17541 (N_17541,N_17225,N_16946);
or U17542 (N_17542,N_16809,N_17458);
xnor U17543 (N_17543,N_17470,N_16886);
and U17544 (N_17544,N_16929,N_16700);
or U17545 (N_17545,N_16347,N_16391);
nand U17546 (N_17546,N_17418,N_17394);
and U17547 (N_17547,N_16734,N_16482);
nand U17548 (N_17548,N_16747,N_16588);
xor U17549 (N_17549,N_16293,N_16657);
nand U17550 (N_17550,N_16399,N_17234);
nor U17551 (N_17551,N_16884,N_16581);
and U17552 (N_17552,N_16757,N_16679);
and U17553 (N_17553,N_17020,N_17106);
or U17554 (N_17554,N_16540,N_17145);
or U17555 (N_17555,N_17050,N_17054);
nor U17556 (N_17556,N_17460,N_17128);
nor U17557 (N_17557,N_16791,N_16409);
xor U17558 (N_17558,N_17297,N_17464);
and U17559 (N_17559,N_16726,N_16453);
and U17560 (N_17560,N_17070,N_16344);
or U17561 (N_17561,N_16745,N_16814);
nor U17562 (N_17562,N_16961,N_16900);
or U17563 (N_17563,N_16656,N_16495);
nand U17564 (N_17564,N_17021,N_16732);
and U17565 (N_17565,N_16950,N_17385);
xor U17566 (N_17566,N_16720,N_16939);
and U17567 (N_17567,N_16964,N_17122);
and U17568 (N_17568,N_17390,N_16694);
nor U17569 (N_17569,N_16284,N_17393);
nor U17570 (N_17570,N_16986,N_16577);
or U17571 (N_17571,N_17146,N_16639);
nand U17572 (N_17572,N_16638,N_16371);
nand U17573 (N_17573,N_16682,N_16306);
or U17574 (N_17574,N_17449,N_17118);
nand U17575 (N_17575,N_16989,N_16760);
and U17576 (N_17576,N_17041,N_16838);
and U17577 (N_17577,N_17262,N_17180);
xnor U17578 (N_17578,N_16583,N_16922);
and U17579 (N_17579,N_17174,N_17402);
or U17580 (N_17580,N_16554,N_16627);
or U17581 (N_17581,N_16778,N_16932);
nand U17582 (N_17582,N_17014,N_16825);
or U17583 (N_17583,N_17271,N_16658);
nor U17584 (N_17584,N_17346,N_16295);
or U17585 (N_17585,N_16290,N_16811);
or U17586 (N_17586,N_16280,N_16992);
xor U17587 (N_17587,N_16792,N_16551);
and U17588 (N_17588,N_16524,N_16525);
nor U17589 (N_17589,N_17367,N_17497);
and U17590 (N_17590,N_16289,N_17104);
or U17591 (N_17591,N_17484,N_16448);
nand U17592 (N_17592,N_17212,N_16535);
and U17593 (N_17593,N_16442,N_17159);
nand U17594 (N_17594,N_16512,N_16851);
nand U17595 (N_17595,N_17119,N_17436);
or U17596 (N_17596,N_16496,N_16541);
xnor U17597 (N_17597,N_17051,N_16710);
and U17598 (N_17598,N_16959,N_16386);
and U17599 (N_17599,N_17334,N_17044);
xor U17600 (N_17600,N_16530,N_16435);
or U17601 (N_17601,N_17179,N_16800);
and U17602 (N_17602,N_16789,N_16816);
xor U17603 (N_17603,N_16984,N_16373);
and U17604 (N_17604,N_16919,N_17454);
nand U17605 (N_17605,N_17332,N_16985);
and U17606 (N_17606,N_17306,N_17152);
or U17607 (N_17607,N_17081,N_16437);
and U17608 (N_17608,N_16897,N_16416);
and U17609 (N_17609,N_16349,N_16340);
and U17610 (N_17610,N_16931,N_16979);
and U17611 (N_17611,N_16870,N_17448);
nand U17612 (N_17612,N_16841,N_16355);
xnor U17613 (N_17613,N_17176,N_17388);
xor U17614 (N_17614,N_16307,N_16605);
xnor U17615 (N_17615,N_17168,N_17030);
xor U17616 (N_17616,N_16441,N_16763);
and U17617 (N_17617,N_16815,N_17006);
nand U17618 (N_17618,N_17072,N_16458);
nand U17619 (N_17619,N_16606,N_16767);
and U17620 (N_17620,N_16904,N_16546);
and U17621 (N_17621,N_16396,N_16936);
or U17622 (N_17622,N_16276,N_16775);
nand U17623 (N_17623,N_16446,N_17164);
or U17624 (N_17624,N_16624,N_16592);
or U17625 (N_17625,N_16364,N_16930);
xor U17626 (N_17626,N_17192,N_16568);
or U17627 (N_17627,N_16372,N_16534);
and U17628 (N_17628,N_16617,N_16927);
xor U17629 (N_17629,N_17236,N_16623);
nand U17630 (N_17630,N_16480,N_16997);
nor U17631 (N_17631,N_16256,N_17127);
nand U17632 (N_17632,N_17300,N_16762);
xnor U17633 (N_17633,N_16252,N_17078);
or U17634 (N_17634,N_16913,N_17170);
nand U17635 (N_17635,N_16558,N_16701);
and U17636 (N_17636,N_17419,N_17304);
nand U17637 (N_17637,N_16713,N_17115);
nor U17638 (N_17638,N_17148,N_17130);
nor U17639 (N_17639,N_16864,N_17075);
or U17640 (N_17640,N_16596,N_16543);
nand U17641 (N_17641,N_16398,N_16263);
or U17642 (N_17642,N_16951,N_16590);
nand U17643 (N_17643,N_17289,N_17424);
nand U17644 (N_17644,N_16803,N_16502);
or U17645 (N_17645,N_16593,N_17079);
nand U17646 (N_17646,N_17026,N_17292);
xor U17647 (N_17647,N_17429,N_16801);
nand U17648 (N_17648,N_17283,N_17347);
or U17649 (N_17649,N_16839,N_16388);
nand U17650 (N_17650,N_16678,N_16664);
nor U17651 (N_17651,N_16444,N_17032);
nand U17652 (N_17652,N_17109,N_17042);
xnor U17653 (N_17653,N_17379,N_17382);
or U17654 (N_17654,N_17417,N_17161);
or U17655 (N_17655,N_17024,N_17392);
or U17656 (N_17656,N_16675,N_16439);
nor U17657 (N_17657,N_16928,N_17206);
and U17658 (N_17658,N_16589,N_16456);
or U17659 (N_17659,N_17219,N_17296);
nand U17660 (N_17660,N_17033,N_17116);
nand U17661 (N_17661,N_17278,N_17434);
nor U17662 (N_17662,N_17453,N_17154);
nand U17663 (N_17663,N_16683,N_17359);
nor U17664 (N_17664,N_16445,N_17077);
or U17665 (N_17665,N_16473,N_17133);
and U17666 (N_17666,N_17428,N_17195);
xor U17667 (N_17667,N_16275,N_16447);
or U17668 (N_17668,N_16423,N_17275);
or U17669 (N_17669,N_16324,N_16807);
and U17670 (N_17670,N_16796,N_17264);
nor U17671 (N_17671,N_16493,N_16844);
or U17672 (N_17672,N_16924,N_17218);
nor U17673 (N_17673,N_17308,N_16722);
nor U17674 (N_17674,N_17113,N_17076);
or U17675 (N_17675,N_16764,N_17114);
or U17676 (N_17676,N_16689,N_17284);
or U17677 (N_17677,N_16836,N_16718);
xor U17678 (N_17678,N_16487,N_17285);
or U17679 (N_17679,N_16335,N_16794);
xnor U17680 (N_17680,N_17047,N_17025);
nor U17681 (N_17681,N_16758,N_16799);
nand U17682 (N_17682,N_16987,N_16649);
or U17683 (N_17683,N_17305,N_17187);
xor U17684 (N_17684,N_16327,N_16390);
or U17685 (N_17685,N_17147,N_16514);
and U17686 (N_17686,N_16771,N_16565);
or U17687 (N_17687,N_16880,N_16268);
or U17688 (N_17688,N_16523,N_17477);
and U17689 (N_17689,N_16746,N_16817);
nor U17690 (N_17690,N_16960,N_17126);
nor U17691 (N_17691,N_16739,N_16608);
xor U17692 (N_17692,N_17173,N_16484);
xnor U17693 (N_17693,N_17446,N_16532);
xor U17694 (N_17694,N_16319,N_16297);
and U17695 (N_17695,N_16359,N_16892);
nor U17696 (N_17696,N_16288,N_16969);
xnor U17697 (N_17697,N_17252,N_16948);
nand U17698 (N_17698,N_16498,N_17403);
or U17699 (N_17699,N_16643,N_17017);
nor U17700 (N_17700,N_16831,N_17309);
xor U17701 (N_17701,N_17228,N_17157);
or U17702 (N_17702,N_16562,N_16395);
nand U17703 (N_17703,N_16559,N_17227);
or U17704 (N_17704,N_17204,N_16915);
or U17705 (N_17705,N_16819,N_16651);
and U17706 (N_17706,N_16321,N_17238);
and U17707 (N_17707,N_16980,N_17494);
or U17708 (N_17708,N_17413,N_16782);
xnor U17709 (N_17709,N_17399,N_17430);
nor U17710 (N_17710,N_16420,N_16888);
and U17711 (N_17711,N_17196,N_17239);
xnor U17712 (N_17712,N_16955,N_16353);
nor U17713 (N_17713,N_17207,N_17053);
nand U17714 (N_17714,N_16647,N_16749);
and U17715 (N_17715,N_16874,N_16323);
nand U17716 (N_17716,N_16538,N_17091);
nand U17717 (N_17717,N_16646,N_16503);
nor U17718 (N_17718,N_16781,N_17019);
nor U17719 (N_17719,N_16850,N_17248);
or U17720 (N_17720,N_17439,N_17261);
nor U17721 (N_17721,N_16696,N_16631);
nand U17722 (N_17722,N_17397,N_16768);
and U17723 (N_17723,N_17172,N_17330);
or U17724 (N_17724,N_17066,N_17451);
nand U17725 (N_17725,N_17216,N_17409);
nand U17726 (N_17726,N_17189,N_17185);
or U17727 (N_17727,N_16873,N_17226);
nand U17728 (N_17728,N_17340,N_16798);
and U17729 (N_17729,N_16882,N_16476);
nand U17730 (N_17730,N_17245,N_16721);
nand U17731 (N_17731,N_16853,N_17443);
and U17732 (N_17732,N_17360,N_17316);
nand U17733 (N_17733,N_16909,N_17230);
nor U17734 (N_17734,N_16277,N_17368);
xor U17735 (N_17735,N_16366,N_16474);
or U17736 (N_17736,N_16468,N_17302);
and U17737 (N_17737,N_16774,N_16414);
and U17738 (N_17738,N_17099,N_16417);
and U17739 (N_17739,N_17229,N_17457);
nor U17740 (N_17740,N_16709,N_16668);
nand U17741 (N_17741,N_16369,N_16697);
xnor U17742 (N_17742,N_16529,N_16871);
and U17743 (N_17743,N_17139,N_17011);
nor U17744 (N_17744,N_17476,N_16993);
or U17745 (N_17745,N_16511,N_17181);
and U17746 (N_17746,N_16443,N_17471);
xnor U17747 (N_17747,N_16410,N_16766);
and U17748 (N_17748,N_17137,N_16343);
nand U17749 (N_17749,N_17103,N_17093);
nand U17750 (N_17750,N_17322,N_17178);
or U17751 (N_17751,N_17043,N_17349);
nor U17752 (N_17752,N_17442,N_16795);
xnor U17753 (N_17753,N_16787,N_17027);
and U17754 (N_17754,N_16526,N_16499);
and U17755 (N_17755,N_17028,N_16925);
nor U17756 (N_17756,N_16515,N_16522);
and U17757 (N_17757,N_17094,N_17186);
nand U17758 (N_17758,N_17062,N_17282);
xor U17759 (N_17759,N_17166,N_17131);
xnor U17760 (N_17760,N_17183,N_17279);
and U17761 (N_17761,N_16478,N_16810);
nor U17762 (N_17762,N_16378,N_16405);
and U17763 (N_17763,N_16744,N_16788);
or U17764 (N_17764,N_16614,N_17215);
or U17765 (N_17765,N_16491,N_16881);
xnor U17766 (N_17766,N_17319,N_16509);
nand U17767 (N_17767,N_16381,N_16477);
xnor U17768 (N_17768,N_16843,N_17410);
nor U17769 (N_17769,N_16849,N_17351);
nand U17770 (N_17770,N_16463,N_16282);
nand U17771 (N_17771,N_17209,N_16751);
nor U17772 (N_17772,N_17329,N_17395);
and U17773 (N_17773,N_16440,N_16629);
xnor U17774 (N_17774,N_16632,N_16501);
xnor U17775 (N_17775,N_17311,N_16464);
nor U17776 (N_17776,N_16361,N_16970);
xnor U17777 (N_17777,N_16963,N_16972);
and U17778 (N_17778,N_16896,N_16578);
or U17779 (N_17779,N_16539,N_16907);
xor U17780 (N_17780,N_17140,N_16784);
nor U17781 (N_17781,N_16572,N_16752);
nand U17782 (N_17782,N_16699,N_16457);
xnor U17783 (N_17783,N_16821,N_16485);
and U17784 (N_17784,N_16753,N_17064);
xor U17785 (N_17785,N_17039,N_16885);
and U17786 (N_17786,N_17325,N_16254);
and U17787 (N_17787,N_17314,N_17008);
and U17788 (N_17788,N_17396,N_17493);
or U17789 (N_17789,N_17376,N_16828);
and U17790 (N_17790,N_16918,N_17004);
nand U17791 (N_17791,N_16314,N_16287);
xor U17792 (N_17792,N_16580,N_16377);
and U17793 (N_17793,N_17433,N_17085);
xor U17794 (N_17794,N_16382,N_17155);
nand U17795 (N_17795,N_16465,N_17057);
nand U17796 (N_17796,N_16899,N_16660);
or U17797 (N_17797,N_16341,N_16641);
xnor U17798 (N_17798,N_17312,N_17022);
nor U17799 (N_17799,N_17235,N_16957);
or U17800 (N_17800,N_16318,N_17391);
nand U17801 (N_17801,N_16645,N_17096);
nand U17802 (N_17802,N_16483,N_16692);
nand U17803 (N_17803,N_16640,N_16889);
or U17804 (N_17804,N_16497,N_16552);
or U17805 (N_17805,N_16404,N_16270);
or U17806 (N_17806,N_16419,N_17374);
nor U17807 (N_17807,N_16348,N_16912);
nand U17808 (N_17808,N_17281,N_17102);
or U17809 (N_17809,N_16737,N_17268);
nor U17810 (N_17810,N_16322,N_16376);
and U17811 (N_17811,N_16595,N_17111);
nand U17812 (N_17812,N_16847,N_17167);
xor U17813 (N_17813,N_16706,N_16308);
or U17814 (N_17814,N_17038,N_16403);
xnor U17815 (N_17815,N_16991,N_17342);
or U17816 (N_17816,N_16990,N_17496);
nor U17817 (N_17817,N_16520,N_17365);
nor U17818 (N_17818,N_16953,N_16567);
and U17819 (N_17819,N_16415,N_16402);
or U17820 (N_17820,N_16835,N_16428);
or U17821 (N_17821,N_16935,N_16848);
nand U17822 (N_17822,N_16506,N_16735);
nand U17823 (N_17823,N_16334,N_16858);
or U17824 (N_17824,N_17052,N_17472);
nor U17825 (N_17825,N_16966,N_16659);
xor U17826 (N_17826,N_17445,N_17208);
nor U17827 (N_17827,N_16427,N_16407);
nand U17828 (N_17828,N_17447,N_17372);
and U17829 (N_17829,N_16891,N_17023);
nor U17830 (N_17830,N_16610,N_16258);
nand U17831 (N_17831,N_16725,N_17068);
xor U17832 (N_17832,N_17369,N_16708);
nand U17833 (N_17833,N_16517,N_17240);
nand U17834 (N_17834,N_17250,N_16429);
or U17835 (N_17835,N_17389,N_17251);
xor U17836 (N_17836,N_16454,N_16728);
or U17837 (N_17837,N_17489,N_17320);
nand U17838 (N_17838,N_16906,N_17135);
nand U17839 (N_17839,N_16422,N_16808);
and U17840 (N_17840,N_17134,N_17406);
and U17841 (N_17841,N_16475,N_17149);
nor U17842 (N_17842,N_16619,N_16703);
and U17843 (N_17843,N_16320,N_17272);
or U17844 (N_17844,N_16545,N_16411);
nand U17845 (N_17845,N_17431,N_17487);
nand U17846 (N_17846,N_16688,N_16298);
and U17847 (N_17847,N_16911,N_16785);
nor U17848 (N_17848,N_16883,N_16820);
or U17849 (N_17849,N_16666,N_17274);
and U17850 (N_17850,N_17307,N_16387);
nor U17851 (N_17851,N_16346,N_17016);
xor U17852 (N_17852,N_17336,N_17202);
and U17853 (N_17853,N_17010,N_17357);
xor U17854 (N_17854,N_16829,N_17467);
nor U17855 (N_17855,N_16470,N_17294);
nor U17856 (N_17856,N_16797,N_16250);
nand U17857 (N_17857,N_16975,N_17498);
xor U17858 (N_17858,N_17129,N_16793);
nand U17859 (N_17859,N_16736,N_16926);
xor U17860 (N_17860,N_16536,N_16269);
or U17861 (N_17861,N_17171,N_17363);
xor U17862 (N_17862,N_16272,N_17378);
xnor U17863 (N_17863,N_17191,N_17060);
xnor U17864 (N_17864,N_17412,N_17232);
or U17865 (N_17865,N_16328,N_16574);
or U17866 (N_17866,N_16504,N_17084);
nor U17867 (N_17867,N_17199,N_16976);
nor U17868 (N_17868,N_17138,N_17401);
or U17869 (N_17869,N_16650,N_16832);
nand U17870 (N_17870,N_16305,N_17040);
nor U17871 (N_17871,N_16644,N_16727);
and U17872 (N_17872,N_17463,N_17354);
and U17873 (N_17873,N_16988,N_16315);
or U17874 (N_17874,N_17254,N_17486);
and U17875 (N_17875,N_17299,N_17092);
or U17876 (N_17876,N_16563,N_16362);
nand U17877 (N_17877,N_16274,N_17277);
and U17878 (N_17878,N_17269,N_16615);
nand U17879 (N_17879,N_17083,N_16622);
nor U17880 (N_17880,N_16566,N_16549);
or U17881 (N_17881,N_16332,N_16418);
or U17882 (N_17882,N_17356,N_17214);
xnor U17883 (N_17883,N_16505,N_16432);
and U17884 (N_17884,N_16352,N_16996);
nand U17885 (N_17885,N_16921,N_17082);
nand U17886 (N_17886,N_16852,N_16867);
or U17887 (N_17887,N_17224,N_16783);
nor U17888 (N_17888,N_17317,N_16356);
nor U17889 (N_17889,N_16947,N_17353);
and U17890 (N_17890,N_16304,N_16374);
xnor U17891 (N_17891,N_17432,N_16621);
and U17892 (N_17892,N_16648,N_17488);
and U17893 (N_17893,N_16833,N_16544);
and U17894 (N_17894,N_16804,N_16861);
nand U17895 (N_17895,N_16695,N_16555);
and U17896 (N_17896,N_16634,N_17177);
nand U17897 (N_17897,N_17175,N_17194);
and U17898 (N_17898,N_16982,N_16743);
and U17899 (N_17899,N_16557,N_17333);
or U17900 (N_17900,N_16680,N_17465);
and U17901 (N_17901,N_17241,N_16652);
nand U17902 (N_17902,N_17063,N_16449);
or U17903 (N_17903,N_17090,N_16337);
nand U17904 (N_17904,N_16901,N_16461);
nand U17905 (N_17905,N_17414,N_16698);
and U17906 (N_17906,N_17125,N_17499);
nand U17907 (N_17907,N_17427,N_16898);
or U17908 (N_17908,N_16253,N_16790);
nor U17909 (N_17909,N_16636,N_16920);
or U17910 (N_17910,N_16508,N_17036);
or U17911 (N_17911,N_16999,N_16940);
or U17912 (N_17912,N_17386,N_16923);
or U17913 (N_17913,N_16902,N_16738);
nand U17914 (N_17914,N_17474,N_16294);
nor U17915 (N_17915,N_17310,N_17404);
and U17916 (N_17916,N_17328,N_17059);
or U17917 (N_17917,N_17303,N_17405);
and U17918 (N_17918,N_17097,N_16759);
xor U17919 (N_17919,N_17015,N_16408);
or U17920 (N_17920,N_16730,N_17415);
xor U17921 (N_17921,N_16301,N_16460);
or U17922 (N_17922,N_16862,N_16375);
nor U17923 (N_17923,N_16585,N_16998);
or U17924 (N_17924,N_17073,N_17045);
and U17925 (N_17925,N_17480,N_16459);
or U17926 (N_17926,N_17244,N_16264);
xor U17927 (N_17927,N_16576,N_17421);
and U17928 (N_17928,N_16714,N_16311);
nor U17929 (N_17929,N_16265,N_17213);
xnor U17930 (N_17930,N_16625,N_17095);
nand U17931 (N_17931,N_17344,N_16575);
or U17932 (N_17932,N_17000,N_16866);
xnor U17933 (N_17933,N_16528,N_16949);
or U17934 (N_17934,N_16471,N_16397);
or U17935 (N_17935,N_16516,N_17364);
xnor U17936 (N_17936,N_16519,N_16724);
nor U17937 (N_17937,N_16662,N_16278);
nand U17938 (N_17938,N_17089,N_17222);
xor U17939 (N_17939,N_17258,N_17398);
and U17940 (N_17940,N_17012,N_17459);
or U17941 (N_17941,N_16661,N_16452);
xor U17942 (N_17942,N_16780,N_16965);
or U17943 (N_17943,N_16518,N_17221);
nor U17944 (N_17944,N_17259,N_16741);
nand U17945 (N_17945,N_17438,N_16942);
and U17946 (N_17946,N_17058,N_16486);
or U17947 (N_17947,N_17383,N_17034);
and U17948 (N_17948,N_17492,N_16261);
nor U17949 (N_17949,N_17203,N_16917);
nand U17950 (N_17950,N_16560,N_16686);
nor U17951 (N_17951,N_16840,N_16612);
or U17952 (N_17952,N_17260,N_16556);
or U17953 (N_17953,N_17256,N_16674);
nor U17954 (N_17954,N_17375,N_17003);
and U17955 (N_17955,N_16956,N_16755);
nand U17956 (N_17956,N_16338,N_16360);
or U17957 (N_17957,N_17142,N_17420);
xnor U17958 (N_17958,N_16393,N_17370);
or U17959 (N_17959,N_17257,N_17188);
or U17960 (N_17960,N_17210,N_17247);
or U17961 (N_17961,N_16351,N_17108);
or U17962 (N_17962,N_17117,N_16494);
or U17963 (N_17963,N_17287,N_16579);
and U17964 (N_17964,N_17141,N_16283);
xor U17965 (N_17965,N_17341,N_17466);
nand U17966 (N_17966,N_17242,N_17456);
or U17967 (N_17967,N_16776,N_16978);
nor U17968 (N_17968,N_16262,N_16531);
and U17969 (N_17969,N_17461,N_16584);
or U17970 (N_17970,N_16877,N_17265);
nand U17971 (N_17971,N_17121,N_16941);
xor U17972 (N_17972,N_16653,N_17035);
or U17973 (N_17973,N_16945,N_16671);
and U17974 (N_17974,N_16628,N_16365);
nand U17975 (N_17975,N_16548,N_17246);
nand U17976 (N_17976,N_16824,N_17495);
nor U17977 (N_17977,N_17074,N_17490);
xnor U17978 (N_17978,N_16601,N_16865);
or U17979 (N_17979,N_16837,N_16756);
nor U17980 (N_17980,N_16333,N_16616);
xnor U17981 (N_17981,N_16302,N_17223);
nor U17982 (N_17982,N_16958,N_16291);
xnor U17983 (N_17983,N_17331,N_17217);
and U17984 (N_17984,N_16687,N_16259);
or U17985 (N_17985,N_16905,N_16303);
or U17986 (N_17986,N_17408,N_17061);
nor U17987 (N_17987,N_16705,N_17120);
xnor U17988 (N_17988,N_16878,N_17361);
nand U17989 (N_17989,N_16573,N_16908);
xor U17990 (N_17990,N_17031,N_17087);
or U17991 (N_17991,N_17144,N_16903);
or U17992 (N_17992,N_17150,N_17253);
or U17993 (N_17993,N_17107,N_16591);
nor U17994 (N_17994,N_16974,N_17352);
nor U17995 (N_17995,N_17483,N_16430);
and U17996 (N_17996,N_16602,N_17491);
nor U17997 (N_17997,N_17007,N_16472);
nand U17998 (N_17998,N_16597,N_16812);
xor U17999 (N_17999,N_17069,N_17205);
nand U18000 (N_18000,N_16251,N_17211);
nor U18001 (N_18001,N_16846,N_17136);
and U18002 (N_18002,N_16586,N_17345);
nand U18003 (N_18003,N_16510,N_16971);
or U18004 (N_18004,N_17324,N_16604);
or U18005 (N_18005,N_16599,N_16934);
or U18006 (N_18006,N_16655,N_16620);
nor U18007 (N_18007,N_16260,N_17243);
nor U18008 (N_18008,N_16451,N_17440);
nand U18009 (N_18009,N_16613,N_16642);
nand U18010 (N_18010,N_17160,N_17156);
nand U18011 (N_18011,N_17037,N_16943);
nand U18012 (N_18012,N_17337,N_16875);
and U18013 (N_18013,N_16711,N_17100);
nand U18014 (N_18014,N_17270,N_17301);
or U18015 (N_18015,N_16587,N_16479);
nand U18016 (N_18016,N_16309,N_16677);
nand U18017 (N_18017,N_16488,N_17273);
nand U18018 (N_18018,N_16569,N_17048);
and U18019 (N_18019,N_17444,N_16462);
nor U18020 (N_18020,N_17373,N_17029);
or U18021 (N_18021,N_16325,N_16553);
and U18022 (N_18022,N_16665,N_16748);
or U18023 (N_18023,N_16895,N_16571);
and U18024 (N_18024,N_17013,N_17056);
or U18025 (N_18025,N_16401,N_17286);
xnor U18026 (N_18026,N_17143,N_17423);
nor U18027 (N_18027,N_16481,N_16630);
and U18028 (N_18028,N_16977,N_17110);
nor U18029 (N_18029,N_17153,N_16354);
nor U18030 (N_18030,N_17086,N_16910);
or U18031 (N_18031,N_17339,N_17482);
or U18032 (N_18032,N_17158,N_16827);
xor U18033 (N_18033,N_16830,N_16300);
nand U18034 (N_18034,N_16715,N_16869);
xnor U18035 (N_18035,N_17298,N_16507);
xnor U18036 (N_18036,N_17362,N_17067);
nand U18037 (N_18037,N_16582,N_17469);
and U18038 (N_18038,N_16933,N_17323);
or U18039 (N_18039,N_16434,N_16707);
xor U18040 (N_18040,N_16754,N_17371);
nor U18041 (N_18041,N_16363,N_17479);
xnor U18042 (N_18042,N_16773,N_17437);
or U18043 (N_18043,N_16712,N_16857);
or U18044 (N_18044,N_17366,N_16533);
xor U18045 (N_18045,N_17112,N_16489);
or U18046 (N_18046,N_16537,N_16859);
and U18047 (N_18047,N_16863,N_16770);
nor U18048 (N_18048,N_17293,N_17350);
nand U18049 (N_18049,N_17295,N_17288);
xor U18050 (N_18050,N_16598,N_17348);
nor U18051 (N_18051,N_16872,N_16550);
xnor U18052 (N_18052,N_17049,N_17197);
xor U18053 (N_18053,N_17267,N_16685);
nand U18054 (N_18054,N_16609,N_16944);
nor U18055 (N_18055,N_17478,N_17425);
xnor U18056 (N_18056,N_17231,N_16425);
nand U18057 (N_18057,N_17276,N_16981);
or U18058 (N_18058,N_16527,N_16255);
or U18059 (N_18059,N_16633,N_16469);
nand U18060 (N_18060,N_16893,N_16693);
xnor U18061 (N_18061,N_16670,N_16761);
nand U18062 (N_18062,N_17315,N_16350);
nand U18063 (N_18063,N_16345,N_16296);
xnor U18064 (N_18064,N_16952,N_17327);
xnor U18065 (N_18065,N_16436,N_16894);
or U18066 (N_18066,N_17400,N_16561);
xor U18067 (N_18067,N_16455,N_16806);
nor U18068 (N_18068,N_16286,N_16370);
xnor U18069 (N_18069,N_17233,N_16383);
or U18070 (N_18070,N_16570,N_17450);
or U18071 (N_18071,N_16772,N_17435);
xnor U18072 (N_18072,N_16983,N_16547);
and U18073 (N_18073,N_17132,N_17018);
or U18074 (N_18074,N_16285,N_17088);
and U18075 (N_18075,N_16513,N_16313);
nor U18076 (N_18076,N_16310,N_17255);
nor U18077 (N_18077,N_17163,N_16702);
xor U18078 (N_18078,N_16635,N_17263);
xnor U18079 (N_18079,N_16968,N_17080);
nor U18080 (N_18080,N_17485,N_17001);
nor U18081 (N_18081,N_16890,N_16731);
xnor U18082 (N_18082,N_16438,N_17182);
and U18083 (N_18083,N_16769,N_16626);
or U18084 (N_18084,N_16413,N_17387);
nor U18085 (N_18085,N_16637,N_16368);
nand U18086 (N_18086,N_17151,N_16331);
nand U18087 (N_18087,N_17411,N_16742);
nor U18088 (N_18088,N_16329,N_17046);
or U18089 (N_18089,N_17055,N_16603);
or U18090 (N_18090,N_16618,N_17101);
or U18091 (N_18091,N_16823,N_17105);
or U18092 (N_18092,N_16876,N_17005);
nor U18093 (N_18093,N_17098,N_17384);
nor U18094 (N_18094,N_16542,N_16684);
nand U18095 (N_18095,N_17426,N_17326);
nor U18096 (N_18096,N_16954,N_16267);
xor U18097 (N_18097,N_16842,N_16717);
xnor U18098 (N_18098,N_16357,N_16879);
and U18099 (N_18099,N_16995,N_16392);
nand U18100 (N_18100,N_16937,N_16854);
nand U18101 (N_18101,N_17169,N_16379);
and U18102 (N_18102,N_16467,N_17452);
xnor U18103 (N_18103,N_17380,N_16938);
nor U18104 (N_18104,N_17190,N_16389);
or U18105 (N_18105,N_16962,N_16669);
and U18106 (N_18106,N_17124,N_16916);
xnor U18107 (N_18107,N_16723,N_17071);
nor U18108 (N_18108,N_16607,N_16521);
or U18109 (N_18109,N_16281,N_16765);
or U18110 (N_18110,N_16600,N_17249);
nand U18111 (N_18111,N_16611,N_17123);
nand U18112 (N_18112,N_16704,N_17355);
nand U18113 (N_18113,N_17184,N_16292);
or U18114 (N_18114,N_17377,N_16672);
and U18115 (N_18115,N_17201,N_16845);
or U18116 (N_18116,N_16433,N_16466);
nand U18117 (N_18117,N_17318,N_16719);
nand U18118 (N_18118,N_16492,N_16421);
xnor U18119 (N_18119,N_17441,N_16367);
xnor U18120 (N_18120,N_16729,N_16273);
nor U18121 (N_18121,N_16312,N_16673);
xnor U18122 (N_18122,N_17065,N_17266);
and U18123 (N_18123,N_17343,N_16716);
and U18124 (N_18124,N_17321,N_16733);
nor U18125 (N_18125,N_17113,N_16590);
nor U18126 (N_18126,N_16602,N_16869);
nor U18127 (N_18127,N_16634,N_17213);
and U18128 (N_18128,N_16982,N_16324);
or U18129 (N_18129,N_16261,N_16369);
nor U18130 (N_18130,N_16865,N_16969);
nor U18131 (N_18131,N_17450,N_17397);
nand U18132 (N_18132,N_17219,N_17064);
or U18133 (N_18133,N_17435,N_16313);
or U18134 (N_18134,N_16921,N_17436);
or U18135 (N_18135,N_16984,N_16923);
or U18136 (N_18136,N_17026,N_16748);
xor U18137 (N_18137,N_17157,N_16262);
or U18138 (N_18138,N_17128,N_17282);
xor U18139 (N_18139,N_16949,N_17105);
nand U18140 (N_18140,N_16827,N_16994);
nand U18141 (N_18141,N_16743,N_17028);
and U18142 (N_18142,N_17170,N_16599);
xor U18143 (N_18143,N_16328,N_16919);
nor U18144 (N_18144,N_16984,N_16296);
and U18145 (N_18145,N_16702,N_17497);
or U18146 (N_18146,N_16463,N_16913);
and U18147 (N_18147,N_16636,N_17025);
and U18148 (N_18148,N_16480,N_16768);
or U18149 (N_18149,N_16675,N_16661);
nand U18150 (N_18150,N_16469,N_16283);
nand U18151 (N_18151,N_16935,N_16932);
nor U18152 (N_18152,N_17189,N_16617);
nor U18153 (N_18153,N_16406,N_17372);
xor U18154 (N_18154,N_17259,N_16858);
nand U18155 (N_18155,N_17240,N_17396);
and U18156 (N_18156,N_17003,N_17355);
and U18157 (N_18157,N_17162,N_17344);
nand U18158 (N_18158,N_16344,N_17207);
and U18159 (N_18159,N_16960,N_16389);
xor U18160 (N_18160,N_17153,N_16661);
nor U18161 (N_18161,N_17172,N_16707);
and U18162 (N_18162,N_16990,N_17235);
nor U18163 (N_18163,N_17370,N_16888);
and U18164 (N_18164,N_17383,N_16361);
nand U18165 (N_18165,N_17452,N_17234);
and U18166 (N_18166,N_16904,N_16581);
nand U18167 (N_18167,N_16566,N_17429);
nand U18168 (N_18168,N_16586,N_16401);
nor U18169 (N_18169,N_16320,N_17136);
or U18170 (N_18170,N_16691,N_16969);
nor U18171 (N_18171,N_17125,N_16613);
or U18172 (N_18172,N_16307,N_16945);
and U18173 (N_18173,N_17488,N_16527);
nand U18174 (N_18174,N_16725,N_16520);
and U18175 (N_18175,N_16314,N_17239);
and U18176 (N_18176,N_16318,N_16367);
nand U18177 (N_18177,N_16375,N_17014);
nand U18178 (N_18178,N_16563,N_16699);
xor U18179 (N_18179,N_17256,N_17087);
and U18180 (N_18180,N_17438,N_17060);
and U18181 (N_18181,N_16532,N_17330);
or U18182 (N_18182,N_17097,N_17248);
nand U18183 (N_18183,N_17211,N_16993);
nand U18184 (N_18184,N_16345,N_16575);
and U18185 (N_18185,N_17196,N_16707);
or U18186 (N_18186,N_16954,N_16622);
nor U18187 (N_18187,N_16872,N_16828);
nand U18188 (N_18188,N_17227,N_16786);
and U18189 (N_18189,N_17124,N_17268);
or U18190 (N_18190,N_17023,N_17342);
xor U18191 (N_18191,N_16734,N_17022);
nand U18192 (N_18192,N_16641,N_16573);
or U18193 (N_18193,N_17420,N_16505);
and U18194 (N_18194,N_16656,N_16320);
or U18195 (N_18195,N_16879,N_16571);
xnor U18196 (N_18196,N_17377,N_17383);
or U18197 (N_18197,N_17455,N_17031);
xor U18198 (N_18198,N_17329,N_17436);
nand U18199 (N_18199,N_17424,N_17143);
nand U18200 (N_18200,N_17457,N_16271);
nor U18201 (N_18201,N_16272,N_16919);
xnor U18202 (N_18202,N_17364,N_16842);
nand U18203 (N_18203,N_16424,N_16694);
and U18204 (N_18204,N_16435,N_17098);
xor U18205 (N_18205,N_17360,N_17046);
nor U18206 (N_18206,N_16792,N_16540);
xor U18207 (N_18207,N_16466,N_16428);
or U18208 (N_18208,N_17216,N_16999);
xor U18209 (N_18209,N_16810,N_16282);
and U18210 (N_18210,N_16972,N_16512);
xnor U18211 (N_18211,N_16447,N_17470);
nor U18212 (N_18212,N_16737,N_16842);
xnor U18213 (N_18213,N_16277,N_16484);
xnor U18214 (N_18214,N_17343,N_17152);
or U18215 (N_18215,N_17105,N_17219);
or U18216 (N_18216,N_17002,N_17413);
xor U18217 (N_18217,N_16702,N_17120);
and U18218 (N_18218,N_16348,N_16516);
or U18219 (N_18219,N_16546,N_16557);
xor U18220 (N_18220,N_16761,N_16955);
nand U18221 (N_18221,N_17406,N_16902);
xor U18222 (N_18222,N_17061,N_17250);
nand U18223 (N_18223,N_17484,N_16488);
and U18224 (N_18224,N_16658,N_16622);
or U18225 (N_18225,N_16837,N_16297);
nor U18226 (N_18226,N_16803,N_16837);
and U18227 (N_18227,N_17473,N_17289);
nand U18228 (N_18228,N_17340,N_16836);
xnor U18229 (N_18229,N_17488,N_16544);
and U18230 (N_18230,N_17299,N_16634);
xnor U18231 (N_18231,N_16304,N_16643);
and U18232 (N_18232,N_16640,N_16418);
nor U18233 (N_18233,N_16492,N_16520);
xor U18234 (N_18234,N_16312,N_16352);
nor U18235 (N_18235,N_16387,N_17305);
or U18236 (N_18236,N_16550,N_17321);
nor U18237 (N_18237,N_17052,N_16553);
and U18238 (N_18238,N_17482,N_17269);
nand U18239 (N_18239,N_16368,N_17371);
xnor U18240 (N_18240,N_17242,N_16414);
and U18241 (N_18241,N_16643,N_16691);
nand U18242 (N_18242,N_16418,N_16259);
or U18243 (N_18243,N_17341,N_17289);
xor U18244 (N_18244,N_17131,N_16920);
and U18245 (N_18245,N_17335,N_17203);
or U18246 (N_18246,N_17383,N_17055);
and U18247 (N_18247,N_16807,N_16924);
or U18248 (N_18248,N_17110,N_16888);
or U18249 (N_18249,N_16317,N_16826);
xor U18250 (N_18250,N_16701,N_16642);
nand U18251 (N_18251,N_16265,N_16678);
nand U18252 (N_18252,N_17482,N_16500);
or U18253 (N_18253,N_16266,N_16477);
and U18254 (N_18254,N_17417,N_17098);
nor U18255 (N_18255,N_17457,N_16365);
nand U18256 (N_18256,N_16398,N_17036);
nand U18257 (N_18257,N_16985,N_17052);
nand U18258 (N_18258,N_16394,N_16710);
xnor U18259 (N_18259,N_16833,N_16268);
nor U18260 (N_18260,N_17125,N_16523);
nand U18261 (N_18261,N_17293,N_16703);
nor U18262 (N_18262,N_16272,N_16264);
xor U18263 (N_18263,N_16781,N_16927);
nor U18264 (N_18264,N_16303,N_16876);
nand U18265 (N_18265,N_16377,N_17471);
xor U18266 (N_18266,N_16561,N_16487);
xnor U18267 (N_18267,N_16958,N_17225);
or U18268 (N_18268,N_16275,N_17449);
xnor U18269 (N_18269,N_16900,N_16332);
xor U18270 (N_18270,N_17279,N_16612);
xor U18271 (N_18271,N_16463,N_16385);
nor U18272 (N_18272,N_17448,N_17426);
nand U18273 (N_18273,N_17483,N_16252);
or U18274 (N_18274,N_16687,N_16785);
xnor U18275 (N_18275,N_16314,N_16442);
or U18276 (N_18276,N_16379,N_16387);
xnor U18277 (N_18277,N_16344,N_16268);
nand U18278 (N_18278,N_16471,N_17123);
or U18279 (N_18279,N_16364,N_16352);
or U18280 (N_18280,N_16832,N_17040);
and U18281 (N_18281,N_17031,N_16783);
nor U18282 (N_18282,N_17043,N_16894);
xor U18283 (N_18283,N_17431,N_16614);
or U18284 (N_18284,N_17341,N_16669);
nor U18285 (N_18285,N_16740,N_16877);
nor U18286 (N_18286,N_16885,N_17401);
nand U18287 (N_18287,N_17330,N_17302);
nand U18288 (N_18288,N_17349,N_17459);
and U18289 (N_18289,N_17458,N_16266);
and U18290 (N_18290,N_16497,N_17359);
xor U18291 (N_18291,N_16300,N_17054);
or U18292 (N_18292,N_16819,N_16892);
and U18293 (N_18293,N_16755,N_16515);
xnor U18294 (N_18294,N_17169,N_16255);
xor U18295 (N_18295,N_16531,N_16309);
xnor U18296 (N_18296,N_17304,N_17492);
nor U18297 (N_18297,N_17278,N_16801);
or U18298 (N_18298,N_16665,N_16615);
xor U18299 (N_18299,N_17087,N_17487);
nand U18300 (N_18300,N_16489,N_17163);
nand U18301 (N_18301,N_16818,N_16387);
nand U18302 (N_18302,N_17360,N_16665);
nor U18303 (N_18303,N_16771,N_17396);
or U18304 (N_18304,N_17044,N_16843);
nand U18305 (N_18305,N_17494,N_16391);
and U18306 (N_18306,N_17378,N_16808);
or U18307 (N_18307,N_16779,N_16760);
and U18308 (N_18308,N_17301,N_16811);
or U18309 (N_18309,N_17084,N_16807);
and U18310 (N_18310,N_16435,N_16785);
nor U18311 (N_18311,N_16602,N_16796);
and U18312 (N_18312,N_17135,N_16336);
and U18313 (N_18313,N_17190,N_16395);
and U18314 (N_18314,N_17280,N_16564);
xor U18315 (N_18315,N_16828,N_16901);
and U18316 (N_18316,N_17244,N_16973);
and U18317 (N_18317,N_16435,N_17118);
xnor U18318 (N_18318,N_17433,N_16361);
or U18319 (N_18319,N_17035,N_16307);
xor U18320 (N_18320,N_16855,N_16597);
or U18321 (N_18321,N_16638,N_17320);
nor U18322 (N_18322,N_16741,N_16438);
nand U18323 (N_18323,N_16737,N_16909);
and U18324 (N_18324,N_17097,N_16912);
xor U18325 (N_18325,N_17227,N_16896);
nor U18326 (N_18326,N_16278,N_17390);
nand U18327 (N_18327,N_17492,N_16654);
nand U18328 (N_18328,N_17231,N_17239);
nor U18329 (N_18329,N_17261,N_17001);
or U18330 (N_18330,N_16383,N_16802);
or U18331 (N_18331,N_17255,N_16446);
nand U18332 (N_18332,N_17367,N_16522);
or U18333 (N_18333,N_16577,N_16466);
or U18334 (N_18334,N_16294,N_16852);
and U18335 (N_18335,N_16327,N_17117);
nor U18336 (N_18336,N_16921,N_17391);
nor U18337 (N_18337,N_16933,N_16936);
xor U18338 (N_18338,N_16653,N_16886);
nand U18339 (N_18339,N_17195,N_17166);
nor U18340 (N_18340,N_16448,N_17014);
nand U18341 (N_18341,N_17306,N_16733);
xor U18342 (N_18342,N_17011,N_16314);
or U18343 (N_18343,N_16643,N_17485);
nor U18344 (N_18344,N_16399,N_17201);
nor U18345 (N_18345,N_17297,N_16785);
xor U18346 (N_18346,N_17389,N_17296);
nor U18347 (N_18347,N_16321,N_17231);
nor U18348 (N_18348,N_16392,N_17289);
or U18349 (N_18349,N_16669,N_16322);
nand U18350 (N_18350,N_16320,N_17295);
nand U18351 (N_18351,N_16730,N_16583);
or U18352 (N_18352,N_17401,N_16988);
nand U18353 (N_18353,N_16695,N_16403);
and U18354 (N_18354,N_17257,N_16979);
and U18355 (N_18355,N_16384,N_16742);
xnor U18356 (N_18356,N_16663,N_17424);
nand U18357 (N_18357,N_17152,N_16920);
xnor U18358 (N_18358,N_17070,N_16988);
or U18359 (N_18359,N_16450,N_17183);
nor U18360 (N_18360,N_16306,N_16405);
and U18361 (N_18361,N_16927,N_16263);
xnor U18362 (N_18362,N_17305,N_16658);
nand U18363 (N_18363,N_16306,N_16590);
or U18364 (N_18364,N_17331,N_16838);
nor U18365 (N_18365,N_16637,N_16301);
and U18366 (N_18366,N_17320,N_16825);
or U18367 (N_18367,N_17264,N_17337);
xnor U18368 (N_18368,N_16508,N_17363);
or U18369 (N_18369,N_17295,N_16749);
nor U18370 (N_18370,N_16269,N_16789);
or U18371 (N_18371,N_16617,N_17149);
nand U18372 (N_18372,N_17473,N_16315);
xnor U18373 (N_18373,N_17265,N_16963);
nor U18374 (N_18374,N_16491,N_16816);
nor U18375 (N_18375,N_16562,N_17402);
xor U18376 (N_18376,N_17355,N_16689);
nand U18377 (N_18377,N_16899,N_16590);
nor U18378 (N_18378,N_17144,N_16581);
or U18379 (N_18379,N_16371,N_16679);
nor U18380 (N_18380,N_17205,N_17496);
and U18381 (N_18381,N_16876,N_17267);
xnor U18382 (N_18382,N_17183,N_17196);
nor U18383 (N_18383,N_16564,N_17277);
xor U18384 (N_18384,N_17128,N_16291);
and U18385 (N_18385,N_17066,N_17414);
xor U18386 (N_18386,N_17440,N_17362);
nor U18387 (N_18387,N_17080,N_16697);
nor U18388 (N_18388,N_16675,N_16644);
or U18389 (N_18389,N_16731,N_16412);
xor U18390 (N_18390,N_16866,N_16552);
nand U18391 (N_18391,N_16471,N_17425);
nand U18392 (N_18392,N_16501,N_16861);
nor U18393 (N_18393,N_16700,N_16966);
xor U18394 (N_18394,N_16754,N_17135);
xnor U18395 (N_18395,N_17111,N_16714);
nor U18396 (N_18396,N_17430,N_16333);
xnor U18397 (N_18397,N_16488,N_17240);
or U18398 (N_18398,N_17444,N_17256);
and U18399 (N_18399,N_16472,N_17171);
nor U18400 (N_18400,N_17329,N_17091);
nor U18401 (N_18401,N_16599,N_17395);
or U18402 (N_18402,N_17129,N_17302);
nand U18403 (N_18403,N_17232,N_16779);
and U18404 (N_18404,N_17333,N_16455);
xor U18405 (N_18405,N_17075,N_16391);
xnor U18406 (N_18406,N_17416,N_17363);
xnor U18407 (N_18407,N_16553,N_16447);
and U18408 (N_18408,N_16787,N_17158);
and U18409 (N_18409,N_17265,N_17257);
nor U18410 (N_18410,N_16807,N_16492);
nand U18411 (N_18411,N_16876,N_17488);
and U18412 (N_18412,N_16407,N_16341);
or U18413 (N_18413,N_17280,N_16824);
xor U18414 (N_18414,N_16499,N_17109);
and U18415 (N_18415,N_16685,N_17088);
xnor U18416 (N_18416,N_17376,N_16623);
nor U18417 (N_18417,N_17004,N_17492);
and U18418 (N_18418,N_16342,N_16494);
nand U18419 (N_18419,N_17068,N_16830);
xnor U18420 (N_18420,N_17291,N_16539);
nand U18421 (N_18421,N_16998,N_16366);
and U18422 (N_18422,N_16843,N_16272);
nand U18423 (N_18423,N_16269,N_17371);
and U18424 (N_18424,N_16832,N_16522);
nand U18425 (N_18425,N_16544,N_17397);
and U18426 (N_18426,N_17190,N_16695);
or U18427 (N_18427,N_16950,N_17394);
and U18428 (N_18428,N_16858,N_16680);
xnor U18429 (N_18429,N_16348,N_17010);
nor U18430 (N_18430,N_16439,N_17464);
xnor U18431 (N_18431,N_16501,N_16571);
nor U18432 (N_18432,N_17369,N_16290);
and U18433 (N_18433,N_16660,N_17322);
and U18434 (N_18434,N_16551,N_17288);
and U18435 (N_18435,N_16903,N_16818);
and U18436 (N_18436,N_17218,N_17388);
and U18437 (N_18437,N_17354,N_17422);
and U18438 (N_18438,N_16334,N_16771);
or U18439 (N_18439,N_16566,N_16474);
xnor U18440 (N_18440,N_16356,N_16415);
or U18441 (N_18441,N_16504,N_16643);
nand U18442 (N_18442,N_16380,N_17394);
and U18443 (N_18443,N_17272,N_17266);
nor U18444 (N_18444,N_17411,N_16594);
nand U18445 (N_18445,N_16786,N_17279);
xor U18446 (N_18446,N_17154,N_16456);
xor U18447 (N_18447,N_17074,N_16310);
nor U18448 (N_18448,N_16808,N_17333);
or U18449 (N_18449,N_16318,N_16903);
and U18450 (N_18450,N_16402,N_17175);
xnor U18451 (N_18451,N_16352,N_16313);
and U18452 (N_18452,N_16332,N_17133);
and U18453 (N_18453,N_16617,N_17045);
and U18454 (N_18454,N_16429,N_16605);
nand U18455 (N_18455,N_17328,N_16347);
and U18456 (N_18456,N_16993,N_17306);
and U18457 (N_18457,N_17047,N_16619);
nor U18458 (N_18458,N_17497,N_16572);
xnor U18459 (N_18459,N_16279,N_16389);
xnor U18460 (N_18460,N_16337,N_16637);
xnor U18461 (N_18461,N_16373,N_17325);
or U18462 (N_18462,N_16400,N_17320);
xnor U18463 (N_18463,N_16982,N_16666);
or U18464 (N_18464,N_17335,N_17434);
and U18465 (N_18465,N_17200,N_16802);
or U18466 (N_18466,N_16647,N_17120);
nand U18467 (N_18467,N_16931,N_17149);
or U18468 (N_18468,N_17120,N_17004);
nor U18469 (N_18469,N_16993,N_16275);
nor U18470 (N_18470,N_16472,N_16639);
nand U18471 (N_18471,N_16750,N_17151);
or U18472 (N_18472,N_16956,N_17305);
nand U18473 (N_18473,N_17293,N_16721);
nand U18474 (N_18474,N_17033,N_16857);
and U18475 (N_18475,N_17381,N_16998);
or U18476 (N_18476,N_17288,N_17013);
xor U18477 (N_18477,N_16342,N_16829);
nor U18478 (N_18478,N_16991,N_16422);
nand U18479 (N_18479,N_16334,N_17348);
nor U18480 (N_18480,N_16762,N_17478);
xnor U18481 (N_18481,N_16639,N_17463);
and U18482 (N_18482,N_17450,N_16606);
and U18483 (N_18483,N_16304,N_16849);
nor U18484 (N_18484,N_16877,N_17011);
or U18485 (N_18485,N_16622,N_16392);
nand U18486 (N_18486,N_16536,N_16287);
or U18487 (N_18487,N_16717,N_17159);
and U18488 (N_18488,N_16927,N_17032);
xor U18489 (N_18489,N_16429,N_16618);
nor U18490 (N_18490,N_17015,N_17231);
and U18491 (N_18491,N_16932,N_17386);
xor U18492 (N_18492,N_17245,N_17361);
nor U18493 (N_18493,N_17272,N_17248);
nand U18494 (N_18494,N_16927,N_16861);
nand U18495 (N_18495,N_17277,N_16269);
nor U18496 (N_18496,N_16908,N_16783);
or U18497 (N_18497,N_16726,N_17095);
nor U18498 (N_18498,N_16447,N_17315);
or U18499 (N_18499,N_17161,N_17357);
and U18500 (N_18500,N_16953,N_17330);
or U18501 (N_18501,N_16288,N_17213);
xnor U18502 (N_18502,N_17454,N_16498);
and U18503 (N_18503,N_17445,N_17496);
xnor U18504 (N_18504,N_16372,N_17146);
nor U18505 (N_18505,N_17208,N_17438);
or U18506 (N_18506,N_17263,N_16590);
and U18507 (N_18507,N_16758,N_16913);
and U18508 (N_18508,N_16875,N_17172);
and U18509 (N_18509,N_16417,N_16989);
nand U18510 (N_18510,N_16767,N_17264);
or U18511 (N_18511,N_17196,N_16361);
xnor U18512 (N_18512,N_17381,N_17457);
or U18513 (N_18513,N_17222,N_16470);
and U18514 (N_18514,N_16712,N_17072);
nor U18515 (N_18515,N_16524,N_16305);
and U18516 (N_18516,N_17436,N_16380);
nand U18517 (N_18517,N_17083,N_17224);
and U18518 (N_18518,N_17409,N_16279);
and U18519 (N_18519,N_16981,N_17308);
nand U18520 (N_18520,N_16628,N_16713);
and U18521 (N_18521,N_16617,N_17119);
nor U18522 (N_18522,N_17308,N_16389);
or U18523 (N_18523,N_16277,N_16649);
and U18524 (N_18524,N_16499,N_16627);
and U18525 (N_18525,N_17432,N_16542);
xor U18526 (N_18526,N_17470,N_17220);
and U18527 (N_18527,N_16491,N_16719);
and U18528 (N_18528,N_17168,N_16464);
or U18529 (N_18529,N_16648,N_16993);
nand U18530 (N_18530,N_17379,N_16486);
and U18531 (N_18531,N_17069,N_16927);
nand U18532 (N_18532,N_16454,N_16576);
xnor U18533 (N_18533,N_16338,N_16435);
and U18534 (N_18534,N_16621,N_17274);
or U18535 (N_18535,N_16269,N_17097);
and U18536 (N_18536,N_17032,N_17437);
xnor U18537 (N_18537,N_16505,N_16300);
or U18538 (N_18538,N_16763,N_16373);
nand U18539 (N_18539,N_17439,N_17413);
nor U18540 (N_18540,N_16974,N_16624);
nor U18541 (N_18541,N_16701,N_17365);
xor U18542 (N_18542,N_16533,N_17316);
or U18543 (N_18543,N_17130,N_16432);
nor U18544 (N_18544,N_16846,N_16575);
nand U18545 (N_18545,N_17253,N_16955);
and U18546 (N_18546,N_17117,N_16893);
xnor U18547 (N_18547,N_17076,N_16587);
or U18548 (N_18548,N_17283,N_16382);
or U18549 (N_18549,N_17207,N_16991);
nand U18550 (N_18550,N_16741,N_16944);
nor U18551 (N_18551,N_16941,N_17231);
nand U18552 (N_18552,N_16455,N_16769);
nor U18553 (N_18553,N_16309,N_17426);
nand U18554 (N_18554,N_16257,N_17462);
nand U18555 (N_18555,N_17354,N_17428);
nor U18556 (N_18556,N_17170,N_16337);
xnor U18557 (N_18557,N_16941,N_16572);
nor U18558 (N_18558,N_17476,N_16269);
nand U18559 (N_18559,N_16483,N_16365);
or U18560 (N_18560,N_17210,N_17225);
nand U18561 (N_18561,N_16881,N_16622);
nand U18562 (N_18562,N_16541,N_17379);
nand U18563 (N_18563,N_17142,N_16572);
or U18564 (N_18564,N_17215,N_17032);
xor U18565 (N_18565,N_17168,N_17180);
xor U18566 (N_18566,N_16983,N_16963);
xor U18567 (N_18567,N_17244,N_16624);
nor U18568 (N_18568,N_17263,N_16739);
or U18569 (N_18569,N_16749,N_16294);
nand U18570 (N_18570,N_16439,N_16669);
nand U18571 (N_18571,N_16331,N_16430);
nor U18572 (N_18572,N_16750,N_16886);
nand U18573 (N_18573,N_16622,N_16703);
or U18574 (N_18574,N_16347,N_17178);
or U18575 (N_18575,N_16350,N_17155);
nor U18576 (N_18576,N_16618,N_16866);
nand U18577 (N_18577,N_16423,N_16586);
and U18578 (N_18578,N_16544,N_16549);
or U18579 (N_18579,N_17125,N_17312);
xnor U18580 (N_18580,N_17160,N_17158);
and U18581 (N_18581,N_17344,N_17498);
or U18582 (N_18582,N_16701,N_17145);
nor U18583 (N_18583,N_16368,N_17293);
xor U18584 (N_18584,N_16297,N_17338);
nor U18585 (N_18585,N_16294,N_16900);
xor U18586 (N_18586,N_16399,N_16283);
nor U18587 (N_18587,N_16653,N_16645);
and U18588 (N_18588,N_17477,N_16737);
or U18589 (N_18589,N_17487,N_16925);
xor U18590 (N_18590,N_17097,N_16784);
nand U18591 (N_18591,N_17460,N_17129);
or U18592 (N_18592,N_17146,N_16286);
nand U18593 (N_18593,N_16262,N_17372);
xor U18594 (N_18594,N_17241,N_16881);
nor U18595 (N_18595,N_16878,N_16344);
or U18596 (N_18596,N_17289,N_17244);
nor U18597 (N_18597,N_16292,N_16936);
or U18598 (N_18598,N_16414,N_16674);
xor U18599 (N_18599,N_16405,N_16429);
nor U18600 (N_18600,N_16972,N_16610);
nor U18601 (N_18601,N_17491,N_16839);
nand U18602 (N_18602,N_16672,N_16465);
nand U18603 (N_18603,N_17308,N_16980);
and U18604 (N_18604,N_17427,N_17129);
and U18605 (N_18605,N_16905,N_17051);
or U18606 (N_18606,N_17327,N_16902);
xor U18607 (N_18607,N_17367,N_16928);
and U18608 (N_18608,N_16555,N_17416);
nand U18609 (N_18609,N_17335,N_17014);
nand U18610 (N_18610,N_17456,N_17321);
and U18611 (N_18611,N_16262,N_16412);
nand U18612 (N_18612,N_17060,N_17072);
and U18613 (N_18613,N_16716,N_17128);
nor U18614 (N_18614,N_16972,N_16334);
xnor U18615 (N_18615,N_16379,N_16338);
xnor U18616 (N_18616,N_17220,N_17173);
and U18617 (N_18617,N_17189,N_16626);
xnor U18618 (N_18618,N_16617,N_16970);
nor U18619 (N_18619,N_16458,N_17218);
or U18620 (N_18620,N_16452,N_17287);
nand U18621 (N_18621,N_17130,N_17288);
and U18622 (N_18622,N_16699,N_16676);
xor U18623 (N_18623,N_16880,N_16781);
nand U18624 (N_18624,N_16931,N_17350);
nor U18625 (N_18625,N_16472,N_16926);
xor U18626 (N_18626,N_17349,N_16634);
and U18627 (N_18627,N_17116,N_16561);
nor U18628 (N_18628,N_16444,N_16620);
xnor U18629 (N_18629,N_17272,N_16599);
nand U18630 (N_18630,N_17329,N_17172);
and U18631 (N_18631,N_16735,N_16710);
and U18632 (N_18632,N_16560,N_17160);
nand U18633 (N_18633,N_16903,N_16866);
xnor U18634 (N_18634,N_17242,N_17073);
nand U18635 (N_18635,N_16811,N_16399);
xor U18636 (N_18636,N_17050,N_17211);
and U18637 (N_18637,N_16521,N_17323);
nor U18638 (N_18638,N_17482,N_17092);
nand U18639 (N_18639,N_16392,N_16929);
nor U18640 (N_18640,N_17002,N_17386);
xor U18641 (N_18641,N_17297,N_17046);
or U18642 (N_18642,N_17191,N_17253);
nor U18643 (N_18643,N_16343,N_16987);
xnor U18644 (N_18644,N_16366,N_16990);
nor U18645 (N_18645,N_16966,N_16622);
nor U18646 (N_18646,N_16432,N_16972);
nand U18647 (N_18647,N_17489,N_16321);
nor U18648 (N_18648,N_16958,N_16430);
and U18649 (N_18649,N_16408,N_16372);
and U18650 (N_18650,N_16807,N_16736);
nand U18651 (N_18651,N_16528,N_16446);
xor U18652 (N_18652,N_16319,N_16676);
nor U18653 (N_18653,N_16352,N_16693);
nand U18654 (N_18654,N_16698,N_17151);
nand U18655 (N_18655,N_17410,N_16463);
and U18656 (N_18656,N_17259,N_16800);
nand U18657 (N_18657,N_17340,N_17219);
and U18658 (N_18658,N_17202,N_16504);
nand U18659 (N_18659,N_16888,N_16316);
xor U18660 (N_18660,N_16481,N_16352);
nand U18661 (N_18661,N_16970,N_17128);
and U18662 (N_18662,N_16428,N_16497);
xor U18663 (N_18663,N_16670,N_17229);
and U18664 (N_18664,N_16590,N_17060);
nand U18665 (N_18665,N_17355,N_16870);
and U18666 (N_18666,N_17461,N_17218);
or U18667 (N_18667,N_16926,N_17305);
and U18668 (N_18668,N_16934,N_17271);
nor U18669 (N_18669,N_16890,N_16716);
or U18670 (N_18670,N_17243,N_16347);
or U18671 (N_18671,N_16801,N_16448);
and U18672 (N_18672,N_17469,N_16553);
xnor U18673 (N_18673,N_17478,N_16586);
or U18674 (N_18674,N_16837,N_16574);
and U18675 (N_18675,N_16529,N_16304);
nor U18676 (N_18676,N_16668,N_17358);
xnor U18677 (N_18677,N_17395,N_17291);
xor U18678 (N_18678,N_16968,N_16571);
or U18679 (N_18679,N_16687,N_16361);
nand U18680 (N_18680,N_16518,N_17484);
xor U18681 (N_18681,N_16394,N_16872);
and U18682 (N_18682,N_17325,N_16274);
nor U18683 (N_18683,N_17272,N_17280);
and U18684 (N_18684,N_17205,N_16608);
xor U18685 (N_18685,N_16361,N_17287);
nand U18686 (N_18686,N_17461,N_16662);
or U18687 (N_18687,N_17260,N_17165);
xnor U18688 (N_18688,N_17142,N_17301);
or U18689 (N_18689,N_17443,N_17170);
xor U18690 (N_18690,N_16920,N_16335);
or U18691 (N_18691,N_17438,N_17122);
nand U18692 (N_18692,N_17497,N_16469);
nand U18693 (N_18693,N_16921,N_17291);
nor U18694 (N_18694,N_17128,N_16610);
xor U18695 (N_18695,N_16717,N_17408);
nand U18696 (N_18696,N_17321,N_16519);
nor U18697 (N_18697,N_16396,N_16490);
and U18698 (N_18698,N_17335,N_16719);
nand U18699 (N_18699,N_17349,N_16464);
or U18700 (N_18700,N_17053,N_17196);
nor U18701 (N_18701,N_17323,N_17256);
and U18702 (N_18702,N_17247,N_17014);
or U18703 (N_18703,N_17351,N_16951);
or U18704 (N_18704,N_17155,N_16695);
or U18705 (N_18705,N_16345,N_16292);
xnor U18706 (N_18706,N_16699,N_17059);
and U18707 (N_18707,N_17466,N_16941);
and U18708 (N_18708,N_17235,N_16844);
or U18709 (N_18709,N_16613,N_16569);
xnor U18710 (N_18710,N_17361,N_17365);
nand U18711 (N_18711,N_17146,N_16484);
or U18712 (N_18712,N_17297,N_17041);
nand U18713 (N_18713,N_16476,N_17393);
nand U18714 (N_18714,N_16607,N_16567);
nor U18715 (N_18715,N_16705,N_17344);
nand U18716 (N_18716,N_17294,N_16382);
or U18717 (N_18717,N_16342,N_16597);
nor U18718 (N_18718,N_17038,N_16825);
or U18719 (N_18719,N_16257,N_16655);
xnor U18720 (N_18720,N_17411,N_16326);
nand U18721 (N_18721,N_16674,N_17092);
nor U18722 (N_18722,N_17114,N_17103);
nor U18723 (N_18723,N_16288,N_16821);
xnor U18724 (N_18724,N_16483,N_17126);
nor U18725 (N_18725,N_16379,N_16752);
nand U18726 (N_18726,N_16963,N_16721);
or U18727 (N_18727,N_17033,N_16758);
nor U18728 (N_18728,N_17177,N_16423);
xor U18729 (N_18729,N_17310,N_17033);
nand U18730 (N_18730,N_17322,N_16394);
and U18731 (N_18731,N_16856,N_16586);
and U18732 (N_18732,N_16262,N_16482);
xnor U18733 (N_18733,N_16647,N_16788);
xor U18734 (N_18734,N_16778,N_16881);
or U18735 (N_18735,N_16702,N_17253);
or U18736 (N_18736,N_16530,N_16494);
and U18737 (N_18737,N_17412,N_16571);
and U18738 (N_18738,N_16572,N_17234);
xnor U18739 (N_18739,N_16477,N_17357);
nand U18740 (N_18740,N_16563,N_16955);
nand U18741 (N_18741,N_16633,N_16719);
and U18742 (N_18742,N_16957,N_16357);
and U18743 (N_18743,N_16342,N_17238);
xnor U18744 (N_18744,N_16519,N_16332);
nand U18745 (N_18745,N_16586,N_17237);
nor U18746 (N_18746,N_16897,N_16943);
and U18747 (N_18747,N_17027,N_16881);
and U18748 (N_18748,N_16869,N_16485);
or U18749 (N_18749,N_17393,N_16412);
or U18750 (N_18750,N_17887,N_18706);
nor U18751 (N_18751,N_17976,N_18558);
nand U18752 (N_18752,N_18180,N_17971);
nor U18753 (N_18753,N_18413,N_18585);
and U18754 (N_18754,N_18130,N_18268);
nor U18755 (N_18755,N_18746,N_17648);
nand U18756 (N_18756,N_18537,N_17566);
and U18757 (N_18757,N_18604,N_18690);
or U18758 (N_18758,N_17684,N_18725);
xor U18759 (N_18759,N_17900,N_18208);
nor U18760 (N_18760,N_17986,N_17657);
or U18761 (N_18761,N_18362,N_17593);
nand U18762 (N_18762,N_18013,N_18552);
and U18763 (N_18763,N_17898,N_18345);
nand U18764 (N_18764,N_18157,N_17987);
nor U18765 (N_18765,N_18113,N_18427);
nor U18766 (N_18766,N_18410,N_18664);
and U18767 (N_18767,N_17542,N_18326);
or U18768 (N_18768,N_17781,N_17868);
and U18769 (N_18769,N_17659,N_17527);
nor U18770 (N_18770,N_18152,N_17520);
xor U18771 (N_18771,N_18512,N_18670);
or U18772 (N_18772,N_18622,N_18490);
nand U18773 (N_18773,N_17760,N_17839);
xnor U18774 (N_18774,N_17553,N_18518);
xor U18775 (N_18775,N_18147,N_17847);
or U18776 (N_18776,N_18112,N_17748);
or U18777 (N_18777,N_18065,N_18545);
or U18778 (N_18778,N_18261,N_18093);
nand U18779 (N_18779,N_18618,N_18574);
and U18780 (N_18780,N_17709,N_17873);
nor U18781 (N_18781,N_17921,N_18207);
and U18782 (N_18782,N_18332,N_18737);
or U18783 (N_18783,N_17942,N_18479);
and U18784 (N_18784,N_18118,N_17766);
and U18785 (N_18785,N_18146,N_18486);
and U18786 (N_18786,N_17687,N_17713);
nor U18787 (N_18787,N_17875,N_17543);
nand U18788 (N_18788,N_17723,N_18262);
and U18789 (N_18789,N_18650,N_17795);
nor U18790 (N_18790,N_17547,N_18662);
and U18791 (N_18791,N_18445,N_18546);
nor U18792 (N_18792,N_17722,N_17886);
nor U18793 (N_18793,N_18695,N_18198);
xor U18794 (N_18794,N_18513,N_18309);
nor U18795 (N_18795,N_18156,N_18425);
xnor U18796 (N_18796,N_17591,N_17779);
nor U18797 (N_18797,N_17843,N_17777);
nor U18798 (N_18798,N_18032,N_17770);
or U18799 (N_18799,N_18615,N_18697);
or U18800 (N_18800,N_18408,N_18699);
or U18801 (N_18801,N_18237,N_17913);
nand U18802 (N_18802,N_17704,N_17824);
and U18803 (N_18803,N_17592,N_18358);
or U18804 (N_18804,N_18224,N_18515);
xor U18805 (N_18805,N_17894,N_18250);
and U18806 (N_18806,N_17644,N_18391);
nand U18807 (N_18807,N_17772,N_18499);
and U18808 (N_18808,N_17915,N_18603);
or U18809 (N_18809,N_17899,N_18483);
or U18810 (N_18810,N_18347,N_18569);
xnor U18811 (N_18811,N_18311,N_18272);
nor U18812 (N_18812,N_18631,N_17934);
nor U18813 (N_18813,N_17833,N_18736);
and U18814 (N_18814,N_18196,N_18641);
xnor U18815 (N_18815,N_17946,N_17743);
and U18816 (N_18816,N_18306,N_17809);
nor U18817 (N_18817,N_18484,N_18243);
and U18818 (N_18818,N_17616,N_18659);
xnor U18819 (N_18819,N_18648,N_17802);
or U18820 (N_18820,N_18307,N_18173);
and U18821 (N_18821,N_17518,N_18142);
or U18822 (N_18822,N_17963,N_18087);
and U18823 (N_18823,N_18133,N_17508);
or U18824 (N_18824,N_18728,N_18097);
xor U18825 (N_18825,N_18556,N_18508);
and U18826 (N_18826,N_18748,N_17874);
or U18827 (N_18827,N_18389,N_18735);
nor U18828 (N_18828,N_17870,N_18566);
nand U18829 (N_18829,N_18459,N_17767);
and U18830 (N_18830,N_18732,N_18608);
and U18831 (N_18831,N_18444,N_18679);
nand U18832 (N_18832,N_17790,N_17500);
and U18833 (N_18833,N_17696,N_18646);
xor U18834 (N_18834,N_17789,N_17736);
xnor U18835 (N_18835,N_18028,N_18671);
xnor U18836 (N_18836,N_17985,N_18709);
or U18837 (N_18837,N_17998,N_18469);
or U18838 (N_18838,N_18205,N_18151);
xor U18839 (N_18839,N_18634,N_18124);
and U18840 (N_18840,N_17679,N_17926);
and U18841 (N_18841,N_17738,N_18015);
nand U18842 (N_18842,N_17923,N_17649);
and U18843 (N_18843,N_18255,N_18046);
nor U18844 (N_18844,N_18303,N_18342);
nor U18845 (N_18845,N_17759,N_18148);
and U18846 (N_18846,N_18242,N_17814);
or U18847 (N_18847,N_17867,N_17594);
or U18848 (N_18848,N_17608,N_18577);
xnor U18849 (N_18849,N_18125,N_17834);
or U18850 (N_18850,N_18005,N_18084);
and U18851 (N_18851,N_18288,N_17561);
and U18852 (N_18852,N_17947,N_18038);
nor U18853 (N_18853,N_17863,N_18526);
xor U18854 (N_18854,N_18098,N_17634);
nor U18855 (N_18855,N_17912,N_18249);
and U18856 (N_18856,N_18052,N_17652);
xnor U18857 (N_18857,N_17981,N_18164);
xor U18858 (N_18858,N_17686,N_17588);
nand U18859 (N_18859,N_18270,N_18562);
nor U18860 (N_18860,N_18683,N_18057);
and U18861 (N_18861,N_18431,N_17851);
nor U18862 (N_18862,N_18007,N_18471);
or U18863 (N_18863,N_18314,N_17600);
and U18864 (N_18864,N_18054,N_17876);
and U18865 (N_18865,N_18467,N_18579);
xor U18866 (N_18866,N_17573,N_17811);
and U18867 (N_18867,N_18397,N_18195);
xor U18868 (N_18868,N_17715,N_17734);
and U18869 (N_18869,N_17504,N_17728);
nor U18870 (N_18870,N_17859,N_17729);
xor U18871 (N_18871,N_17810,N_18589);
nand U18872 (N_18872,N_17521,N_17974);
and U18873 (N_18873,N_18140,N_18300);
and U18874 (N_18874,N_17788,N_18656);
nand U18875 (N_18875,N_18349,N_18139);
and U18876 (N_18876,N_18590,N_18090);
nor U18877 (N_18877,N_17537,N_17852);
nor U18878 (N_18878,N_18310,N_18036);
or U18879 (N_18879,N_18315,N_17975);
xnor U18880 (N_18880,N_17793,N_18000);
nor U18881 (N_18881,N_18259,N_17576);
nand U18882 (N_18882,N_18601,N_17768);
nand U18883 (N_18883,N_17642,N_18570);
nand U18884 (N_18884,N_18060,N_17726);
nor U18885 (N_18885,N_18357,N_18001);
and U18886 (N_18886,N_18014,N_18269);
nand U18887 (N_18887,N_18344,N_17535);
xor U18888 (N_18888,N_18616,N_18406);
nand U18889 (N_18889,N_17840,N_18081);
and U18890 (N_18890,N_18226,N_18210);
and U18891 (N_18891,N_18247,N_17819);
nand U18892 (N_18892,N_17557,N_18305);
or U18893 (N_18893,N_18447,N_18673);
xnor U18894 (N_18894,N_17556,N_17692);
xnor U18895 (N_18895,N_17646,N_17662);
and U18896 (N_18896,N_18131,N_17714);
xnor U18897 (N_18897,N_17994,N_18400);
and U18898 (N_18898,N_18522,N_18366);
nor U18899 (N_18899,N_17671,N_18331);
nor U18900 (N_18900,N_18278,N_18264);
xnor U18901 (N_18901,N_18488,N_17945);
xnor U18902 (N_18902,N_18135,N_17645);
nor U18903 (N_18903,N_18580,N_17820);
or U18904 (N_18904,N_17689,N_18281);
or U18905 (N_18905,N_17961,N_18685);
and U18906 (N_18906,N_17832,N_17702);
nand U18907 (N_18907,N_18030,N_18568);
nor U18908 (N_18908,N_18632,N_18088);
xnor U18909 (N_18909,N_18103,N_18633);
xnor U18910 (N_18910,N_17564,N_18393);
xnor U18911 (N_18911,N_18676,N_18372);
and U18912 (N_18912,N_18394,N_17725);
nor U18913 (N_18913,N_18573,N_18003);
and U18914 (N_18914,N_18635,N_18327);
and U18915 (N_18915,N_18333,N_18064);
nor U18916 (N_18916,N_18402,N_17682);
or U18917 (N_18917,N_17623,N_18168);
xnor U18918 (N_18918,N_18423,N_17904);
and U18919 (N_18919,N_18258,N_17982);
or U18920 (N_18920,N_18544,N_18252);
xnor U18921 (N_18921,N_17812,N_18535);
and U18922 (N_18922,N_17952,N_17813);
and U18923 (N_18923,N_17563,N_17825);
and U18924 (N_18924,N_18026,N_18636);
or U18925 (N_18925,N_17860,N_18598);
or U18926 (N_18926,N_17519,N_17531);
nor U18927 (N_18927,N_18256,N_18630);
nor U18928 (N_18928,N_17602,N_18111);
and U18929 (N_18929,N_18229,N_17619);
nor U18930 (N_18930,N_18215,N_18176);
nand U18931 (N_18931,N_18730,N_17943);
and U18932 (N_18932,N_17651,N_18438);
and U18933 (N_18933,N_17826,N_18285);
nor U18934 (N_18934,N_18586,N_18638);
nor U18935 (N_18935,N_18181,N_17775);
nand U18936 (N_18936,N_18403,N_18099);
nor U18937 (N_18937,N_18409,N_18384);
or U18938 (N_18938,N_17579,N_18387);
and U18939 (N_18939,N_18452,N_18740);
and U18940 (N_18940,N_18405,N_17673);
or U18941 (N_18941,N_18593,N_18025);
or U18942 (N_18942,N_17583,N_18045);
or U18943 (N_18943,N_17685,N_18066);
and U18944 (N_18944,N_18382,N_17621);
nor U18945 (N_18945,N_18612,N_18434);
nand U18946 (N_18946,N_18159,N_18121);
xnor U18947 (N_18947,N_17829,N_18523);
nor U18948 (N_18948,N_18341,N_17567);
nor U18949 (N_18949,N_17895,N_17769);
nor U18950 (N_18950,N_18022,N_18498);
xnor U18951 (N_18951,N_18280,N_18231);
xor U18952 (N_18952,N_17555,N_17710);
or U18953 (N_18953,N_17955,N_17509);
xor U18954 (N_18954,N_18494,N_17925);
nand U18955 (N_18955,N_17808,N_18339);
and U18956 (N_18956,N_17515,N_17750);
and U18957 (N_18957,N_17624,N_17721);
xor U18958 (N_18958,N_18092,N_17718);
nand U18959 (N_18959,N_18031,N_17582);
nand U18960 (N_18960,N_17548,N_18745);
nand U18961 (N_18961,N_17761,N_18693);
nand U18962 (N_18962,N_18435,N_17848);
and U18963 (N_18963,N_17939,N_18448);
xnor U18964 (N_18964,N_18411,N_18719);
nor U18965 (N_18965,N_17916,N_17815);
or U18966 (N_18966,N_17505,N_18338);
or U18967 (N_18967,N_17771,N_18017);
nand U18968 (N_18968,N_18642,N_18596);
nor U18969 (N_18969,N_17636,N_18296);
nand U18970 (N_18970,N_18375,N_18149);
nor U18971 (N_18971,N_17507,N_18449);
and U18972 (N_18972,N_18497,N_17872);
xnor U18973 (N_18973,N_17512,N_17536);
nand U18974 (N_18974,N_17969,N_18716);
nor U18975 (N_18975,N_18298,N_17724);
and U18976 (N_18976,N_17907,N_17892);
or U18977 (N_18977,N_17929,N_18554);
or U18978 (N_18978,N_17617,N_18354);
nor U18979 (N_18979,N_17601,N_18213);
nor U18980 (N_18980,N_17817,N_17575);
nand U18981 (N_18981,N_18378,N_17906);
or U18982 (N_18982,N_17570,N_18487);
nand U18983 (N_18983,N_18398,N_17902);
or U18984 (N_18984,N_18528,N_18591);
nand U18985 (N_18985,N_17711,N_18712);
and U18986 (N_18986,N_18169,N_18478);
nor U18987 (N_18987,N_17574,N_18602);
or U18988 (N_18988,N_17967,N_18192);
xnor U18989 (N_18989,N_18701,N_18502);
xnor U18990 (N_18990,N_17675,N_17676);
or U18991 (N_18991,N_18068,N_18510);
nor U18992 (N_18992,N_18588,N_17691);
nor U18993 (N_18993,N_18455,N_17988);
nor U18994 (N_18994,N_17626,N_17977);
or U18995 (N_18995,N_18276,N_17883);
or U18996 (N_18996,N_18020,N_18238);
or U18997 (N_18997,N_18218,N_17586);
nor U18998 (N_18998,N_18600,N_17694);
nor U18999 (N_18999,N_17745,N_18418);
xor U19000 (N_19000,N_18592,N_18203);
nor U19001 (N_19001,N_18688,N_17911);
and U19002 (N_19002,N_18643,N_17997);
nor U19003 (N_19003,N_18561,N_18110);
and U19004 (N_19004,N_18521,N_17914);
and U19005 (N_19005,N_18419,N_18614);
or U19006 (N_19006,N_18666,N_17803);
nor U19007 (N_19007,N_18658,N_17533);
and U19008 (N_19008,N_18678,N_17910);
nand U19009 (N_19009,N_17908,N_18194);
xor U19010 (N_19010,N_17920,N_17866);
nand U19011 (N_19011,N_18251,N_17558);
xnor U19012 (N_19012,N_18555,N_17855);
nand U19013 (N_19013,N_17854,N_17746);
nor U19014 (N_19014,N_18388,N_18370);
nand U19015 (N_19015,N_17962,N_18514);
nand U19016 (N_19016,N_18334,N_17842);
xor U19017 (N_19017,N_18129,N_17568);
and U19018 (N_19018,N_18325,N_18456);
nor U19019 (N_19019,N_18442,N_18050);
or U19020 (N_19020,N_18532,N_17742);
xnor U19021 (N_19021,N_17554,N_18166);
or U19022 (N_19022,N_18365,N_17927);
nand U19023 (N_19023,N_18233,N_17956);
or U19024 (N_19024,N_17983,N_18086);
nor U19025 (N_19025,N_17990,N_17807);
nor U19026 (N_19026,N_17922,N_17699);
and U19027 (N_19027,N_18669,N_18415);
or U19028 (N_19028,N_18070,N_18077);
or U19029 (N_19029,N_18428,N_18137);
xnor U19030 (N_19030,N_18172,N_18457);
xor U19031 (N_19031,N_18700,N_18677);
or U19032 (N_19032,N_17778,N_18417);
nand U19033 (N_19033,N_18037,N_18346);
nor U19034 (N_19034,N_18282,N_18241);
nand U19035 (N_19035,N_18153,N_18480);
nor U19036 (N_19036,N_18274,N_17841);
nor U19037 (N_19037,N_18421,N_17719);
nand U19038 (N_19038,N_18441,N_17638);
nand U19039 (N_19039,N_18665,N_18012);
nand U19040 (N_19040,N_18254,N_18476);
nor U19041 (N_19041,N_18115,N_17613);
nor U19042 (N_19042,N_17879,N_18074);
xnor U19043 (N_19043,N_18584,N_18234);
or U19044 (N_19044,N_18127,N_18578);
xor U19045 (N_19045,N_17581,N_18175);
nor U19046 (N_19046,N_18067,N_18109);
xnor U19047 (N_19047,N_18043,N_18167);
nand U19048 (N_19048,N_18505,N_17698);
or U19049 (N_19049,N_18379,N_18371);
nor U19050 (N_19050,N_18102,N_17501);
and U19051 (N_19051,N_17791,N_18426);
xnor U19052 (N_19052,N_18197,N_17992);
and U19053 (N_19053,N_18420,N_18011);
nand U19054 (N_19054,N_18609,N_18170);
and U19055 (N_19055,N_18335,N_18707);
xnor U19056 (N_19056,N_17799,N_18684);
nor U19057 (N_19057,N_18567,N_18461);
or U19058 (N_19058,N_17970,N_18155);
or U19059 (N_19059,N_18232,N_17595);
or U19060 (N_19060,N_17656,N_17577);
nor U19061 (N_19061,N_17639,N_17510);
xnor U19062 (N_19062,N_18691,N_18216);
nand U19063 (N_19063,N_17940,N_18481);
or U19064 (N_19064,N_18713,N_18674);
or U19065 (N_19065,N_18248,N_18386);
and U19066 (N_19066,N_18184,N_18524);
nand U19067 (N_19067,N_18714,N_18720);
and U19068 (N_19068,N_17891,N_17610);
nand U19069 (N_19069,N_17516,N_18422);
nand U19070 (N_19070,N_18223,N_17633);
nor U19071 (N_19071,N_17545,N_18516);
and U19072 (N_19072,N_18704,N_18517);
xnor U19073 (N_19073,N_18611,N_18472);
nor U19074 (N_19074,N_18557,N_18308);
or U19075 (N_19075,N_18058,N_18085);
xnor U19076 (N_19076,N_17529,N_18412);
and U19077 (N_19077,N_17950,N_17757);
xnor U19078 (N_19078,N_18451,N_18443);
or U19079 (N_19079,N_18076,N_18289);
nor U19080 (N_19080,N_18655,N_17877);
nor U19081 (N_19081,N_18623,N_18416);
xnor U19082 (N_19082,N_17960,N_18286);
and U19083 (N_19083,N_18396,N_18283);
and U19084 (N_19084,N_17632,N_18343);
xnor U19085 (N_19085,N_18694,N_18385);
xnor U19086 (N_19086,N_18702,N_18163);
nand U19087 (N_19087,N_18477,N_18548);
nand U19088 (N_19088,N_18401,N_17905);
and U19089 (N_19089,N_18436,N_17928);
xnor U19090 (N_19090,N_18547,N_18581);
and U19091 (N_19091,N_17578,N_18189);
nand U19092 (N_19092,N_18267,N_17993);
nor U19093 (N_19093,N_17957,N_17890);
nand U19094 (N_19094,N_18468,N_17631);
xor U19095 (N_19095,N_17753,N_18294);
and U19096 (N_19096,N_17706,N_18539);
nand U19097 (N_19097,N_17612,N_17665);
xor U19098 (N_19098,N_17933,N_18661);
xor U19099 (N_19099,N_17801,N_17917);
and U19100 (N_19100,N_18051,N_18742);
or U19101 (N_19101,N_17805,N_18359);
and U19102 (N_19102,N_17862,N_18575);
nand U19103 (N_19103,N_18473,N_18626);
and U19104 (N_19104,N_18549,N_17739);
xnor U19105 (N_19105,N_17630,N_18246);
or U19106 (N_19106,N_18743,N_18299);
xnor U19107 (N_19107,N_18217,N_18291);
xor U19108 (N_19108,N_18188,N_18221);
and U19109 (N_19109,N_18089,N_18450);
nand U19110 (N_19110,N_18404,N_18531);
nand U19111 (N_19111,N_18744,N_18689);
xnor U19112 (N_19112,N_17944,N_18199);
or U19113 (N_19113,N_18230,N_17680);
xor U19114 (N_19114,N_18747,N_17909);
nor U19115 (N_19115,N_18639,N_17930);
xor U19116 (N_19116,N_17999,N_18640);
or U19117 (N_19117,N_17620,N_18080);
and U19118 (N_19118,N_18733,N_18395);
nor U19119 (N_19119,N_18072,N_18644);
nand U19120 (N_19120,N_18739,N_18543);
nand U19121 (N_19121,N_18317,N_18201);
and U19122 (N_19122,N_18209,N_18474);
or U19123 (N_19123,N_18263,N_18019);
xnor U19124 (N_19124,N_17605,N_17513);
or U19125 (N_19125,N_18200,N_18680);
nand U19126 (N_19126,N_18161,N_17937);
nor U19127 (N_19127,N_18729,N_17749);
nor U19128 (N_19128,N_18062,N_17972);
and U19129 (N_19129,N_18035,N_18492);
and U19130 (N_19130,N_17511,N_18287);
xnor U19131 (N_19131,N_18322,N_17818);
nor U19132 (N_19132,N_18571,N_18185);
and U19133 (N_19133,N_18033,N_18075);
xor U19134 (N_19134,N_18668,N_18667);
or U19135 (N_19135,N_18637,N_17763);
nor U19136 (N_19136,N_18040,N_18039);
or U19137 (N_19137,N_17953,N_17502);
nand U19138 (N_19138,N_17858,N_18144);
and U19139 (N_19139,N_17599,N_17935);
nand U19140 (N_19140,N_17672,N_17526);
and U19141 (N_19141,N_18703,N_18091);
and U19142 (N_19142,N_17762,N_18430);
xor U19143 (N_19143,N_18367,N_18219);
nor U19144 (N_19144,N_18458,N_18078);
and U19145 (N_19145,N_18708,N_18150);
and U19146 (N_19146,N_17727,N_18453);
or U19147 (N_19147,N_17647,N_18493);
or U19148 (N_19148,N_18266,N_18542);
or U19149 (N_19149,N_17755,N_17881);
and U19150 (N_19150,N_18204,N_18337);
nand U19151 (N_19151,N_17845,N_17782);
nor U19152 (N_19152,N_18465,N_17571);
or U19153 (N_19153,N_17517,N_18519);
nand U19154 (N_19154,N_17549,N_17794);
and U19155 (N_19155,N_18016,N_18023);
nor U19156 (N_19156,N_18353,N_18228);
or U19157 (N_19157,N_18122,N_17635);
and U19158 (N_19158,N_18705,N_18594);
or U19159 (N_19159,N_18460,N_17800);
nor U19160 (N_19160,N_17625,N_18120);
xor U19161 (N_19161,N_18654,N_18212);
or U19162 (N_19162,N_17717,N_17544);
nor U19163 (N_19163,N_17798,N_18336);
or U19164 (N_19164,N_18560,N_18466);
and U19165 (N_19165,N_17831,N_18214);
xor U19166 (N_19166,N_17654,N_18304);
nor U19167 (N_19167,N_17756,N_18564);
or U19168 (N_19168,N_18158,N_17850);
xor U19169 (N_19169,N_17965,N_18348);
and U19170 (N_19170,N_17663,N_18463);
and U19171 (N_19171,N_18356,N_18236);
nor U19172 (N_19172,N_18605,N_17783);
nor U19173 (N_19173,N_17597,N_18414);
and U19174 (N_19174,N_17700,N_17754);
nor U19175 (N_19175,N_17655,N_18437);
xor U19176 (N_19176,N_17774,N_17560);
nand U19177 (N_19177,N_18063,N_17747);
nand U19178 (N_19178,N_17524,N_18536);
nor U19179 (N_19179,N_17936,N_18374);
nor U19180 (N_19180,N_18718,N_18597);
nand U19181 (N_19181,N_18491,N_17984);
nand U19182 (N_19182,N_18710,N_18048);
or U19183 (N_19183,N_18530,N_18587);
or U19184 (N_19184,N_18625,N_18407);
nor U19185 (N_19185,N_17784,N_17707);
nor U19186 (N_19186,N_18029,N_18079);
and U19187 (N_19187,N_18565,N_18319);
nor U19188 (N_19188,N_17864,N_17780);
nand U19189 (N_19189,N_17776,N_18101);
xnor U19190 (N_19190,N_18006,N_18541);
and U19191 (N_19191,N_17740,N_17959);
nand U19192 (N_19192,N_18645,N_18100);
nor U19193 (N_19193,N_18056,N_18094);
nor U19194 (N_19194,N_18002,N_18027);
and U19195 (N_19195,N_17951,N_18681);
and U19196 (N_19196,N_18369,N_18190);
or U19197 (N_19197,N_18061,N_17973);
and U19198 (N_19198,N_18318,N_18621);
nor U19199 (N_19199,N_18559,N_18360);
nor U19200 (N_19200,N_18297,N_17844);
and U19201 (N_19201,N_18160,N_17765);
nand U19202 (N_19202,N_18320,N_18350);
xor U19203 (N_19203,N_17585,N_17741);
nor U19204 (N_19204,N_18682,N_18134);
and U19205 (N_19205,N_18138,N_17932);
or U19206 (N_19206,N_18734,N_17628);
xor U19207 (N_19207,N_18741,N_17764);
nand U19208 (N_19208,N_18495,N_17822);
nor U19209 (N_19209,N_17681,N_18328);
nor U19210 (N_19210,N_18106,N_18187);
nor U19211 (N_19211,N_18024,N_18119);
nor U19212 (N_19212,N_17587,N_18145);
nand U19213 (N_19213,N_17835,N_17828);
and U19214 (N_19214,N_17893,N_17562);
nor U19215 (N_19215,N_18227,N_18330);
or U19216 (N_19216,N_18723,N_18186);
nand U19217 (N_19217,N_18538,N_18351);
nand U19218 (N_19218,N_18302,N_18116);
xnor U19219 (N_19219,N_18312,N_17611);
xnor U19220 (N_19220,N_17701,N_17786);
nand U19221 (N_19221,N_17506,N_18222);
nor U19222 (N_19222,N_17958,N_18010);
nand U19223 (N_19223,N_18462,N_18211);
or U19224 (N_19224,N_18533,N_18340);
nor U19225 (N_19225,N_18301,N_17615);
xnor U19226 (N_19226,N_18273,N_18162);
nand U19227 (N_19227,N_17731,N_17806);
or U19228 (N_19228,N_18021,N_17683);
and U19229 (N_19229,N_18323,N_18563);
nand U19230 (N_19230,N_17816,N_18165);
nor U19231 (N_19231,N_18525,N_18154);
nor U19232 (N_19232,N_17532,N_17796);
and U19233 (N_19233,N_18620,N_17996);
nor U19234 (N_19234,N_18657,N_17674);
and U19235 (N_19235,N_18293,N_17903);
nor U19236 (N_19236,N_17804,N_17797);
and U19237 (N_19237,N_18277,N_18202);
nor U19238 (N_19238,N_17751,N_17607);
nand U19239 (N_19239,N_17550,N_18653);
or U19240 (N_19240,N_18649,N_18429);
xnor U19241 (N_19241,N_18380,N_18726);
nor U19242 (N_19242,N_18717,N_17614);
or U19243 (N_19243,N_18117,N_18352);
nor U19244 (N_19244,N_18610,N_17658);
xnor U19245 (N_19245,N_18183,N_18627);
nor U19246 (N_19246,N_17627,N_17735);
nand U19247 (N_19247,N_17565,N_18179);
nor U19248 (N_19248,N_17838,N_18279);
nand U19249 (N_19249,N_17853,N_17618);
nand U19250 (N_19250,N_18324,N_18275);
xnor U19251 (N_19251,N_18253,N_18722);
xnor U19252 (N_19252,N_17871,N_17865);
nor U19253 (N_19253,N_17732,N_18044);
and U19254 (N_19254,N_17737,N_17688);
xor U19255 (N_19255,N_18381,N_17968);
or U19256 (N_19256,N_17604,N_17857);
or U19257 (N_19257,N_17979,N_17534);
nand U19258 (N_19258,N_17643,N_18053);
and U19259 (N_19259,N_17896,N_18440);
nand U19260 (N_19260,N_17606,N_17693);
xnor U19261 (N_19261,N_17569,N_18008);
and U19262 (N_19262,N_17538,N_18143);
nand U19263 (N_19263,N_18599,N_18383);
nor U19264 (N_19264,N_18047,N_18595);
or U19265 (N_19265,N_17880,N_18182);
nor U19266 (N_19266,N_18128,N_18136);
xnor U19267 (N_19267,N_18529,N_18095);
and U19268 (N_19268,N_17572,N_18727);
nor U19269 (N_19269,N_17941,N_18715);
or U19270 (N_19270,N_17677,N_17503);
and U19271 (N_19271,N_18501,N_17637);
or U19272 (N_19272,N_17666,N_18424);
or U19273 (N_19273,N_17954,N_17690);
or U19274 (N_19274,N_17653,N_18041);
xnor U19275 (N_19275,N_18698,N_18049);
nor U19276 (N_19276,N_18009,N_18607);
or U19277 (N_19277,N_18321,N_17661);
and U19278 (N_19278,N_18220,N_17733);
and U19279 (N_19279,N_18141,N_17668);
nand U19280 (N_19280,N_18504,N_17792);
nand U19281 (N_19281,N_17837,N_17664);
or U19282 (N_19282,N_18629,N_17589);
and U19283 (N_19283,N_18177,N_18500);
or U19284 (N_19284,N_18171,N_18193);
or U19285 (N_19285,N_17667,N_18651);
xor U19286 (N_19286,N_18271,N_17629);
nor U19287 (N_19287,N_18108,N_18244);
nand U19288 (N_19288,N_18083,N_17744);
and U19289 (N_19289,N_17670,N_18617);
and U19290 (N_19290,N_18392,N_18105);
nand U19291 (N_19291,N_17949,N_17980);
nand U19292 (N_19292,N_17552,N_17695);
xor U19293 (N_19293,N_18034,N_18576);
xor U19294 (N_19294,N_18511,N_17590);
and U19295 (N_19295,N_17580,N_18647);
nand U19296 (N_19296,N_18316,N_18672);
nor U19297 (N_19297,N_18126,N_18132);
nor U19298 (N_19298,N_18520,N_18313);
nand U19299 (N_19299,N_18206,N_18692);
or U19300 (N_19300,N_17669,N_18628);
nand U19301 (N_19301,N_17931,N_17885);
xnor U19302 (N_19302,N_18004,N_17869);
and U19303 (N_19303,N_18361,N_17978);
and U19304 (N_19304,N_18721,N_18503);
nand U19305 (N_19305,N_18390,N_17730);
or U19306 (N_19306,N_18073,N_18652);
or U19307 (N_19307,N_17787,N_17918);
and U19308 (N_19308,N_17924,N_18675);
or U19309 (N_19309,N_17897,N_17964);
nor U19310 (N_19310,N_18292,N_17528);
or U19311 (N_19311,N_17622,N_18687);
nand U19312 (N_19312,N_17660,N_18454);
and U19313 (N_19313,N_18240,N_18446);
nand U19314 (N_19314,N_18482,N_17603);
xnor U19315 (N_19315,N_17525,N_18619);
nand U19316 (N_19316,N_18355,N_18174);
or U19317 (N_19317,N_18731,N_17785);
or U19318 (N_19318,N_17720,N_18550);
nor U19319 (N_19319,N_18686,N_18096);
or U19320 (N_19320,N_18749,N_17758);
xor U19321 (N_19321,N_18329,N_18540);
xnor U19322 (N_19322,N_18071,N_18696);
nor U19323 (N_19323,N_18059,N_18432);
nand U19324 (N_19324,N_17641,N_17836);
xor U19325 (N_19325,N_18018,N_17716);
nor U19326 (N_19326,N_17938,N_18506);
nor U19327 (N_19327,N_18470,N_18364);
and U19328 (N_19328,N_17609,N_17514);
xor U19329 (N_19329,N_18225,N_17559);
nand U19330 (N_19330,N_18738,N_17827);
and U19331 (N_19331,N_17861,N_18711);
nor U19332 (N_19332,N_17551,N_18069);
xnor U19333 (N_19333,N_18507,N_18260);
and U19334 (N_19334,N_18239,N_17901);
or U19335 (N_19335,N_17856,N_18373);
or U19336 (N_19336,N_18082,N_17539);
and U19337 (N_19337,N_18055,N_18363);
nand U19338 (N_19338,N_17919,N_17650);
or U19339 (N_19339,N_18042,N_18245);
nand U19340 (N_19340,N_18660,N_17823);
nand U19341 (N_19341,N_17598,N_17773);
and U19342 (N_19342,N_17530,N_18265);
nor U19343 (N_19343,N_18235,N_17584);
or U19344 (N_19344,N_18191,N_18613);
nor U19345 (N_19345,N_18624,N_18107);
and U19346 (N_19346,N_17703,N_18433);
and U19347 (N_19347,N_18724,N_18439);
or U19348 (N_19348,N_17540,N_17712);
and U19349 (N_19349,N_17523,N_17878);
nand U19350 (N_19350,N_17991,N_18104);
nand U19351 (N_19351,N_17752,N_17882);
nand U19352 (N_19352,N_18663,N_17830);
xor U19353 (N_19353,N_18123,N_17522);
nor U19354 (N_19354,N_17541,N_18527);
xor U19355 (N_19355,N_17989,N_18489);
and U19356 (N_19356,N_18572,N_18496);
nor U19357 (N_19357,N_18376,N_18377);
nor U19358 (N_19358,N_18290,N_18509);
or U19359 (N_19359,N_17966,N_17596);
nor U19360 (N_19360,N_18606,N_17708);
nand U19361 (N_19361,N_17849,N_17705);
nand U19362 (N_19362,N_18368,N_18114);
or U19363 (N_19363,N_18178,N_18399);
and U19364 (N_19364,N_18295,N_17546);
nor U19365 (N_19365,N_17678,N_18551);
xnor U19366 (N_19366,N_18583,N_17821);
xnor U19367 (N_19367,N_17697,N_17995);
and U19368 (N_19368,N_18553,N_18284);
and U19369 (N_19369,N_18464,N_18582);
nand U19370 (N_19370,N_17640,N_18475);
nand U19371 (N_19371,N_17888,N_17846);
or U19372 (N_19372,N_17884,N_17948);
nand U19373 (N_19373,N_18257,N_18485);
xnor U19374 (N_19374,N_17889,N_18534);
or U19375 (N_19375,N_17562,N_18516);
xnor U19376 (N_19376,N_18157,N_18441);
nor U19377 (N_19377,N_18692,N_18446);
nor U19378 (N_19378,N_17663,N_17703);
and U19379 (N_19379,N_18569,N_18541);
xor U19380 (N_19380,N_17502,N_18097);
nor U19381 (N_19381,N_18178,N_18734);
or U19382 (N_19382,N_18442,N_17661);
xnor U19383 (N_19383,N_17927,N_18141);
nand U19384 (N_19384,N_18051,N_18598);
nor U19385 (N_19385,N_18724,N_18298);
xor U19386 (N_19386,N_18253,N_18592);
or U19387 (N_19387,N_17616,N_17823);
nor U19388 (N_19388,N_17704,N_17657);
nor U19389 (N_19389,N_18443,N_18385);
xnor U19390 (N_19390,N_17997,N_17825);
nor U19391 (N_19391,N_18621,N_17823);
and U19392 (N_19392,N_17802,N_18709);
or U19393 (N_19393,N_18252,N_18715);
nand U19394 (N_19394,N_18038,N_18043);
or U19395 (N_19395,N_17822,N_18142);
nor U19396 (N_19396,N_18498,N_18401);
nor U19397 (N_19397,N_18109,N_18337);
nor U19398 (N_19398,N_18699,N_18036);
nor U19399 (N_19399,N_18545,N_17798);
nand U19400 (N_19400,N_17617,N_18573);
or U19401 (N_19401,N_17593,N_18443);
nand U19402 (N_19402,N_18318,N_18366);
and U19403 (N_19403,N_17737,N_18136);
and U19404 (N_19404,N_17887,N_17744);
nor U19405 (N_19405,N_18290,N_18341);
and U19406 (N_19406,N_18491,N_18381);
nand U19407 (N_19407,N_17860,N_18184);
nand U19408 (N_19408,N_17807,N_18474);
and U19409 (N_19409,N_18567,N_18211);
and U19410 (N_19410,N_17810,N_18247);
or U19411 (N_19411,N_18644,N_18297);
nand U19412 (N_19412,N_18535,N_18683);
or U19413 (N_19413,N_17958,N_18661);
and U19414 (N_19414,N_18656,N_17815);
or U19415 (N_19415,N_18414,N_18219);
nand U19416 (N_19416,N_18639,N_17723);
or U19417 (N_19417,N_18679,N_18291);
or U19418 (N_19418,N_18310,N_18573);
nand U19419 (N_19419,N_18118,N_18632);
nand U19420 (N_19420,N_18272,N_17780);
nand U19421 (N_19421,N_17666,N_17711);
xor U19422 (N_19422,N_17935,N_17719);
nand U19423 (N_19423,N_17544,N_17592);
and U19424 (N_19424,N_18711,N_18718);
nand U19425 (N_19425,N_17585,N_18675);
and U19426 (N_19426,N_18447,N_17574);
nand U19427 (N_19427,N_18079,N_17853);
and U19428 (N_19428,N_18520,N_17695);
nand U19429 (N_19429,N_18641,N_17528);
xor U19430 (N_19430,N_18151,N_17707);
xor U19431 (N_19431,N_18523,N_18702);
xnor U19432 (N_19432,N_18107,N_18400);
xor U19433 (N_19433,N_17892,N_18636);
and U19434 (N_19434,N_18605,N_17934);
and U19435 (N_19435,N_17821,N_17591);
xnor U19436 (N_19436,N_17619,N_18182);
xor U19437 (N_19437,N_17604,N_18431);
nand U19438 (N_19438,N_17523,N_18215);
or U19439 (N_19439,N_17883,N_17688);
and U19440 (N_19440,N_17800,N_18226);
and U19441 (N_19441,N_17585,N_18333);
nor U19442 (N_19442,N_18147,N_18698);
nor U19443 (N_19443,N_18009,N_17612);
or U19444 (N_19444,N_18325,N_18020);
nand U19445 (N_19445,N_18625,N_18326);
or U19446 (N_19446,N_18114,N_18296);
or U19447 (N_19447,N_17612,N_17598);
nor U19448 (N_19448,N_17669,N_17746);
and U19449 (N_19449,N_18620,N_17653);
or U19450 (N_19450,N_17549,N_17642);
nor U19451 (N_19451,N_18022,N_18605);
nor U19452 (N_19452,N_18699,N_17918);
nor U19453 (N_19453,N_18059,N_17817);
nor U19454 (N_19454,N_18250,N_18535);
nand U19455 (N_19455,N_18710,N_17537);
and U19456 (N_19456,N_17885,N_18031);
xor U19457 (N_19457,N_18398,N_18136);
nor U19458 (N_19458,N_17880,N_17995);
nor U19459 (N_19459,N_18135,N_18103);
nand U19460 (N_19460,N_18129,N_17575);
xnor U19461 (N_19461,N_17852,N_17891);
and U19462 (N_19462,N_17990,N_18690);
and U19463 (N_19463,N_17857,N_17509);
nor U19464 (N_19464,N_18143,N_18044);
or U19465 (N_19465,N_18351,N_17980);
or U19466 (N_19466,N_18696,N_17833);
or U19467 (N_19467,N_18329,N_18458);
nand U19468 (N_19468,N_18115,N_18152);
xnor U19469 (N_19469,N_18603,N_18366);
nor U19470 (N_19470,N_17784,N_18392);
nand U19471 (N_19471,N_18566,N_18668);
nand U19472 (N_19472,N_18618,N_17935);
nor U19473 (N_19473,N_18605,N_18076);
xor U19474 (N_19474,N_18503,N_18572);
xor U19475 (N_19475,N_18169,N_18275);
or U19476 (N_19476,N_17845,N_18381);
nor U19477 (N_19477,N_18679,N_18747);
and U19478 (N_19478,N_17970,N_17977);
nor U19479 (N_19479,N_18332,N_18079);
nand U19480 (N_19480,N_17754,N_17650);
or U19481 (N_19481,N_18289,N_18129);
and U19482 (N_19482,N_18368,N_18643);
and U19483 (N_19483,N_18011,N_17703);
xor U19484 (N_19484,N_18095,N_18550);
or U19485 (N_19485,N_18532,N_18710);
and U19486 (N_19486,N_18513,N_18368);
nor U19487 (N_19487,N_17746,N_18484);
or U19488 (N_19488,N_17800,N_17650);
and U19489 (N_19489,N_18051,N_18536);
nand U19490 (N_19490,N_18728,N_17666);
xor U19491 (N_19491,N_17860,N_17658);
nor U19492 (N_19492,N_18705,N_17881);
or U19493 (N_19493,N_18617,N_18120);
nor U19494 (N_19494,N_17938,N_18638);
nor U19495 (N_19495,N_17952,N_18066);
and U19496 (N_19496,N_17550,N_17640);
or U19497 (N_19497,N_18663,N_18342);
nor U19498 (N_19498,N_17644,N_17614);
xnor U19499 (N_19499,N_17983,N_18004);
nand U19500 (N_19500,N_17771,N_18258);
nor U19501 (N_19501,N_17997,N_17753);
or U19502 (N_19502,N_18706,N_18543);
xnor U19503 (N_19503,N_17519,N_18223);
nor U19504 (N_19504,N_17673,N_17875);
or U19505 (N_19505,N_17967,N_18200);
and U19506 (N_19506,N_18531,N_17588);
nor U19507 (N_19507,N_18324,N_18353);
or U19508 (N_19508,N_17563,N_17928);
xor U19509 (N_19509,N_18289,N_18419);
and U19510 (N_19510,N_18360,N_17853);
nor U19511 (N_19511,N_17966,N_18138);
or U19512 (N_19512,N_18571,N_18519);
and U19513 (N_19513,N_18513,N_17791);
and U19514 (N_19514,N_17767,N_17644);
nor U19515 (N_19515,N_18436,N_17568);
xnor U19516 (N_19516,N_17842,N_17567);
nor U19517 (N_19517,N_18631,N_18111);
and U19518 (N_19518,N_18585,N_18677);
nor U19519 (N_19519,N_17598,N_18620);
or U19520 (N_19520,N_17990,N_18074);
nor U19521 (N_19521,N_18214,N_17780);
and U19522 (N_19522,N_17704,N_17633);
nand U19523 (N_19523,N_18151,N_17781);
xnor U19524 (N_19524,N_17663,N_18167);
or U19525 (N_19525,N_17706,N_17521);
or U19526 (N_19526,N_18297,N_18100);
or U19527 (N_19527,N_18679,N_18052);
nand U19528 (N_19528,N_17849,N_18020);
nand U19529 (N_19529,N_17907,N_17596);
nor U19530 (N_19530,N_17549,N_17913);
xor U19531 (N_19531,N_18121,N_17585);
or U19532 (N_19532,N_18237,N_18368);
nand U19533 (N_19533,N_17755,N_18564);
nand U19534 (N_19534,N_18514,N_17788);
nor U19535 (N_19535,N_18168,N_17874);
xnor U19536 (N_19536,N_18743,N_18322);
nor U19537 (N_19537,N_18460,N_17964);
xnor U19538 (N_19538,N_17728,N_18033);
and U19539 (N_19539,N_18113,N_17619);
xor U19540 (N_19540,N_18447,N_18625);
and U19541 (N_19541,N_17923,N_17621);
and U19542 (N_19542,N_17647,N_18575);
nor U19543 (N_19543,N_17931,N_18278);
or U19544 (N_19544,N_17756,N_17684);
or U19545 (N_19545,N_18421,N_18286);
nand U19546 (N_19546,N_18009,N_17709);
and U19547 (N_19547,N_18659,N_17542);
nand U19548 (N_19548,N_18723,N_18161);
xor U19549 (N_19549,N_17666,N_18006);
or U19550 (N_19550,N_18518,N_18659);
xor U19551 (N_19551,N_18352,N_17500);
xor U19552 (N_19552,N_18616,N_18740);
xor U19553 (N_19553,N_18414,N_18040);
and U19554 (N_19554,N_18710,N_18275);
nor U19555 (N_19555,N_18609,N_18037);
xor U19556 (N_19556,N_17538,N_18717);
nor U19557 (N_19557,N_17531,N_17873);
or U19558 (N_19558,N_17946,N_17807);
xnor U19559 (N_19559,N_17952,N_18607);
or U19560 (N_19560,N_17790,N_18066);
nand U19561 (N_19561,N_18293,N_17654);
nand U19562 (N_19562,N_18530,N_18124);
nor U19563 (N_19563,N_18220,N_18230);
and U19564 (N_19564,N_18531,N_17957);
and U19565 (N_19565,N_18280,N_18261);
and U19566 (N_19566,N_18371,N_18314);
and U19567 (N_19567,N_18468,N_18035);
xnor U19568 (N_19568,N_18122,N_18627);
nor U19569 (N_19569,N_18640,N_18445);
xnor U19570 (N_19570,N_17851,N_17899);
nand U19571 (N_19571,N_18544,N_18420);
and U19572 (N_19572,N_18574,N_18700);
and U19573 (N_19573,N_18682,N_17658);
and U19574 (N_19574,N_18640,N_18639);
xor U19575 (N_19575,N_18274,N_18052);
and U19576 (N_19576,N_17569,N_17882);
or U19577 (N_19577,N_18551,N_17637);
nor U19578 (N_19578,N_17719,N_18159);
xnor U19579 (N_19579,N_18439,N_17505);
xor U19580 (N_19580,N_17910,N_18019);
nand U19581 (N_19581,N_18650,N_18533);
nor U19582 (N_19582,N_18119,N_17558);
nand U19583 (N_19583,N_18189,N_18643);
xor U19584 (N_19584,N_18640,N_18225);
or U19585 (N_19585,N_17715,N_18747);
nor U19586 (N_19586,N_17744,N_18036);
or U19587 (N_19587,N_18338,N_18524);
and U19588 (N_19588,N_17786,N_18297);
xnor U19589 (N_19589,N_17913,N_18467);
and U19590 (N_19590,N_18031,N_17585);
nand U19591 (N_19591,N_18582,N_18611);
or U19592 (N_19592,N_17500,N_18575);
and U19593 (N_19593,N_17743,N_18727);
nor U19594 (N_19594,N_17983,N_17642);
or U19595 (N_19595,N_18215,N_17862);
or U19596 (N_19596,N_18457,N_17526);
nor U19597 (N_19597,N_18359,N_18425);
nor U19598 (N_19598,N_18550,N_17961);
and U19599 (N_19599,N_18415,N_17916);
or U19600 (N_19600,N_18634,N_18573);
or U19601 (N_19601,N_17965,N_18183);
xor U19602 (N_19602,N_17701,N_18394);
and U19603 (N_19603,N_17777,N_18646);
or U19604 (N_19604,N_17722,N_18164);
nand U19605 (N_19605,N_18164,N_17686);
or U19606 (N_19606,N_18219,N_18689);
nand U19607 (N_19607,N_17994,N_17726);
nor U19608 (N_19608,N_17778,N_17751);
or U19609 (N_19609,N_17580,N_18658);
nor U19610 (N_19610,N_18622,N_17500);
or U19611 (N_19611,N_18727,N_18310);
or U19612 (N_19612,N_18384,N_17812);
nor U19613 (N_19613,N_18022,N_18393);
and U19614 (N_19614,N_18067,N_17748);
nor U19615 (N_19615,N_17516,N_18229);
nor U19616 (N_19616,N_17688,N_17879);
nor U19617 (N_19617,N_18599,N_18521);
nor U19618 (N_19618,N_17990,N_18384);
nor U19619 (N_19619,N_18671,N_18662);
and U19620 (N_19620,N_18441,N_18317);
and U19621 (N_19621,N_17839,N_18311);
nor U19622 (N_19622,N_18341,N_18554);
nand U19623 (N_19623,N_17861,N_18086);
nor U19624 (N_19624,N_18177,N_18027);
nor U19625 (N_19625,N_17853,N_18406);
xnor U19626 (N_19626,N_18446,N_18177);
xor U19627 (N_19627,N_17598,N_18656);
or U19628 (N_19628,N_17763,N_17708);
nor U19629 (N_19629,N_18362,N_17919);
and U19630 (N_19630,N_17503,N_18616);
xor U19631 (N_19631,N_18625,N_18565);
or U19632 (N_19632,N_18159,N_18570);
or U19633 (N_19633,N_18532,N_18410);
or U19634 (N_19634,N_17649,N_17552);
xnor U19635 (N_19635,N_18631,N_17675);
nand U19636 (N_19636,N_18514,N_17660);
or U19637 (N_19637,N_17803,N_17790);
nor U19638 (N_19638,N_17731,N_18005);
nand U19639 (N_19639,N_18454,N_17524);
xnor U19640 (N_19640,N_17996,N_18626);
and U19641 (N_19641,N_18490,N_18150);
and U19642 (N_19642,N_17720,N_18224);
nor U19643 (N_19643,N_17505,N_17739);
and U19644 (N_19644,N_18098,N_18095);
nor U19645 (N_19645,N_18652,N_17884);
or U19646 (N_19646,N_18686,N_18256);
and U19647 (N_19647,N_17524,N_18364);
nor U19648 (N_19648,N_17677,N_17566);
and U19649 (N_19649,N_18284,N_18079);
xor U19650 (N_19650,N_17848,N_18701);
xnor U19651 (N_19651,N_18460,N_18398);
xor U19652 (N_19652,N_18707,N_17877);
and U19653 (N_19653,N_18448,N_18601);
xnor U19654 (N_19654,N_18587,N_17967);
and U19655 (N_19655,N_17677,N_18704);
nor U19656 (N_19656,N_18467,N_18326);
nor U19657 (N_19657,N_17833,N_17790);
xor U19658 (N_19658,N_18284,N_17765);
and U19659 (N_19659,N_18430,N_17785);
and U19660 (N_19660,N_18511,N_17739);
and U19661 (N_19661,N_18136,N_18056);
and U19662 (N_19662,N_18282,N_17534);
and U19663 (N_19663,N_18404,N_17835);
xor U19664 (N_19664,N_18605,N_17769);
nor U19665 (N_19665,N_17970,N_18245);
nor U19666 (N_19666,N_18591,N_17572);
or U19667 (N_19667,N_18042,N_18351);
or U19668 (N_19668,N_17621,N_18148);
or U19669 (N_19669,N_18442,N_18168);
and U19670 (N_19670,N_18515,N_17509);
xor U19671 (N_19671,N_17639,N_17874);
or U19672 (N_19672,N_18739,N_18401);
xnor U19673 (N_19673,N_18655,N_17740);
or U19674 (N_19674,N_18596,N_18665);
or U19675 (N_19675,N_18081,N_18697);
nand U19676 (N_19676,N_18166,N_17709);
nor U19677 (N_19677,N_18390,N_17921);
or U19678 (N_19678,N_17748,N_18163);
nand U19679 (N_19679,N_18260,N_17577);
and U19680 (N_19680,N_18407,N_18213);
or U19681 (N_19681,N_18614,N_18063);
xor U19682 (N_19682,N_18317,N_17660);
and U19683 (N_19683,N_18267,N_18607);
nand U19684 (N_19684,N_18668,N_18418);
or U19685 (N_19685,N_18726,N_18376);
nand U19686 (N_19686,N_18430,N_18104);
or U19687 (N_19687,N_17872,N_17918);
nor U19688 (N_19688,N_18395,N_18341);
nand U19689 (N_19689,N_17819,N_18142);
and U19690 (N_19690,N_17530,N_17994);
nor U19691 (N_19691,N_17979,N_18634);
and U19692 (N_19692,N_17833,N_17682);
xnor U19693 (N_19693,N_17954,N_18633);
nand U19694 (N_19694,N_18578,N_18387);
or U19695 (N_19695,N_18135,N_18054);
or U19696 (N_19696,N_17985,N_18007);
or U19697 (N_19697,N_17672,N_17596);
xor U19698 (N_19698,N_17745,N_18299);
nand U19699 (N_19699,N_18516,N_18739);
and U19700 (N_19700,N_18365,N_17597);
nand U19701 (N_19701,N_17671,N_18531);
nand U19702 (N_19702,N_18718,N_18633);
and U19703 (N_19703,N_18738,N_18256);
and U19704 (N_19704,N_17613,N_17899);
or U19705 (N_19705,N_18354,N_18316);
or U19706 (N_19706,N_18270,N_18113);
nor U19707 (N_19707,N_17889,N_17828);
or U19708 (N_19708,N_18172,N_17550);
xor U19709 (N_19709,N_18153,N_17542);
xor U19710 (N_19710,N_18028,N_18073);
xor U19711 (N_19711,N_17977,N_17915);
nor U19712 (N_19712,N_18718,N_18332);
nor U19713 (N_19713,N_18269,N_18338);
or U19714 (N_19714,N_18117,N_18682);
nand U19715 (N_19715,N_18238,N_17568);
or U19716 (N_19716,N_18715,N_18262);
nand U19717 (N_19717,N_17767,N_17979);
nor U19718 (N_19718,N_18114,N_17839);
and U19719 (N_19719,N_18603,N_17836);
nand U19720 (N_19720,N_18233,N_18606);
or U19721 (N_19721,N_18255,N_17904);
nand U19722 (N_19722,N_18681,N_18374);
xor U19723 (N_19723,N_17517,N_18653);
xnor U19724 (N_19724,N_18185,N_18037);
xor U19725 (N_19725,N_17986,N_18689);
nand U19726 (N_19726,N_18411,N_17598);
xnor U19727 (N_19727,N_17785,N_18402);
or U19728 (N_19728,N_17794,N_18538);
nand U19729 (N_19729,N_18183,N_18608);
and U19730 (N_19730,N_18169,N_17568);
or U19731 (N_19731,N_18435,N_18315);
and U19732 (N_19732,N_17869,N_17637);
xor U19733 (N_19733,N_17606,N_17803);
and U19734 (N_19734,N_18072,N_17769);
xor U19735 (N_19735,N_18566,N_18403);
nand U19736 (N_19736,N_18597,N_18730);
nor U19737 (N_19737,N_17715,N_18374);
nand U19738 (N_19738,N_18723,N_17999);
xor U19739 (N_19739,N_18666,N_18242);
and U19740 (N_19740,N_17867,N_18560);
nor U19741 (N_19741,N_18650,N_18439);
and U19742 (N_19742,N_18433,N_17906);
or U19743 (N_19743,N_18179,N_17679);
nor U19744 (N_19744,N_18443,N_18326);
nand U19745 (N_19745,N_17623,N_17830);
or U19746 (N_19746,N_18195,N_17723);
or U19747 (N_19747,N_17702,N_18448);
xor U19748 (N_19748,N_17946,N_17512);
or U19749 (N_19749,N_18308,N_18550);
nor U19750 (N_19750,N_18006,N_18225);
nor U19751 (N_19751,N_18401,N_18507);
nor U19752 (N_19752,N_18714,N_17762);
nor U19753 (N_19753,N_18584,N_18148);
and U19754 (N_19754,N_18200,N_18037);
xor U19755 (N_19755,N_18689,N_18020);
xor U19756 (N_19756,N_17821,N_18225);
nor U19757 (N_19757,N_18230,N_18088);
nor U19758 (N_19758,N_18294,N_17810);
or U19759 (N_19759,N_17985,N_18410);
xnor U19760 (N_19760,N_18587,N_17995);
nand U19761 (N_19761,N_17999,N_17640);
xnor U19762 (N_19762,N_17565,N_18520);
or U19763 (N_19763,N_18660,N_18445);
nor U19764 (N_19764,N_18490,N_18175);
nor U19765 (N_19765,N_18643,N_18064);
xor U19766 (N_19766,N_18551,N_18716);
and U19767 (N_19767,N_17678,N_18685);
or U19768 (N_19768,N_17651,N_18303);
xnor U19769 (N_19769,N_18665,N_18611);
or U19770 (N_19770,N_17604,N_18182);
xor U19771 (N_19771,N_17808,N_17714);
nand U19772 (N_19772,N_18575,N_18025);
xnor U19773 (N_19773,N_18631,N_18653);
nor U19774 (N_19774,N_17642,N_18356);
or U19775 (N_19775,N_18251,N_17836);
xnor U19776 (N_19776,N_18115,N_17565);
nor U19777 (N_19777,N_17934,N_18749);
or U19778 (N_19778,N_18527,N_17872);
and U19779 (N_19779,N_18225,N_17591);
and U19780 (N_19780,N_18152,N_17725);
and U19781 (N_19781,N_18613,N_18392);
or U19782 (N_19782,N_17763,N_17654);
nand U19783 (N_19783,N_17843,N_17601);
nand U19784 (N_19784,N_18276,N_17819);
nor U19785 (N_19785,N_17553,N_17798);
or U19786 (N_19786,N_17924,N_18035);
or U19787 (N_19787,N_17777,N_18634);
and U19788 (N_19788,N_17840,N_17745);
xnor U19789 (N_19789,N_17591,N_17515);
nor U19790 (N_19790,N_18316,N_18104);
nand U19791 (N_19791,N_18570,N_17931);
nand U19792 (N_19792,N_18731,N_18293);
or U19793 (N_19793,N_17785,N_18524);
and U19794 (N_19794,N_17714,N_17583);
xor U19795 (N_19795,N_18124,N_18157);
nor U19796 (N_19796,N_17825,N_18205);
and U19797 (N_19797,N_17521,N_17859);
nor U19798 (N_19798,N_18607,N_18481);
nand U19799 (N_19799,N_17884,N_17867);
xor U19800 (N_19800,N_18354,N_18398);
or U19801 (N_19801,N_18491,N_17852);
or U19802 (N_19802,N_18621,N_17805);
nand U19803 (N_19803,N_18251,N_17670);
nor U19804 (N_19804,N_18455,N_18610);
nor U19805 (N_19805,N_18533,N_18611);
xnor U19806 (N_19806,N_18176,N_18637);
nand U19807 (N_19807,N_18312,N_17994);
xor U19808 (N_19808,N_17643,N_18285);
nor U19809 (N_19809,N_17663,N_18356);
and U19810 (N_19810,N_17811,N_17584);
and U19811 (N_19811,N_18201,N_18419);
nand U19812 (N_19812,N_17802,N_17945);
nor U19813 (N_19813,N_18514,N_18352);
nand U19814 (N_19814,N_18260,N_17883);
nand U19815 (N_19815,N_18615,N_17531);
nand U19816 (N_19816,N_18582,N_18055);
nand U19817 (N_19817,N_18644,N_18273);
or U19818 (N_19818,N_18306,N_18363);
nand U19819 (N_19819,N_18168,N_18071);
nor U19820 (N_19820,N_18233,N_18388);
nor U19821 (N_19821,N_18435,N_18390);
and U19822 (N_19822,N_18380,N_18198);
or U19823 (N_19823,N_18085,N_18026);
xnor U19824 (N_19824,N_17631,N_17624);
and U19825 (N_19825,N_18152,N_17970);
xor U19826 (N_19826,N_17711,N_18024);
nand U19827 (N_19827,N_17573,N_17680);
nor U19828 (N_19828,N_18230,N_17535);
or U19829 (N_19829,N_18535,N_18001);
nand U19830 (N_19830,N_17915,N_18307);
nor U19831 (N_19831,N_18601,N_18199);
nand U19832 (N_19832,N_17803,N_18448);
nand U19833 (N_19833,N_18557,N_17521);
nor U19834 (N_19834,N_18492,N_17882);
xnor U19835 (N_19835,N_17500,N_18533);
nor U19836 (N_19836,N_17688,N_17825);
xnor U19837 (N_19837,N_18714,N_18474);
or U19838 (N_19838,N_18251,N_18100);
and U19839 (N_19839,N_17538,N_18065);
or U19840 (N_19840,N_17542,N_18513);
xor U19841 (N_19841,N_18353,N_18560);
and U19842 (N_19842,N_18419,N_17504);
xnor U19843 (N_19843,N_18212,N_18706);
and U19844 (N_19844,N_17586,N_18013);
or U19845 (N_19845,N_18199,N_18502);
nand U19846 (N_19846,N_18670,N_18180);
nor U19847 (N_19847,N_17606,N_18571);
xnor U19848 (N_19848,N_18083,N_17632);
xor U19849 (N_19849,N_18691,N_17879);
nor U19850 (N_19850,N_17662,N_18718);
and U19851 (N_19851,N_18271,N_18453);
xor U19852 (N_19852,N_18326,N_18379);
and U19853 (N_19853,N_18507,N_18057);
or U19854 (N_19854,N_18687,N_17999);
or U19855 (N_19855,N_17935,N_17777);
xnor U19856 (N_19856,N_17624,N_17678);
and U19857 (N_19857,N_17859,N_17636);
nor U19858 (N_19858,N_18721,N_18628);
or U19859 (N_19859,N_18101,N_17956);
nor U19860 (N_19860,N_18689,N_18052);
xor U19861 (N_19861,N_17955,N_18586);
or U19862 (N_19862,N_18322,N_17595);
nor U19863 (N_19863,N_18702,N_18342);
or U19864 (N_19864,N_17946,N_18706);
nor U19865 (N_19865,N_18140,N_18365);
nand U19866 (N_19866,N_17851,N_18239);
nor U19867 (N_19867,N_17593,N_18659);
xnor U19868 (N_19868,N_18272,N_17579);
nor U19869 (N_19869,N_17583,N_17882);
xor U19870 (N_19870,N_17932,N_18703);
nand U19871 (N_19871,N_17627,N_18253);
nand U19872 (N_19872,N_18140,N_17624);
nor U19873 (N_19873,N_17954,N_17559);
and U19874 (N_19874,N_18644,N_18280);
xnor U19875 (N_19875,N_18451,N_17738);
nand U19876 (N_19876,N_18233,N_17926);
nor U19877 (N_19877,N_18601,N_18139);
nor U19878 (N_19878,N_17895,N_18305);
xnor U19879 (N_19879,N_17725,N_18494);
nor U19880 (N_19880,N_18579,N_17904);
and U19881 (N_19881,N_18673,N_17991);
or U19882 (N_19882,N_18014,N_17528);
nor U19883 (N_19883,N_18360,N_17943);
xor U19884 (N_19884,N_17767,N_17585);
or U19885 (N_19885,N_18182,N_18467);
and U19886 (N_19886,N_18516,N_18521);
nor U19887 (N_19887,N_18364,N_17556);
xor U19888 (N_19888,N_18335,N_18701);
nand U19889 (N_19889,N_18243,N_18535);
nor U19890 (N_19890,N_18636,N_18745);
nor U19891 (N_19891,N_17636,N_18334);
nand U19892 (N_19892,N_18530,N_17563);
xnor U19893 (N_19893,N_17995,N_18609);
nor U19894 (N_19894,N_17832,N_18671);
xnor U19895 (N_19895,N_18294,N_17938);
xnor U19896 (N_19896,N_18202,N_17819);
and U19897 (N_19897,N_17922,N_17893);
or U19898 (N_19898,N_17576,N_18426);
nand U19899 (N_19899,N_18369,N_18033);
nand U19900 (N_19900,N_18210,N_17891);
and U19901 (N_19901,N_18353,N_18300);
and U19902 (N_19902,N_18004,N_17534);
xnor U19903 (N_19903,N_17603,N_17615);
xnor U19904 (N_19904,N_18071,N_18187);
xnor U19905 (N_19905,N_18597,N_17626);
or U19906 (N_19906,N_18167,N_18039);
or U19907 (N_19907,N_17759,N_18192);
nand U19908 (N_19908,N_17818,N_18591);
and U19909 (N_19909,N_18442,N_18229);
nand U19910 (N_19910,N_17744,N_17937);
and U19911 (N_19911,N_18584,N_17620);
nor U19912 (N_19912,N_18533,N_18310);
nand U19913 (N_19913,N_17778,N_17858);
nor U19914 (N_19914,N_17972,N_17523);
and U19915 (N_19915,N_17802,N_18592);
and U19916 (N_19916,N_17644,N_18251);
nand U19917 (N_19917,N_17527,N_18326);
xnor U19918 (N_19918,N_17893,N_17998);
nand U19919 (N_19919,N_18694,N_17906);
xnor U19920 (N_19920,N_18032,N_18402);
xnor U19921 (N_19921,N_17944,N_18738);
xor U19922 (N_19922,N_17874,N_17652);
xor U19923 (N_19923,N_17538,N_17761);
and U19924 (N_19924,N_18023,N_17999);
nor U19925 (N_19925,N_17784,N_18158);
or U19926 (N_19926,N_18669,N_18328);
xnor U19927 (N_19927,N_17587,N_17964);
or U19928 (N_19928,N_18430,N_17897);
and U19929 (N_19929,N_18742,N_18666);
nor U19930 (N_19930,N_18352,N_18603);
and U19931 (N_19931,N_17741,N_18560);
and U19932 (N_19932,N_18327,N_17833);
or U19933 (N_19933,N_18631,N_18322);
xnor U19934 (N_19934,N_18492,N_17580);
nand U19935 (N_19935,N_17552,N_18550);
or U19936 (N_19936,N_17577,N_18007);
nand U19937 (N_19937,N_17691,N_18146);
or U19938 (N_19938,N_17789,N_17579);
nand U19939 (N_19939,N_18324,N_18605);
nand U19940 (N_19940,N_17590,N_18231);
nand U19941 (N_19941,N_17507,N_18419);
or U19942 (N_19942,N_17887,N_17576);
nor U19943 (N_19943,N_18658,N_18019);
or U19944 (N_19944,N_18703,N_18307);
or U19945 (N_19945,N_18541,N_18229);
nand U19946 (N_19946,N_17813,N_18736);
xor U19947 (N_19947,N_17968,N_17552);
xnor U19948 (N_19948,N_17531,N_17923);
and U19949 (N_19949,N_18724,N_18207);
nand U19950 (N_19950,N_18318,N_18616);
and U19951 (N_19951,N_18336,N_17963);
nor U19952 (N_19952,N_17884,N_18692);
nand U19953 (N_19953,N_17884,N_17659);
xnor U19954 (N_19954,N_17887,N_17817);
nor U19955 (N_19955,N_18609,N_18001);
nor U19956 (N_19956,N_18614,N_17810);
nand U19957 (N_19957,N_17832,N_18539);
or U19958 (N_19958,N_17509,N_18677);
or U19959 (N_19959,N_18018,N_17547);
nor U19960 (N_19960,N_18464,N_17809);
and U19961 (N_19961,N_17619,N_18279);
or U19962 (N_19962,N_17598,N_18415);
xor U19963 (N_19963,N_17804,N_17521);
nand U19964 (N_19964,N_17782,N_18282);
and U19965 (N_19965,N_18073,N_17990);
and U19966 (N_19966,N_18579,N_18285);
or U19967 (N_19967,N_17584,N_18442);
xor U19968 (N_19968,N_18093,N_17629);
nor U19969 (N_19969,N_18485,N_18083);
or U19970 (N_19970,N_18223,N_17583);
or U19971 (N_19971,N_17848,N_17531);
nand U19972 (N_19972,N_17853,N_18724);
nand U19973 (N_19973,N_18567,N_18723);
nand U19974 (N_19974,N_17821,N_18234);
and U19975 (N_19975,N_17682,N_17936);
or U19976 (N_19976,N_18112,N_17914);
nand U19977 (N_19977,N_18226,N_17705);
nor U19978 (N_19978,N_18687,N_18543);
or U19979 (N_19979,N_18659,N_18363);
or U19980 (N_19980,N_18665,N_18306);
nand U19981 (N_19981,N_17815,N_18661);
and U19982 (N_19982,N_17658,N_17850);
nor U19983 (N_19983,N_18672,N_18600);
nor U19984 (N_19984,N_17888,N_18174);
nor U19985 (N_19985,N_18247,N_17612);
nor U19986 (N_19986,N_18289,N_17748);
nand U19987 (N_19987,N_17839,N_18557);
xnor U19988 (N_19988,N_18313,N_18242);
or U19989 (N_19989,N_17777,N_18563);
or U19990 (N_19990,N_18231,N_17694);
nand U19991 (N_19991,N_17820,N_17960);
nor U19992 (N_19992,N_18307,N_18336);
and U19993 (N_19993,N_18235,N_17625);
xor U19994 (N_19994,N_17866,N_17758);
nor U19995 (N_19995,N_17980,N_18073);
and U19996 (N_19996,N_17831,N_18244);
and U19997 (N_19997,N_18672,N_17954);
nand U19998 (N_19998,N_18422,N_18424);
nand U19999 (N_19999,N_17962,N_18480);
nor U20000 (N_20000,N_19389,N_19255);
xor U20001 (N_20001,N_19239,N_19332);
or U20002 (N_20002,N_19369,N_19230);
nand U20003 (N_20003,N_19450,N_19031);
xnor U20004 (N_20004,N_19334,N_19392);
and U20005 (N_20005,N_19754,N_19678);
and U20006 (N_20006,N_18955,N_19335);
and U20007 (N_20007,N_19275,N_19337);
and U20008 (N_20008,N_19220,N_18965);
and U20009 (N_20009,N_19246,N_18996);
or U20010 (N_20010,N_19304,N_19322);
xor U20011 (N_20011,N_19157,N_19697);
nor U20012 (N_20012,N_19643,N_19736);
xor U20013 (N_20013,N_19807,N_19412);
or U20014 (N_20014,N_19738,N_19829);
or U20015 (N_20015,N_19933,N_19018);
xnor U20016 (N_20016,N_19600,N_19805);
nand U20017 (N_20017,N_19478,N_19890);
or U20018 (N_20018,N_19323,N_19070);
or U20019 (N_20019,N_19102,N_18888);
xor U20020 (N_20020,N_19289,N_18837);
nor U20021 (N_20021,N_19459,N_19139);
and U20022 (N_20022,N_19276,N_19202);
nor U20023 (N_20023,N_19366,N_19005);
nor U20024 (N_20024,N_19204,N_19346);
xor U20025 (N_20025,N_19147,N_19143);
nor U20026 (N_20026,N_19720,N_19299);
or U20027 (N_20027,N_19419,N_19923);
and U20028 (N_20028,N_19254,N_19685);
xor U20029 (N_20029,N_18905,N_19307);
xor U20030 (N_20030,N_19101,N_18854);
xnor U20031 (N_20031,N_19229,N_19327);
nand U20032 (N_20032,N_19818,N_19528);
nand U20033 (N_20033,N_19513,N_19690);
or U20034 (N_20034,N_18946,N_19792);
xor U20035 (N_20035,N_19042,N_19047);
nand U20036 (N_20036,N_19111,N_19226);
xnor U20037 (N_20037,N_19290,N_18917);
or U20038 (N_20038,N_18761,N_19559);
or U20039 (N_20039,N_19415,N_19509);
nand U20040 (N_20040,N_19691,N_19352);
xor U20041 (N_20041,N_19131,N_18977);
nor U20042 (N_20042,N_19731,N_18921);
nand U20043 (N_20043,N_19223,N_19595);
and U20044 (N_20044,N_19750,N_19721);
nor U20045 (N_20045,N_19809,N_19273);
nor U20046 (N_20046,N_19693,N_18932);
xor U20047 (N_20047,N_18887,N_19155);
and U20048 (N_20048,N_19524,N_19427);
nand U20049 (N_20049,N_19786,N_18832);
nand U20050 (N_20050,N_19329,N_18980);
xor U20051 (N_20051,N_19455,N_19873);
and U20052 (N_20052,N_19120,N_19616);
xnor U20053 (N_20053,N_18766,N_19837);
xnor U20054 (N_20054,N_19309,N_18864);
and U20055 (N_20055,N_19638,N_19705);
nor U20056 (N_20056,N_19916,N_19030);
xor U20057 (N_20057,N_19572,N_19312);
nand U20058 (N_20058,N_19972,N_19663);
nand U20059 (N_20059,N_19056,N_19394);
xor U20060 (N_20060,N_18850,N_19353);
or U20061 (N_20061,N_19773,N_19826);
nor U20062 (N_20062,N_18762,N_19507);
xnor U20063 (N_20063,N_19090,N_19103);
and U20064 (N_20064,N_19902,N_19986);
and U20065 (N_20065,N_19015,N_19946);
nor U20066 (N_20066,N_19939,N_19040);
and U20067 (N_20067,N_19658,N_18943);
and U20068 (N_20068,N_19451,N_19424);
nor U20069 (N_20069,N_19183,N_19876);
nand U20070 (N_20070,N_19683,N_18782);
and U20071 (N_20071,N_18776,N_19556);
xor U20072 (N_20072,N_19579,N_19426);
or U20073 (N_20073,N_18990,N_19875);
nand U20074 (N_20074,N_19935,N_18807);
xor U20075 (N_20075,N_19900,N_19248);
and U20076 (N_20076,N_19659,N_19196);
xor U20077 (N_20077,N_19035,N_19630);
xnor U20078 (N_20078,N_19860,N_18803);
and U20079 (N_20079,N_18781,N_19766);
xor U20080 (N_20080,N_19717,N_19043);
xnor U20081 (N_20081,N_19341,N_19260);
xnor U20082 (N_20082,N_19649,N_19184);
xnor U20083 (N_20083,N_19644,N_19227);
xnor U20084 (N_20084,N_19729,N_19636);
and U20085 (N_20085,N_18814,N_19944);
and U20086 (N_20086,N_19533,N_19167);
nand U20087 (N_20087,N_19375,N_19862);
and U20088 (N_20088,N_18936,N_19606);
or U20089 (N_20089,N_18755,N_19990);
and U20090 (N_20090,N_19793,N_19883);
and U20091 (N_20091,N_19970,N_18871);
xor U20092 (N_20092,N_18906,N_19368);
and U20093 (N_20093,N_19719,N_19381);
nor U20094 (N_20094,N_19365,N_19874);
or U20095 (N_20095,N_19940,N_18994);
nor U20096 (N_20096,N_19903,N_19665);
xor U20097 (N_20097,N_18999,N_19980);
xor U20098 (N_20098,N_19495,N_19431);
nand U20099 (N_20099,N_19951,N_19350);
xor U20100 (N_20100,N_19882,N_19928);
or U20101 (N_20101,N_19564,N_19124);
xnor U20102 (N_20102,N_19261,N_19593);
or U20103 (N_20103,N_19727,N_19010);
xnor U20104 (N_20104,N_18752,N_18912);
xor U20105 (N_20105,N_19992,N_19132);
nand U20106 (N_20106,N_19544,N_19856);
nor U20107 (N_20107,N_18821,N_18885);
nor U20108 (N_20108,N_19168,N_19002);
nor U20109 (N_20109,N_18892,N_19075);
nand U20110 (N_20110,N_19583,N_18792);
and U20111 (N_20111,N_18858,N_19608);
xnor U20112 (N_20112,N_19123,N_18979);
nor U20113 (N_20113,N_19137,N_19263);
xor U20114 (N_20114,N_19574,N_19121);
and U20115 (N_20115,N_19619,N_18900);
nand U20116 (N_20116,N_18904,N_19728);
nand U20117 (N_20117,N_19791,N_19479);
nand U20118 (N_20118,N_19449,N_19680);
or U20119 (N_20119,N_19483,N_19588);
xor U20120 (N_20120,N_19490,N_19804);
xnor U20121 (N_20121,N_19404,N_19073);
and U20122 (N_20122,N_19406,N_19247);
or U20123 (N_20123,N_18899,N_18795);
or U20124 (N_20124,N_19019,N_18750);
or U20125 (N_20125,N_19843,N_18877);
nor U20126 (N_20126,N_19909,N_19169);
xor U20127 (N_20127,N_19704,N_18929);
nor U20128 (N_20128,N_18954,N_19840);
nor U20129 (N_20129,N_19417,N_19497);
or U20130 (N_20130,N_19711,N_18879);
nor U20131 (N_20131,N_19821,N_19461);
nor U20132 (N_20132,N_19503,N_18827);
nor U20133 (N_20133,N_19354,N_18866);
and U20134 (N_20134,N_19844,N_18831);
or U20135 (N_20135,N_19812,N_19053);
or U20136 (N_20136,N_18890,N_19112);
nor U20137 (N_20137,N_19995,N_19250);
and U20138 (N_20138,N_19245,N_19560);
xnor U20139 (N_20139,N_19962,N_18845);
xor U20140 (N_20140,N_19025,N_19079);
nor U20141 (N_20141,N_19141,N_18819);
xor U20142 (N_20142,N_19652,N_19463);
xnor U20143 (N_20143,N_19795,N_19577);
nor U20144 (N_20144,N_19531,N_19587);
and U20145 (N_20145,N_18889,N_18869);
xor U20146 (N_20146,N_19489,N_19235);
nand U20147 (N_20147,N_19502,N_19877);
and U20148 (N_20148,N_19470,N_19618);
xnor U20149 (N_20149,N_19467,N_19447);
or U20150 (N_20150,N_19475,N_19893);
xnor U20151 (N_20151,N_18909,N_19632);
nor U20152 (N_20152,N_19622,N_19725);
nor U20153 (N_20153,N_19597,N_19477);
nand U20154 (N_20154,N_19642,N_18896);
nand U20155 (N_20155,N_19095,N_19562);
nand U20156 (N_20156,N_19405,N_19565);
xnor U20157 (N_20157,N_19243,N_19107);
xnor U20158 (N_20158,N_19772,N_18984);
or U20159 (N_20159,N_19889,N_18779);
nand U20160 (N_20160,N_18823,N_19561);
nand U20161 (N_20161,N_19615,N_19915);
nand U20162 (N_20162,N_19592,N_18964);
xor U20163 (N_20163,N_19244,N_19960);
or U20164 (N_20164,N_19491,N_19538);
nor U20165 (N_20165,N_18930,N_18815);
and U20166 (N_20166,N_18966,N_19868);
and U20167 (N_20167,N_19092,N_19534);
xor U20168 (N_20168,N_19819,N_19320);
nand U20169 (N_20169,N_19262,N_19769);
nand U20170 (N_20170,N_19129,N_19468);
xor U20171 (N_20171,N_18751,N_18811);
or U20172 (N_20172,N_19362,N_19788);
xnor U20173 (N_20173,N_18962,N_18852);
xor U20174 (N_20174,N_19462,N_19539);
or U20175 (N_20175,N_19482,N_19096);
xnor U20176 (N_20176,N_19492,N_19037);
and U20177 (N_20177,N_19781,N_18957);
nand U20178 (N_20178,N_19435,N_19080);
and U20179 (N_20179,N_19954,N_19249);
nor U20180 (N_20180,N_18956,N_18771);
nor U20181 (N_20181,N_19127,N_19861);
or U20182 (N_20182,N_19283,N_18758);
and U20183 (N_20183,N_19237,N_19985);
and U20184 (N_20184,N_19535,N_19589);
or U20185 (N_20185,N_19661,N_19373);
nand U20186 (N_20186,N_19163,N_18788);
xor U20187 (N_20187,N_19760,N_19385);
xnor U20188 (N_20188,N_19013,N_19755);
and U20189 (N_20189,N_19317,N_19514);
or U20190 (N_20190,N_19150,N_19635);
xnor U20191 (N_20191,N_19679,N_19747);
nand U20192 (N_20192,N_18881,N_19917);
or U20193 (N_20193,N_19824,N_18993);
nand U20194 (N_20194,N_19950,N_19776);
or U20195 (N_20195,N_19241,N_18953);
xor U20196 (N_20196,N_19498,N_19225);
xor U20197 (N_20197,N_19400,N_18836);
or U20198 (N_20198,N_19425,N_18790);
xnor U20199 (N_20199,N_19599,N_18798);
or U20200 (N_20200,N_19052,N_19575);
and U20201 (N_20201,N_18987,N_19886);
or U20202 (N_20202,N_19897,N_19325);
nor U20203 (N_20203,N_19541,N_19801);
nand U20204 (N_20204,N_19333,N_19188);
nand U20205 (N_20205,N_19789,N_19082);
nand U20206 (N_20206,N_19743,N_19759);
nor U20207 (N_20207,N_19854,N_19446);
or U20208 (N_20208,N_19519,N_18995);
nor U20209 (N_20209,N_19292,N_18915);
nand U20210 (N_20210,N_19997,N_18796);
xnor U20211 (N_20211,N_19979,N_19832);
xor U20212 (N_20212,N_19221,N_19892);
xor U20213 (N_20213,N_19506,N_18969);
nand U20214 (N_20214,N_19557,N_19330);
nand U20215 (N_20215,N_19930,N_19518);
xor U20216 (N_20216,N_19051,N_19386);
xnor U20217 (N_20217,N_19612,N_19913);
xnor U20218 (N_20218,N_19305,N_19765);
xnor U20219 (N_20219,N_19778,N_19396);
nand U20220 (N_20220,N_19857,N_18860);
or U20221 (N_20221,N_19993,N_19285);
and U20222 (N_20222,N_19651,N_19493);
or U20223 (N_20223,N_19085,N_19423);
xor U20224 (N_20224,N_19762,N_18789);
nand U20225 (N_20225,N_19264,N_19814);
or U20226 (N_20226,N_18992,N_19988);
xor U20227 (N_20227,N_18839,N_19418);
or U20228 (N_20228,N_19722,N_19388);
nand U20229 (N_20229,N_19907,N_19379);
xor U20230 (N_20230,N_19228,N_19177);
nand U20231 (N_20231,N_19774,N_18793);
xor U20232 (N_20232,N_19210,N_19949);
nand U20233 (N_20233,N_19000,N_19166);
nor U20234 (N_20234,N_18902,N_19203);
and U20235 (N_20235,N_19674,N_19213);
xor U20236 (N_20236,N_18933,N_19500);
nand U20237 (N_20237,N_19676,N_19740);
xnor U20238 (N_20238,N_19039,N_19991);
or U20239 (N_20239,N_19078,N_19968);
or U20240 (N_20240,N_19757,N_18808);
and U20241 (N_20241,N_19999,N_19623);
nor U20242 (N_20242,N_19232,N_19553);
nand U20243 (N_20243,N_19790,N_19443);
or U20244 (N_20244,N_18922,N_19439);
xor U20245 (N_20245,N_19065,N_19149);
or U20246 (N_20246,N_19233,N_19023);
xnor U20247 (N_20247,N_18981,N_19057);
or U20248 (N_20248,N_19961,N_18786);
or U20249 (N_20249,N_19901,N_19401);
nand U20250 (N_20250,N_18756,N_19054);
nand U20251 (N_20251,N_19512,N_18971);
xnor U20252 (N_20252,N_19300,N_19784);
nor U20253 (N_20253,N_19753,N_19748);
and U20254 (N_20254,N_19938,N_19302);
nand U20255 (N_20255,N_19486,N_19698);
nor U20256 (N_20256,N_18942,N_19214);
xor U20257 (N_20257,N_19794,N_18783);
and U20258 (N_20258,N_19594,N_19105);
nor U20259 (N_20259,N_19783,N_19654);
or U20260 (N_20260,N_19387,N_19521);
xor U20261 (N_20261,N_18872,N_18853);
nand U20262 (N_20262,N_19898,N_19934);
or U20263 (N_20263,N_19675,N_19733);
xor U20264 (N_20264,N_18931,N_19116);
or U20265 (N_20265,N_19816,N_19926);
nor U20266 (N_20266,N_19399,N_18794);
and U20267 (N_20267,N_19218,N_19768);
and U20268 (N_20268,N_19268,N_19339);
and U20269 (N_20269,N_18809,N_19983);
nand U20270 (N_20270,N_18780,N_19957);
nor U20271 (N_20271,N_18753,N_19849);
nand U20272 (N_20272,N_19009,N_18916);
nor U20273 (N_20273,N_19810,N_19029);
and U20274 (N_20274,N_19865,N_18963);
nor U20275 (N_20275,N_19484,N_19971);
nor U20276 (N_20276,N_19068,N_18868);
and U20277 (N_20277,N_19308,N_18947);
or U20278 (N_20278,N_19048,N_19172);
xor U20279 (N_20279,N_19481,N_19540);
xnor U20280 (N_20280,N_19627,N_19667);
and U20281 (N_20281,N_19180,N_19046);
nand U20282 (N_20282,N_18883,N_19620);
nand U20283 (N_20283,N_19707,N_19076);
nor U20284 (N_20284,N_19548,N_18855);
nor U20285 (N_20285,N_19858,N_19282);
or U20286 (N_20286,N_19669,N_18859);
or U20287 (N_20287,N_19165,N_18959);
and U20288 (N_20288,N_19573,N_19195);
or U20289 (N_20289,N_19871,N_19267);
xnor U20290 (N_20290,N_18867,N_19280);
or U20291 (N_20291,N_19409,N_19699);
or U20292 (N_20292,N_19176,N_19071);
and U20293 (N_20293,N_19094,N_19520);
or U20294 (N_20294,N_19660,N_18972);
or U20295 (N_20295,N_19702,N_19716);
nor U20296 (N_20296,N_18914,N_19742);
nand U20297 (N_20297,N_19537,N_18834);
nor U20298 (N_20298,N_19831,N_19173);
nor U20299 (N_20299,N_18870,N_19038);
xor U20300 (N_20300,N_19647,N_19850);
nand U20301 (N_20301,N_19148,N_19115);
or U20302 (N_20302,N_19355,N_18863);
xnor U20303 (N_20303,N_19060,N_19672);
nor U20304 (N_20304,N_19402,N_18759);
xnor U20305 (N_20305,N_18856,N_19393);
nor U20306 (N_20306,N_19639,N_19301);
or U20307 (N_20307,N_18903,N_19842);
nand U20308 (N_20308,N_19628,N_19967);
nor U20309 (N_20309,N_19517,N_19395);
or U20310 (N_20310,N_18934,N_19024);
and U20311 (N_20311,N_19215,N_19884);
and U20312 (N_20312,N_19726,N_19238);
or U20313 (N_20313,N_18754,N_18975);
or U20314 (N_20314,N_19049,N_19887);
nand U20315 (N_20315,N_19252,N_19696);
nand U20316 (N_20316,N_19192,N_19937);
xor U20317 (N_20317,N_18773,N_19523);
xor U20318 (N_20318,N_19356,N_19134);
xnor U20319 (N_20319,N_19912,N_19358);
or U20320 (N_20320,N_19547,N_19434);
nand U20321 (N_20321,N_18760,N_19410);
xnor U20322 (N_20322,N_19552,N_19242);
nor U20323 (N_20323,N_19666,N_18924);
nand U20324 (N_20324,N_19715,N_18826);
nor U20325 (N_20325,N_19190,N_19287);
or U20326 (N_20326,N_19222,N_19212);
nand U20327 (N_20327,N_19723,N_19278);
xor U20328 (N_20328,N_19833,N_19931);
nand U20329 (N_20329,N_18960,N_19117);
and U20330 (N_20330,N_19878,N_19591);
and U20331 (N_20331,N_19182,N_19681);
xor U20332 (N_20332,N_19634,N_19114);
xor U20333 (N_20333,N_19122,N_19870);
or U20334 (N_20334,N_19787,N_19345);
nand U20335 (N_20335,N_19956,N_19596);
or U20336 (N_20336,N_19088,N_19193);
nand U20337 (N_20337,N_19061,N_19151);
nor U20338 (N_20338,N_19872,N_18974);
and U20339 (N_20339,N_19313,N_19847);
or U20340 (N_20340,N_19324,N_19338);
or U20341 (N_20341,N_19421,N_18998);
nor U20342 (N_20342,N_19416,N_19298);
xor U20343 (N_20343,N_19411,N_19511);
and U20344 (N_20344,N_19181,N_19041);
or U20345 (N_20345,N_19852,N_19316);
or U20346 (N_20346,N_19688,N_19779);
xor U20347 (N_20347,N_19808,N_19797);
nand U20348 (N_20348,N_19880,N_19476);
xnor U20349 (N_20349,N_19613,N_19855);
xnor U20350 (N_20350,N_19494,N_19083);
xnor U20351 (N_20351,N_19953,N_19641);
nand U20352 (N_20352,N_19081,N_19867);
and U20353 (N_20353,N_19259,N_19296);
and U20354 (N_20354,N_19234,N_19605);
and U20355 (N_20355,N_18941,N_19929);
xor U20356 (N_20356,N_19996,N_19063);
nand U20357 (N_20357,N_19924,N_19741);
xnor U20358 (N_20358,N_19888,N_19853);
xnor U20359 (N_20359,N_19045,N_19525);
nand U20360 (N_20360,N_19914,N_19969);
and U20361 (N_20361,N_19293,N_19284);
nor U20362 (N_20362,N_19376,N_19098);
xor U20363 (N_20363,N_18989,N_18939);
or U20364 (N_20364,N_18778,N_19380);
and U20365 (N_20365,N_19700,N_18927);
or U20366 (N_20366,N_19413,N_19318);
and U20367 (N_20367,N_19310,N_19135);
nand U20368 (N_20368,N_19251,N_19336);
xnor U20369 (N_20369,N_19558,N_19178);
nand U20370 (N_20370,N_19474,N_19398);
or U20371 (N_20371,N_19058,N_19138);
nor U20372 (N_20372,N_19839,N_18938);
nand U20373 (N_20373,N_19570,N_19994);
xnor U20374 (N_20374,N_19087,N_19274);
nor U20375 (N_20375,N_19822,N_19240);
and U20376 (N_20376,N_19798,N_19637);
or U20377 (N_20377,N_19217,N_18806);
and U20378 (N_20378,N_19104,N_19737);
nor U20379 (N_20379,N_19571,N_19905);
or U20380 (N_20380,N_19429,N_19668);
nand U20381 (N_20381,N_19236,N_18948);
nand U20382 (N_20382,N_19258,N_19331);
xor U20383 (N_20383,N_19016,N_19863);
and U20384 (N_20384,N_19686,N_19982);
and U20385 (N_20385,N_19751,N_19921);
nand U20386 (N_20386,N_18805,N_18884);
nor U20387 (N_20387,N_19932,N_19027);
nand U20388 (N_20388,N_19420,N_19576);
and U20389 (N_20389,N_19209,N_19609);
nor U20390 (N_20390,N_19505,N_19012);
or U20391 (N_20391,N_19319,N_18949);
nand U20392 (N_20392,N_19989,N_18982);
nor U20393 (N_20393,N_19828,N_19294);
nor U20394 (N_20394,N_19767,N_18847);
nand U20395 (N_20395,N_19367,N_19942);
nand U20396 (N_20396,N_18923,N_19692);
or U20397 (N_20397,N_19473,N_19303);
and U20398 (N_20398,N_19361,N_19869);
nand U20399 (N_20399,N_19265,N_19146);
or U20400 (N_20400,N_18777,N_19288);
nor U20401 (N_20401,N_18951,N_18774);
nand U20402 (N_20402,N_19764,N_19626);
nand U20403 (N_20403,N_18841,N_19758);
nor U20404 (N_20404,N_19208,N_19363);
nor U20405 (N_20405,N_19270,N_18973);
or U20406 (N_20406,N_18991,N_19066);
and U20407 (N_20407,N_19445,N_19684);
nor U20408 (N_20408,N_18935,N_19981);
and U20409 (N_20409,N_19133,N_19631);
nand U20410 (N_20410,N_18835,N_19197);
nor U20411 (N_20411,N_19734,N_19677);
or U20412 (N_20412,N_19590,N_19438);
nor U20413 (N_20413,N_18958,N_18926);
nand U20414 (N_20414,N_19200,N_19067);
nor U20415 (N_20415,N_18838,N_19145);
or U20416 (N_20416,N_18976,N_19384);
xnor U20417 (N_20417,N_19689,N_19625);
xor U20418 (N_20418,N_19830,N_19050);
and U20419 (N_20419,N_19430,N_19191);
and U20420 (N_20420,N_19454,N_19378);
and U20421 (N_20421,N_18765,N_18882);
xor U20422 (N_20422,N_19074,N_19359);
nor U20423 (N_20423,N_18875,N_19162);
xor U20424 (N_20424,N_19841,N_19846);
nand U20425 (N_20425,N_19136,N_19827);
and U20426 (N_20426,N_19614,N_19007);
or U20427 (N_20427,N_19959,N_19189);
or U20428 (N_20428,N_18768,N_19910);
nand U20429 (N_20429,N_18876,N_19198);
nor U20430 (N_20430,N_19154,N_18913);
nand U20431 (N_20431,N_19708,N_18844);
xnor U20432 (N_20432,N_19984,N_19109);
xor U20433 (N_20433,N_19977,N_19745);
xnor U20434 (N_20434,N_19171,N_19522);
and U20435 (N_20435,N_19653,N_19496);
nor U20436 (N_20436,N_19391,N_19403);
and U20437 (N_20437,N_19896,N_19501);
nor U20438 (N_20438,N_19448,N_19881);
and U20439 (N_20439,N_19194,N_19253);
nor U20440 (N_20440,N_19633,N_19001);
nand U20441 (N_20441,N_19343,N_19551);
nor U20442 (N_20442,N_19756,N_19752);
or U20443 (N_20443,N_19342,N_19542);
xnor U20444 (N_20444,N_19347,N_19851);
xnor U20445 (N_20445,N_19436,N_19408);
and U20446 (N_20446,N_18944,N_19488);
or U20447 (N_20447,N_18770,N_18886);
and U20448 (N_20448,N_19371,N_19925);
and U20449 (N_20449,N_19291,N_19703);
nor U20450 (N_20450,N_19174,N_19656);
nor U20451 (N_20451,N_19718,N_18775);
xor U20452 (N_20452,N_19281,N_19601);
nand U20453 (N_20453,N_19629,N_19885);
nor U20454 (N_20454,N_19515,N_18791);
or U20455 (N_20455,N_19026,N_19785);
nand U20456 (N_20456,N_18919,N_19687);
nor U20457 (N_20457,N_19550,N_19978);
and U20458 (N_20458,N_19918,N_19709);
nand U20459 (N_20459,N_19510,N_19568);
and U20460 (N_20460,N_19216,N_19125);
xor U20461 (N_20461,N_19306,N_19532);
or U20462 (N_20462,N_19735,N_19266);
or U20463 (N_20463,N_19611,N_19142);
nand U20464 (N_20464,N_19835,N_19671);
and U20465 (N_20465,N_18891,N_19710);
and U20466 (N_20466,N_19179,N_19780);
or U20467 (N_20467,N_19670,N_19975);
or U20468 (N_20468,N_18911,N_19948);
and U20469 (N_20469,N_19279,N_19199);
nand U20470 (N_20470,N_19739,N_19820);
nor U20471 (N_20471,N_19585,N_19803);
nand U20472 (N_20472,N_18893,N_19158);
nand U20473 (N_20473,N_19664,N_19529);
or U20474 (N_20474,N_19032,N_18898);
nor U20475 (N_20475,N_19022,N_19464);
or U20476 (N_20476,N_19543,N_19825);
nand U20477 (N_20477,N_19834,N_19770);
xnor U20478 (N_20478,N_19624,N_19895);
nor U20479 (N_20479,N_19527,N_19811);
xor U20480 (N_20480,N_19185,N_19456);
and U20481 (N_20481,N_18952,N_19315);
and U20482 (N_20482,N_19581,N_19845);
or U20483 (N_20483,N_19504,N_19422);
nand U20484 (N_20484,N_19891,N_19958);
nor U20485 (N_20485,N_19998,N_19836);
nor U20486 (N_20486,N_19920,N_19777);
nand U20487 (N_20487,N_19859,N_19648);
or U20488 (N_20488,N_19894,N_19377);
nand U20489 (N_20489,N_18851,N_19277);
or U20490 (N_20490,N_19091,N_19442);
nand U20491 (N_20491,N_19617,N_19295);
and U20492 (N_20492,N_19546,N_19823);
or U20493 (N_20493,N_19796,N_19578);
and U20494 (N_20494,N_19487,N_19761);
and U20495 (N_20495,N_18818,N_18800);
and U20496 (N_20496,N_19433,N_19440);
or U20497 (N_20497,N_19097,N_19175);
and U20498 (N_20498,N_19349,N_19943);
nor U20499 (N_20499,N_19382,N_19219);
or U20500 (N_20500,N_19113,N_18840);
and U20501 (N_20501,N_19011,N_18968);
and U20502 (N_20502,N_19003,N_19800);
or U20503 (N_20503,N_19034,N_18846);
xnor U20504 (N_20504,N_19952,N_19545);
and U20505 (N_20505,N_18945,N_18785);
nor U20506 (N_20506,N_19706,N_18878);
and U20507 (N_20507,N_18950,N_19469);
xor U20508 (N_20508,N_19701,N_19936);
nand U20509 (N_20509,N_18849,N_18830);
nor U20510 (N_20510,N_18810,N_18828);
and U20511 (N_20511,N_19673,N_19390);
nand U20512 (N_20512,N_19799,N_19963);
and U20513 (N_20513,N_19713,N_19089);
nand U20514 (N_20514,N_19604,N_19062);
xnor U20515 (N_20515,N_18895,N_19580);
nand U20516 (N_20516,N_19607,N_19340);
nor U20517 (N_20517,N_19732,N_18918);
and U20518 (N_20518,N_19044,N_19563);
and U20519 (N_20519,N_18857,N_19118);
xnor U20520 (N_20520,N_18763,N_19976);
nor U20521 (N_20521,N_18940,N_19712);
nand U20522 (N_20522,N_19093,N_19064);
xnor U20523 (N_20523,N_19866,N_18907);
and U20524 (N_20524,N_19694,N_19815);
or U20525 (N_20525,N_19569,N_18967);
nand U20526 (N_20526,N_19775,N_19069);
and U20527 (N_20527,N_19108,N_19110);
or U20528 (N_20528,N_18901,N_19344);
nand U20529 (N_20529,N_19286,N_19006);
and U20530 (N_20530,N_19466,N_19297);
and U20531 (N_20531,N_19206,N_19908);
nand U20532 (N_20532,N_18970,N_19919);
nand U20533 (N_20533,N_19441,N_19771);
nor U20534 (N_20534,N_19549,N_19383);
nor U20535 (N_20535,N_18820,N_19955);
nor U20536 (N_20536,N_19714,N_18997);
nor U20537 (N_20537,N_18961,N_18825);
nand U20538 (N_20538,N_19099,N_19927);
xor U20539 (N_20539,N_19602,N_19257);
xor U20540 (N_20540,N_19100,N_19370);
or U20541 (N_20541,N_19499,N_19077);
or U20542 (N_20542,N_19159,N_19730);
xnor U20543 (N_20543,N_18983,N_19008);
nor U20544 (N_20544,N_18978,N_18824);
nand U20545 (N_20545,N_19156,N_19269);
xnor U20546 (N_20546,N_18769,N_19904);
nor U20547 (N_20547,N_18842,N_18861);
xnor U20548 (N_20548,N_19126,N_19864);
nand U20549 (N_20549,N_18908,N_19458);
xor U20550 (N_20550,N_19724,N_19055);
or U20551 (N_20551,N_19603,N_19207);
xnor U20552 (N_20552,N_18985,N_19256);
xnor U20553 (N_20553,N_19480,N_18787);
nor U20554 (N_20554,N_19945,N_18757);
nand U20555 (N_20555,N_18812,N_19682);
nand U20556 (N_20556,N_19452,N_19879);
xor U20557 (N_20557,N_18865,N_19838);
xor U20558 (N_20558,N_18874,N_19224);
nand U20559 (N_20559,N_19567,N_18799);
and U20560 (N_20560,N_18804,N_19453);
or U20561 (N_20561,N_19211,N_19472);
or U20562 (N_20562,N_19326,N_19164);
and U20563 (N_20563,N_19201,N_19328);
nand U20564 (N_20564,N_19555,N_19351);
nor U20565 (N_20565,N_19621,N_19530);
or U20566 (N_20566,N_18988,N_19059);
xnor U20567 (N_20567,N_19899,N_18797);
or U20568 (N_20568,N_19364,N_19947);
nor U20569 (N_20569,N_19526,N_19153);
nand U20570 (N_20570,N_19397,N_18880);
nor U20571 (N_20571,N_19610,N_19072);
or U20572 (N_20572,N_19372,N_19586);
nand U20573 (N_20573,N_19806,N_18772);
xnor U20574 (N_20574,N_19357,N_19004);
xor U20575 (N_20575,N_18910,N_18873);
nor U20576 (N_20576,N_19428,N_19348);
or U20577 (N_20577,N_19014,N_18848);
or U20578 (N_20578,N_18801,N_19655);
and U20579 (N_20579,N_19128,N_19974);
and U20580 (N_20580,N_19782,N_19020);
or U20581 (N_20581,N_19802,N_19374);
nor U20582 (N_20582,N_18764,N_19187);
nand U20583 (N_20583,N_18784,N_18937);
and U20584 (N_20584,N_19033,N_19460);
or U20585 (N_20585,N_19848,N_19407);
or U20586 (N_20586,N_19911,N_19170);
nand U20587 (N_20587,N_19817,N_19160);
nand U20588 (N_20588,N_19152,N_18925);
nand U20589 (N_20589,N_19271,N_19922);
xnor U20590 (N_20590,N_19205,N_19584);
xnor U20591 (N_20591,N_19311,N_19973);
and U20592 (N_20592,N_19021,N_19941);
or U20593 (N_20593,N_18833,N_19746);
xnor U20594 (N_20594,N_19106,N_19508);
xor U20595 (N_20595,N_19657,N_19749);
nand U20596 (N_20596,N_19272,N_18822);
and U20597 (N_20597,N_19186,N_19084);
xor U20598 (N_20598,N_19144,N_19645);
xor U20599 (N_20599,N_18802,N_19161);
nor U20600 (N_20600,N_19130,N_19744);
xor U20601 (N_20601,N_19414,N_19640);
and U20602 (N_20602,N_19650,N_19485);
and U20603 (N_20603,N_19582,N_18920);
xnor U20604 (N_20604,N_19813,N_19119);
and U20605 (N_20605,N_18862,N_19964);
and U20606 (N_20606,N_18816,N_18843);
and U20607 (N_20607,N_19906,N_19966);
nor U20608 (N_20608,N_19457,N_19017);
or U20609 (N_20609,N_19987,N_18986);
or U20610 (N_20610,N_18928,N_18894);
nand U20611 (N_20611,N_19695,N_18767);
xor U20612 (N_20612,N_19432,N_19444);
or U20613 (N_20613,N_19028,N_19471);
xnor U20614 (N_20614,N_19536,N_19465);
nand U20615 (N_20615,N_19763,N_19662);
xor U20616 (N_20616,N_19321,N_19360);
or U20617 (N_20617,N_19036,N_18897);
nand U20618 (N_20618,N_19965,N_19516);
or U20619 (N_20619,N_18817,N_19598);
nand U20620 (N_20620,N_19231,N_19437);
and U20621 (N_20621,N_18813,N_19314);
and U20622 (N_20622,N_19554,N_18829);
xnor U20623 (N_20623,N_19086,N_19140);
and U20624 (N_20624,N_19646,N_19566);
nor U20625 (N_20625,N_19542,N_19392);
and U20626 (N_20626,N_19964,N_19335);
and U20627 (N_20627,N_19281,N_19117);
nor U20628 (N_20628,N_19926,N_19780);
and U20629 (N_20629,N_19844,N_19911);
nand U20630 (N_20630,N_18808,N_19156);
xor U20631 (N_20631,N_18821,N_19312);
nand U20632 (N_20632,N_19015,N_19533);
or U20633 (N_20633,N_19106,N_19382);
nor U20634 (N_20634,N_19230,N_19367);
and U20635 (N_20635,N_19323,N_19954);
xnor U20636 (N_20636,N_19336,N_19110);
nand U20637 (N_20637,N_19909,N_19866);
nand U20638 (N_20638,N_19125,N_19850);
or U20639 (N_20639,N_19408,N_19918);
xnor U20640 (N_20640,N_19922,N_19782);
xnor U20641 (N_20641,N_19906,N_19393);
and U20642 (N_20642,N_18837,N_19396);
nor U20643 (N_20643,N_19193,N_19866);
nand U20644 (N_20644,N_19652,N_19042);
or U20645 (N_20645,N_19195,N_19911);
nand U20646 (N_20646,N_19030,N_19767);
or U20647 (N_20647,N_19058,N_18827);
and U20648 (N_20648,N_19036,N_19668);
xor U20649 (N_20649,N_18785,N_19815);
xor U20650 (N_20650,N_19905,N_19263);
or U20651 (N_20651,N_19549,N_19206);
xor U20652 (N_20652,N_19241,N_19501);
and U20653 (N_20653,N_19735,N_19183);
xnor U20654 (N_20654,N_19558,N_19265);
nor U20655 (N_20655,N_19296,N_19515);
or U20656 (N_20656,N_19124,N_19294);
or U20657 (N_20657,N_19551,N_19075);
xor U20658 (N_20658,N_19896,N_19366);
nor U20659 (N_20659,N_19335,N_18838);
nor U20660 (N_20660,N_19847,N_18858);
xor U20661 (N_20661,N_19999,N_18877);
and U20662 (N_20662,N_18904,N_19490);
and U20663 (N_20663,N_19504,N_19016);
or U20664 (N_20664,N_19563,N_18987);
nand U20665 (N_20665,N_19616,N_19919);
xnor U20666 (N_20666,N_19034,N_19183);
and U20667 (N_20667,N_19217,N_19309);
or U20668 (N_20668,N_19780,N_19067);
and U20669 (N_20669,N_19522,N_18988);
xnor U20670 (N_20670,N_18923,N_19224);
and U20671 (N_20671,N_19417,N_18835);
or U20672 (N_20672,N_19322,N_18975);
or U20673 (N_20673,N_19864,N_19200);
or U20674 (N_20674,N_19890,N_19115);
or U20675 (N_20675,N_19203,N_19730);
nand U20676 (N_20676,N_19109,N_19681);
xor U20677 (N_20677,N_18957,N_19261);
or U20678 (N_20678,N_18943,N_19700);
or U20679 (N_20679,N_19766,N_19102);
xor U20680 (N_20680,N_19458,N_18846);
nand U20681 (N_20681,N_18865,N_19469);
nand U20682 (N_20682,N_18850,N_18889);
and U20683 (N_20683,N_18756,N_18779);
and U20684 (N_20684,N_19901,N_19037);
nand U20685 (N_20685,N_19589,N_19624);
xor U20686 (N_20686,N_19591,N_18807);
nand U20687 (N_20687,N_19947,N_19821);
nand U20688 (N_20688,N_19063,N_18871);
or U20689 (N_20689,N_19171,N_19084);
xor U20690 (N_20690,N_19036,N_19969);
xor U20691 (N_20691,N_19759,N_19475);
nand U20692 (N_20692,N_19696,N_19593);
and U20693 (N_20693,N_19870,N_19366);
and U20694 (N_20694,N_19697,N_18777);
xnor U20695 (N_20695,N_18998,N_19557);
xor U20696 (N_20696,N_19638,N_19997);
nor U20697 (N_20697,N_18882,N_19341);
and U20698 (N_20698,N_19408,N_19801);
nor U20699 (N_20699,N_18788,N_18985);
and U20700 (N_20700,N_19144,N_19421);
nor U20701 (N_20701,N_19779,N_18985);
xor U20702 (N_20702,N_19190,N_18934);
xor U20703 (N_20703,N_19109,N_18888);
xnor U20704 (N_20704,N_19622,N_18753);
nor U20705 (N_20705,N_18819,N_19719);
nor U20706 (N_20706,N_19124,N_19008);
nor U20707 (N_20707,N_18851,N_19718);
or U20708 (N_20708,N_19972,N_19271);
and U20709 (N_20709,N_19796,N_19763);
xor U20710 (N_20710,N_18860,N_19904);
xnor U20711 (N_20711,N_19994,N_19533);
or U20712 (N_20712,N_19138,N_19909);
and U20713 (N_20713,N_18915,N_19875);
or U20714 (N_20714,N_19548,N_19785);
nor U20715 (N_20715,N_19871,N_19742);
nand U20716 (N_20716,N_19779,N_19427);
and U20717 (N_20717,N_19163,N_19035);
nor U20718 (N_20718,N_19165,N_18917);
nand U20719 (N_20719,N_19722,N_19463);
xor U20720 (N_20720,N_19323,N_19592);
and U20721 (N_20721,N_19469,N_19117);
nand U20722 (N_20722,N_19359,N_18843);
xnor U20723 (N_20723,N_19017,N_19264);
or U20724 (N_20724,N_18955,N_19133);
nor U20725 (N_20725,N_19856,N_19763);
xnor U20726 (N_20726,N_19662,N_18962);
xnor U20727 (N_20727,N_19097,N_19552);
nand U20728 (N_20728,N_19610,N_19792);
or U20729 (N_20729,N_19942,N_19317);
xor U20730 (N_20730,N_18852,N_18860);
or U20731 (N_20731,N_19414,N_19613);
and U20732 (N_20732,N_19715,N_18876);
or U20733 (N_20733,N_18934,N_19676);
and U20734 (N_20734,N_19274,N_19585);
or U20735 (N_20735,N_19768,N_19745);
xor U20736 (N_20736,N_18993,N_19602);
xor U20737 (N_20737,N_19048,N_19176);
xor U20738 (N_20738,N_19229,N_18974);
and U20739 (N_20739,N_19657,N_19439);
nand U20740 (N_20740,N_18906,N_19741);
or U20741 (N_20741,N_19541,N_19039);
nor U20742 (N_20742,N_19481,N_18796);
nand U20743 (N_20743,N_19653,N_18817);
nand U20744 (N_20744,N_19876,N_19067);
xnor U20745 (N_20745,N_19318,N_19525);
nor U20746 (N_20746,N_19083,N_19365);
nor U20747 (N_20747,N_19832,N_19219);
or U20748 (N_20748,N_19318,N_19886);
and U20749 (N_20749,N_19763,N_19788);
nor U20750 (N_20750,N_18966,N_19796);
xnor U20751 (N_20751,N_18750,N_19066);
xor U20752 (N_20752,N_19718,N_19140);
nand U20753 (N_20753,N_19718,N_19018);
xor U20754 (N_20754,N_19684,N_18784);
nand U20755 (N_20755,N_19789,N_19730);
nor U20756 (N_20756,N_19506,N_19548);
xor U20757 (N_20757,N_19397,N_19426);
or U20758 (N_20758,N_19503,N_19249);
or U20759 (N_20759,N_19759,N_19639);
or U20760 (N_20760,N_19821,N_19089);
xnor U20761 (N_20761,N_18877,N_19607);
or U20762 (N_20762,N_18760,N_19867);
xor U20763 (N_20763,N_19882,N_19580);
or U20764 (N_20764,N_19800,N_19539);
and U20765 (N_20765,N_19503,N_18892);
and U20766 (N_20766,N_18861,N_19586);
or U20767 (N_20767,N_19020,N_19716);
nand U20768 (N_20768,N_18776,N_19609);
or U20769 (N_20769,N_19588,N_19309);
nand U20770 (N_20770,N_18955,N_19011);
and U20771 (N_20771,N_19382,N_19347);
or U20772 (N_20772,N_19668,N_19754);
xor U20773 (N_20773,N_19419,N_19819);
nor U20774 (N_20774,N_19338,N_19561);
nand U20775 (N_20775,N_18852,N_18904);
and U20776 (N_20776,N_19062,N_18830);
xnor U20777 (N_20777,N_19030,N_19949);
nand U20778 (N_20778,N_19157,N_19707);
xor U20779 (N_20779,N_19250,N_19834);
nor U20780 (N_20780,N_19023,N_18933);
or U20781 (N_20781,N_19291,N_19978);
or U20782 (N_20782,N_19487,N_19451);
xor U20783 (N_20783,N_19430,N_19842);
nor U20784 (N_20784,N_18990,N_19166);
and U20785 (N_20785,N_18932,N_18802);
nand U20786 (N_20786,N_19973,N_19363);
nor U20787 (N_20787,N_19034,N_18950);
or U20788 (N_20788,N_18843,N_19105);
or U20789 (N_20789,N_19412,N_19710);
nand U20790 (N_20790,N_19323,N_18927);
nor U20791 (N_20791,N_19534,N_19455);
or U20792 (N_20792,N_19618,N_19791);
nand U20793 (N_20793,N_18970,N_19419);
xnor U20794 (N_20794,N_19581,N_19230);
nor U20795 (N_20795,N_19485,N_19677);
nor U20796 (N_20796,N_19722,N_19434);
nor U20797 (N_20797,N_18889,N_19098);
xnor U20798 (N_20798,N_19577,N_19298);
nor U20799 (N_20799,N_19400,N_19363);
nor U20800 (N_20800,N_18832,N_19451);
nand U20801 (N_20801,N_19849,N_19438);
xnor U20802 (N_20802,N_19142,N_19402);
nand U20803 (N_20803,N_19932,N_18972);
xor U20804 (N_20804,N_19284,N_18925);
nor U20805 (N_20805,N_18981,N_19192);
nor U20806 (N_20806,N_18910,N_19746);
and U20807 (N_20807,N_18931,N_19587);
nand U20808 (N_20808,N_19641,N_19709);
or U20809 (N_20809,N_18755,N_18956);
or U20810 (N_20810,N_19871,N_19733);
nand U20811 (N_20811,N_19901,N_19373);
nor U20812 (N_20812,N_19733,N_19815);
nor U20813 (N_20813,N_18845,N_19809);
xor U20814 (N_20814,N_19172,N_19744);
nand U20815 (N_20815,N_19257,N_18921);
nor U20816 (N_20816,N_19162,N_19762);
and U20817 (N_20817,N_19647,N_19516);
nand U20818 (N_20818,N_19687,N_19116);
or U20819 (N_20819,N_19711,N_19215);
xnor U20820 (N_20820,N_19856,N_18944);
xor U20821 (N_20821,N_19727,N_19486);
and U20822 (N_20822,N_19212,N_19132);
or U20823 (N_20823,N_19728,N_19022);
and U20824 (N_20824,N_18959,N_19776);
nand U20825 (N_20825,N_18770,N_19937);
nor U20826 (N_20826,N_19675,N_19765);
xor U20827 (N_20827,N_19644,N_19373);
and U20828 (N_20828,N_19849,N_18979);
nor U20829 (N_20829,N_19500,N_19966);
xor U20830 (N_20830,N_19815,N_19679);
and U20831 (N_20831,N_19751,N_18936);
nor U20832 (N_20832,N_19409,N_18995);
or U20833 (N_20833,N_19382,N_19926);
nand U20834 (N_20834,N_19182,N_19880);
nand U20835 (N_20835,N_18917,N_18974);
or U20836 (N_20836,N_19136,N_19345);
nand U20837 (N_20837,N_18750,N_19465);
and U20838 (N_20838,N_19468,N_19993);
nor U20839 (N_20839,N_19252,N_19797);
or U20840 (N_20840,N_19943,N_19359);
nor U20841 (N_20841,N_19058,N_19889);
and U20842 (N_20842,N_19482,N_19735);
or U20843 (N_20843,N_19450,N_19706);
and U20844 (N_20844,N_19020,N_19358);
nor U20845 (N_20845,N_19691,N_19967);
or U20846 (N_20846,N_19266,N_19566);
nand U20847 (N_20847,N_18958,N_19813);
nor U20848 (N_20848,N_19623,N_19697);
and U20849 (N_20849,N_19954,N_19430);
nand U20850 (N_20850,N_19380,N_19288);
nor U20851 (N_20851,N_19042,N_19658);
xnor U20852 (N_20852,N_19241,N_19219);
and U20853 (N_20853,N_19316,N_19822);
and U20854 (N_20854,N_19683,N_19979);
nor U20855 (N_20855,N_19492,N_18997);
and U20856 (N_20856,N_18867,N_19198);
xnor U20857 (N_20857,N_19293,N_19058);
nor U20858 (N_20858,N_18974,N_19179);
nor U20859 (N_20859,N_19448,N_19977);
nor U20860 (N_20860,N_19038,N_19700);
nor U20861 (N_20861,N_19433,N_19137);
nor U20862 (N_20862,N_18949,N_19643);
and U20863 (N_20863,N_19105,N_19747);
nor U20864 (N_20864,N_19913,N_19897);
or U20865 (N_20865,N_19242,N_18885);
or U20866 (N_20866,N_19805,N_19825);
or U20867 (N_20867,N_19719,N_19804);
nor U20868 (N_20868,N_18855,N_19434);
or U20869 (N_20869,N_19211,N_19413);
xnor U20870 (N_20870,N_19760,N_19763);
and U20871 (N_20871,N_18800,N_19307);
nand U20872 (N_20872,N_19379,N_19537);
xnor U20873 (N_20873,N_19095,N_19829);
nand U20874 (N_20874,N_19088,N_19801);
and U20875 (N_20875,N_19492,N_19533);
or U20876 (N_20876,N_19733,N_19143);
and U20877 (N_20877,N_19763,N_18936);
or U20878 (N_20878,N_19461,N_19563);
or U20879 (N_20879,N_19532,N_19131);
or U20880 (N_20880,N_19970,N_19554);
nor U20881 (N_20881,N_19640,N_19973);
nor U20882 (N_20882,N_18893,N_18780);
nor U20883 (N_20883,N_19038,N_19803);
or U20884 (N_20884,N_19323,N_19062);
nor U20885 (N_20885,N_19032,N_19020);
nand U20886 (N_20886,N_19101,N_18873);
or U20887 (N_20887,N_19393,N_19136);
nand U20888 (N_20888,N_18938,N_19799);
or U20889 (N_20889,N_19102,N_19123);
nand U20890 (N_20890,N_19624,N_19942);
and U20891 (N_20891,N_19680,N_19321);
xnor U20892 (N_20892,N_19940,N_19468);
nand U20893 (N_20893,N_18807,N_19292);
xnor U20894 (N_20894,N_19356,N_19832);
nand U20895 (N_20895,N_19879,N_19239);
nor U20896 (N_20896,N_19699,N_19250);
nor U20897 (N_20897,N_19595,N_19998);
and U20898 (N_20898,N_18961,N_19903);
nand U20899 (N_20899,N_19692,N_19949);
and U20900 (N_20900,N_19906,N_19178);
or U20901 (N_20901,N_19718,N_19784);
xnor U20902 (N_20902,N_19231,N_19101);
or U20903 (N_20903,N_19951,N_19594);
or U20904 (N_20904,N_18836,N_19983);
or U20905 (N_20905,N_18853,N_19006);
and U20906 (N_20906,N_19567,N_18833);
or U20907 (N_20907,N_19722,N_19305);
and U20908 (N_20908,N_19826,N_19298);
xnor U20909 (N_20909,N_19124,N_19040);
or U20910 (N_20910,N_19243,N_18917);
and U20911 (N_20911,N_18845,N_18814);
nand U20912 (N_20912,N_19018,N_19032);
xnor U20913 (N_20913,N_19161,N_19332);
and U20914 (N_20914,N_18899,N_19869);
nor U20915 (N_20915,N_18864,N_19090);
nor U20916 (N_20916,N_19523,N_19662);
and U20917 (N_20917,N_19806,N_19357);
nor U20918 (N_20918,N_19911,N_19601);
or U20919 (N_20919,N_19943,N_19774);
nand U20920 (N_20920,N_18976,N_19013);
or U20921 (N_20921,N_19369,N_18844);
and U20922 (N_20922,N_18970,N_19764);
nor U20923 (N_20923,N_18769,N_19637);
or U20924 (N_20924,N_19736,N_19571);
nor U20925 (N_20925,N_19940,N_19906);
nand U20926 (N_20926,N_19785,N_19258);
nand U20927 (N_20927,N_19723,N_19404);
and U20928 (N_20928,N_19272,N_19349);
and U20929 (N_20929,N_19416,N_19950);
nor U20930 (N_20930,N_19788,N_19748);
nor U20931 (N_20931,N_19018,N_19911);
and U20932 (N_20932,N_19640,N_18867);
nand U20933 (N_20933,N_18848,N_19717);
xor U20934 (N_20934,N_18765,N_18922);
nand U20935 (N_20935,N_19808,N_18983);
nand U20936 (N_20936,N_19268,N_19335);
nor U20937 (N_20937,N_18966,N_19618);
nor U20938 (N_20938,N_19085,N_18843);
nand U20939 (N_20939,N_19394,N_19814);
or U20940 (N_20940,N_19258,N_19017);
or U20941 (N_20941,N_19423,N_18997);
and U20942 (N_20942,N_19395,N_19391);
or U20943 (N_20943,N_19855,N_18794);
and U20944 (N_20944,N_19555,N_19792);
and U20945 (N_20945,N_19658,N_18971);
or U20946 (N_20946,N_19644,N_19329);
and U20947 (N_20947,N_18864,N_19701);
and U20948 (N_20948,N_19557,N_19292);
or U20949 (N_20949,N_19247,N_19329);
or U20950 (N_20950,N_19133,N_19622);
nand U20951 (N_20951,N_19323,N_19629);
and U20952 (N_20952,N_19545,N_19439);
or U20953 (N_20953,N_19802,N_19690);
and U20954 (N_20954,N_19836,N_19498);
and U20955 (N_20955,N_18866,N_19491);
nand U20956 (N_20956,N_18956,N_19058);
or U20957 (N_20957,N_18985,N_18988);
or U20958 (N_20958,N_19973,N_19151);
xnor U20959 (N_20959,N_19263,N_19206);
xnor U20960 (N_20960,N_18958,N_19463);
and U20961 (N_20961,N_18907,N_19984);
or U20962 (N_20962,N_19226,N_19877);
nand U20963 (N_20963,N_19989,N_19654);
nor U20964 (N_20964,N_19094,N_18870);
or U20965 (N_20965,N_18774,N_19024);
or U20966 (N_20966,N_19152,N_19757);
nand U20967 (N_20967,N_19541,N_19935);
xnor U20968 (N_20968,N_18918,N_19184);
nor U20969 (N_20969,N_19389,N_19518);
or U20970 (N_20970,N_19608,N_19169);
and U20971 (N_20971,N_19349,N_19000);
or U20972 (N_20972,N_19745,N_19254);
nand U20973 (N_20973,N_19516,N_19068);
nor U20974 (N_20974,N_19895,N_19791);
or U20975 (N_20975,N_18755,N_18989);
and U20976 (N_20976,N_19842,N_19247);
xor U20977 (N_20977,N_19123,N_18919);
or U20978 (N_20978,N_19934,N_19685);
and U20979 (N_20979,N_19857,N_18783);
xor U20980 (N_20980,N_19505,N_19893);
and U20981 (N_20981,N_19565,N_19560);
nand U20982 (N_20982,N_19921,N_19138);
or U20983 (N_20983,N_19527,N_19123);
xor U20984 (N_20984,N_18854,N_19867);
and U20985 (N_20985,N_19660,N_19695);
xor U20986 (N_20986,N_19589,N_19324);
nand U20987 (N_20987,N_19720,N_19155);
nor U20988 (N_20988,N_19586,N_18849);
or U20989 (N_20989,N_19663,N_19735);
nand U20990 (N_20990,N_19408,N_19466);
xor U20991 (N_20991,N_19996,N_18852);
nand U20992 (N_20992,N_19216,N_19677);
nand U20993 (N_20993,N_19018,N_19864);
nand U20994 (N_20994,N_19096,N_19965);
xor U20995 (N_20995,N_19668,N_19451);
and U20996 (N_20996,N_18810,N_19953);
xnor U20997 (N_20997,N_19047,N_19578);
nand U20998 (N_20998,N_19986,N_18860);
xor U20999 (N_20999,N_19694,N_19398);
nand U21000 (N_21000,N_19992,N_19852);
and U21001 (N_21001,N_19767,N_19633);
nor U21002 (N_21002,N_18988,N_19743);
xor U21003 (N_21003,N_19411,N_19975);
and U21004 (N_21004,N_18945,N_19751);
nand U21005 (N_21005,N_18931,N_19057);
nand U21006 (N_21006,N_19813,N_19374);
or U21007 (N_21007,N_19381,N_18772);
xnor U21008 (N_21008,N_19943,N_18790);
nor U21009 (N_21009,N_19280,N_19291);
or U21010 (N_21010,N_19472,N_18861);
nor U21011 (N_21011,N_18982,N_19629);
xor U21012 (N_21012,N_19048,N_19046);
nand U21013 (N_21013,N_19509,N_19425);
and U21014 (N_21014,N_19335,N_18941);
and U21015 (N_21015,N_19776,N_19917);
nand U21016 (N_21016,N_18865,N_19607);
nand U21017 (N_21017,N_19619,N_19810);
xnor U21018 (N_21018,N_19037,N_19382);
and U21019 (N_21019,N_19005,N_18968);
nor U21020 (N_21020,N_19355,N_19497);
and U21021 (N_21021,N_19119,N_19097);
xnor U21022 (N_21022,N_19461,N_19289);
and U21023 (N_21023,N_19399,N_19669);
or U21024 (N_21024,N_19337,N_19651);
nor U21025 (N_21025,N_19281,N_19728);
nand U21026 (N_21026,N_19871,N_19912);
and U21027 (N_21027,N_19811,N_19172);
and U21028 (N_21028,N_19267,N_19443);
nor U21029 (N_21029,N_19014,N_19948);
or U21030 (N_21030,N_18855,N_19313);
xnor U21031 (N_21031,N_19056,N_19610);
xnor U21032 (N_21032,N_19913,N_18858);
and U21033 (N_21033,N_19685,N_19767);
nand U21034 (N_21034,N_19289,N_18872);
xor U21035 (N_21035,N_19396,N_19446);
nor U21036 (N_21036,N_18947,N_19391);
nor U21037 (N_21037,N_19511,N_19496);
xor U21038 (N_21038,N_18878,N_19987);
and U21039 (N_21039,N_18968,N_18963);
nand U21040 (N_21040,N_18937,N_19044);
xnor U21041 (N_21041,N_19286,N_19940);
nand U21042 (N_21042,N_19545,N_19488);
xnor U21043 (N_21043,N_19726,N_18874);
nor U21044 (N_21044,N_19039,N_19691);
or U21045 (N_21045,N_19949,N_18878);
and U21046 (N_21046,N_18944,N_19186);
nor U21047 (N_21047,N_18857,N_19734);
nor U21048 (N_21048,N_19404,N_19917);
nor U21049 (N_21049,N_18902,N_19064);
and U21050 (N_21050,N_18769,N_19522);
and U21051 (N_21051,N_18900,N_19374);
or U21052 (N_21052,N_19874,N_19907);
or U21053 (N_21053,N_19554,N_18782);
or U21054 (N_21054,N_19991,N_19494);
or U21055 (N_21055,N_18897,N_19532);
nor U21056 (N_21056,N_19240,N_18978);
xnor U21057 (N_21057,N_19357,N_19525);
and U21058 (N_21058,N_19643,N_19177);
nand U21059 (N_21059,N_18918,N_19749);
xor U21060 (N_21060,N_19665,N_19082);
or U21061 (N_21061,N_19697,N_19632);
nand U21062 (N_21062,N_19504,N_19804);
nor U21063 (N_21063,N_18781,N_19461);
and U21064 (N_21064,N_19252,N_19923);
or U21065 (N_21065,N_19732,N_19346);
and U21066 (N_21066,N_18816,N_19964);
nor U21067 (N_21067,N_19696,N_19110);
or U21068 (N_21068,N_19623,N_19147);
nor U21069 (N_21069,N_19922,N_18754);
xnor U21070 (N_21070,N_19870,N_19302);
nand U21071 (N_21071,N_19404,N_19855);
and U21072 (N_21072,N_19613,N_19722);
xor U21073 (N_21073,N_19832,N_19659);
or U21074 (N_21074,N_18838,N_19788);
nand U21075 (N_21075,N_19596,N_18802);
xnor U21076 (N_21076,N_19623,N_19614);
and U21077 (N_21077,N_18869,N_19507);
and U21078 (N_21078,N_19450,N_18782);
nand U21079 (N_21079,N_19398,N_18918);
nand U21080 (N_21080,N_18842,N_19225);
nor U21081 (N_21081,N_19868,N_19224);
nor U21082 (N_21082,N_19171,N_19933);
nor U21083 (N_21083,N_19128,N_19323);
and U21084 (N_21084,N_19212,N_19334);
or U21085 (N_21085,N_19674,N_19415);
and U21086 (N_21086,N_19694,N_19192);
or U21087 (N_21087,N_19661,N_19563);
xor U21088 (N_21088,N_19769,N_19276);
xnor U21089 (N_21089,N_18792,N_18772);
or U21090 (N_21090,N_19688,N_19634);
or U21091 (N_21091,N_19707,N_19689);
xnor U21092 (N_21092,N_19046,N_19357);
xor U21093 (N_21093,N_19956,N_19179);
and U21094 (N_21094,N_19505,N_19872);
or U21095 (N_21095,N_18910,N_19227);
and U21096 (N_21096,N_18837,N_19959);
or U21097 (N_21097,N_19439,N_19357);
nor U21098 (N_21098,N_19702,N_18841);
nand U21099 (N_21099,N_19981,N_19644);
nand U21100 (N_21100,N_19036,N_18794);
nor U21101 (N_21101,N_19708,N_19432);
nand U21102 (N_21102,N_19372,N_18850);
nor U21103 (N_21103,N_19200,N_19054);
nand U21104 (N_21104,N_18955,N_19374);
xnor U21105 (N_21105,N_19081,N_18809);
nor U21106 (N_21106,N_19886,N_19591);
nor U21107 (N_21107,N_19595,N_19964);
nor U21108 (N_21108,N_19773,N_18911);
nand U21109 (N_21109,N_19671,N_19872);
xnor U21110 (N_21110,N_18806,N_19235);
nor U21111 (N_21111,N_19658,N_19442);
or U21112 (N_21112,N_19290,N_18930);
nor U21113 (N_21113,N_19121,N_19789);
nand U21114 (N_21114,N_19523,N_19626);
and U21115 (N_21115,N_19952,N_19657);
nand U21116 (N_21116,N_19611,N_18983);
nor U21117 (N_21117,N_19296,N_18826);
xnor U21118 (N_21118,N_19611,N_18993);
xnor U21119 (N_21119,N_18863,N_19270);
or U21120 (N_21120,N_18844,N_19967);
and U21121 (N_21121,N_19459,N_19027);
nor U21122 (N_21122,N_18782,N_19185);
nand U21123 (N_21123,N_19850,N_19417);
xor U21124 (N_21124,N_19918,N_19520);
xor U21125 (N_21125,N_19389,N_19868);
and U21126 (N_21126,N_19850,N_19196);
or U21127 (N_21127,N_19623,N_19933);
and U21128 (N_21128,N_19990,N_18973);
and U21129 (N_21129,N_19455,N_19365);
and U21130 (N_21130,N_19801,N_18790);
nand U21131 (N_21131,N_19141,N_18811);
and U21132 (N_21132,N_18901,N_19655);
nand U21133 (N_21133,N_19570,N_18940);
nand U21134 (N_21134,N_18825,N_19288);
xnor U21135 (N_21135,N_19616,N_19145);
or U21136 (N_21136,N_19664,N_19107);
nand U21137 (N_21137,N_19726,N_18936);
xor U21138 (N_21138,N_19852,N_19860);
nor U21139 (N_21139,N_19362,N_19311);
xor U21140 (N_21140,N_18819,N_18809);
nand U21141 (N_21141,N_19664,N_19643);
and U21142 (N_21142,N_19276,N_18863);
xnor U21143 (N_21143,N_19912,N_18857);
or U21144 (N_21144,N_19304,N_18926);
or U21145 (N_21145,N_18939,N_19281);
nor U21146 (N_21146,N_19633,N_19866);
nand U21147 (N_21147,N_19694,N_19925);
and U21148 (N_21148,N_18767,N_19005);
nand U21149 (N_21149,N_19349,N_19208);
xor U21150 (N_21150,N_19247,N_19296);
xor U21151 (N_21151,N_19188,N_19845);
nand U21152 (N_21152,N_19924,N_19494);
or U21153 (N_21153,N_19712,N_19842);
nor U21154 (N_21154,N_19935,N_19603);
and U21155 (N_21155,N_19135,N_19950);
nor U21156 (N_21156,N_19699,N_19020);
and U21157 (N_21157,N_19858,N_19570);
nor U21158 (N_21158,N_19075,N_19435);
nor U21159 (N_21159,N_19956,N_19572);
and U21160 (N_21160,N_18789,N_18809);
nand U21161 (N_21161,N_19423,N_19826);
and U21162 (N_21162,N_19733,N_18923);
or U21163 (N_21163,N_19283,N_19501);
and U21164 (N_21164,N_19464,N_19344);
nor U21165 (N_21165,N_19136,N_19611);
nor U21166 (N_21166,N_19051,N_18980);
nor U21167 (N_21167,N_19220,N_19436);
nor U21168 (N_21168,N_19633,N_19498);
nand U21169 (N_21169,N_18956,N_19895);
or U21170 (N_21170,N_19930,N_19694);
nand U21171 (N_21171,N_19212,N_19344);
xor U21172 (N_21172,N_18756,N_19128);
nor U21173 (N_21173,N_18808,N_19685);
nand U21174 (N_21174,N_19699,N_19214);
xor U21175 (N_21175,N_19811,N_18762);
nand U21176 (N_21176,N_18933,N_18985);
and U21177 (N_21177,N_19317,N_19816);
xnor U21178 (N_21178,N_19852,N_19302);
xor U21179 (N_21179,N_19439,N_19661);
nand U21180 (N_21180,N_19219,N_19894);
nor U21181 (N_21181,N_19356,N_19956);
and U21182 (N_21182,N_19834,N_19935);
and U21183 (N_21183,N_18871,N_19939);
nor U21184 (N_21184,N_19807,N_19897);
and U21185 (N_21185,N_19195,N_19076);
nand U21186 (N_21186,N_18978,N_19343);
or U21187 (N_21187,N_18896,N_19104);
and U21188 (N_21188,N_19530,N_19004);
nand U21189 (N_21189,N_19142,N_18962);
nand U21190 (N_21190,N_19905,N_19434);
nand U21191 (N_21191,N_19683,N_19529);
xnor U21192 (N_21192,N_18991,N_19074);
nand U21193 (N_21193,N_19736,N_19772);
xnor U21194 (N_21194,N_19936,N_19982);
and U21195 (N_21195,N_18959,N_19909);
and U21196 (N_21196,N_19466,N_19895);
xor U21197 (N_21197,N_19838,N_19327);
xnor U21198 (N_21198,N_19913,N_19697);
or U21199 (N_21199,N_19158,N_19526);
or U21200 (N_21200,N_19005,N_19119);
nand U21201 (N_21201,N_19050,N_19440);
and U21202 (N_21202,N_19922,N_19309);
xor U21203 (N_21203,N_19039,N_19970);
xnor U21204 (N_21204,N_19537,N_19804);
xor U21205 (N_21205,N_19303,N_19619);
or U21206 (N_21206,N_19366,N_18992);
and U21207 (N_21207,N_19149,N_18842);
or U21208 (N_21208,N_19148,N_19516);
nand U21209 (N_21209,N_19033,N_18979);
or U21210 (N_21210,N_19925,N_18939);
nor U21211 (N_21211,N_19652,N_19186);
xor U21212 (N_21212,N_19481,N_19260);
nand U21213 (N_21213,N_19260,N_19578);
xor U21214 (N_21214,N_19373,N_19875);
and U21215 (N_21215,N_19086,N_18768);
and U21216 (N_21216,N_19984,N_19694);
and U21217 (N_21217,N_19437,N_18755);
xnor U21218 (N_21218,N_18984,N_18879);
nor U21219 (N_21219,N_19100,N_19223);
nor U21220 (N_21220,N_19951,N_18854);
or U21221 (N_21221,N_18964,N_18808);
and U21222 (N_21222,N_19558,N_19130);
xor U21223 (N_21223,N_19652,N_18845);
nand U21224 (N_21224,N_19678,N_19578);
xnor U21225 (N_21225,N_19948,N_19959);
xor U21226 (N_21226,N_19583,N_18787);
and U21227 (N_21227,N_19573,N_19504);
or U21228 (N_21228,N_19348,N_19866);
and U21229 (N_21229,N_19286,N_18883);
or U21230 (N_21230,N_18964,N_18929);
xor U21231 (N_21231,N_19158,N_19944);
or U21232 (N_21232,N_19448,N_19406);
or U21233 (N_21233,N_19435,N_18958);
xor U21234 (N_21234,N_19797,N_19699);
or U21235 (N_21235,N_19325,N_19875);
and U21236 (N_21236,N_18998,N_18939);
and U21237 (N_21237,N_19643,N_19842);
nand U21238 (N_21238,N_18754,N_19354);
and U21239 (N_21239,N_19668,N_19368);
xor U21240 (N_21240,N_19663,N_19670);
and U21241 (N_21241,N_19476,N_19491);
or U21242 (N_21242,N_19640,N_19506);
nand U21243 (N_21243,N_19083,N_18793);
nor U21244 (N_21244,N_19704,N_19267);
xnor U21245 (N_21245,N_19594,N_18851);
and U21246 (N_21246,N_19428,N_19514);
nand U21247 (N_21247,N_19273,N_19173);
nor U21248 (N_21248,N_18839,N_19489);
xor U21249 (N_21249,N_19980,N_19637);
xnor U21250 (N_21250,N_20132,N_20412);
xor U21251 (N_21251,N_20750,N_21241);
nand U21252 (N_21252,N_20595,N_20910);
or U21253 (N_21253,N_20361,N_20809);
xor U21254 (N_21254,N_20548,N_20453);
nor U21255 (N_21255,N_20919,N_20095);
nor U21256 (N_21256,N_20534,N_20449);
and U21257 (N_21257,N_20835,N_21240);
nor U21258 (N_21258,N_20188,N_20732);
and U21259 (N_21259,N_20200,N_20345);
or U21260 (N_21260,N_21045,N_21246);
nor U21261 (N_21261,N_21162,N_20621);
nor U21262 (N_21262,N_20185,N_20176);
nand U21263 (N_21263,N_20522,N_20603);
nand U21264 (N_21264,N_20652,N_20695);
xor U21265 (N_21265,N_20861,N_20944);
nor U21266 (N_21266,N_20414,N_20799);
or U21267 (N_21267,N_20300,N_21029);
nor U21268 (N_21268,N_21225,N_20630);
xnor U21269 (N_21269,N_20313,N_21199);
and U21270 (N_21270,N_20633,N_20273);
nor U21271 (N_21271,N_20860,N_20417);
nand U21272 (N_21272,N_21100,N_20821);
or U21273 (N_21273,N_20933,N_20625);
nand U21274 (N_21274,N_20426,N_20685);
nand U21275 (N_21275,N_21202,N_20715);
nand U21276 (N_21276,N_20438,N_20015);
xor U21277 (N_21277,N_20986,N_20464);
or U21278 (N_21278,N_20932,N_20100);
xnor U21279 (N_21279,N_21012,N_21083);
or U21280 (N_21280,N_20960,N_21026);
nor U21281 (N_21281,N_21006,N_20131);
xor U21282 (N_21282,N_21076,N_20640);
xnor U21283 (N_21283,N_21066,N_21082);
nor U21284 (N_21284,N_20628,N_20043);
and U21285 (N_21285,N_20853,N_20612);
or U21286 (N_21286,N_20653,N_20891);
nand U21287 (N_21287,N_20526,N_20509);
and U21288 (N_21288,N_21158,N_20018);
nand U21289 (N_21289,N_20487,N_20316);
xnor U21290 (N_21290,N_20339,N_20463);
nor U21291 (N_21291,N_21098,N_20287);
xnor U21292 (N_21292,N_20848,N_20767);
nor U21293 (N_21293,N_20253,N_21064);
xnor U21294 (N_21294,N_20145,N_20571);
nor U21295 (N_21295,N_20052,N_20855);
nand U21296 (N_21296,N_20752,N_20322);
xor U21297 (N_21297,N_20122,N_20817);
or U21298 (N_21298,N_20574,N_20366);
nor U21299 (N_21299,N_20056,N_20275);
or U21300 (N_21300,N_20274,N_20500);
nand U21301 (N_21301,N_20777,N_20539);
nor U21302 (N_21302,N_20223,N_20538);
nor U21303 (N_21303,N_20250,N_20302);
nand U21304 (N_21304,N_20849,N_21192);
nand U21305 (N_21305,N_20121,N_20887);
nor U21306 (N_21306,N_20573,N_20111);
or U21307 (N_21307,N_20743,N_20189);
nor U21308 (N_21308,N_21173,N_20565);
xor U21309 (N_21309,N_21102,N_20995);
xnor U21310 (N_21310,N_20459,N_20832);
nor U21311 (N_21311,N_20976,N_20657);
or U21312 (N_21312,N_20577,N_20237);
nor U21313 (N_21313,N_20139,N_20785);
xor U21314 (N_21314,N_20601,N_20165);
nor U21315 (N_21315,N_20264,N_20478);
nor U21316 (N_21316,N_20896,N_20602);
or U21317 (N_21317,N_21129,N_20157);
xnor U21318 (N_21318,N_20590,N_20374);
or U21319 (N_21319,N_20702,N_20551);
nor U21320 (N_21320,N_21016,N_21092);
nand U21321 (N_21321,N_20135,N_20649);
or U21322 (N_21322,N_20061,N_20899);
nand U21323 (N_21323,N_20626,N_20928);
xnor U21324 (N_21324,N_20292,N_20236);
nand U21325 (N_21325,N_20248,N_20701);
xnor U21326 (N_21326,N_21094,N_21048);
nor U21327 (N_21327,N_20376,N_20040);
nand U21328 (N_21328,N_20498,N_20836);
nor U21329 (N_21329,N_20457,N_20915);
or U21330 (N_21330,N_20177,N_20941);
or U21331 (N_21331,N_21133,N_20337);
and U21332 (N_21332,N_20984,N_20954);
or U21333 (N_21333,N_20789,N_20619);
and U21334 (N_21334,N_20768,N_21034);
nor U21335 (N_21335,N_20399,N_20494);
xnor U21336 (N_21336,N_20639,N_21180);
and U21337 (N_21337,N_20097,N_21175);
nor U21338 (N_21338,N_20277,N_20142);
nor U21339 (N_21339,N_20021,N_20623);
nand U21340 (N_21340,N_20419,N_20053);
or U21341 (N_21341,N_20576,N_20323);
nor U21342 (N_21342,N_21024,N_21038);
xnor U21343 (N_21343,N_20301,N_21183);
or U21344 (N_21344,N_21090,N_20970);
and U21345 (N_21345,N_20925,N_20786);
or U21346 (N_21346,N_20327,N_20609);
and U21347 (N_21347,N_20181,N_20044);
and U21348 (N_21348,N_20811,N_20644);
nor U21349 (N_21349,N_20158,N_20171);
or U21350 (N_21350,N_20367,N_21197);
xnor U21351 (N_21351,N_20684,N_20369);
xor U21352 (N_21352,N_21109,N_20330);
nor U21353 (N_21353,N_20774,N_20807);
nor U21354 (N_21354,N_20133,N_20024);
and U21355 (N_21355,N_20047,N_20725);
xnor U21356 (N_21356,N_21243,N_20967);
nor U21357 (N_21357,N_20872,N_21237);
or U21358 (N_21358,N_21206,N_20069);
and U21359 (N_21359,N_20547,N_20077);
or U21360 (N_21360,N_20679,N_20140);
xnor U21361 (N_21361,N_20094,N_20445);
nor U21362 (N_21362,N_20583,N_20137);
nor U21363 (N_21363,N_20656,N_21155);
and U21364 (N_21364,N_20697,N_20898);
xnor U21365 (N_21365,N_20519,N_21138);
nand U21366 (N_21366,N_20813,N_20654);
nor U21367 (N_21367,N_20761,N_20863);
and U21368 (N_21368,N_20229,N_20895);
xor U21369 (N_21369,N_20477,N_20616);
or U21370 (N_21370,N_21063,N_20035);
nand U21371 (N_21371,N_21157,N_21084);
and U21372 (N_21372,N_20845,N_20969);
nor U21373 (N_21373,N_20627,N_20127);
and U21374 (N_21374,N_20674,N_20672);
nand U21375 (N_21375,N_20398,N_20224);
and U21376 (N_21376,N_20029,N_20413);
or U21377 (N_21377,N_20942,N_20671);
xor U21378 (N_21378,N_20559,N_21242);
or U21379 (N_21379,N_20308,N_20461);
and U21380 (N_21380,N_21010,N_21214);
nor U21381 (N_21381,N_20001,N_21050);
nand U21382 (N_21382,N_20924,N_20387);
nor U21383 (N_21383,N_20496,N_20349);
and U21384 (N_21384,N_21247,N_20102);
xnor U21385 (N_21385,N_20825,N_20113);
and U21386 (N_21386,N_20246,N_21115);
or U21387 (N_21387,N_21211,N_21161);
and U21388 (N_21388,N_20989,N_20422);
and U21389 (N_21389,N_20578,N_20555);
or U21390 (N_21390,N_20878,N_21233);
or U21391 (N_21391,N_21124,N_20546);
xnor U21392 (N_21392,N_20691,N_20085);
xor U21393 (N_21393,N_21198,N_20631);
nand U21394 (N_21394,N_20260,N_20110);
or U21395 (N_21395,N_20869,N_20641);
or U21396 (N_21396,N_20472,N_20421);
or U21397 (N_21397,N_20103,N_20004);
nand U21398 (N_21398,N_20938,N_21120);
and U21399 (N_21399,N_20501,N_20937);
or U21400 (N_21400,N_20713,N_20823);
nor U21401 (N_21401,N_20981,N_21108);
nand U21402 (N_21402,N_20884,N_21135);
nor U21403 (N_21403,N_21139,N_20202);
nand U21404 (N_21404,N_20549,N_20356);
nor U21405 (N_21405,N_20288,N_21014);
nand U21406 (N_21406,N_20267,N_20770);
and U21407 (N_21407,N_20423,N_20411);
or U21408 (N_21408,N_20726,N_20124);
and U21409 (N_21409,N_20152,N_20829);
nor U21410 (N_21410,N_20531,N_20658);
or U21411 (N_21411,N_20585,N_20739);
nor U21412 (N_21412,N_20076,N_20544);
or U21413 (N_21413,N_20050,N_20673);
nand U21414 (N_21414,N_20067,N_20384);
nor U21415 (N_21415,N_21223,N_20675);
nand U21416 (N_21416,N_21193,N_20561);
nand U21417 (N_21417,N_20988,N_20580);
xnor U21418 (N_21418,N_20192,N_20473);
and U21419 (N_21419,N_21166,N_20827);
nor U21420 (N_21420,N_20241,N_20587);
nand U21421 (N_21421,N_20305,N_20800);
and U21422 (N_21422,N_20866,N_21191);
xor U21423 (N_21423,N_20998,N_20940);
xor U21424 (N_21424,N_20416,N_20014);
and U21425 (N_21425,N_20705,N_20234);
xor U21426 (N_21426,N_20003,N_20523);
nor U21427 (N_21427,N_20407,N_20424);
and U21428 (N_21428,N_20430,N_20450);
or U21429 (N_21429,N_20146,N_20824);
xor U21430 (N_21430,N_20734,N_21232);
and U21431 (N_21431,N_20930,N_20517);
nor U21432 (N_21432,N_20272,N_20092);
nand U21433 (N_21433,N_20155,N_20346);
nor U21434 (N_21434,N_20638,N_20106);
and U21435 (N_21435,N_20208,N_20452);
and U21436 (N_21436,N_20364,N_20900);
or U21437 (N_21437,N_21196,N_20291);
nand U21438 (N_21438,N_20530,N_20432);
nand U21439 (N_21439,N_21058,N_20741);
or U21440 (N_21440,N_20048,N_20012);
xnor U21441 (N_21441,N_21235,N_20889);
or U21442 (N_21442,N_20022,N_20391);
nor U21443 (N_21443,N_20947,N_20843);
xnor U21444 (N_21444,N_21176,N_20475);
xnor U21445 (N_21445,N_20107,N_20826);
nor U21446 (N_21446,N_20228,N_21207);
xnor U21447 (N_21447,N_20607,N_20041);
xor U21448 (N_21448,N_20214,N_21087);
or U21449 (N_21449,N_20147,N_20591);
or U21450 (N_21450,N_20286,N_20666);
and U21451 (N_21451,N_20222,N_20920);
or U21452 (N_21452,N_20632,N_20386);
nand U21453 (N_21453,N_21230,N_20525);
nand U21454 (N_21454,N_20502,N_20730);
nor U21455 (N_21455,N_21085,N_21042);
or U21456 (N_21456,N_20762,N_21226);
xor U21457 (N_21457,N_20328,N_20815);
nor U21458 (N_21458,N_20667,N_20303);
nand U21459 (N_21459,N_20117,N_20388);
and U21460 (N_21460,N_20819,N_21143);
nor U21461 (N_21461,N_21080,N_20045);
nand U21462 (N_21462,N_20299,N_21031);
or U21463 (N_21463,N_21132,N_20447);
and U21464 (N_21464,N_20440,N_20216);
xor U21465 (N_21465,N_21041,N_20678);
or U21466 (N_21466,N_20212,N_20569);
xnor U21467 (N_21467,N_20535,N_20245);
xnor U21468 (N_21468,N_20233,N_20252);
and U21469 (N_21469,N_20199,N_20646);
or U21470 (N_21470,N_20467,N_20443);
and U21471 (N_21471,N_20870,N_20518);
and U21472 (N_21472,N_21249,N_20304);
nor U21473 (N_21473,N_20007,N_20629);
and U21474 (N_21474,N_20926,N_20951);
nand U21475 (N_21475,N_20722,N_20642);
or U21476 (N_21476,N_20842,N_20894);
xnor U21477 (N_21477,N_20793,N_20972);
nand U21478 (N_21478,N_20383,N_20125);
or U21479 (N_21479,N_20284,N_20016);
or U21480 (N_21480,N_21178,N_21224);
nor U21481 (N_21481,N_20348,N_20008);
xor U21482 (N_21482,N_20660,N_20936);
or U21483 (N_21483,N_21111,N_21156);
or U21484 (N_21484,N_20822,N_20462);
xnor U21485 (N_21485,N_20737,N_20070);
xor U21486 (N_21486,N_20352,N_20394);
and U21487 (N_21487,N_20655,N_21027);
and U21488 (N_21488,N_20903,N_20074);
and U21489 (N_21489,N_20586,N_20410);
xor U21490 (N_21490,N_20027,N_21163);
nand U21491 (N_21491,N_20227,N_20271);
or U21492 (N_21492,N_20888,N_20039);
xor U21493 (N_21493,N_20957,N_20448);
and U21494 (N_21494,N_20451,N_20792);
nand U21495 (N_21495,N_20818,N_20584);
and U21496 (N_21496,N_20688,N_20243);
xor U21497 (N_21497,N_20484,N_20321);
xnor U21498 (N_21498,N_20690,N_21072);
or U21499 (N_21499,N_21073,N_21051);
nand U21500 (N_21500,N_20203,N_20643);
or U21501 (N_21501,N_20508,N_20195);
nor U21502 (N_21502,N_20921,N_20814);
or U21503 (N_21503,N_20446,N_20144);
or U21504 (N_21504,N_21053,N_21079);
and U21505 (N_21505,N_20808,N_21170);
and U21506 (N_21506,N_20992,N_21150);
and U21507 (N_21507,N_21062,N_21218);
or U21508 (N_21508,N_20901,N_20317);
nor U21509 (N_21509,N_21043,N_20439);
nor U21510 (N_21510,N_20949,N_21127);
nand U21511 (N_21511,N_20648,N_20908);
nor U21512 (N_21512,N_20834,N_20733);
nor U21513 (N_21513,N_20444,N_20128);
nor U21514 (N_21514,N_21236,N_20686);
and U21515 (N_21515,N_20120,N_20182);
xor U21516 (N_21516,N_21091,N_20917);
xnor U21517 (N_21517,N_20326,N_20180);
xor U21518 (N_21518,N_20075,N_20063);
or U21519 (N_21519,N_20210,N_20226);
or U21520 (N_21520,N_20716,N_20060);
nor U21521 (N_21521,N_20592,N_20804);
nand U21522 (N_21522,N_20886,N_20955);
nand U21523 (N_21523,N_21118,N_20184);
and U21524 (N_21524,N_21044,N_20454);
nand U21525 (N_21525,N_20282,N_20495);
xor U21526 (N_21526,N_21131,N_20026);
nand U21527 (N_21527,N_20347,N_20794);
nor U21528 (N_21528,N_20400,N_20588);
xnor U21529 (N_21529,N_20997,N_20706);
nor U21530 (N_21530,N_21159,N_20542);
nand U21531 (N_21531,N_21033,N_21106);
nor U21532 (N_21532,N_20086,N_21081);
nor U21533 (N_21533,N_20953,N_20456);
nor U21534 (N_21534,N_20709,N_20885);
or U21535 (N_21535,N_20359,N_20033);
and U21536 (N_21536,N_20693,N_20806);
xnor U21537 (N_21537,N_20516,N_21182);
nand U21538 (N_21538,N_20431,N_21149);
xor U21539 (N_21539,N_20636,N_20711);
xor U21540 (N_21540,N_20563,N_20665);
xor U21541 (N_21541,N_20554,N_21221);
nor U21542 (N_21542,N_20880,N_21007);
nand U21543 (N_21543,N_20193,N_20064);
nor U21544 (N_21544,N_20011,N_20134);
xnor U21545 (N_21545,N_20186,N_21037);
nor U21546 (N_21546,N_20831,N_20882);
xnor U21547 (N_21547,N_20093,N_20335);
and U21548 (N_21548,N_21171,N_20999);
nor U21549 (N_21549,N_20079,N_20281);
and U21550 (N_21550,N_20010,N_20468);
nand U21551 (N_21551,N_20916,N_21018);
nor U21552 (N_21552,N_20191,N_20763);
or U21553 (N_21553,N_20433,N_20482);
nor U21554 (N_21554,N_20857,N_20506);
nand U21555 (N_21555,N_21238,N_21035);
and U21556 (N_21556,N_21056,N_20707);
nor U21557 (N_21557,N_20676,N_20279);
nand U21558 (N_21558,N_20381,N_20036);
nand U21559 (N_21559,N_20511,N_20718);
or U21560 (N_21560,N_20395,N_20694);
nand U21561 (N_21561,N_20973,N_21105);
or U21562 (N_21562,N_20278,N_20594);
and U21563 (N_21563,N_20390,N_20820);
nor U21564 (N_21564,N_20298,N_20854);
or U21565 (N_21565,N_20748,N_21144);
nor U21566 (N_21566,N_20909,N_20119);
nand U21567 (N_21567,N_21104,N_20727);
xnor U21568 (N_21568,N_21172,N_20049);
xnor U21569 (N_21569,N_20261,N_21039);
nand U21570 (N_21570,N_20368,N_20315);
and U21571 (N_21571,N_20198,N_20662);
or U21572 (N_21572,N_20168,N_20558);
xnor U21573 (N_21573,N_20507,N_20084);
nand U21574 (N_21574,N_21187,N_21119);
nand U21575 (N_21575,N_21055,N_20950);
or U21576 (N_21576,N_20114,N_20745);
and U21577 (N_21577,N_21116,N_20377);
nor U21578 (N_21578,N_20054,N_20217);
nor U21579 (N_21579,N_20780,N_20797);
and U21580 (N_21580,N_20108,N_20276);
nand U21581 (N_21581,N_21030,N_20397);
nand U21582 (N_21582,N_20991,N_20392);
xnor U21583 (N_21583,N_20087,N_20977);
nand U21584 (N_21584,N_20159,N_20597);
and U21585 (N_21585,N_20204,N_20721);
nor U21586 (N_21586,N_20669,N_20408);
or U21587 (N_21587,N_20828,N_20002);
nand U21588 (N_21588,N_20247,N_20295);
nor U21589 (N_21589,N_20615,N_20744);
and U21590 (N_21590,N_20309,N_21239);
and U21591 (N_21591,N_20689,N_21220);
nor U21592 (N_21592,N_20329,N_20883);
xnor U21593 (N_21593,N_20428,N_20375);
and U21594 (N_21594,N_20757,N_20393);
nand U21595 (N_21595,N_20194,N_20251);
nor U21596 (N_21596,N_20486,N_21216);
and U21597 (N_21597,N_20668,N_21137);
nand U21598 (N_21598,N_21074,N_21046);
nor U21599 (N_21599,N_20164,N_20455);
xnor U21600 (N_21600,N_20196,N_20927);
nor U21601 (N_21601,N_20283,N_20324);
or U21602 (N_21602,N_20850,N_20028);
or U21603 (N_21603,N_20610,N_21164);
nand U21604 (N_21604,N_20332,N_20256);
and U21605 (N_21605,N_20471,N_20751);
nor U21606 (N_21606,N_20810,N_20837);
xor U21607 (N_21607,N_20982,N_20425);
or U21608 (N_21608,N_20240,N_20568);
or U21609 (N_21609,N_20442,N_20116);
nand U21610 (N_21610,N_21068,N_20754);
nand U21611 (N_21611,N_21101,N_21141);
or U21612 (N_21612,N_20065,N_21205);
and U21613 (N_21613,N_20218,N_20851);
nand U21614 (N_21614,N_21152,N_20469);
nor U21615 (N_21615,N_20362,N_20781);
xor U21616 (N_21616,N_21126,N_20118);
xor U21617 (N_21617,N_21169,N_20696);
nor U21618 (N_21618,N_21017,N_21234);
nand U21619 (N_21619,N_21036,N_20966);
xor U21620 (N_21620,N_20728,N_20876);
and U21621 (N_21621,N_20358,N_21165);
xnor U21622 (N_21622,N_20081,N_20841);
and U21623 (N_21623,N_20839,N_20401);
nand U21624 (N_21624,N_20746,N_21136);
or U21625 (N_21625,N_20952,N_21013);
and U21626 (N_21626,N_21028,N_20692);
nor U21627 (N_21627,N_20700,N_20929);
or U21628 (N_21628,N_20080,N_20360);
nor U21629 (N_21629,N_21107,N_21020);
or U21630 (N_21630,N_20071,N_20566);
and U21631 (N_21631,N_20101,N_20156);
nand U21632 (N_21632,N_21059,N_20460);
or U21633 (N_21633,N_20520,N_20123);
and U21634 (N_21634,N_20637,N_21248);
nand U21635 (N_21635,N_20138,N_20167);
xnor U21636 (N_21636,N_20230,N_20338);
nor U21637 (N_21637,N_21130,N_20766);
and U21638 (N_21638,N_20310,N_20906);
or U21639 (N_21639,N_21004,N_20923);
xor U21640 (N_21640,N_20357,N_20319);
or U21641 (N_21641,N_20334,N_21002);
nand U21642 (N_21642,N_20914,N_20971);
xnor U21643 (N_21643,N_20801,N_20046);
nor U21644 (N_21644,N_20088,N_20557);
nor U21645 (N_21645,N_20205,N_20773);
nand U21646 (N_21646,N_20805,N_20765);
and U21647 (N_21647,N_20622,N_20979);
xnor U21648 (N_21648,N_21145,N_21070);
or U21649 (N_21649,N_21114,N_21154);
nor U21650 (N_21650,N_20847,N_20042);
nand U21651 (N_21651,N_20651,N_20680);
nand U21652 (N_21652,N_20232,N_20055);
or U21653 (N_21653,N_21209,N_20758);
and U21654 (N_21654,N_21177,N_21009);
xnor U21655 (N_21655,N_20211,N_20596);
xor U21656 (N_21656,N_20254,N_20497);
nand U21657 (N_21657,N_21054,N_20796);
nand U21658 (N_21658,N_20434,N_21121);
xor U21659 (N_21659,N_20013,N_20403);
nor U21660 (N_21660,N_20710,N_20527);
nor U21661 (N_21661,N_20025,N_20150);
xnor U21662 (N_21662,N_20803,N_20488);
nor U21663 (N_21663,N_20239,N_20838);
xnor U21664 (N_21664,N_20479,N_20840);
or U21665 (N_21665,N_20354,N_20420);
nor U21666 (N_21666,N_20220,N_20066);
xor U21667 (N_21667,N_20183,N_20249);
nor U21668 (N_21668,N_20436,N_20545);
or U21669 (N_21669,N_20373,N_20405);
or U21670 (N_21670,N_20023,N_20723);
nor U21671 (N_21671,N_20173,N_20537);
nand U21672 (N_21672,N_20570,N_20513);
xnor U21673 (N_21673,N_20599,N_21174);
xnor U21674 (N_21674,N_20959,N_20489);
or U21675 (N_21675,N_20802,N_21201);
xnor U21676 (N_21676,N_20058,N_20474);
and U21677 (N_21677,N_20130,N_20149);
or U21678 (N_21678,N_20485,N_20409);
or U21679 (N_21679,N_20020,N_20956);
and U21680 (N_21680,N_21067,N_21060);
or U21681 (N_21681,N_20795,N_21231);
or U21682 (N_21682,N_20491,N_21204);
nand U21683 (N_21683,N_20415,N_20670);
or U21684 (N_21684,N_20681,N_21000);
xnor U21685 (N_21685,N_21244,N_20983);
and U21686 (N_21686,N_20148,N_21167);
nand U21687 (N_21687,N_20550,N_20975);
xor U21688 (N_21688,N_21122,N_21003);
and U21689 (N_21689,N_20017,N_20962);
xnor U21690 (N_21690,N_20564,N_20790);
nand U21691 (N_21691,N_21185,N_20812);
nor U21692 (N_21692,N_20890,N_20037);
and U21693 (N_21693,N_21179,N_20963);
or U21694 (N_21694,N_20618,N_20704);
and U21695 (N_21695,N_21181,N_20858);
xnor U21696 (N_21696,N_20109,N_20179);
nor U21697 (N_21697,N_20242,N_20892);
xor U21698 (N_21698,N_20816,N_20904);
nor U21699 (N_21699,N_20141,N_21065);
nand U21700 (N_21700,N_20871,N_21245);
nand U21701 (N_21701,N_20213,N_20342);
nor U21702 (N_21702,N_21140,N_20783);
nand U21703 (N_21703,N_21194,N_20160);
nor U21704 (N_21704,N_20856,N_20782);
xor U21705 (N_21705,N_20572,N_20378);
nor U21706 (N_21706,N_21147,N_20905);
or U21707 (N_21707,N_20257,N_20867);
xnor U21708 (N_21708,N_20073,N_21021);
nand U21709 (N_21709,N_20922,N_20505);
xnor U21710 (N_21710,N_20533,N_21215);
xor U21711 (N_21711,N_21189,N_20404);
nor U21712 (N_21712,N_20169,N_20661);
and U21713 (N_21713,N_21015,N_20980);
nand U21714 (N_21714,N_20089,N_20083);
nand U21715 (N_21715,N_21123,N_20514);
and U21716 (N_21716,N_20787,N_21168);
or U21717 (N_21717,N_20262,N_20943);
xor U21718 (N_21718,N_21151,N_21184);
or U21719 (N_21719,N_21097,N_20510);
nand U21720 (N_21720,N_21103,N_20747);
or U21721 (N_21721,N_20593,N_20833);
and U21722 (N_21722,N_20504,N_20341);
nand U21723 (N_21723,N_20325,N_20552);
xnor U21724 (N_21724,N_21160,N_20206);
or U21725 (N_21725,N_21093,N_20540);
nand U21726 (N_21726,N_21228,N_21019);
nand U21727 (N_21727,N_20624,N_20515);
xnor U21728 (N_21728,N_21110,N_21089);
nand U21729 (N_21729,N_20389,N_20994);
and U21730 (N_21730,N_20598,N_20340);
nand U21731 (N_21731,N_21069,N_20483);
xor U21732 (N_21732,N_20659,N_20082);
nand U21733 (N_21733,N_20296,N_20788);
and U21734 (N_21734,N_20311,N_20996);
or U21735 (N_21735,N_20865,N_20215);
xnor U21736 (N_21736,N_20458,N_21217);
nand U21737 (N_21737,N_20503,N_21047);
xnor U21738 (N_21738,N_20990,N_21210);
and U21739 (N_21739,N_21057,N_20611);
xnor U21740 (N_21740,N_20059,N_20019);
and U21741 (N_21741,N_20154,N_20553);
nand U21742 (N_21742,N_20427,N_21148);
nor U21743 (N_21743,N_20562,N_20532);
nand U21744 (N_21744,N_21208,N_20269);
nand U21745 (N_21745,N_21146,N_20371);
and U21746 (N_21746,N_20351,N_20143);
and U21747 (N_21747,N_20556,N_20604);
or U21748 (N_21748,N_20355,N_21061);
or U21749 (N_21749,N_20703,N_20776);
xnor U21750 (N_21750,N_20480,N_20072);
or U21751 (N_21751,N_20978,N_20172);
xor U21752 (N_21752,N_20779,N_20099);
nor U21753 (N_21753,N_20965,N_21190);
nor U21754 (N_21754,N_20034,N_20698);
or U21755 (N_21755,N_20333,N_20492);
nand U21756 (N_21756,N_21032,N_20353);
nand U21757 (N_21757,N_20499,N_20778);
or U21758 (N_21758,N_21203,N_21112);
or U21759 (N_21759,N_20062,N_20740);
nand U21760 (N_21760,N_20945,N_20129);
nor U21761 (N_21761,N_20879,N_20589);
or U21762 (N_21762,N_20005,N_21005);
nor U21763 (N_21763,N_20372,N_20466);
nor U21764 (N_21764,N_20418,N_20582);
nand U21765 (N_21765,N_20717,N_20235);
nor U21766 (N_21766,N_20755,N_20798);
or U21767 (N_21767,N_20512,N_21142);
and U21768 (N_21768,N_20529,N_20528);
xnor U21769 (N_21769,N_20859,N_21071);
nor U21770 (N_21770,N_20521,N_21212);
nand U21771 (N_21771,N_21095,N_20687);
nand U21772 (N_21772,N_20314,N_20536);
or U21773 (N_21773,N_20365,N_20197);
nand U21774 (N_21774,N_21113,N_20280);
xor U21775 (N_21775,N_20724,N_20363);
and U21776 (N_21776,N_20096,N_21025);
xor U21777 (N_21777,N_20575,N_21040);
xnor U21778 (N_21778,N_20151,N_20429);
xnor U21779 (N_21779,N_20320,N_20201);
and U21780 (N_21780,N_20470,N_20907);
xor U21781 (N_21781,N_20613,N_21052);
nor U21782 (N_21782,N_20078,N_20958);
xor U21783 (N_21783,N_20465,N_20712);
or U21784 (N_21784,N_20009,N_20875);
nor U21785 (N_21785,N_20476,N_20708);
nand U21786 (N_21786,N_20581,N_21075);
nor U21787 (N_21787,N_20350,N_20178);
and U21788 (N_21788,N_20560,N_20961);
or U21789 (N_21789,N_20830,N_20221);
xor U21790 (N_21790,N_20934,N_21229);
nor U21791 (N_21791,N_20968,N_20153);
or U21792 (N_21792,N_21200,N_20030);
xor U21793 (N_21793,N_20608,N_20862);
xor U21794 (N_21794,N_21077,N_20864);
or U21795 (N_21795,N_20911,N_21011);
or U21796 (N_21796,N_20162,N_20606);
and U21797 (N_21797,N_20974,N_21186);
or U21798 (N_21798,N_20791,N_20370);
nor U21799 (N_21799,N_20231,N_20614);
or U21800 (N_21800,N_20759,N_20948);
nor U21801 (N_21801,N_20174,N_20756);
and U21802 (N_21802,N_20844,N_21188);
nor U21803 (N_21803,N_21227,N_20306);
or U21804 (N_21804,N_20382,N_20912);
nor U21805 (N_21805,N_20285,N_20946);
or U21806 (N_21806,N_21128,N_20935);
and U21807 (N_21807,N_20881,N_20207);
nand U21808 (N_21808,N_20993,N_20318);
nor U21809 (N_21809,N_20719,N_20209);
nand U21810 (N_21810,N_20913,N_20939);
nor U21811 (N_21811,N_20259,N_20775);
nand U21812 (N_21812,N_20057,N_21088);
xnor U21813 (N_21813,N_20493,N_20105);
and U21814 (N_21814,N_20380,N_20987);
or U21815 (N_21815,N_20931,N_20297);
xnor U21816 (N_21816,N_20255,N_20406);
nor U21817 (N_21817,N_20006,N_21022);
or U21818 (N_21818,N_20543,N_20266);
and U21819 (N_21819,N_20343,N_20112);
and U21820 (N_21820,N_20481,N_20735);
nand U21821 (N_21821,N_20714,N_20238);
and U21822 (N_21822,N_20868,N_20163);
and U21823 (N_21823,N_20225,N_20265);
xnor U21824 (N_21824,N_20000,N_21134);
or U21825 (N_21825,N_20720,N_20038);
nor U21826 (N_21826,N_21078,N_20290);
or U21827 (N_21827,N_20031,N_20874);
nor U21828 (N_21828,N_20769,N_21086);
nand U21829 (N_21829,N_20051,N_20270);
nor U21830 (N_21830,N_20902,N_20136);
nor U21831 (N_21831,N_20258,N_20682);
xor U21832 (N_21832,N_20873,N_20918);
nand U21833 (N_21833,N_20650,N_20579);
or U21834 (N_21834,N_20749,N_20645);
nand U21835 (N_21835,N_20396,N_21023);
and U21836 (N_21836,N_20091,N_20731);
or U21837 (N_21837,N_20032,N_20312);
and U21838 (N_21838,N_20664,N_20647);
or U21839 (N_21839,N_20336,N_20760);
or U21840 (N_21840,N_21096,N_20736);
and U21841 (N_21841,N_20772,N_20897);
or U21842 (N_21842,N_21099,N_21125);
or U21843 (N_21843,N_20683,N_20437);
nand U21844 (N_21844,N_21195,N_20634);
nor U21845 (N_21845,N_20090,N_20379);
xnor U21846 (N_21846,N_20753,N_20244);
or U21847 (N_21847,N_21049,N_20729);
and U21848 (N_21848,N_20742,N_20764);
nand U21849 (N_21849,N_21117,N_20605);
or U21850 (N_21850,N_20490,N_20293);
or U21851 (N_21851,N_20964,N_20846);
nor U21852 (N_21852,N_20263,N_20541);
and U21853 (N_21853,N_20784,N_20600);
nand U21854 (N_21854,N_20268,N_20175);
nor U21855 (N_21855,N_20877,N_20187);
and U21856 (N_21856,N_21222,N_20677);
nor U21857 (N_21857,N_20190,N_21008);
or U21858 (N_21858,N_20771,N_20289);
or U21859 (N_21859,N_20441,N_20617);
or U21860 (N_21860,N_20294,N_20567);
and U21861 (N_21861,N_21153,N_20635);
and U21862 (N_21862,N_20985,N_20402);
nand U21863 (N_21863,N_20435,N_20385);
or U21864 (N_21864,N_20170,N_20344);
nand U21865 (N_21865,N_20663,N_20620);
nand U21866 (N_21866,N_20098,N_21213);
xor U21867 (N_21867,N_20068,N_20307);
and U21868 (N_21868,N_20524,N_20852);
and U21869 (N_21869,N_20738,N_21219);
nor U21870 (N_21870,N_20104,N_21001);
xor U21871 (N_21871,N_20219,N_20115);
nand U21872 (N_21872,N_20126,N_20331);
xnor U21873 (N_21873,N_20699,N_20161);
and U21874 (N_21874,N_20166,N_20893);
nor U21875 (N_21875,N_20902,N_20627);
and U21876 (N_21876,N_21167,N_20030);
or U21877 (N_21877,N_21049,N_20119);
nor U21878 (N_21878,N_20206,N_20010);
and U21879 (N_21879,N_20929,N_20423);
and U21880 (N_21880,N_20730,N_21142);
nor U21881 (N_21881,N_20324,N_20331);
and U21882 (N_21882,N_20554,N_20686);
and U21883 (N_21883,N_20986,N_20293);
nand U21884 (N_21884,N_20817,N_20523);
and U21885 (N_21885,N_20381,N_20331);
and U21886 (N_21886,N_20805,N_20057);
and U21887 (N_21887,N_20734,N_20186);
or U21888 (N_21888,N_20387,N_21207);
xor U21889 (N_21889,N_20880,N_20850);
xor U21890 (N_21890,N_20711,N_21140);
or U21891 (N_21891,N_20592,N_21163);
xnor U21892 (N_21892,N_21017,N_20567);
nand U21893 (N_21893,N_20970,N_20243);
or U21894 (N_21894,N_20496,N_20059);
nand U21895 (N_21895,N_20496,N_20702);
and U21896 (N_21896,N_20032,N_20178);
xnor U21897 (N_21897,N_20317,N_20852);
nand U21898 (N_21898,N_20713,N_20854);
xor U21899 (N_21899,N_20184,N_20662);
and U21900 (N_21900,N_20175,N_20467);
nand U21901 (N_21901,N_20036,N_20747);
nor U21902 (N_21902,N_20648,N_20718);
nand U21903 (N_21903,N_20461,N_21093);
nand U21904 (N_21904,N_21179,N_20391);
or U21905 (N_21905,N_21139,N_21144);
and U21906 (N_21906,N_20375,N_20121);
nand U21907 (N_21907,N_20443,N_20273);
and U21908 (N_21908,N_20991,N_20699);
nand U21909 (N_21909,N_20774,N_20337);
nand U21910 (N_21910,N_20716,N_20027);
nor U21911 (N_21911,N_20317,N_20446);
xor U21912 (N_21912,N_20929,N_20908);
or U21913 (N_21913,N_20546,N_20499);
xor U21914 (N_21914,N_21085,N_20199);
nor U21915 (N_21915,N_20683,N_21076);
and U21916 (N_21916,N_20354,N_20928);
xnor U21917 (N_21917,N_21124,N_20602);
or U21918 (N_21918,N_20303,N_20740);
and U21919 (N_21919,N_20605,N_20251);
or U21920 (N_21920,N_21102,N_21005);
and U21921 (N_21921,N_21029,N_20139);
nor U21922 (N_21922,N_20775,N_20011);
or U21923 (N_21923,N_21177,N_20464);
or U21924 (N_21924,N_20085,N_20278);
nor U21925 (N_21925,N_20938,N_21104);
or U21926 (N_21926,N_21137,N_20625);
and U21927 (N_21927,N_20746,N_21113);
nand U21928 (N_21928,N_20805,N_20415);
nor U21929 (N_21929,N_20862,N_20978);
nand U21930 (N_21930,N_20513,N_21083);
nor U21931 (N_21931,N_20230,N_20911);
xnor U21932 (N_21932,N_20393,N_20325);
or U21933 (N_21933,N_20713,N_21144);
nor U21934 (N_21934,N_20944,N_20400);
nand U21935 (N_21935,N_20168,N_20933);
xor U21936 (N_21936,N_20213,N_21164);
xnor U21937 (N_21937,N_20613,N_20136);
xnor U21938 (N_21938,N_20393,N_20070);
and U21939 (N_21939,N_20723,N_20974);
and U21940 (N_21940,N_20271,N_20881);
xor U21941 (N_21941,N_20978,N_20629);
nor U21942 (N_21942,N_20545,N_20019);
nor U21943 (N_21943,N_20529,N_20525);
nor U21944 (N_21944,N_20187,N_20546);
and U21945 (N_21945,N_20532,N_20554);
or U21946 (N_21946,N_21235,N_20536);
and U21947 (N_21947,N_20857,N_20460);
or U21948 (N_21948,N_20420,N_20408);
nor U21949 (N_21949,N_20741,N_20341);
nand U21950 (N_21950,N_20293,N_20963);
and U21951 (N_21951,N_20253,N_21165);
nand U21952 (N_21952,N_21167,N_20441);
xor U21953 (N_21953,N_20752,N_20125);
xor U21954 (N_21954,N_20040,N_20889);
xor U21955 (N_21955,N_20104,N_20714);
nand U21956 (N_21956,N_20653,N_21205);
and U21957 (N_21957,N_20012,N_20546);
or U21958 (N_21958,N_20084,N_20642);
nor U21959 (N_21959,N_20253,N_20104);
xnor U21960 (N_21960,N_20530,N_20459);
nand U21961 (N_21961,N_20917,N_21151);
xnor U21962 (N_21962,N_20470,N_21094);
xnor U21963 (N_21963,N_20880,N_20315);
or U21964 (N_21964,N_20966,N_21022);
nor U21965 (N_21965,N_20424,N_20651);
or U21966 (N_21966,N_21052,N_20046);
or U21967 (N_21967,N_20837,N_20003);
and U21968 (N_21968,N_20471,N_20563);
nor U21969 (N_21969,N_21065,N_20514);
or U21970 (N_21970,N_21229,N_20157);
or U21971 (N_21971,N_20130,N_20160);
nand U21972 (N_21972,N_20988,N_20235);
xor U21973 (N_21973,N_21216,N_20888);
and U21974 (N_21974,N_20440,N_20486);
xor U21975 (N_21975,N_20691,N_20805);
or U21976 (N_21976,N_20935,N_20565);
nor U21977 (N_21977,N_20139,N_20118);
xor U21978 (N_21978,N_20358,N_20017);
and U21979 (N_21979,N_20523,N_20732);
xor U21980 (N_21980,N_20957,N_20009);
nand U21981 (N_21981,N_20278,N_20481);
xnor U21982 (N_21982,N_20796,N_20728);
xnor U21983 (N_21983,N_20536,N_20809);
and U21984 (N_21984,N_20743,N_21210);
nor U21985 (N_21985,N_21170,N_20853);
xor U21986 (N_21986,N_21010,N_20101);
xnor U21987 (N_21987,N_20677,N_20322);
nor U21988 (N_21988,N_20086,N_20846);
and U21989 (N_21989,N_20246,N_20971);
nor U21990 (N_21990,N_20760,N_20311);
nand U21991 (N_21991,N_20775,N_21095);
nor U21992 (N_21992,N_20148,N_20565);
xor U21993 (N_21993,N_20775,N_20018);
xor U21994 (N_21994,N_20700,N_20196);
nand U21995 (N_21995,N_20997,N_20527);
xnor U21996 (N_21996,N_20141,N_20423);
and U21997 (N_21997,N_20487,N_20699);
nand U21998 (N_21998,N_21149,N_20135);
nor U21999 (N_21999,N_20569,N_20171);
nor U22000 (N_22000,N_20630,N_20003);
nand U22001 (N_22001,N_20301,N_20855);
nand U22002 (N_22002,N_20246,N_20470);
nor U22003 (N_22003,N_21005,N_20907);
nor U22004 (N_22004,N_20686,N_20151);
xor U22005 (N_22005,N_21029,N_20860);
xnor U22006 (N_22006,N_21138,N_21050);
xor U22007 (N_22007,N_20441,N_20864);
and U22008 (N_22008,N_21103,N_21066);
or U22009 (N_22009,N_20703,N_21037);
or U22010 (N_22010,N_20885,N_21103);
xnor U22011 (N_22011,N_20137,N_20946);
xnor U22012 (N_22012,N_20345,N_20396);
and U22013 (N_22013,N_20101,N_20091);
nand U22014 (N_22014,N_20326,N_21100);
and U22015 (N_22015,N_20099,N_21215);
nand U22016 (N_22016,N_20467,N_20092);
or U22017 (N_22017,N_20875,N_20636);
xor U22018 (N_22018,N_20569,N_20434);
or U22019 (N_22019,N_21005,N_20714);
nor U22020 (N_22020,N_20509,N_20109);
and U22021 (N_22021,N_21080,N_20026);
and U22022 (N_22022,N_20222,N_20332);
or U22023 (N_22023,N_20570,N_20592);
xor U22024 (N_22024,N_20421,N_21061);
and U22025 (N_22025,N_21215,N_21130);
nand U22026 (N_22026,N_20710,N_20627);
nor U22027 (N_22027,N_20583,N_21019);
or U22028 (N_22028,N_20379,N_20976);
and U22029 (N_22029,N_20879,N_20390);
or U22030 (N_22030,N_21056,N_20997);
or U22031 (N_22031,N_21222,N_20789);
or U22032 (N_22032,N_20003,N_20027);
or U22033 (N_22033,N_20141,N_20197);
xnor U22034 (N_22034,N_20515,N_20328);
nand U22035 (N_22035,N_20959,N_20421);
nand U22036 (N_22036,N_20853,N_20450);
xnor U22037 (N_22037,N_20096,N_20457);
nand U22038 (N_22038,N_21138,N_21094);
nor U22039 (N_22039,N_20229,N_20591);
or U22040 (N_22040,N_20636,N_20562);
or U22041 (N_22041,N_20744,N_20898);
or U22042 (N_22042,N_20283,N_21029);
or U22043 (N_22043,N_20980,N_20833);
and U22044 (N_22044,N_20502,N_20063);
nor U22045 (N_22045,N_20880,N_21102);
nand U22046 (N_22046,N_20355,N_20075);
nand U22047 (N_22047,N_21119,N_20684);
nor U22048 (N_22048,N_20429,N_20201);
nor U22049 (N_22049,N_20132,N_20319);
nor U22050 (N_22050,N_20171,N_20949);
and U22051 (N_22051,N_20789,N_20525);
or U22052 (N_22052,N_21233,N_20664);
or U22053 (N_22053,N_20481,N_20227);
and U22054 (N_22054,N_20055,N_20265);
xnor U22055 (N_22055,N_20685,N_20753);
and U22056 (N_22056,N_21235,N_20881);
nor U22057 (N_22057,N_20209,N_20778);
nand U22058 (N_22058,N_20574,N_20159);
nor U22059 (N_22059,N_20584,N_20825);
nand U22060 (N_22060,N_20001,N_20595);
and U22061 (N_22061,N_20848,N_20353);
nor U22062 (N_22062,N_20707,N_20264);
nor U22063 (N_22063,N_20815,N_20267);
nand U22064 (N_22064,N_21214,N_20209);
nor U22065 (N_22065,N_20463,N_20856);
and U22066 (N_22066,N_20307,N_20973);
xnor U22067 (N_22067,N_20896,N_20980);
and U22068 (N_22068,N_21088,N_20444);
nand U22069 (N_22069,N_21095,N_20887);
nand U22070 (N_22070,N_20102,N_20089);
xnor U22071 (N_22071,N_20352,N_20006);
or U22072 (N_22072,N_20654,N_20195);
nor U22073 (N_22073,N_21092,N_20204);
or U22074 (N_22074,N_20846,N_20146);
and U22075 (N_22075,N_20141,N_20958);
nor U22076 (N_22076,N_20833,N_20442);
or U22077 (N_22077,N_20797,N_20353);
xor U22078 (N_22078,N_21013,N_20106);
xnor U22079 (N_22079,N_20389,N_20732);
or U22080 (N_22080,N_20543,N_20513);
nand U22081 (N_22081,N_20899,N_20560);
or U22082 (N_22082,N_20748,N_20796);
xor U22083 (N_22083,N_20542,N_20029);
xnor U22084 (N_22084,N_21052,N_20131);
or U22085 (N_22085,N_21190,N_21074);
nand U22086 (N_22086,N_20509,N_21179);
or U22087 (N_22087,N_21018,N_20398);
or U22088 (N_22088,N_21247,N_21129);
and U22089 (N_22089,N_20912,N_20590);
xor U22090 (N_22090,N_20293,N_20156);
nand U22091 (N_22091,N_20352,N_21002);
xnor U22092 (N_22092,N_21156,N_20574);
and U22093 (N_22093,N_21025,N_20106);
or U22094 (N_22094,N_21193,N_21057);
and U22095 (N_22095,N_20448,N_20105);
nor U22096 (N_22096,N_20721,N_20732);
nor U22097 (N_22097,N_20750,N_20185);
xor U22098 (N_22098,N_20298,N_20548);
xnor U22099 (N_22099,N_20373,N_20621);
nand U22100 (N_22100,N_20562,N_21092);
xor U22101 (N_22101,N_21249,N_20179);
or U22102 (N_22102,N_20022,N_20630);
and U22103 (N_22103,N_20229,N_20646);
xor U22104 (N_22104,N_20863,N_20076);
nand U22105 (N_22105,N_20627,N_20275);
or U22106 (N_22106,N_21024,N_20454);
nand U22107 (N_22107,N_21128,N_20972);
xor U22108 (N_22108,N_20000,N_20962);
xor U22109 (N_22109,N_21104,N_20848);
nand U22110 (N_22110,N_20001,N_20687);
or U22111 (N_22111,N_20455,N_20169);
and U22112 (N_22112,N_20076,N_20308);
nor U22113 (N_22113,N_20624,N_20996);
or U22114 (N_22114,N_20954,N_20091);
xnor U22115 (N_22115,N_20181,N_20439);
nand U22116 (N_22116,N_20623,N_21129);
and U22117 (N_22117,N_21138,N_21130);
or U22118 (N_22118,N_20795,N_20633);
and U22119 (N_22119,N_21171,N_20816);
xnor U22120 (N_22120,N_21025,N_20872);
nand U22121 (N_22121,N_20548,N_20295);
nor U22122 (N_22122,N_21015,N_20714);
or U22123 (N_22123,N_20645,N_20921);
or U22124 (N_22124,N_20646,N_21062);
and U22125 (N_22125,N_20121,N_20835);
or U22126 (N_22126,N_21031,N_21081);
xor U22127 (N_22127,N_20423,N_20633);
nor U22128 (N_22128,N_20605,N_20924);
and U22129 (N_22129,N_20971,N_20233);
nor U22130 (N_22130,N_20309,N_20143);
and U22131 (N_22131,N_20544,N_20568);
nor U22132 (N_22132,N_21015,N_21120);
nand U22133 (N_22133,N_20761,N_21034);
nor U22134 (N_22134,N_21185,N_21186);
or U22135 (N_22135,N_21005,N_20391);
and U22136 (N_22136,N_20659,N_20958);
or U22137 (N_22137,N_21200,N_21233);
xor U22138 (N_22138,N_21125,N_20252);
nor U22139 (N_22139,N_20625,N_20739);
or U22140 (N_22140,N_20664,N_20660);
or U22141 (N_22141,N_20166,N_20121);
nand U22142 (N_22142,N_21006,N_20476);
or U22143 (N_22143,N_20242,N_20956);
nand U22144 (N_22144,N_20970,N_20171);
and U22145 (N_22145,N_20956,N_20235);
and U22146 (N_22146,N_20680,N_20149);
and U22147 (N_22147,N_20443,N_20837);
xor U22148 (N_22148,N_20953,N_20322);
nor U22149 (N_22149,N_20073,N_20731);
or U22150 (N_22150,N_21160,N_20259);
and U22151 (N_22151,N_20644,N_20691);
or U22152 (N_22152,N_20945,N_20233);
nand U22153 (N_22153,N_20571,N_20675);
nor U22154 (N_22154,N_20744,N_20596);
or U22155 (N_22155,N_20748,N_20944);
or U22156 (N_22156,N_20250,N_20593);
nand U22157 (N_22157,N_20398,N_21044);
or U22158 (N_22158,N_20351,N_20353);
nor U22159 (N_22159,N_20931,N_20386);
xnor U22160 (N_22160,N_21102,N_21067);
nor U22161 (N_22161,N_20510,N_20914);
nand U22162 (N_22162,N_20361,N_20571);
nand U22163 (N_22163,N_20319,N_20386);
nor U22164 (N_22164,N_20500,N_21207);
nand U22165 (N_22165,N_20843,N_21085);
xor U22166 (N_22166,N_20018,N_20333);
and U22167 (N_22167,N_20957,N_20627);
nand U22168 (N_22168,N_20474,N_20882);
and U22169 (N_22169,N_20305,N_20939);
or U22170 (N_22170,N_20978,N_21093);
nand U22171 (N_22171,N_20219,N_20515);
nand U22172 (N_22172,N_20338,N_20137);
or U22173 (N_22173,N_20401,N_21157);
and U22174 (N_22174,N_21120,N_20138);
and U22175 (N_22175,N_21075,N_20283);
xor U22176 (N_22176,N_21057,N_21209);
nand U22177 (N_22177,N_20891,N_20635);
and U22178 (N_22178,N_20156,N_20468);
xnor U22179 (N_22179,N_20325,N_20091);
nand U22180 (N_22180,N_20816,N_20363);
or U22181 (N_22181,N_21083,N_20773);
nor U22182 (N_22182,N_20178,N_20828);
xnor U22183 (N_22183,N_20529,N_20103);
and U22184 (N_22184,N_20144,N_20993);
nand U22185 (N_22185,N_20172,N_20902);
and U22186 (N_22186,N_20191,N_20615);
nor U22187 (N_22187,N_20063,N_21202);
nand U22188 (N_22188,N_20813,N_20028);
xor U22189 (N_22189,N_20441,N_20685);
nor U22190 (N_22190,N_20049,N_20828);
and U22191 (N_22191,N_20432,N_21099);
nand U22192 (N_22192,N_21205,N_21087);
xor U22193 (N_22193,N_20730,N_20548);
nor U22194 (N_22194,N_21139,N_20403);
xnor U22195 (N_22195,N_20449,N_20884);
nand U22196 (N_22196,N_20553,N_20172);
or U22197 (N_22197,N_20828,N_20048);
xnor U22198 (N_22198,N_20994,N_20963);
nand U22199 (N_22199,N_20159,N_20623);
or U22200 (N_22200,N_20700,N_20152);
or U22201 (N_22201,N_20950,N_20017);
nand U22202 (N_22202,N_20733,N_20601);
xor U22203 (N_22203,N_21183,N_20932);
and U22204 (N_22204,N_20910,N_21119);
nand U22205 (N_22205,N_20396,N_20211);
nand U22206 (N_22206,N_20551,N_21100);
nand U22207 (N_22207,N_20366,N_20969);
nor U22208 (N_22208,N_20044,N_20870);
nor U22209 (N_22209,N_20637,N_20618);
nand U22210 (N_22210,N_20606,N_20882);
nor U22211 (N_22211,N_20970,N_21244);
or U22212 (N_22212,N_21201,N_21071);
or U22213 (N_22213,N_20867,N_20506);
and U22214 (N_22214,N_21038,N_20032);
xnor U22215 (N_22215,N_21243,N_20489);
and U22216 (N_22216,N_20644,N_21086);
and U22217 (N_22217,N_20610,N_20516);
and U22218 (N_22218,N_21182,N_20518);
nand U22219 (N_22219,N_20372,N_20734);
or U22220 (N_22220,N_20652,N_20843);
or U22221 (N_22221,N_20227,N_20665);
and U22222 (N_22222,N_20005,N_20654);
and U22223 (N_22223,N_20449,N_20289);
and U22224 (N_22224,N_20041,N_20495);
xnor U22225 (N_22225,N_20038,N_20454);
and U22226 (N_22226,N_20986,N_20627);
nand U22227 (N_22227,N_20510,N_20527);
nand U22228 (N_22228,N_20039,N_21020);
xor U22229 (N_22229,N_20437,N_20556);
and U22230 (N_22230,N_20016,N_20475);
and U22231 (N_22231,N_20594,N_20589);
nor U22232 (N_22232,N_20507,N_20249);
nand U22233 (N_22233,N_21119,N_20444);
nor U22234 (N_22234,N_20726,N_20056);
and U22235 (N_22235,N_20440,N_20625);
xor U22236 (N_22236,N_21233,N_20928);
nor U22237 (N_22237,N_20278,N_20338);
xnor U22238 (N_22238,N_20720,N_20821);
nand U22239 (N_22239,N_20551,N_20919);
xnor U22240 (N_22240,N_21169,N_20029);
and U22241 (N_22241,N_21112,N_20169);
nand U22242 (N_22242,N_20788,N_20294);
or U22243 (N_22243,N_20038,N_20321);
xor U22244 (N_22244,N_21228,N_20620);
nor U22245 (N_22245,N_20346,N_20541);
nand U22246 (N_22246,N_20551,N_20331);
nor U22247 (N_22247,N_21135,N_20627);
or U22248 (N_22248,N_20990,N_21029);
xnor U22249 (N_22249,N_20790,N_20763);
or U22250 (N_22250,N_20555,N_21241);
and U22251 (N_22251,N_20750,N_20966);
or U22252 (N_22252,N_20152,N_20884);
xnor U22253 (N_22253,N_20228,N_20437);
and U22254 (N_22254,N_20209,N_20363);
and U22255 (N_22255,N_20183,N_20775);
nand U22256 (N_22256,N_21224,N_20736);
and U22257 (N_22257,N_20482,N_20962);
and U22258 (N_22258,N_20254,N_20433);
and U22259 (N_22259,N_20165,N_20400);
and U22260 (N_22260,N_21021,N_20881);
or U22261 (N_22261,N_20937,N_20191);
or U22262 (N_22262,N_20232,N_21100);
and U22263 (N_22263,N_20317,N_20010);
and U22264 (N_22264,N_21115,N_20718);
and U22265 (N_22265,N_20158,N_20210);
or U22266 (N_22266,N_20128,N_20429);
and U22267 (N_22267,N_20774,N_20328);
xor U22268 (N_22268,N_20604,N_20921);
and U22269 (N_22269,N_21108,N_20010);
nand U22270 (N_22270,N_21208,N_20125);
nand U22271 (N_22271,N_20691,N_20028);
xor U22272 (N_22272,N_21055,N_20598);
or U22273 (N_22273,N_20484,N_20925);
or U22274 (N_22274,N_20981,N_20293);
and U22275 (N_22275,N_21099,N_20916);
nand U22276 (N_22276,N_20150,N_21113);
and U22277 (N_22277,N_21236,N_20285);
xor U22278 (N_22278,N_21113,N_20011);
nor U22279 (N_22279,N_20598,N_20579);
nor U22280 (N_22280,N_20662,N_20171);
and U22281 (N_22281,N_20457,N_20123);
nand U22282 (N_22282,N_21050,N_20442);
or U22283 (N_22283,N_20619,N_20937);
nand U22284 (N_22284,N_20836,N_20889);
and U22285 (N_22285,N_20348,N_21195);
and U22286 (N_22286,N_20765,N_20138);
xnor U22287 (N_22287,N_20732,N_20568);
nand U22288 (N_22288,N_21156,N_21225);
xor U22289 (N_22289,N_20722,N_21222);
xnor U22290 (N_22290,N_20979,N_21174);
nand U22291 (N_22291,N_20636,N_20850);
nand U22292 (N_22292,N_20948,N_20045);
xnor U22293 (N_22293,N_20922,N_20454);
xnor U22294 (N_22294,N_20741,N_20453);
or U22295 (N_22295,N_20375,N_20059);
nand U22296 (N_22296,N_20061,N_20707);
or U22297 (N_22297,N_20753,N_20843);
nor U22298 (N_22298,N_20270,N_20789);
or U22299 (N_22299,N_21179,N_20683);
and U22300 (N_22300,N_20247,N_21054);
nand U22301 (N_22301,N_20170,N_20965);
xnor U22302 (N_22302,N_20623,N_21082);
or U22303 (N_22303,N_21129,N_20711);
or U22304 (N_22304,N_20789,N_20111);
nor U22305 (N_22305,N_20317,N_20659);
nor U22306 (N_22306,N_20651,N_20540);
xnor U22307 (N_22307,N_21043,N_20854);
and U22308 (N_22308,N_20522,N_20593);
and U22309 (N_22309,N_20327,N_20009);
or U22310 (N_22310,N_20761,N_20687);
nand U22311 (N_22311,N_20197,N_20232);
and U22312 (N_22312,N_20371,N_21051);
nor U22313 (N_22313,N_20546,N_20202);
and U22314 (N_22314,N_20165,N_20761);
xnor U22315 (N_22315,N_20922,N_20014);
nor U22316 (N_22316,N_20770,N_20778);
nand U22317 (N_22317,N_21037,N_20438);
nand U22318 (N_22318,N_20371,N_20921);
nand U22319 (N_22319,N_20711,N_20800);
nand U22320 (N_22320,N_21140,N_20454);
and U22321 (N_22321,N_20171,N_20123);
nand U22322 (N_22322,N_20542,N_21158);
or U22323 (N_22323,N_20317,N_21153);
nand U22324 (N_22324,N_21033,N_20170);
xor U22325 (N_22325,N_20970,N_20216);
nor U22326 (N_22326,N_20255,N_20730);
xor U22327 (N_22327,N_20828,N_20840);
xnor U22328 (N_22328,N_20333,N_20807);
nor U22329 (N_22329,N_20169,N_20079);
nand U22330 (N_22330,N_21107,N_20183);
xnor U22331 (N_22331,N_20538,N_21234);
xor U22332 (N_22332,N_20440,N_20706);
xor U22333 (N_22333,N_20743,N_20994);
nor U22334 (N_22334,N_20871,N_20345);
or U22335 (N_22335,N_20634,N_20712);
and U22336 (N_22336,N_20796,N_20179);
and U22337 (N_22337,N_20258,N_20922);
xnor U22338 (N_22338,N_20823,N_21126);
or U22339 (N_22339,N_20355,N_21036);
and U22340 (N_22340,N_20458,N_20746);
nor U22341 (N_22341,N_21052,N_20885);
nor U22342 (N_22342,N_20694,N_20035);
xor U22343 (N_22343,N_20400,N_21044);
nor U22344 (N_22344,N_20679,N_20716);
nor U22345 (N_22345,N_20976,N_21090);
nor U22346 (N_22346,N_20216,N_20327);
and U22347 (N_22347,N_21093,N_20434);
xnor U22348 (N_22348,N_20213,N_20192);
nor U22349 (N_22349,N_20025,N_20442);
nand U22350 (N_22350,N_21034,N_20952);
nand U22351 (N_22351,N_20756,N_21027);
or U22352 (N_22352,N_21025,N_20212);
and U22353 (N_22353,N_20211,N_20023);
and U22354 (N_22354,N_21004,N_20636);
and U22355 (N_22355,N_20997,N_20552);
nor U22356 (N_22356,N_20274,N_21000);
xor U22357 (N_22357,N_20425,N_20655);
or U22358 (N_22358,N_21028,N_20508);
xor U22359 (N_22359,N_20007,N_20635);
or U22360 (N_22360,N_20306,N_20790);
xnor U22361 (N_22361,N_21133,N_20217);
nor U22362 (N_22362,N_20217,N_21143);
or U22363 (N_22363,N_20526,N_20033);
and U22364 (N_22364,N_20503,N_20537);
xnor U22365 (N_22365,N_20309,N_20513);
and U22366 (N_22366,N_21043,N_21168);
xnor U22367 (N_22367,N_20451,N_20043);
nor U22368 (N_22368,N_20992,N_20946);
or U22369 (N_22369,N_21163,N_20948);
nor U22370 (N_22370,N_20702,N_20558);
nand U22371 (N_22371,N_20695,N_20956);
xnor U22372 (N_22372,N_20050,N_20477);
xnor U22373 (N_22373,N_21035,N_21149);
and U22374 (N_22374,N_20490,N_20119);
and U22375 (N_22375,N_20148,N_20888);
and U22376 (N_22376,N_21230,N_20091);
or U22377 (N_22377,N_20381,N_20667);
nor U22378 (N_22378,N_20397,N_20534);
or U22379 (N_22379,N_20373,N_21158);
or U22380 (N_22380,N_21239,N_21117);
or U22381 (N_22381,N_20135,N_20341);
xnor U22382 (N_22382,N_20504,N_21007);
and U22383 (N_22383,N_20800,N_20902);
xnor U22384 (N_22384,N_20123,N_20668);
nand U22385 (N_22385,N_21019,N_20671);
nor U22386 (N_22386,N_21059,N_20109);
or U22387 (N_22387,N_20358,N_21053);
nand U22388 (N_22388,N_20891,N_20574);
and U22389 (N_22389,N_20703,N_20464);
xor U22390 (N_22390,N_20255,N_20697);
and U22391 (N_22391,N_21098,N_20047);
nor U22392 (N_22392,N_20991,N_20015);
xor U22393 (N_22393,N_20565,N_20682);
or U22394 (N_22394,N_20040,N_21155);
xor U22395 (N_22395,N_20321,N_20147);
and U22396 (N_22396,N_20907,N_20093);
and U22397 (N_22397,N_20603,N_20588);
or U22398 (N_22398,N_20878,N_20843);
nand U22399 (N_22399,N_20215,N_20236);
nand U22400 (N_22400,N_21022,N_20840);
or U22401 (N_22401,N_20956,N_20327);
nor U22402 (N_22402,N_20682,N_21027);
xnor U22403 (N_22403,N_20856,N_20943);
xor U22404 (N_22404,N_20090,N_20412);
or U22405 (N_22405,N_20743,N_20133);
nand U22406 (N_22406,N_21031,N_20831);
and U22407 (N_22407,N_20806,N_20723);
and U22408 (N_22408,N_21039,N_20366);
or U22409 (N_22409,N_20540,N_21050);
and U22410 (N_22410,N_20643,N_20150);
nor U22411 (N_22411,N_20980,N_21201);
nor U22412 (N_22412,N_20221,N_20474);
and U22413 (N_22413,N_21210,N_20267);
nand U22414 (N_22414,N_20112,N_21215);
nor U22415 (N_22415,N_20109,N_20122);
or U22416 (N_22416,N_20423,N_21078);
or U22417 (N_22417,N_21121,N_20771);
nand U22418 (N_22418,N_20720,N_20124);
or U22419 (N_22419,N_21093,N_20911);
xor U22420 (N_22420,N_20279,N_21249);
nor U22421 (N_22421,N_20185,N_20463);
or U22422 (N_22422,N_20163,N_20339);
and U22423 (N_22423,N_20168,N_20030);
xnor U22424 (N_22424,N_20098,N_20067);
nand U22425 (N_22425,N_20421,N_21035);
nand U22426 (N_22426,N_20188,N_20489);
nor U22427 (N_22427,N_20191,N_20230);
or U22428 (N_22428,N_20775,N_21146);
or U22429 (N_22429,N_20757,N_20158);
xnor U22430 (N_22430,N_20205,N_20067);
or U22431 (N_22431,N_20569,N_20896);
xor U22432 (N_22432,N_20958,N_20363);
nand U22433 (N_22433,N_20121,N_20541);
and U22434 (N_22434,N_20492,N_20138);
or U22435 (N_22435,N_20593,N_20702);
nor U22436 (N_22436,N_20558,N_20495);
nand U22437 (N_22437,N_20454,N_21133);
or U22438 (N_22438,N_20694,N_20240);
xor U22439 (N_22439,N_20063,N_20969);
nor U22440 (N_22440,N_20371,N_20635);
nand U22441 (N_22441,N_20829,N_20215);
nor U22442 (N_22442,N_20236,N_20013);
xor U22443 (N_22443,N_20658,N_20599);
nor U22444 (N_22444,N_20372,N_20985);
xor U22445 (N_22445,N_20205,N_20536);
and U22446 (N_22446,N_20537,N_21153);
nor U22447 (N_22447,N_20189,N_21032);
nor U22448 (N_22448,N_20230,N_20831);
nor U22449 (N_22449,N_20516,N_20498);
and U22450 (N_22450,N_20344,N_20011);
nand U22451 (N_22451,N_20911,N_20027);
and U22452 (N_22452,N_20465,N_20709);
nor U22453 (N_22453,N_20743,N_20965);
and U22454 (N_22454,N_20811,N_20962);
xor U22455 (N_22455,N_20968,N_21043);
nand U22456 (N_22456,N_20157,N_20126);
and U22457 (N_22457,N_20459,N_21019);
nand U22458 (N_22458,N_20875,N_21185);
nor U22459 (N_22459,N_21007,N_20526);
nor U22460 (N_22460,N_20912,N_20763);
and U22461 (N_22461,N_21091,N_20744);
and U22462 (N_22462,N_20865,N_21082);
xor U22463 (N_22463,N_20241,N_20453);
and U22464 (N_22464,N_20052,N_20518);
and U22465 (N_22465,N_21208,N_20900);
and U22466 (N_22466,N_20352,N_20144);
and U22467 (N_22467,N_20825,N_20341);
nand U22468 (N_22468,N_20416,N_20904);
or U22469 (N_22469,N_20920,N_20933);
or U22470 (N_22470,N_20593,N_20416);
and U22471 (N_22471,N_20751,N_20112);
and U22472 (N_22472,N_20441,N_21034);
nor U22473 (N_22473,N_20552,N_20459);
xnor U22474 (N_22474,N_20137,N_21053);
or U22475 (N_22475,N_21049,N_20316);
or U22476 (N_22476,N_20094,N_20000);
xor U22477 (N_22477,N_21235,N_20742);
and U22478 (N_22478,N_20460,N_20050);
xor U22479 (N_22479,N_21024,N_20197);
and U22480 (N_22480,N_20195,N_20604);
xnor U22481 (N_22481,N_20338,N_20688);
xor U22482 (N_22482,N_20854,N_20012);
and U22483 (N_22483,N_20078,N_20921);
and U22484 (N_22484,N_21007,N_20835);
nand U22485 (N_22485,N_20608,N_20793);
and U22486 (N_22486,N_20520,N_20548);
and U22487 (N_22487,N_20116,N_21119);
or U22488 (N_22488,N_20834,N_21181);
nand U22489 (N_22489,N_20108,N_20678);
nand U22490 (N_22490,N_20407,N_20125);
xnor U22491 (N_22491,N_21237,N_20028);
nor U22492 (N_22492,N_21028,N_20156);
nand U22493 (N_22493,N_20403,N_20890);
and U22494 (N_22494,N_20159,N_20559);
nor U22495 (N_22495,N_20609,N_20023);
xor U22496 (N_22496,N_21114,N_20634);
nand U22497 (N_22497,N_20253,N_21216);
nand U22498 (N_22498,N_20033,N_20078);
nand U22499 (N_22499,N_20196,N_20484);
and U22500 (N_22500,N_21801,N_21583);
or U22501 (N_22501,N_21279,N_22210);
nor U22502 (N_22502,N_21383,N_21266);
and U22503 (N_22503,N_22304,N_21844);
nor U22504 (N_22504,N_22228,N_21866);
nand U22505 (N_22505,N_21586,N_21918);
and U22506 (N_22506,N_21566,N_21865);
and U22507 (N_22507,N_22201,N_22482);
nor U22508 (N_22508,N_21517,N_22025);
nor U22509 (N_22509,N_22348,N_21397);
nor U22510 (N_22510,N_21968,N_21936);
nand U22511 (N_22511,N_21490,N_21278);
nor U22512 (N_22512,N_21701,N_21996);
and U22513 (N_22513,N_21914,N_21412);
or U22514 (N_22514,N_21427,N_21598);
and U22515 (N_22515,N_21420,N_22462);
or U22516 (N_22516,N_21474,N_22254);
nand U22517 (N_22517,N_21469,N_21609);
and U22518 (N_22518,N_21476,N_22143);
nor U22519 (N_22519,N_21599,N_22172);
and U22520 (N_22520,N_21819,N_22111);
and U22521 (N_22521,N_21899,N_21753);
xor U22522 (N_22522,N_22182,N_22427);
or U22523 (N_22523,N_22132,N_21313);
and U22524 (N_22524,N_21995,N_21700);
or U22525 (N_22525,N_21465,N_22493);
and U22526 (N_22526,N_21937,N_22035);
xnor U22527 (N_22527,N_22485,N_21990);
nand U22528 (N_22528,N_22224,N_22423);
or U22529 (N_22529,N_21394,N_21509);
nor U22530 (N_22530,N_21822,N_21354);
nor U22531 (N_22531,N_21662,N_21897);
or U22532 (N_22532,N_22108,N_22439);
xnor U22533 (N_22533,N_21518,N_21468);
or U22534 (N_22534,N_21893,N_22457);
and U22535 (N_22535,N_22019,N_21967);
and U22536 (N_22536,N_21386,N_21972);
and U22537 (N_22537,N_22225,N_21624);
nor U22538 (N_22538,N_21280,N_21614);
nor U22539 (N_22539,N_21842,N_21933);
or U22540 (N_22540,N_22494,N_21776);
and U22541 (N_22541,N_22222,N_21352);
nor U22542 (N_22542,N_22384,N_21876);
and U22543 (N_22543,N_22118,N_22286);
and U22544 (N_22544,N_22281,N_21551);
and U22545 (N_22545,N_22474,N_22327);
nand U22546 (N_22546,N_21548,N_22296);
nand U22547 (N_22547,N_21959,N_21514);
or U22548 (N_22548,N_22029,N_22006);
nor U22549 (N_22549,N_22455,N_22047);
xnor U22550 (N_22550,N_21447,N_22101);
or U22551 (N_22551,N_21319,N_21962);
and U22552 (N_22552,N_22215,N_21411);
xor U22553 (N_22553,N_21724,N_22151);
or U22554 (N_22554,N_21450,N_22186);
nor U22555 (N_22555,N_22200,N_22026);
xor U22556 (N_22556,N_22305,N_21326);
xor U22557 (N_22557,N_21963,N_22115);
nand U22558 (N_22558,N_22272,N_21917);
or U22559 (N_22559,N_22220,N_21414);
or U22560 (N_22560,N_21732,N_21454);
nand U22561 (N_22561,N_21846,N_21760);
xnor U22562 (N_22562,N_21888,N_22290);
xnor U22563 (N_22563,N_21303,N_21610);
nor U22564 (N_22564,N_22445,N_22013);
nand U22565 (N_22565,N_22161,N_22011);
xor U22566 (N_22566,N_21814,N_22422);
and U22567 (N_22567,N_21339,N_22017);
or U22568 (N_22568,N_22377,N_22027);
nand U22569 (N_22569,N_21558,N_21683);
nand U22570 (N_22570,N_21520,N_22269);
and U22571 (N_22571,N_22004,N_21422);
xnor U22572 (N_22572,N_21634,N_21878);
or U22573 (N_22573,N_21541,N_22072);
or U22574 (N_22574,N_21991,N_22406);
and U22575 (N_22575,N_21674,N_21883);
and U22576 (N_22576,N_21739,N_21401);
nor U22577 (N_22577,N_22226,N_22120);
or U22578 (N_22578,N_22358,N_21672);
and U22579 (N_22579,N_22033,N_21938);
nand U22580 (N_22580,N_22233,N_21591);
xor U22581 (N_22581,N_21980,N_21628);
xnor U22582 (N_22582,N_21418,N_22175);
nand U22583 (N_22583,N_21443,N_21781);
nand U22584 (N_22584,N_21742,N_21253);
and U22585 (N_22585,N_21799,N_21324);
or U22586 (N_22586,N_22402,N_21976);
or U22587 (N_22587,N_22399,N_22478);
or U22588 (N_22588,N_21793,N_21941);
xnor U22589 (N_22589,N_22472,N_21851);
or U22590 (N_22590,N_22070,N_21746);
and U22591 (N_22591,N_21578,N_22274);
nand U22592 (N_22592,N_21853,N_22360);
nor U22593 (N_22593,N_21925,N_21633);
or U22594 (N_22594,N_21540,N_21791);
nand U22595 (N_22595,N_21960,N_21794);
or U22596 (N_22596,N_22163,N_22202);
and U22597 (N_22597,N_21834,N_21954);
xor U22598 (N_22598,N_22337,N_21913);
xor U22599 (N_22599,N_21749,N_21657);
and U22600 (N_22600,N_21951,N_22090);
and U22601 (N_22601,N_22287,N_21434);
and U22602 (N_22602,N_21758,N_21796);
nand U22603 (N_22603,N_21765,N_21511);
nor U22604 (N_22604,N_22336,N_21727);
nor U22605 (N_22605,N_21625,N_21478);
xor U22606 (N_22606,N_22002,N_21573);
and U22607 (N_22607,N_21986,N_21903);
nor U22608 (N_22608,N_22446,N_21259);
or U22609 (N_22609,N_22203,N_21812);
nor U22610 (N_22610,N_21989,N_21644);
or U22611 (N_22611,N_21515,N_22429);
nor U22612 (N_22612,N_22345,N_21309);
nor U22613 (N_22613,N_21716,N_22189);
nand U22614 (N_22614,N_22039,N_21790);
xnor U22615 (N_22615,N_21704,N_21652);
xor U22616 (N_22616,N_21463,N_22448);
nor U22617 (N_22617,N_22040,N_21286);
or U22618 (N_22618,N_21364,N_21587);
and U22619 (N_22619,N_22407,N_21432);
xor U22620 (N_22620,N_21366,N_22204);
and U22621 (N_22621,N_22372,N_21815);
nor U22622 (N_22622,N_21305,N_21696);
and U22623 (N_22623,N_22251,N_22467);
nand U22624 (N_22624,N_22037,N_21983);
or U22625 (N_22625,N_21916,N_22431);
xor U22626 (N_22626,N_21671,N_21600);
xor U22627 (N_22627,N_22420,N_21969);
and U22628 (N_22628,N_21332,N_21906);
and U22629 (N_22629,N_21529,N_22425);
or U22630 (N_22630,N_22408,N_21594);
xor U22631 (N_22631,N_21330,N_22321);
and U22632 (N_22632,N_21627,N_21729);
and U22633 (N_22633,N_22401,N_21905);
nand U22634 (N_22634,N_21543,N_21966);
and U22635 (N_22635,N_22009,N_21948);
nor U22636 (N_22636,N_21268,N_21698);
nor U22637 (N_22637,N_21409,N_22165);
or U22638 (N_22638,N_21784,N_21390);
and U22639 (N_22639,N_21283,N_21863);
nor U22640 (N_22640,N_22329,N_21340);
xor U22641 (N_22641,N_21538,N_22044);
nand U22642 (N_22642,N_22173,N_22032);
or U22643 (N_22643,N_21975,N_21690);
nor U22644 (N_22644,N_21838,N_22308);
nor U22645 (N_22645,N_21449,N_21856);
and U22646 (N_22646,N_22307,N_22428);
and U22647 (N_22647,N_21568,N_22332);
nand U22648 (N_22648,N_22323,N_21754);
or U22649 (N_22649,N_21717,N_21590);
nor U22650 (N_22650,N_22417,N_21785);
and U22651 (N_22651,N_22415,N_21445);
and U22652 (N_22652,N_21579,N_21389);
and U22653 (N_22653,N_21441,N_21398);
nor U22654 (N_22654,N_21743,N_21949);
nand U22655 (N_22655,N_21329,N_21284);
and U22656 (N_22656,N_21800,N_21741);
nand U22657 (N_22657,N_22125,N_21787);
or U22658 (N_22658,N_21519,N_21378);
and U22659 (N_22659,N_22020,N_21521);
nor U22660 (N_22660,N_21502,N_22082);
xnor U22661 (N_22661,N_21604,N_21929);
nand U22662 (N_22662,N_22442,N_21821);
or U22663 (N_22663,N_21258,N_22043);
xor U22664 (N_22664,N_21885,N_21769);
nor U22665 (N_22665,N_22418,N_21531);
and U22666 (N_22666,N_21553,N_21461);
nor U22667 (N_22667,N_21556,N_22054);
or U22668 (N_22668,N_22324,N_21699);
xor U22669 (N_22669,N_21486,N_21348);
or U22670 (N_22670,N_22400,N_22346);
nor U22671 (N_22671,N_22350,N_22405);
and U22672 (N_22672,N_21525,N_21823);
xnor U22673 (N_22673,N_22190,N_22005);
xor U22674 (N_22674,N_22370,N_22241);
xnor U22675 (N_22675,N_21431,N_22266);
nor U22676 (N_22676,N_22158,N_22052);
nor U22677 (N_22677,N_22320,N_21417);
xor U22678 (N_22678,N_22261,N_22007);
or U22679 (N_22679,N_21372,N_21275);
or U22680 (N_22680,N_21909,N_22456);
and U22681 (N_22681,N_21680,N_21872);
xnor U22682 (N_22682,N_21676,N_21289);
nor U22683 (N_22683,N_21798,N_21988);
and U22684 (N_22684,N_21410,N_22131);
nand U22685 (N_22685,N_22084,N_22010);
or U22686 (N_22686,N_21934,N_22343);
or U22687 (N_22687,N_21589,N_22475);
or U22688 (N_22688,N_21595,N_22335);
and U22689 (N_22689,N_21462,N_21645);
nor U22690 (N_22690,N_21255,N_21351);
xnor U22691 (N_22691,N_21890,N_22303);
nand U22692 (N_22692,N_22310,N_21408);
xnor U22693 (N_22693,N_21764,N_21251);
or U22694 (N_22694,N_22312,N_22382);
or U22695 (N_22695,N_22127,N_22065);
xor U22696 (N_22696,N_22022,N_21320);
xnor U22697 (N_22697,N_21261,N_21726);
xor U22698 (N_22698,N_21868,N_22443);
or U22699 (N_22699,N_21361,N_21947);
xor U22700 (N_22700,N_22096,N_22205);
nand U22701 (N_22701,N_22124,N_22162);
xor U22702 (N_22702,N_21612,N_21564);
xor U22703 (N_22703,N_21272,N_22036);
nor U22704 (N_22704,N_22444,N_22438);
nand U22705 (N_22705,N_21267,N_22489);
nand U22706 (N_22706,N_21257,N_22480);
nand U22707 (N_22707,N_21779,N_21508);
and U22708 (N_22708,N_21880,N_21659);
and U22709 (N_22709,N_21342,N_21608);
xnor U22710 (N_22710,N_21360,N_21935);
nand U22711 (N_22711,N_22318,N_21611);
and U22712 (N_22712,N_22486,N_21596);
nor U22713 (N_22713,N_21423,N_21281);
xnor U22714 (N_22714,N_21945,N_21537);
nand U22715 (N_22715,N_21260,N_21648);
and U22716 (N_22716,N_21854,N_21384);
or U22717 (N_22717,N_22471,N_21887);
xor U22718 (N_22718,N_22255,N_21536);
nor U22719 (N_22719,N_22347,N_22057);
and U22720 (N_22720,N_21734,N_21295);
nor U22721 (N_22721,N_21273,N_21831);
or U22722 (N_22722,N_21315,N_22387);
or U22723 (N_22723,N_21370,N_21557);
nand U22724 (N_22724,N_21481,N_21436);
or U22725 (N_22725,N_21451,N_22366);
nor U22726 (N_22726,N_21448,N_21617);
nor U22727 (N_22727,N_21839,N_21381);
nor U22728 (N_22728,N_21359,N_21982);
or U22729 (N_22729,N_21747,N_22106);
and U22730 (N_22730,N_21421,N_21848);
nor U22731 (N_22731,N_22453,N_21722);
or U22732 (N_22732,N_22338,N_21483);
and U22733 (N_22733,N_21382,N_22081);
nand U22734 (N_22734,N_22000,N_21879);
xor U22735 (N_22735,N_21923,N_22207);
and U22736 (N_22736,N_21884,N_21736);
xor U22737 (N_22737,N_22061,N_22459);
xor U22738 (N_22738,N_22099,N_22153);
xor U22739 (N_22739,N_22376,N_21631);
or U22740 (N_22740,N_21419,N_21569);
or U22741 (N_22741,N_22130,N_22160);
or U22742 (N_22742,N_21882,N_21789);
nor U22743 (N_22743,N_21555,N_22353);
and U22744 (N_22744,N_21416,N_22264);
nor U22745 (N_22745,N_22028,N_21953);
and U22746 (N_22746,N_21928,N_21770);
or U22747 (N_22747,N_22188,N_21867);
nor U22748 (N_22748,N_21697,N_21932);
nand U22749 (N_22749,N_22156,N_21321);
nand U22750 (N_22750,N_21994,N_21271);
and U22751 (N_22751,N_22123,N_21997);
nand U22752 (N_22752,N_22253,N_22314);
and U22753 (N_22753,N_21919,N_21585);
nor U22754 (N_22754,N_22379,N_21830);
xnor U22755 (N_22755,N_21908,N_22293);
xnor U22756 (N_22756,N_22497,N_22479);
nor U22757 (N_22757,N_21797,N_21495);
and U22758 (N_22758,N_21792,N_21488);
nor U22759 (N_22759,N_21775,N_22426);
and U22760 (N_22760,N_21325,N_21973);
nand U22761 (N_22761,N_21355,N_21300);
and U22762 (N_22762,N_22359,N_22289);
nand U22763 (N_22763,N_21547,N_22239);
and U22764 (N_22764,N_21402,N_21889);
nand U22765 (N_22765,N_22212,N_22381);
nor U22766 (N_22766,N_22144,N_22045);
nand U22767 (N_22767,N_22258,N_21357);
and U22768 (N_22768,N_21626,N_21593);
or U22769 (N_22769,N_21510,N_22034);
or U22770 (N_22770,N_21745,N_21827);
nand U22771 (N_22771,N_21719,N_21387);
and U22772 (N_22772,N_21522,N_21670);
or U22773 (N_22773,N_22041,N_21686);
nand U22774 (N_22774,N_21424,N_21689);
or U22775 (N_22775,N_21497,N_22016);
xnor U22776 (N_22776,N_21274,N_22317);
nor U22777 (N_22777,N_21570,N_21350);
nor U22778 (N_22778,N_21504,N_21847);
xor U22779 (N_22779,N_22285,N_21773);
or U22780 (N_22780,N_22473,N_21597);
or U22781 (N_22781,N_22491,N_22363);
or U22782 (N_22782,N_21377,N_21438);
and U22783 (N_22783,N_21649,N_21344);
or U22784 (N_22784,N_21860,N_21376);
xnor U22785 (N_22785,N_21407,N_22257);
or U22786 (N_22786,N_21493,N_22280);
nor U22787 (N_22787,N_22227,N_21318);
xnor U22788 (N_22788,N_21310,N_22492);
and U22789 (N_22789,N_21458,N_21588);
and U22790 (N_22790,N_21992,N_22167);
nand U22791 (N_22791,N_21946,N_21693);
and U22792 (N_22792,N_22394,N_21312);
nand U22793 (N_22793,N_21506,N_21491);
xor U22794 (N_22794,N_21858,N_21406);
or U22795 (N_22795,N_21345,N_21824);
or U22796 (N_22796,N_21459,N_21825);
or U22797 (N_22797,N_21282,N_21641);
nand U22798 (N_22798,N_22416,N_22369);
nand U22799 (N_22799,N_22012,N_21895);
nand U22800 (N_22800,N_21560,N_21503);
nor U22801 (N_22801,N_21681,N_21804);
and U22802 (N_22802,N_22196,N_22171);
nand U22803 (N_22803,N_22062,N_22383);
xnor U22804 (N_22804,N_21400,N_21496);
nor U22805 (N_22805,N_21592,N_22184);
nor U22806 (N_22806,N_21924,N_21613);
nor U22807 (N_22807,N_21964,N_21554);
nor U22808 (N_22808,N_21263,N_21550);
and U22809 (N_22809,N_21635,N_21262);
nor U22810 (N_22810,N_22100,N_22334);
and U22811 (N_22811,N_22078,N_22192);
or U22812 (N_22812,N_22242,N_21256);
or U22813 (N_22813,N_22015,N_21703);
or U22814 (N_22814,N_21678,N_22488);
or U22815 (N_22815,N_22050,N_21971);
xnor U22816 (N_22816,N_21661,N_21668);
and U22817 (N_22817,N_22234,N_21806);
nor U22818 (N_22818,N_21655,N_21766);
nor U22819 (N_22819,N_22481,N_21285);
or U22820 (N_22820,N_22447,N_22465);
xor U22821 (N_22821,N_22271,N_21264);
or U22822 (N_22822,N_21841,N_21930);
and U22823 (N_22823,N_22169,N_21892);
nor U22824 (N_22824,N_22409,N_22107);
nor U22825 (N_22825,N_21299,N_21979);
nand U22826 (N_22826,N_21582,N_21388);
xnor U22827 (N_22827,N_21473,N_22299);
and U22828 (N_22828,N_21396,N_22424);
nand U22829 (N_22829,N_22077,N_22146);
nor U22830 (N_22830,N_21639,N_21833);
and U22831 (N_22831,N_22326,N_21545);
nor U22832 (N_22832,N_22176,N_22378);
nor U22833 (N_22833,N_21565,N_22080);
xnor U22834 (N_22834,N_22325,N_21926);
xnor U22835 (N_22835,N_21437,N_21759);
xor U22836 (N_22836,N_21978,N_22351);
nand U22837 (N_22837,N_22391,N_22380);
and U22838 (N_22838,N_21720,N_21981);
nor U22839 (N_22839,N_21638,N_22086);
xor U22840 (N_22840,N_22244,N_22421);
or U22841 (N_22841,N_21290,N_21780);
nand U22842 (N_22842,N_21673,N_22278);
and U22843 (N_22843,N_21763,N_22235);
nor U22844 (N_22844,N_21415,N_21998);
and U22845 (N_22845,N_21685,N_21642);
xor U22846 (N_22846,N_22279,N_22075);
and U22847 (N_22847,N_22354,N_22059);
xnor U22848 (N_22848,N_21873,N_22436);
nor U22849 (N_22849,N_22149,N_21316);
nand U22850 (N_22850,N_21306,N_22470);
and U22851 (N_22851,N_22483,N_21651);
and U22852 (N_22852,N_21296,N_21666);
nand U22853 (N_22853,N_22216,N_21314);
or U22854 (N_22854,N_22198,N_21921);
nor U22855 (N_22855,N_21363,N_22051);
and U22856 (N_22856,N_21786,N_21311);
or U22857 (N_22857,N_21563,N_22435);
nand U22858 (N_22858,N_22259,N_21901);
xor U22859 (N_22859,N_21512,N_21492);
xor U22860 (N_22860,N_22294,N_21692);
nand U22861 (N_22861,N_21489,N_21532);
xor U22862 (N_22862,N_21869,N_21485);
and U22863 (N_22863,N_21664,N_22135);
and U22864 (N_22864,N_21805,N_21466);
xor U22865 (N_22865,N_21694,N_21970);
nand U22866 (N_22866,N_22454,N_21961);
nor U22867 (N_22867,N_21871,N_21737);
or U22868 (N_22868,N_21446,N_21721);
xnor U22869 (N_22869,N_21898,N_22484);
and U22870 (N_22870,N_22058,N_22433);
xnor U22871 (N_22871,N_21751,N_21323);
or U22872 (N_22872,N_21710,N_22451);
nor U22873 (N_22873,N_22340,N_21528);
nor U22874 (N_22874,N_22122,N_22066);
nand U22875 (N_22875,N_21439,N_21931);
or U22876 (N_22876,N_21516,N_22396);
and U22877 (N_22877,N_21304,N_22373);
or U22878 (N_22878,N_22141,N_21471);
nor U22879 (N_22879,N_22440,N_22148);
nand U22880 (N_22880,N_22432,N_22461);
nand U22881 (N_22881,N_21457,N_22275);
nor U22882 (N_22882,N_22008,N_21752);
and U22883 (N_22883,N_22083,N_22460);
nor U22884 (N_22884,N_21276,N_22450);
nor U22885 (N_22885,N_21499,N_22055);
or U22886 (N_22886,N_21857,N_21336);
nand U22887 (N_22887,N_21373,N_21475);
nor U22888 (N_22888,N_21429,N_21920);
xnor U22889 (N_22889,N_21803,N_22468);
or U22890 (N_22890,N_21544,N_22330);
or U22891 (N_22891,N_22398,N_21993);
nand U22892 (N_22892,N_21298,N_21709);
or U22893 (N_22893,N_22046,N_22194);
nor U22894 (N_22894,N_22223,N_21813);
xor U22895 (N_22895,N_21603,N_21413);
and U22896 (N_22896,N_21718,N_21480);
xor U22897 (N_22897,N_21912,N_22395);
xnor U22898 (N_22898,N_21356,N_21728);
xor U22899 (N_22899,N_21404,N_22300);
nand U22900 (N_22900,N_22282,N_21392);
xor U22901 (N_22901,N_21894,N_22221);
and U22902 (N_22902,N_22024,N_22397);
nand U22903 (N_22903,N_21395,N_22076);
nand U22904 (N_22904,N_21712,N_21622);
xor U22905 (N_22905,N_21607,N_22134);
xnor U22906 (N_22906,N_22362,N_21533);
and U22907 (N_22907,N_21380,N_21393);
nor U22908 (N_22908,N_22085,N_22230);
xor U22909 (N_22909,N_21574,N_21322);
xnor U22910 (N_22910,N_21498,N_21654);
or U22911 (N_22911,N_21761,N_21774);
and U22912 (N_22912,N_22097,N_21886);
nand U22913 (N_22913,N_22413,N_22208);
nor U22914 (N_22914,N_21524,N_21647);
nand U22915 (N_22915,N_21818,N_22157);
nor U22916 (N_22916,N_22177,N_21270);
or U22917 (N_22917,N_21552,N_21840);
nand U22918 (N_22918,N_21957,N_21811);
nand U22919 (N_22919,N_22056,N_22098);
nand U22920 (N_22920,N_21881,N_22419);
nor U22921 (N_22921,N_22183,N_22137);
nand U22922 (N_22922,N_22231,N_21505);
nor U22923 (N_22923,N_22277,N_22364);
nand U22924 (N_22924,N_22357,N_21367);
or U22925 (N_22925,N_21369,N_21810);
or U22926 (N_22926,N_21714,N_22352);
and U22927 (N_22927,N_21845,N_21985);
nand U22928 (N_22928,N_21379,N_21559);
nor U22929 (N_22929,N_21850,N_22498);
xor U22930 (N_22930,N_21861,N_21927);
or U22931 (N_22931,N_22119,N_22138);
or U22932 (N_22932,N_22038,N_22499);
nand U22933 (N_22933,N_22064,N_21755);
nand U22934 (N_22934,N_22191,N_21669);
and U22935 (N_22935,N_22328,N_22238);
xor U22936 (N_22936,N_22114,N_21293);
nand U22937 (N_22937,N_21679,N_21606);
nor U22938 (N_22938,N_21942,N_21535);
and U22939 (N_22939,N_22218,N_22030);
xnor U22940 (N_22940,N_22365,N_22349);
nor U22941 (N_22941,N_21277,N_21494);
xnor U22942 (N_22942,N_21731,N_21965);
xor U22943 (N_22943,N_21795,N_21615);
and U22944 (N_22944,N_22302,N_21534);
nor U22945 (N_22945,N_22063,N_21621);
or U22946 (N_22946,N_21526,N_21605);
nor U22947 (N_22947,N_21630,N_21308);
nor U22948 (N_22948,N_21723,N_21460);
nand U22949 (N_22949,N_21337,N_22333);
nand U22950 (N_22950,N_21733,N_21952);
and U22951 (N_22951,N_22168,N_21768);
nand U22952 (N_22952,N_22344,N_21750);
and U22953 (N_22953,N_22109,N_22089);
xnor U22954 (N_22954,N_21353,N_21837);
nor U22955 (N_22955,N_21771,N_22095);
and U22956 (N_22956,N_21744,N_21287);
nor U22957 (N_22957,N_21829,N_21391);
xnor U22958 (N_22958,N_21832,N_21984);
nand U22959 (N_22959,N_21619,N_21629);
nand U22960 (N_22960,N_22023,N_22139);
nand U22961 (N_22961,N_22411,N_21523);
xnor U22962 (N_22962,N_21835,N_22103);
nand U22963 (N_22963,N_22256,N_21684);
xor U22964 (N_22964,N_21341,N_22219);
nor U22965 (N_22965,N_22339,N_22178);
nand U22966 (N_22966,N_22265,N_21616);
and U22967 (N_22967,N_22113,N_21513);
nand U22968 (N_22968,N_22414,N_21862);
nand U22969 (N_22969,N_21808,N_21371);
or U22970 (N_22970,N_21826,N_21358);
xor U22971 (N_22971,N_22211,N_22068);
and U22972 (N_22972,N_22262,N_21375);
nor U22973 (N_22973,N_21782,N_22246);
xor U22974 (N_22974,N_22049,N_21580);
and U22975 (N_22975,N_21294,N_21501);
and U22976 (N_22976,N_21487,N_21956);
and U22977 (N_22977,N_21444,N_21870);
nand U22978 (N_22978,N_22487,N_22126);
nand U22979 (N_22979,N_21292,N_21656);
nand U22980 (N_22980,N_21405,N_21650);
xor U22981 (N_22981,N_21328,N_21730);
and U22982 (N_22982,N_21762,N_22389);
or U22983 (N_22983,N_22434,N_22374);
nor U22984 (N_22984,N_22386,N_22232);
xor U22985 (N_22985,N_22209,N_21456);
or U22986 (N_22986,N_21362,N_22297);
nor U22987 (N_22987,N_21665,N_21385);
xnor U22988 (N_22988,N_22368,N_21777);
nor U22989 (N_22989,N_21660,N_22371);
xnor U22990 (N_22990,N_21561,N_22104);
or U22991 (N_22991,N_22430,N_22147);
and U22992 (N_22992,N_22133,N_21425);
nand U22993 (N_22993,N_22315,N_22306);
nor U22994 (N_22994,N_22385,N_22140);
nand U22995 (N_22995,N_21875,N_21738);
and U22996 (N_22996,N_22392,N_21859);
or U22997 (N_22997,N_21572,N_22464);
or U22998 (N_22998,N_21705,N_21706);
and U22999 (N_22999,N_21950,N_22154);
nand U23000 (N_23000,N_21467,N_21331);
nor U23001 (N_23001,N_22187,N_21708);
nand U23002 (N_23002,N_22313,N_21542);
nand U23003 (N_23003,N_22110,N_22309);
nor U23004 (N_23004,N_22283,N_22490);
xor U23005 (N_23005,N_22117,N_21843);
nor U23006 (N_23006,N_22495,N_21484);
nand U23007 (N_23007,N_22361,N_21302);
nor U23008 (N_23008,N_21955,N_22136);
nor U23009 (N_23009,N_22476,N_21577);
nand U23010 (N_23010,N_21430,N_22087);
nand U23011 (N_23011,N_22129,N_22316);
and U23012 (N_23012,N_21757,N_22213);
or U23013 (N_23013,N_22245,N_21333);
and U23014 (N_23014,N_22268,N_21479);
nand U23015 (N_23015,N_21620,N_22079);
xnor U23016 (N_23016,N_21939,N_22252);
or U23017 (N_23017,N_22074,N_21707);
or U23018 (N_23018,N_21269,N_22458);
and U23019 (N_23019,N_21907,N_22437);
nand U23020 (N_23020,N_21575,N_21977);
nor U23021 (N_23021,N_22179,N_22128);
nand U23022 (N_23022,N_21327,N_22250);
nor U23023 (N_23023,N_22088,N_21452);
xnor U23024 (N_23024,N_21640,N_22199);
xor U23025 (N_23025,N_21944,N_21549);
and U23026 (N_23026,N_22121,N_22248);
and U23027 (N_23027,N_21455,N_22243);
or U23028 (N_23028,N_21864,N_21500);
nor U23029 (N_23029,N_22375,N_21688);
or U23030 (N_23030,N_21756,N_21748);
and U23031 (N_23031,N_21507,N_22092);
and U23032 (N_23032,N_21426,N_22229);
xor U23033 (N_23033,N_21675,N_22267);
nor U23034 (N_23034,N_21677,N_22247);
nor U23035 (N_23035,N_22150,N_22237);
nand U23036 (N_23036,N_22270,N_22159);
nand U23037 (N_23037,N_21334,N_21338);
nand U23038 (N_23038,N_22071,N_21576);
xnor U23039 (N_23039,N_21653,N_22441);
or U23040 (N_23040,N_22195,N_21349);
nor U23041 (N_23041,N_21618,N_21735);
nand U23042 (N_23042,N_22341,N_22193);
xor U23043 (N_23043,N_21802,N_21403);
xor U23044 (N_23044,N_21877,N_21399);
xnor U23045 (N_23045,N_21632,N_22060);
or U23046 (N_23046,N_21974,N_21428);
or U23047 (N_23047,N_21301,N_22463);
and U23048 (N_23048,N_22001,N_22412);
or U23049 (N_23049,N_21546,N_22449);
nor U23050 (N_23050,N_22236,N_21783);
or U23051 (N_23051,N_21254,N_21852);
xnor U23052 (N_23052,N_22145,N_21911);
nor U23053 (N_23053,N_21482,N_22311);
nand U23054 (N_23054,N_21778,N_21347);
nand U23055 (N_23055,N_21682,N_21915);
nand U23056 (N_23056,N_21435,N_22295);
nor U23057 (N_23057,N_21291,N_22276);
nor U23058 (N_23058,N_22042,N_21904);
or U23059 (N_23059,N_22185,N_22367);
xnor U23060 (N_23060,N_22331,N_21836);
nor U23061 (N_23061,N_21374,N_21816);
nand U23062 (N_23062,N_22073,N_21442);
xnor U23063 (N_23063,N_22031,N_21828);
and U23064 (N_23064,N_21317,N_21581);
nand U23065 (N_23065,N_22021,N_22142);
nor U23066 (N_23066,N_21477,N_22197);
and U23067 (N_23067,N_21922,N_22214);
or U23068 (N_23068,N_21725,N_22018);
or U23069 (N_23069,N_21250,N_21646);
xor U23070 (N_23070,N_22048,N_21849);
and U23071 (N_23071,N_22390,N_22102);
and U23072 (N_23072,N_21896,N_22404);
and U23073 (N_23073,N_22410,N_21623);
xnor U23074 (N_23074,N_21472,N_21772);
nand U23075 (N_23075,N_22355,N_21713);
nor U23076 (N_23076,N_21702,N_22356);
and U23077 (N_23077,N_22284,N_22249);
xor U23078 (N_23078,N_21297,N_21335);
or U23079 (N_23079,N_21368,N_22069);
or U23080 (N_23080,N_21855,N_21307);
or U23081 (N_23081,N_22112,N_22067);
xor U23082 (N_23082,N_22053,N_22466);
nand U23083 (N_23083,N_21453,N_21910);
nor U23084 (N_23084,N_21584,N_21695);
and U23085 (N_23085,N_22260,N_21365);
xnor U23086 (N_23086,N_22155,N_21265);
and U23087 (N_23087,N_22164,N_22288);
nor U23088 (N_23088,N_21562,N_22116);
nand U23089 (N_23089,N_22273,N_22292);
or U23090 (N_23090,N_21891,N_22263);
nor U23091 (N_23091,N_21252,N_22291);
xor U23092 (N_23092,N_22452,N_21900);
or U23093 (N_23093,N_22477,N_21658);
or U23094 (N_23094,N_22014,N_22342);
nor U23095 (N_23095,N_21820,N_22322);
nand U23096 (N_23096,N_21464,N_22393);
and U23097 (N_23097,N_21637,N_21788);
and U23098 (N_23098,N_21943,N_21470);
nand U23099 (N_23099,N_21691,N_21288);
or U23100 (N_23100,N_22301,N_22319);
or U23101 (N_23101,N_21527,N_22217);
nor U23102 (N_23102,N_21940,N_21874);
nand U23103 (N_23103,N_22094,N_22180);
xor U23104 (N_23104,N_21667,N_21687);
and U23105 (N_23105,N_22240,N_21987);
or U23106 (N_23106,N_21343,N_22003);
or U23107 (N_23107,N_21433,N_22181);
nor U23108 (N_23108,N_22206,N_21711);
nand U23109 (N_23109,N_21440,N_21817);
or U23110 (N_23110,N_22166,N_21539);
nor U23111 (N_23111,N_22496,N_21567);
xor U23112 (N_23112,N_22469,N_21636);
or U23113 (N_23113,N_21571,N_21807);
nand U23114 (N_23114,N_21643,N_21902);
or U23115 (N_23115,N_21715,N_21601);
nor U23116 (N_23116,N_21530,N_22152);
xnor U23117 (N_23117,N_21346,N_22091);
and U23118 (N_23118,N_21602,N_22105);
xor U23119 (N_23119,N_21958,N_22170);
nor U23120 (N_23120,N_21999,N_22388);
and U23121 (N_23121,N_21663,N_21740);
nand U23122 (N_23122,N_22403,N_21767);
or U23123 (N_23123,N_22093,N_21809);
nand U23124 (N_23124,N_22298,N_22174);
or U23125 (N_23125,N_21734,N_21726);
nor U23126 (N_23126,N_22480,N_21623);
nor U23127 (N_23127,N_22051,N_22144);
nor U23128 (N_23128,N_22272,N_21416);
nor U23129 (N_23129,N_22206,N_21942);
and U23130 (N_23130,N_21815,N_22374);
and U23131 (N_23131,N_22404,N_21520);
or U23132 (N_23132,N_21825,N_22268);
or U23133 (N_23133,N_21660,N_21272);
and U23134 (N_23134,N_21767,N_21854);
or U23135 (N_23135,N_22468,N_21989);
nor U23136 (N_23136,N_22285,N_21437);
and U23137 (N_23137,N_22401,N_21932);
nor U23138 (N_23138,N_21681,N_22082);
xor U23139 (N_23139,N_22164,N_22254);
xnor U23140 (N_23140,N_22300,N_22169);
and U23141 (N_23141,N_21700,N_21556);
xnor U23142 (N_23142,N_21963,N_21950);
nor U23143 (N_23143,N_22002,N_21958);
nor U23144 (N_23144,N_21297,N_21756);
xor U23145 (N_23145,N_21649,N_22493);
or U23146 (N_23146,N_22069,N_21804);
nor U23147 (N_23147,N_21841,N_22066);
or U23148 (N_23148,N_22295,N_21657);
and U23149 (N_23149,N_21932,N_21635);
and U23150 (N_23150,N_21476,N_21356);
xnor U23151 (N_23151,N_22319,N_21768);
xnor U23152 (N_23152,N_21390,N_22384);
nor U23153 (N_23153,N_21735,N_22462);
nor U23154 (N_23154,N_22489,N_21956);
or U23155 (N_23155,N_22393,N_21403);
nor U23156 (N_23156,N_22163,N_21390);
nor U23157 (N_23157,N_22365,N_21713);
nand U23158 (N_23158,N_21347,N_21946);
or U23159 (N_23159,N_21878,N_21870);
and U23160 (N_23160,N_21558,N_22118);
nand U23161 (N_23161,N_22030,N_21412);
nor U23162 (N_23162,N_22305,N_21608);
and U23163 (N_23163,N_21771,N_21521);
xor U23164 (N_23164,N_21986,N_22328);
nor U23165 (N_23165,N_21391,N_22262);
or U23166 (N_23166,N_21615,N_21523);
or U23167 (N_23167,N_22200,N_21914);
nand U23168 (N_23168,N_22186,N_22010);
nand U23169 (N_23169,N_22030,N_21723);
and U23170 (N_23170,N_21913,N_21626);
and U23171 (N_23171,N_21799,N_22006);
xor U23172 (N_23172,N_21946,N_22233);
or U23173 (N_23173,N_22018,N_21433);
and U23174 (N_23174,N_22342,N_22344);
nor U23175 (N_23175,N_22096,N_21757);
or U23176 (N_23176,N_21837,N_22010);
and U23177 (N_23177,N_21791,N_22176);
nand U23178 (N_23178,N_21895,N_21669);
xnor U23179 (N_23179,N_21492,N_21946);
xnor U23180 (N_23180,N_22339,N_21320);
xnor U23181 (N_23181,N_21276,N_22305);
nand U23182 (N_23182,N_22060,N_21576);
nand U23183 (N_23183,N_22341,N_21882);
nor U23184 (N_23184,N_21523,N_22155);
xor U23185 (N_23185,N_21984,N_21314);
nand U23186 (N_23186,N_21953,N_22012);
and U23187 (N_23187,N_22003,N_21446);
or U23188 (N_23188,N_21936,N_22204);
or U23189 (N_23189,N_21516,N_21997);
nand U23190 (N_23190,N_22071,N_21418);
nor U23191 (N_23191,N_22392,N_21391);
nor U23192 (N_23192,N_22053,N_21789);
nor U23193 (N_23193,N_22184,N_21779);
xor U23194 (N_23194,N_22222,N_21985);
nor U23195 (N_23195,N_21620,N_22341);
nor U23196 (N_23196,N_21477,N_22183);
nand U23197 (N_23197,N_22307,N_21311);
nand U23198 (N_23198,N_22380,N_21624);
xnor U23199 (N_23199,N_21432,N_22291);
nor U23200 (N_23200,N_21838,N_21938);
and U23201 (N_23201,N_21743,N_21363);
xor U23202 (N_23202,N_21459,N_22071);
and U23203 (N_23203,N_22366,N_21369);
xnor U23204 (N_23204,N_22413,N_22233);
or U23205 (N_23205,N_22076,N_22235);
nor U23206 (N_23206,N_22101,N_22447);
or U23207 (N_23207,N_21556,N_22022);
or U23208 (N_23208,N_21345,N_22045);
and U23209 (N_23209,N_21553,N_21970);
nor U23210 (N_23210,N_22024,N_22455);
nor U23211 (N_23211,N_21709,N_22333);
or U23212 (N_23212,N_22071,N_22401);
xnor U23213 (N_23213,N_21482,N_22406);
and U23214 (N_23214,N_21778,N_21387);
nor U23215 (N_23215,N_21409,N_21632);
xor U23216 (N_23216,N_21578,N_21553);
and U23217 (N_23217,N_22403,N_22349);
nand U23218 (N_23218,N_22350,N_22300);
and U23219 (N_23219,N_21672,N_22053);
and U23220 (N_23220,N_21611,N_21281);
xor U23221 (N_23221,N_21785,N_22179);
xnor U23222 (N_23222,N_21930,N_21640);
or U23223 (N_23223,N_21924,N_21606);
nor U23224 (N_23224,N_21614,N_22145);
and U23225 (N_23225,N_22349,N_21273);
and U23226 (N_23226,N_22111,N_22060);
and U23227 (N_23227,N_21589,N_21553);
and U23228 (N_23228,N_21577,N_21560);
nor U23229 (N_23229,N_22300,N_21463);
and U23230 (N_23230,N_21586,N_22318);
and U23231 (N_23231,N_21676,N_21869);
and U23232 (N_23232,N_21264,N_22214);
or U23233 (N_23233,N_21661,N_21730);
or U23234 (N_23234,N_21761,N_22086);
or U23235 (N_23235,N_22191,N_22089);
nand U23236 (N_23236,N_22044,N_21560);
or U23237 (N_23237,N_21909,N_21289);
xnor U23238 (N_23238,N_22441,N_21641);
nand U23239 (N_23239,N_22157,N_21699);
nand U23240 (N_23240,N_21907,N_21797);
nand U23241 (N_23241,N_22026,N_22088);
nand U23242 (N_23242,N_22199,N_21580);
nor U23243 (N_23243,N_22147,N_21509);
and U23244 (N_23244,N_22411,N_21556);
nor U23245 (N_23245,N_22347,N_21367);
nand U23246 (N_23246,N_21410,N_22461);
or U23247 (N_23247,N_21888,N_22498);
or U23248 (N_23248,N_22323,N_21262);
xnor U23249 (N_23249,N_21533,N_22270);
and U23250 (N_23250,N_21432,N_21538);
nor U23251 (N_23251,N_21847,N_21587);
nor U23252 (N_23252,N_21917,N_21469);
xor U23253 (N_23253,N_21552,N_22124);
nand U23254 (N_23254,N_21780,N_21513);
nand U23255 (N_23255,N_22273,N_21800);
and U23256 (N_23256,N_21578,N_22106);
and U23257 (N_23257,N_21350,N_21306);
nand U23258 (N_23258,N_21859,N_21650);
nand U23259 (N_23259,N_22360,N_21719);
and U23260 (N_23260,N_21665,N_21910);
xor U23261 (N_23261,N_21256,N_21613);
xor U23262 (N_23262,N_21679,N_21600);
xor U23263 (N_23263,N_21856,N_21758);
nand U23264 (N_23264,N_21947,N_21573);
nand U23265 (N_23265,N_22005,N_22050);
nand U23266 (N_23266,N_22240,N_22347);
xnor U23267 (N_23267,N_21369,N_21463);
or U23268 (N_23268,N_21621,N_22013);
xnor U23269 (N_23269,N_21391,N_21468);
and U23270 (N_23270,N_21934,N_21747);
or U23271 (N_23271,N_22057,N_22343);
xor U23272 (N_23272,N_21691,N_21493);
nand U23273 (N_23273,N_21630,N_21911);
nand U23274 (N_23274,N_21991,N_22404);
xnor U23275 (N_23275,N_21841,N_22431);
nand U23276 (N_23276,N_22431,N_22023);
nor U23277 (N_23277,N_21396,N_22084);
nor U23278 (N_23278,N_21338,N_22067);
xor U23279 (N_23279,N_22302,N_22217);
or U23280 (N_23280,N_21352,N_21828);
nand U23281 (N_23281,N_21602,N_22216);
nor U23282 (N_23282,N_21293,N_21920);
xor U23283 (N_23283,N_21708,N_21436);
and U23284 (N_23284,N_21385,N_22090);
nand U23285 (N_23285,N_21786,N_21760);
nand U23286 (N_23286,N_22109,N_22266);
nor U23287 (N_23287,N_21388,N_22165);
and U23288 (N_23288,N_22478,N_22084);
nor U23289 (N_23289,N_22174,N_21546);
nor U23290 (N_23290,N_21914,N_22091);
or U23291 (N_23291,N_22492,N_22244);
xor U23292 (N_23292,N_21756,N_22176);
or U23293 (N_23293,N_21309,N_22062);
nor U23294 (N_23294,N_21406,N_21580);
nor U23295 (N_23295,N_21761,N_21341);
nor U23296 (N_23296,N_21770,N_21851);
nor U23297 (N_23297,N_22252,N_21501);
nor U23298 (N_23298,N_21961,N_21746);
nor U23299 (N_23299,N_21319,N_21614);
nand U23300 (N_23300,N_21635,N_21568);
and U23301 (N_23301,N_21937,N_21512);
and U23302 (N_23302,N_22074,N_21481);
nor U23303 (N_23303,N_21534,N_21490);
xnor U23304 (N_23304,N_21283,N_21774);
xor U23305 (N_23305,N_21476,N_21300);
nor U23306 (N_23306,N_21970,N_22486);
nor U23307 (N_23307,N_21924,N_21422);
or U23308 (N_23308,N_21302,N_22415);
nor U23309 (N_23309,N_22232,N_22262);
or U23310 (N_23310,N_22359,N_21494);
xnor U23311 (N_23311,N_22215,N_21595);
xor U23312 (N_23312,N_21999,N_22469);
nand U23313 (N_23313,N_21628,N_22444);
and U23314 (N_23314,N_22215,N_21822);
nand U23315 (N_23315,N_21456,N_22044);
or U23316 (N_23316,N_22016,N_22454);
nor U23317 (N_23317,N_21999,N_22311);
nor U23318 (N_23318,N_22272,N_21289);
and U23319 (N_23319,N_21485,N_22309);
nor U23320 (N_23320,N_21507,N_21514);
xnor U23321 (N_23321,N_21657,N_21574);
and U23322 (N_23322,N_22199,N_22111);
xor U23323 (N_23323,N_21433,N_21447);
nor U23324 (N_23324,N_21460,N_22475);
or U23325 (N_23325,N_21669,N_21951);
or U23326 (N_23326,N_21803,N_22297);
or U23327 (N_23327,N_22484,N_22028);
nand U23328 (N_23328,N_21461,N_22094);
nand U23329 (N_23329,N_22213,N_21814);
and U23330 (N_23330,N_22228,N_21712);
or U23331 (N_23331,N_21841,N_21431);
xor U23332 (N_23332,N_21761,N_21524);
nand U23333 (N_23333,N_21426,N_21988);
xnor U23334 (N_23334,N_21699,N_22334);
xor U23335 (N_23335,N_21787,N_22416);
or U23336 (N_23336,N_22018,N_21872);
or U23337 (N_23337,N_22386,N_22331);
xnor U23338 (N_23338,N_21675,N_21478);
nor U23339 (N_23339,N_21381,N_21909);
or U23340 (N_23340,N_21962,N_22040);
xor U23341 (N_23341,N_22473,N_21328);
nand U23342 (N_23342,N_22401,N_22266);
or U23343 (N_23343,N_21371,N_21490);
nor U23344 (N_23344,N_22013,N_22298);
xor U23345 (N_23345,N_21920,N_22326);
nor U23346 (N_23346,N_22366,N_22303);
or U23347 (N_23347,N_21385,N_21611);
nand U23348 (N_23348,N_22007,N_22182);
xnor U23349 (N_23349,N_22091,N_21946);
and U23350 (N_23350,N_21976,N_22183);
nor U23351 (N_23351,N_21621,N_22017);
nand U23352 (N_23352,N_22368,N_22224);
and U23353 (N_23353,N_22460,N_21290);
nand U23354 (N_23354,N_21991,N_21529);
nor U23355 (N_23355,N_22469,N_22495);
and U23356 (N_23356,N_21421,N_21333);
nand U23357 (N_23357,N_21594,N_21345);
nand U23358 (N_23358,N_21833,N_21308);
nand U23359 (N_23359,N_21451,N_21849);
nand U23360 (N_23360,N_21431,N_21930);
and U23361 (N_23361,N_22397,N_22292);
xnor U23362 (N_23362,N_22054,N_21762);
nand U23363 (N_23363,N_22030,N_21652);
xor U23364 (N_23364,N_21684,N_21269);
nand U23365 (N_23365,N_22315,N_21320);
or U23366 (N_23366,N_22426,N_21341);
or U23367 (N_23367,N_22009,N_22233);
nand U23368 (N_23368,N_21272,N_21851);
nor U23369 (N_23369,N_21626,N_21298);
nand U23370 (N_23370,N_21809,N_22145);
nor U23371 (N_23371,N_21494,N_21597);
and U23372 (N_23372,N_22309,N_21990);
nand U23373 (N_23373,N_21861,N_22387);
and U23374 (N_23374,N_22455,N_21357);
or U23375 (N_23375,N_21441,N_21470);
and U23376 (N_23376,N_22217,N_21628);
nand U23377 (N_23377,N_22030,N_22341);
nand U23378 (N_23378,N_22081,N_21302);
and U23379 (N_23379,N_21350,N_21874);
or U23380 (N_23380,N_21958,N_21903);
xnor U23381 (N_23381,N_21738,N_21294);
nand U23382 (N_23382,N_22405,N_22135);
xor U23383 (N_23383,N_21596,N_21822);
nor U23384 (N_23384,N_21984,N_22412);
nor U23385 (N_23385,N_22442,N_21641);
xnor U23386 (N_23386,N_21434,N_22412);
or U23387 (N_23387,N_21597,N_21312);
nor U23388 (N_23388,N_21772,N_22376);
nor U23389 (N_23389,N_21300,N_21591);
nand U23390 (N_23390,N_21413,N_22304);
nor U23391 (N_23391,N_22017,N_21852);
or U23392 (N_23392,N_22296,N_21921);
or U23393 (N_23393,N_22347,N_21510);
and U23394 (N_23394,N_21616,N_21678);
or U23395 (N_23395,N_22139,N_21589);
nor U23396 (N_23396,N_21562,N_21804);
or U23397 (N_23397,N_21576,N_21537);
nor U23398 (N_23398,N_22233,N_21614);
xor U23399 (N_23399,N_22365,N_21928);
and U23400 (N_23400,N_22254,N_22018);
nand U23401 (N_23401,N_21312,N_21766);
and U23402 (N_23402,N_22499,N_21889);
nor U23403 (N_23403,N_22456,N_21603);
and U23404 (N_23404,N_21363,N_22347);
or U23405 (N_23405,N_21356,N_21452);
xnor U23406 (N_23406,N_21579,N_21370);
and U23407 (N_23407,N_21693,N_21302);
or U23408 (N_23408,N_21870,N_22336);
nor U23409 (N_23409,N_21475,N_22368);
nor U23410 (N_23410,N_21253,N_21405);
nand U23411 (N_23411,N_21642,N_22059);
xor U23412 (N_23412,N_22018,N_22292);
xnor U23413 (N_23413,N_21730,N_22481);
nand U23414 (N_23414,N_21937,N_21924);
xor U23415 (N_23415,N_21739,N_21680);
or U23416 (N_23416,N_22071,N_21426);
or U23417 (N_23417,N_22115,N_21576);
and U23418 (N_23418,N_21309,N_21524);
xnor U23419 (N_23419,N_21877,N_22341);
nand U23420 (N_23420,N_22268,N_21767);
nand U23421 (N_23421,N_22361,N_21369);
or U23422 (N_23422,N_22342,N_22392);
or U23423 (N_23423,N_21846,N_22315);
or U23424 (N_23424,N_21546,N_21948);
and U23425 (N_23425,N_22273,N_22387);
and U23426 (N_23426,N_21795,N_22484);
xnor U23427 (N_23427,N_22321,N_22126);
nor U23428 (N_23428,N_21350,N_22275);
nand U23429 (N_23429,N_22446,N_22401);
nor U23430 (N_23430,N_22170,N_21435);
xor U23431 (N_23431,N_22092,N_21266);
nand U23432 (N_23432,N_22145,N_21553);
or U23433 (N_23433,N_22302,N_22448);
xnor U23434 (N_23434,N_21982,N_22108);
or U23435 (N_23435,N_21575,N_21860);
or U23436 (N_23436,N_22223,N_21985);
and U23437 (N_23437,N_22486,N_21837);
xnor U23438 (N_23438,N_22486,N_22344);
and U23439 (N_23439,N_22443,N_21998);
nand U23440 (N_23440,N_22200,N_22149);
nor U23441 (N_23441,N_22034,N_21511);
nor U23442 (N_23442,N_22099,N_21874);
and U23443 (N_23443,N_22157,N_22463);
or U23444 (N_23444,N_21622,N_21566);
xor U23445 (N_23445,N_21253,N_22270);
nand U23446 (N_23446,N_21971,N_22280);
nand U23447 (N_23447,N_21306,N_21967);
nand U23448 (N_23448,N_22149,N_21453);
xnor U23449 (N_23449,N_22216,N_22250);
nand U23450 (N_23450,N_21840,N_21466);
nand U23451 (N_23451,N_21663,N_22286);
or U23452 (N_23452,N_22344,N_21746);
nor U23453 (N_23453,N_22075,N_21826);
nand U23454 (N_23454,N_21448,N_22315);
and U23455 (N_23455,N_22103,N_22388);
nor U23456 (N_23456,N_22164,N_22446);
xor U23457 (N_23457,N_21960,N_22148);
nand U23458 (N_23458,N_22368,N_22019);
and U23459 (N_23459,N_22472,N_21605);
and U23460 (N_23460,N_21904,N_21850);
xnor U23461 (N_23461,N_22401,N_22022);
or U23462 (N_23462,N_21818,N_22446);
xor U23463 (N_23463,N_21477,N_22342);
or U23464 (N_23464,N_22113,N_21697);
nand U23465 (N_23465,N_21960,N_21927);
nor U23466 (N_23466,N_21493,N_21607);
or U23467 (N_23467,N_21934,N_21977);
or U23468 (N_23468,N_22007,N_21724);
nor U23469 (N_23469,N_21259,N_21662);
or U23470 (N_23470,N_22034,N_22215);
nand U23471 (N_23471,N_21607,N_21382);
and U23472 (N_23472,N_22039,N_21572);
xor U23473 (N_23473,N_21287,N_21329);
and U23474 (N_23474,N_21533,N_22095);
xnor U23475 (N_23475,N_22204,N_21461);
and U23476 (N_23476,N_21908,N_21301);
nor U23477 (N_23477,N_22498,N_22167);
nand U23478 (N_23478,N_22408,N_21904);
and U23479 (N_23479,N_21824,N_21898);
nor U23480 (N_23480,N_21264,N_21643);
nor U23481 (N_23481,N_22241,N_21757);
and U23482 (N_23482,N_21623,N_22460);
nand U23483 (N_23483,N_21603,N_21627);
nand U23484 (N_23484,N_21952,N_22183);
nand U23485 (N_23485,N_21416,N_21798);
or U23486 (N_23486,N_22111,N_22150);
nor U23487 (N_23487,N_22010,N_22165);
nand U23488 (N_23488,N_22335,N_22150);
nor U23489 (N_23489,N_21933,N_21721);
nor U23490 (N_23490,N_21528,N_21445);
and U23491 (N_23491,N_22419,N_22354);
or U23492 (N_23492,N_22167,N_21495);
or U23493 (N_23493,N_21668,N_22136);
nor U23494 (N_23494,N_21345,N_21370);
nor U23495 (N_23495,N_21313,N_22105);
xor U23496 (N_23496,N_21392,N_21450);
or U23497 (N_23497,N_21804,N_21492);
or U23498 (N_23498,N_21415,N_22253);
xnor U23499 (N_23499,N_22483,N_21547);
nand U23500 (N_23500,N_21812,N_22085);
nor U23501 (N_23501,N_21816,N_22000);
or U23502 (N_23502,N_22387,N_21311);
and U23503 (N_23503,N_22444,N_21301);
nand U23504 (N_23504,N_22232,N_21999);
or U23505 (N_23505,N_21863,N_21907);
or U23506 (N_23506,N_21952,N_21811);
and U23507 (N_23507,N_22024,N_22051);
xnor U23508 (N_23508,N_21729,N_21629);
xnor U23509 (N_23509,N_22318,N_21671);
nand U23510 (N_23510,N_22153,N_22126);
or U23511 (N_23511,N_21993,N_21297);
nor U23512 (N_23512,N_22326,N_22170);
xor U23513 (N_23513,N_22282,N_21814);
nor U23514 (N_23514,N_21472,N_21406);
or U23515 (N_23515,N_22105,N_21263);
nand U23516 (N_23516,N_22389,N_21796);
nor U23517 (N_23517,N_21676,N_21627);
xor U23518 (N_23518,N_22349,N_22482);
nand U23519 (N_23519,N_22458,N_21398);
nand U23520 (N_23520,N_22006,N_22202);
or U23521 (N_23521,N_21645,N_21264);
nand U23522 (N_23522,N_21432,N_21425);
and U23523 (N_23523,N_21981,N_22273);
nand U23524 (N_23524,N_22340,N_21986);
or U23525 (N_23525,N_21939,N_22456);
xnor U23526 (N_23526,N_22302,N_21845);
xnor U23527 (N_23527,N_21956,N_22480);
nor U23528 (N_23528,N_22152,N_21827);
nor U23529 (N_23529,N_21668,N_21446);
and U23530 (N_23530,N_22066,N_21551);
nand U23531 (N_23531,N_22049,N_21318);
nand U23532 (N_23532,N_22427,N_22474);
xnor U23533 (N_23533,N_21537,N_22161);
and U23534 (N_23534,N_22283,N_22184);
nor U23535 (N_23535,N_22456,N_22486);
or U23536 (N_23536,N_21905,N_22266);
and U23537 (N_23537,N_21952,N_22364);
or U23538 (N_23538,N_22112,N_21978);
and U23539 (N_23539,N_22198,N_21665);
nand U23540 (N_23540,N_21691,N_22347);
or U23541 (N_23541,N_21537,N_21513);
xor U23542 (N_23542,N_21821,N_21626);
or U23543 (N_23543,N_21656,N_21593);
nor U23544 (N_23544,N_22137,N_21402);
nor U23545 (N_23545,N_21776,N_22277);
or U23546 (N_23546,N_22498,N_21336);
and U23547 (N_23547,N_22496,N_22006);
nand U23548 (N_23548,N_22001,N_21304);
and U23549 (N_23549,N_22420,N_22241);
or U23550 (N_23550,N_21488,N_22126);
nor U23551 (N_23551,N_21706,N_21380);
and U23552 (N_23552,N_21392,N_21754);
and U23553 (N_23553,N_21374,N_21809);
or U23554 (N_23554,N_21465,N_22260);
and U23555 (N_23555,N_21282,N_22002);
xor U23556 (N_23556,N_21992,N_22229);
and U23557 (N_23557,N_21687,N_21466);
nand U23558 (N_23558,N_21737,N_22491);
xnor U23559 (N_23559,N_21479,N_22086);
and U23560 (N_23560,N_22392,N_21418);
xnor U23561 (N_23561,N_22251,N_21677);
nor U23562 (N_23562,N_21952,N_22271);
or U23563 (N_23563,N_21685,N_21663);
or U23564 (N_23564,N_22170,N_22024);
nand U23565 (N_23565,N_21940,N_22411);
nand U23566 (N_23566,N_21277,N_21616);
xnor U23567 (N_23567,N_21708,N_21759);
and U23568 (N_23568,N_21903,N_22371);
and U23569 (N_23569,N_22263,N_21499);
and U23570 (N_23570,N_22191,N_22351);
and U23571 (N_23571,N_21278,N_21501);
or U23572 (N_23572,N_21762,N_21503);
nand U23573 (N_23573,N_22045,N_21734);
nor U23574 (N_23574,N_22379,N_21412);
nor U23575 (N_23575,N_21775,N_22311);
nor U23576 (N_23576,N_21340,N_21923);
and U23577 (N_23577,N_22377,N_21839);
and U23578 (N_23578,N_21612,N_22179);
nand U23579 (N_23579,N_21266,N_21642);
xnor U23580 (N_23580,N_21680,N_22060);
xor U23581 (N_23581,N_22287,N_22422);
or U23582 (N_23582,N_21829,N_22376);
and U23583 (N_23583,N_21944,N_21498);
nor U23584 (N_23584,N_21689,N_21784);
and U23585 (N_23585,N_22298,N_22302);
xor U23586 (N_23586,N_21701,N_21570);
nand U23587 (N_23587,N_22360,N_21729);
nand U23588 (N_23588,N_21917,N_22240);
nand U23589 (N_23589,N_21907,N_21275);
xor U23590 (N_23590,N_21745,N_22300);
nor U23591 (N_23591,N_21359,N_21522);
nor U23592 (N_23592,N_21526,N_21303);
or U23593 (N_23593,N_21782,N_21353);
or U23594 (N_23594,N_21900,N_21727);
and U23595 (N_23595,N_21483,N_21509);
xor U23596 (N_23596,N_21751,N_21289);
nand U23597 (N_23597,N_21631,N_21965);
xnor U23598 (N_23598,N_21619,N_21945);
nand U23599 (N_23599,N_22115,N_21831);
nand U23600 (N_23600,N_22161,N_22017);
nor U23601 (N_23601,N_21728,N_21946);
or U23602 (N_23602,N_21706,N_21711);
nor U23603 (N_23603,N_21415,N_21418);
nor U23604 (N_23604,N_21555,N_21473);
and U23605 (N_23605,N_22316,N_22360);
xnor U23606 (N_23606,N_21717,N_21788);
or U23607 (N_23607,N_22350,N_22348);
xnor U23608 (N_23608,N_21296,N_22407);
xnor U23609 (N_23609,N_22082,N_22132);
or U23610 (N_23610,N_21564,N_22061);
and U23611 (N_23611,N_21854,N_21305);
xor U23612 (N_23612,N_21647,N_21502);
xnor U23613 (N_23613,N_22424,N_21832);
xor U23614 (N_23614,N_22370,N_22196);
nor U23615 (N_23615,N_22314,N_22425);
or U23616 (N_23616,N_21792,N_21346);
nor U23617 (N_23617,N_21933,N_22231);
nand U23618 (N_23618,N_22403,N_22186);
xor U23619 (N_23619,N_22272,N_21308);
or U23620 (N_23620,N_21858,N_22499);
xor U23621 (N_23621,N_21652,N_21725);
and U23622 (N_23622,N_21322,N_21554);
or U23623 (N_23623,N_21688,N_21548);
xor U23624 (N_23624,N_21528,N_22488);
and U23625 (N_23625,N_22305,N_21889);
nand U23626 (N_23626,N_22031,N_21600);
nand U23627 (N_23627,N_21472,N_21705);
xnor U23628 (N_23628,N_21758,N_22059);
nor U23629 (N_23629,N_21710,N_21913);
nand U23630 (N_23630,N_22010,N_21900);
xor U23631 (N_23631,N_22345,N_21825);
nand U23632 (N_23632,N_21456,N_21352);
xor U23633 (N_23633,N_21805,N_21710);
and U23634 (N_23634,N_21667,N_21788);
and U23635 (N_23635,N_21801,N_22038);
nand U23636 (N_23636,N_21362,N_21646);
nor U23637 (N_23637,N_21571,N_21822);
nand U23638 (N_23638,N_22224,N_22341);
nand U23639 (N_23639,N_21963,N_21714);
xor U23640 (N_23640,N_22021,N_22076);
or U23641 (N_23641,N_21633,N_22450);
nand U23642 (N_23642,N_21927,N_22494);
or U23643 (N_23643,N_21931,N_21886);
xor U23644 (N_23644,N_22231,N_21493);
xor U23645 (N_23645,N_21616,N_21670);
xnor U23646 (N_23646,N_22455,N_22413);
nand U23647 (N_23647,N_21386,N_22376);
or U23648 (N_23648,N_21916,N_22446);
nand U23649 (N_23649,N_21725,N_21680);
nand U23650 (N_23650,N_22367,N_22468);
and U23651 (N_23651,N_21784,N_21579);
or U23652 (N_23652,N_21266,N_22293);
nand U23653 (N_23653,N_21753,N_22238);
nand U23654 (N_23654,N_22384,N_21702);
and U23655 (N_23655,N_21618,N_21682);
nand U23656 (N_23656,N_22094,N_21530);
or U23657 (N_23657,N_21545,N_22129);
nor U23658 (N_23658,N_21769,N_22147);
xnor U23659 (N_23659,N_21880,N_22133);
or U23660 (N_23660,N_21508,N_22031);
or U23661 (N_23661,N_21408,N_22338);
and U23662 (N_23662,N_21336,N_22276);
and U23663 (N_23663,N_21546,N_22235);
xor U23664 (N_23664,N_22369,N_22002);
nand U23665 (N_23665,N_21412,N_21415);
xnor U23666 (N_23666,N_22432,N_21986);
nand U23667 (N_23667,N_21368,N_21448);
and U23668 (N_23668,N_21455,N_21471);
and U23669 (N_23669,N_22000,N_21266);
and U23670 (N_23670,N_21518,N_21652);
nand U23671 (N_23671,N_21502,N_21613);
or U23672 (N_23672,N_21624,N_22072);
nand U23673 (N_23673,N_21966,N_21688);
xor U23674 (N_23674,N_21479,N_21383);
nor U23675 (N_23675,N_21417,N_22176);
or U23676 (N_23676,N_22125,N_22484);
or U23677 (N_23677,N_21315,N_22486);
nand U23678 (N_23678,N_22441,N_21846);
nand U23679 (N_23679,N_21666,N_21446);
nand U23680 (N_23680,N_22093,N_21802);
and U23681 (N_23681,N_22386,N_21602);
nand U23682 (N_23682,N_21441,N_21653);
and U23683 (N_23683,N_21688,N_21800);
or U23684 (N_23684,N_21451,N_21708);
nand U23685 (N_23685,N_22363,N_21456);
nand U23686 (N_23686,N_21560,N_21254);
nand U23687 (N_23687,N_21629,N_22020);
and U23688 (N_23688,N_22027,N_21988);
xor U23689 (N_23689,N_21613,N_21884);
nor U23690 (N_23690,N_21309,N_21395);
nand U23691 (N_23691,N_21980,N_22296);
nand U23692 (N_23692,N_21983,N_21592);
nor U23693 (N_23693,N_21565,N_22293);
nand U23694 (N_23694,N_21574,N_22302);
and U23695 (N_23695,N_21292,N_21496);
xor U23696 (N_23696,N_22354,N_21867);
nand U23697 (N_23697,N_22081,N_21854);
and U23698 (N_23698,N_22042,N_22377);
xnor U23699 (N_23699,N_21487,N_21400);
nand U23700 (N_23700,N_21295,N_22050);
nand U23701 (N_23701,N_21365,N_22253);
xnor U23702 (N_23702,N_21307,N_22172);
nor U23703 (N_23703,N_21435,N_22094);
nand U23704 (N_23704,N_22446,N_21891);
xnor U23705 (N_23705,N_22469,N_21751);
or U23706 (N_23706,N_22461,N_22479);
xor U23707 (N_23707,N_22251,N_22343);
xnor U23708 (N_23708,N_21356,N_22369);
nand U23709 (N_23709,N_22210,N_22190);
nor U23710 (N_23710,N_22222,N_21831);
and U23711 (N_23711,N_21978,N_22095);
or U23712 (N_23712,N_22256,N_21673);
and U23713 (N_23713,N_22347,N_21963);
nor U23714 (N_23714,N_22117,N_22388);
xor U23715 (N_23715,N_21379,N_21306);
nand U23716 (N_23716,N_21486,N_22002);
or U23717 (N_23717,N_22039,N_22309);
or U23718 (N_23718,N_21720,N_22227);
xnor U23719 (N_23719,N_21432,N_21504);
and U23720 (N_23720,N_22418,N_21631);
nand U23721 (N_23721,N_22175,N_21849);
xor U23722 (N_23722,N_21299,N_22458);
nor U23723 (N_23723,N_21912,N_21325);
or U23724 (N_23724,N_21533,N_21464);
nor U23725 (N_23725,N_22078,N_22052);
nand U23726 (N_23726,N_21555,N_21602);
and U23727 (N_23727,N_22397,N_22019);
or U23728 (N_23728,N_22016,N_22114);
xor U23729 (N_23729,N_21574,N_21910);
and U23730 (N_23730,N_21735,N_21566);
xnor U23731 (N_23731,N_21827,N_22168);
nor U23732 (N_23732,N_22460,N_22252);
or U23733 (N_23733,N_21867,N_22448);
and U23734 (N_23734,N_21681,N_22347);
or U23735 (N_23735,N_22434,N_22363);
nand U23736 (N_23736,N_21703,N_21511);
nor U23737 (N_23737,N_21491,N_22252);
or U23738 (N_23738,N_21984,N_22437);
xnor U23739 (N_23739,N_21831,N_22225);
and U23740 (N_23740,N_21929,N_21566);
and U23741 (N_23741,N_21583,N_21899);
xor U23742 (N_23742,N_21576,N_22439);
or U23743 (N_23743,N_21803,N_21394);
nand U23744 (N_23744,N_22458,N_22413);
or U23745 (N_23745,N_21886,N_21481);
nand U23746 (N_23746,N_21884,N_21916);
or U23747 (N_23747,N_22022,N_21272);
nor U23748 (N_23748,N_21278,N_22212);
nand U23749 (N_23749,N_22351,N_22456);
nor U23750 (N_23750,N_22815,N_23596);
xor U23751 (N_23751,N_23686,N_22810);
xnor U23752 (N_23752,N_23463,N_23280);
nor U23753 (N_23753,N_22833,N_23152);
or U23754 (N_23754,N_22874,N_22883);
nand U23755 (N_23755,N_23481,N_23292);
xor U23756 (N_23756,N_23681,N_22727);
nand U23757 (N_23757,N_22732,N_22812);
xnor U23758 (N_23758,N_22929,N_23005);
xor U23759 (N_23759,N_22843,N_22565);
and U23760 (N_23760,N_22733,N_23546);
and U23761 (N_23761,N_23267,N_23568);
and U23762 (N_23762,N_22749,N_23637);
nor U23763 (N_23763,N_23294,N_22726);
and U23764 (N_23764,N_22731,N_22647);
nor U23765 (N_23765,N_22816,N_22662);
or U23766 (N_23766,N_23213,N_23226);
and U23767 (N_23767,N_22899,N_22796);
nand U23768 (N_23768,N_22854,N_23203);
and U23769 (N_23769,N_23003,N_23034);
or U23770 (N_23770,N_22673,N_23235);
and U23771 (N_23771,N_23351,N_23160);
and U23772 (N_23772,N_23636,N_23266);
or U23773 (N_23773,N_23653,N_23166);
and U23774 (N_23774,N_23474,N_23106);
or U23775 (N_23775,N_22898,N_22533);
nor U23776 (N_23776,N_23286,N_22504);
xnor U23777 (N_23777,N_23397,N_23483);
nor U23778 (N_23778,N_23317,N_23308);
nand U23779 (N_23779,N_23642,N_23009);
and U23780 (N_23780,N_23222,N_22893);
and U23781 (N_23781,N_23214,N_22592);
and U23782 (N_23782,N_22572,N_22758);
xnor U23783 (N_23783,N_22763,N_23279);
or U23784 (N_23784,N_23219,N_23053);
or U23785 (N_23785,N_23320,N_22997);
or U23786 (N_23786,N_23698,N_23412);
and U23787 (N_23787,N_22665,N_22743);
nor U23788 (N_23788,N_23526,N_23158);
or U23789 (N_23789,N_22660,N_23103);
nor U23790 (N_23790,N_23418,N_22806);
and U23791 (N_23791,N_22531,N_23440);
or U23792 (N_23792,N_23304,N_22922);
xor U23793 (N_23793,N_23259,N_22503);
nand U23794 (N_23794,N_23366,N_23101);
xnor U23795 (N_23795,N_22719,N_23002);
and U23796 (N_23796,N_23480,N_22517);
nand U23797 (N_23797,N_22721,N_22961);
nand U23798 (N_23798,N_23287,N_22516);
xor U23799 (N_23799,N_23610,N_22829);
xor U23800 (N_23800,N_23169,N_23689);
xor U23801 (N_23801,N_23515,N_23123);
xor U23802 (N_23802,N_23690,N_22996);
nor U23803 (N_23803,N_23665,N_22539);
nand U23804 (N_23804,N_22958,N_22973);
or U23805 (N_23805,N_23254,N_22663);
or U23806 (N_23806,N_23477,N_23371);
xnor U23807 (N_23807,N_23672,N_22793);
xor U23808 (N_23808,N_23110,N_22571);
and U23809 (N_23809,N_23640,N_22676);
nor U23810 (N_23810,N_22638,N_23726);
nand U23811 (N_23811,N_23602,N_22677);
or U23812 (N_23812,N_23116,N_22813);
nor U23813 (N_23813,N_23673,N_23646);
xnor U23814 (N_23814,N_22937,N_23413);
or U23815 (N_23815,N_23291,N_22604);
and U23816 (N_23816,N_22881,N_23422);
or U23817 (N_23817,N_23258,N_23746);
nand U23818 (N_23818,N_22701,N_22695);
and U23819 (N_23819,N_22532,N_23056);
or U23820 (N_23820,N_22779,N_22931);
and U23821 (N_23821,N_23576,N_23693);
nand U23822 (N_23822,N_22993,N_22505);
or U23823 (N_23823,N_23098,N_23078);
and U23824 (N_23824,N_23299,N_22560);
or U23825 (N_23825,N_22784,N_22549);
nor U23826 (N_23826,N_23582,N_23608);
xor U23827 (N_23827,N_22752,N_22842);
nand U23828 (N_23828,N_23485,N_23595);
xor U23829 (N_23829,N_23269,N_23617);
xnor U23830 (N_23830,N_23468,N_23414);
xor U23831 (N_23831,N_22740,N_23641);
xor U23832 (N_23832,N_23679,N_23189);
and U23833 (N_23833,N_22500,N_22579);
and U23834 (N_23834,N_22915,N_23668);
or U23835 (N_23835,N_22906,N_23441);
nand U23836 (N_23836,N_23523,N_22823);
and U23837 (N_23837,N_22844,N_23611);
nor U23838 (N_23838,N_22746,N_22644);
xor U23839 (N_23839,N_23389,N_22876);
or U23840 (N_23840,N_23251,N_23648);
and U23841 (N_23841,N_23352,N_22613);
and U23842 (N_23842,N_23570,N_23001);
or U23843 (N_23843,N_23540,N_22841);
nor U23844 (N_23844,N_22583,N_22608);
and U23845 (N_23845,N_23639,N_23651);
and U23846 (N_23846,N_22845,N_22798);
nor U23847 (N_23847,N_23255,N_22928);
nand U23848 (N_23848,N_23402,N_23091);
nand U23849 (N_23849,N_22641,N_23343);
xor U23850 (N_23850,N_23271,N_23211);
and U23851 (N_23851,N_23633,N_22974);
nor U23852 (N_23852,N_22822,N_23702);
or U23853 (N_23853,N_22821,N_22629);
xor U23854 (N_23854,N_22771,N_23499);
xnor U23855 (N_23855,N_23156,N_23227);
xnor U23856 (N_23856,N_23071,N_23416);
nor U23857 (N_23857,N_23135,N_23454);
nor U23858 (N_23858,N_22766,N_23554);
or U23859 (N_23859,N_22912,N_22683);
xor U23860 (N_23860,N_23504,N_22949);
nand U23861 (N_23861,N_22610,N_23423);
or U23862 (N_23862,N_23631,N_22741);
nand U23863 (N_23863,N_22634,N_23186);
xor U23864 (N_23864,N_22801,N_23121);
nor U23865 (N_23865,N_22824,N_23150);
nand U23866 (N_23866,N_23612,N_22728);
xor U23867 (N_23867,N_23486,N_23507);
xor U23868 (N_23868,N_23401,N_22692);
or U23869 (N_23869,N_22675,N_23006);
and U23870 (N_23870,N_23586,N_23293);
nand U23871 (N_23871,N_22696,N_23667);
xor U23872 (N_23872,N_22544,N_23566);
nor U23873 (N_23873,N_22980,N_22976);
and U23874 (N_23874,N_23603,N_22836);
or U23875 (N_23875,N_23248,N_22910);
xor U23876 (N_23876,N_22697,N_23747);
nor U23877 (N_23877,N_22878,N_22865);
nand U23878 (N_23878,N_23205,N_23577);
xnor U23879 (N_23879,N_22770,N_23239);
nand U23880 (N_23880,N_23119,N_23177);
xor U23881 (N_23881,N_23503,N_23398);
nor U23882 (N_23882,N_23174,N_23193);
nand U23883 (N_23883,N_22927,N_22867);
nor U23884 (N_23884,N_22554,N_23144);
and U23885 (N_23885,N_22742,N_23041);
nor U23886 (N_23886,N_23021,N_23562);
nor U23887 (N_23887,N_22888,N_23217);
or U23888 (N_23888,N_23490,N_23198);
nor U23889 (N_23889,N_23126,N_23601);
xor U23890 (N_23890,N_23115,N_22671);
or U23891 (N_23891,N_22884,N_22512);
xor U23892 (N_23892,N_22591,N_22636);
nor U23893 (N_23893,N_23060,N_22751);
and U23894 (N_23894,N_23708,N_23488);
nand U23895 (N_23895,N_22564,N_22744);
or U23896 (N_23896,N_22757,N_22902);
nor U23897 (N_23897,N_23072,N_23088);
xor U23898 (N_23898,N_22879,N_22627);
and U23899 (N_23899,N_23334,N_23043);
xnor U23900 (N_23900,N_22814,N_23388);
nand U23901 (N_23901,N_22945,N_22525);
and U23902 (N_23902,N_23729,N_23544);
nand U23903 (N_23903,N_23212,N_22938);
nand U23904 (N_23904,N_23404,N_23065);
nand U23905 (N_23905,N_23310,N_23457);
nand U23906 (N_23906,N_23319,N_23229);
nor U23907 (N_23907,N_23661,N_23359);
xor U23908 (N_23908,N_23709,N_23495);
or U23909 (N_23909,N_23378,N_22904);
and U23910 (N_23910,N_22611,N_23233);
xor U23911 (N_23911,N_22971,N_23700);
and U23912 (N_23912,N_22959,N_23433);
nand U23913 (N_23913,N_22578,N_23647);
xnor U23914 (N_23914,N_23068,N_23737);
nand U23915 (N_23915,N_22817,N_22605);
nand U23916 (N_23916,N_23369,N_23296);
or U23917 (N_23917,N_23335,N_23687);
or U23918 (N_23918,N_22656,N_23232);
nand U23919 (N_23919,N_22913,N_23536);
nor U23920 (N_23920,N_22556,N_22552);
xor U23921 (N_23921,N_23087,N_22767);
xnor U23922 (N_23922,N_23183,N_22620);
nor U23923 (N_23923,N_22970,N_22777);
nand U23924 (N_23924,N_23151,N_23120);
and U23925 (N_23925,N_22700,N_23460);
xnor U23926 (N_23926,N_23318,N_22690);
nor U23927 (N_23927,N_22940,N_23367);
or U23928 (N_23928,N_22640,N_23428);
xor U23929 (N_23929,N_22541,N_23011);
or U23930 (N_23930,N_23218,N_23430);
nand U23931 (N_23931,N_23305,N_22772);
xor U23932 (N_23932,N_22964,N_22890);
nand U23933 (N_23933,N_22599,N_23528);
and U23934 (N_23934,N_23128,N_23519);
nand U23935 (N_23935,N_23663,N_22750);
xor U23936 (N_23936,N_22606,N_23386);
or U23937 (N_23937,N_23331,N_23656);
or U23938 (N_23938,N_23598,N_23724);
nand U23939 (N_23939,N_22587,N_22828);
nand U23940 (N_23940,N_22586,N_23462);
or U23941 (N_23941,N_22725,N_23506);
nand U23942 (N_23942,N_23032,N_23132);
or U23943 (N_23943,N_23036,N_23525);
or U23944 (N_23944,N_23524,N_22705);
nand U23945 (N_23945,N_23345,N_23244);
nor U23946 (N_23946,N_23316,N_23671);
nor U23947 (N_23947,N_22914,N_23394);
xor U23948 (N_23948,N_22827,N_23408);
nand U23949 (N_23949,N_22911,N_22624);
nand U23950 (N_23950,N_23230,N_22901);
nand U23951 (N_23951,N_22569,N_23044);
and U23952 (N_23952,N_23253,N_23122);
and U23953 (N_23953,N_22684,N_23374);
and U23954 (N_23954,N_22559,N_23234);
nand U23955 (N_23955,N_23315,N_23583);
nand U23956 (N_23956,N_22753,N_23487);
nor U23957 (N_23957,N_22698,N_22601);
nor U23958 (N_23958,N_23215,N_22612);
xor U23959 (N_23959,N_22711,N_23199);
or U23960 (N_23960,N_23471,N_23246);
and U23961 (N_23961,N_23237,N_22943);
nor U23962 (N_23962,N_23497,N_23715);
nand U23963 (N_23963,N_22946,N_22905);
and U23964 (N_23964,N_23114,N_22639);
or U23965 (N_23965,N_23455,N_22524);
and U23966 (N_23966,N_22773,N_22693);
nor U23967 (N_23967,N_22619,N_23125);
or U23968 (N_23968,N_22942,N_22966);
nor U23969 (N_23969,N_23252,N_22745);
and U23970 (N_23970,N_23094,N_23442);
nor U23971 (N_23971,N_23739,N_23138);
nand U23972 (N_23972,N_22680,N_22618);
xnor U23973 (N_23973,N_23384,N_22666);
xnor U23974 (N_23974,N_22764,N_23734);
and U23975 (N_23975,N_23243,N_23161);
or U23976 (N_23976,N_22809,N_23621);
xnor U23977 (N_23977,N_23410,N_22602);
and U23978 (N_23978,N_23680,N_23339);
xnor U23979 (N_23979,N_23469,N_23084);
nor U23980 (N_23980,N_23713,N_23730);
nor U23981 (N_23981,N_23728,N_22628);
xor U23982 (N_23982,N_22584,N_22593);
nor U23983 (N_23983,N_23284,N_23531);
or U23984 (N_23984,N_23081,N_23623);
nand U23985 (N_23985,N_23015,N_23417);
nor U23986 (N_23986,N_23321,N_23511);
or U23987 (N_23987,N_23721,N_23675);
and U23988 (N_23988,N_23185,N_23159);
xor U23989 (N_23989,N_22655,N_23645);
nor U23990 (N_23990,N_23664,N_23019);
xor U23991 (N_23991,N_22858,N_22668);
nand U23992 (N_23992,N_22546,N_23385);
xnor U23993 (N_23993,N_23619,N_23741);
and U23994 (N_23994,N_22775,N_23250);
xor U23995 (N_23995,N_23659,N_23146);
xnor U23996 (N_23996,N_23090,N_23551);
nand U23997 (N_23997,N_23437,N_22820);
or U23998 (N_23998,N_23521,N_23446);
xor U23999 (N_23999,N_23192,N_23124);
and U24000 (N_24000,N_22871,N_23163);
or U24001 (N_24001,N_23558,N_23626);
xor U24002 (N_24002,N_23140,N_23373);
or U24003 (N_24003,N_23375,N_23644);
nand U24004 (N_24004,N_23592,N_22921);
nand U24005 (N_24005,N_23364,N_23200);
or U24006 (N_24006,N_22986,N_23075);
and U24007 (N_24007,N_23607,N_23396);
xnor U24008 (N_24008,N_23306,N_22955);
nand U24009 (N_24009,N_23154,N_23591);
nor U24010 (N_24010,N_22849,N_23033);
nand U24011 (N_24011,N_23048,N_23434);
or U24012 (N_24012,N_22625,N_23247);
nor U24013 (N_24013,N_23275,N_23658);
and U24014 (N_24014,N_23013,N_22632);
nor U24015 (N_24015,N_22839,N_22713);
xnor U24016 (N_24016,N_23482,N_23415);
nor U24017 (N_24017,N_23421,N_22536);
or U24018 (N_24018,N_23133,N_23445);
and U24019 (N_24019,N_22846,N_23743);
nor U24020 (N_24020,N_22778,N_23694);
or U24021 (N_24021,N_23061,N_22831);
nor U24022 (N_24022,N_23338,N_23684);
nand U24023 (N_24023,N_22851,N_23261);
or U24024 (N_24024,N_22794,N_22664);
xor U24025 (N_24025,N_23155,N_23093);
or U24026 (N_24026,N_23676,N_22689);
xor U24027 (N_24027,N_22535,N_23249);
nand U24028 (N_24028,N_23173,N_23701);
or U24029 (N_24029,N_23092,N_23660);
and U24030 (N_24030,N_22573,N_23311);
nand U24031 (N_24031,N_23387,N_23175);
or U24032 (N_24032,N_22835,N_22838);
nor U24033 (N_24033,N_23360,N_23476);
nor U24034 (N_24034,N_23555,N_22581);
or U24035 (N_24035,N_23240,N_23472);
nor U24036 (N_24036,N_22596,N_23587);
xnor U24037 (N_24037,N_23731,N_23014);
nand U24038 (N_24038,N_23265,N_23270);
or U24039 (N_24039,N_23543,N_23738);
and U24040 (N_24040,N_22607,N_23228);
xor U24041 (N_24041,N_22954,N_22894);
xnor U24042 (N_24042,N_22519,N_23662);
nor U24043 (N_24043,N_23560,N_23539);
or U24044 (N_24044,N_23298,N_23632);
and U24045 (N_24045,N_23597,N_23100);
nor U24046 (N_24046,N_23438,N_23111);
xnor U24047 (N_24047,N_22678,N_23039);
or U24048 (N_24048,N_23614,N_23363);
nor U24049 (N_24049,N_23357,N_23004);
and U24050 (N_24050,N_23031,N_23403);
xnor U24051 (N_24051,N_22513,N_23104);
nor U24052 (N_24052,N_23399,N_23030);
nor U24053 (N_24053,N_23066,N_23372);
and U24054 (N_24054,N_22534,N_23341);
nand U24055 (N_24055,N_22716,N_22896);
nand U24056 (N_24056,N_23337,N_22975);
nand U24057 (N_24057,N_23706,N_23083);
xor U24058 (N_24058,N_23085,N_22868);
nor U24059 (N_24059,N_22585,N_23353);
or U24060 (N_24060,N_23565,N_23447);
nand U24061 (N_24061,N_23431,N_23594);
and U24062 (N_24062,N_23720,N_23350);
xor U24063 (N_24063,N_22995,N_22999);
and U24064 (N_24064,N_23107,N_22590);
and U24065 (N_24065,N_23137,N_23262);
or U24066 (N_24066,N_22941,N_22568);
xor U24067 (N_24067,N_22595,N_23492);
nor U24068 (N_24068,N_23307,N_23049);
nor U24069 (N_24069,N_23281,N_22880);
xnor U24070 (N_24070,N_22977,N_23567);
nor U24071 (N_24071,N_22521,N_23038);
nand U24072 (N_24072,N_22681,N_23439);
xnor U24073 (N_24073,N_22501,N_23277);
and U24074 (N_24074,N_23725,N_23047);
nor U24075 (N_24075,N_22551,N_22670);
and U24076 (N_24076,N_22537,N_23392);
nor U24077 (N_24077,N_22708,N_23405);
xnor U24078 (N_24078,N_22704,N_23581);
and U24079 (N_24079,N_23593,N_22738);
nand U24080 (N_24080,N_22991,N_23470);
nand U24081 (N_24081,N_22807,N_22953);
nor U24082 (N_24082,N_23742,N_23530);
or U24083 (N_24083,N_23278,N_22866);
nand U24084 (N_24084,N_22870,N_23564);
xor U24085 (N_24085,N_22661,N_23297);
and U24086 (N_24086,N_23629,N_23527);
and U24087 (N_24087,N_23052,N_22756);
nand U24088 (N_24088,N_23697,N_22555);
nand U24089 (N_24089,N_23395,N_23452);
or U24090 (N_24090,N_23609,N_22957);
nand U24091 (N_24091,N_22998,N_22570);
nand U24092 (N_24092,N_22860,N_23178);
or U24093 (N_24093,N_23427,N_22787);
nor U24094 (N_24094,N_22789,N_23578);
nand U24095 (N_24095,N_23201,N_23326);
nand U24096 (N_24096,N_22774,N_22598);
nand U24097 (N_24097,N_23181,N_23303);
nand U24098 (N_24098,N_23196,N_22561);
and U24099 (N_24099,N_23346,N_22710);
xor U24100 (N_24100,N_22654,N_22686);
or U24101 (N_24101,N_22873,N_22968);
nor U24102 (N_24102,N_22859,N_23309);
or U24103 (N_24103,N_23134,N_23236);
and U24104 (N_24104,N_23444,N_23541);
xor U24105 (N_24105,N_23585,N_22735);
nand U24106 (N_24106,N_22754,N_22985);
xnor U24107 (N_24107,N_22930,N_23348);
nand U24108 (N_24108,N_23669,N_23145);
xnor U24109 (N_24109,N_23207,N_23020);
or U24110 (N_24110,N_22972,N_23710);
and U24111 (N_24111,N_22635,N_23187);
and U24112 (N_24112,N_22780,N_23569);
nor U24113 (N_24113,N_22783,N_23678);
nand U24114 (N_24114,N_23055,N_23618);
or U24115 (N_24115,N_22630,N_23361);
xnor U24116 (N_24116,N_23139,N_23493);
nor U24117 (N_24117,N_23025,N_22545);
or U24118 (N_24118,N_23699,N_23074);
or U24119 (N_24119,N_22651,N_22631);
xor U24120 (N_24120,N_23024,N_23195);
or U24121 (N_24121,N_22540,N_23086);
xnor U24122 (N_24122,N_23475,N_23282);
nor U24123 (N_24123,N_23131,N_22863);
nand U24124 (N_24124,N_23368,N_23096);
xor U24125 (N_24125,N_22803,N_23026);
and U24126 (N_24126,N_22615,N_22908);
or U24127 (N_24127,N_23008,N_22952);
and U24128 (N_24128,N_23448,N_22520);
nor U24129 (N_24129,N_22761,N_23257);
and U24130 (N_24130,N_23142,N_23172);
or U24131 (N_24131,N_22553,N_23443);
nor U24132 (N_24132,N_22933,N_23238);
and U24133 (N_24133,N_22724,N_23574);
nand U24134 (N_24134,N_23208,N_23391);
and U24135 (N_24135,N_23242,N_23322);
xor U24136 (N_24136,N_23657,N_23022);
xor U24137 (N_24137,N_22886,N_23285);
or U24138 (N_24138,N_23210,N_23102);
nand U24139 (N_24139,N_23589,N_23168);
and U24140 (N_24140,N_22808,N_23127);
or U24141 (N_24141,N_23740,N_23718);
and U24142 (N_24142,N_23624,N_23188);
or U24143 (N_24143,N_22588,N_23010);
nor U24144 (N_24144,N_23670,N_23029);
and U24145 (N_24145,N_22786,N_23007);
nor U24146 (N_24146,N_22633,N_22776);
or U24147 (N_24147,N_22717,N_22652);
xor U24148 (N_24148,N_23654,N_22748);
or U24149 (N_24149,N_22514,N_22543);
nand U24150 (N_24150,N_23615,N_23108);
and U24151 (N_24151,N_22643,N_22892);
nor U24152 (N_24152,N_23512,N_23620);
xnor U24153 (N_24153,N_22963,N_23067);
and U24154 (N_24154,N_23016,N_22855);
or U24155 (N_24155,N_22547,N_22785);
nor U24156 (N_24156,N_22760,N_22759);
nor U24157 (N_24157,N_23625,N_22617);
or U24158 (N_24158,N_23535,N_23516);
and U24159 (N_24159,N_22730,N_23736);
nor U24160 (N_24160,N_22694,N_23023);
nand U24161 (N_24161,N_23382,N_23484);
xnor U24162 (N_24162,N_23157,N_23241);
nor U24163 (N_24163,N_23748,N_23162);
and U24164 (N_24164,N_23143,N_23514);
or U24165 (N_24165,N_23064,N_23069);
nand U24166 (N_24166,N_23424,N_22687);
and U24167 (N_24167,N_22511,N_23561);
or U24168 (N_24168,N_22818,N_23079);
nor U24169 (N_24169,N_23508,N_23356);
and U24170 (N_24170,N_23202,N_23037);
xnor U24171 (N_24171,N_23695,N_23141);
and U24172 (N_24172,N_23688,N_22739);
or U24173 (N_24173,N_23590,N_23046);
nor U24174 (N_24174,N_22850,N_23354);
nor U24175 (N_24175,N_23638,N_22548);
nand U24176 (N_24176,N_22674,N_23510);
nor U24177 (N_24177,N_23409,N_23349);
xor U24178 (N_24178,N_23379,N_22934);
nor U24179 (N_24179,N_23563,N_22984);
and U24180 (N_24180,N_22988,N_23420);
and U24181 (N_24181,N_22982,N_23347);
and U24182 (N_24182,N_22538,N_23453);
and U24183 (N_24183,N_23522,N_22576);
xnor U24184 (N_24184,N_23179,N_23082);
xnor U24185 (N_24185,N_22609,N_22916);
nor U24186 (N_24186,N_22889,N_22557);
and U24187 (N_24187,N_23537,N_23666);
or U24188 (N_24188,N_22788,N_23426);
nor U24189 (N_24189,N_23149,N_23707);
and U24190 (N_24190,N_23190,N_23573);
xnor U24191 (N_24191,N_23459,N_23622);
or U24192 (N_24192,N_22669,N_23312);
nand U24193 (N_24193,N_23073,N_23324);
nand U24194 (N_24194,N_23606,N_22507);
nand U24195 (N_24195,N_22682,N_22826);
and U24196 (N_24196,N_23704,N_23456);
xnor U24197 (N_24197,N_23600,N_23571);
xnor U24198 (N_24198,N_22603,N_22990);
nand U24199 (N_24199,N_23628,N_23411);
nor U24200 (N_24200,N_22979,N_23095);
nor U24201 (N_24201,N_22582,N_22566);
xnor U24202 (N_24202,N_23216,N_22802);
and U24203 (N_24203,N_22506,N_22965);
xor U24204 (N_24204,N_23520,N_22800);
xor U24205 (N_24205,N_23529,N_22550);
xnor U24206 (N_24206,N_22718,N_23327);
xnor U24207 (N_24207,N_22909,N_22948);
nand U24208 (N_24208,N_22936,N_22685);
xor U24209 (N_24209,N_23498,N_22992);
nand U24210 (N_24210,N_22597,N_23027);
and U24211 (N_24211,N_22747,N_23501);
nand U24212 (N_24212,N_23148,N_22623);
xor U24213 (N_24213,N_22667,N_22811);
or U24214 (N_24214,N_23225,N_23342);
nand U24215 (N_24215,N_23376,N_23370);
xor U24216 (N_24216,N_22900,N_23605);
or U24217 (N_24217,N_23652,N_23276);
xnor U24218 (N_24218,N_23650,N_22869);
and U24219 (N_24219,N_22939,N_23330);
nor U24220 (N_24220,N_22580,N_22600);
and U24221 (N_24221,N_23076,N_23496);
nand U24222 (N_24222,N_22653,N_22994);
xor U24223 (N_24223,N_22649,N_22672);
nor U24224 (N_24224,N_22518,N_22659);
nor U24225 (N_24225,N_23494,N_23491);
or U24226 (N_24226,N_22920,N_23696);
nand U24227 (N_24227,N_23473,N_23272);
and U24228 (N_24228,N_22526,N_22791);
nor U24229 (N_24229,N_23118,N_23209);
xor U24230 (N_24230,N_22956,N_22962);
or U24231 (N_24231,N_22797,N_22523);
nand U24232 (N_24232,N_23451,N_23129);
nand U24233 (N_24233,N_23466,N_22837);
and U24234 (N_24234,N_23197,N_23509);
xnor U24235 (N_24235,N_23517,N_23170);
nand U24236 (N_24236,N_23532,N_23732);
nand U24237 (N_24237,N_23542,N_22804);
nor U24238 (N_24238,N_23735,N_23171);
nor U24239 (N_24239,N_23549,N_22950);
nand U24240 (N_24240,N_22530,N_22594);
xor U24241 (N_24241,N_23579,N_22567);
nor U24242 (N_24242,N_23333,N_23040);
and U24243 (N_24243,N_22897,N_22637);
xnor U24244 (N_24244,N_23634,N_22691);
or U24245 (N_24245,N_22558,N_23429);
nand U24246 (N_24246,N_22885,N_22877);
xnor U24247 (N_24247,N_23450,N_23406);
xor U24248 (N_24248,N_23325,N_23458);
nor U24249 (N_24249,N_23051,N_22528);
xnor U24250 (N_24250,N_23518,N_23547);
or U24251 (N_24251,N_23683,N_23604);
nand U24252 (N_24252,N_23393,N_22907);
nor U24253 (N_24253,N_22737,N_22935);
nor U24254 (N_24254,N_23099,N_22706);
or U24255 (N_24255,N_23245,N_23290);
xor U24256 (N_24256,N_22720,N_22562);
nor U24257 (N_24257,N_22947,N_23165);
nand U24258 (N_24258,N_22852,N_23054);
or U24259 (N_24259,N_22702,N_23655);
or U24260 (N_24260,N_22862,N_23077);
nand U24261 (N_24261,N_23635,N_23545);
and U24262 (N_24262,N_23464,N_23616);
and U24263 (N_24263,N_23176,N_22795);
or U24264 (N_24264,N_23674,N_22527);
nand U24265 (N_24265,N_23691,N_23314);
nor U24266 (N_24266,N_23714,N_23182);
nor U24267 (N_24267,N_22923,N_22577);
nor U24268 (N_24268,N_23381,N_22768);
xor U24269 (N_24269,N_23643,N_23112);
and U24270 (N_24270,N_23295,N_23419);
nor U24271 (N_24271,N_23184,N_23336);
xor U24272 (N_24272,N_22769,N_22951);
nor U24273 (N_24273,N_22614,N_22574);
nand U24274 (N_24274,N_22734,N_22709);
or U24275 (N_24275,N_22699,N_23588);
xnor U24276 (N_24276,N_23575,N_23113);
nand U24277 (N_24277,N_22522,N_22825);
or U24278 (N_24278,N_23400,N_23449);
and U24279 (N_24279,N_22542,N_22903);
and U24280 (N_24280,N_23062,N_23153);
or U24281 (N_24281,N_22857,N_22864);
xor U24282 (N_24282,N_22515,N_23572);
nor U24283 (N_24283,N_23692,N_23167);
or U24284 (N_24284,N_23513,N_22853);
or U24285 (N_24285,N_22819,N_23070);
nor U24286 (N_24286,N_22714,N_23028);
and U24287 (N_24287,N_22755,N_23012);
nor U24288 (N_24288,N_22658,N_23329);
xor U24289 (N_24289,N_22781,N_22882);
xor U24290 (N_24290,N_23705,N_22895);
nand U24291 (N_24291,N_23407,N_23649);
nand U24292 (N_24292,N_22925,N_22729);
and U24293 (N_24293,N_22723,N_22861);
nor U24294 (N_24294,N_23548,N_22650);
nand U24295 (N_24295,N_22765,N_23256);
nor U24296 (N_24296,N_23344,N_22926);
nor U24297 (N_24297,N_22622,N_23744);
or U24298 (N_24298,N_22799,N_22762);
and U24299 (N_24299,N_23425,N_23058);
xor U24300 (N_24300,N_22529,N_22840);
nor U24301 (N_24301,N_23500,N_23436);
nor U24302 (N_24302,N_23220,N_23553);
xnor U24303 (N_24303,N_23613,N_23097);
nor U24304 (N_24304,N_23313,N_23323);
and U24305 (N_24305,N_22987,N_23147);
nand U24306 (N_24306,N_22679,N_22830);
nand U24307 (N_24307,N_23677,N_22891);
xnor U24308 (N_24308,N_22924,N_22944);
and U24309 (N_24309,N_22510,N_23050);
nor U24310 (N_24310,N_23264,N_23489);
nand U24311 (N_24311,N_22688,N_23383);
or U24312 (N_24312,N_23063,N_23206);
nand U24313 (N_24313,N_23355,N_23231);
nor U24314 (N_24314,N_23749,N_23461);
or U24315 (N_24315,N_23733,N_23722);
and U24316 (N_24316,N_23550,N_23719);
nor U24317 (N_24317,N_22872,N_23105);
nand U24318 (N_24318,N_22657,N_22960);
xnor U24319 (N_24319,N_23042,N_23059);
nand U24320 (N_24320,N_22805,N_22848);
nand U24321 (N_24321,N_23502,N_23057);
and U24322 (N_24322,N_23283,N_23377);
and U24323 (N_24323,N_22782,N_23556);
nand U24324 (N_24324,N_23682,N_23358);
or U24325 (N_24325,N_22917,N_22978);
xor U24326 (N_24326,N_23727,N_23260);
nor U24327 (N_24327,N_23273,N_23018);
nor U24328 (N_24328,N_23362,N_22575);
or U24329 (N_24329,N_22918,N_23533);
and U24330 (N_24330,N_23017,N_23559);
xor U24331 (N_24331,N_23117,N_22969);
nand U24332 (N_24332,N_23467,N_23380);
nand U24333 (N_24333,N_23274,N_23328);
and U24334 (N_24334,N_23221,N_22646);
and U24335 (N_24335,N_22645,N_23505);
and U24336 (N_24336,N_23301,N_23089);
and U24337 (N_24337,N_23045,N_23194);
nand U24338 (N_24338,N_22642,N_22989);
nor U24339 (N_24339,N_23130,N_22648);
and U24340 (N_24340,N_23580,N_23584);
xor U24341 (N_24341,N_22792,N_23340);
xor U24342 (N_24342,N_23365,N_23534);
nor U24343 (N_24343,N_23300,N_23745);
xor U24344 (N_24344,N_22626,N_23288);
nand U24345 (N_24345,N_22856,N_23599);
and U24346 (N_24346,N_22832,N_23432);
nor U24347 (N_24347,N_23552,N_23332);
nor U24348 (N_24348,N_23465,N_23080);
and U24349 (N_24349,N_23716,N_22983);
nor U24350 (N_24350,N_23302,N_23703);
nand U24351 (N_24351,N_23711,N_22919);
nor U24352 (N_24352,N_22722,N_23390);
nor U24353 (N_24353,N_22509,N_23224);
or U24354 (N_24354,N_23263,N_23435);
nand U24355 (N_24355,N_23191,N_23723);
xor U24356 (N_24356,N_22981,N_22712);
nand U24357 (N_24357,N_23223,N_23685);
xor U24358 (N_24358,N_22875,N_22834);
nor U24359 (N_24359,N_23109,N_23712);
or U24360 (N_24360,N_22932,N_22508);
xor U24361 (N_24361,N_23478,N_22967);
nand U24362 (N_24362,N_23289,N_22736);
nor U24363 (N_24363,N_23204,N_23627);
and U24364 (N_24364,N_23136,N_23538);
and U24365 (N_24365,N_23000,N_22715);
and U24366 (N_24366,N_23268,N_23479);
and U24367 (N_24367,N_22847,N_22790);
and U24368 (N_24368,N_22616,N_22589);
nand U24369 (N_24369,N_22703,N_23557);
nor U24370 (N_24370,N_22502,N_22621);
nand U24371 (N_24371,N_22563,N_23630);
or U24372 (N_24372,N_23180,N_23164);
xor U24373 (N_24373,N_22887,N_22707);
or U24374 (N_24374,N_23717,N_23035);
and U24375 (N_24375,N_22833,N_22629);
and U24376 (N_24376,N_22556,N_23149);
xnor U24377 (N_24377,N_23456,N_23030);
and U24378 (N_24378,N_22917,N_22775);
nand U24379 (N_24379,N_23737,N_23439);
xor U24380 (N_24380,N_22561,N_23564);
nor U24381 (N_24381,N_22972,N_22790);
nand U24382 (N_24382,N_23506,N_22898);
and U24383 (N_24383,N_22879,N_22890);
nor U24384 (N_24384,N_23444,N_22915);
nor U24385 (N_24385,N_22671,N_23448);
nor U24386 (N_24386,N_22851,N_23139);
or U24387 (N_24387,N_23335,N_22772);
nand U24388 (N_24388,N_23343,N_23450);
nor U24389 (N_24389,N_23739,N_23309);
xor U24390 (N_24390,N_23298,N_23499);
nor U24391 (N_24391,N_22835,N_23430);
xnor U24392 (N_24392,N_23422,N_22599);
xor U24393 (N_24393,N_23415,N_23540);
nor U24394 (N_24394,N_23423,N_23005);
or U24395 (N_24395,N_22985,N_23187);
xnor U24396 (N_24396,N_22630,N_23397);
nand U24397 (N_24397,N_22907,N_23040);
nor U24398 (N_24398,N_23337,N_22552);
xnor U24399 (N_24399,N_22872,N_23668);
xnor U24400 (N_24400,N_22660,N_23177);
nand U24401 (N_24401,N_23625,N_23267);
and U24402 (N_24402,N_23262,N_22540);
or U24403 (N_24403,N_23497,N_22774);
nand U24404 (N_24404,N_22800,N_23072);
nand U24405 (N_24405,N_23672,N_22791);
xor U24406 (N_24406,N_22645,N_23353);
or U24407 (N_24407,N_23303,N_23329);
or U24408 (N_24408,N_23740,N_22512);
and U24409 (N_24409,N_22899,N_23189);
nand U24410 (N_24410,N_23699,N_23463);
nor U24411 (N_24411,N_22648,N_23710);
nand U24412 (N_24412,N_22649,N_22968);
and U24413 (N_24413,N_23632,N_22737);
nand U24414 (N_24414,N_22844,N_23271);
and U24415 (N_24415,N_22868,N_23563);
nor U24416 (N_24416,N_23649,N_23503);
xnor U24417 (N_24417,N_22523,N_23232);
and U24418 (N_24418,N_23188,N_23088);
or U24419 (N_24419,N_23677,N_22961);
nand U24420 (N_24420,N_23521,N_23612);
nand U24421 (N_24421,N_23472,N_23545);
nand U24422 (N_24422,N_23510,N_23073);
nor U24423 (N_24423,N_23154,N_23414);
and U24424 (N_24424,N_23734,N_23475);
xnor U24425 (N_24425,N_23582,N_22647);
or U24426 (N_24426,N_23299,N_23698);
nor U24427 (N_24427,N_23304,N_23749);
xnor U24428 (N_24428,N_23414,N_23192);
and U24429 (N_24429,N_23243,N_22610);
or U24430 (N_24430,N_23110,N_23452);
nor U24431 (N_24431,N_23575,N_23309);
nand U24432 (N_24432,N_23191,N_23673);
nand U24433 (N_24433,N_23695,N_23498);
nor U24434 (N_24434,N_23114,N_23205);
nand U24435 (N_24435,N_22827,N_23364);
nor U24436 (N_24436,N_22538,N_22961);
and U24437 (N_24437,N_23003,N_22523);
nor U24438 (N_24438,N_23387,N_22994);
and U24439 (N_24439,N_23437,N_23155);
nor U24440 (N_24440,N_23688,N_23723);
or U24441 (N_24441,N_22814,N_23318);
or U24442 (N_24442,N_23096,N_23744);
nor U24443 (N_24443,N_23236,N_22819);
or U24444 (N_24444,N_22563,N_22902);
and U24445 (N_24445,N_22929,N_22876);
and U24446 (N_24446,N_23119,N_22553);
nor U24447 (N_24447,N_23431,N_23157);
xor U24448 (N_24448,N_22729,N_23685);
nand U24449 (N_24449,N_22597,N_22633);
and U24450 (N_24450,N_22710,N_23719);
xnor U24451 (N_24451,N_23171,N_23550);
xor U24452 (N_24452,N_23597,N_22793);
xor U24453 (N_24453,N_23577,N_22656);
nand U24454 (N_24454,N_23213,N_23375);
nor U24455 (N_24455,N_23327,N_23223);
nor U24456 (N_24456,N_23671,N_22540);
xor U24457 (N_24457,N_23542,N_22505);
nor U24458 (N_24458,N_22772,N_23685);
nand U24459 (N_24459,N_23029,N_22900);
nand U24460 (N_24460,N_23213,N_23668);
nand U24461 (N_24461,N_22652,N_23419);
xor U24462 (N_24462,N_23240,N_22824);
nand U24463 (N_24463,N_23410,N_22641);
nand U24464 (N_24464,N_22821,N_22800);
nor U24465 (N_24465,N_22996,N_23610);
xor U24466 (N_24466,N_22513,N_22858);
and U24467 (N_24467,N_22803,N_23219);
nor U24468 (N_24468,N_23469,N_23161);
nand U24469 (N_24469,N_23354,N_23225);
nor U24470 (N_24470,N_22740,N_22868);
nor U24471 (N_24471,N_23301,N_22992);
or U24472 (N_24472,N_23373,N_22702);
xor U24473 (N_24473,N_22527,N_22805);
xnor U24474 (N_24474,N_22918,N_23463);
nand U24475 (N_24475,N_22969,N_23703);
nor U24476 (N_24476,N_22911,N_22716);
or U24477 (N_24477,N_23727,N_22852);
xor U24478 (N_24478,N_22960,N_22990);
nand U24479 (N_24479,N_23088,N_23116);
and U24480 (N_24480,N_23337,N_22743);
nand U24481 (N_24481,N_22895,N_23312);
nand U24482 (N_24482,N_22692,N_22663);
and U24483 (N_24483,N_23191,N_23294);
or U24484 (N_24484,N_22652,N_23286);
and U24485 (N_24485,N_23132,N_23271);
nand U24486 (N_24486,N_22651,N_23473);
xor U24487 (N_24487,N_22513,N_22533);
nor U24488 (N_24488,N_22505,N_23072);
xor U24489 (N_24489,N_23295,N_23377);
or U24490 (N_24490,N_23053,N_23394);
or U24491 (N_24491,N_22982,N_22792);
or U24492 (N_24492,N_23676,N_22700);
and U24493 (N_24493,N_22622,N_22982);
xnor U24494 (N_24494,N_22613,N_22659);
and U24495 (N_24495,N_22893,N_23668);
or U24496 (N_24496,N_23728,N_23055);
xnor U24497 (N_24497,N_22601,N_22897);
nand U24498 (N_24498,N_23041,N_23309);
nand U24499 (N_24499,N_23310,N_23728);
nor U24500 (N_24500,N_22793,N_23247);
nor U24501 (N_24501,N_23126,N_23559);
nand U24502 (N_24502,N_23628,N_22598);
xnor U24503 (N_24503,N_23188,N_22898);
nor U24504 (N_24504,N_22964,N_23082);
nand U24505 (N_24505,N_22848,N_22984);
xor U24506 (N_24506,N_22998,N_23708);
nand U24507 (N_24507,N_22715,N_23351);
or U24508 (N_24508,N_22626,N_23291);
or U24509 (N_24509,N_23097,N_23168);
or U24510 (N_24510,N_22932,N_23004);
or U24511 (N_24511,N_23114,N_23282);
nand U24512 (N_24512,N_23540,N_22693);
or U24513 (N_24513,N_22564,N_22887);
xnor U24514 (N_24514,N_23281,N_23710);
xnor U24515 (N_24515,N_22773,N_23412);
nand U24516 (N_24516,N_22830,N_22971);
or U24517 (N_24517,N_23300,N_23739);
or U24518 (N_24518,N_22522,N_22919);
xor U24519 (N_24519,N_23689,N_23037);
nor U24520 (N_24520,N_23188,N_23496);
xor U24521 (N_24521,N_23552,N_23212);
nor U24522 (N_24522,N_23479,N_22668);
xor U24523 (N_24523,N_23123,N_22772);
xor U24524 (N_24524,N_22587,N_23465);
or U24525 (N_24525,N_23240,N_22527);
nor U24526 (N_24526,N_22818,N_22663);
or U24527 (N_24527,N_22528,N_23531);
and U24528 (N_24528,N_22879,N_22587);
or U24529 (N_24529,N_22551,N_23566);
xnor U24530 (N_24530,N_23420,N_23026);
or U24531 (N_24531,N_23278,N_22585);
nand U24532 (N_24532,N_22809,N_23292);
xor U24533 (N_24533,N_22621,N_23189);
and U24534 (N_24534,N_23082,N_22812);
nor U24535 (N_24535,N_23254,N_22578);
nor U24536 (N_24536,N_23621,N_23078);
xnor U24537 (N_24537,N_22883,N_23415);
nor U24538 (N_24538,N_22820,N_23108);
nand U24539 (N_24539,N_22975,N_23492);
nand U24540 (N_24540,N_23019,N_23117);
and U24541 (N_24541,N_23047,N_23606);
nand U24542 (N_24542,N_22614,N_22934);
xnor U24543 (N_24543,N_23091,N_22550);
xor U24544 (N_24544,N_22503,N_22924);
or U24545 (N_24545,N_23597,N_23296);
or U24546 (N_24546,N_23279,N_23110);
xnor U24547 (N_24547,N_22884,N_23344);
and U24548 (N_24548,N_23367,N_22546);
and U24549 (N_24549,N_23339,N_23069);
nand U24550 (N_24550,N_23253,N_23028);
xnor U24551 (N_24551,N_23446,N_22814);
and U24552 (N_24552,N_22718,N_23657);
or U24553 (N_24553,N_23024,N_22735);
nand U24554 (N_24554,N_23130,N_22548);
xor U24555 (N_24555,N_23143,N_22573);
nand U24556 (N_24556,N_23125,N_22600);
nor U24557 (N_24557,N_22962,N_23614);
or U24558 (N_24558,N_22710,N_22735);
nand U24559 (N_24559,N_23489,N_23637);
nand U24560 (N_24560,N_23132,N_22898);
xnor U24561 (N_24561,N_22766,N_23699);
and U24562 (N_24562,N_23747,N_23602);
nor U24563 (N_24563,N_22855,N_23241);
nand U24564 (N_24564,N_23330,N_23495);
nand U24565 (N_24565,N_23239,N_23520);
nor U24566 (N_24566,N_22891,N_23307);
or U24567 (N_24567,N_22728,N_22851);
xnor U24568 (N_24568,N_23524,N_23018);
or U24569 (N_24569,N_22884,N_22870);
nor U24570 (N_24570,N_23729,N_23508);
or U24571 (N_24571,N_23069,N_23514);
or U24572 (N_24572,N_23075,N_23375);
nand U24573 (N_24573,N_23362,N_23501);
and U24574 (N_24574,N_23280,N_23635);
nand U24575 (N_24575,N_23539,N_23477);
nor U24576 (N_24576,N_22921,N_22537);
and U24577 (N_24577,N_22563,N_22696);
nor U24578 (N_24578,N_22943,N_22863);
nor U24579 (N_24579,N_23060,N_22684);
nor U24580 (N_24580,N_23300,N_23504);
nand U24581 (N_24581,N_22781,N_23589);
and U24582 (N_24582,N_23409,N_23703);
xor U24583 (N_24583,N_23535,N_22727);
or U24584 (N_24584,N_23319,N_23584);
or U24585 (N_24585,N_23029,N_23235);
or U24586 (N_24586,N_23562,N_23101);
and U24587 (N_24587,N_23305,N_23159);
nand U24588 (N_24588,N_23103,N_23712);
xor U24589 (N_24589,N_22660,N_22996);
nor U24590 (N_24590,N_23031,N_23237);
nand U24591 (N_24591,N_23393,N_23592);
nand U24592 (N_24592,N_22792,N_23187);
nand U24593 (N_24593,N_23668,N_22793);
or U24594 (N_24594,N_23267,N_23116);
nand U24595 (N_24595,N_22521,N_23155);
nor U24596 (N_24596,N_23672,N_22975);
nand U24597 (N_24597,N_22513,N_22742);
nand U24598 (N_24598,N_23507,N_23624);
or U24599 (N_24599,N_23547,N_22940);
xor U24600 (N_24600,N_22638,N_23503);
nor U24601 (N_24601,N_23451,N_23283);
nand U24602 (N_24602,N_23236,N_23397);
xor U24603 (N_24603,N_23293,N_23571);
or U24604 (N_24604,N_22629,N_23102);
xor U24605 (N_24605,N_23536,N_22663);
or U24606 (N_24606,N_22791,N_23500);
and U24607 (N_24607,N_23567,N_23127);
or U24608 (N_24608,N_22684,N_22754);
nand U24609 (N_24609,N_23660,N_23119);
nor U24610 (N_24610,N_23180,N_23053);
nor U24611 (N_24611,N_22624,N_23188);
xnor U24612 (N_24612,N_23463,N_23038);
nand U24613 (N_24613,N_22530,N_22821);
or U24614 (N_24614,N_22793,N_22909);
or U24615 (N_24615,N_23296,N_22938);
and U24616 (N_24616,N_23099,N_22596);
and U24617 (N_24617,N_23723,N_23628);
xor U24618 (N_24618,N_23441,N_22890);
xnor U24619 (N_24619,N_23355,N_22813);
nor U24620 (N_24620,N_23690,N_23011);
and U24621 (N_24621,N_23707,N_22654);
nor U24622 (N_24622,N_23176,N_23698);
nor U24623 (N_24623,N_23526,N_22718);
or U24624 (N_24624,N_23154,N_22975);
nor U24625 (N_24625,N_22819,N_22871);
and U24626 (N_24626,N_23413,N_22504);
or U24627 (N_24627,N_22779,N_23248);
xor U24628 (N_24628,N_22629,N_22633);
nor U24629 (N_24629,N_23012,N_23532);
xor U24630 (N_24630,N_23328,N_23165);
nand U24631 (N_24631,N_23659,N_22735);
nor U24632 (N_24632,N_23019,N_23342);
nor U24633 (N_24633,N_23250,N_23580);
nand U24634 (N_24634,N_23589,N_23637);
nor U24635 (N_24635,N_23730,N_23620);
nor U24636 (N_24636,N_23205,N_22553);
xor U24637 (N_24637,N_23595,N_23725);
nor U24638 (N_24638,N_23568,N_22692);
and U24639 (N_24639,N_22896,N_22676);
xor U24640 (N_24640,N_23228,N_23417);
nand U24641 (N_24641,N_22795,N_23667);
xor U24642 (N_24642,N_23117,N_22513);
or U24643 (N_24643,N_23632,N_22633);
nor U24644 (N_24644,N_23471,N_22720);
xnor U24645 (N_24645,N_22500,N_23700);
xor U24646 (N_24646,N_22531,N_23382);
and U24647 (N_24647,N_23723,N_23471);
nor U24648 (N_24648,N_23314,N_22649);
nor U24649 (N_24649,N_23438,N_23626);
nor U24650 (N_24650,N_23221,N_22871);
or U24651 (N_24651,N_23645,N_22872);
and U24652 (N_24652,N_23498,N_23664);
nor U24653 (N_24653,N_22667,N_22722);
nor U24654 (N_24654,N_23279,N_23641);
nor U24655 (N_24655,N_23010,N_22615);
nor U24656 (N_24656,N_22742,N_23393);
xor U24657 (N_24657,N_23591,N_23603);
nand U24658 (N_24658,N_23215,N_22600);
nor U24659 (N_24659,N_23664,N_23334);
and U24660 (N_24660,N_23095,N_23136);
or U24661 (N_24661,N_22854,N_22606);
nand U24662 (N_24662,N_22836,N_23073);
nor U24663 (N_24663,N_23055,N_23027);
or U24664 (N_24664,N_22953,N_23159);
or U24665 (N_24665,N_23071,N_23349);
or U24666 (N_24666,N_22935,N_23289);
nor U24667 (N_24667,N_23610,N_23387);
nor U24668 (N_24668,N_23020,N_23496);
or U24669 (N_24669,N_23084,N_23696);
and U24670 (N_24670,N_23035,N_22913);
nand U24671 (N_24671,N_23368,N_22818);
xnor U24672 (N_24672,N_23163,N_23287);
nor U24673 (N_24673,N_22924,N_23105);
and U24674 (N_24674,N_23465,N_23536);
nor U24675 (N_24675,N_22941,N_23651);
nor U24676 (N_24676,N_23583,N_23685);
nor U24677 (N_24677,N_23372,N_23385);
nor U24678 (N_24678,N_22811,N_23315);
nor U24679 (N_24679,N_22644,N_22558);
and U24680 (N_24680,N_23131,N_22664);
or U24681 (N_24681,N_23206,N_22628);
nor U24682 (N_24682,N_22588,N_23637);
and U24683 (N_24683,N_23392,N_22531);
or U24684 (N_24684,N_23279,N_23288);
or U24685 (N_24685,N_22749,N_23407);
xnor U24686 (N_24686,N_23256,N_23674);
or U24687 (N_24687,N_23634,N_22782);
xnor U24688 (N_24688,N_22712,N_23696);
xnor U24689 (N_24689,N_23080,N_23316);
or U24690 (N_24690,N_23728,N_23513);
and U24691 (N_24691,N_23222,N_22683);
xor U24692 (N_24692,N_23171,N_23566);
or U24693 (N_24693,N_22689,N_22523);
xnor U24694 (N_24694,N_22819,N_22634);
xnor U24695 (N_24695,N_22503,N_22651);
xnor U24696 (N_24696,N_23679,N_23076);
nor U24697 (N_24697,N_22842,N_23422);
nor U24698 (N_24698,N_23135,N_22715);
nor U24699 (N_24699,N_22803,N_22511);
xnor U24700 (N_24700,N_23506,N_22926);
or U24701 (N_24701,N_22700,N_22778);
and U24702 (N_24702,N_23732,N_23232);
nor U24703 (N_24703,N_23461,N_23123);
nand U24704 (N_24704,N_22918,N_23023);
xnor U24705 (N_24705,N_23690,N_22734);
and U24706 (N_24706,N_23402,N_23185);
and U24707 (N_24707,N_22636,N_22814);
or U24708 (N_24708,N_23660,N_23685);
nor U24709 (N_24709,N_23450,N_22778);
xnor U24710 (N_24710,N_23335,N_22756);
or U24711 (N_24711,N_23490,N_23650);
or U24712 (N_24712,N_22882,N_23099);
nand U24713 (N_24713,N_22806,N_23173);
nand U24714 (N_24714,N_22918,N_22978);
or U24715 (N_24715,N_23098,N_23248);
or U24716 (N_24716,N_23128,N_22862);
and U24717 (N_24717,N_23064,N_23382);
nand U24718 (N_24718,N_22703,N_23209);
and U24719 (N_24719,N_23456,N_22519);
and U24720 (N_24720,N_23465,N_23141);
nand U24721 (N_24721,N_23524,N_23740);
xnor U24722 (N_24722,N_23715,N_23348);
or U24723 (N_24723,N_23492,N_22984);
nor U24724 (N_24724,N_23266,N_22504);
xor U24725 (N_24725,N_23381,N_22782);
xor U24726 (N_24726,N_23015,N_23687);
or U24727 (N_24727,N_23354,N_23305);
nand U24728 (N_24728,N_23551,N_22588);
nor U24729 (N_24729,N_22647,N_22523);
xnor U24730 (N_24730,N_23148,N_22527);
or U24731 (N_24731,N_23698,N_23126);
and U24732 (N_24732,N_22654,N_23487);
nand U24733 (N_24733,N_23510,N_22530);
xor U24734 (N_24734,N_23064,N_23117);
nor U24735 (N_24735,N_22990,N_22764);
or U24736 (N_24736,N_23368,N_23105);
nor U24737 (N_24737,N_23371,N_22663);
nand U24738 (N_24738,N_23192,N_23170);
xnor U24739 (N_24739,N_23411,N_23179);
nor U24740 (N_24740,N_23372,N_22652);
xnor U24741 (N_24741,N_23499,N_22778);
or U24742 (N_24742,N_22590,N_22605);
or U24743 (N_24743,N_23567,N_22825);
nor U24744 (N_24744,N_23230,N_23632);
and U24745 (N_24745,N_23317,N_23044);
and U24746 (N_24746,N_23596,N_23637);
xnor U24747 (N_24747,N_23298,N_23713);
nand U24748 (N_24748,N_22522,N_22713);
nor U24749 (N_24749,N_22842,N_22836);
xor U24750 (N_24750,N_23380,N_23029);
xor U24751 (N_24751,N_23362,N_23518);
and U24752 (N_24752,N_22878,N_22735);
nor U24753 (N_24753,N_23461,N_23246);
nand U24754 (N_24754,N_23043,N_23635);
nor U24755 (N_24755,N_22792,N_22655);
nand U24756 (N_24756,N_23030,N_23700);
nor U24757 (N_24757,N_23555,N_23582);
nor U24758 (N_24758,N_22727,N_23401);
xor U24759 (N_24759,N_23733,N_23055);
nand U24760 (N_24760,N_23354,N_23069);
and U24761 (N_24761,N_23105,N_23366);
nor U24762 (N_24762,N_22630,N_23305);
nor U24763 (N_24763,N_23494,N_23184);
nor U24764 (N_24764,N_22967,N_22730);
nor U24765 (N_24765,N_22820,N_23196);
or U24766 (N_24766,N_22707,N_22689);
nor U24767 (N_24767,N_22930,N_23539);
nand U24768 (N_24768,N_22707,N_23732);
and U24769 (N_24769,N_22994,N_22706);
or U24770 (N_24770,N_23452,N_23081);
nand U24771 (N_24771,N_23177,N_22941);
and U24772 (N_24772,N_23099,N_23175);
nor U24773 (N_24773,N_22629,N_23531);
nand U24774 (N_24774,N_22639,N_23416);
and U24775 (N_24775,N_23135,N_23167);
or U24776 (N_24776,N_23138,N_23182);
xor U24777 (N_24777,N_22844,N_23176);
or U24778 (N_24778,N_23527,N_22911);
nand U24779 (N_24779,N_23184,N_23206);
xor U24780 (N_24780,N_22960,N_23048);
or U24781 (N_24781,N_22713,N_22810);
nand U24782 (N_24782,N_22610,N_23501);
or U24783 (N_24783,N_23468,N_22683);
nor U24784 (N_24784,N_23347,N_23568);
nand U24785 (N_24785,N_23644,N_23249);
nor U24786 (N_24786,N_23277,N_22689);
and U24787 (N_24787,N_22924,N_23710);
nand U24788 (N_24788,N_23260,N_23069);
xor U24789 (N_24789,N_23742,N_23585);
xnor U24790 (N_24790,N_23204,N_23360);
nand U24791 (N_24791,N_22941,N_23243);
nor U24792 (N_24792,N_22894,N_22614);
xor U24793 (N_24793,N_23390,N_23582);
nor U24794 (N_24794,N_22762,N_23543);
nor U24795 (N_24795,N_23522,N_23385);
nor U24796 (N_24796,N_22934,N_23400);
or U24797 (N_24797,N_23326,N_23286);
nand U24798 (N_24798,N_22526,N_22996);
and U24799 (N_24799,N_22841,N_22709);
nand U24800 (N_24800,N_22576,N_22832);
xor U24801 (N_24801,N_23055,N_22650);
or U24802 (N_24802,N_23076,N_22737);
xor U24803 (N_24803,N_22657,N_23571);
xnor U24804 (N_24804,N_23700,N_22519);
nand U24805 (N_24805,N_23025,N_22876);
or U24806 (N_24806,N_22984,N_22636);
xor U24807 (N_24807,N_22840,N_23127);
nor U24808 (N_24808,N_23385,N_23640);
xnor U24809 (N_24809,N_22684,N_23483);
and U24810 (N_24810,N_23746,N_22801);
and U24811 (N_24811,N_23038,N_23715);
and U24812 (N_24812,N_22971,N_22531);
nand U24813 (N_24813,N_22973,N_22673);
and U24814 (N_24814,N_22799,N_23636);
and U24815 (N_24815,N_23743,N_22670);
nor U24816 (N_24816,N_22873,N_23656);
nand U24817 (N_24817,N_23039,N_23570);
or U24818 (N_24818,N_23215,N_23482);
or U24819 (N_24819,N_22842,N_23106);
or U24820 (N_24820,N_23598,N_23268);
and U24821 (N_24821,N_22969,N_22942);
or U24822 (N_24822,N_23659,N_23398);
nand U24823 (N_24823,N_22848,N_23673);
and U24824 (N_24824,N_23043,N_22978);
and U24825 (N_24825,N_22508,N_23096);
or U24826 (N_24826,N_22751,N_23582);
xnor U24827 (N_24827,N_23732,N_22812);
xor U24828 (N_24828,N_22905,N_23403);
nor U24829 (N_24829,N_23474,N_22527);
or U24830 (N_24830,N_23726,N_23382);
xnor U24831 (N_24831,N_22981,N_23736);
or U24832 (N_24832,N_22696,N_22791);
xor U24833 (N_24833,N_22520,N_23649);
and U24834 (N_24834,N_22587,N_22727);
nand U24835 (N_24835,N_23687,N_23432);
xnor U24836 (N_24836,N_23250,N_22637);
xnor U24837 (N_24837,N_22517,N_23688);
nor U24838 (N_24838,N_23333,N_23089);
or U24839 (N_24839,N_22547,N_22686);
and U24840 (N_24840,N_22989,N_22681);
nand U24841 (N_24841,N_23043,N_22660);
and U24842 (N_24842,N_23321,N_23133);
or U24843 (N_24843,N_22537,N_22508);
and U24844 (N_24844,N_23388,N_22674);
or U24845 (N_24845,N_23206,N_22599);
and U24846 (N_24846,N_23216,N_22998);
nand U24847 (N_24847,N_23212,N_22726);
nor U24848 (N_24848,N_22775,N_23433);
xor U24849 (N_24849,N_22817,N_23323);
and U24850 (N_24850,N_22682,N_23473);
and U24851 (N_24851,N_23089,N_22881);
nor U24852 (N_24852,N_23076,N_22708);
xnor U24853 (N_24853,N_23345,N_23185);
or U24854 (N_24854,N_23383,N_22866);
or U24855 (N_24855,N_22605,N_23660);
nand U24856 (N_24856,N_22941,N_23283);
xnor U24857 (N_24857,N_22925,N_22619);
and U24858 (N_24858,N_23628,N_23527);
and U24859 (N_24859,N_22987,N_23134);
xor U24860 (N_24860,N_23046,N_22615);
and U24861 (N_24861,N_23598,N_23539);
xor U24862 (N_24862,N_23419,N_23726);
and U24863 (N_24863,N_23372,N_23685);
nor U24864 (N_24864,N_23517,N_22638);
nor U24865 (N_24865,N_22739,N_22666);
xnor U24866 (N_24866,N_23426,N_23386);
xor U24867 (N_24867,N_22872,N_22611);
and U24868 (N_24868,N_22568,N_22811);
nand U24869 (N_24869,N_22899,N_22539);
xnor U24870 (N_24870,N_23466,N_23459);
or U24871 (N_24871,N_23161,N_22587);
or U24872 (N_24872,N_23094,N_23692);
or U24873 (N_24873,N_22698,N_23334);
or U24874 (N_24874,N_22861,N_22914);
and U24875 (N_24875,N_22516,N_23729);
nor U24876 (N_24876,N_22763,N_23113);
and U24877 (N_24877,N_23322,N_22520);
or U24878 (N_24878,N_23091,N_22554);
xor U24879 (N_24879,N_22803,N_23699);
nand U24880 (N_24880,N_22713,N_23531);
and U24881 (N_24881,N_22589,N_23228);
nor U24882 (N_24882,N_22900,N_22549);
nand U24883 (N_24883,N_22627,N_22812);
nor U24884 (N_24884,N_23491,N_23376);
or U24885 (N_24885,N_22747,N_22908);
or U24886 (N_24886,N_23481,N_22648);
xor U24887 (N_24887,N_23254,N_23057);
and U24888 (N_24888,N_22522,N_23558);
nand U24889 (N_24889,N_22506,N_22713);
or U24890 (N_24890,N_23114,N_23300);
nand U24891 (N_24891,N_23454,N_22580);
or U24892 (N_24892,N_23749,N_23131);
and U24893 (N_24893,N_22779,N_22718);
xnor U24894 (N_24894,N_22559,N_22627);
and U24895 (N_24895,N_23688,N_23236);
xor U24896 (N_24896,N_22952,N_22529);
or U24897 (N_24897,N_23454,N_22765);
nand U24898 (N_24898,N_23103,N_23420);
or U24899 (N_24899,N_22676,N_22877);
or U24900 (N_24900,N_22611,N_22886);
and U24901 (N_24901,N_23377,N_23276);
xor U24902 (N_24902,N_23138,N_23674);
or U24903 (N_24903,N_23384,N_22891);
nor U24904 (N_24904,N_22887,N_22796);
xor U24905 (N_24905,N_23079,N_22642);
nor U24906 (N_24906,N_22776,N_22877);
xor U24907 (N_24907,N_22896,N_22909);
or U24908 (N_24908,N_23007,N_22874);
or U24909 (N_24909,N_22556,N_23523);
nor U24910 (N_24910,N_23292,N_23607);
nor U24911 (N_24911,N_22751,N_23643);
xor U24912 (N_24912,N_23072,N_23015);
nor U24913 (N_24913,N_23184,N_22741);
nor U24914 (N_24914,N_22649,N_23214);
and U24915 (N_24915,N_23409,N_22948);
xor U24916 (N_24916,N_23569,N_22693);
and U24917 (N_24917,N_23373,N_23141);
and U24918 (N_24918,N_22660,N_23264);
nor U24919 (N_24919,N_23660,N_23087);
xnor U24920 (N_24920,N_23385,N_23195);
xor U24921 (N_24921,N_22609,N_22515);
nand U24922 (N_24922,N_22699,N_22628);
nor U24923 (N_24923,N_22711,N_23420);
xnor U24924 (N_24924,N_22528,N_23345);
and U24925 (N_24925,N_23037,N_23036);
or U24926 (N_24926,N_23215,N_23096);
xor U24927 (N_24927,N_22927,N_23527);
and U24928 (N_24928,N_22949,N_22533);
and U24929 (N_24929,N_22558,N_23462);
nand U24930 (N_24930,N_22785,N_22880);
nand U24931 (N_24931,N_22612,N_22905);
nor U24932 (N_24932,N_23474,N_23436);
nand U24933 (N_24933,N_23105,N_22966);
nor U24934 (N_24934,N_23487,N_22608);
or U24935 (N_24935,N_23693,N_23605);
xnor U24936 (N_24936,N_23052,N_22961);
and U24937 (N_24937,N_23455,N_22520);
nor U24938 (N_24938,N_23143,N_22995);
nand U24939 (N_24939,N_22826,N_23123);
and U24940 (N_24940,N_23594,N_22652);
or U24941 (N_24941,N_23267,N_23224);
or U24942 (N_24942,N_23681,N_23302);
and U24943 (N_24943,N_22709,N_23150);
nand U24944 (N_24944,N_23606,N_23355);
nor U24945 (N_24945,N_23105,N_23237);
xnor U24946 (N_24946,N_23183,N_23091);
nor U24947 (N_24947,N_22752,N_23014);
nor U24948 (N_24948,N_23606,N_23464);
nor U24949 (N_24949,N_22822,N_23138);
nor U24950 (N_24950,N_23538,N_23349);
nor U24951 (N_24951,N_23157,N_23693);
xnor U24952 (N_24952,N_23134,N_23372);
nor U24953 (N_24953,N_22700,N_23069);
nor U24954 (N_24954,N_23564,N_22733);
nand U24955 (N_24955,N_22889,N_22738);
or U24956 (N_24956,N_22718,N_23498);
nor U24957 (N_24957,N_23028,N_22632);
xor U24958 (N_24958,N_23067,N_22827);
or U24959 (N_24959,N_22997,N_22888);
xor U24960 (N_24960,N_22598,N_22626);
or U24961 (N_24961,N_23217,N_23477);
xor U24962 (N_24962,N_22743,N_23552);
nand U24963 (N_24963,N_23585,N_23151);
xor U24964 (N_24964,N_23132,N_23447);
nand U24965 (N_24965,N_22557,N_23434);
nor U24966 (N_24966,N_23632,N_23328);
nand U24967 (N_24967,N_22906,N_23193);
nand U24968 (N_24968,N_22689,N_23138);
nor U24969 (N_24969,N_23714,N_23127);
nor U24970 (N_24970,N_23086,N_22565);
and U24971 (N_24971,N_22504,N_23629);
xor U24972 (N_24972,N_23198,N_23319);
xor U24973 (N_24973,N_23114,N_23450);
xnor U24974 (N_24974,N_23384,N_23388);
xnor U24975 (N_24975,N_22746,N_23617);
nand U24976 (N_24976,N_22861,N_22675);
nor U24977 (N_24977,N_23077,N_23243);
and U24978 (N_24978,N_22987,N_22632);
or U24979 (N_24979,N_23605,N_22691);
nand U24980 (N_24980,N_23109,N_23709);
and U24981 (N_24981,N_23154,N_23200);
and U24982 (N_24982,N_23532,N_22967);
and U24983 (N_24983,N_22547,N_23043);
or U24984 (N_24984,N_23110,N_22984);
nor U24985 (N_24985,N_23275,N_22530);
xor U24986 (N_24986,N_23231,N_23001);
and U24987 (N_24987,N_22806,N_23577);
nand U24988 (N_24988,N_23165,N_22586);
nand U24989 (N_24989,N_23269,N_23680);
xor U24990 (N_24990,N_23481,N_22651);
nor U24991 (N_24991,N_23106,N_22879);
and U24992 (N_24992,N_23302,N_23203);
and U24993 (N_24993,N_23230,N_23580);
nand U24994 (N_24994,N_22917,N_22738);
nor U24995 (N_24995,N_23538,N_22860);
xnor U24996 (N_24996,N_23235,N_23021);
or U24997 (N_24997,N_23142,N_22550);
nand U24998 (N_24998,N_23161,N_23453);
nand U24999 (N_24999,N_23647,N_23369);
or UO_0 (O_0,N_24436,N_23889);
nand UO_1 (O_1,N_24228,N_24994);
or UO_2 (O_2,N_24226,N_24669);
nor UO_3 (O_3,N_24772,N_24018);
nand UO_4 (O_4,N_24380,N_24538);
and UO_5 (O_5,N_24584,N_24204);
nor UO_6 (O_6,N_24271,N_24555);
xnor UO_7 (O_7,N_24747,N_24510);
xor UO_8 (O_8,N_24280,N_24536);
and UO_9 (O_9,N_24615,N_23803);
and UO_10 (O_10,N_24451,N_23960);
nor UO_11 (O_11,N_24567,N_24983);
nor UO_12 (O_12,N_24409,N_24320);
xnor UO_13 (O_13,N_24800,N_24680);
and UO_14 (O_14,N_24743,N_24394);
or UO_15 (O_15,N_24633,N_24992);
nor UO_16 (O_16,N_24617,N_24864);
and UO_17 (O_17,N_24110,N_24881);
and UO_18 (O_18,N_24890,N_24739);
and UO_19 (O_19,N_23865,N_24420);
xnor UO_20 (O_20,N_24075,N_24533);
or UO_21 (O_21,N_24054,N_24612);
or UO_22 (O_22,N_24738,N_24735);
nor UO_23 (O_23,N_24951,N_24687);
xnor UO_24 (O_24,N_24919,N_24129);
xor UO_25 (O_25,N_24091,N_24435);
or UO_26 (O_26,N_24767,N_24643);
xnor UO_27 (O_27,N_24608,N_24681);
nand UO_28 (O_28,N_23918,N_24086);
and UO_29 (O_29,N_24816,N_24067);
or UO_30 (O_30,N_24064,N_24469);
nor UO_31 (O_31,N_24880,N_24684);
and UO_32 (O_32,N_24381,N_24023);
or UO_33 (O_33,N_24166,N_24857);
or UO_34 (O_34,N_24611,N_24480);
and UO_35 (O_35,N_24526,N_24786);
xor UO_36 (O_36,N_24289,N_24809);
nand UO_37 (O_37,N_24205,N_24286);
nand UO_38 (O_38,N_24902,N_24970);
nand UO_39 (O_39,N_24182,N_24984);
xnor UO_40 (O_40,N_24486,N_24917);
or UO_41 (O_41,N_24155,N_24650);
or UO_42 (O_42,N_24832,N_24465);
and UO_43 (O_43,N_24327,N_24231);
and UO_44 (O_44,N_24516,N_24243);
nor UO_45 (O_45,N_24683,N_24980);
xor UO_46 (O_46,N_24833,N_24920);
or UO_47 (O_47,N_24063,N_24041);
nand UO_48 (O_48,N_24493,N_24393);
nor UO_49 (O_49,N_24597,N_23826);
nor UO_50 (O_50,N_24167,N_23975);
nor UO_51 (O_51,N_24214,N_24048);
xnor UO_52 (O_52,N_24812,N_23951);
or UO_53 (O_53,N_24095,N_24802);
xnor UO_54 (O_54,N_24246,N_24413);
nor UO_55 (O_55,N_24066,N_23804);
or UO_56 (O_56,N_24093,N_24478);
nor UO_57 (O_57,N_24736,N_24944);
nand UO_58 (O_58,N_23989,N_24826);
nor UO_59 (O_59,N_23993,N_24689);
or UO_60 (O_60,N_24838,N_24887);
nand UO_61 (O_61,N_24532,N_23780);
nand UO_62 (O_62,N_24116,N_23832);
nand UO_63 (O_63,N_24117,N_24047);
nor UO_64 (O_64,N_24755,N_24400);
or UO_65 (O_65,N_23793,N_24468);
and UO_66 (O_66,N_24235,N_24589);
xor UO_67 (O_67,N_24343,N_24044);
nand UO_68 (O_68,N_24607,N_24457);
nor UO_69 (O_69,N_24730,N_24834);
and UO_70 (O_70,N_24808,N_24978);
or UO_71 (O_71,N_23927,N_24200);
nand UO_72 (O_72,N_24520,N_24998);
nor UO_73 (O_73,N_24446,N_24931);
xnor UO_74 (O_74,N_24153,N_23882);
xor UO_75 (O_75,N_24550,N_23773);
xnor UO_76 (O_76,N_24562,N_24316);
nand UO_77 (O_77,N_24328,N_23753);
and UO_78 (O_78,N_24258,N_24215);
nand UO_79 (O_79,N_24563,N_23892);
and UO_80 (O_80,N_24311,N_24999);
and UO_81 (O_81,N_24752,N_24412);
xnor UO_82 (O_82,N_24481,N_24038);
and UO_83 (O_83,N_23774,N_24933);
and UO_84 (O_84,N_24025,N_23905);
or UO_85 (O_85,N_24028,N_24804);
nor UO_86 (O_86,N_24350,N_24900);
nor UO_87 (O_87,N_23788,N_23762);
nand UO_88 (O_88,N_24768,N_24169);
nor UO_89 (O_89,N_24896,N_24453);
nand UO_90 (O_90,N_24461,N_24694);
nand UO_91 (O_91,N_24337,N_24947);
xor UO_92 (O_92,N_23974,N_24954);
xor UO_93 (O_93,N_24644,N_24097);
or UO_94 (O_94,N_24924,N_24484);
nand UO_95 (O_95,N_23833,N_23821);
nand UO_96 (O_96,N_24438,N_24870);
nor UO_97 (O_97,N_24294,N_24572);
or UO_98 (O_98,N_23890,N_24418);
nand UO_99 (O_99,N_24784,N_24189);
and UO_100 (O_100,N_24259,N_24729);
nor UO_101 (O_101,N_24385,N_24460);
xnor UO_102 (O_102,N_24073,N_24770);
or UO_103 (O_103,N_24679,N_23866);
xnor UO_104 (O_104,N_23979,N_24988);
or UO_105 (O_105,N_24540,N_23840);
and UO_106 (O_106,N_23783,N_24108);
nor UO_107 (O_107,N_24524,N_24839);
xor UO_108 (O_108,N_24444,N_24569);
nand UO_109 (O_109,N_24886,N_24514);
or UO_110 (O_110,N_24213,N_23913);
and UO_111 (O_111,N_24766,N_24971);
and UO_112 (O_112,N_23864,N_24317);
and UO_113 (O_113,N_24973,N_24100);
and UO_114 (O_114,N_23873,N_23926);
nand UO_115 (O_115,N_24270,N_24255);
or UO_116 (O_116,N_24244,N_23942);
or UO_117 (O_117,N_24375,N_24570);
or UO_118 (O_118,N_23827,N_24969);
and UO_119 (O_119,N_24163,N_23949);
xnor UO_120 (O_120,N_23921,N_23966);
nand UO_121 (O_121,N_24358,N_24898);
or UO_122 (O_122,N_23895,N_24665);
xnor UO_123 (O_123,N_24421,N_24130);
xor UO_124 (O_124,N_24821,N_24009);
nor UO_125 (O_125,N_24829,N_24267);
nor UO_126 (O_126,N_24657,N_24642);
xnor UO_127 (O_127,N_23811,N_24002);
or UO_128 (O_128,N_24362,N_24485);
nand UO_129 (O_129,N_24856,N_23983);
xor UO_130 (O_130,N_23829,N_23992);
or UO_131 (O_131,N_23964,N_24703);
and UO_132 (O_132,N_23845,N_23883);
and UO_133 (O_133,N_23950,N_23815);
xor UO_134 (O_134,N_23791,N_23984);
nor UO_135 (O_135,N_24777,N_24348);
nand UO_136 (O_136,N_24525,N_24915);
and UO_137 (O_137,N_23901,N_24760);
and UO_138 (O_138,N_24692,N_24387);
nor UO_139 (O_139,N_24245,N_24952);
xor UO_140 (O_140,N_24033,N_24434);
nor UO_141 (O_141,N_24197,N_24489);
and UO_142 (O_142,N_24397,N_24229);
xnor UO_143 (O_143,N_24728,N_23777);
and UO_144 (O_144,N_24552,N_23999);
or UO_145 (O_145,N_24551,N_24654);
and UO_146 (O_146,N_24256,N_24930);
xnor UO_147 (O_147,N_24504,N_24344);
and UO_148 (O_148,N_24123,N_23917);
and UO_149 (O_149,N_23981,N_24875);
or UO_150 (O_150,N_24517,N_24744);
nand UO_151 (O_151,N_24714,N_24899);
or UO_152 (O_152,N_24844,N_24748);
nor UO_153 (O_153,N_24141,N_24353);
nand UO_154 (O_154,N_24989,N_24072);
xnor UO_155 (O_155,N_24771,N_24577);
nor UO_156 (O_156,N_24906,N_23785);
nand UO_157 (O_157,N_24008,N_24871);
nand UO_158 (O_158,N_24634,N_23766);
nand UO_159 (O_159,N_24962,N_24691);
nor UO_160 (O_160,N_24174,N_24233);
xor UO_161 (O_161,N_23795,N_23779);
xnor UO_162 (O_162,N_23843,N_24805);
xnor UO_163 (O_163,N_24170,N_23904);
and UO_164 (O_164,N_24333,N_24661);
xor UO_165 (O_165,N_24836,N_24125);
nor UO_166 (O_166,N_24464,N_23976);
nor UO_167 (O_167,N_24195,N_24712);
and UO_168 (O_168,N_23899,N_24997);
or UO_169 (O_169,N_24212,N_23813);
nand UO_170 (O_170,N_23805,N_24807);
or UO_171 (O_171,N_24721,N_24926);
xnor UO_172 (O_172,N_24053,N_23969);
or UO_173 (O_173,N_23959,N_24945);
nand UO_174 (O_174,N_24151,N_24279);
or UO_175 (O_175,N_23887,N_24144);
nand UO_176 (O_176,N_24559,N_24827);
and UO_177 (O_177,N_24003,N_24496);
nor UO_178 (O_178,N_24892,N_24012);
nor UO_179 (O_179,N_24290,N_23879);
xor UO_180 (O_180,N_24699,N_24234);
and UO_181 (O_181,N_24720,N_24456);
xnor UO_182 (O_182,N_24395,N_24031);
or UO_183 (O_183,N_24943,N_24627);
or UO_184 (O_184,N_23770,N_24210);
xor UO_185 (O_185,N_24713,N_23799);
or UO_186 (O_186,N_24872,N_24863);
nand UO_187 (O_187,N_24056,N_23838);
nand UO_188 (O_188,N_24284,N_23877);
nand UO_189 (O_189,N_24495,N_24102);
nand UO_190 (O_190,N_24652,N_24869);
nand UO_191 (O_191,N_24599,N_24614);
nor UO_192 (O_192,N_24977,N_23851);
nor UO_193 (O_193,N_24512,N_24842);
and UO_194 (O_194,N_23776,N_23841);
xor UO_195 (O_195,N_24027,N_24806);
nand UO_196 (O_196,N_24554,N_24497);
xnor UO_197 (O_197,N_24884,N_24542);
nor UO_198 (O_198,N_24249,N_24430);
xnor UO_199 (O_199,N_23856,N_23825);
and UO_200 (O_200,N_24587,N_24660);
and UO_201 (O_201,N_24410,N_23800);
xnor UO_202 (O_202,N_24157,N_24172);
xnor UO_203 (O_203,N_24326,N_24301);
xnor UO_204 (O_204,N_24849,N_24648);
or UO_205 (O_205,N_24052,N_24447);
or UO_206 (O_206,N_24773,N_23850);
xnor UO_207 (O_207,N_24603,N_24574);
and UO_208 (O_208,N_24678,N_24077);
and UO_209 (O_209,N_24814,N_24787);
and UO_210 (O_210,N_24579,N_23757);
or UO_211 (O_211,N_23947,N_24422);
or UO_212 (O_212,N_24291,N_24257);
and UO_213 (O_213,N_24855,N_24145);
or UO_214 (O_214,N_23937,N_24763);
nand UO_215 (O_215,N_24113,N_23994);
or UO_216 (O_216,N_24960,N_24873);
or UO_217 (O_217,N_24349,N_24238);
nand UO_218 (O_218,N_24490,N_24363);
or UO_219 (O_219,N_23962,N_24639);
and UO_220 (O_220,N_24181,N_24606);
xor UO_221 (O_221,N_24758,N_24019);
nand UO_222 (O_222,N_24336,N_23908);
nor UO_223 (O_223,N_24148,N_23941);
nor UO_224 (O_224,N_24891,N_24283);
xor UO_225 (O_225,N_24993,N_24180);
xnor UO_226 (O_226,N_23798,N_23853);
nor UO_227 (O_227,N_23818,N_24521);
nand UO_228 (O_228,N_24860,N_24641);
xnor UO_229 (O_229,N_23836,N_24368);
xor UO_230 (O_230,N_24726,N_24621);
nand UO_231 (O_231,N_24000,N_24741);
nor UO_232 (O_232,N_24927,N_24663);
nor UO_233 (O_233,N_24079,N_24548);
xnor UO_234 (O_234,N_24414,N_24794);
and UO_235 (O_235,N_24094,N_24841);
nand UO_236 (O_236,N_24136,N_24357);
or UO_237 (O_237,N_23857,N_24388);
nand UO_238 (O_238,N_24390,N_24107);
or UO_239 (O_239,N_24408,N_23801);
xor UO_240 (O_240,N_24923,N_24928);
nand UO_241 (O_241,N_24737,N_24037);
xnor UO_242 (O_242,N_24757,N_24274);
and UO_243 (O_243,N_24640,N_23953);
nand UO_244 (O_244,N_24754,N_24433);
nand UO_245 (O_245,N_23973,N_24275);
and UO_246 (O_246,N_24901,N_24137);
nand UO_247 (O_247,N_24454,N_24261);
xnor UO_248 (O_248,N_24253,N_24017);
nand UO_249 (O_249,N_24304,N_24076);
xor UO_250 (O_250,N_24840,N_24964);
nor UO_251 (O_251,N_23823,N_24020);
xor UO_252 (O_252,N_24473,N_24178);
and UO_253 (O_253,N_24658,N_24146);
nor UO_254 (O_254,N_24985,N_24475);
and UO_255 (O_255,N_24043,N_24698);
nor UO_256 (O_256,N_24143,N_24693);
xor UO_257 (O_257,N_24345,N_24332);
and UO_258 (O_258,N_24734,N_24491);
nand UO_259 (O_259,N_24957,N_24785);
nand UO_260 (O_260,N_24531,N_24329);
xnor UO_261 (O_261,N_24553,N_24398);
nor UO_262 (O_262,N_24188,N_24903);
nand UO_263 (O_263,N_23971,N_24049);
nand UO_264 (O_264,N_23876,N_23920);
and UO_265 (O_265,N_24797,N_23977);
nor UO_266 (O_266,N_24470,N_24585);
and UO_267 (O_267,N_23824,N_24401);
nor UO_268 (O_268,N_24556,N_24050);
xnor UO_269 (O_269,N_24426,N_24583);
xnor UO_270 (O_270,N_23986,N_24668);
xnor UO_271 (O_271,N_24367,N_24407);
and UO_272 (O_272,N_24600,N_24528);
xor UO_273 (O_273,N_24352,N_23752);
and UO_274 (O_274,N_24742,N_24651);
nand UO_275 (O_275,N_24152,N_24222);
or UO_276 (O_276,N_24177,N_24011);
or UO_277 (O_277,N_24783,N_24365);
nor UO_278 (O_278,N_24040,N_24030);
nor UO_279 (O_279,N_24934,N_24402);
nor UO_280 (O_280,N_24288,N_24529);
xnor UO_281 (O_281,N_23781,N_24282);
or UO_282 (O_282,N_24618,N_24431);
nand UO_283 (O_283,N_24990,N_24662);
or UO_284 (O_284,N_23846,N_24090);
nand UO_285 (O_285,N_24069,N_24711);
or UO_286 (O_286,N_24637,N_24013);
nor UO_287 (O_287,N_23807,N_24450);
xor UO_288 (O_288,N_24192,N_24124);
nand UO_289 (O_289,N_24087,N_23855);
nand UO_290 (O_290,N_24299,N_24005);
and UO_291 (O_291,N_24498,N_24789);
nand UO_292 (O_292,N_24740,N_24428);
nand UO_293 (O_293,N_23810,N_23784);
and UO_294 (O_294,N_24686,N_24974);
xnor UO_295 (O_295,N_23884,N_24996);
nand UO_296 (O_296,N_24967,N_24287);
nor UO_297 (O_297,N_24494,N_24265);
and UO_298 (O_298,N_24126,N_24861);
or UO_299 (O_299,N_24061,N_24946);
nor UO_300 (O_300,N_24191,N_24846);
nor UO_301 (O_301,N_24883,N_24396);
nor UO_302 (O_302,N_24732,N_23998);
nor UO_303 (O_303,N_24968,N_23952);
and UO_304 (O_304,N_24937,N_24975);
or UO_305 (O_305,N_24549,N_24057);
nor UO_306 (O_306,N_24866,N_23933);
and UO_307 (O_307,N_24862,N_24035);
xnor UO_308 (O_308,N_24399,N_24092);
or UO_309 (O_309,N_24466,N_24753);
and UO_310 (O_310,N_24854,N_24254);
xor UO_311 (O_311,N_24297,N_24708);
nand UO_312 (O_312,N_24459,N_24196);
and UO_313 (O_313,N_24893,N_24389);
xor UO_314 (O_314,N_23914,N_24488);
and UO_315 (O_315,N_24697,N_24194);
or UO_316 (O_316,N_24798,N_24360);
nand UO_317 (O_317,N_24622,N_24543);
nor UO_318 (O_318,N_24750,N_23754);
xnor UO_319 (O_319,N_24929,N_23852);
xor UO_320 (O_320,N_24058,N_24247);
xnor UO_321 (O_321,N_24472,N_24340);
or UO_322 (O_322,N_24670,N_24305);
nor UO_323 (O_323,N_24649,N_24746);
nand UO_324 (O_324,N_23764,N_24266);
or UO_325 (O_325,N_24576,N_24822);
and UO_326 (O_326,N_23861,N_23980);
and UO_327 (O_327,N_24628,N_24239);
xnor UO_328 (O_328,N_23844,N_24404);
or UO_329 (O_329,N_24103,N_24625);
and UO_330 (O_330,N_24101,N_24021);
nand UO_331 (O_331,N_24935,N_24225);
nor UO_332 (O_332,N_24309,N_24133);
or UO_333 (O_333,N_24879,N_23787);
or UO_334 (O_334,N_24016,N_23871);
and UO_335 (O_335,N_24190,N_23909);
and UO_336 (O_336,N_24185,N_24306);
and UO_337 (O_337,N_24448,N_24825);
or UO_338 (O_338,N_24765,N_23830);
and UO_339 (O_339,N_24251,N_24582);
and UO_340 (O_340,N_24815,N_24843);
and UO_341 (O_341,N_24965,N_24014);
and UO_342 (O_342,N_24232,N_23847);
xnor UO_343 (O_343,N_24314,N_24132);
nand UO_344 (O_344,N_24573,N_23790);
or UO_345 (O_345,N_24847,N_24034);
nand UO_346 (O_346,N_23802,N_24590);
or UO_347 (O_347,N_23831,N_24745);
nand UO_348 (O_348,N_24307,N_23988);
and UO_349 (O_349,N_24281,N_23771);
or UO_350 (O_350,N_24509,N_23842);
xnor UO_351 (O_351,N_24122,N_23996);
and UO_352 (O_352,N_24636,N_23903);
xor UO_353 (O_353,N_24082,N_24706);
xnor UO_354 (O_354,N_24791,N_23859);
nand UO_355 (O_355,N_24359,N_24515);
nor UO_356 (O_356,N_24346,N_24913);
nand UO_357 (O_357,N_24723,N_24260);
nand UO_358 (O_358,N_24790,N_24386);
and UO_359 (O_359,N_24564,N_24131);
or UO_360 (O_360,N_24492,N_24065);
or UO_361 (O_361,N_24593,N_24487);
or UO_362 (O_362,N_24263,N_24149);
nor UO_363 (O_363,N_24823,N_23778);
nor UO_364 (O_364,N_24764,N_24318);
and UO_365 (O_365,N_24756,N_24010);
nand UO_366 (O_366,N_24972,N_23751);
and UO_367 (O_367,N_24793,N_23990);
xor UO_368 (O_368,N_23849,N_23970);
xnor UO_369 (O_369,N_24114,N_23911);
nand UO_370 (O_370,N_24904,N_23796);
nand UO_371 (O_371,N_24949,N_24530);
and UO_372 (O_372,N_24656,N_24203);
and UO_373 (O_373,N_23935,N_24848);
or UO_374 (O_374,N_23944,N_24221);
and UO_375 (O_375,N_23956,N_24334);
nand UO_376 (O_376,N_24032,N_24922);
and UO_377 (O_377,N_24704,N_24276);
and UO_378 (O_378,N_24458,N_24961);
and UO_379 (O_379,N_23880,N_24323);
nand UO_380 (O_380,N_24685,N_23888);
and UO_381 (O_381,N_23972,N_24119);
nand UO_382 (O_382,N_23875,N_24505);
xor UO_383 (O_383,N_24819,N_24779);
nand UO_384 (O_384,N_24331,N_24128);
and UO_385 (O_385,N_24022,N_24051);
or UO_386 (O_386,N_24004,N_24070);
nand UO_387 (O_387,N_24580,N_24074);
or UO_388 (O_388,N_24595,N_24199);
or UO_389 (O_389,N_24026,N_24987);
or UO_390 (O_390,N_24632,N_24546);
nand UO_391 (O_391,N_24293,N_23997);
or UO_392 (O_392,N_24731,N_23878);
xor UO_393 (O_393,N_24184,N_24820);
nor UO_394 (O_394,N_24780,N_24921);
nor UO_395 (O_395,N_24059,N_24262);
or UO_396 (O_396,N_24162,N_24217);
nor UO_397 (O_397,N_23794,N_24361);
or UO_398 (O_398,N_24725,N_24224);
and UO_399 (O_399,N_24046,N_23822);
or UO_400 (O_400,N_24912,N_24139);
nand UO_401 (O_401,N_23835,N_23806);
nor UO_402 (O_402,N_24853,N_24384);
or UO_403 (O_403,N_24624,N_23946);
or UO_404 (O_404,N_23934,N_24609);
nand UO_405 (O_405,N_24068,N_24187);
xor UO_406 (O_406,N_24062,N_24308);
xor UO_407 (O_407,N_24324,N_23967);
xor UO_408 (O_408,N_24558,N_24635);
nand UO_409 (O_409,N_24575,N_24581);
nor UO_410 (O_410,N_24613,N_24701);
xor UO_411 (O_411,N_23812,N_24941);
or UO_412 (O_412,N_24541,N_24586);
xnor UO_413 (O_413,N_24700,N_23965);
and UO_414 (O_414,N_23902,N_24423);
nand UO_415 (O_415,N_24695,N_24845);
or UO_416 (O_416,N_24278,N_24227);
nor UO_417 (O_417,N_24707,N_23943);
or UO_418 (O_418,N_24950,N_24598);
and UO_419 (O_419,N_24120,N_24769);
nand UO_420 (O_420,N_24751,N_24476);
xnor UO_421 (O_421,N_24623,N_24594);
or UO_422 (O_422,N_24277,N_24201);
or UO_423 (O_423,N_24591,N_24406);
nand UO_424 (O_424,N_24939,N_24905);
xor UO_425 (O_425,N_24440,N_24437);
nor UO_426 (O_426,N_24302,N_24813);
xnor UO_427 (O_427,N_24338,N_24672);
nand UO_428 (O_428,N_24150,N_24015);
and UO_429 (O_429,N_24176,N_24925);
xor UO_430 (O_430,N_24682,N_24981);
or UO_431 (O_431,N_24183,N_24909);
nand UO_432 (O_432,N_24850,N_24868);
or UO_433 (O_433,N_23995,N_23928);
or UO_434 (O_434,N_24330,N_24718);
or UO_435 (O_435,N_24801,N_24976);
xnor UO_436 (O_436,N_23936,N_24852);
nor UO_437 (O_437,N_24006,N_24571);
nand UO_438 (O_438,N_24055,N_24513);
nand UO_439 (O_439,N_24370,N_24303);
xor UO_440 (O_440,N_24932,N_24830);
or UO_441 (O_441,N_24715,N_24664);
xor UO_442 (O_442,N_24774,N_23894);
nor UO_443 (O_443,N_24508,N_24161);
or UO_444 (O_444,N_24001,N_24310);
or UO_445 (O_445,N_23828,N_23767);
nand UO_446 (O_446,N_23867,N_24121);
nand UO_447 (O_447,N_23819,N_24206);
or UO_448 (O_448,N_24667,N_24722);
nor UO_449 (O_449,N_24429,N_24795);
and UO_450 (O_450,N_24717,N_24817);
and UO_451 (O_451,N_24631,N_23820);
and UO_452 (O_452,N_23958,N_24938);
nand UO_453 (O_453,N_23915,N_24544);
nor UO_454 (O_454,N_23991,N_23925);
or UO_455 (O_455,N_24874,N_24749);
and UO_456 (O_456,N_24218,N_24250);
nor UO_457 (O_457,N_24273,N_24193);
nand UO_458 (O_458,N_24354,N_24710);
xor UO_459 (O_459,N_23924,N_24953);
xor UO_460 (O_460,N_24036,N_23982);
or UO_461 (O_461,N_23870,N_24986);
and UO_462 (O_462,N_23931,N_24759);
and UO_463 (O_463,N_24118,N_24566);
and UO_464 (O_464,N_23987,N_24106);
and UO_465 (O_465,N_24878,N_24078);
and UO_466 (O_466,N_24810,N_24319);
or UO_467 (O_467,N_23922,N_24539);
nand UO_468 (O_468,N_24392,N_24391);
and UO_469 (O_469,N_24455,N_23860);
nor UO_470 (O_470,N_24379,N_23816);
xnor UO_471 (O_471,N_24463,N_23814);
and UO_472 (O_472,N_24241,N_24138);
xor UO_473 (O_473,N_24604,N_24963);
and UO_474 (O_474,N_24676,N_24557);
and UO_475 (O_475,N_24500,N_24154);
and UO_476 (O_476,N_24762,N_24364);
xor UO_477 (O_477,N_24376,N_24479);
and UO_478 (O_478,N_23885,N_24089);
nand UO_479 (O_479,N_23863,N_24907);
nand UO_480 (O_480,N_24503,N_24220);
xnor UO_481 (O_481,N_24216,N_24502);
xnor UO_482 (O_482,N_24776,N_24709);
xor UO_483 (O_483,N_24518,N_24778);
xor UO_484 (O_484,N_24104,N_24111);
xnor UO_485 (O_485,N_23869,N_24908);
xnor UO_486 (O_486,N_24824,N_24351);
or UO_487 (O_487,N_24596,N_24877);
nor UO_488 (O_488,N_24335,N_24171);
nand UO_489 (O_489,N_24416,N_24702);
and UO_490 (O_490,N_23961,N_24948);
and UO_491 (O_491,N_24208,N_24083);
nor UO_492 (O_492,N_24527,N_24207);
nor UO_493 (O_493,N_24135,N_24115);
or UO_494 (O_494,N_24382,N_24088);
xor UO_495 (O_495,N_24647,N_24888);
and UO_496 (O_496,N_23797,N_24084);
and UO_497 (O_497,N_24782,N_23769);
nand UO_498 (O_498,N_24230,N_24638);
nor UO_499 (O_499,N_23916,N_24383);
and UO_500 (O_500,N_24158,N_24347);
xnor UO_501 (O_501,N_24796,N_24911);
xnor UO_502 (O_502,N_23763,N_24705);
and UO_503 (O_503,N_24610,N_23930);
nor UO_504 (O_504,N_24405,N_24958);
or UO_505 (O_505,N_24173,N_23868);
xor UO_506 (O_506,N_23848,N_23837);
xnor UO_507 (O_507,N_24507,N_24630);
nor UO_508 (O_508,N_24858,N_24042);
or UO_509 (O_509,N_24865,N_24837);
nor UO_510 (O_510,N_24415,N_24372);
nand UO_511 (O_511,N_24355,N_24443);
or UO_512 (O_512,N_23910,N_24240);
and UO_513 (O_513,N_23782,N_23808);
nor UO_514 (O_514,N_24325,N_23896);
nand UO_515 (O_515,N_24522,N_24223);
nor UO_516 (O_516,N_24105,N_24356);
xnor UO_517 (O_517,N_24168,N_23758);
or UO_518 (O_518,N_23765,N_24897);
nor UO_519 (O_519,N_24164,N_24688);
nor UO_520 (O_520,N_23900,N_23862);
and UO_521 (O_521,N_24198,N_24403);
or UO_522 (O_522,N_23929,N_24761);
xor UO_523 (O_523,N_23755,N_24727);
nor UO_524 (O_524,N_24537,N_24202);
xnor UO_525 (O_525,N_24775,N_24876);
and UO_526 (O_526,N_24620,N_24236);
nand UO_527 (O_527,N_23940,N_24442);
nor UO_528 (O_528,N_24237,N_24675);
xnor UO_529 (O_529,N_23954,N_24080);
nor UO_530 (O_530,N_23945,N_24646);
and UO_531 (O_531,N_24616,N_24313);
xnor UO_532 (O_532,N_24673,N_24109);
or UO_533 (O_533,N_24535,N_24578);
nand UO_534 (O_534,N_24272,N_23839);
nand UO_535 (O_535,N_24916,N_24966);
and UO_536 (O_536,N_24506,N_24483);
nor UO_537 (O_537,N_24499,N_23874);
and UO_538 (O_538,N_24373,N_24671);
and UO_539 (O_539,N_23919,N_23817);
xnor UO_540 (O_540,N_24914,N_24955);
and UO_541 (O_541,N_24142,N_24296);
or UO_542 (O_542,N_24165,N_24096);
or UO_543 (O_543,N_24565,N_24127);
nor UO_544 (O_544,N_23760,N_24264);
nor UO_545 (O_545,N_24523,N_24645);
and UO_546 (O_546,N_24602,N_24605);
nand UO_547 (O_547,N_23768,N_23759);
nand UO_548 (O_548,N_24534,N_24690);
nand UO_549 (O_549,N_24482,N_23939);
nand UO_550 (O_550,N_24979,N_24099);
and UO_551 (O_551,N_24268,N_24071);
nand UO_552 (O_552,N_24219,N_24991);
or UO_553 (O_553,N_24098,N_24894);
or UO_554 (O_554,N_24285,N_24186);
or UO_555 (O_555,N_24369,N_24792);
nand UO_556 (O_556,N_24511,N_24248);
nor UO_557 (O_557,N_24432,N_24885);
or UO_558 (O_558,N_24147,N_24321);
xnor UO_559 (O_559,N_24024,N_24159);
or UO_560 (O_560,N_24995,N_24462);
xor UO_561 (O_561,N_24209,N_24788);
nor UO_562 (O_562,N_23978,N_24677);
xnor UO_563 (O_563,N_24910,N_24439);
nand UO_564 (O_564,N_24867,N_24477);
xor UO_565 (O_565,N_24659,N_24724);
nand UO_566 (O_566,N_24242,N_23750);
xor UO_567 (O_567,N_24085,N_24889);
and UO_568 (O_568,N_24269,N_24560);
and UO_569 (O_569,N_23834,N_24882);
nand UO_570 (O_570,N_24851,N_24696);
nand UO_571 (O_571,N_24547,N_24942);
and UO_572 (O_572,N_23858,N_24377);
nor UO_573 (O_573,N_24959,N_24342);
nand UO_574 (O_574,N_24471,N_24211);
nand UO_575 (O_575,N_23985,N_24561);
nor UO_576 (O_576,N_23938,N_24982);
or UO_577 (O_577,N_23775,N_24626);
nand UO_578 (O_578,N_24039,N_24179);
nor UO_579 (O_579,N_24341,N_24315);
xor UO_580 (O_580,N_23761,N_24588);
and UO_581 (O_581,N_24060,N_23772);
or UO_582 (O_582,N_23756,N_24956);
nor UO_583 (O_583,N_23897,N_24918);
nand UO_584 (O_584,N_24859,N_24936);
nor UO_585 (O_585,N_23968,N_23881);
nor UO_586 (O_586,N_24295,N_23906);
nor UO_587 (O_587,N_24160,N_24568);
xnor UO_588 (O_588,N_24417,N_24474);
and UO_589 (O_589,N_23809,N_24029);
nor UO_590 (O_590,N_24449,N_24501);
nor UO_591 (O_591,N_24629,N_24424);
and UO_592 (O_592,N_24411,N_24895);
nor UO_593 (O_593,N_23891,N_24339);
nor UO_594 (O_594,N_23893,N_24175);
nand UO_595 (O_595,N_24467,N_23872);
xnor UO_596 (O_596,N_24156,N_24045);
and UO_597 (O_597,N_24298,N_24371);
or UO_598 (O_598,N_24312,N_24445);
or UO_599 (O_599,N_24378,N_23955);
nor UO_600 (O_600,N_24716,N_24140);
or UO_601 (O_601,N_24427,N_24666);
nand UO_602 (O_602,N_24835,N_24799);
nand UO_603 (O_603,N_23854,N_23963);
xnor UO_604 (O_604,N_24007,N_24322);
or UO_605 (O_605,N_24803,N_24134);
xnor UO_606 (O_606,N_24619,N_24940);
nand UO_607 (O_607,N_24818,N_24831);
nand UO_608 (O_608,N_24081,N_23789);
and UO_609 (O_609,N_24733,N_23912);
nand UO_610 (O_610,N_24252,N_24828);
nor UO_611 (O_611,N_24781,N_24811);
and UO_612 (O_612,N_24655,N_24441);
nor UO_613 (O_613,N_23792,N_24425);
and UO_614 (O_614,N_23923,N_24366);
or UO_615 (O_615,N_24601,N_24419);
nor UO_616 (O_616,N_24292,N_24519);
nand UO_617 (O_617,N_23957,N_24452);
and UO_618 (O_618,N_23948,N_24592);
nand UO_619 (O_619,N_24674,N_23898);
and UO_620 (O_620,N_23886,N_24719);
and UO_621 (O_621,N_24300,N_24374);
xor UO_622 (O_622,N_23932,N_24545);
and UO_623 (O_623,N_23907,N_24112);
xnor UO_624 (O_624,N_23786,N_24653);
or UO_625 (O_625,N_23944,N_24378);
nand UO_626 (O_626,N_24808,N_23993);
or UO_627 (O_627,N_24462,N_24602);
xor UO_628 (O_628,N_24457,N_24351);
xnor UO_629 (O_629,N_24440,N_24675);
xor UO_630 (O_630,N_24593,N_24473);
xnor UO_631 (O_631,N_24460,N_23948);
nor UO_632 (O_632,N_24274,N_24960);
and UO_633 (O_633,N_24579,N_24978);
xnor UO_634 (O_634,N_24265,N_24854);
nand UO_635 (O_635,N_24335,N_23786);
nor UO_636 (O_636,N_24922,N_24493);
and UO_637 (O_637,N_23753,N_23887);
xor UO_638 (O_638,N_24047,N_24013);
nand UO_639 (O_639,N_24867,N_24590);
nand UO_640 (O_640,N_24613,N_24381);
nand UO_641 (O_641,N_24417,N_24466);
nor UO_642 (O_642,N_24969,N_24413);
xor UO_643 (O_643,N_24269,N_23784);
nor UO_644 (O_644,N_24034,N_24556);
nand UO_645 (O_645,N_24121,N_24287);
nand UO_646 (O_646,N_24114,N_24416);
or UO_647 (O_647,N_24569,N_24491);
nand UO_648 (O_648,N_23995,N_24852);
and UO_649 (O_649,N_24347,N_23912);
nor UO_650 (O_650,N_23770,N_24254);
xor UO_651 (O_651,N_24306,N_23879);
or UO_652 (O_652,N_24882,N_23837);
or UO_653 (O_653,N_24534,N_24879);
or UO_654 (O_654,N_24956,N_24611);
nor UO_655 (O_655,N_24192,N_24131);
and UO_656 (O_656,N_24650,N_24222);
or UO_657 (O_657,N_24636,N_24423);
xor UO_658 (O_658,N_24416,N_24332);
nor UO_659 (O_659,N_24309,N_24628);
nand UO_660 (O_660,N_23883,N_24188);
nor UO_661 (O_661,N_24624,N_24968);
or UO_662 (O_662,N_24804,N_24935);
or UO_663 (O_663,N_23806,N_24945);
nor UO_664 (O_664,N_24236,N_24934);
and UO_665 (O_665,N_24241,N_24759);
xnor UO_666 (O_666,N_23791,N_24169);
xor UO_667 (O_667,N_23884,N_24934);
nor UO_668 (O_668,N_24892,N_24017);
xor UO_669 (O_669,N_24644,N_24677);
or UO_670 (O_670,N_24379,N_24578);
or UO_671 (O_671,N_24908,N_24841);
and UO_672 (O_672,N_24368,N_24217);
xor UO_673 (O_673,N_24083,N_24983);
nor UO_674 (O_674,N_24638,N_24137);
and UO_675 (O_675,N_24459,N_24848);
or UO_676 (O_676,N_24511,N_23908);
and UO_677 (O_677,N_24010,N_24888);
or UO_678 (O_678,N_23804,N_23821);
xor UO_679 (O_679,N_24674,N_23816);
xnor UO_680 (O_680,N_23859,N_24131);
or UO_681 (O_681,N_24596,N_24762);
nand UO_682 (O_682,N_24802,N_24213);
and UO_683 (O_683,N_24868,N_24356);
nand UO_684 (O_684,N_24059,N_24856);
nor UO_685 (O_685,N_24975,N_24549);
or UO_686 (O_686,N_24887,N_24798);
nand UO_687 (O_687,N_23992,N_24940);
nor UO_688 (O_688,N_23882,N_24044);
and UO_689 (O_689,N_23841,N_24618);
or UO_690 (O_690,N_24735,N_24605);
and UO_691 (O_691,N_24260,N_24475);
xor UO_692 (O_692,N_23972,N_24594);
nor UO_693 (O_693,N_24825,N_24525);
nand UO_694 (O_694,N_24914,N_24086);
nand UO_695 (O_695,N_24420,N_23974);
nor UO_696 (O_696,N_23758,N_23890);
and UO_697 (O_697,N_24699,N_24057);
or UO_698 (O_698,N_24485,N_24428);
and UO_699 (O_699,N_24833,N_24107);
xnor UO_700 (O_700,N_24788,N_23826);
and UO_701 (O_701,N_24916,N_24157);
or UO_702 (O_702,N_24634,N_24179);
xnor UO_703 (O_703,N_24786,N_24288);
nand UO_704 (O_704,N_24976,N_24186);
xnor UO_705 (O_705,N_24434,N_23958);
nor UO_706 (O_706,N_24500,N_23754);
and UO_707 (O_707,N_24892,N_24609);
nor UO_708 (O_708,N_24798,N_24772);
nor UO_709 (O_709,N_24661,N_24817);
and UO_710 (O_710,N_24774,N_24479);
nand UO_711 (O_711,N_24549,N_24824);
xnor UO_712 (O_712,N_24942,N_24238);
and UO_713 (O_713,N_24458,N_24170);
xor UO_714 (O_714,N_24751,N_24157);
nand UO_715 (O_715,N_24872,N_24027);
xnor UO_716 (O_716,N_24664,N_24085);
and UO_717 (O_717,N_23838,N_24999);
xor UO_718 (O_718,N_24817,N_24176);
or UO_719 (O_719,N_24909,N_24741);
or UO_720 (O_720,N_24715,N_24780);
or UO_721 (O_721,N_23916,N_24782);
nor UO_722 (O_722,N_24446,N_24168);
nand UO_723 (O_723,N_24037,N_23766);
xor UO_724 (O_724,N_24424,N_24456);
or UO_725 (O_725,N_24130,N_24990);
xor UO_726 (O_726,N_24956,N_24907);
nor UO_727 (O_727,N_24329,N_23931);
xor UO_728 (O_728,N_23992,N_24442);
xor UO_729 (O_729,N_24967,N_24884);
and UO_730 (O_730,N_24680,N_23758);
xnor UO_731 (O_731,N_24400,N_23986);
xor UO_732 (O_732,N_23779,N_23947);
and UO_733 (O_733,N_24591,N_23958);
xnor UO_734 (O_734,N_24541,N_24620);
xor UO_735 (O_735,N_23808,N_24222);
xnor UO_736 (O_736,N_24123,N_24608);
nor UO_737 (O_737,N_24573,N_24281);
nor UO_738 (O_738,N_24194,N_23954);
nand UO_739 (O_739,N_24560,N_24537);
xor UO_740 (O_740,N_23790,N_24920);
and UO_741 (O_741,N_24569,N_23855);
nor UO_742 (O_742,N_24294,N_24813);
and UO_743 (O_743,N_23974,N_24050);
nor UO_744 (O_744,N_24276,N_23992);
and UO_745 (O_745,N_24122,N_24406);
nand UO_746 (O_746,N_24344,N_24780);
nor UO_747 (O_747,N_24228,N_24355);
or UO_748 (O_748,N_24930,N_24959);
xor UO_749 (O_749,N_24840,N_23756);
xor UO_750 (O_750,N_24121,N_23887);
or UO_751 (O_751,N_23934,N_24742);
nand UO_752 (O_752,N_24488,N_24145);
and UO_753 (O_753,N_23992,N_24535);
and UO_754 (O_754,N_24531,N_24677);
nor UO_755 (O_755,N_24351,N_23920);
nor UO_756 (O_756,N_24788,N_23801);
xor UO_757 (O_757,N_24635,N_24035);
nor UO_758 (O_758,N_23861,N_23944);
and UO_759 (O_759,N_24805,N_23885);
or UO_760 (O_760,N_23985,N_24564);
or UO_761 (O_761,N_24975,N_24217);
nand UO_762 (O_762,N_24231,N_24801);
nand UO_763 (O_763,N_24635,N_24070);
xor UO_764 (O_764,N_24482,N_24121);
xnor UO_765 (O_765,N_24461,N_24757);
and UO_766 (O_766,N_23872,N_23805);
and UO_767 (O_767,N_24383,N_24632);
xnor UO_768 (O_768,N_24311,N_24603);
nor UO_769 (O_769,N_23989,N_24199);
xnor UO_770 (O_770,N_24565,N_23978);
or UO_771 (O_771,N_24319,N_24042);
nor UO_772 (O_772,N_23897,N_23994);
nand UO_773 (O_773,N_24269,N_24246);
xnor UO_774 (O_774,N_24149,N_24260);
nand UO_775 (O_775,N_24218,N_24013);
xnor UO_776 (O_776,N_24775,N_24100);
nor UO_777 (O_777,N_24037,N_24077);
and UO_778 (O_778,N_24427,N_24580);
and UO_779 (O_779,N_24349,N_23821);
or UO_780 (O_780,N_24994,N_24772);
or UO_781 (O_781,N_24105,N_24025);
nor UO_782 (O_782,N_24832,N_23883);
xor UO_783 (O_783,N_24523,N_23836);
nor UO_784 (O_784,N_24058,N_24395);
xor UO_785 (O_785,N_24323,N_24766);
nor UO_786 (O_786,N_24603,N_24667);
xor UO_787 (O_787,N_24255,N_24101);
or UO_788 (O_788,N_23976,N_24263);
nor UO_789 (O_789,N_24653,N_24676);
nor UO_790 (O_790,N_24486,N_24806);
xor UO_791 (O_791,N_23871,N_24794);
or UO_792 (O_792,N_24310,N_24451);
or UO_793 (O_793,N_24333,N_24203);
or UO_794 (O_794,N_24804,N_24031);
xor UO_795 (O_795,N_24713,N_24782);
xor UO_796 (O_796,N_24514,N_24933);
or UO_797 (O_797,N_23960,N_24894);
and UO_798 (O_798,N_24865,N_24765);
nand UO_799 (O_799,N_24103,N_24956);
and UO_800 (O_800,N_24516,N_24780);
nand UO_801 (O_801,N_24609,N_24716);
nand UO_802 (O_802,N_24704,N_23762);
and UO_803 (O_803,N_24828,N_23949);
or UO_804 (O_804,N_24127,N_24179);
and UO_805 (O_805,N_24799,N_23807);
nor UO_806 (O_806,N_24646,N_24682);
or UO_807 (O_807,N_24355,N_23875);
nor UO_808 (O_808,N_24105,N_24240);
or UO_809 (O_809,N_24452,N_23850);
nand UO_810 (O_810,N_24236,N_23938);
or UO_811 (O_811,N_23759,N_24891);
nand UO_812 (O_812,N_24175,N_24871);
or UO_813 (O_813,N_24279,N_24823);
nor UO_814 (O_814,N_24875,N_24423);
or UO_815 (O_815,N_23828,N_24608);
nand UO_816 (O_816,N_24251,N_23929);
xor UO_817 (O_817,N_24736,N_24410);
nand UO_818 (O_818,N_24468,N_24647);
xor UO_819 (O_819,N_24776,N_23754);
and UO_820 (O_820,N_24317,N_24957);
nand UO_821 (O_821,N_23935,N_24663);
xnor UO_822 (O_822,N_24459,N_24688);
nand UO_823 (O_823,N_23797,N_23922);
and UO_824 (O_824,N_23784,N_24127);
nand UO_825 (O_825,N_23880,N_24684);
or UO_826 (O_826,N_24316,N_24479);
and UO_827 (O_827,N_24294,N_23852);
xnor UO_828 (O_828,N_24672,N_24626);
xor UO_829 (O_829,N_24043,N_23796);
nand UO_830 (O_830,N_24484,N_24861);
and UO_831 (O_831,N_24336,N_24396);
and UO_832 (O_832,N_24423,N_24018);
and UO_833 (O_833,N_24123,N_24340);
xnor UO_834 (O_834,N_23876,N_24202);
and UO_835 (O_835,N_24435,N_24764);
nor UO_836 (O_836,N_24037,N_24822);
xor UO_837 (O_837,N_24469,N_24905);
xor UO_838 (O_838,N_24884,N_24416);
nor UO_839 (O_839,N_24256,N_24478);
nor UO_840 (O_840,N_24008,N_23894);
or UO_841 (O_841,N_24427,N_23912);
or UO_842 (O_842,N_24124,N_24903);
nand UO_843 (O_843,N_24540,N_24004);
nand UO_844 (O_844,N_24109,N_24971);
and UO_845 (O_845,N_24103,N_24608);
xor UO_846 (O_846,N_24880,N_24824);
or UO_847 (O_847,N_24530,N_24060);
nand UO_848 (O_848,N_24541,N_24471);
or UO_849 (O_849,N_24524,N_24759);
nand UO_850 (O_850,N_24531,N_24775);
and UO_851 (O_851,N_24444,N_24883);
and UO_852 (O_852,N_23904,N_24148);
nor UO_853 (O_853,N_24032,N_24976);
xnor UO_854 (O_854,N_24943,N_24390);
and UO_855 (O_855,N_24015,N_23916);
nand UO_856 (O_856,N_24205,N_24398);
nor UO_857 (O_857,N_24258,N_24118);
nor UO_858 (O_858,N_23861,N_23858);
nand UO_859 (O_859,N_24551,N_24882);
nor UO_860 (O_860,N_24249,N_24885);
nand UO_861 (O_861,N_24690,N_24368);
xor UO_862 (O_862,N_24609,N_24976);
or UO_863 (O_863,N_24968,N_24938);
nand UO_864 (O_864,N_24177,N_24729);
nand UO_865 (O_865,N_24750,N_24152);
nor UO_866 (O_866,N_24231,N_23822);
and UO_867 (O_867,N_24357,N_24678);
nand UO_868 (O_868,N_24420,N_24306);
nor UO_869 (O_869,N_24159,N_24160);
or UO_870 (O_870,N_24094,N_24850);
xor UO_871 (O_871,N_24702,N_24326);
and UO_872 (O_872,N_24712,N_23891);
and UO_873 (O_873,N_24281,N_23754);
and UO_874 (O_874,N_24461,N_23765);
xnor UO_875 (O_875,N_24452,N_24480);
nor UO_876 (O_876,N_24013,N_24764);
xnor UO_877 (O_877,N_24754,N_24312);
and UO_878 (O_878,N_24983,N_24214);
nand UO_879 (O_879,N_24562,N_24165);
and UO_880 (O_880,N_24297,N_24446);
and UO_881 (O_881,N_24223,N_24987);
nor UO_882 (O_882,N_24770,N_24247);
nor UO_883 (O_883,N_23898,N_24362);
or UO_884 (O_884,N_24097,N_23951);
and UO_885 (O_885,N_24666,N_24507);
nor UO_886 (O_886,N_24335,N_23941);
xor UO_887 (O_887,N_23959,N_24792);
or UO_888 (O_888,N_24041,N_23973);
nor UO_889 (O_889,N_24285,N_24036);
xor UO_890 (O_890,N_24068,N_23768);
or UO_891 (O_891,N_24152,N_24700);
and UO_892 (O_892,N_23834,N_24231);
xnor UO_893 (O_893,N_24659,N_23926);
nand UO_894 (O_894,N_24673,N_24532);
xor UO_895 (O_895,N_24171,N_23996);
nand UO_896 (O_896,N_24636,N_24631);
xor UO_897 (O_897,N_24853,N_24076);
and UO_898 (O_898,N_24980,N_24174);
xor UO_899 (O_899,N_24730,N_24011);
nand UO_900 (O_900,N_24532,N_24716);
and UO_901 (O_901,N_24874,N_24767);
xnor UO_902 (O_902,N_24245,N_24757);
xor UO_903 (O_903,N_24892,N_24614);
and UO_904 (O_904,N_24643,N_24166);
or UO_905 (O_905,N_24447,N_24417);
nand UO_906 (O_906,N_23914,N_24931);
and UO_907 (O_907,N_24275,N_24492);
xnor UO_908 (O_908,N_23858,N_24276);
nor UO_909 (O_909,N_23879,N_24138);
nand UO_910 (O_910,N_24770,N_24978);
nor UO_911 (O_911,N_24421,N_23835);
or UO_912 (O_912,N_24887,N_24480);
or UO_913 (O_913,N_24543,N_24555);
and UO_914 (O_914,N_24364,N_23987);
nand UO_915 (O_915,N_23908,N_24840);
nor UO_916 (O_916,N_23771,N_24319);
nand UO_917 (O_917,N_23879,N_24948);
and UO_918 (O_918,N_23909,N_24914);
or UO_919 (O_919,N_24700,N_24510);
xnor UO_920 (O_920,N_24738,N_23793);
nor UO_921 (O_921,N_23891,N_24473);
and UO_922 (O_922,N_24194,N_23855);
or UO_923 (O_923,N_24161,N_24448);
nand UO_924 (O_924,N_24808,N_23997);
or UO_925 (O_925,N_24572,N_24214);
or UO_926 (O_926,N_24908,N_24226);
nand UO_927 (O_927,N_23900,N_24375);
nand UO_928 (O_928,N_24938,N_24435);
xnor UO_929 (O_929,N_23908,N_24829);
and UO_930 (O_930,N_24664,N_24333);
or UO_931 (O_931,N_24151,N_23972);
nor UO_932 (O_932,N_24005,N_24561);
nor UO_933 (O_933,N_24981,N_24629);
nor UO_934 (O_934,N_24532,N_23752);
and UO_935 (O_935,N_24737,N_23824);
and UO_936 (O_936,N_24150,N_24227);
or UO_937 (O_937,N_24958,N_24629);
nand UO_938 (O_938,N_24927,N_24187);
nor UO_939 (O_939,N_24452,N_24535);
or UO_940 (O_940,N_24790,N_24417);
or UO_941 (O_941,N_24351,N_23952);
or UO_942 (O_942,N_24663,N_24255);
nor UO_943 (O_943,N_24775,N_24356);
xor UO_944 (O_944,N_24187,N_23882);
nor UO_945 (O_945,N_23974,N_24552);
and UO_946 (O_946,N_24407,N_24964);
and UO_947 (O_947,N_23779,N_23996);
nor UO_948 (O_948,N_23993,N_24252);
nand UO_949 (O_949,N_24543,N_23754);
nand UO_950 (O_950,N_24261,N_23989);
nor UO_951 (O_951,N_24585,N_24320);
or UO_952 (O_952,N_24246,N_24359);
xnor UO_953 (O_953,N_24630,N_23908);
and UO_954 (O_954,N_24163,N_23930);
xnor UO_955 (O_955,N_23769,N_24294);
nand UO_956 (O_956,N_24819,N_24930);
or UO_957 (O_957,N_24067,N_24887);
nand UO_958 (O_958,N_24321,N_24626);
xor UO_959 (O_959,N_24662,N_24270);
xnor UO_960 (O_960,N_23795,N_23772);
xnor UO_961 (O_961,N_24711,N_24883);
nand UO_962 (O_962,N_23881,N_24244);
or UO_963 (O_963,N_24062,N_24944);
nor UO_964 (O_964,N_23755,N_24862);
xor UO_965 (O_965,N_24846,N_24087);
and UO_966 (O_966,N_23854,N_24510);
nand UO_967 (O_967,N_23999,N_23812);
nor UO_968 (O_968,N_24504,N_23855);
nor UO_969 (O_969,N_23908,N_24467);
nor UO_970 (O_970,N_24704,N_23925);
xnor UO_971 (O_971,N_24653,N_24575);
and UO_972 (O_972,N_24421,N_24369);
and UO_973 (O_973,N_23903,N_24716);
nor UO_974 (O_974,N_24337,N_24008);
and UO_975 (O_975,N_23801,N_23918);
nor UO_976 (O_976,N_24814,N_24753);
and UO_977 (O_977,N_24790,N_24193);
or UO_978 (O_978,N_24625,N_24812);
or UO_979 (O_979,N_24487,N_23914);
or UO_980 (O_980,N_24992,N_24474);
nand UO_981 (O_981,N_24260,N_24435);
and UO_982 (O_982,N_23998,N_24049);
or UO_983 (O_983,N_23771,N_24609);
nor UO_984 (O_984,N_24814,N_24635);
and UO_985 (O_985,N_23836,N_24182);
and UO_986 (O_986,N_24538,N_24473);
nand UO_987 (O_987,N_24006,N_24389);
or UO_988 (O_988,N_23771,N_24284);
nor UO_989 (O_989,N_24066,N_24393);
and UO_990 (O_990,N_24509,N_24787);
nor UO_991 (O_991,N_24482,N_24598);
and UO_992 (O_992,N_23934,N_24184);
xnor UO_993 (O_993,N_24071,N_24264);
nand UO_994 (O_994,N_24036,N_24030);
or UO_995 (O_995,N_24157,N_24874);
or UO_996 (O_996,N_24973,N_24057);
xnor UO_997 (O_997,N_24448,N_24837);
xnor UO_998 (O_998,N_23816,N_24937);
nor UO_999 (O_999,N_24274,N_24701);
or UO_1000 (O_1000,N_24856,N_24481);
and UO_1001 (O_1001,N_24435,N_23953);
nand UO_1002 (O_1002,N_24250,N_24162);
or UO_1003 (O_1003,N_24116,N_23859);
nand UO_1004 (O_1004,N_24752,N_24640);
nand UO_1005 (O_1005,N_23898,N_24325);
xnor UO_1006 (O_1006,N_24036,N_24352);
or UO_1007 (O_1007,N_23938,N_24111);
xor UO_1008 (O_1008,N_23963,N_24121);
and UO_1009 (O_1009,N_24671,N_24009);
or UO_1010 (O_1010,N_23764,N_24912);
or UO_1011 (O_1011,N_24807,N_23807);
or UO_1012 (O_1012,N_23777,N_24495);
nor UO_1013 (O_1013,N_24548,N_24240);
nand UO_1014 (O_1014,N_24276,N_23876);
nor UO_1015 (O_1015,N_23801,N_24584);
and UO_1016 (O_1016,N_24835,N_24357);
and UO_1017 (O_1017,N_23943,N_24003);
nor UO_1018 (O_1018,N_24685,N_24872);
xor UO_1019 (O_1019,N_23941,N_24186);
and UO_1020 (O_1020,N_24796,N_24314);
nand UO_1021 (O_1021,N_23926,N_24018);
nor UO_1022 (O_1022,N_23755,N_24934);
and UO_1023 (O_1023,N_24559,N_24522);
nor UO_1024 (O_1024,N_24467,N_24051);
and UO_1025 (O_1025,N_24632,N_24379);
nor UO_1026 (O_1026,N_24926,N_23801);
nor UO_1027 (O_1027,N_24935,N_24102);
xnor UO_1028 (O_1028,N_23891,N_23798);
nand UO_1029 (O_1029,N_24340,N_24212);
and UO_1030 (O_1030,N_24649,N_23904);
xor UO_1031 (O_1031,N_24523,N_24341);
and UO_1032 (O_1032,N_24582,N_24062);
or UO_1033 (O_1033,N_23993,N_24455);
and UO_1034 (O_1034,N_23774,N_24638);
nand UO_1035 (O_1035,N_24647,N_24859);
or UO_1036 (O_1036,N_24459,N_24199);
nor UO_1037 (O_1037,N_24848,N_24242);
nand UO_1038 (O_1038,N_24467,N_24359);
and UO_1039 (O_1039,N_24113,N_23791);
and UO_1040 (O_1040,N_24190,N_24111);
xnor UO_1041 (O_1041,N_24160,N_24228);
nor UO_1042 (O_1042,N_24489,N_24164);
xor UO_1043 (O_1043,N_23983,N_24067);
nand UO_1044 (O_1044,N_24583,N_23760);
nor UO_1045 (O_1045,N_24009,N_24950);
nor UO_1046 (O_1046,N_23797,N_24357);
or UO_1047 (O_1047,N_24363,N_24589);
nand UO_1048 (O_1048,N_23972,N_24035);
xor UO_1049 (O_1049,N_23822,N_24604);
or UO_1050 (O_1050,N_24302,N_24549);
or UO_1051 (O_1051,N_24347,N_24027);
xor UO_1052 (O_1052,N_24202,N_24143);
xnor UO_1053 (O_1053,N_24891,N_24476);
nand UO_1054 (O_1054,N_24122,N_24790);
xor UO_1055 (O_1055,N_24604,N_24702);
nand UO_1056 (O_1056,N_23966,N_24432);
nor UO_1057 (O_1057,N_24439,N_23968);
xor UO_1058 (O_1058,N_24797,N_24358);
nand UO_1059 (O_1059,N_24921,N_23865);
xnor UO_1060 (O_1060,N_24155,N_24920);
nand UO_1061 (O_1061,N_23934,N_23929);
and UO_1062 (O_1062,N_24999,N_24747);
nor UO_1063 (O_1063,N_23914,N_24833);
nor UO_1064 (O_1064,N_24373,N_24035);
and UO_1065 (O_1065,N_24161,N_24282);
xnor UO_1066 (O_1066,N_24210,N_24243);
xor UO_1067 (O_1067,N_24470,N_24444);
or UO_1068 (O_1068,N_23802,N_23965);
and UO_1069 (O_1069,N_23950,N_24710);
or UO_1070 (O_1070,N_23933,N_24922);
nor UO_1071 (O_1071,N_23893,N_24967);
nand UO_1072 (O_1072,N_24150,N_24790);
nor UO_1073 (O_1073,N_24061,N_24179);
xnor UO_1074 (O_1074,N_24390,N_24130);
or UO_1075 (O_1075,N_23807,N_24284);
xor UO_1076 (O_1076,N_24799,N_24806);
or UO_1077 (O_1077,N_24747,N_24457);
or UO_1078 (O_1078,N_23841,N_24101);
and UO_1079 (O_1079,N_24132,N_23770);
and UO_1080 (O_1080,N_24977,N_24514);
nand UO_1081 (O_1081,N_24216,N_24466);
nor UO_1082 (O_1082,N_24591,N_24285);
or UO_1083 (O_1083,N_24472,N_23852);
or UO_1084 (O_1084,N_23961,N_24770);
or UO_1085 (O_1085,N_24802,N_24109);
xnor UO_1086 (O_1086,N_24582,N_24607);
and UO_1087 (O_1087,N_24764,N_24137);
or UO_1088 (O_1088,N_24783,N_24909);
and UO_1089 (O_1089,N_24564,N_24289);
xnor UO_1090 (O_1090,N_24635,N_23805);
nor UO_1091 (O_1091,N_24104,N_23986);
nor UO_1092 (O_1092,N_24893,N_24486);
nand UO_1093 (O_1093,N_24927,N_24052);
and UO_1094 (O_1094,N_24530,N_23947);
nor UO_1095 (O_1095,N_24409,N_23866);
or UO_1096 (O_1096,N_23782,N_24740);
xor UO_1097 (O_1097,N_24984,N_24476);
or UO_1098 (O_1098,N_24033,N_24023);
nand UO_1099 (O_1099,N_24496,N_24392);
nand UO_1100 (O_1100,N_24269,N_24829);
nor UO_1101 (O_1101,N_23777,N_23898);
xor UO_1102 (O_1102,N_24953,N_24036);
xnor UO_1103 (O_1103,N_24593,N_24467);
nor UO_1104 (O_1104,N_24639,N_24533);
nor UO_1105 (O_1105,N_24206,N_24919);
xor UO_1106 (O_1106,N_24725,N_24479);
nand UO_1107 (O_1107,N_24386,N_24266);
and UO_1108 (O_1108,N_24853,N_23999);
nand UO_1109 (O_1109,N_24061,N_24708);
xor UO_1110 (O_1110,N_24680,N_23905);
xor UO_1111 (O_1111,N_24413,N_24540);
and UO_1112 (O_1112,N_24622,N_24142);
or UO_1113 (O_1113,N_24976,N_24268);
or UO_1114 (O_1114,N_24326,N_24560);
or UO_1115 (O_1115,N_24604,N_24631);
or UO_1116 (O_1116,N_24913,N_24138);
xnor UO_1117 (O_1117,N_24016,N_23808);
and UO_1118 (O_1118,N_24731,N_23973);
or UO_1119 (O_1119,N_24414,N_24547);
xor UO_1120 (O_1120,N_23989,N_23980);
nand UO_1121 (O_1121,N_24920,N_23813);
xnor UO_1122 (O_1122,N_24055,N_24516);
or UO_1123 (O_1123,N_24627,N_23813);
nor UO_1124 (O_1124,N_24145,N_24940);
nand UO_1125 (O_1125,N_24139,N_24535);
nor UO_1126 (O_1126,N_24162,N_23889);
xnor UO_1127 (O_1127,N_24817,N_24839);
xnor UO_1128 (O_1128,N_24116,N_24637);
nor UO_1129 (O_1129,N_23934,N_24005);
or UO_1130 (O_1130,N_23938,N_23929);
nand UO_1131 (O_1131,N_23988,N_24699);
nor UO_1132 (O_1132,N_24189,N_24394);
nor UO_1133 (O_1133,N_23880,N_24064);
nor UO_1134 (O_1134,N_24219,N_24398);
and UO_1135 (O_1135,N_24970,N_23979);
or UO_1136 (O_1136,N_24406,N_24744);
nor UO_1137 (O_1137,N_23964,N_24742);
or UO_1138 (O_1138,N_24919,N_24533);
nor UO_1139 (O_1139,N_23935,N_23799);
xor UO_1140 (O_1140,N_24771,N_23997);
nor UO_1141 (O_1141,N_24037,N_24808);
nand UO_1142 (O_1142,N_24679,N_24493);
or UO_1143 (O_1143,N_24519,N_23828);
xnor UO_1144 (O_1144,N_23914,N_24857);
and UO_1145 (O_1145,N_23932,N_24725);
or UO_1146 (O_1146,N_24409,N_24382);
nor UO_1147 (O_1147,N_24696,N_23824);
nor UO_1148 (O_1148,N_24738,N_24670);
nor UO_1149 (O_1149,N_23793,N_24751);
nand UO_1150 (O_1150,N_24222,N_24368);
xnor UO_1151 (O_1151,N_24006,N_24670);
xor UO_1152 (O_1152,N_23922,N_24542);
and UO_1153 (O_1153,N_23926,N_24012);
xor UO_1154 (O_1154,N_24231,N_24660);
and UO_1155 (O_1155,N_24750,N_23950);
and UO_1156 (O_1156,N_24110,N_23918);
and UO_1157 (O_1157,N_24184,N_24495);
nand UO_1158 (O_1158,N_23808,N_23765);
nor UO_1159 (O_1159,N_24949,N_24272);
xnor UO_1160 (O_1160,N_24507,N_24801);
nor UO_1161 (O_1161,N_24800,N_24486);
xor UO_1162 (O_1162,N_23802,N_24815);
and UO_1163 (O_1163,N_24536,N_24292);
or UO_1164 (O_1164,N_23984,N_24499);
xnor UO_1165 (O_1165,N_24873,N_24654);
nand UO_1166 (O_1166,N_24070,N_24293);
or UO_1167 (O_1167,N_23868,N_24100);
and UO_1168 (O_1168,N_24303,N_24070);
nor UO_1169 (O_1169,N_23780,N_24142);
and UO_1170 (O_1170,N_24745,N_23809);
xor UO_1171 (O_1171,N_24492,N_24566);
nor UO_1172 (O_1172,N_24442,N_24739);
or UO_1173 (O_1173,N_24378,N_24469);
nand UO_1174 (O_1174,N_24783,N_24945);
or UO_1175 (O_1175,N_24565,N_24774);
and UO_1176 (O_1176,N_24066,N_24719);
nor UO_1177 (O_1177,N_24639,N_24332);
nor UO_1178 (O_1178,N_24305,N_23809);
nand UO_1179 (O_1179,N_24922,N_23963);
nor UO_1180 (O_1180,N_24461,N_24568);
nor UO_1181 (O_1181,N_24709,N_24737);
nor UO_1182 (O_1182,N_24936,N_24694);
nand UO_1183 (O_1183,N_24741,N_24605);
xor UO_1184 (O_1184,N_23889,N_23856);
and UO_1185 (O_1185,N_24152,N_24341);
nand UO_1186 (O_1186,N_24670,N_24543);
nand UO_1187 (O_1187,N_24066,N_24688);
xor UO_1188 (O_1188,N_23901,N_24562);
nand UO_1189 (O_1189,N_24270,N_24189);
and UO_1190 (O_1190,N_24459,N_23807);
or UO_1191 (O_1191,N_24840,N_24167);
xnor UO_1192 (O_1192,N_23974,N_23803);
or UO_1193 (O_1193,N_24511,N_24347);
or UO_1194 (O_1194,N_24662,N_24371);
and UO_1195 (O_1195,N_24688,N_24235);
and UO_1196 (O_1196,N_24908,N_24079);
xnor UO_1197 (O_1197,N_24176,N_23791);
xor UO_1198 (O_1198,N_24014,N_23792);
xor UO_1199 (O_1199,N_23937,N_24852);
or UO_1200 (O_1200,N_23877,N_24326);
or UO_1201 (O_1201,N_24863,N_24251);
and UO_1202 (O_1202,N_24425,N_24160);
xor UO_1203 (O_1203,N_24965,N_24492);
xnor UO_1204 (O_1204,N_24994,N_24825);
xnor UO_1205 (O_1205,N_24641,N_24161);
nor UO_1206 (O_1206,N_24098,N_24133);
or UO_1207 (O_1207,N_24270,N_24480);
xnor UO_1208 (O_1208,N_23929,N_24443);
nor UO_1209 (O_1209,N_24948,N_23787);
and UO_1210 (O_1210,N_24679,N_23898);
xor UO_1211 (O_1211,N_23913,N_23965);
and UO_1212 (O_1212,N_24938,N_24794);
nor UO_1213 (O_1213,N_24210,N_24986);
and UO_1214 (O_1214,N_24767,N_24962);
xor UO_1215 (O_1215,N_24309,N_24797);
xor UO_1216 (O_1216,N_24163,N_24112);
nand UO_1217 (O_1217,N_24455,N_24268);
and UO_1218 (O_1218,N_24681,N_24665);
and UO_1219 (O_1219,N_24472,N_24975);
nor UO_1220 (O_1220,N_24817,N_23917);
and UO_1221 (O_1221,N_24050,N_23851);
xor UO_1222 (O_1222,N_24047,N_24752);
nand UO_1223 (O_1223,N_24245,N_23912);
nor UO_1224 (O_1224,N_24513,N_24299);
or UO_1225 (O_1225,N_24541,N_23873);
or UO_1226 (O_1226,N_24601,N_24768);
or UO_1227 (O_1227,N_24569,N_24677);
nand UO_1228 (O_1228,N_24483,N_23819);
nor UO_1229 (O_1229,N_24391,N_24372);
or UO_1230 (O_1230,N_24500,N_24311);
or UO_1231 (O_1231,N_24794,N_24017);
or UO_1232 (O_1232,N_24490,N_23903);
or UO_1233 (O_1233,N_23948,N_24043);
nor UO_1234 (O_1234,N_24386,N_24529);
and UO_1235 (O_1235,N_24422,N_24360);
and UO_1236 (O_1236,N_24910,N_23998);
or UO_1237 (O_1237,N_24644,N_23793);
nand UO_1238 (O_1238,N_24027,N_24742);
xnor UO_1239 (O_1239,N_24557,N_24546);
or UO_1240 (O_1240,N_24947,N_24346);
xor UO_1241 (O_1241,N_24254,N_24954);
xnor UO_1242 (O_1242,N_23974,N_24811);
or UO_1243 (O_1243,N_23805,N_24926);
xor UO_1244 (O_1244,N_24749,N_23932);
nor UO_1245 (O_1245,N_24043,N_24536);
nand UO_1246 (O_1246,N_24879,N_24483);
and UO_1247 (O_1247,N_24891,N_24163);
xor UO_1248 (O_1248,N_24877,N_24294);
xor UO_1249 (O_1249,N_24443,N_24712);
xnor UO_1250 (O_1250,N_24058,N_24639);
xnor UO_1251 (O_1251,N_23824,N_24668);
and UO_1252 (O_1252,N_24584,N_24963);
xnor UO_1253 (O_1253,N_23923,N_23758);
xnor UO_1254 (O_1254,N_24608,N_24676);
xor UO_1255 (O_1255,N_24190,N_23874);
or UO_1256 (O_1256,N_24344,N_24633);
xor UO_1257 (O_1257,N_23774,N_24853);
or UO_1258 (O_1258,N_24357,N_24296);
nand UO_1259 (O_1259,N_24090,N_24460);
and UO_1260 (O_1260,N_24419,N_24738);
xnor UO_1261 (O_1261,N_23810,N_24567);
nor UO_1262 (O_1262,N_23886,N_24026);
nor UO_1263 (O_1263,N_23846,N_24823);
nor UO_1264 (O_1264,N_23853,N_24340);
or UO_1265 (O_1265,N_24179,N_24454);
nand UO_1266 (O_1266,N_23750,N_24739);
xnor UO_1267 (O_1267,N_23901,N_24611);
or UO_1268 (O_1268,N_24597,N_24689);
or UO_1269 (O_1269,N_24974,N_24269);
nand UO_1270 (O_1270,N_24580,N_24950);
nand UO_1271 (O_1271,N_24618,N_23869);
or UO_1272 (O_1272,N_24783,N_24592);
or UO_1273 (O_1273,N_24683,N_23767);
and UO_1274 (O_1274,N_23928,N_24030);
or UO_1275 (O_1275,N_24398,N_24597);
nand UO_1276 (O_1276,N_24035,N_24727);
nor UO_1277 (O_1277,N_24984,N_23898);
xnor UO_1278 (O_1278,N_24891,N_24965);
and UO_1279 (O_1279,N_24202,N_24383);
or UO_1280 (O_1280,N_24551,N_24787);
and UO_1281 (O_1281,N_24217,N_23772);
nor UO_1282 (O_1282,N_24869,N_24781);
and UO_1283 (O_1283,N_23797,N_23933);
or UO_1284 (O_1284,N_24645,N_23971);
xor UO_1285 (O_1285,N_24419,N_24829);
nand UO_1286 (O_1286,N_24486,N_24590);
and UO_1287 (O_1287,N_24921,N_24399);
nand UO_1288 (O_1288,N_24115,N_24820);
xor UO_1289 (O_1289,N_24606,N_24098);
xor UO_1290 (O_1290,N_24380,N_23874);
xnor UO_1291 (O_1291,N_23750,N_24609);
nor UO_1292 (O_1292,N_24950,N_23935);
and UO_1293 (O_1293,N_24594,N_24063);
xnor UO_1294 (O_1294,N_24007,N_24954);
nand UO_1295 (O_1295,N_24127,N_23982);
and UO_1296 (O_1296,N_24237,N_24323);
nor UO_1297 (O_1297,N_24000,N_24567);
or UO_1298 (O_1298,N_24535,N_24817);
xnor UO_1299 (O_1299,N_24563,N_24735);
xnor UO_1300 (O_1300,N_24387,N_24577);
or UO_1301 (O_1301,N_23902,N_23935);
or UO_1302 (O_1302,N_23907,N_24604);
nand UO_1303 (O_1303,N_23807,N_24485);
or UO_1304 (O_1304,N_24107,N_24789);
or UO_1305 (O_1305,N_24938,N_24797);
or UO_1306 (O_1306,N_23789,N_23762);
xnor UO_1307 (O_1307,N_24582,N_24002);
or UO_1308 (O_1308,N_24784,N_24735);
or UO_1309 (O_1309,N_24926,N_24859);
and UO_1310 (O_1310,N_24163,N_23860);
or UO_1311 (O_1311,N_24283,N_24701);
xor UO_1312 (O_1312,N_24021,N_23774);
and UO_1313 (O_1313,N_24691,N_24529);
or UO_1314 (O_1314,N_23881,N_24741);
nand UO_1315 (O_1315,N_24087,N_24093);
or UO_1316 (O_1316,N_24180,N_24871);
xor UO_1317 (O_1317,N_24957,N_24239);
xnor UO_1318 (O_1318,N_24917,N_23824);
and UO_1319 (O_1319,N_24652,N_24587);
nor UO_1320 (O_1320,N_24494,N_24452);
xor UO_1321 (O_1321,N_24827,N_24772);
nand UO_1322 (O_1322,N_24385,N_24863);
nand UO_1323 (O_1323,N_24454,N_24887);
xor UO_1324 (O_1324,N_24693,N_24023);
nand UO_1325 (O_1325,N_24228,N_24768);
nand UO_1326 (O_1326,N_24280,N_24236);
nor UO_1327 (O_1327,N_23810,N_24986);
and UO_1328 (O_1328,N_23973,N_24461);
nand UO_1329 (O_1329,N_24336,N_24828);
nand UO_1330 (O_1330,N_24443,N_24439);
nor UO_1331 (O_1331,N_23865,N_24101);
xnor UO_1332 (O_1332,N_24821,N_24377);
xor UO_1333 (O_1333,N_24923,N_24873);
or UO_1334 (O_1334,N_24923,N_23884);
or UO_1335 (O_1335,N_24963,N_24474);
xnor UO_1336 (O_1336,N_24308,N_24645);
nor UO_1337 (O_1337,N_24471,N_24764);
nand UO_1338 (O_1338,N_24748,N_24475);
and UO_1339 (O_1339,N_23975,N_24326);
xnor UO_1340 (O_1340,N_24849,N_24138);
nand UO_1341 (O_1341,N_24912,N_24198);
nor UO_1342 (O_1342,N_24074,N_24734);
nor UO_1343 (O_1343,N_24480,N_24876);
and UO_1344 (O_1344,N_24224,N_24984);
nor UO_1345 (O_1345,N_24275,N_24791);
or UO_1346 (O_1346,N_24093,N_23823);
nor UO_1347 (O_1347,N_24220,N_24147);
nand UO_1348 (O_1348,N_23888,N_23770);
nor UO_1349 (O_1349,N_24377,N_23806);
xor UO_1350 (O_1350,N_24765,N_23920);
xor UO_1351 (O_1351,N_23760,N_24837);
and UO_1352 (O_1352,N_24584,N_23785);
or UO_1353 (O_1353,N_24823,N_23969);
nand UO_1354 (O_1354,N_24940,N_24169);
nor UO_1355 (O_1355,N_24473,N_24270);
nand UO_1356 (O_1356,N_23959,N_24145);
or UO_1357 (O_1357,N_24357,N_23957);
nor UO_1358 (O_1358,N_23981,N_23890);
or UO_1359 (O_1359,N_23942,N_24940);
or UO_1360 (O_1360,N_24930,N_23938);
xor UO_1361 (O_1361,N_24513,N_23908);
or UO_1362 (O_1362,N_23868,N_24356);
and UO_1363 (O_1363,N_24023,N_24489);
xnor UO_1364 (O_1364,N_24159,N_23906);
nor UO_1365 (O_1365,N_24747,N_23766);
and UO_1366 (O_1366,N_24947,N_24087);
nor UO_1367 (O_1367,N_24664,N_23989);
nor UO_1368 (O_1368,N_23924,N_24710);
nand UO_1369 (O_1369,N_23945,N_24657);
nand UO_1370 (O_1370,N_23791,N_24748);
nor UO_1371 (O_1371,N_24534,N_24108);
nand UO_1372 (O_1372,N_24894,N_23968);
nor UO_1373 (O_1373,N_24069,N_24198);
nand UO_1374 (O_1374,N_24430,N_24569);
nand UO_1375 (O_1375,N_24099,N_24519);
nand UO_1376 (O_1376,N_23868,N_24269);
nand UO_1377 (O_1377,N_24679,N_23868);
and UO_1378 (O_1378,N_24735,N_24926);
nor UO_1379 (O_1379,N_24585,N_23757);
nand UO_1380 (O_1380,N_24268,N_24913);
nor UO_1381 (O_1381,N_24221,N_24618);
nand UO_1382 (O_1382,N_24885,N_24052);
nand UO_1383 (O_1383,N_24033,N_23927);
or UO_1384 (O_1384,N_24811,N_23847);
nor UO_1385 (O_1385,N_24310,N_24519);
and UO_1386 (O_1386,N_24681,N_24045);
or UO_1387 (O_1387,N_24119,N_24720);
nand UO_1388 (O_1388,N_24566,N_24885);
nand UO_1389 (O_1389,N_24782,N_23984);
or UO_1390 (O_1390,N_24893,N_24414);
nor UO_1391 (O_1391,N_24964,N_24215);
and UO_1392 (O_1392,N_24327,N_24461);
nor UO_1393 (O_1393,N_24735,N_24690);
and UO_1394 (O_1394,N_24249,N_24991);
or UO_1395 (O_1395,N_24384,N_24685);
xnor UO_1396 (O_1396,N_24153,N_24962);
nor UO_1397 (O_1397,N_24284,N_24388);
nor UO_1398 (O_1398,N_24054,N_24518);
and UO_1399 (O_1399,N_24538,N_23983);
and UO_1400 (O_1400,N_24027,N_23869);
nand UO_1401 (O_1401,N_24884,N_24082);
nor UO_1402 (O_1402,N_24374,N_24750);
xor UO_1403 (O_1403,N_24966,N_24504);
nor UO_1404 (O_1404,N_23802,N_24542);
nand UO_1405 (O_1405,N_24002,N_24773);
xor UO_1406 (O_1406,N_24219,N_24270);
xnor UO_1407 (O_1407,N_23944,N_23919);
nand UO_1408 (O_1408,N_24545,N_24337);
and UO_1409 (O_1409,N_24191,N_24071);
nand UO_1410 (O_1410,N_24317,N_24717);
xor UO_1411 (O_1411,N_23847,N_23825);
or UO_1412 (O_1412,N_24183,N_24345);
and UO_1413 (O_1413,N_24854,N_23823);
nand UO_1414 (O_1414,N_24247,N_24854);
nor UO_1415 (O_1415,N_24818,N_24767);
and UO_1416 (O_1416,N_24613,N_24689);
nand UO_1417 (O_1417,N_24145,N_24329);
and UO_1418 (O_1418,N_24673,N_24479);
nor UO_1419 (O_1419,N_24381,N_24940);
nor UO_1420 (O_1420,N_24637,N_24587);
nand UO_1421 (O_1421,N_23769,N_24596);
nand UO_1422 (O_1422,N_23858,N_23796);
and UO_1423 (O_1423,N_24760,N_24172);
and UO_1424 (O_1424,N_23907,N_23882);
xnor UO_1425 (O_1425,N_24209,N_23770);
and UO_1426 (O_1426,N_24389,N_24747);
xnor UO_1427 (O_1427,N_24451,N_24167);
nand UO_1428 (O_1428,N_24857,N_24145);
nand UO_1429 (O_1429,N_23981,N_23781);
nand UO_1430 (O_1430,N_24388,N_24746);
nor UO_1431 (O_1431,N_24371,N_23807);
nor UO_1432 (O_1432,N_24228,N_24960);
nand UO_1433 (O_1433,N_24449,N_23827);
and UO_1434 (O_1434,N_24171,N_24160);
xor UO_1435 (O_1435,N_24095,N_24839);
nand UO_1436 (O_1436,N_24849,N_24076);
or UO_1437 (O_1437,N_24451,N_24258);
nand UO_1438 (O_1438,N_24504,N_24434);
nor UO_1439 (O_1439,N_24795,N_24523);
or UO_1440 (O_1440,N_23888,N_24763);
nor UO_1441 (O_1441,N_23981,N_24416);
nand UO_1442 (O_1442,N_23944,N_24637);
nor UO_1443 (O_1443,N_24731,N_24363);
xnor UO_1444 (O_1444,N_24321,N_24738);
nor UO_1445 (O_1445,N_24705,N_24727);
nand UO_1446 (O_1446,N_24429,N_24755);
or UO_1447 (O_1447,N_24200,N_24982);
nor UO_1448 (O_1448,N_23906,N_24661);
and UO_1449 (O_1449,N_24859,N_23771);
nor UO_1450 (O_1450,N_24453,N_24315);
xor UO_1451 (O_1451,N_24190,N_24172);
and UO_1452 (O_1452,N_23975,N_23859);
xor UO_1453 (O_1453,N_24611,N_23895);
xnor UO_1454 (O_1454,N_24776,N_24837);
nand UO_1455 (O_1455,N_24484,N_24610);
xor UO_1456 (O_1456,N_24059,N_24009);
nor UO_1457 (O_1457,N_24009,N_23857);
xnor UO_1458 (O_1458,N_24402,N_24296);
xor UO_1459 (O_1459,N_24951,N_24613);
nor UO_1460 (O_1460,N_24579,N_24112);
xnor UO_1461 (O_1461,N_24141,N_24184);
xnor UO_1462 (O_1462,N_24064,N_24488);
or UO_1463 (O_1463,N_24032,N_23957);
nor UO_1464 (O_1464,N_24452,N_24774);
xnor UO_1465 (O_1465,N_24776,N_24294);
xor UO_1466 (O_1466,N_24017,N_23968);
nor UO_1467 (O_1467,N_24102,N_24604);
and UO_1468 (O_1468,N_23849,N_24749);
nand UO_1469 (O_1469,N_24719,N_24548);
nor UO_1470 (O_1470,N_23974,N_24194);
and UO_1471 (O_1471,N_23974,N_24232);
nor UO_1472 (O_1472,N_23792,N_24545);
nor UO_1473 (O_1473,N_23756,N_24366);
nand UO_1474 (O_1474,N_24309,N_24629);
xor UO_1475 (O_1475,N_23873,N_24995);
and UO_1476 (O_1476,N_24522,N_23932);
xnor UO_1477 (O_1477,N_23997,N_24856);
nor UO_1478 (O_1478,N_24403,N_24890);
nand UO_1479 (O_1479,N_24422,N_23996);
nor UO_1480 (O_1480,N_24656,N_24435);
or UO_1481 (O_1481,N_23773,N_24921);
or UO_1482 (O_1482,N_24888,N_23852);
nor UO_1483 (O_1483,N_23869,N_24187);
nand UO_1484 (O_1484,N_24058,N_23755);
nor UO_1485 (O_1485,N_24102,N_24612);
nor UO_1486 (O_1486,N_24861,N_24698);
nor UO_1487 (O_1487,N_24925,N_23761);
or UO_1488 (O_1488,N_24821,N_23961);
and UO_1489 (O_1489,N_24423,N_24509);
nor UO_1490 (O_1490,N_24864,N_24316);
nor UO_1491 (O_1491,N_24401,N_23830);
and UO_1492 (O_1492,N_24763,N_24640);
nand UO_1493 (O_1493,N_24068,N_24099);
or UO_1494 (O_1494,N_24577,N_23892);
nor UO_1495 (O_1495,N_23939,N_24451);
nand UO_1496 (O_1496,N_24599,N_24004);
and UO_1497 (O_1497,N_24251,N_24912);
nor UO_1498 (O_1498,N_24174,N_23888);
or UO_1499 (O_1499,N_24457,N_24167);
xor UO_1500 (O_1500,N_24495,N_24734);
and UO_1501 (O_1501,N_24651,N_24454);
nor UO_1502 (O_1502,N_24211,N_24162);
nand UO_1503 (O_1503,N_24561,N_24148);
xnor UO_1504 (O_1504,N_24759,N_24713);
nor UO_1505 (O_1505,N_24641,N_24863);
and UO_1506 (O_1506,N_24795,N_23825);
xor UO_1507 (O_1507,N_24499,N_24612);
and UO_1508 (O_1508,N_23913,N_24044);
or UO_1509 (O_1509,N_24726,N_23795);
or UO_1510 (O_1510,N_24834,N_24923);
and UO_1511 (O_1511,N_24783,N_24271);
xnor UO_1512 (O_1512,N_24615,N_24183);
nor UO_1513 (O_1513,N_24228,N_24930);
and UO_1514 (O_1514,N_23886,N_24966);
or UO_1515 (O_1515,N_23846,N_24191);
and UO_1516 (O_1516,N_24558,N_23780);
xor UO_1517 (O_1517,N_24555,N_24375);
xnor UO_1518 (O_1518,N_23952,N_24074);
nor UO_1519 (O_1519,N_23968,N_24618);
and UO_1520 (O_1520,N_24144,N_24426);
xor UO_1521 (O_1521,N_23760,N_24153);
nor UO_1522 (O_1522,N_24577,N_24297);
nand UO_1523 (O_1523,N_24801,N_23834);
nor UO_1524 (O_1524,N_23795,N_24497);
or UO_1525 (O_1525,N_24156,N_24687);
nand UO_1526 (O_1526,N_24103,N_24421);
nor UO_1527 (O_1527,N_24794,N_24035);
or UO_1528 (O_1528,N_24702,N_24916);
and UO_1529 (O_1529,N_24766,N_24528);
nand UO_1530 (O_1530,N_24518,N_24074);
and UO_1531 (O_1531,N_23791,N_24751);
nand UO_1532 (O_1532,N_24612,N_23823);
nor UO_1533 (O_1533,N_23842,N_24558);
nor UO_1534 (O_1534,N_24529,N_24249);
and UO_1535 (O_1535,N_24209,N_24896);
or UO_1536 (O_1536,N_24607,N_24815);
nand UO_1537 (O_1537,N_23849,N_23871);
xor UO_1538 (O_1538,N_24799,N_24586);
nor UO_1539 (O_1539,N_24204,N_24876);
nand UO_1540 (O_1540,N_24359,N_23967);
or UO_1541 (O_1541,N_24489,N_24274);
or UO_1542 (O_1542,N_24591,N_24670);
and UO_1543 (O_1543,N_24891,N_23792);
and UO_1544 (O_1544,N_24990,N_24054);
nand UO_1545 (O_1545,N_24871,N_23973);
and UO_1546 (O_1546,N_24211,N_23951);
nand UO_1547 (O_1547,N_24372,N_23792);
or UO_1548 (O_1548,N_24893,N_24307);
xnor UO_1549 (O_1549,N_24983,N_24598);
nand UO_1550 (O_1550,N_24214,N_24972);
or UO_1551 (O_1551,N_24435,N_24151);
nor UO_1552 (O_1552,N_23888,N_24689);
and UO_1553 (O_1553,N_23763,N_24403);
nor UO_1554 (O_1554,N_24819,N_24063);
nor UO_1555 (O_1555,N_24015,N_24047);
and UO_1556 (O_1556,N_24446,N_23838);
xor UO_1557 (O_1557,N_24401,N_24428);
nor UO_1558 (O_1558,N_23950,N_24910);
and UO_1559 (O_1559,N_24605,N_24300);
xnor UO_1560 (O_1560,N_24172,N_24979);
nor UO_1561 (O_1561,N_24712,N_24728);
nor UO_1562 (O_1562,N_24437,N_24865);
xnor UO_1563 (O_1563,N_24541,N_24970);
xnor UO_1564 (O_1564,N_24489,N_24352);
and UO_1565 (O_1565,N_24768,N_24659);
nor UO_1566 (O_1566,N_24498,N_23862);
nor UO_1567 (O_1567,N_24807,N_24401);
or UO_1568 (O_1568,N_23806,N_24170);
xor UO_1569 (O_1569,N_24996,N_24486);
xnor UO_1570 (O_1570,N_24076,N_24789);
nor UO_1571 (O_1571,N_24397,N_24658);
nor UO_1572 (O_1572,N_23854,N_23914);
or UO_1573 (O_1573,N_24953,N_24183);
nand UO_1574 (O_1574,N_24674,N_24402);
xor UO_1575 (O_1575,N_24196,N_23783);
nand UO_1576 (O_1576,N_24411,N_24898);
nor UO_1577 (O_1577,N_24808,N_24182);
and UO_1578 (O_1578,N_23995,N_24633);
and UO_1579 (O_1579,N_24180,N_24953);
nand UO_1580 (O_1580,N_23927,N_24073);
xor UO_1581 (O_1581,N_23842,N_23827);
nand UO_1582 (O_1582,N_24504,N_24878);
nor UO_1583 (O_1583,N_24132,N_24954);
or UO_1584 (O_1584,N_24738,N_24923);
xnor UO_1585 (O_1585,N_24382,N_24270);
xor UO_1586 (O_1586,N_24562,N_24523);
nand UO_1587 (O_1587,N_23847,N_23879);
or UO_1588 (O_1588,N_24510,N_23964);
nand UO_1589 (O_1589,N_23856,N_24244);
or UO_1590 (O_1590,N_24953,N_24627);
and UO_1591 (O_1591,N_24103,N_24911);
or UO_1592 (O_1592,N_24120,N_24070);
or UO_1593 (O_1593,N_23919,N_24086);
xnor UO_1594 (O_1594,N_24670,N_24057);
or UO_1595 (O_1595,N_24013,N_24724);
xor UO_1596 (O_1596,N_24232,N_24233);
and UO_1597 (O_1597,N_24002,N_24116);
or UO_1598 (O_1598,N_23942,N_24182);
or UO_1599 (O_1599,N_24374,N_23868);
xnor UO_1600 (O_1600,N_24205,N_24182);
xor UO_1601 (O_1601,N_24322,N_24246);
xor UO_1602 (O_1602,N_23993,N_23843);
xor UO_1603 (O_1603,N_24349,N_23928);
or UO_1604 (O_1604,N_24956,N_24934);
nor UO_1605 (O_1605,N_24836,N_24035);
nor UO_1606 (O_1606,N_24652,N_24116);
nand UO_1607 (O_1607,N_23822,N_24764);
and UO_1608 (O_1608,N_24061,N_23755);
and UO_1609 (O_1609,N_24119,N_24057);
xor UO_1610 (O_1610,N_24887,N_24337);
or UO_1611 (O_1611,N_24087,N_24318);
nor UO_1612 (O_1612,N_24849,N_24118);
nor UO_1613 (O_1613,N_24236,N_24034);
or UO_1614 (O_1614,N_23898,N_24427);
xor UO_1615 (O_1615,N_23940,N_24324);
or UO_1616 (O_1616,N_23833,N_24521);
xnor UO_1617 (O_1617,N_24010,N_24490);
or UO_1618 (O_1618,N_24975,N_24505);
xor UO_1619 (O_1619,N_24831,N_23988);
xnor UO_1620 (O_1620,N_23970,N_24725);
or UO_1621 (O_1621,N_24239,N_24561);
or UO_1622 (O_1622,N_24519,N_24381);
xnor UO_1623 (O_1623,N_24479,N_24910);
nand UO_1624 (O_1624,N_24078,N_24256);
nand UO_1625 (O_1625,N_24222,N_23862);
nor UO_1626 (O_1626,N_24434,N_24222);
nand UO_1627 (O_1627,N_24508,N_23961);
xor UO_1628 (O_1628,N_24327,N_24653);
xor UO_1629 (O_1629,N_23901,N_24747);
nand UO_1630 (O_1630,N_24098,N_24022);
and UO_1631 (O_1631,N_24044,N_24409);
or UO_1632 (O_1632,N_24782,N_24669);
xor UO_1633 (O_1633,N_24865,N_24575);
or UO_1634 (O_1634,N_24245,N_24555);
nor UO_1635 (O_1635,N_24226,N_24645);
xor UO_1636 (O_1636,N_24114,N_24750);
nand UO_1637 (O_1637,N_23853,N_24201);
nand UO_1638 (O_1638,N_24177,N_24267);
or UO_1639 (O_1639,N_23794,N_24759);
nand UO_1640 (O_1640,N_24956,N_24412);
and UO_1641 (O_1641,N_23830,N_24930);
nor UO_1642 (O_1642,N_24395,N_24100);
and UO_1643 (O_1643,N_23928,N_23866);
and UO_1644 (O_1644,N_24793,N_24387);
nor UO_1645 (O_1645,N_24630,N_24470);
xnor UO_1646 (O_1646,N_23870,N_24414);
nor UO_1647 (O_1647,N_24475,N_24709);
xnor UO_1648 (O_1648,N_24282,N_24399);
and UO_1649 (O_1649,N_24624,N_23764);
nor UO_1650 (O_1650,N_24134,N_24702);
nor UO_1651 (O_1651,N_24878,N_24478);
or UO_1652 (O_1652,N_24503,N_24823);
nor UO_1653 (O_1653,N_24702,N_24644);
xnor UO_1654 (O_1654,N_24327,N_24695);
xor UO_1655 (O_1655,N_24779,N_24207);
and UO_1656 (O_1656,N_23911,N_24193);
nand UO_1657 (O_1657,N_24744,N_23752);
and UO_1658 (O_1658,N_24717,N_24563);
and UO_1659 (O_1659,N_24933,N_24503);
or UO_1660 (O_1660,N_24366,N_24083);
nor UO_1661 (O_1661,N_24125,N_24650);
or UO_1662 (O_1662,N_24991,N_24414);
xor UO_1663 (O_1663,N_24692,N_24648);
nor UO_1664 (O_1664,N_24945,N_24684);
nand UO_1665 (O_1665,N_23862,N_24907);
and UO_1666 (O_1666,N_24224,N_23924);
nor UO_1667 (O_1667,N_23806,N_24542);
and UO_1668 (O_1668,N_24787,N_24276);
nand UO_1669 (O_1669,N_24704,N_23822);
nand UO_1670 (O_1670,N_24961,N_23804);
and UO_1671 (O_1671,N_24374,N_24978);
nor UO_1672 (O_1672,N_24953,N_24857);
or UO_1673 (O_1673,N_24073,N_24924);
or UO_1674 (O_1674,N_24803,N_24440);
nor UO_1675 (O_1675,N_23752,N_23889);
xnor UO_1676 (O_1676,N_23775,N_24828);
and UO_1677 (O_1677,N_24981,N_24847);
nand UO_1678 (O_1678,N_24851,N_24313);
nand UO_1679 (O_1679,N_24092,N_24917);
or UO_1680 (O_1680,N_24390,N_24090);
or UO_1681 (O_1681,N_24793,N_24629);
nand UO_1682 (O_1682,N_24558,N_24633);
nor UO_1683 (O_1683,N_24883,N_24458);
or UO_1684 (O_1684,N_24607,N_24183);
and UO_1685 (O_1685,N_23933,N_24153);
or UO_1686 (O_1686,N_24809,N_24118);
nor UO_1687 (O_1687,N_24501,N_24683);
and UO_1688 (O_1688,N_24600,N_24870);
xor UO_1689 (O_1689,N_24661,N_24415);
or UO_1690 (O_1690,N_24059,N_23860);
nor UO_1691 (O_1691,N_24763,N_24930);
and UO_1692 (O_1692,N_24315,N_24254);
xor UO_1693 (O_1693,N_23844,N_24856);
nor UO_1694 (O_1694,N_24122,N_24167);
nand UO_1695 (O_1695,N_24011,N_24787);
and UO_1696 (O_1696,N_24521,N_24759);
and UO_1697 (O_1697,N_23750,N_24997);
and UO_1698 (O_1698,N_24896,N_24648);
or UO_1699 (O_1699,N_24116,N_23817);
nand UO_1700 (O_1700,N_24971,N_24750);
nand UO_1701 (O_1701,N_24795,N_24868);
and UO_1702 (O_1702,N_24600,N_24851);
and UO_1703 (O_1703,N_23839,N_24075);
or UO_1704 (O_1704,N_24188,N_24151);
or UO_1705 (O_1705,N_24083,N_24954);
xor UO_1706 (O_1706,N_24268,N_23962);
xnor UO_1707 (O_1707,N_24353,N_24893);
or UO_1708 (O_1708,N_24334,N_24521);
and UO_1709 (O_1709,N_24386,N_24060);
xor UO_1710 (O_1710,N_24822,N_24171);
xor UO_1711 (O_1711,N_24137,N_23955);
or UO_1712 (O_1712,N_24829,N_23950);
nor UO_1713 (O_1713,N_24435,N_23867);
and UO_1714 (O_1714,N_24217,N_24331);
nand UO_1715 (O_1715,N_24066,N_24341);
nand UO_1716 (O_1716,N_24475,N_23835);
nand UO_1717 (O_1717,N_23823,N_24267);
and UO_1718 (O_1718,N_24298,N_24951);
and UO_1719 (O_1719,N_23972,N_24421);
or UO_1720 (O_1720,N_24723,N_23798);
xnor UO_1721 (O_1721,N_24318,N_24127);
nand UO_1722 (O_1722,N_24626,N_24345);
nor UO_1723 (O_1723,N_24668,N_24504);
nor UO_1724 (O_1724,N_24423,N_24083);
nor UO_1725 (O_1725,N_24766,N_24652);
nand UO_1726 (O_1726,N_24858,N_24773);
or UO_1727 (O_1727,N_24473,N_24711);
and UO_1728 (O_1728,N_24419,N_24741);
and UO_1729 (O_1729,N_24306,N_24864);
and UO_1730 (O_1730,N_24920,N_24216);
or UO_1731 (O_1731,N_23753,N_23811);
and UO_1732 (O_1732,N_24947,N_23759);
nand UO_1733 (O_1733,N_24896,N_24490);
xnor UO_1734 (O_1734,N_24944,N_24648);
or UO_1735 (O_1735,N_23878,N_24766);
xnor UO_1736 (O_1736,N_24929,N_24577);
nand UO_1737 (O_1737,N_23911,N_24229);
nor UO_1738 (O_1738,N_24161,N_24621);
and UO_1739 (O_1739,N_24663,N_24891);
or UO_1740 (O_1740,N_24309,N_24455);
xnor UO_1741 (O_1741,N_24156,N_24328);
nand UO_1742 (O_1742,N_24232,N_24620);
or UO_1743 (O_1743,N_23926,N_24692);
and UO_1744 (O_1744,N_24222,N_24230);
and UO_1745 (O_1745,N_24565,N_24766);
nand UO_1746 (O_1746,N_24719,N_23825);
or UO_1747 (O_1747,N_24361,N_23970);
nor UO_1748 (O_1748,N_24119,N_24174);
nor UO_1749 (O_1749,N_24688,N_24281);
nand UO_1750 (O_1750,N_24630,N_24738);
nor UO_1751 (O_1751,N_24640,N_24901);
nand UO_1752 (O_1752,N_24333,N_23958);
nor UO_1753 (O_1753,N_23854,N_23935);
nor UO_1754 (O_1754,N_24206,N_24621);
or UO_1755 (O_1755,N_24711,N_23799);
nand UO_1756 (O_1756,N_24604,N_24100);
and UO_1757 (O_1757,N_24429,N_24365);
nor UO_1758 (O_1758,N_24113,N_24535);
nand UO_1759 (O_1759,N_24097,N_24937);
nor UO_1760 (O_1760,N_24077,N_24687);
or UO_1761 (O_1761,N_24716,N_24552);
nor UO_1762 (O_1762,N_24715,N_23942);
or UO_1763 (O_1763,N_24747,N_24815);
or UO_1764 (O_1764,N_24274,N_24432);
and UO_1765 (O_1765,N_24444,N_24696);
nor UO_1766 (O_1766,N_23782,N_24869);
and UO_1767 (O_1767,N_24085,N_24047);
and UO_1768 (O_1768,N_24156,N_24894);
and UO_1769 (O_1769,N_24730,N_23761);
nand UO_1770 (O_1770,N_24648,N_24379);
xnor UO_1771 (O_1771,N_23773,N_24039);
xnor UO_1772 (O_1772,N_24337,N_23898);
and UO_1773 (O_1773,N_24704,N_24154);
nor UO_1774 (O_1774,N_23810,N_24514);
nor UO_1775 (O_1775,N_24332,N_24696);
nor UO_1776 (O_1776,N_23813,N_23879);
and UO_1777 (O_1777,N_24340,N_24823);
or UO_1778 (O_1778,N_24254,N_23999);
or UO_1779 (O_1779,N_24593,N_24753);
or UO_1780 (O_1780,N_24531,N_23942);
or UO_1781 (O_1781,N_24303,N_23947);
and UO_1782 (O_1782,N_23813,N_24743);
nor UO_1783 (O_1783,N_23939,N_24181);
nand UO_1784 (O_1784,N_23776,N_24083);
or UO_1785 (O_1785,N_24360,N_24237);
nor UO_1786 (O_1786,N_24744,N_24354);
nand UO_1787 (O_1787,N_24184,N_24388);
and UO_1788 (O_1788,N_23782,N_24078);
nand UO_1789 (O_1789,N_24338,N_23992);
nor UO_1790 (O_1790,N_23818,N_24899);
nor UO_1791 (O_1791,N_24589,N_23841);
and UO_1792 (O_1792,N_24721,N_23970);
or UO_1793 (O_1793,N_24007,N_24803);
nor UO_1794 (O_1794,N_24720,N_24574);
and UO_1795 (O_1795,N_23917,N_23942);
or UO_1796 (O_1796,N_24709,N_24094);
nand UO_1797 (O_1797,N_24098,N_23855);
or UO_1798 (O_1798,N_23774,N_24476);
nor UO_1799 (O_1799,N_23958,N_24964);
nor UO_1800 (O_1800,N_23881,N_23835);
nor UO_1801 (O_1801,N_24484,N_24860);
nand UO_1802 (O_1802,N_23759,N_24140);
or UO_1803 (O_1803,N_24404,N_23983);
xor UO_1804 (O_1804,N_24470,N_24162);
or UO_1805 (O_1805,N_24912,N_23833);
nand UO_1806 (O_1806,N_24854,N_24990);
xor UO_1807 (O_1807,N_24857,N_24527);
nor UO_1808 (O_1808,N_24138,N_24872);
or UO_1809 (O_1809,N_24183,N_24257);
xor UO_1810 (O_1810,N_24486,N_24498);
and UO_1811 (O_1811,N_24460,N_24202);
nand UO_1812 (O_1812,N_23814,N_23811);
and UO_1813 (O_1813,N_24501,N_24760);
nor UO_1814 (O_1814,N_24243,N_24872);
xor UO_1815 (O_1815,N_24480,N_24645);
xnor UO_1816 (O_1816,N_23982,N_24076);
and UO_1817 (O_1817,N_24172,N_24378);
nor UO_1818 (O_1818,N_24035,N_23985);
nor UO_1819 (O_1819,N_24735,N_24739);
xnor UO_1820 (O_1820,N_23907,N_24696);
nand UO_1821 (O_1821,N_24196,N_24756);
or UO_1822 (O_1822,N_24939,N_24333);
nor UO_1823 (O_1823,N_24049,N_24070);
or UO_1824 (O_1824,N_23893,N_24608);
or UO_1825 (O_1825,N_24614,N_24013);
and UO_1826 (O_1826,N_23801,N_24976);
and UO_1827 (O_1827,N_24927,N_23823);
nor UO_1828 (O_1828,N_24697,N_24588);
xor UO_1829 (O_1829,N_24726,N_24813);
and UO_1830 (O_1830,N_24108,N_24702);
and UO_1831 (O_1831,N_24710,N_24443);
or UO_1832 (O_1832,N_23835,N_24518);
nor UO_1833 (O_1833,N_23774,N_24198);
xor UO_1834 (O_1834,N_24868,N_24023);
and UO_1835 (O_1835,N_24820,N_24392);
or UO_1836 (O_1836,N_24574,N_24157);
or UO_1837 (O_1837,N_24226,N_23918);
and UO_1838 (O_1838,N_24414,N_23992);
xor UO_1839 (O_1839,N_24330,N_24381);
xnor UO_1840 (O_1840,N_24223,N_24972);
and UO_1841 (O_1841,N_23877,N_24451);
or UO_1842 (O_1842,N_24082,N_24299);
nor UO_1843 (O_1843,N_24953,N_24886);
xor UO_1844 (O_1844,N_24982,N_24208);
nor UO_1845 (O_1845,N_24028,N_24317);
and UO_1846 (O_1846,N_24021,N_24114);
nand UO_1847 (O_1847,N_24974,N_24653);
nor UO_1848 (O_1848,N_23926,N_24619);
xor UO_1849 (O_1849,N_24115,N_24408);
and UO_1850 (O_1850,N_24513,N_24489);
and UO_1851 (O_1851,N_23926,N_24208);
or UO_1852 (O_1852,N_24261,N_24455);
xor UO_1853 (O_1853,N_24751,N_24242);
xor UO_1854 (O_1854,N_24635,N_24561);
xor UO_1855 (O_1855,N_24338,N_24868);
nand UO_1856 (O_1856,N_23906,N_24934);
and UO_1857 (O_1857,N_24921,N_24069);
nor UO_1858 (O_1858,N_24183,N_24403);
nor UO_1859 (O_1859,N_24578,N_24347);
nand UO_1860 (O_1860,N_23785,N_23759);
nand UO_1861 (O_1861,N_24726,N_24840);
and UO_1862 (O_1862,N_23837,N_24564);
or UO_1863 (O_1863,N_23983,N_23825);
or UO_1864 (O_1864,N_24914,N_24370);
and UO_1865 (O_1865,N_24801,N_24293);
and UO_1866 (O_1866,N_24336,N_24446);
or UO_1867 (O_1867,N_24420,N_24916);
or UO_1868 (O_1868,N_24376,N_24491);
xnor UO_1869 (O_1869,N_23989,N_24735);
nor UO_1870 (O_1870,N_24261,N_24794);
xor UO_1871 (O_1871,N_24561,N_24912);
nor UO_1872 (O_1872,N_24266,N_24686);
or UO_1873 (O_1873,N_24379,N_24179);
xnor UO_1874 (O_1874,N_24654,N_23961);
or UO_1875 (O_1875,N_24446,N_24482);
or UO_1876 (O_1876,N_24113,N_24396);
and UO_1877 (O_1877,N_24104,N_24041);
or UO_1878 (O_1878,N_24739,N_23833);
and UO_1879 (O_1879,N_24841,N_24164);
nor UO_1880 (O_1880,N_24793,N_24267);
and UO_1881 (O_1881,N_24658,N_24900);
xnor UO_1882 (O_1882,N_24954,N_24142);
nor UO_1883 (O_1883,N_24449,N_23844);
or UO_1884 (O_1884,N_24510,N_23973);
xor UO_1885 (O_1885,N_24523,N_24349);
or UO_1886 (O_1886,N_24776,N_24802);
and UO_1887 (O_1887,N_23795,N_23805);
nor UO_1888 (O_1888,N_24960,N_24596);
nor UO_1889 (O_1889,N_24290,N_24180);
and UO_1890 (O_1890,N_24554,N_24328);
xnor UO_1891 (O_1891,N_24381,N_24690);
nor UO_1892 (O_1892,N_24466,N_23958);
and UO_1893 (O_1893,N_24047,N_24880);
nand UO_1894 (O_1894,N_23865,N_24853);
or UO_1895 (O_1895,N_24768,N_24310);
xor UO_1896 (O_1896,N_24717,N_24727);
nand UO_1897 (O_1897,N_24332,N_24457);
nand UO_1898 (O_1898,N_24775,N_24482);
nand UO_1899 (O_1899,N_24949,N_24676);
xnor UO_1900 (O_1900,N_24920,N_24148);
and UO_1901 (O_1901,N_24378,N_24815);
or UO_1902 (O_1902,N_24791,N_24315);
nor UO_1903 (O_1903,N_24645,N_24824);
nand UO_1904 (O_1904,N_24050,N_23886);
and UO_1905 (O_1905,N_23824,N_24118);
and UO_1906 (O_1906,N_24786,N_24908);
and UO_1907 (O_1907,N_24937,N_24241);
and UO_1908 (O_1908,N_24672,N_24948);
nor UO_1909 (O_1909,N_24299,N_24702);
nor UO_1910 (O_1910,N_23827,N_24923);
and UO_1911 (O_1911,N_23903,N_24183);
nand UO_1912 (O_1912,N_24659,N_24171);
and UO_1913 (O_1913,N_24665,N_24982);
nor UO_1914 (O_1914,N_24719,N_24981);
and UO_1915 (O_1915,N_24611,N_24349);
or UO_1916 (O_1916,N_24269,N_23934);
xor UO_1917 (O_1917,N_24496,N_24696);
and UO_1918 (O_1918,N_24429,N_23919);
xor UO_1919 (O_1919,N_24308,N_24266);
or UO_1920 (O_1920,N_24241,N_23926);
xnor UO_1921 (O_1921,N_24859,N_24769);
nand UO_1922 (O_1922,N_24309,N_24289);
or UO_1923 (O_1923,N_24411,N_24742);
xnor UO_1924 (O_1924,N_24640,N_24803);
xor UO_1925 (O_1925,N_24179,N_23751);
nor UO_1926 (O_1926,N_24920,N_23863);
and UO_1927 (O_1927,N_23755,N_23787);
or UO_1928 (O_1928,N_23792,N_24503);
or UO_1929 (O_1929,N_24954,N_24904);
and UO_1930 (O_1930,N_23780,N_24579);
and UO_1931 (O_1931,N_24678,N_24265);
nand UO_1932 (O_1932,N_24147,N_24791);
xor UO_1933 (O_1933,N_24467,N_23893);
or UO_1934 (O_1934,N_24108,N_24952);
nand UO_1935 (O_1935,N_24724,N_23865);
and UO_1936 (O_1936,N_24541,N_24405);
xor UO_1937 (O_1937,N_23876,N_24310);
or UO_1938 (O_1938,N_23856,N_23756);
nor UO_1939 (O_1939,N_24597,N_24617);
or UO_1940 (O_1940,N_24447,N_24591);
or UO_1941 (O_1941,N_24933,N_24964);
xor UO_1942 (O_1942,N_23888,N_23791);
and UO_1943 (O_1943,N_24918,N_24876);
nand UO_1944 (O_1944,N_24135,N_24740);
or UO_1945 (O_1945,N_24541,N_24482);
nand UO_1946 (O_1946,N_24209,N_23963);
nor UO_1947 (O_1947,N_24188,N_24916);
nand UO_1948 (O_1948,N_24155,N_24811);
nand UO_1949 (O_1949,N_23979,N_23869);
nand UO_1950 (O_1950,N_24945,N_24869);
xor UO_1951 (O_1951,N_23864,N_24673);
and UO_1952 (O_1952,N_23778,N_24612);
nand UO_1953 (O_1953,N_24318,N_24101);
nor UO_1954 (O_1954,N_23960,N_24579);
and UO_1955 (O_1955,N_24649,N_24626);
nor UO_1956 (O_1956,N_24912,N_24354);
nand UO_1957 (O_1957,N_24008,N_24020);
nand UO_1958 (O_1958,N_24546,N_23862);
nand UO_1959 (O_1959,N_24809,N_24063);
or UO_1960 (O_1960,N_23960,N_24306);
and UO_1961 (O_1961,N_24095,N_24479);
and UO_1962 (O_1962,N_24339,N_24792);
nor UO_1963 (O_1963,N_24816,N_23795);
or UO_1964 (O_1964,N_24281,N_24305);
nor UO_1965 (O_1965,N_23892,N_23945);
nor UO_1966 (O_1966,N_24329,N_24912);
xnor UO_1967 (O_1967,N_24851,N_24794);
and UO_1968 (O_1968,N_23785,N_24267);
nor UO_1969 (O_1969,N_24155,N_24661);
nand UO_1970 (O_1970,N_24817,N_24810);
or UO_1971 (O_1971,N_24994,N_24432);
or UO_1972 (O_1972,N_24403,N_24730);
nor UO_1973 (O_1973,N_24359,N_23865);
or UO_1974 (O_1974,N_24127,N_23769);
and UO_1975 (O_1975,N_24146,N_23888);
nand UO_1976 (O_1976,N_24130,N_23978);
nand UO_1977 (O_1977,N_23936,N_24050);
xor UO_1978 (O_1978,N_24154,N_24936);
nor UO_1979 (O_1979,N_24747,N_24980);
nor UO_1980 (O_1980,N_23846,N_23841);
or UO_1981 (O_1981,N_24800,N_24975);
xnor UO_1982 (O_1982,N_24156,N_24269);
or UO_1983 (O_1983,N_24311,N_24754);
xor UO_1984 (O_1984,N_24413,N_23836);
xnor UO_1985 (O_1985,N_24399,N_24928);
nand UO_1986 (O_1986,N_24026,N_24288);
and UO_1987 (O_1987,N_24631,N_24419);
nor UO_1988 (O_1988,N_24893,N_24632);
or UO_1989 (O_1989,N_24120,N_24283);
or UO_1990 (O_1990,N_24565,N_24269);
xnor UO_1991 (O_1991,N_24029,N_24203);
or UO_1992 (O_1992,N_23751,N_24474);
or UO_1993 (O_1993,N_24256,N_24962);
nor UO_1994 (O_1994,N_24040,N_24631);
or UO_1995 (O_1995,N_23958,N_24283);
nor UO_1996 (O_1996,N_24400,N_24123);
or UO_1997 (O_1997,N_24861,N_24724);
and UO_1998 (O_1998,N_24709,N_24976);
and UO_1999 (O_1999,N_24726,N_24017);
or UO_2000 (O_2000,N_24561,N_23758);
or UO_2001 (O_2001,N_24549,N_24252);
or UO_2002 (O_2002,N_24403,N_23769);
nand UO_2003 (O_2003,N_23855,N_24546);
nor UO_2004 (O_2004,N_24294,N_23939);
and UO_2005 (O_2005,N_24034,N_24182);
nor UO_2006 (O_2006,N_23825,N_24014);
or UO_2007 (O_2007,N_24124,N_23987);
nand UO_2008 (O_2008,N_24918,N_24482);
nand UO_2009 (O_2009,N_24300,N_24680);
and UO_2010 (O_2010,N_24332,N_24941);
nand UO_2011 (O_2011,N_24681,N_24191);
or UO_2012 (O_2012,N_23973,N_23792);
or UO_2013 (O_2013,N_24211,N_24235);
nand UO_2014 (O_2014,N_24894,N_23950);
xor UO_2015 (O_2015,N_23867,N_24366);
xnor UO_2016 (O_2016,N_24775,N_24020);
nand UO_2017 (O_2017,N_23920,N_24260);
or UO_2018 (O_2018,N_24453,N_23942);
or UO_2019 (O_2019,N_24252,N_24337);
and UO_2020 (O_2020,N_23790,N_23855);
or UO_2021 (O_2021,N_24906,N_24478);
nand UO_2022 (O_2022,N_24085,N_24970);
nor UO_2023 (O_2023,N_24596,N_24166);
nand UO_2024 (O_2024,N_23766,N_24728);
xnor UO_2025 (O_2025,N_24273,N_23920);
and UO_2026 (O_2026,N_23890,N_24944);
xnor UO_2027 (O_2027,N_24992,N_24885);
xnor UO_2028 (O_2028,N_24566,N_23784);
and UO_2029 (O_2029,N_24334,N_24137);
nor UO_2030 (O_2030,N_24120,N_24598);
nand UO_2031 (O_2031,N_24660,N_24098);
nor UO_2032 (O_2032,N_24332,N_24898);
nand UO_2033 (O_2033,N_24273,N_24137);
nand UO_2034 (O_2034,N_23923,N_24378);
or UO_2035 (O_2035,N_24071,N_23850);
nand UO_2036 (O_2036,N_24248,N_24206);
and UO_2037 (O_2037,N_23953,N_24936);
and UO_2038 (O_2038,N_24933,N_24762);
nand UO_2039 (O_2039,N_24666,N_23808);
nor UO_2040 (O_2040,N_24750,N_24761);
and UO_2041 (O_2041,N_24202,N_24641);
xnor UO_2042 (O_2042,N_24819,N_24571);
and UO_2043 (O_2043,N_24627,N_24543);
nor UO_2044 (O_2044,N_24762,N_24496);
or UO_2045 (O_2045,N_24740,N_23942);
and UO_2046 (O_2046,N_24893,N_23875);
or UO_2047 (O_2047,N_24094,N_23840);
nor UO_2048 (O_2048,N_23860,N_23891);
and UO_2049 (O_2049,N_24410,N_24790);
xor UO_2050 (O_2050,N_24742,N_24904);
nand UO_2051 (O_2051,N_23852,N_23781);
and UO_2052 (O_2052,N_23971,N_24737);
nand UO_2053 (O_2053,N_24930,N_23925);
nand UO_2054 (O_2054,N_24410,N_24769);
and UO_2055 (O_2055,N_24844,N_24298);
nand UO_2056 (O_2056,N_24458,N_24674);
and UO_2057 (O_2057,N_24295,N_24458);
xor UO_2058 (O_2058,N_24409,N_24779);
or UO_2059 (O_2059,N_24305,N_24456);
or UO_2060 (O_2060,N_24182,N_24702);
nor UO_2061 (O_2061,N_24522,N_24620);
nand UO_2062 (O_2062,N_24058,N_24355);
nor UO_2063 (O_2063,N_24969,N_24693);
xnor UO_2064 (O_2064,N_24004,N_24556);
xnor UO_2065 (O_2065,N_24273,N_24423);
or UO_2066 (O_2066,N_24699,N_24828);
and UO_2067 (O_2067,N_24847,N_24365);
nand UO_2068 (O_2068,N_23992,N_24808);
xnor UO_2069 (O_2069,N_24449,N_24270);
xnor UO_2070 (O_2070,N_24746,N_23970);
nand UO_2071 (O_2071,N_23999,N_23762);
or UO_2072 (O_2072,N_24173,N_24769);
xnor UO_2073 (O_2073,N_24958,N_24325);
nand UO_2074 (O_2074,N_24817,N_23932);
nor UO_2075 (O_2075,N_24327,N_24752);
or UO_2076 (O_2076,N_24830,N_24657);
or UO_2077 (O_2077,N_24823,N_23939);
xnor UO_2078 (O_2078,N_23995,N_24241);
nor UO_2079 (O_2079,N_23820,N_24447);
nand UO_2080 (O_2080,N_24331,N_23994);
and UO_2081 (O_2081,N_24625,N_23938);
nor UO_2082 (O_2082,N_24833,N_24466);
or UO_2083 (O_2083,N_24522,N_23883);
xnor UO_2084 (O_2084,N_24578,N_23831);
nand UO_2085 (O_2085,N_24458,N_23925);
nand UO_2086 (O_2086,N_23873,N_24998);
or UO_2087 (O_2087,N_24940,N_23820);
and UO_2088 (O_2088,N_24564,N_24453);
or UO_2089 (O_2089,N_24822,N_24357);
or UO_2090 (O_2090,N_24847,N_24548);
xor UO_2091 (O_2091,N_24381,N_24471);
and UO_2092 (O_2092,N_23790,N_23879);
nor UO_2093 (O_2093,N_24373,N_23879);
or UO_2094 (O_2094,N_24210,N_24350);
or UO_2095 (O_2095,N_24892,N_24597);
nor UO_2096 (O_2096,N_24111,N_24047);
and UO_2097 (O_2097,N_24542,N_24429);
and UO_2098 (O_2098,N_24981,N_24437);
and UO_2099 (O_2099,N_24612,N_23799);
and UO_2100 (O_2100,N_23790,N_23994);
xor UO_2101 (O_2101,N_24989,N_24917);
or UO_2102 (O_2102,N_24862,N_24683);
nand UO_2103 (O_2103,N_24649,N_23890);
and UO_2104 (O_2104,N_24020,N_24012);
xor UO_2105 (O_2105,N_24500,N_23760);
xor UO_2106 (O_2106,N_24267,N_23964);
nand UO_2107 (O_2107,N_24631,N_23771);
nor UO_2108 (O_2108,N_24773,N_24752);
xor UO_2109 (O_2109,N_24003,N_24326);
and UO_2110 (O_2110,N_24416,N_24026);
and UO_2111 (O_2111,N_24612,N_23771);
nand UO_2112 (O_2112,N_24949,N_23930);
or UO_2113 (O_2113,N_24471,N_24507);
and UO_2114 (O_2114,N_24751,N_24307);
and UO_2115 (O_2115,N_24605,N_24961);
or UO_2116 (O_2116,N_24393,N_24569);
nor UO_2117 (O_2117,N_24442,N_24302);
nand UO_2118 (O_2118,N_24578,N_24027);
xnor UO_2119 (O_2119,N_24501,N_24322);
nand UO_2120 (O_2120,N_24631,N_24803);
or UO_2121 (O_2121,N_24755,N_24420);
nand UO_2122 (O_2122,N_23909,N_24291);
xor UO_2123 (O_2123,N_23759,N_24382);
or UO_2124 (O_2124,N_24349,N_24032);
nor UO_2125 (O_2125,N_23874,N_24574);
or UO_2126 (O_2126,N_23887,N_24816);
and UO_2127 (O_2127,N_24397,N_24863);
nor UO_2128 (O_2128,N_24459,N_24981);
nor UO_2129 (O_2129,N_23766,N_24982);
or UO_2130 (O_2130,N_24121,N_23871);
and UO_2131 (O_2131,N_24248,N_24865);
and UO_2132 (O_2132,N_24186,N_24891);
nand UO_2133 (O_2133,N_23825,N_23888);
and UO_2134 (O_2134,N_24199,N_24212);
nand UO_2135 (O_2135,N_24994,N_24311);
nor UO_2136 (O_2136,N_24810,N_24107);
and UO_2137 (O_2137,N_24909,N_24753);
and UO_2138 (O_2138,N_23834,N_24812);
nand UO_2139 (O_2139,N_24515,N_24725);
nor UO_2140 (O_2140,N_23988,N_24220);
xnor UO_2141 (O_2141,N_24406,N_23979);
nor UO_2142 (O_2142,N_24456,N_23788);
nand UO_2143 (O_2143,N_24886,N_24596);
xnor UO_2144 (O_2144,N_24668,N_23952);
or UO_2145 (O_2145,N_23896,N_24018);
and UO_2146 (O_2146,N_24190,N_24246);
nor UO_2147 (O_2147,N_24593,N_24084);
and UO_2148 (O_2148,N_24334,N_23894);
xor UO_2149 (O_2149,N_24874,N_24649);
xnor UO_2150 (O_2150,N_24644,N_24792);
nand UO_2151 (O_2151,N_24874,N_23992);
nor UO_2152 (O_2152,N_23853,N_23943);
xnor UO_2153 (O_2153,N_24655,N_24048);
or UO_2154 (O_2154,N_24161,N_24895);
or UO_2155 (O_2155,N_24223,N_24284);
nand UO_2156 (O_2156,N_24603,N_24830);
or UO_2157 (O_2157,N_24608,N_24497);
xor UO_2158 (O_2158,N_23844,N_23823);
xnor UO_2159 (O_2159,N_24996,N_24314);
xor UO_2160 (O_2160,N_24016,N_24663);
or UO_2161 (O_2161,N_23801,N_23853);
xor UO_2162 (O_2162,N_24984,N_24311);
or UO_2163 (O_2163,N_24652,N_24129);
xor UO_2164 (O_2164,N_23832,N_24905);
nor UO_2165 (O_2165,N_24646,N_24114);
nor UO_2166 (O_2166,N_24346,N_24402);
nor UO_2167 (O_2167,N_24715,N_24218);
or UO_2168 (O_2168,N_24999,N_23765);
nand UO_2169 (O_2169,N_24036,N_23903);
and UO_2170 (O_2170,N_23957,N_24466);
or UO_2171 (O_2171,N_24336,N_24397);
nor UO_2172 (O_2172,N_24322,N_24166);
nor UO_2173 (O_2173,N_24248,N_24422);
and UO_2174 (O_2174,N_24675,N_24702);
or UO_2175 (O_2175,N_24294,N_24260);
or UO_2176 (O_2176,N_24533,N_24671);
xnor UO_2177 (O_2177,N_24598,N_24720);
nor UO_2178 (O_2178,N_24184,N_24545);
nor UO_2179 (O_2179,N_24662,N_23898);
xor UO_2180 (O_2180,N_24693,N_24680);
xnor UO_2181 (O_2181,N_23865,N_23864);
and UO_2182 (O_2182,N_24580,N_24290);
xnor UO_2183 (O_2183,N_23993,N_24500);
and UO_2184 (O_2184,N_23822,N_24779);
nand UO_2185 (O_2185,N_24273,N_24305);
nor UO_2186 (O_2186,N_24220,N_24629);
nand UO_2187 (O_2187,N_23912,N_23858);
xnor UO_2188 (O_2188,N_24081,N_24769);
xnor UO_2189 (O_2189,N_23753,N_24836);
nor UO_2190 (O_2190,N_23754,N_24720);
nor UO_2191 (O_2191,N_24134,N_24564);
nor UO_2192 (O_2192,N_24966,N_24406);
nor UO_2193 (O_2193,N_24691,N_24223);
and UO_2194 (O_2194,N_24201,N_23978);
and UO_2195 (O_2195,N_24620,N_24312);
nand UO_2196 (O_2196,N_23809,N_24145);
nor UO_2197 (O_2197,N_24039,N_24154);
nand UO_2198 (O_2198,N_24443,N_23885);
nor UO_2199 (O_2199,N_24058,N_24574);
nor UO_2200 (O_2200,N_23910,N_24017);
and UO_2201 (O_2201,N_24263,N_24359);
nor UO_2202 (O_2202,N_24585,N_23889);
nand UO_2203 (O_2203,N_24116,N_24161);
or UO_2204 (O_2204,N_23962,N_23949);
nor UO_2205 (O_2205,N_23857,N_24781);
nor UO_2206 (O_2206,N_24276,N_24487);
xnor UO_2207 (O_2207,N_24254,N_24024);
xnor UO_2208 (O_2208,N_24483,N_23937);
nand UO_2209 (O_2209,N_24839,N_23849);
nand UO_2210 (O_2210,N_24541,N_24942);
nor UO_2211 (O_2211,N_24082,N_23925);
and UO_2212 (O_2212,N_24917,N_24405);
or UO_2213 (O_2213,N_24650,N_24952);
nand UO_2214 (O_2214,N_23880,N_24745);
xor UO_2215 (O_2215,N_24404,N_24877);
and UO_2216 (O_2216,N_24041,N_24457);
or UO_2217 (O_2217,N_24101,N_24420);
xor UO_2218 (O_2218,N_23816,N_23792);
xnor UO_2219 (O_2219,N_24852,N_24670);
xor UO_2220 (O_2220,N_24906,N_24706);
xnor UO_2221 (O_2221,N_24645,N_24563);
xor UO_2222 (O_2222,N_23902,N_23830);
or UO_2223 (O_2223,N_24929,N_24637);
and UO_2224 (O_2224,N_24238,N_24232);
and UO_2225 (O_2225,N_24951,N_24694);
nand UO_2226 (O_2226,N_24280,N_24339);
xnor UO_2227 (O_2227,N_24105,N_24316);
xor UO_2228 (O_2228,N_23849,N_24549);
or UO_2229 (O_2229,N_24409,N_23765);
or UO_2230 (O_2230,N_24266,N_23925);
nand UO_2231 (O_2231,N_23945,N_23754);
and UO_2232 (O_2232,N_24988,N_24405);
and UO_2233 (O_2233,N_23932,N_23798);
xnor UO_2234 (O_2234,N_23779,N_24649);
and UO_2235 (O_2235,N_24131,N_24867);
xor UO_2236 (O_2236,N_23877,N_23853);
and UO_2237 (O_2237,N_24317,N_24979);
or UO_2238 (O_2238,N_24205,N_24809);
nor UO_2239 (O_2239,N_24365,N_24084);
and UO_2240 (O_2240,N_23901,N_24705);
or UO_2241 (O_2241,N_24743,N_24034);
nor UO_2242 (O_2242,N_24749,N_24269);
or UO_2243 (O_2243,N_24494,N_24295);
nor UO_2244 (O_2244,N_24181,N_23781);
nand UO_2245 (O_2245,N_24987,N_24313);
xnor UO_2246 (O_2246,N_24293,N_23993);
nand UO_2247 (O_2247,N_23755,N_24197);
and UO_2248 (O_2248,N_24042,N_23953);
xor UO_2249 (O_2249,N_24937,N_24459);
or UO_2250 (O_2250,N_24725,N_24973);
nor UO_2251 (O_2251,N_24352,N_24913);
nand UO_2252 (O_2252,N_24370,N_24512);
nor UO_2253 (O_2253,N_23849,N_24811);
or UO_2254 (O_2254,N_24496,N_24362);
and UO_2255 (O_2255,N_24671,N_24518);
nand UO_2256 (O_2256,N_24887,N_24307);
nand UO_2257 (O_2257,N_24684,N_24966);
or UO_2258 (O_2258,N_23765,N_24192);
or UO_2259 (O_2259,N_23941,N_24578);
or UO_2260 (O_2260,N_23756,N_24886);
or UO_2261 (O_2261,N_24746,N_23787);
nand UO_2262 (O_2262,N_24260,N_24376);
or UO_2263 (O_2263,N_24999,N_23822);
and UO_2264 (O_2264,N_24707,N_24019);
or UO_2265 (O_2265,N_24826,N_24768);
xor UO_2266 (O_2266,N_24921,N_24062);
or UO_2267 (O_2267,N_24229,N_24256);
xor UO_2268 (O_2268,N_23845,N_23947);
or UO_2269 (O_2269,N_24269,N_24105);
nand UO_2270 (O_2270,N_24321,N_23996);
and UO_2271 (O_2271,N_24909,N_23807);
nor UO_2272 (O_2272,N_24610,N_24540);
xor UO_2273 (O_2273,N_24444,N_24889);
xor UO_2274 (O_2274,N_24989,N_24650);
nand UO_2275 (O_2275,N_23851,N_24082);
xor UO_2276 (O_2276,N_24210,N_23961);
nor UO_2277 (O_2277,N_24920,N_24311);
or UO_2278 (O_2278,N_24256,N_24899);
and UO_2279 (O_2279,N_24169,N_24392);
and UO_2280 (O_2280,N_24264,N_24524);
or UO_2281 (O_2281,N_24002,N_24161);
nor UO_2282 (O_2282,N_23921,N_23863);
nor UO_2283 (O_2283,N_23832,N_24993);
and UO_2284 (O_2284,N_24766,N_24842);
and UO_2285 (O_2285,N_24418,N_24032);
xor UO_2286 (O_2286,N_24122,N_24439);
nor UO_2287 (O_2287,N_24210,N_24689);
nor UO_2288 (O_2288,N_24094,N_23782);
xnor UO_2289 (O_2289,N_24124,N_23842);
nor UO_2290 (O_2290,N_24289,N_24285);
and UO_2291 (O_2291,N_24410,N_24696);
xnor UO_2292 (O_2292,N_24900,N_24666);
nand UO_2293 (O_2293,N_23836,N_24813);
and UO_2294 (O_2294,N_24030,N_24892);
xor UO_2295 (O_2295,N_23927,N_23762);
nor UO_2296 (O_2296,N_24750,N_24797);
or UO_2297 (O_2297,N_24538,N_24843);
or UO_2298 (O_2298,N_24227,N_24497);
or UO_2299 (O_2299,N_24077,N_24712);
nor UO_2300 (O_2300,N_24367,N_24529);
or UO_2301 (O_2301,N_24617,N_23755);
nor UO_2302 (O_2302,N_24289,N_23928);
or UO_2303 (O_2303,N_23827,N_24635);
and UO_2304 (O_2304,N_24165,N_23941);
nand UO_2305 (O_2305,N_24153,N_24782);
and UO_2306 (O_2306,N_23843,N_24496);
nor UO_2307 (O_2307,N_24221,N_24666);
xor UO_2308 (O_2308,N_24892,N_23928);
nand UO_2309 (O_2309,N_24658,N_24469);
nor UO_2310 (O_2310,N_24408,N_24492);
xor UO_2311 (O_2311,N_24724,N_23904);
xnor UO_2312 (O_2312,N_23827,N_23918);
nor UO_2313 (O_2313,N_23881,N_24952);
nand UO_2314 (O_2314,N_24143,N_24790);
or UO_2315 (O_2315,N_24298,N_24119);
nand UO_2316 (O_2316,N_24494,N_24355);
nor UO_2317 (O_2317,N_24981,N_23782);
nand UO_2318 (O_2318,N_23957,N_23984);
nand UO_2319 (O_2319,N_24650,N_24136);
and UO_2320 (O_2320,N_24648,N_24007);
nor UO_2321 (O_2321,N_24924,N_24195);
or UO_2322 (O_2322,N_24186,N_24308);
nor UO_2323 (O_2323,N_23751,N_24814);
nand UO_2324 (O_2324,N_23957,N_24734);
nand UO_2325 (O_2325,N_24588,N_24243);
nand UO_2326 (O_2326,N_24704,N_23975);
xnor UO_2327 (O_2327,N_23815,N_24971);
xor UO_2328 (O_2328,N_23883,N_24888);
nand UO_2329 (O_2329,N_24214,N_24684);
xnor UO_2330 (O_2330,N_24365,N_24364);
and UO_2331 (O_2331,N_24531,N_23951);
or UO_2332 (O_2332,N_24952,N_24906);
xor UO_2333 (O_2333,N_24022,N_23764);
nand UO_2334 (O_2334,N_24382,N_23809);
nor UO_2335 (O_2335,N_23954,N_24563);
nor UO_2336 (O_2336,N_24519,N_24762);
or UO_2337 (O_2337,N_24964,N_24458);
and UO_2338 (O_2338,N_24403,N_24129);
and UO_2339 (O_2339,N_24500,N_24812);
nand UO_2340 (O_2340,N_23984,N_24678);
or UO_2341 (O_2341,N_24154,N_24544);
nand UO_2342 (O_2342,N_24830,N_23870);
nand UO_2343 (O_2343,N_24364,N_23808);
or UO_2344 (O_2344,N_24246,N_23969);
nor UO_2345 (O_2345,N_23841,N_23873);
nor UO_2346 (O_2346,N_24963,N_23811);
xor UO_2347 (O_2347,N_24897,N_24893);
nand UO_2348 (O_2348,N_23913,N_24364);
or UO_2349 (O_2349,N_24905,N_24427);
or UO_2350 (O_2350,N_23974,N_24116);
and UO_2351 (O_2351,N_24459,N_24326);
nand UO_2352 (O_2352,N_24386,N_24420);
xnor UO_2353 (O_2353,N_23842,N_24616);
nor UO_2354 (O_2354,N_23898,N_23939);
nor UO_2355 (O_2355,N_24998,N_24724);
or UO_2356 (O_2356,N_24089,N_23754);
xor UO_2357 (O_2357,N_24738,N_24970);
nand UO_2358 (O_2358,N_24206,N_24453);
or UO_2359 (O_2359,N_24162,N_23787);
nor UO_2360 (O_2360,N_23753,N_23936);
nor UO_2361 (O_2361,N_24711,N_24203);
xnor UO_2362 (O_2362,N_24398,N_24176);
and UO_2363 (O_2363,N_24519,N_24027);
xnor UO_2364 (O_2364,N_24385,N_24368);
xor UO_2365 (O_2365,N_24235,N_24675);
nand UO_2366 (O_2366,N_24656,N_24738);
and UO_2367 (O_2367,N_24755,N_24357);
xnor UO_2368 (O_2368,N_24196,N_23836);
xor UO_2369 (O_2369,N_24952,N_24587);
and UO_2370 (O_2370,N_23859,N_24813);
nand UO_2371 (O_2371,N_24695,N_24405);
xnor UO_2372 (O_2372,N_23804,N_24748);
xnor UO_2373 (O_2373,N_24400,N_24723);
or UO_2374 (O_2374,N_24186,N_24531);
xnor UO_2375 (O_2375,N_24264,N_24573);
nand UO_2376 (O_2376,N_24793,N_24081);
and UO_2377 (O_2377,N_23858,N_23822);
or UO_2378 (O_2378,N_24917,N_24440);
nor UO_2379 (O_2379,N_23893,N_23979);
xor UO_2380 (O_2380,N_24438,N_24050);
nor UO_2381 (O_2381,N_24404,N_24801);
nand UO_2382 (O_2382,N_24696,N_24161);
or UO_2383 (O_2383,N_24306,N_24598);
and UO_2384 (O_2384,N_24200,N_23782);
nand UO_2385 (O_2385,N_23938,N_24877);
nand UO_2386 (O_2386,N_23842,N_24504);
nor UO_2387 (O_2387,N_24763,N_24466);
nor UO_2388 (O_2388,N_23937,N_24846);
or UO_2389 (O_2389,N_24878,N_24477);
and UO_2390 (O_2390,N_24661,N_24353);
nor UO_2391 (O_2391,N_24717,N_23939);
nand UO_2392 (O_2392,N_23771,N_23772);
and UO_2393 (O_2393,N_24573,N_24931);
nand UO_2394 (O_2394,N_24769,N_24375);
nor UO_2395 (O_2395,N_24039,N_24077);
xor UO_2396 (O_2396,N_24997,N_24939);
or UO_2397 (O_2397,N_24959,N_23763);
nor UO_2398 (O_2398,N_23947,N_24140);
or UO_2399 (O_2399,N_24325,N_24419);
or UO_2400 (O_2400,N_23841,N_24948);
nor UO_2401 (O_2401,N_23981,N_24394);
xnor UO_2402 (O_2402,N_24228,N_23999);
and UO_2403 (O_2403,N_24697,N_24064);
nor UO_2404 (O_2404,N_23781,N_24855);
xor UO_2405 (O_2405,N_24220,N_23842);
and UO_2406 (O_2406,N_24287,N_23853);
and UO_2407 (O_2407,N_23777,N_24874);
nor UO_2408 (O_2408,N_24802,N_24305);
nor UO_2409 (O_2409,N_24905,N_24067);
or UO_2410 (O_2410,N_23882,N_24001);
xnor UO_2411 (O_2411,N_24689,N_24225);
or UO_2412 (O_2412,N_24247,N_23891);
nor UO_2413 (O_2413,N_24732,N_24209);
nor UO_2414 (O_2414,N_24035,N_24249);
nor UO_2415 (O_2415,N_23929,N_24742);
xor UO_2416 (O_2416,N_23912,N_23881);
or UO_2417 (O_2417,N_24420,N_24611);
or UO_2418 (O_2418,N_24510,N_24311);
xnor UO_2419 (O_2419,N_24555,N_24208);
xnor UO_2420 (O_2420,N_24013,N_24572);
nand UO_2421 (O_2421,N_24813,N_23955);
xor UO_2422 (O_2422,N_24244,N_23781);
and UO_2423 (O_2423,N_23891,N_23820);
or UO_2424 (O_2424,N_24366,N_24662);
nand UO_2425 (O_2425,N_24955,N_24392);
and UO_2426 (O_2426,N_24664,N_23978);
or UO_2427 (O_2427,N_24628,N_24506);
nor UO_2428 (O_2428,N_24397,N_24637);
and UO_2429 (O_2429,N_24777,N_24355);
and UO_2430 (O_2430,N_23845,N_24316);
or UO_2431 (O_2431,N_24592,N_24498);
xnor UO_2432 (O_2432,N_24559,N_24226);
or UO_2433 (O_2433,N_24859,N_24699);
or UO_2434 (O_2434,N_24234,N_23750);
or UO_2435 (O_2435,N_24290,N_24920);
xor UO_2436 (O_2436,N_24351,N_23928);
or UO_2437 (O_2437,N_24144,N_24925);
xnor UO_2438 (O_2438,N_24359,N_24883);
and UO_2439 (O_2439,N_24183,N_24980);
nand UO_2440 (O_2440,N_24197,N_24776);
nor UO_2441 (O_2441,N_24199,N_24869);
and UO_2442 (O_2442,N_24119,N_24281);
and UO_2443 (O_2443,N_24479,N_23787);
or UO_2444 (O_2444,N_24326,N_24219);
xor UO_2445 (O_2445,N_24076,N_24470);
or UO_2446 (O_2446,N_24322,N_24095);
and UO_2447 (O_2447,N_23780,N_24066);
nand UO_2448 (O_2448,N_24624,N_23897);
nand UO_2449 (O_2449,N_24977,N_23850);
nand UO_2450 (O_2450,N_24641,N_24937);
and UO_2451 (O_2451,N_24404,N_24019);
or UO_2452 (O_2452,N_24133,N_24716);
or UO_2453 (O_2453,N_24386,N_24541);
nand UO_2454 (O_2454,N_24527,N_24691);
and UO_2455 (O_2455,N_24445,N_24321);
nor UO_2456 (O_2456,N_24143,N_24268);
xnor UO_2457 (O_2457,N_24544,N_23783);
or UO_2458 (O_2458,N_24001,N_24827);
nand UO_2459 (O_2459,N_23877,N_24062);
xnor UO_2460 (O_2460,N_24132,N_23779);
and UO_2461 (O_2461,N_24676,N_24066);
nand UO_2462 (O_2462,N_24272,N_23892);
and UO_2463 (O_2463,N_24879,N_24953);
nand UO_2464 (O_2464,N_23786,N_24832);
and UO_2465 (O_2465,N_24090,N_23934);
nand UO_2466 (O_2466,N_23958,N_24369);
xnor UO_2467 (O_2467,N_24288,N_24565);
and UO_2468 (O_2468,N_24087,N_23967);
xnor UO_2469 (O_2469,N_24831,N_24576);
xor UO_2470 (O_2470,N_24845,N_23913);
xnor UO_2471 (O_2471,N_24995,N_24286);
or UO_2472 (O_2472,N_23773,N_23760);
nor UO_2473 (O_2473,N_24910,N_23999);
or UO_2474 (O_2474,N_24257,N_24545);
nand UO_2475 (O_2475,N_24359,N_23790);
or UO_2476 (O_2476,N_23842,N_24310);
nor UO_2477 (O_2477,N_24871,N_24327);
nor UO_2478 (O_2478,N_24889,N_23817);
nor UO_2479 (O_2479,N_24207,N_24595);
xor UO_2480 (O_2480,N_24289,N_23778);
nand UO_2481 (O_2481,N_24000,N_24580);
nor UO_2482 (O_2482,N_23812,N_24181);
nand UO_2483 (O_2483,N_24819,N_24509);
nor UO_2484 (O_2484,N_24031,N_23789);
nor UO_2485 (O_2485,N_24131,N_24778);
or UO_2486 (O_2486,N_24918,N_24513);
and UO_2487 (O_2487,N_24398,N_24912);
nor UO_2488 (O_2488,N_24553,N_24168);
nor UO_2489 (O_2489,N_24215,N_23971);
nor UO_2490 (O_2490,N_24558,N_24970);
nor UO_2491 (O_2491,N_24351,N_24134);
and UO_2492 (O_2492,N_24929,N_24922);
nor UO_2493 (O_2493,N_24617,N_24987);
nor UO_2494 (O_2494,N_24105,N_24552);
or UO_2495 (O_2495,N_24769,N_24266);
nand UO_2496 (O_2496,N_24860,N_24254);
or UO_2497 (O_2497,N_24461,N_24646);
nor UO_2498 (O_2498,N_24579,N_24858);
and UO_2499 (O_2499,N_23927,N_24576);
nor UO_2500 (O_2500,N_24708,N_24912);
xnor UO_2501 (O_2501,N_24305,N_24669);
xnor UO_2502 (O_2502,N_24061,N_24006);
and UO_2503 (O_2503,N_23783,N_23950);
xnor UO_2504 (O_2504,N_24881,N_24609);
or UO_2505 (O_2505,N_24518,N_23903);
or UO_2506 (O_2506,N_24543,N_23942);
nor UO_2507 (O_2507,N_24557,N_24477);
and UO_2508 (O_2508,N_24344,N_24413);
or UO_2509 (O_2509,N_24485,N_24634);
and UO_2510 (O_2510,N_24523,N_24489);
and UO_2511 (O_2511,N_24057,N_24898);
and UO_2512 (O_2512,N_24730,N_24534);
and UO_2513 (O_2513,N_23821,N_24038);
and UO_2514 (O_2514,N_23886,N_24313);
nor UO_2515 (O_2515,N_24913,N_24382);
and UO_2516 (O_2516,N_24088,N_24319);
nand UO_2517 (O_2517,N_24892,N_24363);
or UO_2518 (O_2518,N_24753,N_24728);
and UO_2519 (O_2519,N_24879,N_24323);
xor UO_2520 (O_2520,N_23756,N_23983);
nand UO_2521 (O_2521,N_23991,N_24115);
nand UO_2522 (O_2522,N_24916,N_24733);
xor UO_2523 (O_2523,N_24166,N_24396);
nand UO_2524 (O_2524,N_23829,N_24116);
and UO_2525 (O_2525,N_24206,N_23992);
or UO_2526 (O_2526,N_23755,N_24423);
nand UO_2527 (O_2527,N_24935,N_23773);
nor UO_2528 (O_2528,N_24192,N_24959);
nand UO_2529 (O_2529,N_24252,N_23959);
nor UO_2530 (O_2530,N_24101,N_24286);
or UO_2531 (O_2531,N_24057,N_23967);
or UO_2532 (O_2532,N_24219,N_24315);
xnor UO_2533 (O_2533,N_24930,N_24013);
xnor UO_2534 (O_2534,N_24735,N_24543);
and UO_2535 (O_2535,N_24517,N_24918);
nor UO_2536 (O_2536,N_24215,N_23896);
nand UO_2537 (O_2537,N_23801,N_24723);
nor UO_2538 (O_2538,N_24089,N_24284);
xor UO_2539 (O_2539,N_24976,N_24869);
and UO_2540 (O_2540,N_23978,N_24290);
and UO_2541 (O_2541,N_24436,N_24408);
nand UO_2542 (O_2542,N_24496,N_24013);
or UO_2543 (O_2543,N_24545,N_24941);
nand UO_2544 (O_2544,N_24100,N_24138);
or UO_2545 (O_2545,N_24942,N_24505);
nor UO_2546 (O_2546,N_23961,N_24388);
or UO_2547 (O_2547,N_24301,N_24023);
nand UO_2548 (O_2548,N_24574,N_24219);
nor UO_2549 (O_2549,N_24528,N_24481);
nand UO_2550 (O_2550,N_24928,N_24725);
or UO_2551 (O_2551,N_24234,N_24121);
and UO_2552 (O_2552,N_23956,N_24976);
nand UO_2553 (O_2553,N_24622,N_24734);
or UO_2554 (O_2554,N_24983,N_24389);
or UO_2555 (O_2555,N_24799,N_24788);
or UO_2556 (O_2556,N_23784,N_24980);
or UO_2557 (O_2557,N_24281,N_24763);
nor UO_2558 (O_2558,N_24604,N_24039);
and UO_2559 (O_2559,N_24726,N_24300);
xor UO_2560 (O_2560,N_24575,N_24582);
nor UO_2561 (O_2561,N_24444,N_24969);
and UO_2562 (O_2562,N_24101,N_24251);
and UO_2563 (O_2563,N_24082,N_23856);
or UO_2564 (O_2564,N_24768,N_24773);
nand UO_2565 (O_2565,N_23884,N_23953);
nor UO_2566 (O_2566,N_24441,N_23957);
or UO_2567 (O_2567,N_23962,N_24575);
and UO_2568 (O_2568,N_24063,N_24988);
nand UO_2569 (O_2569,N_24015,N_24296);
xnor UO_2570 (O_2570,N_24698,N_23880);
nand UO_2571 (O_2571,N_24549,N_23966);
xor UO_2572 (O_2572,N_23810,N_24461);
xnor UO_2573 (O_2573,N_24936,N_23845);
nor UO_2574 (O_2574,N_24823,N_24530);
and UO_2575 (O_2575,N_23982,N_24202);
nand UO_2576 (O_2576,N_23869,N_24852);
nor UO_2577 (O_2577,N_24711,N_24451);
nor UO_2578 (O_2578,N_24982,N_24762);
nor UO_2579 (O_2579,N_24620,N_24724);
nor UO_2580 (O_2580,N_23991,N_24660);
nor UO_2581 (O_2581,N_24827,N_24142);
nor UO_2582 (O_2582,N_24973,N_23992);
or UO_2583 (O_2583,N_24652,N_23924);
nor UO_2584 (O_2584,N_24316,N_24547);
nor UO_2585 (O_2585,N_24282,N_24675);
nor UO_2586 (O_2586,N_24440,N_24367);
xnor UO_2587 (O_2587,N_24021,N_24869);
and UO_2588 (O_2588,N_24648,N_24982);
or UO_2589 (O_2589,N_24554,N_24960);
or UO_2590 (O_2590,N_24319,N_24120);
and UO_2591 (O_2591,N_23780,N_24496);
nand UO_2592 (O_2592,N_24176,N_23752);
and UO_2593 (O_2593,N_24469,N_24793);
nor UO_2594 (O_2594,N_24412,N_24728);
nand UO_2595 (O_2595,N_24277,N_24168);
nor UO_2596 (O_2596,N_24818,N_24133);
and UO_2597 (O_2597,N_24748,N_24195);
and UO_2598 (O_2598,N_23915,N_24471);
xnor UO_2599 (O_2599,N_24138,N_24899);
nor UO_2600 (O_2600,N_24987,N_24183);
and UO_2601 (O_2601,N_24423,N_23892);
nand UO_2602 (O_2602,N_24527,N_23781);
and UO_2603 (O_2603,N_24923,N_24912);
or UO_2604 (O_2604,N_24821,N_23958);
and UO_2605 (O_2605,N_24578,N_23755);
xor UO_2606 (O_2606,N_24073,N_23943);
nor UO_2607 (O_2607,N_23913,N_24254);
nor UO_2608 (O_2608,N_24229,N_23793);
or UO_2609 (O_2609,N_23926,N_24974);
nor UO_2610 (O_2610,N_24884,N_23752);
and UO_2611 (O_2611,N_24126,N_24501);
xnor UO_2612 (O_2612,N_23887,N_24142);
and UO_2613 (O_2613,N_23841,N_24939);
or UO_2614 (O_2614,N_24837,N_24876);
nor UO_2615 (O_2615,N_24901,N_24828);
nand UO_2616 (O_2616,N_24649,N_23912);
or UO_2617 (O_2617,N_24017,N_24965);
or UO_2618 (O_2618,N_24910,N_24256);
nor UO_2619 (O_2619,N_23855,N_24735);
nor UO_2620 (O_2620,N_23896,N_24715);
or UO_2621 (O_2621,N_24651,N_24959);
nor UO_2622 (O_2622,N_24395,N_24890);
nand UO_2623 (O_2623,N_24809,N_23895);
nand UO_2624 (O_2624,N_24514,N_24081);
or UO_2625 (O_2625,N_24360,N_24629);
and UO_2626 (O_2626,N_24946,N_24571);
or UO_2627 (O_2627,N_24984,N_24466);
nand UO_2628 (O_2628,N_24921,N_24056);
and UO_2629 (O_2629,N_24463,N_24842);
xnor UO_2630 (O_2630,N_24179,N_24947);
or UO_2631 (O_2631,N_24482,N_24899);
nand UO_2632 (O_2632,N_24981,N_24503);
nor UO_2633 (O_2633,N_23781,N_24820);
xor UO_2634 (O_2634,N_24289,N_24626);
or UO_2635 (O_2635,N_23933,N_24603);
or UO_2636 (O_2636,N_24184,N_23966);
nor UO_2637 (O_2637,N_24569,N_24741);
or UO_2638 (O_2638,N_23767,N_24913);
xnor UO_2639 (O_2639,N_23978,N_24327);
xor UO_2640 (O_2640,N_24783,N_24619);
nor UO_2641 (O_2641,N_24373,N_24686);
or UO_2642 (O_2642,N_24752,N_24155);
and UO_2643 (O_2643,N_24207,N_24497);
and UO_2644 (O_2644,N_23972,N_24588);
or UO_2645 (O_2645,N_23929,N_24651);
and UO_2646 (O_2646,N_24644,N_24879);
nor UO_2647 (O_2647,N_24367,N_24013);
nand UO_2648 (O_2648,N_24084,N_24351);
nor UO_2649 (O_2649,N_24490,N_24874);
or UO_2650 (O_2650,N_24952,N_24148);
or UO_2651 (O_2651,N_23966,N_23940);
nand UO_2652 (O_2652,N_24319,N_24738);
nand UO_2653 (O_2653,N_23975,N_24181);
and UO_2654 (O_2654,N_24233,N_23897);
or UO_2655 (O_2655,N_24882,N_23967);
nand UO_2656 (O_2656,N_23832,N_24819);
or UO_2657 (O_2657,N_24011,N_24710);
xor UO_2658 (O_2658,N_23942,N_24085);
nand UO_2659 (O_2659,N_23872,N_24922);
xor UO_2660 (O_2660,N_24782,N_24276);
nand UO_2661 (O_2661,N_23887,N_24348);
xor UO_2662 (O_2662,N_24092,N_24424);
and UO_2663 (O_2663,N_24215,N_24594);
nand UO_2664 (O_2664,N_24256,N_24374);
nand UO_2665 (O_2665,N_24604,N_23897);
nor UO_2666 (O_2666,N_23779,N_24514);
xor UO_2667 (O_2667,N_24476,N_24571);
xor UO_2668 (O_2668,N_23873,N_24508);
xnor UO_2669 (O_2669,N_23875,N_24970);
and UO_2670 (O_2670,N_23875,N_24419);
nor UO_2671 (O_2671,N_24539,N_23882);
nor UO_2672 (O_2672,N_24385,N_24213);
and UO_2673 (O_2673,N_24161,N_24775);
nor UO_2674 (O_2674,N_24881,N_24540);
or UO_2675 (O_2675,N_24162,N_24837);
and UO_2676 (O_2676,N_24925,N_24947);
nand UO_2677 (O_2677,N_24734,N_24337);
or UO_2678 (O_2678,N_24273,N_24520);
xnor UO_2679 (O_2679,N_24385,N_24654);
or UO_2680 (O_2680,N_24979,N_24076);
nor UO_2681 (O_2681,N_24140,N_24088);
xor UO_2682 (O_2682,N_24349,N_24284);
and UO_2683 (O_2683,N_24090,N_24326);
or UO_2684 (O_2684,N_23836,N_23811);
xnor UO_2685 (O_2685,N_23822,N_24669);
or UO_2686 (O_2686,N_24948,N_24915);
nor UO_2687 (O_2687,N_24826,N_24948);
nand UO_2688 (O_2688,N_24133,N_24316);
and UO_2689 (O_2689,N_24604,N_24721);
nand UO_2690 (O_2690,N_24596,N_24309);
nor UO_2691 (O_2691,N_24048,N_24435);
or UO_2692 (O_2692,N_24971,N_24177);
and UO_2693 (O_2693,N_24797,N_24091);
or UO_2694 (O_2694,N_24915,N_24505);
or UO_2695 (O_2695,N_24409,N_24271);
nor UO_2696 (O_2696,N_24103,N_24754);
xnor UO_2697 (O_2697,N_23821,N_23973);
and UO_2698 (O_2698,N_24086,N_24036);
nand UO_2699 (O_2699,N_23987,N_24309);
nand UO_2700 (O_2700,N_24762,N_24505);
xnor UO_2701 (O_2701,N_24593,N_24262);
or UO_2702 (O_2702,N_24628,N_23862);
or UO_2703 (O_2703,N_24824,N_24001);
nor UO_2704 (O_2704,N_24817,N_24639);
or UO_2705 (O_2705,N_24726,N_24194);
nand UO_2706 (O_2706,N_24076,N_24779);
or UO_2707 (O_2707,N_24260,N_24062);
and UO_2708 (O_2708,N_24356,N_24282);
nor UO_2709 (O_2709,N_24342,N_24581);
and UO_2710 (O_2710,N_24994,N_24967);
and UO_2711 (O_2711,N_24872,N_24668);
xnor UO_2712 (O_2712,N_24767,N_24527);
or UO_2713 (O_2713,N_24686,N_24174);
nor UO_2714 (O_2714,N_24038,N_24502);
nand UO_2715 (O_2715,N_24790,N_24741);
nor UO_2716 (O_2716,N_24787,N_24550);
xor UO_2717 (O_2717,N_24043,N_24469);
and UO_2718 (O_2718,N_24548,N_24891);
nor UO_2719 (O_2719,N_24488,N_24472);
nor UO_2720 (O_2720,N_24438,N_24603);
and UO_2721 (O_2721,N_23981,N_24120);
nand UO_2722 (O_2722,N_24283,N_24046);
or UO_2723 (O_2723,N_23887,N_24082);
xnor UO_2724 (O_2724,N_24944,N_24778);
xor UO_2725 (O_2725,N_23924,N_23800);
xnor UO_2726 (O_2726,N_24036,N_24963);
nand UO_2727 (O_2727,N_24105,N_24580);
nor UO_2728 (O_2728,N_24952,N_24976);
or UO_2729 (O_2729,N_24970,N_24500);
nand UO_2730 (O_2730,N_24236,N_23807);
and UO_2731 (O_2731,N_23763,N_23910);
nor UO_2732 (O_2732,N_24052,N_24653);
and UO_2733 (O_2733,N_23781,N_24727);
and UO_2734 (O_2734,N_24041,N_23902);
and UO_2735 (O_2735,N_24273,N_24060);
or UO_2736 (O_2736,N_23848,N_23752);
or UO_2737 (O_2737,N_24108,N_24033);
nor UO_2738 (O_2738,N_23898,N_23913);
nand UO_2739 (O_2739,N_23758,N_24962);
nand UO_2740 (O_2740,N_23915,N_24614);
and UO_2741 (O_2741,N_23753,N_24623);
or UO_2742 (O_2742,N_23841,N_23877);
nor UO_2743 (O_2743,N_24076,N_24609);
nor UO_2744 (O_2744,N_23959,N_24814);
and UO_2745 (O_2745,N_23829,N_24618);
or UO_2746 (O_2746,N_24577,N_24801);
xnor UO_2747 (O_2747,N_24345,N_23904);
and UO_2748 (O_2748,N_23769,N_24865);
xnor UO_2749 (O_2749,N_24636,N_24719);
nor UO_2750 (O_2750,N_24275,N_24518);
xnor UO_2751 (O_2751,N_24327,N_24456);
xnor UO_2752 (O_2752,N_23835,N_24990);
or UO_2753 (O_2753,N_24990,N_24352);
or UO_2754 (O_2754,N_24688,N_23835);
or UO_2755 (O_2755,N_24664,N_24501);
or UO_2756 (O_2756,N_24313,N_24849);
nor UO_2757 (O_2757,N_24463,N_24664);
nor UO_2758 (O_2758,N_24767,N_24902);
and UO_2759 (O_2759,N_24814,N_23754);
nor UO_2760 (O_2760,N_24454,N_24322);
or UO_2761 (O_2761,N_23806,N_23814);
nand UO_2762 (O_2762,N_23973,N_23770);
nand UO_2763 (O_2763,N_24047,N_24588);
xnor UO_2764 (O_2764,N_24238,N_24593);
xor UO_2765 (O_2765,N_24761,N_24705);
and UO_2766 (O_2766,N_23958,N_24310);
or UO_2767 (O_2767,N_23876,N_24853);
nand UO_2768 (O_2768,N_24715,N_24597);
nand UO_2769 (O_2769,N_24049,N_24670);
or UO_2770 (O_2770,N_24313,N_24528);
or UO_2771 (O_2771,N_24221,N_24025);
nor UO_2772 (O_2772,N_24168,N_24913);
and UO_2773 (O_2773,N_24221,N_23871);
xor UO_2774 (O_2774,N_23769,N_24930);
xor UO_2775 (O_2775,N_24742,N_23753);
nor UO_2776 (O_2776,N_24544,N_24066);
xor UO_2777 (O_2777,N_24905,N_24161);
nand UO_2778 (O_2778,N_24502,N_24060);
xnor UO_2779 (O_2779,N_24123,N_24809);
nand UO_2780 (O_2780,N_24234,N_24127);
and UO_2781 (O_2781,N_24824,N_24892);
nand UO_2782 (O_2782,N_24832,N_24114);
nor UO_2783 (O_2783,N_24018,N_24542);
nor UO_2784 (O_2784,N_23832,N_23872);
xnor UO_2785 (O_2785,N_24524,N_24621);
xnor UO_2786 (O_2786,N_24370,N_23853);
nor UO_2787 (O_2787,N_24260,N_23927);
and UO_2788 (O_2788,N_24752,N_24961);
or UO_2789 (O_2789,N_23763,N_24695);
xor UO_2790 (O_2790,N_24393,N_24055);
nand UO_2791 (O_2791,N_24875,N_24736);
and UO_2792 (O_2792,N_23847,N_24500);
or UO_2793 (O_2793,N_24834,N_23765);
and UO_2794 (O_2794,N_23968,N_23788);
nor UO_2795 (O_2795,N_24528,N_23760);
xor UO_2796 (O_2796,N_24898,N_24773);
and UO_2797 (O_2797,N_24501,N_24028);
or UO_2798 (O_2798,N_24403,N_23811);
xor UO_2799 (O_2799,N_24709,N_23969);
nand UO_2800 (O_2800,N_23800,N_24553);
xor UO_2801 (O_2801,N_24256,N_24148);
xor UO_2802 (O_2802,N_24904,N_24810);
and UO_2803 (O_2803,N_24446,N_24941);
and UO_2804 (O_2804,N_23868,N_24724);
xor UO_2805 (O_2805,N_24313,N_24578);
xor UO_2806 (O_2806,N_24292,N_23923);
nand UO_2807 (O_2807,N_24168,N_24468);
nor UO_2808 (O_2808,N_24661,N_24174);
nand UO_2809 (O_2809,N_24290,N_24992);
xor UO_2810 (O_2810,N_24296,N_24877);
xnor UO_2811 (O_2811,N_24373,N_24694);
xnor UO_2812 (O_2812,N_24232,N_24660);
xor UO_2813 (O_2813,N_24512,N_24071);
and UO_2814 (O_2814,N_24850,N_24751);
nand UO_2815 (O_2815,N_24943,N_24855);
nand UO_2816 (O_2816,N_24961,N_24885);
xor UO_2817 (O_2817,N_23987,N_24777);
xor UO_2818 (O_2818,N_24807,N_24997);
or UO_2819 (O_2819,N_24619,N_24558);
or UO_2820 (O_2820,N_24417,N_24101);
or UO_2821 (O_2821,N_24625,N_24172);
nand UO_2822 (O_2822,N_23959,N_24034);
nand UO_2823 (O_2823,N_24958,N_23808);
or UO_2824 (O_2824,N_23763,N_24558);
and UO_2825 (O_2825,N_24821,N_24301);
nor UO_2826 (O_2826,N_24140,N_24315);
nand UO_2827 (O_2827,N_23911,N_24197);
xor UO_2828 (O_2828,N_24659,N_23852);
nor UO_2829 (O_2829,N_24719,N_24733);
xor UO_2830 (O_2830,N_24193,N_23888);
or UO_2831 (O_2831,N_24283,N_24620);
xor UO_2832 (O_2832,N_24342,N_24162);
or UO_2833 (O_2833,N_23928,N_24711);
nor UO_2834 (O_2834,N_24161,N_24587);
or UO_2835 (O_2835,N_23857,N_24603);
nand UO_2836 (O_2836,N_23999,N_24282);
and UO_2837 (O_2837,N_24312,N_23957);
nor UO_2838 (O_2838,N_24669,N_24433);
or UO_2839 (O_2839,N_24598,N_24992);
nand UO_2840 (O_2840,N_24166,N_23834);
nand UO_2841 (O_2841,N_24518,N_24550);
nand UO_2842 (O_2842,N_24127,N_24660);
nand UO_2843 (O_2843,N_24017,N_24150);
xor UO_2844 (O_2844,N_24991,N_23981);
and UO_2845 (O_2845,N_24812,N_24179);
and UO_2846 (O_2846,N_24217,N_24346);
nor UO_2847 (O_2847,N_24255,N_24343);
nand UO_2848 (O_2848,N_24845,N_24162);
nand UO_2849 (O_2849,N_24605,N_24823);
xor UO_2850 (O_2850,N_23802,N_24573);
or UO_2851 (O_2851,N_24682,N_24336);
nor UO_2852 (O_2852,N_24732,N_23894);
nor UO_2853 (O_2853,N_24750,N_24986);
or UO_2854 (O_2854,N_24812,N_24902);
xor UO_2855 (O_2855,N_24460,N_24759);
nand UO_2856 (O_2856,N_23943,N_24269);
nor UO_2857 (O_2857,N_24248,N_24547);
nand UO_2858 (O_2858,N_24452,N_23961);
xor UO_2859 (O_2859,N_23791,N_24439);
nor UO_2860 (O_2860,N_24687,N_24766);
and UO_2861 (O_2861,N_23991,N_24940);
nand UO_2862 (O_2862,N_24364,N_24823);
xnor UO_2863 (O_2863,N_24801,N_24771);
and UO_2864 (O_2864,N_24001,N_24006);
or UO_2865 (O_2865,N_24923,N_24899);
or UO_2866 (O_2866,N_24241,N_24473);
xor UO_2867 (O_2867,N_23952,N_24444);
and UO_2868 (O_2868,N_24399,N_24575);
and UO_2869 (O_2869,N_24780,N_24261);
and UO_2870 (O_2870,N_24546,N_24222);
or UO_2871 (O_2871,N_24276,N_24016);
nor UO_2872 (O_2872,N_24379,N_23795);
and UO_2873 (O_2873,N_23977,N_23989);
and UO_2874 (O_2874,N_24943,N_24514);
and UO_2875 (O_2875,N_24837,N_24573);
and UO_2876 (O_2876,N_23818,N_24641);
and UO_2877 (O_2877,N_24200,N_24251);
nand UO_2878 (O_2878,N_24093,N_24554);
nand UO_2879 (O_2879,N_24132,N_24267);
nand UO_2880 (O_2880,N_24620,N_24609);
or UO_2881 (O_2881,N_24278,N_24520);
xor UO_2882 (O_2882,N_24335,N_24824);
nor UO_2883 (O_2883,N_24746,N_24782);
nor UO_2884 (O_2884,N_23765,N_24960);
and UO_2885 (O_2885,N_24831,N_24632);
nor UO_2886 (O_2886,N_23830,N_23770);
nor UO_2887 (O_2887,N_24337,N_24770);
xor UO_2888 (O_2888,N_24400,N_23835);
or UO_2889 (O_2889,N_24833,N_24352);
and UO_2890 (O_2890,N_24534,N_24085);
or UO_2891 (O_2891,N_24756,N_23898);
xnor UO_2892 (O_2892,N_24546,N_24983);
nand UO_2893 (O_2893,N_24242,N_24602);
nor UO_2894 (O_2894,N_24998,N_23775);
xor UO_2895 (O_2895,N_23774,N_24692);
and UO_2896 (O_2896,N_24230,N_24557);
or UO_2897 (O_2897,N_24801,N_24246);
xnor UO_2898 (O_2898,N_24410,N_24908);
nor UO_2899 (O_2899,N_24082,N_24309);
nand UO_2900 (O_2900,N_24851,N_24411);
or UO_2901 (O_2901,N_24720,N_24504);
nand UO_2902 (O_2902,N_24479,N_24679);
nand UO_2903 (O_2903,N_24418,N_23838);
or UO_2904 (O_2904,N_24140,N_24043);
nor UO_2905 (O_2905,N_24972,N_24518);
nor UO_2906 (O_2906,N_23817,N_24393);
or UO_2907 (O_2907,N_24100,N_24669);
xor UO_2908 (O_2908,N_24361,N_24873);
xnor UO_2909 (O_2909,N_24653,N_24085);
or UO_2910 (O_2910,N_24447,N_24322);
xnor UO_2911 (O_2911,N_24836,N_24599);
xnor UO_2912 (O_2912,N_24271,N_24820);
and UO_2913 (O_2913,N_24706,N_24109);
and UO_2914 (O_2914,N_24478,N_24832);
or UO_2915 (O_2915,N_24144,N_23901);
or UO_2916 (O_2916,N_24169,N_23853);
nor UO_2917 (O_2917,N_23879,N_24806);
nand UO_2918 (O_2918,N_24991,N_24932);
xor UO_2919 (O_2919,N_24914,N_24800);
nor UO_2920 (O_2920,N_24410,N_24690);
nand UO_2921 (O_2921,N_24984,N_24973);
nand UO_2922 (O_2922,N_24243,N_24895);
nand UO_2923 (O_2923,N_24342,N_24756);
nor UO_2924 (O_2924,N_24152,N_24709);
or UO_2925 (O_2925,N_24873,N_23833);
xnor UO_2926 (O_2926,N_23963,N_24261);
xor UO_2927 (O_2927,N_23858,N_23771);
and UO_2928 (O_2928,N_24934,N_23824);
nand UO_2929 (O_2929,N_24558,N_24127);
xor UO_2930 (O_2930,N_24197,N_24606);
or UO_2931 (O_2931,N_24010,N_24038);
and UO_2932 (O_2932,N_24116,N_24360);
nand UO_2933 (O_2933,N_24492,N_23756);
xnor UO_2934 (O_2934,N_24720,N_24709);
nor UO_2935 (O_2935,N_24664,N_24047);
and UO_2936 (O_2936,N_24320,N_24358);
xor UO_2937 (O_2937,N_24312,N_24529);
nor UO_2938 (O_2938,N_24501,N_24109);
or UO_2939 (O_2939,N_24600,N_24277);
xor UO_2940 (O_2940,N_24564,N_23760);
nand UO_2941 (O_2941,N_24089,N_23973);
xnor UO_2942 (O_2942,N_24855,N_24197);
and UO_2943 (O_2943,N_24374,N_24176);
xor UO_2944 (O_2944,N_24254,N_24641);
nor UO_2945 (O_2945,N_24558,N_24438);
xnor UO_2946 (O_2946,N_24562,N_24997);
or UO_2947 (O_2947,N_23996,N_24143);
nor UO_2948 (O_2948,N_24165,N_24561);
xnor UO_2949 (O_2949,N_24365,N_24534);
nand UO_2950 (O_2950,N_24298,N_24969);
and UO_2951 (O_2951,N_24317,N_23795);
or UO_2952 (O_2952,N_24049,N_24985);
and UO_2953 (O_2953,N_24497,N_24503);
and UO_2954 (O_2954,N_24180,N_24172);
nor UO_2955 (O_2955,N_24071,N_24384);
or UO_2956 (O_2956,N_24855,N_24779);
and UO_2957 (O_2957,N_24461,N_24641);
xnor UO_2958 (O_2958,N_24225,N_24736);
and UO_2959 (O_2959,N_24938,N_24366);
and UO_2960 (O_2960,N_24071,N_24663);
or UO_2961 (O_2961,N_24081,N_23799);
nor UO_2962 (O_2962,N_24437,N_24242);
nand UO_2963 (O_2963,N_23769,N_24713);
xnor UO_2964 (O_2964,N_24230,N_23982);
or UO_2965 (O_2965,N_24541,N_24719);
nor UO_2966 (O_2966,N_24614,N_23983);
and UO_2967 (O_2967,N_24016,N_24548);
nand UO_2968 (O_2968,N_24151,N_24248);
or UO_2969 (O_2969,N_24693,N_24790);
nand UO_2970 (O_2970,N_23995,N_23945);
or UO_2971 (O_2971,N_24924,N_23782);
nor UO_2972 (O_2972,N_24844,N_24188);
nor UO_2973 (O_2973,N_24854,N_24911);
and UO_2974 (O_2974,N_24922,N_23801);
nand UO_2975 (O_2975,N_24301,N_24166);
or UO_2976 (O_2976,N_24334,N_24078);
or UO_2977 (O_2977,N_24958,N_24094);
and UO_2978 (O_2978,N_24048,N_24707);
and UO_2979 (O_2979,N_24263,N_24171);
xor UO_2980 (O_2980,N_23829,N_24589);
and UO_2981 (O_2981,N_23767,N_24423);
nand UO_2982 (O_2982,N_24264,N_24531);
nor UO_2983 (O_2983,N_24381,N_24140);
nor UO_2984 (O_2984,N_24854,N_24735);
and UO_2985 (O_2985,N_24233,N_24443);
or UO_2986 (O_2986,N_23883,N_24065);
and UO_2987 (O_2987,N_24776,N_24495);
xnor UO_2988 (O_2988,N_24153,N_24025);
or UO_2989 (O_2989,N_24917,N_24044);
nand UO_2990 (O_2990,N_24902,N_23767);
nand UO_2991 (O_2991,N_24284,N_24230);
nor UO_2992 (O_2992,N_24391,N_24351);
or UO_2993 (O_2993,N_24414,N_24932);
nor UO_2994 (O_2994,N_24419,N_24353);
xor UO_2995 (O_2995,N_23795,N_24401);
nand UO_2996 (O_2996,N_24592,N_24109);
or UO_2997 (O_2997,N_24088,N_24341);
nand UO_2998 (O_2998,N_23987,N_24707);
nor UO_2999 (O_2999,N_24523,N_24071);
endmodule