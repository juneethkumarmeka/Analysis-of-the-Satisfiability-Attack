module basic_1500_15000_2000_3_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10003,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10013,N_10015,N_10018,N_10019,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10050,N_10051,N_10053,N_10054,N_10056,N_10058,N_10059,N_10060,N_10061,N_10062,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10076,N_10077,N_10079,N_10080,N_10081,N_10082,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10136,N_10137,N_10138,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10168,N_10170,N_10171,N_10172,N_10173,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10185,N_10186,N_10187,N_10189,N_10190,N_10192,N_10193,N_10194,N_10195,N_10196,N_10198,N_10199,N_10200,N_10201,N_10202,N_10204,N_10205,N_10206,N_10207,N_10208,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10238,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10247,N_10248,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10272,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10281,N_10283,N_10284,N_10285,N_10287,N_10288,N_10290,N_10291,N_10294,N_10295,N_10296,N_10297,N_10299,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10318,N_10321,N_10322,N_10323,N_10325,N_10327,N_10329,N_10330,N_10331,N_10332,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10342,N_10344,N_10345,N_10346,N_10348,N_10349,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10358,N_10359,N_10360,N_10361,N_10362,N_10365,N_10366,N_10367,N_10368,N_10369,N_10371,N_10372,N_10373,N_10374,N_10375,N_10377,N_10378,N_10381,N_10382,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10393,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10403,N_10406,N_10407,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10443,N_10444,N_10445,N_10447,N_10448,N_10449,N_10450,N_10452,N_10453,N_10454,N_10455,N_10456,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10469,N_10470,N_10471,N_10473,N_10474,N_10477,N_10478,N_10479,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10493,N_10494,N_10495,N_10498,N_10499,N_10500,N_10502,N_10503,N_10504,N_10505,N_10507,N_10508,N_10509,N_10512,N_10513,N_10514,N_10515,N_10517,N_10518,N_10519,N_10520,N_10522,N_10525,N_10526,N_10527,N_10529,N_10532,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10544,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10555,N_10557,N_10558,N_10560,N_10561,N_10562,N_10564,N_10565,N_10566,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10586,N_10587,N_10588,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10620,N_10621,N_10622,N_10623,N_10625,N_10629,N_10630,N_10632,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10642,N_10643,N_10646,N_10647,N_10650,N_10651,N_10653,N_10654,N_10655,N_10656,N_10657,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10667,N_10668,N_10669,N_10671,N_10672,N_10673,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10692,N_10693,N_10694,N_10695,N_10696,N_10699,N_10700,N_10701,N_10702,N_10703,N_10705,N_10706,N_10707,N_10708,N_10711,N_10712,N_10713,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10734,N_10735,N_10736,N_10737,N_10739,N_10741,N_10742,N_10743,N_10744,N_10745,N_10749,N_10751,N_10752,N_10753,N_10755,N_10757,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10774,N_10775,N_10776,N_10777,N_10778,N_10780,N_10781,N_10782,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10802,N_10803,N_10804,N_10805,N_10808,N_10810,N_10812,N_10814,N_10815,N_10816,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10846,N_10849,N_10851,N_10852,N_10853,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10903,N_10904,N_10905,N_10906,N_10908,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10923,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10950,N_10952,N_10953,N_10954,N_10955,N_10957,N_10958,N_10959,N_10960,N_10962,N_10965,N_10966,N_10967,N_10969,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10978,N_10979,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11010,N_11011,N_11012,N_11013,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11032,N_11033,N_11034,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11051,N_11053,N_11054,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11083,N_11084,N_11085,N_11086,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11104,N_11105,N_11106,N_11108,N_11111,N_11112,N_11113,N_11114,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11168,N_11169,N_11170,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11180,N_11181,N_11182,N_11184,N_11185,N_11186,N_11187,N_11188,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11205,N_11207,N_11208,N_11209,N_11211,N_11212,N_11213,N_11215,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11230,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11249,N_11251,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11262,N_11263,N_11264,N_11266,N_11267,N_11268,N_11270,N_11271,N_11272,N_11273,N_11276,N_11278,N_11279,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11299,N_11300,N_11301,N_11302,N_11303,N_11305,N_11306,N_11307,N_11308,N_11309,N_11311,N_11313,N_11315,N_11316,N_11317,N_11318,N_11319,N_11321,N_11322,N_11324,N_11326,N_11327,N_11329,N_11332,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11355,N_11357,N_11358,N_11360,N_11361,N_11362,N_11363,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11376,N_11377,N_11378,N_11380,N_11381,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11392,N_11393,N_11394,N_11395,N_11396,N_11400,N_11404,N_11405,N_11406,N_11407,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11442,N_11443,N_11444,N_11445,N_11446,N_11448,N_11449,N_11450,N_11451,N_11453,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11519,N_11520,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11532,N_11533,N_11534,N_11535,N_11539,N_11541,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11592,N_11593,N_11595,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11629,N_11630,N_11631,N_11632,N_11634,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11644,N_11645,N_11646,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11660,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11669,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11679,N_11680,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11727,N_11729,N_11730,N_11732,N_11735,N_11737,N_11738,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11747,N_11750,N_11751,N_11752,N_11754,N_11755,N_11757,N_11760,N_11762,N_11764,N_11765,N_11767,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11792,N_11793,N_11794,N_11796,N_11797,N_11800,N_11801,N_11803,N_11804,N_11807,N_11808,N_11809,N_11810,N_11812,N_11813,N_11814,N_11815,N_11816,N_11818,N_11819,N_11821,N_11823,N_11824,N_11825,N_11826,N_11828,N_11829,N_11830,N_11831,N_11833,N_11835,N_11836,N_11837,N_11838,N_11840,N_11842,N_11843,N_11846,N_11847,N_11848,N_11849,N_11851,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11862,N_11863,N_11864,N_11866,N_11867,N_11868,N_11869,N_11872,N_11873,N_11874,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11886,N_11887,N_11888,N_11889,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11899,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11909,N_11910,N_11913,N_11914,N_11916,N_11917,N_11918,N_11921,N_11922,N_11925,N_11926,N_11927,N_11930,N_11931,N_11932,N_11934,N_11936,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11953,N_11955,N_11956,N_11958,N_11959,N_11962,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12007,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12024,N_12025,N_12027,N_12028,N_12031,N_12032,N_12034,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12057,N_12058,N_12059,N_12060,N_12061,N_12063,N_12066,N_12067,N_12069,N_12070,N_12072,N_12073,N_12074,N_12076,N_12077,N_12078,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12103,N_12104,N_12105,N_12106,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12117,N_12119,N_12120,N_12121,N_12122,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12166,N_12167,N_12168,N_12169,N_12171,N_12172,N_12173,N_12174,N_12175,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12185,N_12186,N_12188,N_12189,N_12191,N_12192,N_12194,N_12195,N_12196,N_12199,N_12200,N_12202,N_12203,N_12204,N_12206,N_12207,N_12208,N_12210,N_12211,N_12213,N_12215,N_12216,N_12217,N_12218,N_12219,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12232,N_12233,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12257,N_12258,N_12259,N_12260,N_12261,N_12264,N_12266,N_12267,N_12268,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12283,N_12284,N_12287,N_12288,N_12291,N_12292,N_12293,N_12294,N_12296,N_12298,N_12299,N_12300,N_12301,N_12302,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12315,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12325,N_12328,N_12329,N_12330,N_12332,N_12333,N_12334,N_12335,N_12338,N_12339,N_12342,N_12343,N_12344,N_12346,N_12348,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12372,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12384,N_12385,N_12388,N_12389,N_12390,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12409,N_12410,N_12412,N_12414,N_12416,N_12417,N_12419,N_12420,N_12421,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12432,N_12435,N_12436,N_12437,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12452,N_12453,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12497,N_12498,N_12499,N_12500,N_12502,N_12503,N_12504,N_12505,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12515,N_12516,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12542,N_12543,N_12544,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12555,N_12556,N_12559,N_12560,N_12562,N_12563,N_12564,N_12567,N_12569,N_12570,N_12572,N_12573,N_12574,N_12575,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12589,N_12590,N_12591,N_12592,N_12594,N_12595,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12604,N_12605,N_12606,N_12607,N_12608,N_12610,N_12611,N_12612,N_12613,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12639,N_12641,N_12642,N_12643,N_12644,N_12646,N_12647,N_12648,N_12649,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12660,N_12661,N_12663,N_12664,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12702,N_12704,N_12705,N_12707,N_12710,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12757,N_12758,N_12760,N_12762,N_12763,N_12764,N_12766,N_12767,N_12768,N_12769,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12783,N_12784,N_12785,N_12786,N_12788,N_12791,N_12792,N_12793,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12809,N_12810,N_12811,N_12812,N_12813,N_12817,N_12818,N_12820,N_12821,N_12822,N_12824,N_12825,N_12826,N_12828,N_12829,N_12830,N_12832,N_12833,N_12834,N_12837,N_12838,N_12840,N_12841,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12857,N_12858,N_12859,N_12860,N_12862,N_12863,N_12864,N_12866,N_12868,N_12869,N_12870,N_12872,N_12873,N_12874,N_12875,N_12877,N_12878,N_12879,N_12880,N_12881,N_12885,N_12886,N_12887,N_12888,N_12889,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12928,N_12930,N_12931,N_12932,N_12934,N_12936,N_12937,N_12938,N_12939,N_12941,N_12942,N_12944,N_12945,N_12948,N_12949,N_12950,N_12951,N_12953,N_12954,N_12956,N_12957,N_12958,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12982,N_12983,N_12984,N_12985,N_12986,N_12988,N_12989,N_12991,N_12994,N_12996,N_12997,N_12998,N_12999,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13033,N_13035,N_13037,N_13038,N_13040,N_13041,N_13042,N_13044,N_13045,N_13046,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13095,N_13096,N_13097,N_13099,N_13100,N_13101,N_13105,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13128,N_13129,N_13130,N_13131,N_13132,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13157,N_13159,N_13160,N_13161,N_13162,N_13163,N_13166,N_13167,N_13168,N_13169,N_13171,N_13172,N_13173,N_13175,N_13176,N_13177,N_13179,N_13180,N_13181,N_13182,N_13183,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13211,N_13212,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13247,N_13248,N_13249,N_13250,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13265,N_13266,N_13268,N_13269,N_13270,N_13271,N_13272,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13281,N_13283,N_13284,N_13285,N_13287,N_13288,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13299,N_13300,N_13301,N_13303,N_13304,N_13305,N_13307,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13324,N_13325,N_13326,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13337,N_13339,N_13340,N_13341,N_13343,N_13344,N_13345,N_13346,N_13347,N_13349,N_13350,N_13352,N_13353,N_13354,N_13355,N_13357,N_13359,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13374,N_13375,N_13376,N_13378,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13392,N_13393,N_13394,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13411,N_13412,N_13414,N_13415,N_13416,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13432,N_13433,N_13434,N_13435,N_13436,N_13438,N_13440,N_13441,N_13442,N_13443,N_13444,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13492,N_13493,N_13494,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13512,N_13513,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13526,N_13527,N_13528,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13541,N_13542,N_13544,N_13545,N_13547,N_13549,N_13550,N_13551,N_13552,N_13553,N_13555,N_13556,N_13557,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13573,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13582,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13599,N_13603,N_13605,N_13606,N_13607,N_13609,N_13610,N_13612,N_13613,N_13614,N_13618,N_13619,N_13621,N_13624,N_13625,N_13627,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13656,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13671,N_13673,N_13675,N_13677,N_13678,N_13679,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13688,N_13689,N_13690,N_13691,N_13695,N_13696,N_13697,N_13699,N_13701,N_13702,N_13703,N_13704,N_13706,N_13707,N_13708,N_13711,N_13712,N_13713,N_13714,N_13715,N_13717,N_13718,N_13719,N_13720,N_13722,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13737,N_13740,N_13742,N_13743,N_13744,N_13745,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13760,N_13761,N_13762,N_13763,N_13765,N_13766,N_13767,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13778,N_13779,N_13780,N_13781,N_13783,N_13784,N_13785,N_13788,N_13789,N_13790,N_13794,N_13795,N_13796,N_13799,N_13800,N_13801,N_13802,N_13804,N_13805,N_13806,N_13808,N_13809,N_13811,N_13812,N_13813,N_13814,N_13815,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13824,N_13825,N_13826,N_13827,N_13830,N_13831,N_13832,N_13833,N_13834,N_13836,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13852,N_13853,N_13854,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13877,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13899,N_13900,N_13901,N_13902,N_13903,N_13905,N_13906,N_13908,N_13909,N_13910,N_13911,N_13914,N_13915,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13926,N_13927,N_13928,N_13929,N_13930,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13951,N_13952,N_13954,N_13955,N_13956,N_13957,N_13959,N_13960,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13993,N_13994,N_13995,N_13997,N_13998,N_13999,N_14000,N_14002,N_14004,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14016,N_14017,N_14019,N_14020,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14043,N_14044,N_14045,N_14047,N_14048,N_14049,N_14050,N_14051,N_14054,N_14055,N_14056,N_14057,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14071,N_14072,N_14073,N_14075,N_14076,N_14077,N_14080,N_14081,N_14082,N_14083,N_14084,N_14086,N_14087,N_14089,N_14090,N_14091,N_14092,N_14094,N_14096,N_14097,N_14099,N_14100,N_14101,N_14102,N_14103,N_14106,N_14107,N_14108,N_14109,N_14111,N_14112,N_14114,N_14115,N_14116,N_14117,N_14119,N_14120,N_14121,N_14122,N_14124,N_14125,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14168,N_14169,N_14171,N_14172,N_14173,N_14174,N_14176,N_14177,N_14178,N_14180,N_14181,N_14182,N_14183,N_14184,N_14186,N_14187,N_14189,N_14190,N_14192,N_14193,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14216,N_14217,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14241,N_14242,N_14244,N_14246,N_14248,N_14249,N_14250,N_14251,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14262,N_14263,N_14264,N_14266,N_14267,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14296,N_14297,N_14298,N_14299,N_14301,N_14302,N_14303,N_14304,N_14306,N_14307,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14317,N_14318,N_14319,N_14320,N_14321,N_14323,N_14325,N_14326,N_14327,N_14329,N_14330,N_14331,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14359,N_14362,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14381,N_14383,N_14385,N_14386,N_14388,N_14389,N_14390,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14400,N_14401,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14413,N_14414,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14432,N_14433,N_14434,N_14435,N_14437,N_14438,N_14439,N_14440,N_14443,N_14444,N_14446,N_14447,N_14449,N_14451,N_14452,N_14454,N_14455,N_14456,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14465,N_14466,N_14467,N_14468,N_14469,N_14471,N_14472,N_14473,N_14475,N_14476,N_14477,N_14478,N_14479,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14488,N_14489,N_14491,N_14492,N_14493,N_14494,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14537,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14565,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14579,N_14580,N_14581,N_14582,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14594,N_14595,N_14596,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14626,N_14627,N_14628,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14642,N_14643,N_14644,N_14645,N_14647,N_14648,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14660,N_14662,N_14663,N_14665,N_14666,N_14667,N_14668,N_14669,N_14672,N_14673,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14719,N_14720,N_14722,N_14723,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14735,N_14736,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14761,N_14762,N_14763,N_14764,N_14766,N_14767,N_14768,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14780,N_14783,N_14785,N_14786,N_14787,N_14788,N_14790,N_14791,N_14793,N_14794,N_14795,N_14796,N_14797,N_14799,N_14800,N_14801,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14837,N_14838,N_14840,N_14841,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14852,N_14854,N_14855,N_14856,N_14858,N_14861,N_14862,N_14863,N_14865,N_14866,N_14868,N_14869,N_14872,N_14873,N_14874,N_14875,N_14876,N_14879,N_14880,N_14882,N_14883,N_14884,N_14885,N_14886,N_14888,N_14889,N_14890,N_14891,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14914,N_14916,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14953,N_14954,N_14955,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14979,N_14980,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14989,N_14990,N_14991,N_14993,N_14995,N_14996,N_14997,N_14998;
nor U0 (N_0,In_347,In_382);
nand U1 (N_1,In_1399,In_607);
or U2 (N_2,In_462,In_1124);
and U3 (N_3,In_1389,In_744);
and U4 (N_4,In_1337,In_412);
nand U5 (N_5,In_1446,In_82);
nand U6 (N_6,In_123,In_1054);
nor U7 (N_7,In_118,In_863);
xor U8 (N_8,In_1155,In_1191);
nand U9 (N_9,In_513,In_1128);
or U10 (N_10,In_618,In_1434);
or U11 (N_11,In_1484,In_1037);
nand U12 (N_12,In_1022,In_1391);
and U13 (N_13,In_989,In_910);
and U14 (N_14,In_242,In_272);
or U15 (N_15,In_1060,In_569);
or U16 (N_16,In_348,In_909);
nor U17 (N_17,In_802,In_192);
or U18 (N_18,In_460,In_1439);
or U19 (N_19,In_851,In_1348);
nand U20 (N_20,In_938,In_1221);
nor U21 (N_21,In_270,In_817);
xnor U22 (N_22,In_93,In_772);
or U23 (N_23,In_905,In_1438);
nand U24 (N_24,In_1219,In_960);
or U25 (N_25,In_1359,In_1415);
xnor U26 (N_26,In_92,In_41);
or U27 (N_27,In_177,In_627);
nand U28 (N_28,In_346,In_1175);
nand U29 (N_29,In_1169,In_1338);
nor U30 (N_30,In_1021,In_444);
xnor U31 (N_31,In_259,In_117);
nand U32 (N_32,In_1067,In_266);
nand U33 (N_33,In_185,In_777);
and U34 (N_34,In_998,In_629);
or U35 (N_35,In_726,In_655);
nor U36 (N_36,In_367,In_1051);
and U37 (N_37,In_249,In_1308);
and U38 (N_38,In_958,In_856);
nor U39 (N_39,In_996,In_1422);
and U40 (N_40,In_575,In_309);
and U41 (N_41,In_1103,In_646);
nand U42 (N_42,In_790,In_49);
and U43 (N_43,In_1216,In_574);
or U44 (N_44,In_76,In_263);
and U45 (N_45,In_718,In_827);
and U46 (N_46,In_141,In_567);
xnor U47 (N_47,In_321,In_840);
nor U48 (N_48,In_1453,In_88);
nor U49 (N_49,In_872,In_690);
nand U50 (N_50,In_650,In_37);
xor U51 (N_51,In_12,In_68);
and U52 (N_52,In_787,In_763);
nor U53 (N_53,In_454,In_814);
or U54 (N_54,In_296,In_73);
nor U55 (N_55,In_605,In_1294);
and U56 (N_56,In_1218,In_286);
nor U57 (N_57,In_131,In_583);
and U58 (N_58,In_1290,In_712);
nor U59 (N_59,In_595,In_518);
or U60 (N_60,In_857,In_928);
or U61 (N_61,In_325,In_44);
nand U62 (N_62,In_868,In_694);
nand U63 (N_63,In_887,In_1233);
nand U64 (N_64,In_239,In_1393);
and U65 (N_65,In_1043,In_7);
and U66 (N_66,In_522,In_426);
nor U67 (N_67,In_1312,In_854);
or U68 (N_68,In_416,In_630);
nor U69 (N_69,In_870,In_1176);
and U70 (N_70,In_861,In_353);
and U71 (N_71,In_220,In_28);
and U72 (N_72,In_586,In_1072);
and U73 (N_73,In_838,In_734);
xnor U74 (N_74,In_439,In_1153);
and U75 (N_75,In_912,In_1199);
and U76 (N_76,In_788,In_1024);
nand U77 (N_77,In_980,In_431);
and U78 (N_78,In_722,In_458);
nand U79 (N_79,In_762,In_1227);
nand U80 (N_80,In_708,In_102);
and U81 (N_81,In_633,In_1088);
or U82 (N_82,In_1373,In_1419);
and U83 (N_83,In_893,In_1084);
nor U84 (N_84,In_1028,In_776);
nand U85 (N_85,In_1265,In_1397);
or U86 (N_86,In_359,In_810);
or U87 (N_87,In_345,In_297);
and U88 (N_88,In_1086,In_1135);
nor U89 (N_89,In_528,In_901);
or U90 (N_90,In_816,In_1421);
nand U91 (N_91,In_534,In_465);
nor U92 (N_92,In_248,In_149);
nand U93 (N_93,In_1098,In_157);
nor U94 (N_94,In_1363,In_723);
nand U95 (N_95,In_446,In_435);
and U96 (N_96,In_97,In_969);
nand U97 (N_97,In_16,In_742);
nand U98 (N_98,In_351,In_997);
nand U99 (N_99,In_1215,In_152);
nand U100 (N_100,In_1095,In_667);
and U101 (N_101,In_1370,In_1401);
nand U102 (N_102,In_873,In_1120);
nand U103 (N_103,In_1442,In_303);
nand U104 (N_104,In_70,In_882);
and U105 (N_105,In_393,In_933);
nor U106 (N_106,In_780,In_1466);
nand U107 (N_107,In_372,In_791);
and U108 (N_108,In_1435,In_792);
nor U109 (N_109,In_232,In_1297);
or U110 (N_110,In_1376,In_1033);
nand U111 (N_111,In_1092,In_251);
nor U112 (N_112,In_548,In_753);
nor U113 (N_113,In_1039,In_1230);
or U114 (N_114,In_824,In_294);
xnor U115 (N_115,In_908,In_778);
nor U116 (N_116,In_930,In_1057);
nand U117 (N_117,In_1104,In_927);
nand U118 (N_118,In_1427,In_561);
and U119 (N_119,In_1475,In_1240);
nor U120 (N_120,In_191,In_1330);
nand U121 (N_121,In_1300,In_628);
nor U122 (N_122,In_198,In_532);
nand U123 (N_123,In_622,In_413);
nand U124 (N_124,In_85,In_1059);
or U125 (N_125,In_179,In_1044);
and U126 (N_126,In_254,In_767);
xor U127 (N_127,In_1009,In_305);
or U128 (N_128,In_394,In_926);
nand U129 (N_129,In_1125,In_79);
nor U130 (N_130,In_890,In_621);
or U131 (N_131,In_965,In_992);
nand U132 (N_132,In_207,In_65);
or U133 (N_133,In_132,In_831);
nand U134 (N_134,In_13,In_530);
nand U135 (N_135,In_428,In_190);
nor U136 (N_136,In_836,In_715);
or U137 (N_137,In_150,In_1335);
nand U138 (N_138,In_1056,In_427);
nand U139 (N_139,In_658,In_830);
and U140 (N_140,In_1148,In_509);
and U141 (N_141,In_580,In_136);
nor U142 (N_142,In_611,In_91);
and U143 (N_143,In_373,In_1478);
nand U144 (N_144,In_707,In_119);
nand U145 (N_145,In_314,In_95);
and U146 (N_146,In_1274,In_1001);
or U147 (N_147,In_434,In_1226);
nand U148 (N_148,In_732,In_1350);
or U149 (N_149,In_892,In_1323);
or U150 (N_150,In_846,In_471);
or U151 (N_151,In_918,In_1333);
nor U152 (N_152,In_335,In_1203);
nor U153 (N_153,In_96,In_937);
nor U154 (N_154,In_796,In_1211);
and U155 (N_155,In_1400,In_649);
nand U156 (N_156,In_357,In_1412);
nand U157 (N_157,In_1473,In_915);
nor U158 (N_158,In_1096,In_1004);
and U159 (N_159,In_921,In_919);
or U160 (N_160,In_282,In_225);
xor U161 (N_161,In_120,In_1298);
and U162 (N_162,In_1161,In_1418);
nand U163 (N_163,In_779,In_1075);
nor U164 (N_164,In_758,In_109);
and U165 (N_165,In_663,In_344);
and U166 (N_166,In_8,In_299);
or U167 (N_167,In_875,In_1118);
and U168 (N_168,In_1015,In_236);
xor U169 (N_169,In_1186,In_645);
xnor U170 (N_170,In_542,In_1451);
and U171 (N_171,In_932,In_804);
nand U172 (N_172,In_57,In_322);
nor U173 (N_173,In_1137,In_1185);
nor U174 (N_174,In_1388,In_565);
or U175 (N_175,In_167,In_702);
xor U176 (N_176,In_420,In_80);
or U177 (N_177,In_525,In_886);
and U178 (N_178,In_1055,In_1027);
or U179 (N_179,In_175,In_328);
and U180 (N_180,In_67,In_963);
nor U181 (N_181,In_124,In_404);
or U182 (N_182,In_623,In_964);
nand U183 (N_183,In_337,In_637);
nor U184 (N_184,In_809,In_409);
or U185 (N_185,In_324,In_769);
xor U186 (N_186,In_793,In_1117);
nand U187 (N_187,In_255,In_436);
and U188 (N_188,In_631,In_51);
nor U189 (N_189,In_539,In_237);
nand U190 (N_190,In_484,In_1487);
and U191 (N_191,In_1119,In_724);
nor U192 (N_192,In_1102,In_1229);
nand U193 (N_193,In_654,In_62);
nand U194 (N_194,In_20,In_288);
nor U195 (N_195,In_46,In_1132);
nor U196 (N_196,In_601,In_292);
or U197 (N_197,In_1005,In_23);
nand U198 (N_198,In_1089,In_786);
nor U199 (N_199,In_1485,In_799);
nor U200 (N_200,In_293,In_1481);
nor U201 (N_201,In_1077,In_1101);
nand U202 (N_202,In_1193,In_1319);
or U203 (N_203,In_826,In_1352);
or U204 (N_204,In_774,In_544);
nor U205 (N_205,In_1177,In_839);
and U206 (N_206,In_449,In_1408);
nand U207 (N_207,In_1224,In_1301);
or U208 (N_208,In_201,In_952);
nand U209 (N_209,In_1020,In_706);
or U210 (N_210,In_163,In_1204);
and U211 (N_211,In_193,In_1431);
nor U212 (N_212,In_1303,In_1188);
nand U213 (N_213,In_865,In_822);
nor U214 (N_214,In_1242,In_476);
or U215 (N_215,In_538,In_835);
nor U216 (N_216,In_593,In_990);
nand U217 (N_217,In_140,In_687);
and U218 (N_218,In_129,In_1183);
and U219 (N_219,In_273,In_1390);
nor U220 (N_220,In_1375,In_456);
nor U221 (N_221,In_447,In_130);
nand U222 (N_222,In_874,In_1074);
xnor U223 (N_223,In_766,In_159);
nand U224 (N_224,In_966,In_913);
or U225 (N_225,In_1450,In_1404);
or U226 (N_226,In_470,In_626);
nand U227 (N_227,In_589,In_747);
nand U228 (N_228,In_323,In_664);
and U229 (N_229,In_1269,In_222);
and U230 (N_230,In_1272,In_1430);
or U231 (N_231,In_1029,In_1209);
nor U232 (N_232,In_699,In_356);
nand U233 (N_233,In_1249,In_741);
and U234 (N_234,In_1355,In_1336);
nand U235 (N_235,In_160,In_659);
and U236 (N_236,In_1257,In_98);
or U237 (N_237,In_227,In_11);
or U238 (N_238,In_591,In_620);
or U239 (N_239,In_155,In_1049);
nor U240 (N_240,In_1491,In_1220);
nor U241 (N_241,In_986,In_1315);
and U242 (N_242,In_147,In_1472);
or U243 (N_243,In_78,In_1267);
and U244 (N_244,In_452,In_939);
and U245 (N_245,In_527,In_1141);
or U246 (N_246,In_955,In_579);
nand U247 (N_247,In_582,In_541);
nand U248 (N_248,In_504,In_704);
or U249 (N_249,In_729,In_1144);
and U250 (N_250,In_257,In_594);
or U251 (N_251,In_1392,In_494);
nor U252 (N_252,In_405,In_1032);
or U253 (N_253,In_1261,In_615);
nand U254 (N_254,In_445,In_858);
and U255 (N_255,In_376,In_738);
nand U256 (N_256,In_543,In_843);
or U257 (N_257,In_540,In_492);
or U258 (N_258,In_670,In_1405);
nand U259 (N_259,In_1202,In_1052);
or U260 (N_260,In_829,In_716);
nand U261 (N_261,In_1073,In_1357);
xnor U262 (N_262,In_570,In_949);
or U263 (N_263,In_896,In_226);
and U264 (N_264,In_230,In_14);
and U265 (N_265,In_987,In_978);
nor U266 (N_266,In_678,In_54);
or U267 (N_267,In_1429,In_246);
and U268 (N_268,In_110,In_1035);
and U269 (N_269,In_925,In_1080);
and U270 (N_270,In_21,In_186);
nor U271 (N_271,In_338,In_339);
or U272 (N_272,In_1413,In_797);
nor U273 (N_273,In_250,In_180);
and U274 (N_274,In_2,In_1443);
nor U275 (N_275,In_847,In_1011);
and U276 (N_276,In_154,In_508);
nor U277 (N_277,In_1150,In_114);
or U278 (N_278,In_1234,In_64);
nor U279 (N_279,In_52,In_1156);
xnor U280 (N_280,In_768,In_22);
and U281 (N_281,In_1471,In_1470);
nor U282 (N_282,In_889,In_1034);
and U283 (N_283,In_143,In_825);
nor U284 (N_284,In_69,In_247);
nor U285 (N_285,In_1332,In_173);
nor U286 (N_286,In_648,In_1414);
nor U287 (N_287,In_1147,In_184);
nand U288 (N_288,In_264,In_1048);
and U289 (N_289,In_602,In_811);
xnor U290 (N_290,In_521,In_1174);
nand U291 (N_291,In_1255,In_1476);
and U292 (N_292,In_1007,In_488);
nor U293 (N_293,In_940,In_1127);
nand U294 (N_294,In_318,In_657);
nor U295 (N_295,In_461,In_695);
and U296 (N_296,In_1152,In_1016);
and U297 (N_297,In_1410,In_1146);
or U298 (N_298,In_312,In_578);
nor U299 (N_299,In_487,In_1163);
xnor U300 (N_300,In_1126,In_1154);
nand U301 (N_301,In_832,In_1407);
nor U302 (N_302,In_782,In_951);
and U303 (N_303,In_1469,In_481);
and U304 (N_304,In_438,In_343);
and U305 (N_305,In_676,In_402);
and U306 (N_306,In_24,In_174);
or U307 (N_307,In_677,In_950);
or U308 (N_308,In_877,In_453);
nand U309 (N_309,In_210,In_153);
nand U310 (N_310,In_441,In_166);
and U311 (N_311,In_641,In_619);
and U312 (N_312,In_25,In_1441);
and U313 (N_313,In_585,In_1142);
nand U314 (N_314,In_17,In_27);
or U315 (N_315,In_517,In_1346);
and U316 (N_316,In_979,In_970);
nor U317 (N_317,In_243,In_26);
and U318 (N_318,In_1479,In_1483);
nor U319 (N_319,In_466,In_475);
and U320 (N_320,In_422,In_1395);
nand U321 (N_321,In_1061,In_1214);
nor U322 (N_322,In_924,In_479);
nor U323 (N_323,In_599,In_410);
nor U324 (N_324,In_756,In_1110);
and U325 (N_325,In_505,In_498);
nor U326 (N_326,In_1396,In_515);
xor U327 (N_327,In_1107,In_168);
and U328 (N_328,In_137,In_1365);
or U329 (N_329,In_1166,In_821);
or U330 (N_330,In_386,In_1480);
and U331 (N_331,In_789,In_749);
nor U332 (N_332,In_1258,In_682);
and U333 (N_333,In_1090,In_1256);
and U334 (N_334,In_581,In_467);
nand U335 (N_335,In_472,In_423);
or U336 (N_336,In_1381,In_943);
nor U337 (N_337,In_898,In_904);
and U338 (N_338,In_134,In_1378);
and U339 (N_339,In_1030,In_1010);
and U340 (N_340,In_418,In_770);
nand U341 (N_341,In_976,In_1130);
nor U342 (N_342,In_1042,In_1490);
nor U343 (N_343,In_1179,In_746);
and U344 (N_344,In_956,In_946);
nand U345 (N_345,In_361,In_1322);
nand U346 (N_346,In_30,In_1235);
and U347 (N_347,In_354,In_1063);
nand U348 (N_348,In_430,In_1239);
nand U349 (N_349,In_1444,In_1122);
nand U350 (N_350,In_1069,In_665);
and U351 (N_351,In_944,In_316);
nor U352 (N_352,In_1356,In_662);
or U353 (N_353,In_1428,In_1138);
nand U354 (N_354,In_1496,In_995);
nand U355 (N_355,In_135,In_278);
xor U356 (N_356,In_693,In_375);
or U357 (N_357,In_634,In_233);
and U358 (N_358,In_358,In_1078);
nor U359 (N_359,In_692,In_116);
and U360 (N_360,In_100,In_1313);
or U361 (N_361,In_698,In_823);
or U362 (N_362,In_514,In_1447);
and U363 (N_363,In_1279,In_537);
or U364 (N_364,In_231,In_75);
or U365 (N_365,In_1133,In_878);
nor U366 (N_366,In_884,In_1123);
and U367 (N_367,In_1082,In_1171);
nand U368 (N_368,In_568,In_1286);
and U369 (N_369,In_267,In_253);
nor U370 (N_370,In_1053,In_176);
and U371 (N_371,In_837,In_397);
nor U372 (N_372,In_326,In_962);
nor U373 (N_373,In_72,In_258);
nand U374 (N_374,In_696,In_374);
nand U375 (N_375,In_262,In_571);
and U376 (N_376,In_240,In_604);
or U377 (N_377,In_674,In_1454);
or U378 (N_378,In_99,In_1276);
xor U379 (N_379,In_371,In_188);
xor U380 (N_380,In_1423,In_564);
or U381 (N_381,In_686,In_108);
nor U382 (N_382,In_573,In_871);
nand U383 (N_383,In_614,In_32);
or U384 (N_384,In_355,In_761);
and U385 (N_385,In_590,In_365);
nor U386 (N_386,In_603,In_833);
nor U387 (N_387,In_562,In_388);
and U388 (N_388,In_883,In_828);
nand U389 (N_389,In_1383,In_274);
or U390 (N_390,In_547,In_598);
or U391 (N_391,In_1231,In_384);
xnor U392 (N_392,In_380,In_464);
nand U393 (N_393,In_608,In_636);
nor U394 (N_394,In_881,In_1246);
nor U395 (N_395,In_1417,In_9);
and U396 (N_396,In_477,In_1482);
or U397 (N_397,In_1071,In_1262);
or U398 (N_398,In_496,In_1099);
nand U399 (N_399,In_94,In_256);
nand U400 (N_400,In_1266,In_731);
or U401 (N_401,In_424,In_760);
nor U402 (N_402,In_1145,In_317);
nand U403 (N_403,In_34,In_442);
or U404 (N_404,In_204,In_1081);
nor U405 (N_405,In_183,In_531);
nand U406 (N_406,In_480,In_1302);
or U407 (N_407,In_957,In_1164);
xnor U408 (N_408,In_443,In_209);
nor U409 (N_409,In_1468,In_647);
nand U410 (N_410,In_87,In_31);
or U411 (N_411,In_35,In_1380);
nand U412 (N_412,In_511,In_350);
or U413 (N_413,In_15,In_377);
and U414 (N_414,In_985,In_178);
and U415 (N_415,In_50,In_869);
or U416 (N_416,In_879,In_369);
nand U417 (N_417,In_1025,In_1304);
nand U418 (N_418,In_287,In_224);
nor U419 (N_419,In_917,In_818);
or U420 (N_420,In_520,In_228);
nor U421 (N_421,In_500,In_425);
or U422 (N_422,In_3,In_281);
or U423 (N_423,In_406,In_1345);
and U424 (N_424,In_523,In_302);
nor U425 (N_425,In_429,In_74);
nor U426 (N_426,In_1361,In_1498);
nand U427 (N_427,In_205,In_1244);
and U428 (N_428,In_490,In_971);
and U429 (N_429,In_1046,In_360);
and U430 (N_430,In_922,In_491);
nand U431 (N_431,In_945,In_66);
and U432 (N_432,In_680,In_319);
and U433 (N_433,In_5,In_1349);
nand U434 (N_434,In_988,In_592);
nor U435 (N_435,In_1283,In_1343);
and U436 (N_436,In_625,In_895);
nor U437 (N_437,In_493,In_679);
nand U438 (N_438,In_1190,In_151);
nand U439 (N_439,In_867,In_300);
or U440 (N_440,In_333,In_862);
or U441 (N_441,In_1178,In_284);
nor U442 (N_442,In_550,In_1003);
nand U443 (N_443,In_1347,In_39);
and U444 (N_444,In_1328,In_666);
nand U445 (N_445,In_1091,In_1317);
nor U446 (N_446,In_553,In_414);
nor U447 (N_447,In_451,In_991);
or U448 (N_448,In_165,In_1432);
and U449 (N_449,In_701,In_1288);
nor U450 (N_450,In_310,In_1206);
or U451 (N_451,In_398,In_203);
and U452 (N_452,In_391,In_1426);
nand U453 (N_453,In_880,In_1452);
nand U454 (N_454,In_888,In_936);
nand U455 (N_455,In_58,In_735);
nand U456 (N_456,In_145,In_171);
nor U457 (N_457,In_463,In_1050);
nor U458 (N_458,In_1372,In_983);
and U459 (N_459,In_1340,In_1253);
nand U460 (N_460,In_215,In_1382);
and U461 (N_461,In_685,In_1094);
nand U462 (N_462,In_489,In_1192);
nor U463 (N_463,In_683,In_967);
nor U464 (N_464,In_1324,In_751);
nor U465 (N_465,In_211,In_162);
or U466 (N_466,In_390,In_408);
nor U467 (N_467,In_59,In_352);
nor U468 (N_468,In_1109,In_1486);
nor U469 (N_469,In_334,In_1411);
nand U470 (N_470,In_1305,In_813);
nand U471 (N_471,In_546,In_1275);
nand U472 (N_472,In_1116,In_221);
nor U473 (N_473,In_1198,In_387);
nor U474 (N_474,In_276,In_340);
and U475 (N_475,In_557,In_1263);
or U476 (N_476,In_1284,In_703);
or U477 (N_477,In_617,In_1160);
and U478 (N_478,In_1097,In_1217);
or U479 (N_479,In_1368,In_241);
nor U480 (N_480,In_808,In_1331);
nor U481 (N_481,In_1207,In_364);
nor U482 (N_482,In_600,In_947);
or U483 (N_483,In_1321,In_512);
xor U484 (N_484,In_849,In_697);
and U485 (N_485,In_19,In_1247);
nor U486 (N_486,In_954,In_1031);
or U487 (N_487,In_53,In_1318);
and U488 (N_488,In_1165,In_757);
and U489 (N_489,In_1248,In_1225);
or U490 (N_490,In_238,In_745);
or U491 (N_491,In_1041,In_469);
nor U492 (N_492,In_642,In_1136);
nand U493 (N_493,In_1477,In_1433);
or U494 (N_494,In_1111,In_497);
and U495 (N_495,In_681,In_612);
nor U496 (N_496,In_56,In_1344);
or U497 (N_497,In_781,In_771);
nor U498 (N_498,In_315,In_473);
nor U499 (N_499,In_1013,In_725);
nor U500 (N_500,In_60,In_349);
nand U501 (N_501,In_1377,In_1366);
and U502 (N_502,In_1351,In_639);
nor U503 (N_503,In_1083,In_336);
and U504 (N_504,In_651,In_805);
nor U505 (N_505,In_653,In_311);
or U506 (N_506,In_122,In_214);
and U507 (N_507,In_440,In_1341);
and U508 (N_508,In_306,In_1353);
nand U509 (N_509,In_320,In_342);
or U510 (N_510,In_914,In_169);
nand U511 (N_511,In_803,In_40);
or U512 (N_512,In_545,In_529);
nor U513 (N_513,In_616,In_1173);
and U514 (N_514,In_133,In_717);
or U515 (N_515,In_411,In_448);
and U516 (N_516,In_216,In_399);
nor U517 (N_517,In_164,In_977);
nand U518 (N_518,In_268,In_610);
nand U519 (N_519,In_111,In_1222);
or U520 (N_520,In_982,In_968);
nand U521 (N_521,In_18,In_1062);
nor U522 (N_522,In_219,In_999);
nand U523 (N_523,In_125,In_891);
and U524 (N_524,In_644,In_669);
nand U525 (N_525,In_1131,In_172);
nor U526 (N_526,In_1306,In_860);
nor U527 (N_527,In_450,In_42);
and U528 (N_528,In_554,In_127);
or U529 (N_529,In_1232,In_1384);
nand U530 (N_530,In_55,In_1162);
nand U531 (N_531,In_672,In_1108);
or U532 (N_532,In_486,In_392);
nand U533 (N_533,In_533,In_1014);
nand U534 (N_534,In_596,In_1143);
nor U535 (N_535,In_1311,In_126);
nand U536 (N_536,In_104,In_43);
or U537 (N_537,In_1100,In_6);
and U538 (N_538,In_820,In_1236);
or U539 (N_539,In_283,In_1364);
nor U540 (N_540,In_1445,In_1342);
nor U541 (N_541,In_1440,In_229);
and U542 (N_542,In_1181,In_588);
or U543 (N_543,In_743,In_1189);
and U544 (N_544,In_506,In_510);
nand U545 (N_545,In_1325,In_1187);
and U546 (N_546,In_437,In_298);
or U547 (N_547,In_1403,In_916);
or U548 (N_548,In_1065,In_848);
nor U549 (N_549,In_139,In_1172);
nor U550 (N_550,In_341,In_1168);
and U551 (N_551,In_265,In_0);
or U552 (N_552,In_923,In_1458);
and U553 (N_553,In_332,In_313);
and U554 (N_554,In_1245,In_1197);
xnor U555 (N_555,In_714,In_536);
and U556 (N_556,In_483,In_417);
and U557 (N_557,In_107,In_1134);
and U558 (N_558,In_535,In_502);
or U559 (N_559,In_948,In_555);
nor U560 (N_560,In_1070,In_941);
and U561 (N_561,In_785,In_841);
nand U562 (N_562,In_1437,In_584);
or U563 (N_563,In_1006,In_81);
nand U564 (N_564,In_395,In_208);
nor U565 (N_565,In_721,In_433);
nor U566 (N_566,In_1281,In_700);
nand U567 (N_567,In_212,In_1296);
nor U568 (N_568,In_1292,In_689);
or U569 (N_569,In_223,In_1264);
or U570 (N_570,In_806,In_113);
nand U571 (N_571,In_1260,In_1406);
or U572 (N_572,In_89,In_245);
nor U573 (N_573,In_834,In_606);
or U574 (N_574,In_1316,In_1463);
nor U575 (N_575,In_432,In_482);
and U576 (N_576,In_260,In_736);
nor U577 (N_577,In_1114,In_684);
nand U578 (N_578,In_170,In_876);
or U579 (N_579,In_1358,In_269);
and U580 (N_580,In_773,In_552);
and U581 (N_581,In_844,In_643);
nand U582 (N_582,In_1492,In_984);
nor U583 (N_583,In_1210,In_1494);
nor U584 (N_584,In_1208,In_934);
nand U585 (N_585,In_1314,In_1259);
nand U586 (N_586,In_1295,In_800);
or U587 (N_587,In_1309,In_187);
nand U588 (N_588,In_711,In_289);
nor U589 (N_589,In_457,In_1310);
nand U590 (N_590,In_194,In_1008);
and U591 (N_591,In_556,In_1115);
or U592 (N_592,In_688,In_519);
nand U593 (N_593,In_279,In_362);
or U594 (N_594,In_1416,In_1019);
nand U595 (N_595,In_71,In_327);
nand U596 (N_596,In_1238,In_1237);
nor U597 (N_597,In_1170,In_1448);
and U598 (N_598,In_400,In_1002);
and U599 (N_599,In_572,In_1398);
nand U600 (N_600,In_727,In_271);
nor U601 (N_601,In_1273,In_29);
or U602 (N_602,In_981,In_1461);
xnor U603 (N_603,In_1385,In_1113);
nor U604 (N_604,In_1,In_182);
or U605 (N_605,In_752,In_739);
and U606 (N_606,In_864,In_795);
nor U607 (N_607,In_842,In_304);
and U608 (N_608,In_1277,In_624);
nor U609 (N_609,In_640,In_115);
nor U610 (N_610,In_1299,In_1334);
nor U611 (N_611,In_244,In_911);
nor U612 (N_612,In_1287,In_558);
nand U613 (N_613,In_1394,In_161);
and U614 (N_614,In_1449,In_1205);
nor U615 (N_615,In_1038,In_1149);
nor U616 (N_616,In_1329,In_1360);
or U617 (N_617,In_368,In_801);
nand U618 (N_618,In_784,In_1252);
nor U619 (N_619,In_1326,In_112);
or U620 (N_620,In_1018,In_994);
and U621 (N_621,In_1106,In_1497);
and U622 (N_622,In_524,In_366);
nand U623 (N_623,In_798,In_10);
nor U624 (N_624,In_705,In_48);
nand U625 (N_625,In_1036,In_755);
nor U626 (N_626,In_1362,In_1489);
nand U627 (N_627,In_1464,In_1420);
and U628 (N_628,In_907,In_1462);
nor U629 (N_629,In_106,In_148);
or U630 (N_630,In_1465,In_559);
nand U631 (N_631,In_195,In_485);
nor U632 (N_632,In_128,In_47);
nand U633 (N_633,In_993,In_507);
or U634 (N_634,In_855,In_903);
and U635 (N_635,In_1369,In_403);
and U636 (N_636,In_459,In_894);
and U637 (N_637,In_1167,In_121);
nor U638 (N_638,In_859,In_455);
nand U639 (N_639,In_206,In_549);
nand U640 (N_640,In_261,In_577);
or U641 (N_641,In_1327,In_144);
nor U642 (N_642,In_710,In_635);
and U643 (N_643,In_381,In_45);
nor U644 (N_644,In_199,In_83);
nor U645 (N_645,In_234,In_1047);
or U646 (N_646,In_1271,In_733);
nor U647 (N_647,In_217,In_1139);
and U648 (N_648,In_526,In_1474);
nor U649 (N_649,In_363,In_389);
nand U650 (N_650,In_1243,In_1387);
nand U651 (N_651,In_1158,In_33);
or U652 (N_652,In_906,In_419);
and U653 (N_653,In_61,In_942);
and U654 (N_654,In_301,In_807);
nor U655 (N_655,In_407,In_560);
and U656 (N_656,In_501,In_218);
and U657 (N_657,In_90,In_421);
xor U658 (N_658,In_1354,In_675);
and U659 (N_659,In_295,In_1251);
nor U660 (N_660,In_385,In_516);
nor U661 (N_661,In_1112,In_1409);
and U662 (N_662,In_1129,In_1012);
nand U663 (N_663,In_158,In_973);
and U664 (N_664,In_1105,In_379);
nand U665 (N_665,In_728,In_1068);
or U666 (N_666,In_1157,In_4);
and U667 (N_667,In_401,In_931);
or U668 (N_668,In_638,In_36);
or U669 (N_669,In_1087,In_783);
xor U670 (N_670,In_1402,In_1184);
nor U671 (N_671,In_897,In_1307);
nand U672 (N_672,In_1151,In_920);
or U673 (N_673,In_1223,In_63);
nand U674 (N_674,In_1201,In_566);
and U675 (N_675,In_1268,In_1250);
or U676 (N_676,In_1140,In_1459);
nand U677 (N_677,In_1093,In_331);
nor U678 (N_678,In_415,In_748);
nor U679 (N_679,In_576,In_754);
nand U680 (N_680,In_101,In_750);
nand U681 (N_681,In_972,In_277);
or U682 (N_682,In_252,In_759);
or U683 (N_683,In_1159,In_1493);
nand U684 (N_684,In_656,In_866);
or U685 (N_685,In_961,In_77);
nor U686 (N_686,In_899,In_1495);
nor U687 (N_687,In_1456,In_935);
nand U688 (N_688,In_1371,In_142);
nand U689 (N_689,In_1291,In_1285);
nor U690 (N_690,In_1064,In_885);
and U691 (N_691,In_765,In_1289);
or U692 (N_692,In_671,In_474);
or U693 (N_693,In_1499,In_730);
and U694 (N_694,In_138,In_383);
or U695 (N_695,In_1367,In_551);
nor U696 (N_696,In_953,In_1079);
or U697 (N_697,In_202,In_563);
or U698 (N_698,In_1200,In_1282);
or U699 (N_699,In_1374,In_632);
nand U700 (N_700,In_673,In_329);
or U701 (N_701,In_1436,In_86);
and U702 (N_702,In_38,In_1066);
nor U703 (N_703,In_396,In_613);
and U704 (N_704,In_1085,In_275);
or U705 (N_705,In_1040,In_290);
nor U706 (N_706,In_587,In_1241);
nor U707 (N_707,In_609,In_850);
xnor U708 (N_708,In_189,In_1467);
and U709 (N_709,In_815,In_196);
and U710 (N_710,In_794,In_975);
and U711 (N_711,In_291,In_1212);
nand U712 (N_712,In_330,In_1339);
and U713 (N_713,In_929,In_959);
nand U714 (N_714,In_1195,In_495);
nor U715 (N_715,In_307,In_1228);
and U716 (N_716,In_285,In_974);
and U717 (N_717,In_764,In_853);
nand U718 (N_718,In_845,In_1000);
and U719 (N_719,In_280,In_308);
or U720 (N_720,In_1278,In_105);
or U721 (N_721,In_235,In_1424);
and U722 (N_722,In_1488,In_819);
nor U723 (N_723,In_197,In_103);
or U724 (N_724,In_740,In_503);
nor U725 (N_725,In_737,In_1058);
nand U726 (N_726,In_156,In_478);
nor U727 (N_727,In_1213,In_84);
or U728 (N_728,In_1076,In_370);
and U729 (N_729,In_1045,In_661);
or U730 (N_730,In_181,In_1121);
nand U731 (N_731,In_146,In_709);
and U732 (N_732,In_691,In_1457);
or U733 (N_733,In_852,In_378);
or U734 (N_734,In_1460,In_1023);
nand U735 (N_735,In_812,In_597);
nor U736 (N_736,In_668,In_1386);
nand U737 (N_737,In_468,In_499);
or U738 (N_738,In_1182,In_652);
and U739 (N_739,In_1280,In_1320);
nor U740 (N_740,In_1425,In_900);
nand U741 (N_741,In_775,In_1196);
xor U742 (N_742,In_660,In_1026);
or U743 (N_743,In_1017,In_1293);
or U744 (N_744,In_1455,In_720);
nand U745 (N_745,In_1270,In_213);
and U746 (N_746,In_719,In_1194);
or U747 (N_747,In_1254,In_713);
nor U748 (N_748,In_200,In_1180);
or U749 (N_749,In_902,In_1379);
nand U750 (N_750,In_690,In_149);
or U751 (N_751,In_1025,In_36);
or U752 (N_752,In_1154,In_149);
xor U753 (N_753,In_502,In_650);
or U754 (N_754,In_31,In_1145);
xnor U755 (N_755,In_601,In_1223);
nand U756 (N_756,In_1275,In_141);
nor U757 (N_757,In_287,In_676);
or U758 (N_758,In_406,In_1201);
or U759 (N_759,In_334,In_627);
nand U760 (N_760,In_43,In_648);
nor U761 (N_761,In_1494,In_727);
or U762 (N_762,In_1056,In_414);
nand U763 (N_763,In_286,In_728);
and U764 (N_764,In_1362,In_1225);
nand U765 (N_765,In_1421,In_472);
or U766 (N_766,In_566,In_98);
nor U767 (N_767,In_461,In_178);
nor U768 (N_768,In_552,In_418);
nor U769 (N_769,In_970,In_260);
nor U770 (N_770,In_95,In_164);
and U771 (N_771,In_872,In_532);
nand U772 (N_772,In_520,In_193);
and U773 (N_773,In_802,In_238);
nor U774 (N_774,In_411,In_701);
nor U775 (N_775,In_1184,In_1112);
or U776 (N_776,In_1260,In_1277);
and U777 (N_777,In_1419,In_1187);
nor U778 (N_778,In_291,In_1317);
and U779 (N_779,In_1269,In_599);
nor U780 (N_780,In_1463,In_111);
nand U781 (N_781,In_1360,In_260);
nor U782 (N_782,In_893,In_454);
nor U783 (N_783,In_1167,In_1166);
or U784 (N_784,In_453,In_733);
nor U785 (N_785,In_863,In_1097);
or U786 (N_786,In_327,In_680);
nor U787 (N_787,In_199,In_225);
and U788 (N_788,In_504,In_692);
and U789 (N_789,In_1394,In_426);
nand U790 (N_790,In_1331,In_463);
and U791 (N_791,In_1403,In_498);
and U792 (N_792,In_876,In_889);
or U793 (N_793,In_663,In_485);
nor U794 (N_794,In_1277,In_1170);
nand U795 (N_795,In_400,In_588);
nor U796 (N_796,In_1099,In_1168);
nand U797 (N_797,In_1352,In_1079);
and U798 (N_798,In_900,In_983);
xnor U799 (N_799,In_1178,In_1059);
nand U800 (N_800,In_735,In_138);
or U801 (N_801,In_521,In_1461);
nand U802 (N_802,In_1290,In_159);
and U803 (N_803,In_1075,In_307);
and U804 (N_804,In_613,In_178);
nand U805 (N_805,In_355,In_1379);
nand U806 (N_806,In_902,In_800);
nand U807 (N_807,In_1147,In_120);
nand U808 (N_808,In_1211,In_651);
nor U809 (N_809,In_769,In_1193);
or U810 (N_810,In_190,In_1074);
nor U811 (N_811,In_1472,In_1060);
nand U812 (N_812,In_1139,In_874);
or U813 (N_813,In_852,In_271);
nand U814 (N_814,In_1033,In_979);
and U815 (N_815,In_1461,In_221);
nand U816 (N_816,In_330,In_1331);
or U817 (N_817,In_687,In_427);
nand U818 (N_818,In_434,In_1340);
and U819 (N_819,In_534,In_160);
nor U820 (N_820,In_364,In_913);
or U821 (N_821,In_930,In_1160);
or U822 (N_822,In_1459,In_1296);
or U823 (N_823,In_708,In_1210);
or U824 (N_824,In_1477,In_967);
nor U825 (N_825,In_569,In_976);
nor U826 (N_826,In_771,In_328);
or U827 (N_827,In_1012,In_404);
or U828 (N_828,In_147,In_426);
nor U829 (N_829,In_1213,In_50);
or U830 (N_830,In_83,In_53);
nand U831 (N_831,In_1412,In_1484);
nand U832 (N_832,In_208,In_784);
nand U833 (N_833,In_1166,In_205);
and U834 (N_834,In_1245,In_224);
nor U835 (N_835,In_933,In_28);
or U836 (N_836,In_1082,In_436);
or U837 (N_837,In_231,In_840);
and U838 (N_838,In_642,In_551);
or U839 (N_839,In_710,In_469);
and U840 (N_840,In_691,In_252);
or U841 (N_841,In_803,In_168);
and U842 (N_842,In_262,In_1126);
nand U843 (N_843,In_140,In_577);
nand U844 (N_844,In_1255,In_746);
nand U845 (N_845,In_547,In_763);
or U846 (N_846,In_1424,In_671);
nand U847 (N_847,In_720,In_700);
nor U848 (N_848,In_1222,In_1389);
or U849 (N_849,In_289,In_895);
nor U850 (N_850,In_762,In_635);
and U851 (N_851,In_312,In_87);
nand U852 (N_852,In_1137,In_312);
or U853 (N_853,In_1404,In_500);
nand U854 (N_854,In_938,In_284);
and U855 (N_855,In_391,In_637);
and U856 (N_856,In_1467,In_990);
and U857 (N_857,In_1186,In_1333);
nor U858 (N_858,In_1374,In_887);
nor U859 (N_859,In_664,In_799);
nand U860 (N_860,In_1092,In_564);
and U861 (N_861,In_1100,In_897);
nand U862 (N_862,In_1113,In_33);
and U863 (N_863,In_1298,In_251);
or U864 (N_864,In_206,In_986);
and U865 (N_865,In_186,In_377);
nor U866 (N_866,In_838,In_1069);
or U867 (N_867,In_1112,In_1089);
nand U868 (N_868,In_979,In_23);
nor U869 (N_869,In_1460,In_749);
nand U870 (N_870,In_1418,In_990);
or U871 (N_871,In_515,In_316);
or U872 (N_872,In_948,In_363);
or U873 (N_873,In_1383,In_949);
xnor U874 (N_874,In_1296,In_1188);
or U875 (N_875,In_1248,In_347);
nor U876 (N_876,In_1291,In_307);
nor U877 (N_877,In_1335,In_1423);
nor U878 (N_878,In_313,In_864);
or U879 (N_879,In_166,In_688);
and U880 (N_880,In_583,In_963);
nand U881 (N_881,In_1092,In_1238);
nand U882 (N_882,In_207,In_137);
nand U883 (N_883,In_366,In_499);
or U884 (N_884,In_17,In_439);
and U885 (N_885,In_136,In_77);
nand U886 (N_886,In_1139,In_1236);
nand U887 (N_887,In_415,In_1435);
nor U888 (N_888,In_621,In_166);
nand U889 (N_889,In_1284,In_1192);
or U890 (N_890,In_925,In_1216);
nor U891 (N_891,In_990,In_55);
nor U892 (N_892,In_1035,In_1125);
nor U893 (N_893,In_608,In_1433);
and U894 (N_894,In_1122,In_516);
or U895 (N_895,In_1291,In_395);
and U896 (N_896,In_76,In_1377);
nor U897 (N_897,In_687,In_317);
nor U898 (N_898,In_1135,In_1318);
nor U899 (N_899,In_829,In_1383);
nand U900 (N_900,In_1440,In_1454);
nor U901 (N_901,In_382,In_1192);
nor U902 (N_902,In_661,In_1285);
nand U903 (N_903,In_1403,In_483);
nor U904 (N_904,In_547,In_1459);
or U905 (N_905,In_855,In_908);
nor U906 (N_906,In_594,In_132);
and U907 (N_907,In_914,In_976);
xor U908 (N_908,In_1144,In_1307);
and U909 (N_909,In_1097,In_691);
or U910 (N_910,In_147,In_252);
nand U911 (N_911,In_844,In_850);
nor U912 (N_912,In_549,In_746);
nor U913 (N_913,In_467,In_1428);
nor U914 (N_914,In_1447,In_808);
and U915 (N_915,In_467,In_468);
or U916 (N_916,In_800,In_980);
xnor U917 (N_917,In_1374,In_665);
nor U918 (N_918,In_266,In_763);
and U919 (N_919,In_579,In_1478);
and U920 (N_920,In_701,In_109);
and U921 (N_921,In_57,In_1284);
and U922 (N_922,In_626,In_1374);
and U923 (N_923,In_1118,In_386);
nor U924 (N_924,In_1039,In_1302);
and U925 (N_925,In_266,In_700);
and U926 (N_926,In_376,In_283);
nand U927 (N_927,In_1057,In_940);
and U928 (N_928,In_508,In_1368);
nand U929 (N_929,In_447,In_1231);
or U930 (N_930,In_1349,In_403);
or U931 (N_931,In_662,In_552);
nand U932 (N_932,In_400,In_40);
or U933 (N_933,In_101,In_297);
nor U934 (N_934,In_1212,In_532);
or U935 (N_935,In_964,In_188);
and U936 (N_936,In_714,In_684);
or U937 (N_937,In_1470,In_508);
and U938 (N_938,In_1112,In_963);
or U939 (N_939,In_473,In_1034);
and U940 (N_940,In_642,In_1070);
or U941 (N_941,In_880,In_1267);
or U942 (N_942,In_1132,In_309);
or U943 (N_943,In_192,In_1440);
or U944 (N_944,In_1411,In_1480);
nor U945 (N_945,In_1172,In_66);
or U946 (N_946,In_647,In_716);
and U947 (N_947,In_1297,In_1063);
and U948 (N_948,In_1083,In_297);
and U949 (N_949,In_1392,In_1414);
nor U950 (N_950,In_1474,In_7);
nand U951 (N_951,In_332,In_193);
or U952 (N_952,In_890,In_614);
nor U953 (N_953,In_1312,In_67);
nor U954 (N_954,In_1314,In_395);
or U955 (N_955,In_1469,In_1179);
nand U956 (N_956,In_188,In_1477);
or U957 (N_957,In_217,In_837);
and U958 (N_958,In_501,In_1209);
nand U959 (N_959,In_263,In_1285);
nand U960 (N_960,In_129,In_674);
and U961 (N_961,In_538,In_875);
or U962 (N_962,In_708,In_616);
and U963 (N_963,In_625,In_677);
nand U964 (N_964,In_938,In_1374);
and U965 (N_965,In_431,In_1364);
and U966 (N_966,In_564,In_1274);
and U967 (N_967,In_1226,In_524);
nand U968 (N_968,In_318,In_167);
xor U969 (N_969,In_760,In_787);
or U970 (N_970,In_1249,In_264);
or U971 (N_971,In_1340,In_1087);
nand U972 (N_972,In_1053,In_251);
nor U973 (N_973,In_220,In_995);
or U974 (N_974,In_646,In_1207);
nand U975 (N_975,In_1167,In_208);
nor U976 (N_976,In_1043,In_1205);
nor U977 (N_977,In_705,In_915);
or U978 (N_978,In_1171,In_916);
and U979 (N_979,In_79,In_740);
and U980 (N_980,In_1232,In_898);
or U981 (N_981,In_216,In_1307);
and U982 (N_982,In_885,In_903);
nor U983 (N_983,In_834,In_1237);
or U984 (N_984,In_180,In_1495);
and U985 (N_985,In_1274,In_751);
nand U986 (N_986,In_911,In_869);
and U987 (N_987,In_32,In_372);
and U988 (N_988,In_1417,In_879);
nand U989 (N_989,In_846,In_1136);
xnor U990 (N_990,In_694,In_466);
nand U991 (N_991,In_158,In_665);
and U992 (N_992,In_471,In_201);
nor U993 (N_993,In_1418,In_205);
nor U994 (N_994,In_479,In_1039);
nor U995 (N_995,In_929,In_805);
xor U996 (N_996,In_18,In_76);
and U997 (N_997,In_928,In_1487);
and U998 (N_998,In_334,In_1295);
nor U999 (N_999,In_1252,In_1116);
nand U1000 (N_1000,In_255,In_202);
and U1001 (N_1001,In_156,In_692);
and U1002 (N_1002,In_708,In_449);
and U1003 (N_1003,In_843,In_503);
nand U1004 (N_1004,In_808,In_908);
and U1005 (N_1005,In_356,In_713);
nor U1006 (N_1006,In_1285,In_320);
or U1007 (N_1007,In_1106,In_604);
xor U1008 (N_1008,In_1109,In_137);
nor U1009 (N_1009,In_176,In_425);
or U1010 (N_1010,In_468,In_130);
and U1011 (N_1011,In_625,In_1141);
nor U1012 (N_1012,In_734,In_78);
and U1013 (N_1013,In_123,In_917);
nand U1014 (N_1014,In_367,In_89);
nor U1015 (N_1015,In_138,In_402);
or U1016 (N_1016,In_1402,In_1326);
and U1017 (N_1017,In_485,In_847);
and U1018 (N_1018,In_228,In_943);
nor U1019 (N_1019,In_325,In_871);
nand U1020 (N_1020,In_1340,In_904);
nor U1021 (N_1021,In_448,In_739);
or U1022 (N_1022,In_585,In_1140);
nor U1023 (N_1023,In_1142,In_392);
and U1024 (N_1024,In_1185,In_1164);
or U1025 (N_1025,In_94,In_1416);
and U1026 (N_1026,In_729,In_1319);
nor U1027 (N_1027,In_380,In_695);
nand U1028 (N_1028,In_566,In_1445);
nor U1029 (N_1029,In_696,In_87);
or U1030 (N_1030,In_149,In_408);
and U1031 (N_1031,In_1291,In_116);
and U1032 (N_1032,In_1220,In_159);
nand U1033 (N_1033,In_376,In_1175);
nand U1034 (N_1034,In_717,In_758);
or U1035 (N_1035,In_1182,In_706);
or U1036 (N_1036,In_225,In_706);
xor U1037 (N_1037,In_5,In_929);
or U1038 (N_1038,In_148,In_219);
nand U1039 (N_1039,In_1086,In_348);
and U1040 (N_1040,In_674,In_73);
or U1041 (N_1041,In_648,In_446);
or U1042 (N_1042,In_673,In_166);
and U1043 (N_1043,In_386,In_394);
nand U1044 (N_1044,In_842,In_930);
nand U1045 (N_1045,In_3,In_1194);
and U1046 (N_1046,In_1454,In_367);
or U1047 (N_1047,In_1048,In_1174);
and U1048 (N_1048,In_348,In_1114);
and U1049 (N_1049,In_729,In_911);
or U1050 (N_1050,In_414,In_630);
nand U1051 (N_1051,In_1215,In_260);
and U1052 (N_1052,In_1164,In_348);
or U1053 (N_1053,In_84,In_546);
or U1054 (N_1054,In_654,In_1264);
nor U1055 (N_1055,In_1401,In_854);
xor U1056 (N_1056,In_1054,In_896);
or U1057 (N_1057,In_956,In_1021);
or U1058 (N_1058,In_1171,In_64);
nand U1059 (N_1059,In_1286,In_398);
nor U1060 (N_1060,In_401,In_349);
nor U1061 (N_1061,In_26,In_45);
nor U1062 (N_1062,In_1030,In_1350);
or U1063 (N_1063,In_1274,In_1087);
nand U1064 (N_1064,In_498,In_973);
and U1065 (N_1065,In_502,In_660);
nor U1066 (N_1066,In_367,In_281);
and U1067 (N_1067,In_434,In_509);
nand U1068 (N_1068,In_519,In_913);
nand U1069 (N_1069,In_1080,In_1230);
and U1070 (N_1070,In_629,In_850);
xnor U1071 (N_1071,In_837,In_1495);
and U1072 (N_1072,In_1418,In_1283);
nor U1073 (N_1073,In_519,In_348);
nand U1074 (N_1074,In_1481,In_9);
and U1075 (N_1075,In_1398,In_1335);
and U1076 (N_1076,In_263,In_1409);
nand U1077 (N_1077,In_1314,In_799);
or U1078 (N_1078,In_992,In_1138);
and U1079 (N_1079,In_865,In_1478);
nand U1080 (N_1080,In_130,In_865);
nand U1081 (N_1081,In_1210,In_1361);
nor U1082 (N_1082,In_963,In_1297);
and U1083 (N_1083,In_318,In_645);
nor U1084 (N_1084,In_319,In_475);
nand U1085 (N_1085,In_588,In_99);
nor U1086 (N_1086,In_327,In_693);
nand U1087 (N_1087,In_537,In_373);
and U1088 (N_1088,In_695,In_169);
nor U1089 (N_1089,In_467,In_630);
xor U1090 (N_1090,In_641,In_1263);
and U1091 (N_1091,In_896,In_337);
or U1092 (N_1092,In_244,In_833);
or U1093 (N_1093,In_692,In_1302);
and U1094 (N_1094,In_968,In_326);
xor U1095 (N_1095,In_1088,In_1492);
nor U1096 (N_1096,In_159,In_1264);
nor U1097 (N_1097,In_443,In_899);
nor U1098 (N_1098,In_624,In_812);
nand U1099 (N_1099,In_1312,In_113);
and U1100 (N_1100,In_456,In_873);
nor U1101 (N_1101,In_198,In_1207);
or U1102 (N_1102,In_861,In_1168);
nor U1103 (N_1103,In_669,In_504);
or U1104 (N_1104,In_37,In_813);
nor U1105 (N_1105,In_1140,In_1288);
nand U1106 (N_1106,In_1407,In_1049);
nand U1107 (N_1107,In_1121,In_515);
or U1108 (N_1108,In_270,In_340);
or U1109 (N_1109,In_1376,In_1253);
and U1110 (N_1110,In_1065,In_456);
nor U1111 (N_1111,In_1098,In_1015);
nand U1112 (N_1112,In_578,In_1395);
nand U1113 (N_1113,In_22,In_979);
or U1114 (N_1114,In_441,In_324);
nor U1115 (N_1115,In_363,In_498);
or U1116 (N_1116,In_359,In_984);
nor U1117 (N_1117,In_51,In_92);
nand U1118 (N_1118,In_1070,In_968);
nand U1119 (N_1119,In_535,In_1031);
nor U1120 (N_1120,In_591,In_883);
xor U1121 (N_1121,In_1470,In_1056);
and U1122 (N_1122,In_1477,In_629);
nand U1123 (N_1123,In_33,In_535);
and U1124 (N_1124,In_807,In_809);
nand U1125 (N_1125,In_756,In_960);
or U1126 (N_1126,In_786,In_602);
nand U1127 (N_1127,In_1479,In_1095);
nand U1128 (N_1128,In_1098,In_1114);
nor U1129 (N_1129,In_578,In_1342);
nand U1130 (N_1130,In_1275,In_1417);
nand U1131 (N_1131,In_977,In_1331);
or U1132 (N_1132,In_1291,In_711);
nor U1133 (N_1133,In_105,In_151);
nor U1134 (N_1134,In_23,In_157);
or U1135 (N_1135,In_702,In_1474);
nand U1136 (N_1136,In_369,In_1022);
nand U1137 (N_1137,In_601,In_575);
and U1138 (N_1138,In_4,In_97);
nand U1139 (N_1139,In_1016,In_781);
or U1140 (N_1140,In_99,In_1446);
and U1141 (N_1141,In_217,In_1485);
and U1142 (N_1142,In_1062,In_1447);
nand U1143 (N_1143,In_533,In_400);
nand U1144 (N_1144,In_802,In_564);
or U1145 (N_1145,In_70,In_1488);
nand U1146 (N_1146,In_1020,In_1361);
and U1147 (N_1147,In_1238,In_143);
nand U1148 (N_1148,In_463,In_1158);
nor U1149 (N_1149,In_367,In_617);
or U1150 (N_1150,In_1240,In_466);
or U1151 (N_1151,In_245,In_1458);
or U1152 (N_1152,In_930,In_827);
nor U1153 (N_1153,In_434,In_796);
and U1154 (N_1154,In_201,In_73);
or U1155 (N_1155,In_1142,In_324);
and U1156 (N_1156,In_372,In_862);
or U1157 (N_1157,In_1454,In_237);
nand U1158 (N_1158,In_117,In_335);
and U1159 (N_1159,In_306,In_1381);
xor U1160 (N_1160,In_881,In_1171);
nor U1161 (N_1161,In_867,In_258);
nand U1162 (N_1162,In_552,In_913);
xor U1163 (N_1163,In_989,In_1119);
nand U1164 (N_1164,In_139,In_283);
nand U1165 (N_1165,In_377,In_332);
nor U1166 (N_1166,In_458,In_1333);
nor U1167 (N_1167,In_1079,In_691);
and U1168 (N_1168,In_917,In_956);
and U1169 (N_1169,In_508,In_1445);
nand U1170 (N_1170,In_646,In_568);
nor U1171 (N_1171,In_200,In_1154);
or U1172 (N_1172,In_1398,In_134);
or U1173 (N_1173,In_209,In_1004);
nand U1174 (N_1174,In_1087,In_536);
and U1175 (N_1175,In_323,In_573);
nor U1176 (N_1176,In_1405,In_250);
nor U1177 (N_1177,In_1142,In_445);
nand U1178 (N_1178,In_1129,In_246);
or U1179 (N_1179,In_108,In_963);
nand U1180 (N_1180,In_1365,In_444);
nor U1181 (N_1181,In_1120,In_1223);
nand U1182 (N_1182,In_1051,In_423);
nand U1183 (N_1183,In_417,In_789);
nand U1184 (N_1184,In_399,In_140);
or U1185 (N_1185,In_959,In_664);
nor U1186 (N_1186,In_1419,In_1077);
xor U1187 (N_1187,In_316,In_522);
nor U1188 (N_1188,In_636,In_274);
or U1189 (N_1189,In_932,In_376);
nor U1190 (N_1190,In_778,In_554);
nand U1191 (N_1191,In_178,In_1347);
nand U1192 (N_1192,In_974,In_875);
nor U1193 (N_1193,In_805,In_820);
xnor U1194 (N_1194,In_680,In_624);
nor U1195 (N_1195,In_146,In_358);
nand U1196 (N_1196,In_967,In_1009);
and U1197 (N_1197,In_458,In_165);
nand U1198 (N_1198,In_1337,In_318);
xnor U1199 (N_1199,In_789,In_250);
nor U1200 (N_1200,In_1449,In_967);
and U1201 (N_1201,In_739,In_46);
nand U1202 (N_1202,In_1277,In_71);
or U1203 (N_1203,In_1420,In_1319);
and U1204 (N_1204,In_620,In_976);
nor U1205 (N_1205,In_868,In_1143);
nor U1206 (N_1206,In_835,In_845);
or U1207 (N_1207,In_452,In_734);
nand U1208 (N_1208,In_1033,In_237);
nand U1209 (N_1209,In_861,In_588);
nor U1210 (N_1210,In_847,In_1465);
or U1211 (N_1211,In_450,In_823);
and U1212 (N_1212,In_337,In_1083);
and U1213 (N_1213,In_668,In_1185);
and U1214 (N_1214,In_519,In_871);
nor U1215 (N_1215,In_1305,In_20);
and U1216 (N_1216,In_344,In_300);
xnor U1217 (N_1217,In_80,In_389);
nor U1218 (N_1218,In_1063,In_194);
nor U1219 (N_1219,In_340,In_375);
nand U1220 (N_1220,In_730,In_532);
nor U1221 (N_1221,In_840,In_612);
nand U1222 (N_1222,In_639,In_720);
nor U1223 (N_1223,In_982,In_458);
xor U1224 (N_1224,In_1042,In_116);
and U1225 (N_1225,In_1047,In_1062);
or U1226 (N_1226,In_1031,In_545);
nand U1227 (N_1227,In_377,In_628);
nor U1228 (N_1228,In_796,In_395);
and U1229 (N_1229,In_1124,In_67);
or U1230 (N_1230,In_419,In_1116);
or U1231 (N_1231,In_1246,In_277);
nand U1232 (N_1232,In_688,In_867);
nand U1233 (N_1233,In_1181,In_1309);
nor U1234 (N_1234,In_306,In_150);
nor U1235 (N_1235,In_1246,In_552);
and U1236 (N_1236,In_553,In_1441);
and U1237 (N_1237,In_499,In_1099);
nand U1238 (N_1238,In_452,In_671);
and U1239 (N_1239,In_871,In_146);
nand U1240 (N_1240,In_389,In_905);
xnor U1241 (N_1241,In_1389,In_898);
and U1242 (N_1242,In_396,In_370);
nor U1243 (N_1243,In_553,In_904);
and U1244 (N_1244,In_1426,In_306);
nor U1245 (N_1245,In_965,In_925);
and U1246 (N_1246,In_220,In_149);
nor U1247 (N_1247,In_420,In_671);
and U1248 (N_1248,In_64,In_87);
or U1249 (N_1249,In_1436,In_215);
nand U1250 (N_1250,In_899,In_1191);
nand U1251 (N_1251,In_529,In_1344);
or U1252 (N_1252,In_427,In_84);
and U1253 (N_1253,In_1333,In_681);
nand U1254 (N_1254,In_867,In_1318);
nor U1255 (N_1255,In_1363,In_1358);
or U1256 (N_1256,In_1224,In_618);
nor U1257 (N_1257,In_1016,In_371);
xnor U1258 (N_1258,In_186,In_1156);
nor U1259 (N_1259,In_998,In_337);
and U1260 (N_1260,In_171,In_1262);
or U1261 (N_1261,In_241,In_541);
or U1262 (N_1262,In_1025,In_1371);
nor U1263 (N_1263,In_1373,In_298);
and U1264 (N_1264,In_893,In_487);
or U1265 (N_1265,In_905,In_314);
nor U1266 (N_1266,In_475,In_415);
nor U1267 (N_1267,In_252,In_780);
nor U1268 (N_1268,In_1223,In_1347);
nand U1269 (N_1269,In_836,In_1324);
nand U1270 (N_1270,In_794,In_1036);
nand U1271 (N_1271,In_1459,In_238);
nand U1272 (N_1272,In_102,In_24);
nand U1273 (N_1273,In_738,In_486);
nor U1274 (N_1274,In_1068,In_180);
nor U1275 (N_1275,In_1255,In_659);
nand U1276 (N_1276,In_835,In_1265);
or U1277 (N_1277,In_1494,In_1282);
and U1278 (N_1278,In_1148,In_872);
and U1279 (N_1279,In_622,In_964);
or U1280 (N_1280,In_399,In_1281);
nand U1281 (N_1281,In_118,In_318);
nand U1282 (N_1282,In_124,In_1096);
nand U1283 (N_1283,In_884,In_1338);
nand U1284 (N_1284,In_1284,In_436);
nor U1285 (N_1285,In_99,In_12);
nand U1286 (N_1286,In_1007,In_75);
nand U1287 (N_1287,In_1309,In_475);
nor U1288 (N_1288,In_42,In_1012);
or U1289 (N_1289,In_691,In_447);
or U1290 (N_1290,In_755,In_179);
and U1291 (N_1291,In_1430,In_423);
or U1292 (N_1292,In_1476,In_987);
nor U1293 (N_1293,In_1399,In_807);
and U1294 (N_1294,In_1465,In_130);
or U1295 (N_1295,In_651,In_666);
nand U1296 (N_1296,In_308,In_1468);
nor U1297 (N_1297,In_498,In_371);
xor U1298 (N_1298,In_866,In_834);
nor U1299 (N_1299,In_1302,In_869);
and U1300 (N_1300,In_433,In_91);
nand U1301 (N_1301,In_633,In_332);
nor U1302 (N_1302,In_1170,In_246);
or U1303 (N_1303,In_69,In_649);
nor U1304 (N_1304,In_714,In_309);
nand U1305 (N_1305,In_180,In_451);
nor U1306 (N_1306,In_749,In_292);
or U1307 (N_1307,In_1024,In_530);
and U1308 (N_1308,In_469,In_864);
nor U1309 (N_1309,In_722,In_971);
nor U1310 (N_1310,In_641,In_533);
nand U1311 (N_1311,In_788,In_375);
and U1312 (N_1312,In_1122,In_1003);
and U1313 (N_1313,In_1496,In_1387);
nor U1314 (N_1314,In_1396,In_239);
or U1315 (N_1315,In_650,In_599);
and U1316 (N_1316,In_223,In_744);
or U1317 (N_1317,In_1023,In_77);
nand U1318 (N_1318,In_82,In_1148);
nand U1319 (N_1319,In_25,In_1112);
and U1320 (N_1320,In_1175,In_583);
nand U1321 (N_1321,In_53,In_1293);
nand U1322 (N_1322,In_1286,In_754);
nand U1323 (N_1323,In_31,In_1371);
and U1324 (N_1324,In_11,In_690);
nand U1325 (N_1325,In_651,In_401);
or U1326 (N_1326,In_341,In_106);
nor U1327 (N_1327,In_617,In_1055);
nor U1328 (N_1328,In_792,In_197);
nand U1329 (N_1329,In_1205,In_279);
or U1330 (N_1330,In_1110,In_185);
or U1331 (N_1331,In_966,In_531);
nor U1332 (N_1332,In_829,In_857);
nor U1333 (N_1333,In_888,In_74);
and U1334 (N_1334,In_1316,In_45);
nor U1335 (N_1335,In_376,In_1369);
nand U1336 (N_1336,In_1376,In_847);
or U1337 (N_1337,In_500,In_802);
or U1338 (N_1338,In_414,In_1203);
or U1339 (N_1339,In_1319,In_159);
nand U1340 (N_1340,In_880,In_1476);
nor U1341 (N_1341,In_1377,In_869);
or U1342 (N_1342,In_1257,In_637);
nand U1343 (N_1343,In_671,In_1197);
and U1344 (N_1344,In_140,In_1445);
nand U1345 (N_1345,In_971,In_131);
or U1346 (N_1346,In_1000,In_1266);
or U1347 (N_1347,In_471,In_649);
nor U1348 (N_1348,In_281,In_1494);
nand U1349 (N_1349,In_1099,In_449);
and U1350 (N_1350,In_80,In_1116);
or U1351 (N_1351,In_497,In_180);
nor U1352 (N_1352,In_1047,In_940);
nand U1353 (N_1353,In_665,In_751);
nand U1354 (N_1354,In_626,In_654);
or U1355 (N_1355,In_1305,In_49);
nand U1356 (N_1356,In_356,In_850);
and U1357 (N_1357,In_661,In_508);
or U1358 (N_1358,In_920,In_461);
and U1359 (N_1359,In_1187,In_641);
xor U1360 (N_1360,In_478,In_493);
nor U1361 (N_1361,In_769,In_130);
or U1362 (N_1362,In_517,In_858);
and U1363 (N_1363,In_82,In_523);
and U1364 (N_1364,In_562,In_1408);
or U1365 (N_1365,In_200,In_920);
nor U1366 (N_1366,In_0,In_1090);
and U1367 (N_1367,In_899,In_123);
and U1368 (N_1368,In_205,In_624);
nand U1369 (N_1369,In_1481,In_799);
or U1370 (N_1370,In_150,In_145);
nor U1371 (N_1371,In_240,In_1295);
nand U1372 (N_1372,In_322,In_488);
xor U1373 (N_1373,In_267,In_508);
or U1374 (N_1374,In_283,In_285);
nor U1375 (N_1375,In_800,In_637);
nor U1376 (N_1376,In_585,In_125);
or U1377 (N_1377,In_357,In_516);
nor U1378 (N_1378,In_720,In_771);
nor U1379 (N_1379,In_769,In_268);
and U1380 (N_1380,In_779,In_1245);
nor U1381 (N_1381,In_181,In_618);
or U1382 (N_1382,In_929,In_1396);
nand U1383 (N_1383,In_879,In_41);
nor U1384 (N_1384,In_769,In_423);
and U1385 (N_1385,In_1465,In_1370);
or U1386 (N_1386,In_92,In_1103);
nand U1387 (N_1387,In_428,In_1463);
and U1388 (N_1388,In_104,In_117);
nand U1389 (N_1389,In_274,In_567);
xor U1390 (N_1390,In_1416,In_615);
nor U1391 (N_1391,In_1430,In_600);
and U1392 (N_1392,In_204,In_1279);
and U1393 (N_1393,In_1133,In_907);
or U1394 (N_1394,In_786,In_1473);
nor U1395 (N_1395,In_967,In_1148);
nor U1396 (N_1396,In_450,In_1413);
and U1397 (N_1397,In_761,In_210);
or U1398 (N_1398,In_1490,In_1403);
or U1399 (N_1399,In_1296,In_1051);
nor U1400 (N_1400,In_1317,In_1089);
and U1401 (N_1401,In_1329,In_843);
or U1402 (N_1402,In_1060,In_309);
and U1403 (N_1403,In_46,In_877);
nand U1404 (N_1404,In_314,In_477);
nor U1405 (N_1405,In_482,In_472);
and U1406 (N_1406,In_853,In_636);
nor U1407 (N_1407,In_168,In_293);
nor U1408 (N_1408,In_1040,In_558);
or U1409 (N_1409,In_21,In_887);
nor U1410 (N_1410,In_178,In_129);
nor U1411 (N_1411,In_914,In_262);
or U1412 (N_1412,In_585,In_1301);
nor U1413 (N_1413,In_329,In_1267);
and U1414 (N_1414,In_1068,In_900);
nand U1415 (N_1415,In_1167,In_1436);
nand U1416 (N_1416,In_85,In_1154);
nor U1417 (N_1417,In_47,In_1447);
or U1418 (N_1418,In_177,In_710);
nor U1419 (N_1419,In_590,In_851);
and U1420 (N_1420,In_1022,In_527);
and U1421 (N_1421,In_509,In_66);
and U1422 (N_1422,In_1316,In_1095);
nand U1423 (N_1423,In_1439,In_115);
or U1424 (N_1424,In_1452,In_425);
and U1425 (N_1425,In_713,In_487);
and U1426 (N_1426,In_1162,In_1009);
and U1427 (N_1427,In_1331,In_502);
nor U1428 (N_1428,In_262,In_1272);
nor U1429 (N_1429,In_857,In_650);
nand U1430 (N_1430,In_217,In_124);
nor U1431 (N_1431,In_723,In_970);
or U1432 (N_1432,In_603,In_30);
nand U1433 (N_1433,In_461,In_1104);
and U1434 (N_1434,In_488,In_366);
or U1435 (N_1435,In_1300,In_1404);
or U1436 (N_1436,In_15,In_1127);
nor U1437 (N_1437,In_983,In_86);
nor U1438 (N_1438,In_1470,In_822);
or U1439 (N_1439,In_99,In_102);
nor U1440 (N_1440,In_1266,In_302);
nor U1441 (N_1441,In_1315,In_679);
or U1442 (N_1442,In_231,In_802);
nor U1443 (N_1443,In_767,In_251);
or U1444 (N_1444,In_115,In_10);
nand U1445 (N_1445,In_266,In_290);
and U1446 (N_1446,In_52,In_315);
nor U1447 (N_1447,In_155,In_1233);
nor U1448 (N_1448,In_1088,In_696);
or U1449 (N_1449,In_876,In_4);
nor U1450 (N_1450,In_800,In_827);
and U1451 (N_1451,In_721,In_704);
and U1452 (N_1452,In_1200,In_1437);
or U1453 (N_1453,In_1038,In_544);
and U1454 (N_1454,In_937,In_740);
nor U1455 (N_1455,In_1445,In_1012);
nand U1456 (N_1456,In_217,In_238);
nand U1457 (N_1457,In_873,In_929);
nand U1458 (N_1458,In_1026,In_816);
and U1459 (N_1459,In_990,In_69);
nand U1460 (N_1460,In_479,In_250);
or U1461 (N_1461,In_706,In_668);
xor U1462 (N_1462,In_904,In_1296);
nor U1463 (N_1463,In_380,In_1031);
nor U1464 (N_1464,In_1039,In_1084);
nand U1465 (N_1465,In_1330,In_1100);
nor U1466 (N_1466,In_1279,In_162);
or U1467 (N_1467,In_398,In_193);
and U1468 (N_1468,In_585,In_727);
and U1469 (N_1469,In_549,In_502);
or U1470 (N_1470,In_237,In_1110);
nor U1471 (N_1471,In_454,In_852);
nor U1472 (N_1472,In_321,In_476);
nand U1473 (N_1473,In_777,In_105);
and U1474 (N_1474,In_1271,In_604);
and U1475 (N_1475,In_868,In_1487);
or U1476 (N_1476,In_944,In_624);
nor U1477 (N_1477,In_1232,In_1386);
and U1478 (N_1478,In_94,In_288);
nand U1479 (N_1479,In_338,In_851);
nor U1480 (N_1480,In_1285,In_1102);
or U1481 (N_1481,In_528,In_731);
and U1482 (N_1482,In_1264,In_128);
or U1483 (N_1483,In_888,In_765);
or U1484 (N_1484,In_384,In_1254);
or U1485 (N_1485,In_658,In_331);
nor U1486 (N_1486,In_1169,In_283);
or U1487 (N_1487,In_1237,In_461);
nor U1488 (N_1488,In_1300,In_1195);
xnor U1489 (N_1489,In_293,In_963);
or U1490 (N_1490,In_247,In_1106);
and U1491 (N_1491,In_183,In_1257);
nor U1492 (N_1492,In_750,In_799);
and U1493 (N_1493,In_315,In_1275);
nor U1494 (N_1494,In_778,In_353);
nor U1495 (N_1495,In_816,In_57);
nand U1496 (N_1496,In_559,In_520);
nor U1497 (N_1497,In_467,In_189);
or U1498 (N_1498,In_1338,In_211);
nor U1499 (N_1499,In_1447,In_502);
or U1500 (N_1500,In_542,In_490);
and U1501 (N_1501,In_979,In_456);
or U1502 (N_1502,In_802,In_1268);
nand U1503 (N_1503,In_718,In_603);
nor U1504 (N_1504,In_1305,In_338);
and U1505 (N_1505,In_536,In_935);
or U1506 (N_1506,In_404,In_914);
nand U1507 (N_1507,In_573,In_473);
nor U1508 (N_1508,In_791,In_817);
nor U1509 (N_1509,In_933,In_100);
xnor U1510 (N_1510,In_167,In_504);
nand U1511 (N_1511,In_1224,In_704);
nand U1512 (N_1512,In_1096,In_231);
or U1513 (N_1513,In_811,In_969);
nor U1514 (N_1514,In_740,In_30);
and U1515 (N_1515,In_1318,In_46);
and U1516 (N_1516,In_668,In_1213);
nand U1517 (N_1517,In_313,In_265);
nor U1518 (N_1518,In_557,In_279);
or U1519 (N_1519,In_1154,In_49);
or U1520 (N_1520,In_1188,In_1318);
and U1521 (N_1521,In_523,In_44);
nand U1522 (N_1522,In_128,In_42);
and U1523 (N_1523,In_810,In_646);
nand U1524 (N_1524,In_779,In_591);
and U1525 (N_1525,In_322,In_279);
or U1526 (N_1526,In_710,In_777);
nor U1527 (N_1527,In_1054,In_256);
or U1528 (N_1528,In_980,In_893);
and U1529 (N_1529,In_3,In_348);
or U1530 (N_1530,In_747,In_875);
nor U1531 (N_1531,In_180,In_556);
nor U1532 (N_1532,In_290,In_207);
or U1533 (N_1533,In_845,In_818);
nand U1534 (N_1534,In_1262,In_7);
or U1535 (N_1535,In_529,In_1196);
nor U1536 (N_1536,In_1496,In_68);
and U1537 (N_1537,In_925,In_1378);
and U1538 (N_1538,In_1360,In_1016);
nor U1539 (N_1539,In_855,In_602);
nand U1540 (N_1540,In_1158,In_1361);
nor U1541 (N_1541,In_812,In_211);
and U1542 (N_1542,In_1112,In_427);
xnor U1543 (N_1543,In_588,In_1492);
nand U1544 (N_1544,In_493,In_1171);
nand U1545 (N_1545,In_202,In_169);
nor U1546 (N_1546,In_1455,In_762);
or U1547 (N_1547,In_1146,In_965);
nor U1548 (N_1548,In_367,In_147);
or U1549 (N_1549,In_185,In_548);
nor U1550 (N_1550,In_790,In_873);
nand U1551 (N_1551,In_646,In_499);
or U1552 (N_1552,In_1221,In_1304);
and U1553 (N_1553,In_1099,In_874);
or U1554 (N_1554,In_731,In_753);
and U1555 (N_1555,In_888,In_1243);
and U1556 (N_1556,In_560,In_816);
or U1557 (N_1557,In_465,In_242);
and U1558 (N_1558,In_1174,In_1419);
or U1559 (N_1559,In_90,In_482);
or U1560 (N_1560,In_514,In_777);
nor U1561 (N_1561,In_1334,In_497);
nor U1562 (N_1562,In_1220,In_815);
or U1563 (N_1563,In_520,In_181);
nand U1564 (N_1564,In_712,In_548);
nand U1565 (N_1565,In_47,In_6);
nor U1566 (N_1566,In_121,In_715);
nand U1567 (N_1567,In_595,In_520);
or U1568 (N_1568,In_183,In_532);
nand U1569 (N_1569,In_1482,In_392);
nor U1570 (N_1570,In_679,In_592);
nand U1571 (N_1571,In_1061,In_431);
nor U1572 (N_1572,In_5,In_438);
and U1573 (N_1573,In_149,In_963);
nor U1574 (N_1574,In_1467,In_1003);
nand U1575 (N_1575,In_221,In_52);
and U1576 (N_1576,In_142,In_1272);
nor U1577 (N_1577,In_1152,In_69);
nand U1578 (N_1578,In_645,In_1346);
nor U1579 (N_1579,In_1466,In_305);
nor U1580 (N_1580,In_419,In_1260);
nor U1581 (N_1581,In_640,In_451);
nand U1582 (N_1582,In_584,In_493);
nor U1583 (N_1583,In_162,In_937);
or U1584 (N_1584,In_149,In_219);
and U1585 (N_1585,In_267,In_984);
or U1586 (N_1586,In_1371,In_362);
nand U1587 (N_1587,In_707,In_362);
and U1588 (N_1588,In_820,In_151);
or U1589 (N_1589,In_476,In_958);
nor U1590 (N_1590,In_223,In_246);
xor U1591 (N_1591,In_88,In_1268);
or U1592 (N_1592,In_457,In_947);
nor U1593 (N_1593,In_434,In_1213);
nand U1594 (N_1594,In_919,In_1099);
nand U1595 (N_1595,In_850,In_968);
nor U1596 (N_1596,In_1196,In_1423);
and U1597 (N_1597,In_730,In_733);
nor U1598 (N_1598,In_1138,In_683);
or U1599 (N_1599,In_446,In_1104);
and U1600 (N_1600,In_117,In_173);
nor U1601 (N_1601,In_1439,In_1208);
or U1602 (N_1602,In_658,In_1479);
xnor U1603 (N_1603,In_710,In_1487);
and U1604 (N_1604,In_1204,In_205);
nand U1605 (N_1605,In_47,In_988);
or U1606 (N_1606,In_403,In_140);
or U1607 (N_1607,In_177,In_643);
nor U1608 (N_1608,In_437,In_1325);
nand U1609 (N_1609,In_231,In_667);
nand U1610 (N_1610,In_394,In_606);
and U1611 (N_1611,In_777,In_586);
nand U1612 (N_1612,In_827,In_1463);
nor U1613 (N_1613,In_1137,In_194);
or U1614 (N_1614,In_502,In_1271);
nand U1615 (N_1615,In_994,In_4);
and U1616 (N_1616,In_1080,In_1289);
or U1617 (N_1617,In_158,In_1378);
nand U1618 (N_1618,In_47,In_468);
nor U1619 (N_1619,In_1320,In_866);
nand U1620 (N_1620,In_108,In_465);
nand U1621 (N_1621,In_683,In_1202);
nand U1622 (N_1622,In_120,In_1464);
or U1623 (N_1623,In_217,In_914);
or U1624 (N_1624,In_713,In_1497);
xnor U1625 (N_1625,In_161,In_1017);
or U1626 (N_1626,In_597,In_376);
or U1627 (N_1627,In_860,In_771);
or U1628 (N_1628,In_383,In_36);
nand U1629 (N_1629,In_276,In_55);
nor U1630 (N_1630,In_344,In_857);
or U1631 (N_1631,In_1044,In_551);
nor U1632 (N_1632,In_393,In_1092);
or U1633 (N_1633,In_1273,In_999);
nor U1634 (N_1634,In_1369,In_905);
and U1635 (N_1635,In_1431,In_755);
nor U1636 (N_1636,In_457,In_154);
and U1637 (N_1637,In_1281,In_1311);
nor U1638 (N_1638,In_423,In_355);
nor U1639 (N_1639,In_1010,In_798);
or U1640 (N_1640,In_411,In_95);
or U1641 (N_1641,In_1010,In_1332);
or U1642 (N_1642,In_788,In_1465);
nor U1643 (N_1643,In_971,In_67);
nor U1644 (N_1644,In_778,In_973);
or U1645 (N_1645,In_119,In_1095);
or U1646 (N_1646,In_416,In_838);
nand U1647 (N_1647,In_293,In_1090);
or U1648 (N_1648,In_479,In_962);
nor U1649 (N_1649,In_826,In_386);
and U1650 (N_1650,In_1342,In_685);
nand U1651 (N_1651,In_564,In_488);
nor U1652 (N_1652,In_1477,In_95);
and U1653 (N_1653,In_799,In_775);
nand U1654 (N_1654,In_39,In_1402);
nor U1655 (N_1655,In_738,In_1466);
nand U1656 (N_1656,In_96,In_828);
nor U1657 (N_1657,In_1145,In_586);
and U1658 (N_1658,In_211,In_1100);
and U1659 (N_1659,In_170,In_1437);
and U1660 (N_1660,In_31,In_1166);
and U1661 (N_1661,In_390,In_1373);
and U1662 (N_1662,In_291,In_1143);
or U1663 (N_1663,In_311,In_642);
or U1664 (N_1664,In_521,In_1049);
nand U1665 (N_1665,In_1074,In_763);
nor U1666 (N_1666,In_731,In_390);
nor U1667 (N_1667,In_1408,In_383);
nor U1668 (N_1668,In_1371,In_1477);
nor U1669 (N_1669,In_817,In_1463);
and U1670 (N_1670,In_1007,In_1161);
nand U1671 (N_1671,In_433,In_1251);
nor U1672 (N_1672,In_1033,In_749);
nor U1673 (N_1673,In_1147,In_474);
or U1674 (N_1674,In_752,In_304);
nor U1675 (N_1675,In_589,In_163);
nor U1676 (N_1676,In_1329,In_1097);
nor U1677 (N_1677,In_1291,In_981);
or U1678 (N_1678,In_549,In_1405);
nand U1679 (N_1679,In_628,In_72);
and U1680 (N_1680,In_1399,In_422);
nor U1681 (N_1681,In_266,In_544);
nand U1682 (N_1682,In_263,In_811);
nor U1683 (N_1683,In_558,In_1108);
nand U1684 (N_1684,In_754,In_1204);
nor U1685 (N_1685,In_1176,In_867);
or U1686 (N_1686,In_696,In_785);
nor U1687 (N_1687,In_1015,In_1085);
nand U1688 (N_1688,In_1027,In_169);
or U1689 (N_1689,In_1034,In_1020);
nand U1690 (N_1690,In_682,In_119);
or U1691 (N_1691,In_48,In_111);
or U1692 (N_1692,In_483,In_225);
or U1693 (N_1693,In_40,In_475);
nand U1694 (N_1694,In_1374,In_842);
nor U1695 (N_1695,In_291,In_941);
nor U1696 (N_1696,In_1386,In_29);
or U1697 (N_1697,In_854,In_362);
and U1698 (N_1698,In_354,In_1206);
nand U1699 (N_1699,In_1412,In_90);
or U1700 (N_1700,In_753,In_76);
and U1701 (N_1701,In_328,In_270);
or U1702 (N_1702,In_526,In_1312);
and U1703 (N_1703,In_20,In_123);
or U1704 (N_1704,In_187,In_593);
or U1705 (N_1705,In_1481,In_1360);
nor U1706 (N_1706,In_1321,In_714);
and U1707 (N_1707,In_1113,In_1188);
nor U1708 (N_1708,In_74,In_1443);
or U1709 (N_1709,In_1349,In_561);
nand U1710 (N_1710,In_478,In_981);
nor U1711 (N_1711,In_776,In_1145);
or U1712 (N_1712,In_483,In_1366);
nor U1713 (N_1713,In_900,In_1479);
nand U1714 (N_1714,In_870,In_625);
and U1715 (N_1715,In_434,In_851);
or U1716 (N_1716,In_370,In_275);
nand U1717 (N_1717,In_492,In_1108);
or U1718 (N_1718,In_1005,In_1285);
or U1719 (N_1719,In_375,In_1154);
and U1720 (N_1720,In_243,In_1394);
and U1721 (N_1721,In_142,In_1258);
and U1722 (N_1722,In_439,In_1348);
xnor U1723 (N_1723,In_1086,In_912);
nor U1724 (N_1724,In_301,In_75);
nand U1725 (N_1725,In_955,In_11);
and U1726 (N_1726,In_532,In_1460);
or U1727 (N_1727,In_665,In_51);
nand U1728 (N_1728,In_400,In_728);
or U1729 (N_1729,In_1089,In_29);
nor U1730 (N_1730,In_371,In_128);
nor U1731 (N_1731,In_727,In_406);
nor U1732 (N_1732,In_942,In_1264);
and U1733 (N_1733,In_611,In_644);
or U1734 (N_1734,In_531,In_1053);
nor U1735 (N_1735,In_216,In_115);
or U1736 (N_1736,In_370,In_375);
nor U1737 (N_1737,In_1434,In_962);
nor U1738 (N_1738,In_139,In_233);
nor U1739 (N_1739,In_128,In_63);
nand U1740 (N_1740,In_480,In_743);
nor U1741 (N_1741,In_854,In_55);
and U1742 (N_1742,In_1304,In_892);
nor U1743 (N_1743,In_255,In_1285);
nor U1744 (N_1744,In_1284,In_1349);
or U1745 (N_1745,In_1461,In_706);
or U1746 (N_1746,In_28,In_452);
and U1747 (N_1747,In_154,In_1240);
or U1748 (N_1748,In_1028,In_222);
or U1749 (N_1749,In_144,In_1239);
and U1750 (N_1750,In_231,In_982);
xnor U1751 (N_1751,In_537,In_513);
nand U1752 (N_1752,In_1408,In_1336);
nor U1753 (N_1753,In_335,In_1050);
or U1754 (N_1754,In_1289,In_903);
nand U1755 (N_1755,In_1249,In_427);
nor U1756 (N_1756,In_596,In_1458);
or U1757 (N_1757,In_410,In_539);
nand U1758 (N_1758,In_847,In_789);
and U1759 (N_1759,In_711,In_642);
and U1760 (N_1760,In_861,In_447);
and U1761 (N_1761,In_940,In_643);
nand U1762 (N_1762,In_1198,In_1482);
or U1763 (N_1763,In_1417,In_1201);
and U1764 (N_1764,In_809,In_266);
or U1765 (N_1765,In_957,In_912);
and U1766 (N_1766,In_330,In_1205);
or U1767 (N_1767,In_959,In_1338);
and U1768 (N_1768,In_257,In_94);
nand U1769 (N_1769,In_64,In_53);
nor U1770 (N_1770,In_813,In_1333);
nor U1771 (N_1771,In_947,In_1495);
and U1772 (N_1772,In_498,In_132);
nor U1773 (N_1773,In_208,In_626);
nor U1774 (N_1774,In_262,In_199);
nand U1775 (N_1775,In_799,In_616);
and U1776 (N_1776,In_1001,In_606);
and U1777 (N_1777,In_1292,In_1394);
or U1778 (N_1778,In_792,In_850);
and U1779 (N_1779,In_1003,In_365);
or U1780 (N_1780,In_403,In_273);
nor U1781 (N_1781,In_850,In_702);
and U1782 (N_1782,In_465,In_1331);
nor U1783 (N_1783,In_515,In_1032);
nand U1784 (N_1784,In_936,In_871);
or U1785 (N_1785,In_1353,In_476);
and U1786 (N_1786,In_574,In_1441);
or U1787 (N_1787,In_264,In_917);
nor U1788 (N_1788,In_1309,In_730);
and U1789 (N_1789,In_1481,In_761);
and U1790 (N_1790,In_225,In_1320);
nand U1791 (N_1791,In_1253,In_645);
and U1792 (N_1792,In_1156,In_1197);
or U1793 (N_1793,In_424,In_1267);
or U1794 (N_1794,In_525,In_222);
and U1795 (N_1795,In_1202,In_32);
nand U1796 (N_1796,In_660,In_651);
or U1797 (N_1797,In_30,In_64);
and U1798 (N_1798,In_543,In_873);
and U1799 (N_1799,In_968,In_1480);
nand U1800 (N_1800,In_1160,In_850);
or U1801 (N_1801,In_407,In_195);
nand U1802 (N_1802,In_1255,In_726);
nand U1803 (N_1803,In_581,In_686);
nor U1804 (N_1804,In_794,In_617);
or U1805 (N_1805,In_322,In_303);
nor U1806 (N_1806,In_1002,In_1385);
and U1807 (N_1807,In_460,In_1193);
nor U1808 (N_1808,In_727,In_1139);
or U1809 (N_1809,In_69,In_1073);
nand U1810 (N_1810,In_728,In_1237);
nor U1811 (N_1811,In_1140,In_1039);
and U1812 (N_1812,In_187,In_289);
or U1813 (N_1813,In_405,In_333);
nand U1814 (N_1814,In_531,In_748);
and U1815 (N_1815,In_570,In_1409);
nor U1816 (N_1816,In_1137,In_1471);
nor U1817 (N_1817,In_93,In_1190);
or U1818 (N_1818,In_823,In_1434);
nand U1819 (N_1819,In_464,In_166);
or U1820 (N_1820,In_1031,In_365);
nor U1821 (N_1821,In_670,In_1286);
or U1822 (N_1822,In_23,In_179);
and U1823 (N_1823,In_1052,In_1312);
or U1824 (N_1824,In_418,In_61);
nor U1825 (N_1825,In_870,In_860);
nor U1826 (N_1826,In_525,In_472);
and U1827 (N_1827,In_421,In_1132);
and U1828 (N_1828,In_193,In_1482);
nor U1829 (N_1829,In_151,In_37);
xor U1830 (N_1830,In_766,In_997);
and U1831 (N_1831,In_778,In_1359);
nor U1832 (N_1832,In_634,In_108);
nand U1833 (N_1833,In_1409,In_190);
nor U1834 (N_1834,In_146,In_1257);
nor U1835 (N_1835,In_717,In_713);
and U1836 (N_1836,In_659,In_976);
or U1837 (N_1837,In_1321,In_537);
or U1838 (N_1838,In_831,In_189);
and U1839 (N_1839,In_228,In_1469);
or U1840 (N_1840,In_1305,In_109);
nor U1841 (N_1841,In_834,In_1254);
and U1842 (N_1842,In_25,In_382);
nand U1843 (N_1843,In_395,In_774);
nor U1844 (N_1844,In_1050,In_343);
nand U1845 (N_1845,In_795,In_1015);
nor U1846 (N_1846,In_967,In_1211);
nand U1847 (N_1847,In_218,In_388);
and U1848 (N_1848,In_107,In_872);
or U1849 (N_1849,In_1453,In_574);
nor U1850 (N_1850,In_866,In_998);
and U1851 (N_1851,In_1377,In_271);
or U1852 (N_1852,In_771,In_1332);
or U1853 (N_1853,In_1399,In_1283);
nand U1854 (N_1854,In_253,In_197);
nand U1855 (N_1855,In_931,In_814);
nor U1856 (N_1856,In_521,In_1399);
nand U1857 (N_1857,In_344,In_1382);
nand U1858 (N_1858,In_1065,In_1490);
or U1859 (N_1859,In_927,In_262);
nor U1860 (N_1860,In_1394,In_1449);
nor U1861 (N_1861,In_981,In_94);
and U1862 (N_1862,In_463,In_737);
nor U1863 (N_1863,In_571,In_952);
and U1864 (N_1864,In_1230,In_102);
or U1865 (N_1865,In_1393,In_602);
or U1866 (N_1866,In_1166,In_424);
nand U1867 (N_1867,In_891,In_510);
nor U1868 (N_1868,In_803,In_617);
nor U1869 (N_1869,In_535,In_607);
nand U1870 (N_1870,In_42,In_136);
and U1871 (N_1871,In_434,In_137);
or U1872 (N_1872,In_1029,In_277);
nand U1873 (N_1873,In_916,In_479);
and U1874 (N_1874,In_900,In_909);
nor U1875 (N_1875,In_1412,In_180);
nand U1876 (N_1876,In_701,In_1433);
nand U1877 (N_1877,In_656,In_1391);
nor U1878 (N_1878,In_916,In_1430);
nand U1879 (N_1879,In_1348,In_1182);
and U1880 (N_1880,In_335,In_1240);
nand U1881 (N_1881,In_1305,In_274);
and U1882 (N_1882,In_683,In_302);
xor U1883 (N_1883,In_1458,In_759);
nand U1884 (N_1884,In_57,In_172);
nand U1885 (N_1885,In_742,In_901);
or U1886 (N_1886,In_538,In_343);
or U1887 (N_1887,In_720,In_1365);
and U1888 (N_1888,In_1445,In_1246);
or U1889 (N_1889,In_1219,In_1340);
and U1890 (N_1890,In_158,In_11);
nand U1891 (N_1891,In_1182,In_694);
nor U1892 (N_1892,In_235,In_394);
or U1893 (N_1893,In_1256,In_291);
or U1894 (N_1894,In_950,In_680);
or U1895 (N_1895,In_229,In_176);
nand U1896 (N_1896,In_1002,In_1181);
and U1897 (N_1897,In_1298,In_148);
xnor U1898 (N_1898,In_1096,In_1046);
nor U1899 (N_1899,In_190,In_694);
nand U1900 (N_1900,In_932,In_781);
and U1901 (N_1901,In_568,In_1345);
and U1902 (N_1902,In_1357,In_353);
or U1903 (N_1903,In_46,In_531);
or U1904 (N_1904,In_845,In_1160);
and U1905 (N_1905,In_1113,In_596);
nand U1906 (N_1906,In_545,In_1349);
and U1907 (N_1907,In_1425,In_1307);
or U1908 (N_1908,In_248,In_1374);
and U1909 (N_1909,In_1228,In_110);
nor U1910 (N_1910,In_119,In_1152);
xor U1911 (N_1911,In_746,In_442);
nor U1912 (N_1912,In_251,In_132);
or U1913 (N_1913,In_1374,In_189);
and U1914 (N_1914,In_1233,In_850);
or U1915 (N_1915,In_616,In_1377);
or U1916 (N_1916,In_1028,In_854);
nand U1917 (N_1917,In_1324,In_599);
xnor U1918 (N_1918,In_1039,In_385);
nor U1919 (N_1919,In_53,In_1276);
nor U1920 (N_1920,In_1457,In_168);
xor U1921 (N_1921,In_1188,In_887);
nand U1922 (N_1922,In_899,In_431);
nand U1923 (N_1923,In_14,In_483);
nor U1924 (N_1924,In_1172,In_962);
xor U1925 (N_1925,In_710,In_143);
nand U1926 (N_1926,In_428,In_1274);
or U1927 (N_1927,In_840,In_906);
or U1928 (N_1928,In_749,In_680);
nand U1929 (N_1929,In_346,In_582);
nand U1930 (N_1930,In_865,In_291);
and U1931 (N_1931,In_1345,In_1225);
and U1932 (N_1932,In_564,In_231);
or U1933 (N_1933,In_951,In_1110);
and U1934 (N_1934,In_731,In_670);
nand U1935 (N_1935,In_45,In_352);
or U1936 (N_1936,In_899,In_1153);
nand U1937 (N_1937,In_1181,In_262);
or U1938 (N_1938,In_1498,In_1086);
or U1939 (N_1939,In_681,In_196);
nand U1940 (N_1940,In_764,In_930);
and U1941 (N_1941,In_677,In_79);
and U1942 (N_1942,In_476,In_1017);
or U1943 (N_1943,In_795,In_631);
or U1944 (N_1944,In_656,In_755);
nand U1945 (N_1945,In_1201,In_620);
and U1946 (N_1946,In_665,In_697);
and U1947 (N_1947,In_1388,In_791);
or U1948 (N_1948,In_603,In_1457);
nor U1949 (N_1949,In_718,In_1174);
or U1950 (N_1950,In_433,In_509);
or U1951 (N_1951,In_673,In_258);
or U1952 (N_1952,In_758,In_372);
nand U1953 (N_1953,In_35,In_1110);
and U1954 (N_1954,In_411,In_1272);
nor U1955 (N_1955,In_555,In_736);
and U1956 (N_1956,In_1387,In_211);
nor U1957 (N_1957,In_262,In_1217);
or U1958 (N_1958,In_939,In_231);
nand U1959 (N_1959,In_328,In_1395);
and U1960 (N_1960,In_922,In_1359);
nor U1961 (N_1961,In_352,In_1306);
or U1962 (N_1962,In_210,In_463);
and U1963 (N_1963,In_417,In_279);
nand U1964 (N_1964,In_106,In_644);
nand U1965 (N_1965,In_806,In_1387);
nand U1966 (N_1966,In_172,In_1336);
nor U1967 (N_1967,In_298,In_593);
xor U1968 (N_1968,In_1423,In_74);
nor U1969 (N_1969,In_1057,In_627);
nor U1970 (N_1970,In_1237,In_339);
or U1971 (N_1971,In_51,In_1243);
nor U1972 (N_1972,In_1474,In_716);
nand U1973 (N_1973,In_85,In_1102);
and U1974 (N_1974,In_515,In_86);
or U1975 (N_1975,In_296,In_754);
or U1976 (N_1976,In_1311,In_290);
and U1977 (N_1977,In_724,In_321);
or U1978 (N_1978,In_696,In_899);
nand U1979 (N_1979,In_902,In_1019);
nand U1980 (N_1980,In_278,In_450);
nand U1981 (N_1981,In_985,In_1330);
nand U1982 (N_1982,In_1389,In_582);
and U1983 (N_1983,In_1469,In_1204);
xor U1984 (N_1984,In_903,In_952);
nor U1985 (N_1985,In_780,In_478);
nand U1986 (N_1986,In_529,In_704);
and U1987 (N_1987,In_1250,In_566);
nand U1988 (N_1988,In_270,In_1031);
nand U1989 (N_1989,In_1433,In_976);
and U1990 (N_1990,In_16,In_1132);
or U1991 (N_1991,In_842,In_805);
and U1992 (N_1992,In_756,In_1045);
nand U1993 (N_1993,In_194,In_294);
and U1994 (N_1994,In_868,In_141);
nor U1995 (N_1995,In_1421,In_1213);
nand U1996 (N_1996,In_251,In_827);
and U1997 (N_1997,In_166,In_596);
and U1998 (N_1998,In_483,In_209);
and U1999 (N_1999,In_221,In_674);
nand U2000 (N_2000,In_1467,In_867);
or U2001 (N_2001,In_338,In_1389);
nand U2002 (N_2002,In_1228,In_769);
nand U2003 (N_2003,In_1175,In_764);
xnor U2004 (N_2004,In_410,In_1366);
nor U2005 (N_2005,In_394,In_1137);
nor U2006 (N_2006,In_120,In_784);
xor U2007 (N_2007,In_1237,In_357);
nand U2008 (N_2008,In_1056,In_108);
and U2009 (N_2009,In_558,In_1397);
or U2010 (N_2010,In_302,In_1481);
nand U2011 (N_2011,In_438,In_421);
or U2012 (N_2012,In_1210,In_1378);
or U2013 (N_2013,In_739,In_645);
and U2014 (N_2014,In_816,In_242);
or U2015 (N_2015,In_481,In_766);
nand U2016 (N_2016,In_1139,In_810);
nor U2017 (N_2017,In_336,In_1005);
xor U2018 (N_2018,In_1023,In_670);
nor U2019 (N_2019,In_581,In_620);
or U2020 (N_2020,In_928,In_1052);
and U2021 (N_2021,In_220,In_1423);
and U2022 (N_2022,In_200,In_1124);
nor U2023 (N_2023,In_580,In_167);
nor U2024 (N_2024,In_364,In_730);
nand U2025 (N_2025,In_671,In_413);
and U2026 (N_2026,In_1494,In_75);
nor U2027 (N_2027,In_142,In_430);
or U2028 (N_2028,In_251,In_435);
or U2029 (N_2029,In_1425,In_1151);
or U2030 (N_2030,In_1383,In_696);
nand U2031 (N_2031,In_67,In_907);
and U2032 (N_2032,In_1112,In_1359);
or U2033 (N_2033,In_292,In_371);
and U2034 (N_2034,In_690,In_871);
or U2035 (N_2035,In_335,In_1424);
nor U2036 (N_2036,In_1459,In_37);
and U2037 (N_2037,In_802,In_1341);
or U2038 (N_2038,In_707,In_1160);
and U2039 (N_2039,In_1253,In_1385);
nor U2040 (N_2040,In_962,In_1183);
and U2041 (N_2041,In_360,In_802);
and U2042 (N_2042,In_728,In_578);
or U2043 (N_2043,In_1258,In_1166);
nand U2044 (N_2044,In_245,In_164);
nand U2045 (N_2045,In_132,In_1274);
and U2046 (N_2046,In_906,In_1496);
nor U2047 (N_2047,In_1434,In_672);
xnor U2048 (N_2048,In_924,In_1139);
nand U2049 (N_2049,In_492,In_785);
nor U2050 (N_2050,In_105,In_382);
or U2051 (N_2051,In_43,In_702);
or U2052 (N_2052,In_748,In_637);
nand U2053 (N_2053,In_1066,In_375);
or U2054 (N_2054,In_698,In_436);
nor U2055 (N_2055,In_191,In_1051);
nand U2056 (N_2056,In_938,In_1062);
xnor U2057 (N_2057,In_415,In_414);
nand U2058 (N_2058,In_148,In_793);
and U2059 (N_2059,In_840,In_273);
nand U2060 (N_2060,In_431,In_1074);
and U2061 (N_2061,In_886,In_749);
or U2062 (N_2062,In_1243,In_405);
or U2063 (N_2063,In_926,In_200);
nand U2064 (N_2064,In_927,In_20);
or U2065 (N_2065,In_33,In_962);
or U2066 (N_2066,In_221,In_1092);
or U2067 (N_2067,In_1418,In_402);
or U2068 (N_2068,In_240,In_1263);
nor U2069 (N_2069,In_414,In_302);
nand U2070 (N_2070,In_706,In_812);
nand U2071 (N_2071,In_923,In_128);
nor U2072 (N_2072,In_54,In_1454);
and U2073 (N_2073,In_882,In_304);
nand U2074 (N_2074,In_1444,In_570);
nor U2075 (N_2075,In_1422,In_1063);
or U2076 (N_2076,In_1385,In_1335);
nor U2077 (N_2077,In_1238,In_840);
or U2078 (N_2078,In_1228,In_91);
and U2079 (N_2079,In_687,In_90);
and U2080 (N_2080,In_980,In_1475);
nor U2081 (N_2081,In_153,In_1300);
or U2082 (N_2082,In_1327,In_1173);
nand U2083 (N_2083,In_152,In_207);
or U2084 (N_2084,In_1463,In_186);
nor U2085 (N_2085,In_777,In_1102);
and U2086 (N_2086,In_976,In_1241);
or U2087 (N_2087,In_755,In_576);
and U2088 (N_2088,In_1101,In_785);
nand U2089 (N_2089,In_724,In_1029);
nand U2090 (N_2090,In_920,In_396);
or U2091 (N_2091,In_391,In_73);
or U2092 (N_2092,In_555,In_1035);
nand U2093 (N_2093,In_1389,In_622);
or U2094 (N_2094,In_455,In_936);
nor U2095 (N_2095,In_80,In_605);
and U2096 (N_2096,In_887,In_498);
nor U2097 (N_2097,In_893,In_466);
nand U2098 (N_2098,In_368,In_1186);
nand U2099 (N_2099,In_449,In_206);
nand U2100 (N_2100,In_794,In_1382);
and U2101 (N_2101,In_681,In_985);
and U2102 (N_2102,In_1153,In_1157);
nor U2103 (N_2103,In_1416,In_544);
and U2104 (N_2104,In_935,In_788);
nor U2105 (N_2105,In_781,In_773);
xor U2106 (N_2106,In_315,In_205);
or U2107 (N_2107,In_1294,In_1239);
nand U2108 (N_2108,In_517,In_357);
or U2109 (N_2109,In_1413,In_260);
and U2110 (N_2110,In_619,In_1002);
or U2111 (N_2111,In_1065,In_453);
xor U2112 (N_2112,In_174,In_1497);
nand U2113 (N_2113,In_1035,In_1213);
or U2114 (N_2114,In_998,In_231);
nor U2115 (N_2115,In_1459,In_1483);
nor U2116 (N_2116,In_3,In_215);
nor U2117 (N_2117,In_1392,In_988);
nor U2118 (N_2118,In_344,In_683);
nand U2119 (N_2119,In_986,In_88);
xor U2120 (N_2120,In_211,In_497);
or U2121 (N_2121,In_638,In_960);
or U2122 (N_2122,In_595,In_928);
or U2123 (N_2123,In_872,In_1120);
nor U2124 (N_2124,In_462,In_1217);
and U2125 (N_2125,In_1376,In_91);
or U2126 (N_2126,In_858,In_1386);
or U2127 (N_2127,In_1257,In_103);
or U2128 (N_2128,In_1283,In_1024);
nand U2129 (N_2129,In_1134,In_1274);
and U2130 (N_2130,In_1445,In_98);
xor U2131 (N_2131,In_413,In_1246);
or U2132 (N_2132,In_164,In_784);
and U2133 (N_2133,In_28,In_518);
and U2134 (N_2134,In_731,In_825);
or U2135 (N_2135,In_1075,In_1148);
nand U2136 (N_2136,In_1369,In_1300);
and U2137 (N_2137,In_301,In_564);
nor U2138 (N_2138,In_453,In_121);
and U2139 (N_2139,In_929,In_616);
or U2140 (N_2140,In_978,In_778);
and U2141 (N_2141,In_1379,In_406);
xnor U2142 (N_2142,In_458,In_76);
or U2143 (N_2143,In_320,In_675);
nor U2144 (N_2144,In_872,In_858);
nor U2145 (N_2145,In_812,In_693);
and U2146 (N_2146,In_448,In_52);
nor U2147 (N_2147,In_610,In_778);
nand U2148 (N_2148,In_996,In_729);
nor U2149 (N_2149,In_506,In_399);
or U2150 (N_2150,In_749,In_698);
and U2151 (N_2151,In_106,In_1214);
or U2152 (N_2152,In_348,In_1260);
and U2153 (N_2153,In_1218,In_231);
or U2154 (N_2154,In_494,In_625);
xor U2155 (N_2155,In_878,In_399);
and U2156 (N_2156,In_967,In_1459);
nand U2157 (N_2157,In_968,In_404);
nor U2158 (N_2158,In_979,In_1283);
and U2159 (N_2159,In_246,In_1436);
nand U2160 (N_2160,In_68,In_661);
or U2161 (N_2161,In_580,In_727);
nand U2162 (N_2162,In_327,In_870);
or U2163 (N_2163,In_786,In_940);
nor U2164 (N_2164,In_22,In_707);
nor U2165 (N_2165,In_722,In_725);
and U2166 (N_2166,In_97,In_812);
and U2167 (N_2167,In_888,In_242);
nor U2168 (N_2168,In_1300,In_98);
and U2169 (N_2169,In_663,In_957);
nand U2170 (N_2170,In_441,In_548);
nand U2171 (N_2171,In_929,In_1264);
nand U2172 (N_2172,In_357,In_265);
nor U2173 (N_2173,In_1073,In_1427);
nand U2174 (N_2174,In_1285,In_1193);
and U2175 (N_2175,In_409,In_601);
nor U2176 (N_2176,In_49,In_1278);
nand U2177 (N_2177,In_998,In_818);
and U2178 (N_2178,In_694,In_347);
or U2179 (N_2179,In_1417,In_154);
nand U2180 (N_2180,In_290,In_709);
nor U2181 (N_2181,In_939,In_120);
or U2182 (N_2182,In_560,In_1272);
or U2183 (N_2183,In_190,In_1273);
or U2184 (N_2184,In_743,In_186);
nand U2185 (N_2185,In_748,In_27);
nand U2186 (N_2186,In_1109,In_1122);
and U2187 (N_2187,In_374,In_38);
or U2188 (N_2188,In_242,In_1120);
and U2189 (N_2189,In_1028,In_862);
nand U2190 (N_2190,In_867,In_1390);
nor U2191 (N_2191,In_883,In_386);
or U2192 (N_2192,In_514,In_477);
nand U2193 (N_2193,In_378,In_682);
nor U2194 (N_2194,In_157,In_1023);
nor U2195 (N_2195,In_811,In_837);
and U2196 (N_2196,In_1201,In_739);
or U2197 (N_2197,In_603,In_992);
and U2198 (N_2198,In_1073,In_334);
nor U2199 (N_2199,In_1263,In_355);
or U2200 (N_2200,In_604,In_183);
or U2201 (N_2201,In_957,In_637);
nor U2202 (N_2202,In_345,In_1057);
nand U2203 (N_2203,In_669,In_931);
or U2204 (N_2204,In_412,In_436);
and U2205 (N_2205,In_702,In_123);
nor U2206 (N_2206,In_1301,In_21);
or U2207 (N_2207,In_15,In_1482);
or U2208 (N_2208,In_972,In_51);
and U2209 (N_2209,In_1283,In_531);
or U2210 (N_2210,In_1133,In_777);
nor U2211 (N_2211,In_336,In_1244);
nor U2212 (N_2212,In_1454,In_191);
nand U2213 (N_2213,In_620,In_606);
nor U2214 (N_2214,In_126,In_54);
nand U2215 (N_2215,In_1030,In_926);
and U2216 (N_2216,In_593,In_1014);
and U2217 (N_2217,In_266,In_1074);
or U2218 (N_2218,In_1308,In_541);
and U2219 (N_2219,In_1176,In_466);
and U2220 (N_2220,In_373,In_1430);
nor U2221 (N_2221,In_705,In_856);
nand U2222 (N_2222,In_793,In_49);
nand U2223 (N_2223,In_457,In_391);
nor U2224 (N_2224,In_1463,In_1442);
or U2225 (N_2225,In_486,In_1295);
and U2226 (N_2226,In_917,In_1320);
nor U2227 (N_2227,In_1017,In_904);
and U2228 (N_2228,In_1041,In_262);
nand U2229 (N_2229,In_788,In_1072);
and U2230 (N_2230,In_1016,In_823);
nand U2231 (N_2231,In_967,In_94);
or U2232 (N_2232,In_493,In_1223);
nor U2233 (N_2233,In_1263,In_929);
and U2234 (N_2234,In_913,In_251);
and U2235 (N_2235,In_574,In_1315);
xnor U2236 (N_2236,In_33,In_1118);
and U2237 (N_2237,In_819,In_814);
nor U2238 (N_2238,In_455,In_1433);
and U2239 (N_2239,In_522,In_631);
and U2240 (N_2240,In_310,In_47);
nor U2241 (N_2241,In_933,In_730);
nand U2242 (N_2242,In_1395,In_1232);
xnor U2243 (N_2243,In_306,In_1125);
nor U2244 (N_2244,In_5,In_111);
nor U2245 (N_2245,In_131,In_1117);
and U2246 (N_2246,In_263,In_316);
and U2247 (N_2247,In_594,In_1426);
and U2248 (N_2248,In_1252,In_364);
or U2249 (N_2249,In_803,In_729);
nor U2250 (N_2250,In_29,In_1298);
nor U2251 (N_2251,In_589,In_823);
or U2252 (N_2252,In_275,In_1309);
and U2253 (N_2253,In_878,In_1300);
nand U2254 (N_2254,In_1386,In_1055);
or U2255 (N_2255,In_4,In_1146);
or U2256 (N_2256,In_219,In_1036);
nor U2257 (N_2257,In_945,In_517);
and U2258 (N_2258,In_339,In_590);
nor U2259 (N_2259,In_1147,In_176);
and U2260 (N_2260,In_1016,In_44);
nand U2261 (N_2261,In_1181,In_231);
nor U2262 (N_2262,In_1080,In_753);
nand U2263 (N_2263,In_435,In_1187);
and U2264 (N_2264,In_550,In_727);
xnor U2265 (N_2265,In_1294,In_1029);
nand U2266 (N_2266,In_1216,In_5);
and U2267 (N_2267,In_142,In_235);
or U2268 (N_2268,In_853,In_131);
nand U2269 (N_2269,In_1330,In_1017);
nand U2270 (N_2270,In_953,In_1496);
and U2271 (N_2271,In_1047,In_1270);
nand U2272 (N_2272,In_209,In_1131);
nand U2273 (N_2273,In_893,In_383);
or U2274 (N_2274,In_1245,In_802);
nand U2275 (N_2275,In_928,In_1348);
and U2276 (N_2276,In_1481,In_1028);
nor U2277 (N_2277,In_521,In_1231);
and U2278 (N_2278,In_121,In_734);
nand U2279 (N_2279,In_118,In_731);
or U2280 (N_2280,In_686,In_1325);
and U2281 (N_2281,In_439,In_1283);
nor U2282 (N_2282,In_173,In_1343);
xor U2283 (N_2283,In_653,In_132);
or U2284 (N_2284,In_194,In_803);
nor U2285 (N_2285,In_785,In_1118);
nor U2286 (N_2286,In_1290,In_601);
and U2287 (N_2287,In_13,In_453);
nor U2288 (N_2288,In_1006,In_591);
or U2289 (N_2289,In_1053,In_862);
or U2290 (N_2290,In_171,In_667);
and U2291 (N_2291,In_1022,In_1275);
nor U2292 (N_2292,In_1093,In_336);
nand U2293 (N_2293,In_789,In_1279);
nand U2294 (N_2294,In_879,In_240);
or U2295 (N_2295,In_1084,In_1051);
nor U2296 (N_2296,In_1372,In_31);
or U2297 (N_2297,In_543,In_1058);
or U2298 (N_2298,In_3,In_506);
nand U2299 (N_2299,In_393,In_940);
and U2300 (N_2300,In_742,In_1327);
nand U2301 (N_2301,In_715,In_1479);
nand U2302 (N_2302,In_1378,In_1277);
nand U2303 (N_2303,In_958,In_248);
or U2304 (N_2304,In_480,In_221);
nand U2305 (N_2305,In_1204,In_501);
nand U2306 (N_2306,In_578,In_288);
and U2307 (N_2307,In_721,In_390);
and U2308 (N_2308,In_700,In_807);
or U2309 (N_2309,In_795,In_1269);
or U2310 (N_2310,In_760,In_1092);
and U2311 (N_2311,In_479,In_279);
nand U2312 (N_2312,In_1164,In_273);
nor U2313 (N_2313,In_380,In_499);
and U2314 (N_2314,In_77,In_304);
xor U2315 (N_2315,In_1267,In_441);
or U2316 (N_2316,In_534,In_49);
xnor U2317 (N_2317,In_1112,In_1117);
nand U2318 (N_2318,In_1145,In_739);
nor U2319 (N_2319,In_240,In_886);
or U2320 (N_2320,In_1218,In_322);
xnor U2321 (N_2321,In_1186,In_311);
xnor U2322 (N_2322,In_1094,In_104);
nor U2323 (N_2323,In_321,In_109);
nand U2324 (N_2324,In_613,In_803);
and U2325 (N_2325,In_672,In_330);
nand U2326 (N_2326,In_80,In_37);
nor U2327 (N_2327,In_1010,In_1458);
nand U2328 (N_2328,In_734,In_1153);
nand U2329 (N_2329,In_821,In_283);
nand U2330 (N_2330,In_1230,In_497);
and U2331 (N_2331,In_109,In_277);
nor U2332 (N_2332,In_1489,In_1075);
nor U2333 (N_2333,In_915,In_1466);
or U2334 (N_2334,In_547,In_744);
or U2335 (N_2335,In_1166,In_1370);
or U2336 (N_2336,In_1019,In_819);
nand U2337 (N_2337,In_646,In_1448);
or U2338 (N_2338,In_893,In_755);
nand U2339 (N_2339,In_745,In_1130);
nor U2340 (N_2340,In_931,In_893);
nor U2341 (N_2341,In_117,In_367);
and U2342 (N_2342,In_900,In_1321);
or U2343 (N_2343,In_1381,In_255);
and U2344 (N_2344,In_629,In_863);
nor U2345 (N_2345,In_129,In_1079);
xnor U2346 (N_2346,In_1194,In_827);
nor U2347 (N_2347,In_1172,In_71);
nor U2348 (N_2348,In_26,In_280);
or U2349 (N_2349,In_1046,In_212);
xor U2350 (N_2350,In_292,In_699);
nand U2351 (N_2351,In_1327,In_609);
nand U2352 (N_2352,In_108,In_1485);
nor U2353 (N_2353,In_1076,In_418);
nor U2354 (N_2354,In_1133,In_210);
and U2355 (N_2355,In_785,In_1468);
nand U2356 (N_2356,In_904,In_811);
xor U2357 (N_2357,In_105,In_45);
or U2358 (N_2358,In_74,In_729);
and U2359 (N_2359,In_635,In_279);
and U2360 (N_2360,In_1216,In_488);
nor U2361 (N_2361,In_17,In_154);
nor U2362 (N_2362,In_319,In_655);
nor U2363 (N_2363,In_713,In_125);
nor U2364 (N_2364,In_1217,In_483);
and U2365 (N_2365,In_187,In_423);
or U2366 (N_2366,In_954,In_1108);
nor U2367 (N_2367,In_967,In_1017);
nand U2368 (N_2368,In_166,In_1069);
and U2369 (N_2369,In_358,In_1240);
or U2370 (N_2370,In_620,In_670);
and U2371 (N_2371,In_726,In_359);
nor U2372 (N_2372,In_1087,In_1146);
and U2373 (N_2373,In_258,In_1010);
and U2374 (N_2374,In_366,In_961);
or U2375 (N_2375,In_1404,In_1220);
nand U2376 (N_2376,In_1083,In_1257);
and U2377 (N_2377,In_1341,In_431);
nand U2378 (N_2378,In_517,In_1440);
nand U2379 (N_2379,In_1226,In_425);
nor U2380 (N_2380,In_967,In_282);
and U2381 (N_2381,In_46,In_814);
nand U2382 (N_2382,In_1181,In_299);
and U2383 (N_2383,In_1241,In_1399);
nand U2384 (N_2384,In_665,In_1394);
nor U2385 (N_2385,In_408,In_901);
and U2386 (N_2386,In_966,In_4);
nand U2387 (N_2387,In_1016,In_718);
nor U2388 (N_2388,In_1248,In_165);
nor U2389 (N_2389,In_278,In_1375);
and U2390 (N_2390,In_449,In_968);
or U2391 (N_2391,In_862,In_1006);
and U2392 (N_2392,In_665,In_498);
nand U2393 (N_2393,In_1384,In_941);
nand U2394 (N_2394,In_248,In_998);
or U2395 (N_2395,In_1403,In_1055);
or U2396 (N_2396,In_217,In_392);
and U2397 (N_2397,In_518,In_271);
nand U2398 (N_2398,In_1250,In_220);
nand U2399 (N_2399,In_444,In_432);
nand U2400 (N_2400,In_894,In_1479);
and U2401 (N_2401,In_1199,In_506);
nor U2402 (N_2402,In_913,In_529);
nor U2403 (N_2403,In_954,In_1307);
or U2404 (N_2404,In_703,In_249);
and U2405 (N_2405,In_1268,In_393);
or U2406 (N_2406,In_942,In_743);
nor U2407 (N_2407,In_19,In_595);
and U2408 (N_2408,In_557,In_551);
and U2409 (N_2409,In_1228,In_797);
nand U2410 (N_2410,In_413,In_680);
and U2411 (N_2411,In_153,In_989);
or U2412 (N_2412,In_370,In_742);
or U2413 (N_2413,In_1037,In_184);
and U2414 (N_2414,In_1225,In_770);
or U2415 (N_2415,In_876,In_1443);
and U2416 (N_2416,In_106,In_874);
nand U2417 (N_2417,In_980,In_1110);
nor U2418 (N_2418,In_1467,In_486);
nand U2419 (N_2419,In_1269,In_1485);
and U2420 (N_2420,In_92,In_517);
nand U2421 (N_2421,In_270,In_659);
nand U2422 (N_2422,In_84,In_897);
nor U2423 (N_2423,In_135,In_762);
and U2424 (N_2424,In_443,In_236);
or U2425 (N_2425,In_47,In_843);
nand U2426 (N_2426,In_1056,In_363);
xnor U2427 (N_2427,In_518,In_1022);
and U2428 (N_2428,In_71,In_1247);
nand U2429 (N_2429,In_944,In_1023);
or U2430 (N_2430,In_959,In_1371);
or U2431 (N_2431,In_855,In_595);
and U2432 (N_2432,In_98,In_1333);
and U2433 (N_2433,In_1221,In_452);
or U2434 (N_2434,In_511,In_794);
nor U2435 (N_2435,In_326,In_1082);
nand U2436 (N_2436,In_222,In_911);
nand U2437 (N_2437,In_919,In_1102);
or U2438 (N_2438,In_1378,In_508);
nor U2439 (N_2439,In_1364,In_354);
nor U2440 (N_2440,In_1010,In_666);
or U2441 (N_2441,In_1413,In_1492);
or U2442 (N_2442,In_1499,In_944);
nor U2443 (N_2443,In_347,In_355);
and U2444 (N_2444,In_332,In_1351);
or U2445 (N_2445,In_853,In_555);
or U2446 (N_2446,In_1407,In_1083);
or U2447 (N_2447,In_157,In_574);
and U2448 (N_2448,In_83,In_1021);
nor U2449 (N_2449,In_619,In_181);
nand U2450 (N_2450,In_392,In_1341);
and U2451 (N_2451,In_1386,In_322);
nand U2452 (N_2452,In_1116,In_872);
nand U2453 (N_2453,In_843,In_753);
and U2454 (N_2454,In_370,In_1134);
nor U2455 (N_2455,In_80,In_1276);
or U2456 (N_2456,In_1281,In_441);
nand U2457 (N_2457,In_124,In_1145);
nor U2458 (N_2458,In_927,In_1110);
or U2459 (N_2459,In_238,In_795);
nor U2460 (N_2460,In_1426,In_697);
or U2461 (N_2461,In_1105,In_1172);
nor U2462 (N_2462,In_823,In_567);
nor U2463 (N_2463,In_1300,In_673);
and U2464 (N_2464,In_159,In_148);
nand U2465 (N_2465,In_1048,In_1300);
and U2466 (N_2466,In_1141,In_857);
or U2467 (N_2467,In_1181,In_1404);
and U2468 (N_2468,In_1176,In_933);
or U2469 (N_2469,In_387,In_689);
nand U2470 (N_2470,In_191,In_33);
xnor U2471 (N_2471,In_1200,In_1128);
nor U2472 (N_2472,In_382,In_1469);
nand U2473 (N_2473,In_710,In_985);
nand U2474 (N_2474,In_1269,In_1311);
xnor U2475 (N_2475,In_1457,In_1448);
and U2476 (N_2476,In_909,In_1414);
nor U2477 (N_2477,In_1052,In_436);
nand U2478 (N_2478,In_1456,In_505);
nand U2479 (N_2479,In_724,In_1329);
nor U2480 (N_2480,In_407,In_1147);
nand U2481 (N_2481,In_847,In_974);
nand U2482 (N_2482,In_1123,In_1212);
or U2483 (N_2483,In_1173,In_487);
and U2484 (N_2484,In_1141,In_922);
or U2485 (N_2485,In_253,In_1160);
and U2486 (N_2486,In_908,In_105);
and U2487 (N_2487,In_197,In_1170);
xor U2488 (N_2488,In_178,In_547);
and U2489 (N_2489,In_947,In_388);
nor U2490 (N_2490,In_1488,In_262);
and U2491 (N_2491,In_721,In_442);
nand U2492 (N_2492,In_153,In_1401);
nor U2493 (N_2493,In_885,In_1123);
nand U2494 (N_2494,In_9,In_78);
and U2495 (N_2495,In_751,In_874);
and U2496 (N_2496,In_1026,In_652);
or U2497 (N_2497,In_1458,In_1232);
nand U2498 (N_2498,In_38,In_81);
or U2499 (N_2499,In_739,In_664);
nand U2500 (N_2500,In_1027,In_345);
or U2501 (N_2501,In_1301,In_301);
and U2502 (N_2502,In_1048,In_409);
or U2503 (N_2503,In_482,In_600);
nor U2504 (N_2504,In_1198,In_1455);
and U2505 (N_2505,In_366,In_182);
nor U2506 (N_2506,In_136,In_56);
xnor U2507 (N_2507,In_1329,In_124);
nor U2508 (N_2508,In_549,In_354);
nor U2509 (N_2509,In_994,In_434);
or U2510 (N_2510,In_1192,In_526);
and U2511 (N_2511,In_657,In_15);
nor U2512 (N_2512,In_811,In_1239);
and U2513 (N_2513,In_1093,In_1392);
and U2514 (N_2514,In_205,In_258);
nor U2515 (N_2515,In_1244,In_745);
and U2516 (N_2516,In_30,In_182);
and U2517 (N_2517,In_369,In_1438);
and U2518 (N_2518,In_596,In_1183);
nor U2519 (N_2519,In_806,In_1134);
nand U2520 (N_2520,In_365,In_106);
nor U2521 (N_2521,In_43,In_490);
and U2522 (N_2522,In_1465,In_319);
nand U2523 (N_2523,In_1098,In_412);
or U2524 (N_2524,In_1488,In_809);
and U2525 (N_2525,In_907,In_83);
or U2526 (N_2526,In_443,In_1115);
or U2527 (N_2527,In_328,In_1321);
or U2528 (N_2528,In_537,In_599);
nand U2529 (N_2529,In_1459,In_844);
nand U2530 (N_2530,In_1403,In_881);
or U2531 (N_2531,In_1300,In_1262);
or U2532 (N_2532,In_1044,In_54);
and U2533 (N_2533,In_839,In_468);
and U2534 (N_2534,In_715,In_1232);
nor U2535 (N_2535,In_1434,In_652);
or U2536 (N_2536,In_253,In_1215);
nand U2537 (N_2537,In_782,In_923);
nor U2538 (N_2538,In_407,In_1458);
nand U2539 (N_2539,In_1073,In_1258);
or U2540 (N_2540,In_1240,In_476);
and U2541 (N_2541,In_1266,In_57);
and U2542 (N_2542,In_290,In_277);
or U2543 (N_2543,In_1028,In_403);
nor U2544 (N_2544,In_286,In_1019);
nand U2545 (N_2545,In_1356,In_1327);
nor U2546 (N_2546,In_691,In_708);
nor U2547 (N_2547,In_989,In_507);
nand U2548 (N_2548,In_363,In_856);
nand U2549 (N_2549,In_870,In_466);
nor U2550 (N_2550,In_291,In_546);
or U2551 (N_2551,In_461,In_1456);
or U2552 (N_2552,In_689,In_864);
and U2553 (N_2553,In_1377,In_175);
nor U2554 (N_2554,In_1230,In_563);
or U2555 (N_2555,In_1140,In_1101);
nor U2556 (N_2556,In_306,In_1313);
nor U2557 (N_2557,In_607,In_659);
nand U2558 (N_2558,In_1166,In_564);
nand U2559 (N_2559,In_82,In_660);
nand U2560 (N_2560,In_347,In_6);
nand U2561 (N_2561,In_790,In_943);
nand U2562 (N_2562,In_1074,In_6);
and U2563 (N_2563,In_658,In_478);
nor U2564 (N_2564,In_808,In_670);
nor U2565 (N_2565,In_1093,In_1097);
nand U2566 (N_2566,In_1416,In_314);
and U2567 (N_2567,In_67,In_900);
or U2568 (N_2568,In_413,In_753);
and U2569 (N_2569,In_1490,In_468);
nand U2570 (N_2570,In_935,In_1485);
nor U2571 (N_2571,In_638,In_74);
nor U2572 (N_2572,In_1089,In_388);
nand U2573 (N_2573,In_1344,In_1339);
nor U2574 (N_2574,In_839,In_424);
or U2575 (N_2575,In_1491,In_519);
or U2576 (N_2576,In_1078,In_318);
and U2577 (N_2577,In_244,In_1032);
nand U2578 (N_2578,In_842,In_489);
nor U2579 (N_2579,In_913,In_810);
and U2580 (N_2580,In_709,In_1215);
or U2581 (N_2581,In_426,In_872);
nand U2582 (N_2582,In_205,In_477);
and U2583 (N_2583,In_1236,In_688);
and U2584 (N_2584,In_7,In_39);
nand U2585 (N_2585,In_760,In_458);
nand U2586 (N_2586,In_1410,In_490);
nand U2587 (N_2587,In_195,In_433);
or U2588 (N_2588,In_751,In_22);
nor U2589 (N_2589,In_225,In_426);
nand U2590 (N_2590,In_1356,In_337);
and U2591 (N_2591,In_963,In_886);
nor U2592 (N_2592,In_635,In_1093);
or U2593 (N_2593,In_1171,In_1054);
or U2594 (N_2594,In_538,In_1206);
nand U2595 (N_2595,In_1189,In_72);
nor U2596 (N_2596,In_620,In_820);
and U2597 (N_2597,In_1055,In_763);
nor U2598 (N_2598,In_490,In_1322);
and U2599 (N_2599,In_509,In_129);
and U2600 (N_2600,In_664,In_458);
or U2601 (N_2601,In_1112,In_1368);
or U2602 (N_2602,In_267,In_413);
nor U2603 (N_2603,In_152,In_446);
and U2604 (N_2604,In_482,In_981);
or U2605 (N_2605,In_680,In_857);
or U2606 (N_2606,In_290,In_580);
or U2607 (N_2607,In_318,In_1400);
xor U2608 (N_2608,In_471,In_592);
and U2609 (N_2609,In_1070,In_573);
nor U2610 (N_2610,In_1400,In_167);
or U2611 (N_2611,In_1454,In_279);
and U2612 (N_2612,In_42,In_1474);
and U2613 (N_2613,In_309,In_442);
and U2614 (N_2614,In_1133,In_656);
nor U2615 (N_2615,In_479,In_1000);
nand U2616 (N_2616,In_420,In_1037);
nor U2617 (N_2617,In_1453,In_301);
and U2618 (N_2618,In_1074,In_34);
nand U2619 (N_2619,In_727,In_602);
nand U2620 (N_2620,In_553,In_1183);
nand U2621 (N_2621,In_787,In_1488);
and U2622 (N_2622,In_462,In_673);
nor U2623 (N_2623,In_1216,In_194);
or U2624 (N_2624,In_1331,In_592);
nand U2625 (N_2625,In_1493,In_1353);
or U2626 (N_2626,In_637,In_498);
nor U2627 (N_2627,In_621,In_1336);
or U2628 (N_2628,In_812,In_616);
xnor U2629 (N_2629,In_1478,In_23);
nor U2630 (N_2630,In_690,In_408);
or U2631 (N_2631,In_991,In_247);
nor U2632 (N_2632,In_812,In_548);
and U2633 (N_2633,In_1479,In_1396);
nand U2634 (N_2634,In_1133,In_1409);
or U2635 (N_2635,In_77,In_772);
nor U2636 (N_2636,In_600,In_723);
and U2637 (N_2637,In_995,In_920);
or U2638 (N_2638,In_797,In_985);
or U2639 (N_2639,In_1180,In_1210);
nand U2640 (N_2640,In_793,In_938);
nand U2641 (N_2641,In_1010,In_353);
nand U2642 (N_2642,In_700,In_553);
nand U2643 (N_2643,In_477,In_884);
nand U2644 (N_2644,In_689,In_914);
and U2645 (N_2645,In_378,In_592);
nor U2646 (N_2646,In_287,In_565);
nand U2647 (N_2647,In_805,In_665);
nor U2648 (N_2648,In_1106,In_1419);
or U2649 (N_2649,In_908,In_457);
nor U2650 (N_2650,In_447,In_121);
and U2651 (N_2651,In_267,In_1436);
or U2652 (N_2652,In_1325,In_614);
or U2653 (N_2653,In_1032,In_734);
or U2654 (N_2654,In_357,In_189);
nand U2655 (N_2655,In_1391,In_191);
nor U2656 (N_2656,In_918,In_1254);
nor U2657 (N_2657,In_58,In_761);
nand U2658 (N_2658,In_325,In_1418);
and U2659 (N_2659,In_558,In_1478);
nand U2660 (N_2660,In_1236,In_405);
nand U2661 (N_2661,In_347,In_1210);
and U2662 (N_2662,In_944,In_757);
and U2663 (N_2663,In_1446,In_636);
nand U2664 (N_2664,In_1153,In_1398);
and U2665 (N_2665,In_76,In_1331);
nor U2666 (N_2666,In_1249,In_1097);
nor U2667 (N_2667,In_1181,In_867);
nand U2668 (N_2668,In_192,In_96);
nor U2669 (N_2669,In_442,In_324);
nand U2670 (N_2670,In_1459,In_948);
nor U2671 (N_2671,In_296,In_1388);
and U2672 (N_2672,In_1172,In_751);
nor U2673 (N_2673,In_420,In_1206);
xnor U2674 (N_2674,In_1111,In_1366);
nor U2675 (N_2675,In_1479,In_1230);
nor U2676 (N_2676,In_40,In_1243);
nor U2677 (N_2677,In_773,In_105);
nor U2678 (N_2678,In_584,In_593);
and U2679 (N_2679,In_1320,In_910);
and U2680 (N_2680,In_803,In_1426);
and U2681 (N_2681,In_575,In_1007);
nand U2682 (N_2682,In_74,In_520);
and U2683 (N_2683,In_867,In_538);
xor U2684 (N_2684,In_85,In_87);
and U2685 (N_2685,In_268,In_1456);
and U2686 (N_2686,In_1152,In_290);
nor U2687 (N_2687,In_528,In_1032);
and U2688 (N_2688,In_581,In_1013);
and U2689 (N_2689,In_320,In_1069);
nand U2690 (N_2690,In_1310,In_1159);
or U2691 (N_2691,In_1252,In_340);
nor U2692 (N_2692,In_1130,In_554);
nor U2693 (N_2693,In_112,In_341);
xor U2694 (N_2694,In_1137,In_308);
nor U2695 (N_2695,In_147,In_284);
and U2696 (N_2696,In_531,In_1059);
nand U2697 (N_2697,In_825,In_1142);
or U2698 (N_2698,In_395,In_1379);
nand U2699 (N_2699,In_773,In_407);
and U2700 (N_2700,In_163,In_870);
nand U2701 (N_2701,In_566,In_354);
and U2702 (N_2702,In_1452,In_410);
nand U2703 (N_2703,In_716,In_1491);
nor U2704 (N_2704,In_466,In_812);
and U2705 (N_2705,In_679,In_636);
and U2706 (N_2706,In_1284,In_257);
nor U2707 (N_2707,In_240,In_1146);
nor U2708 (N_2708,In_119,In_348);
nand U2709 (N_2709,In_236,In_884);
nand U2710 (N_2710,In_382,In_1489);
or U2711 (N_2711,In_1100,In_1169);
or U2712 (N_2712,In_1177,In_557);
or U2713 (N_2713,In_1416,In_122);
or U2714 (N_2714,In_833,In_365);
and U2715 (N_2715,In_667,In_954);
and U2716 (N_2716,In_836,In_440);
or U2717 (N_2717,In_78,In_1423);
or U2718 (N_2718,In_941,In_835);
nand U2719 (N_2719,In_639,In_545);
nand U2720 (N_2720,In_724,In_1319);
nand U2721 (N_2721,In_553,In_862);
nor U2722 (N_2722,In_1445,In_871);
or U2723 (N_2723,In_90,In_215);
or U2724 (N_2724,In_446,In_1418);
or U2725 (N_2725,In_444,In_709);
and U2726 (N_2726,In_1182,In_474);
and U2727 (N_2727,In_1053,In_313);
nand U2728 (N_2728,In_443,In_47);
or U2729 (N_2729,In_1201,In_1182);
or U2730 (N_2730,In_176,In_942);
or U2731 (N_2731,In_1176,In_1408);
nand U2732 (N_2732,In_1198,In_1488);
and U2733 (N_2733,In_739,In_19);
and U2734 (N_2734,In_682,In_531);
nor U2735 (N_2735,In_293,In_860);
and U2736 (N_2736,In_361,In_412);
nor U2737 (N_2737,In_706,In_596);
nor U2738 (N_2738,In_594,In_620);
nor U2739 (N_2739,In_163,In_665);
and U2740 (N_2740,In_521,In_785);
nand U2741 (N_2741,In_668,In_1018);
and U2742 (N_2742,In_1291,In_461);
and U2743 (N_2743,In_630,In_1461);
or U2744 (N_2744,In_749,In_892);
or U2745 (N_2745,In_288,In_860);
nand U2746 (N_2746,In_162,In_1164);
and U2747 (N_2747,In_1442,In_575);
or U2748 (N_2748,In_482,In_1375);
and U2749 (N_2749,In_175,In_288);
nor U2750 (N_2750,In_1019,In_149);
nor U2751 (N_2751,In_47,In_745);
nand U2752 (N_2752,In_5,In_1329);
nor U2753 (N_2753,In_62,In_60);
nand U2754 (N_2754,In_103,In_35);
nor U2755 (N_2755,In_93,In_336);
nor U2756 (N_2756,In_430,In_864);
or U2757 (N_2757,In_1315,In_918);
or U2758 (N_2758,In_358,In_1272);
nor U2759 (N_2759,In_1045,In_234);
and U2760 (N_2760,In_54,In_93);
nor U2761 (N_2761,In_1114,In_1080);
and U2762 (N_2762,In_1475,In_190);
xnor U2763 (N_2763,In_788,In_930);
nor U2764 (N_2764,In_471,In_414);
nor U2765 (N_2765,In_720,In_1349);
nand U2766 (N_2766,In_815,In_635);
nor U2767 (N_2767,In_1411,In_1190);
and U2768 (N_2768,In_713,In_199);
nand U2769 (N_2769,In_994,In_766);
and U2770 (N_2770,In_1409,In_885);
or U2771 (N_2771,In_1236,In_978);
or U2772 (N_2772,In_1269,In_270);
or U2773 (N_2773,In_432,In_1493);
nand U2774 (N_2774,In_1258,In_1443);
nor U2775 (N_2775,In_279,In_521);
nor U2776 (N_2776,In_260,In_820);
or U2777 (N_2777,In_537,In_1134);
or U2778 (N_2778,In_239,In_199);
nand U2779 (N_2779,In_1263,In_736);
or U2780 (N_2780,In_1063,In_335);
or U2781 (N_2781,In_1482,In_648);
nand U2782 (N_2782,In_1111,In_912);
nand U2783 (N_2783,In_1032,In_811);
nor U2784 (N_2784,In_1297,In_1088);
xor U2785 (N_2785,In_686,In_225);
or U2786 (N_2786,In_535,In_980);
nand U2787 (N_2787,In_1441,In_1075);
and U2788 (N_2788,In_1234,In_587);
and U2789 (N_2789,In_393,In_639);
nor U2790 (N_2790,In_1037,In_1235);
and U2791 (N_2791,In_858,In_902);
or U2792 (N_2792,In_126,In_636);
xnor U2793 (N_2793,In_1064,In_71);
nand U2794 (N_2794,In_433,In_565);
nor U2795 (N_2795,In_607,In_1058);
or U2796 (N_2796,In_738,In_832);
nand U2797 (N_2797,In_1306,In_470);
or U2798 (N_2798,In_1121,In_218);
nor U2799 (N_2799,In_387,In_848);
or U2800 (N_2800,In_648,In_337);
and U2801 (N_2801,In_198,In_802);
and U2802 (N_2802,In_806,In_263);
nor U2803 (N_2803,In_1377,In_1420);
nand U2804 (N_2804,In_701,In_1066);
or U2805 (N_2805,In_1140,In_525);
nand U2806 (N_2806,In_949,In_1404);
or U2807 (N_2807,In_415,In_1047);
nand U2808 (N_2808,In_557,In_1353);
nand U2809 (N_2809,In_256,In_1480);
xnor U2810 (N_2810,In_1089,In_1349);
nand U2811 (N_2811,In_30,In_219);
nand U2812 (N_2812,In_1241,In_17);
and U2813 (N_2813,In_320,In_417);
or U2814 (N_2814,In_469,In_154);
or U2815 (N_2815,In_238,In_1304);
nor U2816 (N_2816,In_1113,In_84);
nand U2817 (N_2817,In_1078,In_1160);
nand U2818 (N_2818,In_856,In_948);
nand U2819 (N_2819,In_457,In_460);
and U2820 (N_2820,In_269,In_1470);
and U2821 (N_2821,In_575,In_907);
nand U2822 (N_2822,In_1289,In_381);
nor U2823 (N_2823,In_1098,In_1038);
and U2824 (N_2824,In_1393,In_1479);
and U2825 (N_2825,In_827,In_867);
and U2826 (N_2826,In_861,In_1106);
and U2827 (N_2827,In_1107,In_672);
nor U2828 (N_2828,In_840,In_500);
nor U2829 (N_2829,In_1301,In_797);
or U2830 (N_2830,In_23,In_175);
or U2831 (N_2831,In_1337,In_338);
and U2832 (N_2832,In_578,In_244);
nor U2833 (N_2833,In_201,In_266);
nor U2834 (N_2834,In_64,In_250);
and U2835 (N_2835,In_1020,In_758);
nand U2836 (N_2836,In_1204,In_100);
or U2837 (N_2837,In_983,In_389);
or U2838 (N_2838,In_181,In_861);
nor U2839 (N_2839,In_626,In_992);
nand U2840 (N_2840,In_1134,In_1350);
and U2841 (N_2841,In_710,In_678);
and U2842 (N_2842,In_1250,In_87);
nand U2843 (N_2843,In_854,In_930);
or U2844 (N_2844,In_1447,In_1212);
nor U2845 (N_2845,In_1227,In_1128);
and U2846 (N_2846,In_1081,In_157);
nor U2847 (N_2847,In_502,In_1235);
or U2848 (N_2848,In_666,In_1363);
and U2849 (N_2849,In_1368,In_826);
nand U2850 (N_2850,In_217,In_1311);
nand U2851 (N_2851,In_835,In_855);
or U2852 (N_2852,In_915,In_291);
and U2853 (N_2853,In_1344,In_838);
and U2854 (N_2854,In_173,In_290);
and U2855 (N_2855,In_1279,In_1165);
nand U2856 (N_2856,In_1195,In_655);
nand U2857 (N_2857,In_174,In_1183);
and U2858 (N_2858,In_312,In_1195);
nor U2859 (N_2859,In_1482,In_783);
and U2860 (N_2860,In_170,In_513);
nand U2861 (N_2861,In_1366,In_1189);
nand U2862 (N_2862,In_1456,In_696);
or U2863 (N_2863,In_1321,In_356);
nand U2864 (N_2864,In_409,In_146);
nand U2865 (N_2865,In_218,In_860);
or U2866 (N_2866,In_987,In_870);
nand U2867 (N_2867,In_978,In_1335);
or U2868 (N_2868,In_889,In_1005);
nand U2869 (N_2869,In_665,In_1352);
nor U2870 (N_2870,In_840,In_609);
or U2871 (N_2871,In_528,In_1359);
nor U2872 (N_2872,In_1089,In_278);
xnor U2873 (N_2873,In_1302,In_1321);
xnor U2874 (N_2874,In_982,In_1078);
nor U2875 (N_2875,In_128,In_1181);
xor U2876 (N_2876,In_80,In_1419);
xnor U2877 (N_2877,In_1245,In_320);
or U2878 (N_2878,In_499,In_1470);
and U2879 (N_2879,In_312,In_765);
or U2880 (N_2880,In_1193,In_641);
and U2881 (N_2881,In_815,In_669);
or U2882 (N_2882,In_8,In_1316);
and U2883 (N_2883,In_144,In_425);
nand U2884 (N_2884,In_1206,In_977);
nor U2885 (N_2885,In_453,In_588);
and U2886 (N_2886,In_225,In_844);
or U2887 (N_2887,In_165,In_1302);
or U2888 (N_2888,In_322,In_524);
or U2889 (N_2889,In_355,In_296);
and U2890 (N_2890,In_1203,In_1349);
nor U2891 (N_2891,In_1380,In_1460);
nor U2892 (N_2892,In_1477,In_1251);
or U2893 (N_2893,In_1065,In_1457);
and U2894 (N_2894,In_1370,In_890);
or U2895 (N_2895,In_541,In_291);
and U2896 (N_2896,In_1314,In_1411);
nand U2897 (N_2897,In_563,In_115);
and U2898 (N_2898,In_190,In_1068);
or U2899 (N_2899,In_50,In_440);
or U2900 (N_2900,In_802,In_1243);
nor U2901 (N_2901,In_1219,In_1362);
nand U2902 (N_2902,In_953,In_950);
xor U2903 (N_2903,In_738,In_607);
nand U2904 (N_2904,In_1103,In_1153);
nor U2905 (N_2905,In_1163,In_27);
or U2906 (N_2906,In_106,In_538);
xor U2907 (N_2907,In_608,In_1482);
nand U2908 (N_2908,In_756,In_591);
nor U2909 (N_2909,In_377,In_386);
nor U2910 (N_2910,In_559,In_953);
nand U2911 (N_2911,In_1182,In_1488);
or U2912 (N_2912,In_474,In_665);
and U2913 (N_2913,In_493,In_1425);
nand U2914 (N_2914,In_1224,In_1246);
nand U2915 (N_2915,In_993,In_1165);
nor U2916 (N_2916,In_1187,In_927);
nor U2917 (N_2917,In_323,In_557);
nor U2918 (N_2918,In_250,In_777);
or U2919 (N_2919,In_1077,In_261);
and U2920 (N_2920,In_1402,In_645);
and U2921 (N_2921,In_1457,In_81);
and U2922 (N_2922,In_1025,In_1277);
nand U2923 (N_2923,In_269,In_905);
and U2924 (N_2924,In_172,In_1095);
and U2925 (N_2925,In_578,In_682);
xor U2926 (N_2926,In_1074,In_736);
and U2927 (N_2927,In_100,In_1296);
and U2928 (N_2928,In_1480,In_86);
nor U2929 (N_2929,In_716,In_26);
and U2930 (N_2930,In_200,In_1158);
and U2931 (N_2931,In_980,In_274);
nor U2932 (N_2932,In_31,In_1042);
nor U2933 (N_2933,In_143,In_68);
and U2934 (N_2934,In_406,In_807);
or U2935 (N_2935,In_1468,In_385);
nor U2936 (N_2936,In_301,In_755);
or U2937 (N_2937,In_1028,In_838);
and U2938 (N_2938,In_1106,In_1493);
or U2939 (N_2939,In_668,In_225);
and U2940 (N_2940,In_1425,In_785);
nor U2941 (N_2941,In_900,In_201);
or U2942 (N_2942,In_59,In_361);
nand U2943 (N_2943,In_1198,In_1331);
nand U2944 (N_2944,In_355,In_120);
or U2945 (N_2945,In_738,In_352);
nand U2946 (N_2946,In_704,In_247);
and U2947 (N_2947,In_1338,In_339);
and U2948 (N_2948,In_850,In_200);
nor U2949 (N_2949,In_511,In_298);
nor U2950 (N_2950,In_1318,In_1284);
xnor U2951 (N_2951,In_1049,In_690);
nor U2952 (N_2952,In_968,In_1377);
and U2953 (N_2953,In_279,In_605);
or U2954 (N_2954,In_705,In_996);
or U2955 (N_2955,In_3,In_672);
nand U2956 (N_2956,In_676,In_611);
nor U2957 (N_2957,In_924,In_1286);
or U2958 (N_2958,In_237,In_875);
nand U2959 (N_2959,In_371,In_1369);
nand U2960 (N_2960,In_943,In_1253);
or U2961 (N_2961,In_1175,In_303);
and U2962 (N_2962,In_161,In_74);
nand U2963 (N_2963,In_53,In_547);
xor U2964 (N_2964,In_1337,In_340);
nand U2965 (N_2965,In_917,In_1048);
and U2966 (N_2966,In_808,In_1262);
nand U2967 (N_2967,In_1445,In_760);
nor U2968 (N_2968,In_67,In_1354);
nor U2969 (N_2969,In_473,In_76);
nor U2970 (N_2970,In_884,In_29);
nor U2971 (N_2971,In_348,In_1468);
and U2972 (N_2972,In_1432,In_1252);
nor U2973 (N_2973,In_1442,In_598);
xnor U2974 (N_2974,In_790,In_810);
and U2975 (N_2975,In_448,In_586);
and U2976 (N_2976,In_1250,In_297);
and U2977 (N_2977,In_962,In_1480);
nand U2978 (N_2978,In_629,In_186);
nand U2979 (N_2979,In_669,In_74);
nor U2980 (N_2980,In_536,In_1490);
nor U2981 (N_2981,In_989,In_509);
nand U2982 (N_2982,In_1360,In_308);
and U2983 (N_2983,In_750,In_299);
and U2984 (N_2984,In_68,In_929);
and U2985 (N_2985,In_1057,In_1227);
nand U2986 (N_2986,In_619,In_1422);
and U2987 (N_2987,In_1462,In_851);
xnor U2988 (N_2988,In_26,In_558);
or U2989 (N_2989,In_605,In_1419);
and U2990 (N_2990,In_889,In_349);
xnor U2991 (N_2991,In_1314,In_713);
nor U2992 (N_2992,In_1143,In_591);
nor U2993 (N_2993,In_76,In_1175);
and U2994 (N_2994,In_858,In_198);
nor U2995 (N_2995,In_179,In_1451);
nand U2996 (N_2996,In_1300,In_300);
and U2997 (N_2997,In_1212,In_1450);
xor U2998 (N_2998,In_618,In_737);
nand U2999 (N_2999,In_42,In_1055);
and U3000 (N_3000,In_1112,In_243);
and U3001 (N_3001,In_286,In_730);
nand U3002 (N_3002,In_962,In_1424);
and U3003 (N_3003,In_101,In_730);
nand U3004 (N_3004,In_365,In_337);
nor U3005 (N_3005,In_836,In_741);
and U3006 (N_3006,In_442,In_1072);
and U3007 (N_3007,In_802,In_440);
or U3008 (N_3008,In_544,In_114);
or U3009 (N_3009,In_446,In_39);
or U3010 (N_3010,In_505,In_106);
nor U3011 (N_3011,In_1274,In_281);
or U3012 (N_3012,In_631,In_303);
nand U3013 (N_3013,In_1229,In_560);
or U3014 (N_3014,In_1468,In_383);
nand U3015 (N_3015,In_809,In_1258);
and U3016 (N_3016,In_829,In_1290);
nand U3017 (N_3017,In_389,In_939);
nand U3018 (N_3018,In_88,In_76);
and U3019 (N_3019,In_56,In_57);
nand U3020 (N_3020,In_1241,In_173);
nor U3021 (N_3021,In_544,In_1285);
nand U3022 (N_3022,In_1340,In_175);
and U3023 (N_3023,In_152,In_204);
or U3024 (N_3024,In_316,In_64);
or U3025 (N_3025,In_1489,In_1139);
or U3026 (N_3026,In_406,In_397);
nor U3027 (N_3027,In_1332,In_1378);
nand U3028 (N_3028,In_594,In_1199);
nor U3029 (N_3029,In_7,In_779);
nor U3030 (N_3030,In_83,In_913);
or U3031 (N_3031,In_62,In_1350);
and U3032 (N_3032,In_1343,In_426);
nor U3033 (N_3033,In_356,In_1465);
nand U3034 (N_3034,In_640,In_83);
nor U3035 (N_3035,In_1159,In_533);
nor U3036 (N_3036,In_1312,In_598);
or U3037 (N_3037,In_329,In_1448);
nand U3038 (N_3038,In_383,In_1233);
nor U3039 (N_3039,In_930,In_1470);
nand U3040 (N_3040,In_811,In_613);
and U3041 (N_3041,In_133,In_825);
xnor U3042 (N_3042,In_1267,In_1212);
or U3043 (N_3043,In_149,In_747);
or U3044 (N_3044,In_649,In_1203);
and U3045 (N_3045,In_714,In_89);
and U3046 (N_3046,In_229,In_529);
and U3047 (N_3047,In_96,In_613);
or U3048 (N_3048,In_427,In_102);
nand U3049 (N_3049,In_88,In_251);
and U3050 (N_3050,In_185,In_1231);
nor U3051 (N_3051,In_319,In_913);
or U3052 (N_3052,In_46,In_751);
or U3053 (N_3053,In_408,In_194);
nor U3054 (N_3054,In_269,In_866);
and U3055 (N_3055,In_437,In_51);
and U3056 (N_3056,In_752,In_222);
nor U3057 (N_3057,In_182,In_784);
nand U3058 (N_3058,In_620,In_408);
xnor U3059 (N_3059,In_716,In_1273);
or U3060 (N_3060,In_521,In_1036);
and U3061 (N_3061,In_1369,In_1398);
nor U3062 (N_3062,In_926,In_540);
or U3063 (N_3063,In_566,In_1334);
nand U3064 (N_3064,In_972,In_614);
nand U3065 (N_3065,In_148,In_600);
and U3066 (N_3066,In_194,In_902);
nor U3067 (N_3067,In_576,In_569);
nor U3068 (N_3068,In_520,In_1194);
and U3069 (N_3069,In_1435,In_1347);
and U3070 (N_3070,In_452,In_550);
or U3071 (N_3071,In_1409,In_1132);
nor U3072 (N_3072,In_77,In_17);
nor U3073 (N_3073,In_1419,In_565);
or U3074 (N_3074,In_493,In_158);
nand U3075 (N_3075,In_319,In_568);
and U3076 (N_3076,In_852,In_780);
nor U3077 (N_3077,In_139,In_417);
nand U3078 (N_3078,In_63,In_3);
nand U3079 (N_3079,In_950,In_1160);
or U3080 (N_3080,In_188,In_1292);
nand U3081 (N_3081,In_994,In_1232);
xnor U3082 (N_3082,In_176,In_913);
nor U3083 (N_3083,In_608,In_126);
or U3084 (N_3084,In_1115,In_557);
and U3085 (N_3085,In_350,In_138);
and U3086 (N_3086,In_1400,In_142);
nand U3087 (N_3087,In_1486,In_378);
or U3088 (N_3088,In_568,In_193);
nor U3089 (N_3089,In_1064,In_123);
nand U3090 (N_3090,In_75,In_112);
nor U3091 (N_3091,In_1151,In_296);
nor U3092 (N_3092,In_1468,In_270);
or U3093 (N_3093,In_377,In_1248);
xor U3094 (N_3094,In_235,In_829);
xnor U3095 (N_3095,In_984,In_562);
and U3096 (N_3096,In_960,In_366);
or U3097 (N_3097,In_1001,In_148);
nor U3098 (N_3098,In_139,In_291);
and U3099 (N_3099,In_309,In_1277);
and U3100 (N_3100,In_668,In_1087);
or U3101 (N_3101,In_1174,In_302);
or U3102 (N_3102,In_1240,In_1360);
nor U3103 (N_3103,In_276,In_390);
xor U3104 (N_3104,In_824,In_690);
and U3105 (N_3105,In_678,In_1000);
or U3106 (N_3106,In_238,In_1044);
nand U3107 (N_3107,In_814,In_1082);
nand U3108 (N_3108,In_1025,In_652);
nand U3109 (N_3109,In_1367,In_1410);
or U3110 (N_3110,In_994,In_36);
nor U3111 (N_3111,In_663,In_231);
nand U3112 (N_3112,In_539,In_186);
and U3113 (N_3113,In_301,In_235);
and U3114 (N_3114,In_1355,In_155);
and U3115 (N_3115,In_340,In_297);
nor U3116 (N_3116,In_1400,In_1279);
and U3117 (N_3117,In_399,In_1131);
nor U3118 (N_3118,In_1454,In_74);
and U3119 (N_3119,In_386,In_1437);
or U3120 (N_3120,In_545,In_1272);
and U3121 (N_3121,In_132,In_411);
nand U3122 (N_3122,In_1205,In_1131);
nand U3123 (N_3123,In_88,In_660);
nor U3124 (N_3124,In_516,In_1426);
nor U3125 (N_3125,In_355,In_1210);
and U3126 (N_3126,In_1468,In_586);
or U3127 (N_3127,In_1320,In_537);
nand U3128 (N_3128,In_270,In_455);
nor U3129 (N_3129,In_756,In_390);
nand U3130 (N_3130,In_1228,In_861);
nand U3131 (N_3131,In_317,In_729);
or U3132 (N_3132,In_861,In_245);
nor U3133 (N_3133,In_1454,In_163);
xor U3134 (N_3134,In_364,In_981);
and U3135 (N_3135,In_1409,In_30);
nor U3136 (N_3136,In_986,In_1146);
and U3137 (N_3137,In_32,In_1192);
and U3138 (N_3138,In_330,In_513);
nand U3139 (N_3139,In_690,In_492);
nand U3140 (N_3140,In_12,In_501);
nand U3141 (N_3141,In_965,In_655);
nor U3142 (N_3142,In_693,In_4);
or U3143 (N_3143,In_1424,In_1337);
nor U3144 (N_3144,In_507,In_690);
nand U3145 (N_3145,In_413,In_1297);
or U3146 (N_3146,In_744,In_540);
nand U3147 (N_3147,In_306,In_116);
nand U3148 (N_3148,In_594,In_182);
or U3149 (N_3149,In_1139,In_234);
and U3150 (N_3150,In_185,In_490);
nand U3151 (N_3151,In_823,In_1465);
nor U3152 (N_3152,In_986,In_741);
nor U3153 (N_3153,In_831,In_741);
and U3154 (N_3154,In_133,In_850);
nor U3155 (N_3155,In_1318,In_1245);
and U3156 (N_3156,In_1200,In_1136);
and U3157 (N_3157,In_177,In_383);
nor U3158 (N_3158,In_158,In_632);
nor U3159 (N_3159,In_39,In_380);
nor U3160 (N_3160,In_468,In_1419);
or U3161 (N_3161,In_989,In_1439);
nor U3162 (N_3162,In_651,In_583);
and U3163 (N_3163,In_285,In_239);
nand U3164 (N_3164,In_797,In_362);
and U3165 (N_3165,In_1061,In_92);
nor U3166 (N_3166,In_1367,In_1353);
or U3167 (N_3167,In_176,In_539);
and U3168 (N_3168,In_1008,In_981);
or U3169 (N_3169,In_310,In_279);
nor U3170 (N_3170,In_949,In_922);
xnor U3171 (N_3171,In_1080,In_733);
nand U3172 (N_3172,In_928,In_64);
or U3173 (N_3173,In_842,In_617);
and U3174 (N_3174,In_94,In_1471);
nor U3175 (N_3175,In_113,In_1293);
and U3176 (N_3176,In_1440,In_596);
nor U3177 (N_3177,In_29,In_1105);
or U3178 (N_3178,In_1305,In_1209);
nand U3179 (N_3179,In_1174,In_849);
nor U3180 (N_3180,In_511,In_440);
or U3181 (N_3181,In_1165,In_1237);
and U3182 (N_3182,In_467,In_78);
nor U3183 (N_3183,In_1074,In_515);
nand U3184 (N_3184,In_866,In_455);
nand U3185 (N_3185,In_556,In_388);
nor U3186 (N_3186,In_856,In_262);
nor U3187 (N_3187,In_267,In_1135);
nor U3188 (N_3188,In_438,In_142);
nand U3189 (N_3189,In_415,In_945);
and U3190 (N_3190,In_724,In_1196);
nor U3191 (N_3191,In_221,In_775);
and U3192 (N_3192,In_154,In_33);
and U3193 (N_3193,In_747,In_1229);
nor U3194 (N_3194,In_632,In_240);
nor U3195 (N_3195,In_405,In_1363);
nand U3196 (N_3196,In_1217,In_315);
nand U3197 (N_3197,In_1188,In_767);
or U3198 (N_3198,In_797,In_249);
or U3199 (N_3199,In_714,In_31);
or U3200 (N_3200,In_882,In_1499);
and U3201 (N_3201,In_375,In_200);
nor U3202 (N_3202,In_696,In_1346);
or U3203 (N_3203,In_252,In_917);
nand U3204 (N_3204,In_1365,In_1079);
nand U3205 (N_3205,In_1314,In_198);
and U3206 (N_3206,In_126,In_213);
or U3207 (N_3207,In_855,In_156);
and U3208 (N_3208,In_57,In_467);
nor U3209 (N_3209,In_1162,In_1293);
or U3210 (N_3210,In_178,In_534);
and U3211 (N_3211,In_55,In_1053);
and U3212 (N_3212,In_398,In_798);
and U3213 (N_3213,In_113,In_1203);
nand U3214 (N_3214,In_225,In_494);
or U3215 (N_3215,In_534,In_613);
xnor U3216 (N_3216,In_284,In_341);
nand U3217 (N_3217,In_1491,In_1068);
and U3218 (N_3218,In_896,In_388);
nand U3219 (N_3219,In_970,In_1146);
or U3220 (N_3220,In_1432,In_954);
xnor U3221 (N_3221,In_1339,In_1368);
nand U3222 (N_3222,In_1318,In_573);
and U3223 (N_3223,In_67,In_249);
or U3224 (N_3224,In_1234,In_179);
xnor U3225 (N_3225,In_1445,In_146);
or U3226 (N_3226,In_955,In_669);
and U3227 (N_3227,In_1110,In_1450);
or U3228 (N_3228,In_910,In_36);
nand U3229 (N_3229,In_1094,In_1350);
and U3230 (N_3230,In_1270,In_887);
nand U3231 (N_3231,In_1349,In_1245);
or U3232 (N_3232,In_1310,In_1297);
nor U3233 (N_3233,In_468,In_1412);
nor U3234 (N_3234,In_940,In_1085);
nand U3235 (N_3235,In_343,In_712);
and U3236 (N_3236,In_1154,In_1107);
or U3237 (N_3237,In_1024,In_1263);
nand U3238 (N_3238,In_1084,In_1267);
and U3239 (N_3239,In_666,In_802);
nor U3240 (N_3240,In_1254,In_1309);
and U3241 (N_3241,In_964,In_883);
or U3242 (N_3242,In_1363,In_1055);
nand U3243 (N_3243,In_1002,In_76);
nand U3244 (N_3244,In_1479,In_146);
nand U3245 (N_3245,In_728,In_297);
and U3246 (N_3246,In_167,In_512);
or U3247 (N_3247,In_864,In_137);
or U3248 (N_3248,In_482,In_828);
or U3249 (N_3249,In_1167,In_1126);
and U3250 (N_3250,In_1065,In_1307);
nand U3251 (N_3251,In_644,In_905);
and U3252 (N_3252,In_1397,In_570);
and U3253 (N_3253,In_127,In_47);
and U3254 (N_3254,In_817,In_1079);
nor U3255 (N_3255,In_500,In_1092);
or U3256 (N_3256,In_1154,In_312);
nand U3257 (N_3257,In_1171,In_1042);
nand U3258 (N_3258,In_229,In_878);
or U3259 (N_3259,In_1242,In_1383);
and U3260 (N_3260,In_1238,In_500);
and U3261 (N_3261,In_184,In_1182);
nor U3262 (N_3262,In_432,In_813);
nand U3263 (N_3263,In_1109,In_1465);
or U3264 (N_3264,In_888,In_1329);
nand U3265 (N_3265,In_770,In_109);
or U3266 (N_3266,In_1000,In_1346);
nand U3267 (N_3267,In_574,In_851);
and U3268 (N_3268,In_417,In_1189);
and U3269 (N_3269,In_1027,In_443);
nor U3270 (N_3270,In_860,In_727);
nand U3271 (N_3271,In_120,In_2);
nand U3272 (N_3272,In_955,In_19);
or U3273 (N_3273,In_123,In_378);
and U3274 (N_3274,In_1305,In_113);
or U3275 (N_3275,In_343,In_961);
or U3276 (N_3276,In_37,In_1265);
and U3277 (N_3277,In_1445,In_618);
or U3278 (N_3278,In_1100,In_1232);
nor U3279 (N_3279,In_371,In_68);
and U3280 (N_3280,In_603,In_1441);
nor U3281 (N_3281,In_681,In_589);
nand U3282 (N_3282,In_932,In_1082);
nor U3283 (N_3283,In_455,In_774);
or U3284 (N_3284,In_670,In_1388);
nand U3285 (N_3285,In_1093,In_353);
and U3286 (N_3286,In_645,In_1469);
and U3287 (N_3287,In_557,In_822);
and U3288 (N_3288,In_1064,In_575);
nand U3289 (N_3289,In_832,In_397);
nand U3290 (N_3290,In_94,In_1064);
or U3291 (N_3291,In_1131,In_650);
and U3292 (N_3292,In_258,In_15);
and U3293 (N_3293,In_1416,In_203);
and U3294 (N_3294,In_1303,In_331);
or U3295 (N_3295,In_1082,In_746);
nor U3296 (N_3296,In_17,In_390);
nor U3297 (N_3297,In_1193,In_1480);
nand U3298 (N_3298,In_1076,In_868);
and U3299 (N_3299,In_598,In_449);
and U3300 (N_3300,In_851,In_1189);
nand U3301 (N_3301,In_262,In_1035);
nand U3302 (N_3302,In_1154,In_1153);
or U3303 (N_3303,In_613,In_1001);
nand U3304 (N_3304,In_1490,In_494);
and U3305 (N_3305,In_1298,In_576);
nor U3306 (N_3306,In_312,In_434);
and U3307 (N_3307,In_734,In_960);
nor U3308 (N_3308,In_623,In_1484);
and U3309 (N_3309,In_505,In_1339);
nand U3310 (N_3310,In_878,In_384);
nor U3311 (N_3311,In_260,In_598);
nor U3312 (N_3312,In_841,In_504);
or U3313 (N_3313,In_275,In_795);
nor U3314 (N_3314,In_1307,In_79);
nor U3315 (N_3315,In_523,In_1148);
nor U3316 (N_3316,In_119,In_36);
nand U3317 (N_3317,In_1138,In_40);
or U3318 (N_3318,In_513,In_385);
and U3319 (N_3319,In_1104,In_574);
and U3320 (N_3320,In_755,In_395);
nor U3321 (N_3321,In_1233,In_1261);
nand U3322 (N_3322,In_257,In_541);
and U3323 (N_3323,In_110,In_720);
nand U3324 (N_3324,In_129,In_1011);
or U3325 (N_3325,In_1309,In_826);
nand U3326 (N_3326,In_1408,In_1244);
and U3327 (N_3327,In_1144,In_909);
nand U3328 (N_3328,In_1325,In_717);
nand U3329 (N_3329,In_22,In_138);
or U3330 (N_3330,In_767,In_832);
and U3331 (N_3331,In_459,In_344);
nand U3332 (N_3332,In_1427,In_421);
nand U3333 (N_3333,In_1480,In_679);
or U3334 (N_3334,In_308,In_713);
nor U3335 (N_3335,In_1308,In_163);
nor U3336 (N_3336,In_530,In_977);
nand U3337 (N_3337,In_942,In_803);
and U3338 (N_3338,In_525,In_748);
or U3339 (N_3339,In_362,In_1250);
and U3340 (N_3340,In_294,In_155);
nand U3341 (N_3341,In_1374,In_288);
nor U3342 (N_3342,In_915,In_378);
or U3343 (N_3343,In_1395,In_289);
nand U3344 (N_3344,In_156,In_933);
nor U3345 (N_3345,In_827,In_791);
nand U3346 (N_3346,In_55,In_142);
nand U3347 (N_3347,In_718,In_488);
and U3348 (N_3348,In_755,In_296);
and U3349 (N_3349,In_284,In_1230);
nand U3350 (N_3350,In_1181,In_237);
nor U3351 (N_3351,In_1383,In_103);
or U3352 (N_3352,In_61,In_143);
xnor U3353 (N_3353,In_1123,In_1395);
nor U3354 (N_3354,In_780,In_787);
and U3355 (N_3355,In_1296,In_1163);
nor U3356 (N_3356,In_1027,In_876);
and U3357 (N_3357,In_494,In_567);
and U3358 (N_3358,In_441,In_875);
and U3359 (N_3359,In_1323,In_991);
or U3360 (N_3360,In_84,In_460);
and U3361 (N_3361,In_1166,In_1225);
nand U3362 (N_3362,In_1162,In_507);
nand U3363 (N_3363,In_602,In_660);
nand U3364 (N_3364,In_852,In_1439);
and U3365 (N_3365,In_405,In_1150);
and U3366 (N_3366,In_762,In_361);
nor U3367 (N_3367,In_966,In_1213);
nand U3368 (N_3368,In_565,In_1498);
nor U3369 (N_3369,In_178,In_518);
nor U3370 (N_3370,In_124,In_1213);
nand U3371 (N_3371,In_1342,In_79);
and U3372 (N_3372,In_843,In_1053);
nand U3373 (N_3373,In_642,In_1330);
nor U3374 (N_3374,In_718,In_188);
and U3375 (N_3375,In_1024,In_1198);
nand U3376 (N_3376,In_1042,In_979);
xor U3377 (N_3377,In_720,In_254);
or U3378 (N_3378,In_1038,In_60);
and U3379 (N_3379,In_484,In_389);
nand U3380 (N_3380,In_1144,In_1107);
nor U3381 (N_3381,In_775,In_903);
nor U3382 (N_3382,In_1487,In_373);
nor U3383 (N_3383,In_483,In_85);
nor U3384 (N_3384,In_784,In_564);
nor U3385 (N_3385,In_405,In_209);
nor U3386 (N_3386,In_809,In_525);
nand U3387 (N_3387,In_999,In_863);
or U3388 (N_3388,In_520,In_423);
and U3389 (N_3389,In_148,In_583);
or U3390 (N_3390,In_978,In_556);
nor U3391 (N_3391,In_1128,In_1229);
nand U3392 (N_3392,In_673,In_468);
nand U3393 (N_3393,In_1389,In_1134);
nand U3394 (N_3394,In_48,In_725);
and U3395 (N_3395,In_1405,In_854);
or U3396 (N_3396,In_1352,In_1251);
and U3397 (N_3397,In_672,In_155);
or U3398 (N_3398,In_811,In_997);
nand U3399 (N_3399,In_1210,In_838);
and U3400 (N_3400,In_1257,In_361);
nor U3401 (N_3401,In_1437,In_590);
or U3402 (N_3402,In_556,In_170);
nand U3403 (N_3403,In_820,In_353);
nand U3404 (N_3404,In_882,In_417);
and U3405 (N_3405,In_411,In_741);
or U3406 (N_3406,In_491,In_349);
and U3407 (N_3407,In_682,In_402);
or U3408 (N_3408,In_1418,In_896);
or U3409 (N_3409,In_316,In_1165);
and U3410 (N_3410,In_1040,In_642);
nand U3411 (N_3411,In_917,In_253);
or U3412 (N_3412,In_1290,In_351);
nor U3413 (N_3413,In_1481,In_1391);
and U3414 (N_3414,In_1048,In_627);
xnor U3415 (N_3415,In_226,In_1305);
and U3416 (N_3416,In_1083,In_968);
or U3417 (N_3417,In_1088,In_1374);
nor U3418 (N_3418,In_1229,In_773);
and U3419 (N_3419,In_1084,In_930);
nor U3420 (N_3420,In_260,In_617);
nand U3421 (N_3421,In_1099,In_995);
or U3422 (N_3422,In_1084,In_1281);
and U3423 (N_3423,In_433,In_29);
nor U3424 (N_3424,In_323,In_946);
and U3425 (N_3425,In_1129,In_1373);
xor U3426 (N_3426,In_890,In_1207);
and U3427 (N_3427,In_506,In_697);
nor U3428 (N_3428,In_489,In_1197);
nor U3429 (N_3429,In_953,In_814);
or U3430 (N_3430,In_165,In_256);
or U3431 (N_3431,In_88,In_1155);
nor U3432 (N_3432,In_749,In_97);
nand U3433 (N_3433,In_225,In_1084);
nor U3434 (N_3434,In_0,In_1198);
nand U3435 (N_3435,In_168,In_1121);
xor U3436 (N_3436,In_888,In_1130);
nor U3437 (N_3437,In_1159,In_755);
xnor U3438 (N_3438,In_1220,In_643);
nor U3439 (N_3439,In_1362,In_182);
or U3440 (N_3440,In_515,In_52);
or U3441 (N_3441,In_1011,In_1361);
and U3442 (N_3442,In_243,In_920);
nor U3443 (N_3443,In_274,In_683);
nor U3444 (N_3444,In_137,In_1041);
nand U3445 (N_3445,In_661,In_210);
nor U3446 (N_3446,In_1300,In_1256);
nor U3447 (N_3447,In_629,In_121);
nand U3448 (N_3448,In_734,In_269);
nor U3449 (N_3449,In_1283,In_327);
or U3450 (N_3450,In_197,In_1123);
and U3451 (N_3451,In_639,In_301);
and U3452 (N_3452,In_519,In_1231);
nand U3453 (N_3453,In_549,In_565);
nand U3454 (N_3454,In_37,In_351);
or U3455 (N_3455,In_1451,In_372);
and U3456 (N_3456,In_667,In_1169);
nor U3457 (N_3457,In_598,In_1113);
or U3458 (N_3458,In_238,In_1263);
nand U3459 (N_3459,In_1279,In_1287);
and U3460 (N_3460,In_517,In_1212);
and U3461 (N_3461,In_1334,In_1094);
nor U3462 (N_3462,In_971,In_191);
nor U3463 (N_3463,In_490,In_1227);
nor U3464 (N_3464,In_1447,In_500);
and U3465 (N_3465,In_273,In_537);
nor U3466 (N_3466,In_540,In_87);
or U3467 (N_3467,In_1239,In_222);
xor U3468 (N_3468,In_1356,In_555);
nand U3469 (N_3469,In_365,In_694);
or U3470 (N_3470,In_739,In_1014);
nor U3471 (N_3471,In_1414,In_930);
nand U3472 (N_3472,In_140,In_226);
or U3473 (N_3473,In_50,In_984);
nand U3474 (N_3474,In_869,In_1159);
nor U3475 (N_3475,In_691,In_553);
and U3476 (N_3476,In_1417,In_211);
or U3477 (N_3477,In_1183,In_416);
or U3478 (N_3478,In_108,In_525);
nor U3479 (N_3479,In_1041,In_1497);
and U3480 (N_3480,In_703,In_681);
nor U3481 (N_3481,In_1060,In_722);
nand U3482 (N_3482,In_1133,In_632);
nand U3483 (N_3483,In_494,In_24);
and U3484 (N_3484,In_855,In_687);
and U3485 (N_3485,In_1414,In_130);
and U3486 (N_3486,In_592,In_1443);
or U3487 (N_3487,In_27,In_1421);
nand U3488 (N_3488,In_215,In_1053);
nor U3489 (N_3489,In_258,In_330);
nor U3490 (N_3490,In_314,In_842);
nor U3491 (N_3491,In_622,In_1377);
nand U3492 (N_3492,In_227,In_629);
nor U3493 (N_3493,In_186,In_891);
nand U3494 (N_3494,In_882,In_402);
and U3495 (N_3495,In_823,In_487);
nand U3496 (N_3496,In_755,In_854);
and U3497 (N_3497,In_875,In_573);
nor U3498 (N_3498,In_711,In_609);
and U3499 (N_3499,In_449,In_7);
or U3500 (N_3500,In_410,In_1245);
nand U3501 (N_3501,In_1356,In_1033);
and U3502 (N_3502,In_787,In_1479);
or U3503 (N_3503,In_1196,In_1039);
and U3504 (N_3504,In_73,In_1367);
or U3505 (N_3505,In_1286,In_1342);
xor U3506 (N_3506,In_800,In_44);
nand U3507 (N_3507,In_977,In_97);
nor U3508 (N_3508,In_666,In_111);
nor U3509 (N_3509,In_598,In_273);
nand U3510 (N_3510,In_410,In_1287);
nand U3511 (N_3511,In_456,In_188);
nor U3512 (N_3512,In_326,In_993);
nand U3513 (N_3513,In_839,In_89);
or U3514 (N_3514,In_891,In_928);
nor U3515 (N_3515,In_1125,In_1021);
xnor U3516 (N_3516,In_618,In_643);
or U3517 (N_3517,In_737,In_994);
nand U3518 (N_3518,In_872,In_36);
nor U3519 (N_3519,In_1106,In_1484);
and U3520 (N_3520,In_356,In_65);
and U3521 (N_3521,In_714,In_195);
and U3522 (N_3522,In_942,In_313);
and U3523 (N_3523,In_914,In_1148);
or U3524 (N_3524,In_1171,In_494);
nor U3525 (N_3525,In_1128,In_1280);
nor U3526 (N_3526,In_606,In_143);
nand U3527 (N_3527,In_1110,In_602);
and U3528 (N_3528,In_479,In_1201);
nand U3529 (N_3529,In_1250,In_882);
nor U3530 (N_3530,In_1471,In_102);
or U3531 (N_3531,In_7,In_968);
nand U3532 (N_3532,In_317,In_543);
and U3533 (N_3533,In_579,In_694);
and U3534 (N_3534,In_5,In_697);
nand U3535 (N_3535,In_1446,In_858);
nor U3536 (N_3536,In_759,In_521);
nor U3537 (N_3537,In_1059,In_630);
nor U3538 (N_3538,In_1133,In_757);
and U3539 (N_3539,In_27,In_751);
or U3540 (N_3540,In_1083,In_60);
and U3541 (N_3541,In_680,In_178);
nor U3542 (N_3542,In_253,In_858);
nand U3543 (N_3543,In_551,In_877);
and U3544 (N_3544,In_953,In_1225);
or U3545 (N_3545,In_739,In_605);
nor U3546 (N_3546,In_849,In_1365);
nor U3547 (N_3547,In_1168,In_902);
or U3548 (N_3548,In_395,In_303);
and U3549 (N_3549,In_567,In_1394);
nor U3550 (N_3550,In_1418,In_1173);
nor U3551 (N_3551,In_568,In_838);
or U3552 (N_3552,In_117,In_554);
nand U3553 (N_3553,In_103,In_886);
nand U3554 (N_3554,In_496,In_318);
nand U3555 (N_3555,In_948,In_465);
or U3556 (N_3556,In_339,In_1270);
and U3557 (N_3557,In_348,In_1029);
nor U3558 (N_3558,In_84,In_1404);
and U3559 (N_3559,In_207,In_85);
nor U3560 (N_3560,In_137,In_1163);
nor U3561 (N_3561,In_957,In_314);
or U3562 (N_3562,In_855,In_1211);
nor U3563 (N_3563,In_654,In_286);
nand U3564 (N_3564,In_518,In_453);
or U3565 (N_3565,In_894,In_906);
nor U3566 (N_3566,In_1140,In_1128);
nand U3567 (N_3567,In_138,In_1044);
and U3568 (N_3568,In_689,In_446);
nor U3569 (N_3569,In_1210,In_850);
and U3570 (N_3570,In_170,In_1023);
or U3571 (N_3571,In_546,In_1044);
nor U3572 (N_3572,In_985,In_107);
nand U3573 (N_3573,In_567,In_719);
nand U3574 (N_3574,In_411,In_1231);
nor U3575 (N_3575,In_470,In_1428);
xnor U3576 (N_3576,In_1190,In_342);
nor U3577 (N_3577,In_419,In_124);
and U3578 (N_3578,In_1245,In_734);
nor U3579 (N_3579,In_580,In_442);
and U3580 (N_3580,In_288,In_1207);
and U3581 (N_3581,In_1186,In_747);
or U3582 (N_3582,In_796,In_64);
and U3583 (N_3583,In_752,In_1240);
nor U3584 (N_3584,In_139,In_1468);
nand U3585 (N_3585,In_1043,In_330);
nand U3586 (N_3586,In_1414,In_1198);
and U3587 (N_3587,In_1188,In_708);
and U3588 (N_3588,In_333,In_326);
and U3589 (N_3589,In_1497,In_920);
nor U3590 (N_3590,In_575,In_783);
and U3591 (N_3591,In_765,In_1280);
and U3592 (N_3592,In_557,In_518);
and U3593 (N_3593,In_442,In_395);
or U3594 (N_3594,In_741,In_1079);
and U3595 (N_3595,In_549,In_331);
nand U3596 (N_3596,In_92,In_845);
nor U3597 (N_3597,In_1150,In_285);
and U3598 (N_3598,In_1147,In_74);
nor U3599 (N_3599,In_1209,In_42);
nor U3600 (N_3600,In_657,In_1485);
and U3601 (N_3601,In_894,In_438);
xor U3602 (N_3602,In_1075,In_135);
nor U3603 (N_3603,In_1183,In_536);
nor U3604 (N_3604,In_219,In_1102);
nor U3605 (N_3605,In_499,In_753);
nand U3606 (N_3606,In_1330,In_546);
nand U3607 (N_3607,In_275,In_579);
nor U3608 (N_3608,In_957,In_381);
nor U3609 (N_3609,In_322,In_1294);
nor U3610 (N_3610,In_953,In_151);
and U3611 (N_3611,In_224,In_1369);
xnor U3612 (N_3612,In_1437,In_1131);
or U3613 (N_3613,In_1415,In_873);
nor U3614 (N_3614,In_967,In_765);
or U3615 (N_3615,In_1364,In_449);
nor U3616 (N_3616,In_524,In_1279);
and U3617 (N_3617,In_496,In_1278);
nor U3618 (N_3618,In_325,In_295);
or U3619 (N_3619,In_985,In_1146);
nand U3620 (N_3620,In_743,In_403);
nor U3621 (N_3621,In_1478,In_301);
and U3622 (N_3622,In_784,In_1214);
nand U3623 (N_3623,In_1314,In_297);
or U3624 (N_3624,In_719,In_87);
nor U3625 (N_3625,In_285,In_693);
nand U3626 (N_3626,In_1445,In_487);
nand U3627 (N_3627,In_683,In_335);
and U3628 (N_3628,In_1372,In_186);
or U3629 (N_3629,In_1304,In_253);
xor U3630 (N_3630,In_89,In_1030);
nand U3631 (N_3631,In_267,In_1013);
and U3632 (N_3632,In_642,In_72);
or U3633 (N_3633,In_609,In_793);
and U3634 (N_3634,In_644,In_1375);
and U3635 (N_3635,In_1069,In_1336);
nor U3636 (N_3636,In_680,In_684);
or U3637 (N_3637,In_706,In_1311);
or U3638 (N_3638,In_543,In_1309);
nor U3639 (N_3639,In_1304,In_1152);
and U3640 (N_3640,In_1309,In_1305);
xnor U3641 (N_3641,In_1357,In_1226);
and U3642 (N_3642,In_657,In_1125);
nand U3643 (N_3643,In_1123,In_1479);
and U3644 (N_3644,In_1172,In_211);
or U3645 (N_3645,In_128,In_922);
or U3646 (N_3646,In_773,In_1387);
nand U3647 (N_3647,In_619,In_477);
and U3648 (N_3648,In_427,In_1378);
or U3649 (N_3649,In_1223,In_548);
or U3650 (N_3650,In_1015,In_168);
nand U3651 (N_3651,In_263,In_1476);
or U3652 (N_3652,In_404,In_1391);
nand U3653 (N_3653,In_713,In_781);
nor U3654 (N_3654,In_1099,In_286);
or U3655 (N_3655,In_984,In_328);
nand U3656 (N_3656,In_83,In_629);
nor U3657 (N_3657,In_1179,In_1371);
nand U3658 (N_3658,In_583,In_162);
nand U3659 (N_3659,In_825,In_23);
nor U3660 (N_3660,In_89,In_1295);
nand U3661 (N_3661,In_371,In_1404);
or U3662 (N_3662,In_71,In_519);
and U3663 (N_3663,In_254,In_105);
nor U3664 (N_3664,In_8,In_612);
and U3665 (N_3665,In_12,In_831);
nand U3666 (N_3666,In_626,In_156);
or U3667 (N_3667,In_1018,In_154);
or U3668 (N_3668,In_1300,In_37);
or U3669 (N_3669,In_1021,In_1129);
nor U3670 (N_3670,In_1171,In_1048);
nand U3671 (N_3671,In_672,In_1121);
and U3672 (N_3672,In_175,In_1477);
or U3673 (N_3673,In_251,In_203);
and U3674 (N_3674,In_1341,In_755);
nand U3675 (N_3675,In_712,In_789);
xnor U3676 (N_3676,In_881,In_1466);
or U3677 (N_3677,In_181,In_1303);
and U3678 (N_3678,In_282,In_289);
nand U3679 (N_3679,In_1310,In_1201);
or U3680 (N_3680,In_1206,In_1465);
nor U3681 (N_3681,In_927,In_574);
nand U3682 (N_3682,In_1098,In_495);
nor U3683 (N_3683,In_489,In_862);
nor U3684 (N_3684,In_702,In_177);
and U3685 (N_3685,In_336,In_1138);
nand U3686 (N_3686,In_117,In_884);
and U3687 (N_3687,In_1491,In_1105);
and U3688 (N_3688,In_143,In_992);
nand U3689 (N_3689,In_559,In_45);
or U3690 (N_3690,In_1089,In_606);
nand U3691 (N_3691,In_1381,In_790);
nor U3692 (N_3692,In_435,In_402);
and U3693 (N_3693,In_1371,In_1072);
or U3694 (N_3694,In_134,In_1339);
nor U3695 (N_3695,In_1318,In_1172);
or U3696 (N_3696,In_1069,In_1136);
or U3697 (N_3697,In_1282,In_82);
nor U3698 (N_3698,In_1039,In_252);
or U3699 (N_3699,In_738,In_576);
nand U3700 (N_3700,In_1117,In_593);
nor U3701 (N_3701,In_1296,In_926);
nor U3702 (N_3702,In_386,In_1435);
nor U3703 (N_3703,In_1084,In_399);
nor U3704 (N_3704,In_824,In_242);
nand U3705 (N_3705,In_820,In_54);
or U3706 (N_3706,In_855,In_980);
nand U3707 (N_3707,In_1277,In_1488);
or U3708 (N_3708,In_712,In_675);
nand U3709 (N_3709,In_353,In_1391);
nor U3710 (N_3710,In_133,In_498);
or U3711 (N_3711,In_991,In_1160);
nand U3712 (N_3712,In_425,In_875);
and U3713 (N_3713,In_480,In_989);
and U3714 (N_3714,In_333,In_1350);
nand U3715 (N_3715,In_1193,In_542);
or U3716 (N_3716,In_1150,In_459);
nor U3717 (N_3717,In_773,In_267);
nor U3718 (N_3718,In_1060,In_254);
nand U3719 (N_3719,In_847,In_919);
nand U3720 (N_3720,In_804,In_480);
nand U3721 (N_3721,In_346,In_420);
and U3722 (N_3722,In_500,In_1246);
nor U3723 (N_3723,In_1301,In_67);
and U3724 (N_3724,In_892,In_799);
nor U3725 (N_3725,In_957,In_1128);
nor U3726 (N_3726,In_406,In_712);
nand U3727 (N_3727,In_1084,In_1184);
xnor U3728 (N_3728,In_747,In_1023);
and U3729 (N_3729,In_134,In_799);
and U3730 (N_3730,In_1155,In_929);
nand U3731 (N_3731,In_1273,In_178);
nand U3732 (N_3732,In_368,In_387);
nor U3733 (N_3733,In_994,In_377);
nand U3734 (N_3734,In_1097,In_992);
or U3735 (N_3735,In_857,In_788);
and U3736 (N_3736,In_511,In_337);
nand U3737 (N_3737,In_478,In_600);
and U3738 (N_3738,In_1340,In_1324);
nand U3739 (N_3739,In_995,In_1182);
nand U3740 (N_3740,In_139,In_282);
or U3741 (N_3741,In_1240,In_468);
nor U3742 (N_3742,In_1162,In_390);
and U3743 (N_3743,In_42,In_1256);
or U3744 (N_3744,In_388,In_1425);
nand U3745 (N_3745,In_328,In_1247);
and U3746 (N_3746,In_932,In_1413);
nor U3747 (N_3747,In_1245,In_1175);
and U3748 (N_3748,In_825,In_881);
nor U3749 (N_3749,In_1156,In_924);
nor U3750 (N_3750,In_1354,In_138);
nand U3751 (N_3751,In_113,In_112);
or U3752 (N_3752,In_485,In_1180);
nand U3753 (N_3753,In_423,In_505);
or U3754 (N_3754,In_996,In_805);
nor U3755 (N_3755,In_517,In_609);
and U3756 (N_3756,In_30,In_1246);
or U3757 (N_3757,In_654,In_990);
nand U3758 (N_3758,In_30,In_789);
xor U3759 (N_3759,In_1127,In_261);
nand U3760 (N_3760,In_181,In_969);
nand U3761 (N_3761,In_1084,In_406);
xnor U3762 (N_3762,In_243,In_598);
and U3763 (N_3763,In_740,In_646);
and U3764 (N_3764,In_548,In_845);
nand U3765 (N_3765,In_1314,In_214);
nor U3766 (N_3766,In_849,In_110);
or U3767 (N_3767,In_621,In_1172);
nand U3768 (N_3768,In_1072,In_998);
nor U3769 (N_3769,In_502,In_555);
or U3770 (N_3770,In_448,In_957);
or U3771 (N_3771,In_624,In_595);
nand U3772 (N_3772,In_1495,In_998);
or U3773 (N_3773,In_58,In_341);
nand U3774 (N_3774,In_972,In_441);
nand U3775 (N_3775,In_1490,In_16);
nand U3776 (N_3776,In_401,In_714);
or U3777 (N_3777,In_1102,In_1219);
and U3778 (N_3778,In_155,In_1441);
and U3779 (N_3779,In_411,In_65);
nor U3780 (N_3780,In_832,In_300);
and U3781 (N_3781,In_741,In_1174);
nand U3782 (N_3782,In_43,In_349);
nand U3783 (N_3783,In_26,In_287);
nor U3784 (N_3784,In_998,In_562);
nor U3785 (N_3785,In_900,In_546);
and U3786 (N_3786,In_53,In_882);
or U3787 (N_3787,In_1353,In_182);
and U3788 (N_3788,In_253,In_24);
and U3789 (N_3789,In_1006,In_404);
nor U3790 (N_3790,In_63,In_140);
and U3791 (N_3791,In_918,In_922);
xnor U3792 (N_3792,In_1417,In_63);
nor U3793 (N_3793,In_119,In_1435);
and U3794 (N_3794,In_234,In_1019);
nor U3795 (N_3795,In_259,In_1040);
and U3796 (N_3796,In_1265,In_296);
nor U3797 (N_3797,In_507,In_313);
nor U3798 (N_3798,In_1389,In_1266);
nor U3799 (N_3799,In_576,In_1060);
nor U3800 (N_3800,In_592,In_995);
and U3801 (N_3801,In_331,In_875);
and U3802 (N_3802,In_1136,In_623);
and U3803 (N_3803,In_281,In_596);
nor U3804 (N_3804,In_443,In_1414);
or U3805 (N_3805,In_1350,In_765);
and U3806 (N_3806,In_1004,In_615);
nor U3807 (N_3807,In_366,In_895);
nand U3808 (N_3808,In_1361,In_1201);
and U3809 (N_3809,In_1074,In_1377);
nor U3810 (N_3810,In_122,In_180);
or U3811 (N_3811,In_419,In_694);
nor U3812 (N_3812,In_564,In_841);
and U3813 (N_3813,In_1364,In_882);
nand U3814 (N_3814,In_22,In_330);
nor U3815 (N_3815,In_1133,In_467);
or U3816 (N_3816,In_113,In_68);
or U3817 (N_3817,In_1156,In_1211);
and U3818 (N_3818,In_840,In_141);
nor U3819 (N_3819,In_1146,In_1012);
nor U3820 (N_3820,In_91,In_99);
nand U3821 (N_3821,In_347,In_844);
and U3822 (N_3822,In_1071,In_683);
or U3823 (N_3823,In_80,In_319);
nor U3824 (N_3824,In_90,In_691);
nor U3825 (N_3825,In_972,In_1360);
and U3826 (N_3826,In_1371,In_630);
or U3827 (N_3827,In_223,In_1174);
and U3828 (N_3828,In_561,In_1017);
and U3829 (N_3829,In_441,In_305);
or U3830 (N_3830,In_646,In_157);
nand U3831 (N_3831,In_189,In_588);
nand U3832 (N_3832,In_889,In_262);
nand U3833 (N_3833,In_1442,In_668);
nor U3834 (N_3834,In_537,In_577);
nor U3835 (N_3835,In_1466,In_19);
and U3836 (N_3836,In_1377,In_576);
nand U3837 (N_3837,In_1264,In_391);
nor U3838 (N_3838,In_568,In_1472);
or U3839 (N_3839,In_1081,In_563);
or U3840 (N_3840,In_1095,In_339);
and U3841 (N_3841,In_355,In_1072);
and U3842 (N_3842,In_322,In_1313);
and U3843 (N_3843,In_1196,In_1365);
and U3844 (N_3844,In_1192,In_1087);
and U3845 (N_3845,In_648,In_952);
nand U3846 (N_3846,In_429,In_85);
nor U3847 (N_3847,In_370,In_727);
or U3848 (N_3848,In_797,In_1454);
nand U3849 (N_3849,In_1098,In_636);
nor U3850 (N_3850,In_1380,In_1159);
or U3851 (N_3851,In_1212,In_99);
nor U3852 (N_3852,In_1440,In_1498);
nand U3853 (N_3853,In_726,In_979);
and U3854 (N_3854,In_1383,In_1452);
nand U3855 (N_3855,In_189,In_1139);
or U3856 (N_3856,In_971,In_966);
or U3857 (N_3857,In_1017,In_53);
nor U3858 (N_3858,In_1098,In_1203);
nand U3859 (N_3859,In_1297,In_1434);
xnor U3860 (N_3860,In_1280,In_922);
or U3861 (N_3861,In_1001,In_311);
nand U3862 (N_3862,In_1222,In_545);
or U3863 (N_3863,In_1010,In_95);
or U3864 (N_3864,In_246,In_113);
or U3865 (N_3865,In_1024,In_544);
xor U3866 (N_3866,In_1153,In_1300);
nor U3867 (N_3867,In_1428,In_1036);
and U3868 (N_3868,In_1068,In_659);
or U3869 (N_3869,In_338,In_720);
and U3870 (N_3870,In_1120,In_655);
nand U3871 (N_3871,In_888,In_315);
or U3872 (N_3872,In_708,In_561);
nand U3873 (N_3873,In_912,In_61);
nand U3874 (N_3874,In_1393,In_375);
nor U3875 (N_3875,In_450,In_1190);
nor U3876 (N_3876,In_931,In_445);
or U3877 (N_3877,In_56,In_961);
nor U3878 (N_3878,In_468,In_304);
nand U3879 (N_3879,In_1034,In_999);
nand U3880 (N_3880,In_1080,In_845);
nor U3881 (N_3881,In_483,In_637);
and U3882 (N_3882,In_30,In_108);
and U3883 (N_3883,In_896,In_438);
and U3884 (N_3884,In_368,In_94);
nand U3885 (N_3885,In_378,In_518);
or U3886 (N_3886,In_862,In_68);
and U3887 (N_3887,In_1139,In_852);
nand U3888 (N_3888,In_525,In_528);
nand U3889 (N_3889,In_914,In_746);
xor U3890 (N_3890,In_66,In_1339);
nand U3891 (N_3891,In_476,In_914);
and U3892 (N_3892,In_1099,In_1338);
nand U3893 (N_3893,In_661,In_1495);
or U3894 (N_3894,In_11,In_969);
and U3895 (N_3895,In_1019,In_1264);
or U3896 (N_3896,In_175,In_1241);
or U3897 (N_3897,In_1310,In_1282);
nand U3898 (N_3898,In_1022,In_1412);
xor U3899 (N_3899,In_1298,In_624);
or U3900 (N_3900,In_1386,In_1410);
nor U3901 (N_3901,In_1238,In_90);
nand U3902 (N_3902,In_1303,In_342);
nand U3903 (N_3903,In_257,In_894);
or U3904 (N_3904,In_563,In_998);
nand U3905 (N_3905,In_681,In_1230);
nand U3906 (N_3906,In_486,In_613);
nor U3907 (N_3907,In_747,In_1477);
or U3908 (N_3908,In_1391,In_388);
nand U3909 (N_3909,In_449,In_40);
and U3910 (N_3910,In_177,In_600);
nor U3911 (N_3911,In_1249,In_1285);
and U3912 (N_3912,In_550,In_1235);
nor U3913 (N_3913,In_1014,In_617);
and U3914 (N_3914,In_334,In_845);
nor U3915 (N_3915,In_135,In_111);
or U3916 (N_3916,In_708,In_949);
nand U3917 (N_3917,In_448,In_1373);
nand U3918 (N_3918,In_412,In_1302);
nor U3919 (N_3919,In_784,In_259);
or U3920 (N_3920,In_620,In_254);
and U3921 (N_3921,In_1376,In_1206);
or U3922 (N_3922,In_386,In_56);
nor U3923 (N_3923,In_1155,In_68);
and U3924 (N_3924,In_1005,In_1296);
nand U3925 (N_3925,In_380,In_331);
and U3926 (N_3926,In_216,In_1495);
nand U3927 (N_3927,In_395,In_1177);
or U3928 (N_3928,In_1203,In_1250);
nand U3929 (N_3929,In_889,In_1130);
or U3930 (N_3930,In_248,In_1431);
xnor U3931 (N_3931,In_1314,In_104);
or U3932 (N_3932,In_6,In_443);
nand U3933 (N_3933,In_321,In_442);
xnor U3934 (N_3934,In_437,In_300);
and U3935 (N_3935,In_1126,In_942);
nand U3936 (N_3936,In_556,In_827);
nor U3937 (N_3937,In_682,In_331);
nand U3938 (N_3938,In_279,In_929);
and U3939 (N_3939,In_524,In_1065);
or U3940 (N_3940,In_528,In_1413);
nand U3941 (N_3941,In_1382,In_43);
or U3942 (N_3942,In_54,In_1317);
or U3943 (N_3943,In_1080,In_101);
nand U3944 (N_3944,In_1011,In_520);
nor U3945 (N_3945,In_1041,In_126);
nand U3946 (N_3946,In_1138,In_473);
nor U3947 (N_3947,In_1247,In_1296);
and U3948 (N_3948,In_151,In_46);
nand U3949 (N_3949,In_578,In_1476);
nand U3950 (N_3950,In_572,In_1199);
nor U3951 (N_3951,In_677,In_336);
nand U3952 (N_3952,In_527,In_799);
xnor U3953 (N_3953,In_325,In_577);
and U3954 (N_3954,In_395,In_508);
or U3955 (N_3955,In_179,In_771);
and U3956 (N_3956,In_377,In_422);
nand U3957 (N_3957,In_1059,In_161);
or U3958 (N_3958,In_757,In_1295);
and U3959 (N_3959,In_105,In_1074);
nor U3960 (N_3960,In_1103,In_1321);
or U3961 (N_3961,In_1291,In_781);
and U3962 (N_3962,In_178,In_1376);
nor U3963 (N_3963,In_809,In_1282);
and U3964 (N_3964,In_130,In_977);
or U3965 (N_3965,In_956,In_528);
xnor U3966 (N_3966,In_782,In_139);
nor U3967 (N_3967,In_468,In_788);
nand U3968 (N_3968,In_1051,In_1268);
nor U3969 (N_3969,In_242,In_1113);
or U3970 (N_3970,In_689,In_104);
or U3971 (N_3971,In_949,In_262);
and U3972 (N_3972,In_815,In_386);
nand U3973 (N_3973,In_1109,In_1141);
or U3974 (N_3974,In_527,In_640);
or U3975 (N_3975,In_588,In_583);
xnor U3976 (N_3976,In_687,In_33);
nor U3977 (N_3977,In_295,In_1132);
nor U3978 (N_3978,In_626,In_496);
and U3979 (N_3979,In_747,In_217);
xor U3980 (N_3980,In_256,In_312);
and U3981 (N_3981,In_539,In_747);
and U3982 (N_3982,In_1360,In_64);
and U3983 (N_3983,In_163,In_1146);
nor U3984 (N_3984,In_1171,In_311);
nand U3985 (N_3985,In_215,In_489);
xor U3986 (N_3986,In_1493,In_1022);
nor U3987 (N_3987,In_54,In_1453);
or U3988 (N_3988,In_437,In_612);
or U3989 (N_3989,In_1202,In_184);
nand U3990 (N_3990,In_1482,In_1412);
nor U3991 (N_3991,In_551,In_191);
nand U3992 (N_3992,In_195,In_704);
nand U3993 (N_3993,In_945,In_1214);
and U3994 (N_3994,In_873,In_1340);
or U3995 (N_3995,In_875,In_386);
and U3996 (N_3996,In_1158,In_325);
or U3997 (N_3997,In_14,In_406);
nor U3998 (N_3998,In_635,In_162);
nor U3999 (N_3999,In_1299,In_1011);
or U4000 (N_4000,In_591,In_204);
or U4001 (N_4001,In_609,In_78);
nor U4002 (N_4002,In_1088,In_455);
nand U4003 (N_4003,In_118,In_1311);
or U4004 (N_4004,In_665,In_996);
nor U4005 (N_4005,In_745,In_898);
and U4006 (N_4006,In_633,In_400);
xor U4007 (N_4007,In_354,In_317);
nor U4008 (N_4008,In_1087,In_712);
or U4009 (N_4009,In_200,In_730);
nand U4010 (N_4010,In_1248,In_1468);
nand U4011 (N_4011,In_313,In_231);
xnor U4012 (N_4012,In_1094,In_945);
or U4013 (N_4013,In_356,In_858);
xor U4014 (N_4014,In_231,In_1226);
nand U4015 (N_4015,In_414,In_633);
nor U4016 (N_4016,In_207,In_477);
nand U4017 (N_4017,In_958,In_1344);
and U4018 (N_4018,In_1113,In_263);
or U4019 (N_4019,In_78,In_191);
nor U4020 (N_4020,In_262,In_335);
or U4021 (N_4021,In_439,In_1457);
nor U4022 (N_4022,In_622,In_1241);
or U4023 (N_4023,In_451,In_821);
or U4024 (N_4024,In_663,In_661);
and U4025 (N_4025,In_1193,In_204);
nand U4026 (N_4026,In_461,In_675);
and U4027 (N_4027,In_535,In_665);
or U4028 (N_4028,In_588,In_416);
and U4029 (N_4029,In_391,In_754);
and U4030 (N_4030,In_478,In_920);
nor U4031 (N_4031,In_360,In_400);
nand U4032 (N_4032,In_426,In_382);
and U4033 (N_4033,In_1101,In_973);
nand U4034 (N_4034,In_947,In_271);
and U4035 (N_4035,In_1192,In_576);
nor U4036 (N_4036,In_661,In_838);
nand U4037 (N_4037,In_1129,In_59);
and U4038 (N_4038,In_204,In_140);
nor U4039 (N_4039,In_1029,In_240);
or U4040 (N_4040,In_1294,In_459);
nor U4041 (N_4041,In_391,In_952);
nor U4042 (N_4042,In_1187,In_376);
nor U4043 (N_4043,In_573,In_358);
or U4044 (N_4044,In_766,In_47);
nand U4045 (N_4045,In_914,In_455);
nor U4046 (N_4046,In_350,In_1468);
and U4047 (N_4047,In_1060,In_255);
nand U4048 (N_4048,In_292,In_280);
or U4049 (N_4049,In_61,In_1384);
and U4050 (N_4050,In_91,In_1237);
or U4051 (N_4051,In_292,In_75);
or U4052 (N_4052,In_1449,In_1463);
nor U4053 (N_4053,In_1469,In_1237);
nand U4054 (N_4054,In_815,In_453);
and U4055 (N_4055,In_1410,In_244);
nor U4056 (N_4056,In_168,In_614);
or U4057 (N_4057,In_1113,In_336);
nor U4058 (N_4058,In_774,In_127);
and U4059 (N_4059,In_856,In_959);
nor U4060 (N_4060,In_1180,In_352);
nor U4061 (N_4061,In_1087,In_432);
and U4062 (N_4062,In_558,In_1147);
nand U4063 (N_4063,In_988,In_835);
nand U4064 (N_4064,In_1475,In_327);
or U4065 (N_4065,In_1467,In_1239);
and U4066 (N_4066,In_1473,In_189);
nor U4067 (N_4067,In_464,In_951);
or U4068 (N_4068,In_204,In_575);
nand U4069 (N_4069,In_582,In_271);
nor U4070 (N_4070,In_23,In_740);
nand U4071 (N_4071,In_603,In_740);
nand U4072 (N_4072,In_177,In_1285);
and U4073 (N_4073,In_954,In_1076);
nand U4074 (N_4074,In_633,In_506);
and U4075 (N_4075,In_233,In_653);
and U4076 (N_4076,In_415,In_250);
and U4077 (N_4077,In_1207,In_688);
nor U4078 (N_4078,In_459,In_902);
nor U4079 (N_4079,In_3,In_1357);
or U4080 (N_4080,In_514,In_695);
xnor U4081 (N_4081,In_24,In_617);
or U4082 (N_4082,In_963,In_1432);
nor U4083 (N_4083,In_583,In_319);
nand U4084 (N_4084,In_490,In_1275);
nand U4085 (N_4085,In_884,In_1178);
or U4086 (N_4086,In_635,In_1074);
and U4087 (N_4087,In_379,In_1392);
or U4088 (N_4088,In_542,In_1149);
or U4089 (N_4089,In_203,In_980);
or U4090 (N_4090,In_1032,In_1077);
nor U4091 (N_4091,In_290,In_274);
or U4092 (N_4092,In_956,In_1057);
and U4093 (N_4093,In_928,In_1310);
or U4094 (N_4094,In_302,In_115);
and U4095 (N_4095,In_254,In_60);
and U4096 (N_4096,In_841,In_984);
and U4097 (N_4097,In_260,In_1109);
nor U4098 (N_4098,In_1441,In_952);
or U4099 (N_4099,In_471,In_58);
or U4100 (N_4100,In_1259,In_1448);
nor U4101 (N_4101,In_232,In_993);
nand U4102 (N_4102,In_833,In_800);
or U4103 (N_4103,In_1370,In_1409);
nor U4104 (N_4104,In_372,In_627);
nand U4105 (N_4105,In_1223,In_1276);
or U4106 (N_4106,In_1131,In_754);
and U4107 (N_4107,In_183,In_97);
and U4108 (N_4108,In_1452,In_31);
nand U4109 (N_4109,In_106,In_735);
nor U4110 (N_4110,In_261,In_925);
and U4111 (N_4111,In_1296,In_90);
or U4112 (N_4112,In_539,In_478);
nor U4113 (N_4113,In_294,In_341);
and U4114 (N_4114,In_780,In_347);
nor U4115 (N_4115,In_230,In_372);
nor U4116 (N_4116,In_281,In_1103);
and U4117 (N_4117,In_83,In_785);
nor U4118 (N_4118,In_590,In_1349);
and U4119 (N_4119,In_582,In_990);
or U4120 (N_4120,In_1150,In_1442);
nand U4121 (N_4121,In_1084,In_1243);
and U4122 (N_4122,In_471,In_985);
or U4123 (N_4123,In_439,In_352);
nand U4124 (N_4124,In_670,In_179);
and U4125 (N_4125,In_184,In_1011);
and U4126 (N_4126,In_156,In_815);
nand U4127 (N_4127,In_931,In_600);
nand U4128 (N_4128,In_662,In_1121);
or U4129 (N_4129,In_1239,In_320);
nor U4130 (N_4130,In_966,In_544);
or U4131 (N_4131,In_586,In_807);
nand U4132 (N_4132,In_1476,In_1125);
and U4133 (N_4133,In_1398,In_1497);
or U4134 (N_4134,In_121,In_1181);
or U4135 (N_4135,In_662,In_911);
and U4136 (N_4136,In_145,In_938);
and U4137 (N_4137,In_955,In_279);
nor U4138 (N_4138,In_1399,In_1120);
nand U4139 (N_4139,In_93,In_539);
nand U4140 (N_4140,In_1319,In_388);
nand U4141 (N_4141,In_81,In_1157);
and U4142 (N_4142,In_889,In_404);
or U4143 (N_4143,In_968,In_1403);
nand U4144 (N_4144,In_1157,In_966);
nor U4145 (N_4145,In_968,In_554);
or U4146 (N_4146,In_704,In_507);
nand U4147 (N_4147,In_140,In_1137);
xor U4148 (N_4148,In_1444,In_1267);
and U4149 (N_4149,In_1026,In_1210);
nor U4150 (N_4150,In_880,In_957);
or U4151 (N_4151,In_813,In_1094);
nor U4152 (N_4152,In_1417,In_1001);
nand U4153 (N_4153,In_259,In_655);
or U4154 (N_4154,In_306,In_1295);
and U4155 (N_4155,In_97,In_441);
nand U4156 (N_4156,In_1161,In_1219);
nand U4157 (N_4157,In_358,In_902);
or U4158 (N_4158,In_1460,In_1326);
nor U4159 (N_4159,In_1145,In_392);
nor U4160 (N_4160,In_984,In_1146);
nand U4161 (N_4161,In_248,In_1176);
or U4162 (N_4162,In_211,In_727);
and U4163 (N_4163,In_331,In_626);
or U4164 (N_4164,In_420,In_902);
nand U4165 (N_4165,In_1031,In_1053);
and U4166 (N_4166,In_700,In_236);
nand U4167 (N_4167,In_1345,In_896);
nand U4168 (N_4168,In_1242,In_1394);
and U4169 (N_4169,In_161,In_1178);
nand U4170 (N_4170,In_1317,In_130);
nand U4171 (N_4171,In_49,In_52);
or U4172 (N_4172,In_476,In_657);
nor U4173 (N_4173,In_77,In_1442);
and U4174 (N_4174,In_852,In_400);
and U4175 (N_4175,In_551,In_345);
or U4176 (N_4176,In_294,In_1407);
or U4177 (N_4177,In_27,In_868);
nor U4178 (N_4178,In_920,In_1003);
nand U4179 (N_4179,In_1241,In_1089);
or U4180 (N_4180,In_785,In_885);
and U4181 (N_4181,In_1446,In_629);
or U4182 (N_4182,In_648,In_738);
or U4183 (N_4183,In_728,In_753);
and U4184 (N_4184,In_1266,In_1245);
or U4185 (N_4185,In_1452,In_552);
or U4186 (N_4186,In_304,In_361);
nand U4187 (N_4187,In_1149,In_258);
and U4188 (N_4188,In_1000,In_1047);
xor U4189 (N_4189,In_1198,In_393);
and U4190 (N_4190,In_1046,In_1242);
nand U4191 (N_4191,In_1049,In_1113);
or U4192 (N_4192,In_259,In_86);
xor U4193 (N_4193,In_356,In_48);
xnor U4194 (N_4194,In_863,In_850);
xor U4195 (N_4195,In_177,In_1122);
or U4196 (N_4196,In_1065,In_1211);
or U4197 (N_4197,In_1130,In_47);
nor U4198 (N_4198,In_803,In_1435);
or U4199 (N_4199,In_905,In_1047);
or U4200 (N_4200,In_701,In_1079);
nor U4201 (N_4201,In_845,In_648);
nand U4202 (N_4202,In_387,In_1370);
nand U4203 (N_4203,In_1095,In_1348);
or U4204 (N_4204,In_955,In_1304);
nor U4205 (N_4205,In_659,In_294);
nand U4206 (N_4206,In_720,In_631);
nand U4207 (N_4207,In_381,In_54);
nor U4208 (N_4208,In_232,In_970);
nand U4209 (N_4209,In_137,In_1025);
or U4210 (N_4210,In_1194,In_582);
nand U4211 (N_4211,In_535,In_460);
and U4212 (N_4212,In_1257,In_809);
nor U4213 (N_4213,In_1497,In_650);
or U4214 (N_4214,In_1116,In_840);
nand U4215 (N_4215,In_566,In_79);
or U4216 (N_4216,In_118,In_197);
nor U4217 (N_4217,In_1017,In_870);
and U4218 (N_4218,In_427,In_724);
nor U4219 (N_4219,In_822,In_1469);
or U4220 (N_4220,In_1380,In_751);
and U4221 (N_4221,In_287,In_575);
nand U4222 (N_4222,In_1215,In_231);
nand U4223 (N_4223,In_693,In_1404);
or U4224 (N_4224,In_110,In_842);
or U4225 (N_4225,In_750,In_1211);
and U4226 (N_4226,In_1139,In_154);
nor U4227 (N_4227,In_1236,In_682);
and U4228 (N_4228,In_1016,In_1380);
nand U4229 (N_4229,In_893,In_996);
and U4230 (N_4230,In_545,In_1171);
nor U4231 (N_4231,In_681,In_520);
and U4232 (N_4232,In_338,In_1197);
and U4233 (N_4233,In_644,In_489);
nor U4234 (N_4234,In_534,In_908);
or U4235 (N_4235,In_313,In_107);
nor U4236 (N_4236,In_914,In_629);
xnor U4237 (N_4237,In_1182,In_50);
nor U4238 (N_4238,In_756,In_187);
or U4239 (N_4239,In_265,In_609);
or U4240 (N_4240,In_780,In_864);
or U4241 (N_4241,In_954,In_411);
and U4242 (N_4242,In_414,In_1175);
nand U4243 (N_4243,In_1393,In_1101);
nor U4244 (N_4244,In_218,In_400);
or U4245 (N_4245,In_1236,In_1316);
or U4246 (N_4246,In_389,In_925);
nand U4247 (N_4247,In_1048,In_1383);
nor U4248 (N_4248,In_143,In_387);
nor U4249 (N_4249,In_1337,In_1309);
or U4250 (N_4250,In_501,In_337);
and U4251 (N_4251,In_755,In_864);
or U4252 (N_4252,In_1239,In_448);
and U4253 (N_4253,In_1115,In_1294);
and U4254 (N_4254,In_87,In_882);
and U4255 (N_4255,In_1449,In_933);
nand U4256 (N_4256,In_1167,In_1294);
nor U4257 (N_4257,In_241,In_1135);
or U4258 (N_4258,In_1494,In_881);
or U4259 (N_4259,In_1194,In_1299);
or U4260 (N_4260,In_626,In_800);
nor U4261 (N_4261,In_343,In_237);
nor U4262 (N_4262,In_693,In_1305);
and U4263 (N_4263,In_464,In_424);
or U4264 (N_4264,In_417,In_304);
nand U4265 (N_4265,In_1298,In_113);
or U4266 (N_4266,In_431,In_463);
nor U4267 (N_4267,In_129,In_24);
nor U4268 (N_4268,In_448,In_1497);
or U4269 (N_4269,In_1173,In_696);
nand U4270 (N_4270,In_825,In_566);
or U4271 (N_4271,In_183,In_398);
nand U4272 (N_4272,In_197,In_534);
and U4273 (N_4273,In_1228,In_409);
and U4274 (N_4274,In_1423,In_1481);
or U4275 (N_4275,In_1433,In_1342);
and U4276 (N_4276,In_994,In_22);
xnor U4277 (N_4277,In_552,In_1077);
nand U4278 (N_4278,In_452,In_1459);
or U4279 (N_4279,In_780,In_75);
or U4280 (N_4280,In_569,In_252);
nand U4281 (N_4281,In_636,In_301);
nand U4282 (N_4282,In_1417,In_1467);
and U4283 (N_4283,In_639,In_1478);
and U4284 (N_4284,In_1081,In_458);
or U4285 (N_4285,In_1224,In_1143);
nor U4286 (N_4286,In_1054,In_144);
or U4287 (N_4287,In_970,In_367);
and U4288 (N_4288,In_1077,In_1153);
and U4289 (N_4289,In_1114,In_1416);
xor U4290 (N_4290,In_440,In_1116);
and U4291 (N_4291,In_972,In_1166);
nor U4292 (N_4292,In_47,In_963);
nand U4293 (N_4293,In_689,In_634);
or U4294 (N_4294,In_148,In_673);
nor U4295 (N_4295,In_1471,In_1013);
nor U4296 (N_4296,In_1335,In_1416);
nand U4297 (N_4297,In_538,In_499);
nand U4298 (N_4298,In_916,In_1113);
nand U4299 (N_4299,In_652,In_1079);
or U4300 (N_4300,In_572,In_1271);
nor U4301 (N_4301,In_549,In_700);
or U4302 (N_4302,In_847,In_1161);
nand U4303 (N_4303,In_279,In_850);
nor U4304 (N_4304,In_679,In_845);
and U4305 (N_4305,In_1169,In_431);
nand U4306 (N_4306,In_231,In_1072);
nand U4307 (N_4307,In_171,In_115);
and U4308 (N_4308,In_445,In_200);
nand U4309 (N_4309,In_1076,In_825);
and U4310 (N_4310,In_532,In_398);
nand U4311 (N_4311,In_1206,In_1076);
xor U4312 (N_4312,In_409,In_920);
or U4313 (N_4313,In_1499,In_642);
nand U4314 (N_4314,In_747,In_470);
nand U4315 (N_4315,In_369,In_296);
or U4316 (N_4316,In_129,In_338);
nor U4317 (N_4317,In_704,In_837);
or U4318 (N_4318,In_1126,In_908);
nor U4319 (N_4319,In_834,In_117);
nand U4320 (N_4320,In_1140,In_1138);
nand U4321 (N_4321,In_981,In_828);
nor U4322 (N_4322,In_1012,In_323);
nand U4323 (N_4323,In_1331,In_1285);
or U4324 (N_4324,In_878,In_610);
and U4325 (N_4325,In_932,In_304);
nor U4326 (N_4326,In_142,In_1425);
and U4327 (N_4327,In_1019,In_1466);
nand U4328 (N_4328,In_104,In_160);
and U4329 (N_4329,In_777,In_1093);
xnor U4330 (N_4330,In_1330,In_790);
or U4331 (N_4331,In_1083,In_1262);
nor U4332 (N_4332,In_204,In_1070);
nand U4333 (N_4333,In_755,In_314);
nand U4334 (N_4334,In_1104,In_985);
nand U4335 (N_4335,In_197,In_765);
and U4336 (N_4336,In_27,In_328);
and U4337 (N_4337,In_1415,In_207);
xnor U4338 (N_4338,In_1106,In_703);
and U4339 (N_4339,In_490,In_480);
and U4340 (N_4340,In_930,In_84);
nor U4341 (N_4341,In_499,In_63);
and U4342 (N_4342,In_1349,In_572);
or U4343 (N_4343,In_888,In_641);
or U4344 (N_4344,In_531,In_930);
nand U4345 (N_4345,In_1265,In_1300);
and U4346 (N_4346,In_1379,In_446);
or U4347 (N_4347,In_619,In_958);
xor U4348 (N_4348,In_516,In_1249);
nor U4349 (N_4349,In_519,In_142);
and U4350 (N_4350,In_257,In_127);
nor U4351 (N_4351,In_547,In_21);
or U4352 (N_4352,In_1352,In_851);
nand U4353 (N_4353,In_956,In_766);
nor U4354 (N_4354,In_1176,In_149);
nor U4355 (N_4355,In_71,In_666);
nand U4356 (N_4356,In_469,In_1071);
or U4357 (N_4357,In_374,In_1435);
and U4358 (N_4358,In_1020,In_771);
or U4359 (N_4359,In_577,In_269);
or U4360 (N_4360,In_1068,In_567);
nand U4361 (N_4361,In_835,In_1373);
xor U4362 (N_4362,In_641,In_800);
and U4363 (N_4363,In_1388,In_1095);
nand U4364 (N_4364,In_1213,In_122);
nor U4365 (N_4365,In_105,In_315);
or U4366 (N_4366,In_605,In_1484);
nor U4367 (N_4367,In_1391,In_630);
nor U4368 (N_4368,In_1212,In_100);
and U4369 (N_4369,In_975,In_823);
nor U4370 (N_4370,In_985,In_712);
nand U4371 (N_4371,In_1210,In_899);
and U4372 (N_4372,In_1434,In_541);
and U4373 (N_4373,In_1266,In_1277);
xor U4374 (N_4374,In_694,In_1337);
and U4375 (N_4375,In_176,In_1377);
nor U4376 (N_4376,In_983,In_1072);
and U4377 (N_4377,In_998,In_312);
or U4378 (N_4378,In_491,In_510);
or U4379 (N_4379,In_766,In_1181);
nor U4380 (N_4380,In_1101,In_370);
nor U4381 (N_4381,In_854,In_266);
nor U4382 (N_4382,In_1373,In_1094);
and U4383 (N_4383,In_1459,In_1181);
nor U4384 (N_4384,In_1387,In_615);
nand U4385 (N_4385,In_949,In_1144);
nor U4386 (N_4386,In_1183,In_968);
and U4387 (N_4387,In_1048,In_1423);
and U4388 (N_4388,In_1379,In_147);
and U4389 (N_4389,In_964,In_1110);
or U4390 (N_4390,In_282,In_158);
xor U4391 (N_4391,In_26,In_636);
and U4392 (N_4392,In_1360,In_290);
nor U4393 (N_4393,In_352,In_511);
and U4394 (N_4394,In_235,In_1349);
and U4395 (N_4395,In_1019,In_530);
nor U4396 (N_4396,In_1468,In_1194);
nor U4397 (N_4397,In_1257,In_881);
and U4398 (N_4398,In_1488,In_134);
nor U4399 (N_4399,In_1311,In_531);
nand U4400 (N_4400,In_393,In_248);
nand U4401 (N_4401,In_769,In_1288);
nand U4402 (N_4402,In_1300,In_1251);
nand U4403 (N_4403,In_1397,In_568);
or U4404 (N_4404,In_340,In_505);
nand U4405 (N_4405,In_1076,In_936);
and U4406 (N_4406,In_429,In_1384);
xnor U4407 (N_4407,In_1383,In_220);
or U4408 (N_4408,In_246,In_960);
and U4409 (N_4409,In_755,In_908);
and U4410 (N_4410,In_36,In_740);
nor U4411 (N_4411,In_124,In_624);
nand U4412 (N_4412,In_372,In_841);
nor U4413 (N_4413,In_226,In_525);
nor U4414 (N_4414,In_1328,In_624);
nand U4415 (N_4415,In_786,In_1063);
nand U4416 (N_4416,In_62,In_1418);
nor U4417 (N_4417,In_292,In_527);
nor U4418 (N_4418,In_210,In_5);
and U4419 (N_4419,In_316,In_251);
or U4420 (N_4420,In_384,In_635);
or U4421 (N_4421,In_413,In_1152);
nor U4422 (N_4422,In_816,In_387);
or U4423 (N_4423,In_642,In_423);
nand U4424 (N_4424,In_73,In_1077);
and U4425 (N_4425,In_283,In_585);
nand U4426 (N_4426,In_38,In_990);
nand U4427 (N_4427,In_332,In_990);
or U4428 (N_4428,In_1389,In_1130);
nor U4429 (N_4429,In_1476,In_820);
nand U4430 (N_4430,In_599,In_232);
nor U4431 (N_4431,In_1376,In_755);
nor U4432 (N_4432,In_244,In_215);
nor U4433 (N_4433,In_916,In_1197);
nor U4434 (N_4434,In_223,In_204);
and U4435 (N_4435,In_420,In_1363);
or U4436 (N_4436,In_423,In_1475);
nand U4437 (N_4437,In_395,In_255);
nor U4438 (N_4438,In_1069,In_310);
nand U4439 (N_4439,In_6,In_80);
xnor U4440 (N_4440,In_568,In_776);
or U4441 (N_4441,In_228,In_122);
or U4442 (N_4442,In_387,In_1183);
xor U4443 (N_4443,In_1415,In_910);
nor U4444 (N_4444,In_1088,In_395);
and U4445 (N_4445,In_927,In_500);
nor U4446 (N_4446,In_903,In_30);
or U4447 (N_4447,In_580,In_829);
or U4448 (N_4448,In_546,In_1119);
nor U4449 (N_4449,In_853,In_73);
nand U4450 (N_4450,In_913,In_1318);
nand U4451 (N_4451,In_36,In_1029);
or U4452 (N_4452,In_1304,In_45);
and U4453 (N_4453,In_830,In_1201);
and U4454 (N_4454,In_257,In_693);
and U4455 (N_4455,In_15,In_179);
nand U4456 (N_4456,In_36,In_739);
and U4457 (N_4457,In_1449,In_1249);
or U4458 (N_4458,In_175,In_843);
xor U4459 (N_4459,In_934,In_382);
nor U4460 (N_4460,In_1455,In_617);
nor U4461 (N_4461,In_759,In_1243);
nor U4462 (N_4462,In_222,In_277);
nand U4463 (N_4463,In_452,In_1264);
nor U4464 (N_4464,In_1014,In_111);
and U4465 (N_4465,In_129,In_959);
nand U4466 (N_4466,In_621,In_1284);
xnor U4467 (N_4467,In_1297,In_242);
nor U4468 (N_4468,In_1338,In_119);
or U4469 (N_4469,In_22,In_968);
nand U4470 (N_4470,In_480,In_822);
or U4471 (N_4471,In_711,In_1397);
nor U4472 (N_4472,In_388,In_940);
nor U4473 (N_4473,In_420,In_706);
nand U4474 (N_4474,In_380,In_1140);
nand U4475 (N_4475,In_115,In_1187);
nor U4476 (N_4476,In_820,In_345);
nor U4477 (N_4477,In_690,In_862);
and U4478 (N_4478,In_216,In_238);
nand U4479 (N_4479,In_257,In_1084);
nand U4480 (N_4480,In_1132,In_1126);
and U4481 (N_4481,In_290,In_1002);
and U4482 (N_4482,In_1481,In_1305);
and U4483 (N_4483,In_768,In_798);
nor U4484 (N_4484,In_1021,In_1253);
nand U4485 (N_4485,In_114,In_1209);
or U4486 (N_4486,In_1198,In_977);
nor U4487 (N_4487,In_102,In_377);
or U4488 (N_4488,In_1410,In_454);
nor U4489 (N_4489,In_1402,In_692);
nand U4490 (N_4490,In_804,In_1363);
nor U4491 (N_4491,In_1234,In_372);
nor U4492 (N_4492,In_1424,In_1290);
nand U4493 (N_4493,In_791,In_450);
nor U4494 (N_4494,In_430,In_416);
nor U4495 (N_4495,In_501,In_1057);
or U4496 (N_4496,In_1371,In_995);
or U4497 (N_4497,In_130,In_284);
and U4498 (N_4498,In_179,In_1151);
or U4499 (N_4499,In_812,In_19);
nand U4500 (N_4500,In_216,In_211);
xor U4501 (N_4501,In_458,In_135);
and U4502 (N_4502,In_1084,In_1314);
or U4503 (N_4503,In_165,In_1450);
nand U4504 (N_4504,In_55,In_419);
nor U4505 (N_4505,In_900,In_1277);
or U4506 (N_4506,In_1420,In_1329);
and U4507 (N_4507,In_1496,In_1481);
nor U4508 (N_4508,In_727,In_1279);
or U4509 (N_4509,In_791,In_460);
or U4510 (N_4510,In_394,In_1370);
nand U4511 (N_4511,In_1257,In_879);
nor U4512 (N_4512,In_490,In_590);
nand U4513 (N_4513,In_249,In_551);
or U4514 (N_4514,In_372,In_839);
nor U4515 (N_4515,In_1368,In_346);
or U4516 (N_4516,In_777,In_394);
or U4517 (N_4517,In_998,In_169);
and U4518 (N_4518,In_370,In_1125);
nand U4519 (N_4519,In_1495,In_199);
and U4520 (N_4520,In_491,In_1024);
xnor U4521 (N_4521,In_1017,In_405);
or U4522 (N_4522,In_253,In_576);
or U4523 (N_4523,In_1440,In_511);
and U4524 (N_4524,In_895,In_1286);
nor U4525 (N_4525,In_355,In_1383);
and U4526 (N_4526,In_285,In_633);
nor U4527 (N_4527,In_423,In_640);
nor U4528 (N_4528,In_1436,In_997);
and U4529 (N_4529,In_151,In_385);
nor U4530 (N_4530,In_890,In_1325);
nand U4531 (N_4531,In_100,In_1260);
nor U4532 (N_4532,In_445,In_543);
and U4533 (N_4533,In_985,In_236);
nand U4534 (N_4534,In_797,In_1108);
or U4535 (N_4535,In_123,In_814);
or U4536 (N_4536,In_1062,In_202);
and U4537 (N_4537,In_477,In_828);
nand U4538 (N_4538,In_374,In_923);
nor U4539 (N_4539,In_1376,In_485);
or U4540 (N_4540,In_137,In_1071);
nor U4541 (N_4541,In_1439,In_1453);
nor U4542 (N_4542,In_895,In_467);
nand U4543 (N_4543,In_1471,In_72);
and U4544 (N_4544,In_310,In_430);
nor U4545 (N_4545,In_659,In_1337);
or U4546 (N_4546,In_27,In_1379);
nand U4547 (N_4547,In_71,In_602);
nor U4548 (N_4548,In_1366,In_194);
and U4549 (N_4549,In_750,In_1151);
or U4550 (N_4550,In_972,In_1459);
or U4551 (N_4551,In_463,In_739);
and U4552 (N_4552,In_33,In_541);
nor U4553 (N_4553,In_567,In_1042);
nand U4554 (N_4554,In_958,In_947);
and U4555 (N_4555,In_275,In_1255);
nor U4556 (N_4556,In_1385,In_814);
or U4557 (N_4557,In_1126,In_830);
and U4558 (N_4558,In_1254,In_961);
nor U4559 (N_4559,In_1251,In_1332);
nand U4560 (N_4560,In_708,In_1022);
and U4561 (N_4561,In_90,In_667);
or U4562 (N_4562,In_373,In_736);
or U4563 (N_4563,In_56,In_1329);
nor U4564 (N_4564,In_1232,In_990);
and U4565 (N_4565,In_1492,In_1362);
or U4566 (N_4566,In_315,In_965);
nor U4567 (N_4567,In_1175,In_1045);
nand U4568 (N_4568,In_574,In_866);
or U4569 (N_4569,In_925,In_1411);
or U4570 (N_4570,In_495,In_1192);
nand U4571 (N_4571,In_377,In_216);
nor U4572 (N_4572,In_133,In_1441);
nor U4573 (N_4573,In_232,In_173);
nor U4574 (N_4574,In_1083,In_673);
or U4575 (N_4575,In_169,In_1362);
and U4576 (N_4576,In_1044,In_71);
and U4577 (N_4577,In_92,In_1459);
or U4578 (N_4578,In_672,In_919);
or U4579 (N_4579,In_821,In_45);
nand U4580 (N_4580,In_629,In_421);
or U4581 (N_4581,In_35,In_95);
nor U4582 (N_4582,In_319,In_1357);
nand U4583 (N_4583,In_66,In_430);
and U4584 (N_4584,In_984,In_19);
and U4585 (N_4585,In_768,In_674);
nand U4586 (N_4586,In_1433,In_628);
nand U4587 (N_4587,In_7,In_3);
or U4588 (N_4588,In_244,In_339);
xnor U4589 (N_4589,In_1412,In_896);
nor U4590 (N_4590,In_1092,In_938);
or U4591 (N_4591,In_1471,In_950);
and U4592 (N_4592,In_1067,In_962);
or U4593 (N_4593,In_444,In_1375);
or U4594 (N_4594,In_1472,In_1200);
or U4595 (N_4595,In_1022,In_328);
nor U4596 (N_4596,In_379,In_359);
nor U4597 (N_4597,In_637,In_1495);
or U4598 (N_4598,In_161,In_1126);
and U4599 (N_4599,In_618,In_844);
nor U4600 (N_4600,In_251,In_1282);
or U4601 (N_4601,In_353,In_54);
nand U4602 (N_4602,In_78,In_312);
xnor U4603 (N_4603,In_750,In_864);
nand U4604 (N_4604,In_1041,In_1481);
nand U4605 (N_4605,In_1411,In_1290);
and U4606 (N_4606,In_731,In_86);
nand U4607 (N_4607,In_193,In_638);
or U4608 (N_4608,In_296,In_1203);
and U4609 (N_4609,In_1312,In_592);
nand U4610 (N_4610,In_1271,In_1022);
and U4611 (N_4611,In_1016,In_526);
and U4612 (N_4612,In_8,In_666);
nor U4613 (N_4613,In_316,In_228);
or U4614 (N_4614,In_1017,In_475);
nor U4615 (N_4615,In_1497,In_661);
nand U4616 (N_4616,In_371,In_1044);
and U4617 (N_4617,In_766,In_732);
or U4618 (N_4618,In_383,In_1377);
or U4619 (N_4619,In_618,In_714);
nor U4620 (N_4620,In_603,In_836);
nand U4621 (N_4621,In_809,In_749);
or U4622 (N_4622,In_338,In_1329);
and U4623 (N_4623,In_231,In_969);
or U4624 (N_4624,In_742,In_175);
nand U4625 (N_4625,In_846,In_412);
nor U4626 (N_4626,In_216,In_36);
nand U4627 (N_4627,In_1155,In_1425);
or U4628 (N_4628,In_1279,In_440);
and U4629 (N_4629,In_1259,In_447);
and U4630 (N_4630,In_44,In_456);
nand U4631 (N_4631,In_322,In_701);
or U4632 (N_4632,In_393,In_416);
or U4633 (N_4633,In_588,In_547);
and U4634 (N_4634,In_138,In_1132);
or U4635 (N_4635,In_413,In_713);
nand U4636 (N_4636,In_353,In_713);
and U4637 (N_4637,In_39,In_1388);
xor U4638 (N_4638,In_1445,In_285);
and U4639 (N_4639,In_247,In_992);
nand U4640 (N_4640,In_249,In_1208);
or U4641 (N_4641,In_540,In_746);
or U4642 (N_4642,In_1161,In_1355);
nor U4643 (N_4643,In_1096,In_1477);
or U4644 (N_4644,In_1272,In_1026);
nor U4645 (N_4645,In_1191,In_1357);
or U4646 (N_4646,In_882,In_293);
xor U4647 (N_4647,In_1029,In_1437);
and U4648 (N_4648,In_1420,In_631);
and U4649 (N_4649,In_173,In_1015);
nor U4650 (N_4650,In_1393,In_355);
or U4651 (N_4651,In_1389,In_927);
nor U4652 (N_4652,In_415,In_888);
nor U4653 (N_4653,In_143,In_1490);
nor U4654 (N_4654,In_341,In_886);
and U4655 (N_4655,In_442,In_30);
xnor U4656 (N_4656,In_431,In_144);
or U4657 (N_4657,In_762,In_339);
nor U4658 (N_4658,In_1470,In_5);
nand U4659 (N_4659,In_988,In_1477);
and U4660 (N_4660,In_906,In_1144);
or U4661 (N_4661,In_273,In_1264);
or U4662 (N_4662,In_1155,In_920);
nor U4663 (N_4663,In_1138,In_96);
nor U4664 (N_4664,In_394,In_317);
nor U4665 (N_4665,In_570,In_221);
or U4666 (N_4666,In_744,In_1299);
and U4667 (N_4667,In_1238,In_51);
nor U4668 (N_4668,In_919,In_217);
or U4669 (N_4669,In_578,In_25);
xor U4670 (N_4670,In_1458,In_561);
and U4671 (N_4671,In_1393,In_379);
nand U4672 (N_4672,In_149,In_275);
nand U4673 (N_4673,In_1113,In_1284);
nand U4674 (N_4674,In_145,In_582);
and U4675 (N_4675,In_571,In_1491);
or U4676 (N_4676,In_138,In_1121);
nand U4677 (N_4677,In_1226,In_1496);
and U4678 (N_4678,In_1382,In_1136);
or U4679 (N_4679,In_792,In_1315);
nand U4680 (N_4680,In_689,In_960);
or U4681 (N_4681,In_392,In_39);
or U4682 (N_4682,In_478,In_1487);
nor U4683 (N_4683,In_714,In_1030);
and U4684 (N_4684,In_301,In_231);
and U4685 (N_4685,In_1181,In_931);
nor U4686 (N_4686,In_1401,In_1330);
and U4687 (N_4687,In_127,In_1477);
and U4688 (N_4688,In_633,In_1287);
nand U4689 (N_4689,In_1382,In_285);
nor U4690 (N_4690,In_397,In_907);
or U4691 (N_4691,In_1010,In_1216);
and U4692 (N_4692,In_1339,In_1198);
nor U4693 (N_4693,In_592,In_1038);
nand U4694 (N_4694,In_963,In_736);
nand U4695 (N_4695,In_693,In_337);
and U4696 (N_4696,In_840,In_892);
and U4697 (N_4697,In_1460,In_417);
and U4698 (N_4698,In_358,In_268);
nor U4699 (N_4699,In_1426,In_1379);
or U4700 (N_4700,In_451,In_1243);
and U4701 (N_4701,In_234,In_278);
and U4702 (N_4702,In_1449,In_1315);
or U4703 (N_4703,In_1242,In_1037);
nor U4704 (N_4704,In_645,In_364);
or U4705 (N_4705,In_1310,In_580);
or U4706 (N_4706,In_513,In_845);
nand U4707 (N_4707,In_73,In_16);
and U4708 (N_4708,In_179,In_1367);
or U4709 (N_4709,In_1138,In_1335);
or U4710 (N_4710,In_733,In_919);
nand U4711 (N_4711,In_119,In_207);
and U4712 (N_4712,In_1264,In_629);
nor U4713 (N_4713,In_388,In_296);
xnor U4714 (N_4714,In_1353,In_1188);
nor U4715 (N_4715,In_575,In_938);
and U4716 (N_4716,In_1214,In_373);
or U4717 (N_4717,In_865,In_373);
nand U4718 (N_4718,In_1279,In_704);
and U4719 (N_4719,In_838,In_1295);
nand U4720 (N_4720,In_104,In_497);
and U4721 (N_4721,In_883,In_33);
or U4722 (N_4722,In_739,In_270);
and U4723 (N_4723,In_970,In_57);
nand U4724 (N_4724,In_647,In_1355);
nand U4725 (N_4725,In_305,In_1136);
nand U4726 (N_4726,In_1059,In_365);
nand U4727 (N_4727,In_1217,In_438);
nor U4728 (N_4728,In_1415,In_459);
and U4729 (N_4729,In_1119,In_371);
and U4730 (N_4730,In_752,In_1365);
nand U4731 (N_4731,In_875,In_900);
nand U4732 (N_4732,In_850,In_852);
and U4733 (N_4733,In_301,In_1084);
and U4734 (N_4734,In_589,In_958);
and U4735 (N_4735,In_319,In_959);
and U4736 (N_4736,In_1441,In_738);
and U4737 (N_4737,In_760,In_951);
nand U4738 (N_4738,In_219,In_817);
nor U4739 (N_4739,In_90,In_1375);
nor U4740 (N_4740,In_700,In_501);
nand U4741 (N_4741,In_274,In_29);
or U4742 (N_4742,In_1098,In_241);
and U4743 (N_4743,In_1458,In_570);
or U4744 (N_4744,In_342,In_546);
and U4745 (N_4745,In_1237,In_955);
nand U4746 (N_4746,In_1459,In_1488);
and U4747 (N_4747,In_152,In_1348);
nor U4748 (N_4748,In_616,In_1426);
nand U4749 (N_4749,In_1029,In_1329);
nor U4750 (N_4750,In_129,In_1157);
and U4751 (N_4751,In_576,In_1327);
and U4752 (N_4752,In_1290,In_1066);
nand U4753 (N_4753,In_1324,In_311);
nor U4754 (N_4754,In_688,In_621);
nor U4755 (N_4755,In_63,In_873);
nand U4756 (N_4756,In_1238,In_328);
and U4757 (N_4757,In_609,In_846);
or U4758 (N_4758,In_1443,In_456);
nand U4759 (N_4759,In_1313,In_1112);
and U4760 (N_4760,In_1409,In_672);
nor U4761 (N_4761,In_984,In_277);
or U4762 (N_4762,In_349,In_1485);
nor U4763 (N_4763,In_601,In_520);
nand U4764 (N_4764,In_213,In_721);
nand U4765 (N_4765,In_453,In_447);
nand U4766 (N_4766,In_0,In_736);
and U4767 (N_4767,In_616,In_30);
nand U4768 (N_4768,In_1419,In_88);
nand U4769 (N_4769,In_782,In_972);
and U4770 (N_4770,In_315,In_747);
or U4771 (N_4771,In_135,In_1168);
or U4772 (N_4772,In_884,In_1328);
or U4773 (N_4773,In_1024,In_190);
nand U4774 (N_4774,In_410,In_487);
nand U4775 (N_4775,In_1436,In_540);
and U4776 (N_4776,In_1069,In_553);
nand U4777 (N_4777,In_1129,In_1213);
nand U4778 (N_4778,In_260,In_168);
nand U4779 (N_4779,In_326,In_1005);
xor U4780 (N_4780,In_1015,In_197);
or U4781 (N_4781,In_1181,In_539);
nor U4782 (N_4782,In_1068,In_585);
and U4783 (N_4783,In_790,In_349);
or U4784 (N_4784,In_414,In_720);
and U4785 (N_4785,In_1099,In_201);
or U4786 (N_4786,In_366,In_1225);
and U4787 (N_4787,In_1068,In_65);
and U4788 (N_4788,In_1016,In_544);
nand U4789 (N_4789,In_210,In_162);
and U4790 (N_4790,In_1459,In_669);
nor U4791 (N_4791,In_482,In_275);
or U4792 (N_4792,In_1356,In_1124);
nor U4793 (N_4793,In_1469,In_320);
nor U4794 (N_4794,In_805,In_1163);
and U4795 (N_4795,In_1441,In_1095);
nand U4796 (N_4796,In_181,In_785);
or U4797 (N_4797,In_1232,In_631);
xnor U4798 (N_4798,In_797,In_786);
nor U4799 (N_4799,In_823,In_928);
nand U4800 (N_4800,In_492,In_330);
nand U4801 (N_4801,In_815,In_1133);
nor U4802 (N_4802,In_662,In_964);
or U4803 (N_4803,In_888,In_1196);
nor U4804 (N_4804,In_643,In_1138);
and U4805 (N_4805,In_916,In_1152);
nor U4806 (N_4806,In_526,In_1229);
and U4807 (N_4807,In_1221,In_738);
nand U4808 (N_4808,In_724,In_471);
nand U4809 (N_4809,In_468,In_120);
or U4810 (N_4810,In_866,In_396);
or U4811 (N_4811,In_100,In_756);
nand U4812 (N_4812,In_763,In_1456);
nand U4813 (N_4813,In_1167,In_288);
nand U4814 (N_4814,In_905,In_1400);
nand U4815 (N_4815,In_1062,In_46);
nor U4816 (N_4816,In_962,In_1091);
nand U4817 (N_4817,In_14,In_88);
nand U4818 (N_4818,In_816,In_205);
nand U4819 (N_4819,In_378,In_77);
nand U4820 (N_4820,In_1443,In_742);
nor U4821 (N_4821,In_66,In_1355);
and U4822 (N_4822,In_742,In_1166);
or U4823 (N_4823,In_1017,In_1091);
nor U4824 (N_4824,In_1405,In_507);
nor U4825 (N_4825,In_1013,In_166);
or U4826 (N_4826,In_1454,In_393);
and U4827 (N_4827,In_924,In_1111);
and U4828 (N_4828,In_509,In_1321);
and U4829 (N_4829,In_1070,In_466);
and U4830 (N_4830,In_501,In_1118);
and U4831 (N_4831,In_496,In_40);
or U4832 (N_4832,In_295,In_840);
nand U4833 (N_4833,In_55,In_1299);
or U4834 (N_4834,In_1460,In_635);
and U4835 (N_4835,In_888,In_529);
nand U4836 (N_4836,In_500,In_382);
nand U4837 (N_4837,In_722,In_344);
nor U4838 (N_4838,In_600,In_649);
or U4839 (N_4839,In_823,In_846);
or U4840 (N_4840,In_317,In_613);
nor U4841 (N_4841,In_1256,In_886);
or U4842 (N_4842,In_731,In_1135);
nor U4843 (N_4843,In_918,In_50);
or U4844 (N_4844,In_203,In_1283);
xor U4845 (N_4845,In_735,In_104);
and U4846 (N_4846,In_141,In_1029);
nand U4847 (N_4847,In_778,In_642);
nor U4848 (N_4848,In_159,In_1315);
or U4849 (N_4849,In_419,In_208);
and U4850 (N_4850,In_56,In_1046);
nand U4851 (N_4851,In_490,In_58);
nand U4852 (N_4852,In_918,In_942);
nor U4853 (N_4853,In_877,In_203);
nor U4854 (N_4854,In_739,In_1499);
or U4855 (N_4855,In_1076,In_205);
and U4856 (N_4856,In_299,In_622);
and U4857 (N_4857,In_852,In_964);
nand U4858 (N_4858,In_1063,In_248);
nor U4859 (N_4859,In_1247,In_1099);
nor U4860 (N_4860,In_1308,In_916);
xor U4861 (N_4861,In_844,In_512);
and U4862 (N_4862,In_375,In_713);
nor U4863 (N_4863,In_1036,In_1162);
or U4864 (N_4864,In_886,In_595);
and U4865 (N_4865,In_950,In_646);
or U4866 (N_4866,In_716,In_663);
or U4867 (N_4867,In_1368,In_398);
or U4868 (N_4868,In_566,In_1426);
nand U4869 (N_4869,In_531,In_115);
or U4870 (N_4870,In_1241,In_401);
nor U4871 (N_4871,In_682,In_534);
or U4872 (N_4872,In_1432,In_619);
and U4873 (N_4873,In_812,In_1430);
nand U4874 (N_4874,In_1225,In_730);
nor U4875 (N_4875,In_1148,In_952);
nand U4876 (N_4876,In_1172,In_995);
and U4877 (N_4877,In_1241,In_5);
nand U4878 (N_4878,In_1171,In_1011);
nand U4879 (N_4879,In_594,In_354);
nor U4880 (N_4880,In_996,In_170);
and U4881 (N_4881,In_85,In_183);
or U4882 (N_4882,In_516,In_894);
or U4883 (N_4883,In_349,In_318);
or U4884 (N_4884,In_894,In_327);
and U4885 (N_4885,In_703,In_713);
or U4886 (N_4886,In_539,In_1005);
nor U4887 (N_4887,In_1427,In_1254);
or U4888 (N_4888,In_1006,In_668);
nor U4889 (N_4889,In_558,In_323);
nor U4890 (N_4890,In_1261,In_294);
xor U4891 (N_4891,In_22,In_1436);
nand U4892 (N_4892,In_346,In_1066);
and U4893 (N_4893,In_603,In_111);
or U4894 (N_4894,In_1396,In_288);
nand U4895 (N_4895,In_1499,In_503);
or U4896 (N_4896,In_723,In_1415);
nor U4897 (N_4897,In_123,In_689);
nand U4898 (N_4898,In_554,In_1103);
xnor U4899 (N_4899,In_1444,In_632);
xor U4900 (N_4900,In_1444,In_508);
nor U4901 (N_4901,In_574,In_49);
and U4902 (N_4902,In_1124,In_1155);
and U4903 (N_4903,In_390,In_1215);
and U4904 (N_4904,In_474,In_1314);
and U4905 (N_4905,In_642,In_535);
nor U4906 (N_4906,In_452,In_416);
or U4907 (N_4907,In_1050,In_1381);
nor U4908 (N_4908,In_272,In_1329);
nand U4909 (N_4909,In_1442,In_937);
xnor U4910 (N_4910,In_1006,In_216);
xnor U4911 (N_4911,In_457,In_1314);
nand U4912 (N_4912,In_900,In_889);
nor U4913 (N_4913,In_858,In_1108);
nand U4914 (N_4914,In_705,In_1177);
and U4915 (N_4915,In_442,In_1146);
nor U4916 (N_4916,In_146,In_462);
and U4917 (N_4917,In_756,In_1137);
xor U4918 (N_4918,In_1351,In_570);
or U4919 (N_4919,In_184,In_408);
and U4920 (N_4920,In_509,In_409);
and U4921 (N_4921,In_838,In_1179);
or U4922 (N_4922,In_1070,In_883);
or U4923 (N_4923,In_454,In_53);
or U4924 (N_4924,In_1260,In_603);
or U4925 (N_4925,In_1145,In_997);
nand U4926 (N_4926,In_149,In_265);
nand U4927 (N_4927,In_296,In_80);
or U4928 (N_4928,In_344,In_428);
nor U4929 (N_4929,In_1419,In_613);
nor U4930 (N_4930,In_774,In_371);
or U4931 (N_4931,In_1402,In_24);
nor U4932 (N_4932,In_1157,In_865);
or U4933 (N_4933,In_1456,In_458);
and U4934 (N_4934,In_1056,In_622);
nand U4935 (N_4935,In_1297,In_1077);
nor U4936 (N_4936,In_654,In_4);
nand U4937 (N_4937,In_370,In_1396);
and U4938 (N_4938,In_1372,In_1076);
or U4939 (N_4939,In_294,In_618);
nand U4940 (N_4940,In_758,In_770);
nor U4941 (N_4941,In_1330,In_70);
nand U4942 (N_4942,In_522,In_575);
nand U4943 (N_4943,In_37,In_1042);
nand U4944 (N_4944,In_716,In_415);
and U4945 (N_4945,In_630,In_1093);
or U4946 (N_4946,In_322,In_960);
nor U4947 (N_4947,In_859,In_818);
nand U4948 (N_4948,In_1185,In_225);
nor U4949 (N_4949,In_1043,In_178);
and U4950 (N_4950,In_615,In_859);
nand U4951 (N_4951,In_1089,In_140);
and U4952 (N_4952,In_1493,In_1329);
or U4953 (N_4953,In_1183,In_641);
nor U4954 (N_4954,In_1456,In_1091);
nand U4955 (N_4955,In_551,In_31);
nand U4956 (N_4956,In_1092,In_1311);
nor U4957 (N_4957,In_1473,In_910);
nand U4958 (N_4958,In_238,In_1400);
and U4959 (N_4959,In_139,In_830);
nand U4960 (N_4960,In_1147,In_1153);
nor U4961 (N_4961,In_446,In_712);
or U4962 (N_4962,In_1344,In_1278);
nand U4963 (N_4963,In_706,In_386);
or U4964 (N_4964,In_441,In_278);
or U4965 (N_4965,In_1482,In_383);
nor U4966 (N_4966,In_667,In_1444);
and U4967 (N_4967,In_654,In_225);
or U4968 (N_4968,In_1053,In_849);
or U4969 (N_4969,In_1262,In_880);
or U4970 (N_4970,In_1244,In_1206);
or U4971 (N_4971,In_580,In_308);
or U4972 (N_4972,In_1301,In_1378);
nor U4973 (N_4973,In_1259,In_1156);
or U4974 (N_4974,In_672,In_1002);
nor U4975 (N_4975,In_391,In_119);
or U4976 (N_4976,In_591,In_1329);
nand U4977 (N_4977,In_508,In_643);
or U4978 (N_4978,In_1211,In_1013);
nand U4979 (N_4979,In_1280,In_368);
and U4980 (N_4980,In_483,In_230);
nand U4981 (N_4981,In_744,In_297);
nand U4982 (N_4982,In_643,In_488);
nor U4983 (N_4983,In_857,In_1112);
nand U4984 (N_4984,In_1084,In_681);
or U4985 (N_4985,In_1069,In_312);
and U4986 (N_4986,In_1422,In_686);
and U4987 (N_4987,In_127,In_1298);
or U4988 (N_4988,In_813,In_1237);
nor U4989 (N_4989,In_1132,In_389);
and U4990 (N_4990,In_441,In_1463);
nor U4991 (N_4991,In_1280,In_995);
nor U4992 (N_4992,In_1059,In_594);
or U4993 (N_4993,In_943,In_818);
or U4994 (N_4994,In_812,In_667);
or U4995 (N_4995,In_620,In_301);
and U4996 (N_4996,In_162,In_65);
nand U4997 (N_4997,In_1397,In_1346);
and U4998 (N_4998,In_766,In_879);
or U4999 (N_4999,In_1217,In_540);
or U5000 (N_5000,N_957,N_1985);
and U5001 (N_5001,N_1788,N_1997);
nand U5002 (N_5002,N_4247,N_892);
or U5003 (N_5003,N_1687,N_2195);
nor U5004 (N_5004,N_3445,N_1099);
nor U5005 (N_5005,N_2007,N_1237);
and U5006 (N_5006,N_2864,N_4955);
or U5007 (N_5007,N_4868,N_3886);
nand U5008 (N_5008,N_3453,N_2916);
nor U5009 (N_5009,N_2473,N_4354);
xor U5010 (N_5010,N_1897,N_1545);
nor U5011 (N_5011,N_862,N_1304);
nor U5012 (N_5012,N_1112,N_1274);
or U5013 (N_5013,N_1488,N_679);
nor U5014 (N_5014,N_144,N_4801);
or U5015 (N_5015,N_4001,N_3325);
or U5016 (N_5016,N_3246,N_1937);
or U5017 (N_5017,N_401,N_1700);
nand U5018 (N_5018,N_2614,N_153);
or U5019 (N_5019,N_3153,N_3649);
or U5020 (N_5020,N_1000,N_2305);
nor U5021 (N_5021,N_3286,N_328);
or U5022 (N_5022,N_3574,N_2082);
or U5023 (N_5023,N_1370,N_2901);
or U5024 (N_5024,N_3425,N_4463);
nor U5025 (N_5025,N_3929,N_1460);
nor U5026 (N_5026,N_4461,N_469);
and U5027 (N_5027,N_1577,N_1093);
nor U5028 (N_5028,N_2727,N_2307);
nand U5029 (N_5029,N_4190,N_4958);
and U5030 (N_5030,N_3684,N_4583);
or U5031 (N_5031,N_1121,N_1390);
nand U5032 (N_5032,N_3529,N_4739);
and U5033 (N_5033,N_271,N_3087);
nand U5034 (N_5034,N_3959,N_2593);
nand U5035 (N_5035,N_4092,N_4339);
nor U5036 (N_5036,N_3777,N_4347);
and U5037 (N_5037,N_841,N_657);
nand U5038 (N_5038,N_3285,N_4145);
and U5039 (N_5039,N_3779,N_1914);
nand U5040 (N_5040,N_989,N_1829);
and U5041 (N_5041,N_2596,N_2976);
nor U5042 (N_5042,N_539,N_3981);
nor U5043 (N_5043,N_4249,N_2670);
or U5044 (N_5044,N_2472,N_2642);
nor U5045 (N_5045,N_3015,N_2832);
or U5046 (N_5046,N_1768,N_4512);
nand U5047 (N_5047,N_4074,N_2504);
or U5048 (N_5048,N_1281,N_4416);
and U5049 (N_5049,N_1042,N_1964);
or U5050 (N_5050,N_2722,N_155);
nor U5051 (N_5051,N_3864,N_2479);
or U5052 (N_5052,N_3210,N_2265);
nand U5053 (N_5053,N_935,N_1260);
nor U5054 (N_5054,N_312,N_1936);
xnor U5055 (N_5055,N_4846,N_2729);
nand U5056 (N_5056,N_3622,N_4157);
and U5057 (N_5057,N_3008,N_3914);
nor U5058 (N_5058,N_1570,N_2143);
nor U5059 (N_5059,N_2737,N_4123);
and U5060 (N_5060,N_1194,N_1875);
nor U5061 (N_5061,N_3016,N_3347);
nor U5062 (N_5062,N_4900,N_2322);
nand U5063 (N_5063,N_4112,N_1148);
and U5064 (N_5064,N_1566,N_22);
and U5065 (N_5065,N_2960,N_1809);
nand U5066 (N_5066,N_2277,N_1991);
or U5067 (N_5067,N_4980,N_1192);
and U5068 (N_5068,N_3330,N_4363);
and U5069 (N_5069,N_4834,N_3855);
or U5070 (N_5070,N_79,N_2632);
nand U5071 (N_5071,N_3993,N_3056);
or U5072 (N_5072,N_214,N_2895);
and U5073 (N_5073,N_2657,N_852);
or U5074 (N_5074,N_4518,N_545);
nor U5075 (N_5075,N_3612,N_4838);
or U5076 (N_5076,N_4300,N_3221);
and U5077 (N_5077,N_1317,N_1693);
and U5078 (N_5078,N_1306,N_2073);
or U5079 (N_5079,N_2661,N_350);
nor U5080 (N_5080,N_927,N_3251);
and U5081 (N_5081,N_4978,N_3515);
and U5082 (N_5082,N_3320,N_4965);
nand U5083 (N_5083,N_3434,N_991);
nor U5084 (N_5084,N_4093,N_4195);
nor U5085 (N_5085,N_4820,N_3033);
nor U5086 (N_5086,N_4564,N_3063);
and U5087 (N_5087,N_3472,N_930);
and U5088 (N_5088,N_3339,N_2689);
and U5089 (N_5089,N_2666,N_675);
and U5090 (N_5090,N_1778,N_1691);
nor U5091 (N_5091,N_177,N_4208);
nor U5092 (N_5092,N_950,N_2432);
nor U5093 (N_5093,N_1628,N_1073);
or U5094 (N_5094,N_1839,N_2584);
nand U5095 (N_5095,N_4643,N_4177);
nand U5096 (N_5096,N_1398,N_2550);
or U5097 (N_5097,N_48,N_4813);
nand U5098 (N_5098,N_1689,N_1535);
and U5099 (N_5099,N_2933,N_2868);
or U5100 (N_5100,N_3396,N_1679);
nand U5101 (N_5101,N_4106,N_4165);
or U5102 (N_5102,N_4213,N_4655);
or U5103 (N_5103,N_531,N_15);
and U5104 (N_5104,N_2109,N_4623);
or U5105 (N_5105,N_1650,N_412);
nand U5106 (N_5106,N_2478,N_1155);
nand U5107 (N_5107,N_4052,N_554);
nor U5108 (N_5108,N_3790,N_1838);
nand U5109 (N_5109,N_2886,N_91);
nand U5110 (N_5110,N_2229,N_2664);
nor U5111 (N_5111,N_4714,N_1951);
xor U5112 (N_5112,N_2025,N_2829);
nor U5113 (N_5113,N_3894,N_4443);
or U5114 (N_5114,N_4614,N_1556);
nor U5115 (N_5115,N_3294,N_1568);
nand U5116 (N_5116,N_3494,N_4585);
nor U5117 (N_5117,N_2294,N_3589);
nor U5118 (N_5118,N_3838,N_4959);
and U5119 (N_5119,N_1717,N_1606);
nand U5120 (N_5120,N_1228,N_2574);
nor U5121 (N_5121,N_2761,N_343);
or U5122 (N_5122,N_4149,N_183);
nand U5123 (N_5123,N_1225,N_347);
nor U5124 (N_5124,N_284,N_4857);
or U5125 (N_5125,N_4982,N_1418);
and U5126 (N_5126,N_3224,N_2507);
or U5127 (N_5127,N_4310,N_2370);
and U5128 (N_5128,N_4171,N_905);
nor U5129 (N_5129,N_2672,N_972);
or U5130 (N_5130,N_4881,N_4228);
and U5131 (N_5131,N_360,N_3311);
and U5132 (N_5132,N_4484,N_3922);
or U5133 (N_5133,N_4329,N_3764);
nand U5134 (N_5134,N_87,N_58);
nand U5135 (N_5135,N_3771,N_267);
nand U5136 (N_5136,N_3729,N_3401);
nor U5137 (N_5137,N_1492,N_3484);
or U5138 (N_5138,N_854,N_3551);
nor U5139 (N_5139,N_740,N_3348);
nand U5140 (N_5140,N_3030,N_3991);
or U5141 (N_5141,N_399,N_1822);
nand U5142 (N_5142,N_4648,N_3789);
nor U5143 (N_5143,N_4055,N_1866);
and U5144 (N_5144,N_4712,N_1823);
or U5145 (N_5145,N_566,N_1278);
nor U5146 (N_5146,N_4636,N_650);
nand U5147 (N_5147,N_2788,N_618);
nand U5148 (N_5148,N_4109,N_584);
nand U5149 (N_5149,N_3587,N_2755);
nand U5150 (N_5150,N_834,N_607);
nand U5151 (N_5151,N_644,N_3868);
or U5152 (N_5152,N_2090,N_4121);
nor U5153 (N_5153,N_3882,N_4925);
nor U5154 (N_5154,N_1119,N_2430);
nand U5155 (N_5155,N_151,N_1083);
or U5156 (N_5156,N_2137,N_2845);
nand U5157 (N_5157,N_4624,N_3276);
nor U5158 (N_5158,N_3439,N_2450);
nand U5159 (N_5159,N_3860,N_4462);
and U5160 (N_5160,N_1223,N_435);
nor U5161 (N_5161,N_2088,N_560);
nand U5162 (N_5162,N_1769,N_1142);
nor U5163 (N_5163,N_1308,N_816);
or U5164 (N_5164,N_3140,N_4967);
nor U5165 (N_5165,N_2493,N_1157);
nor U5166 (N_5166,N_3787,N_3360);
or U5167 (N_5167,N_217,N_132);
or U5168 (N_5168,N_1078,N_770);
nor U5169 (N_5169,N_4550,N_2454);
nor U5170 (N_5170,N_3700,N_1865);
nor U5171 (N_5171,N_3531,N_4571);
nand U5172 (N_5172,N_3756,N_1893);
nor U5173 (N_5173,N_419,N_1319);
or U5174 (N_5174,N_4546,N_2070);
and U5175 (N_5175,N_2249,N_215);
nor U5176 (N_5176,N_1071,N_1444);
or U5177 (N_5177,N_3436,N_586);
nor U5178 (N_5178,N_4283,N_1002);
and U5179 (N_5179,N_2847,N_4498);
and U5180 (N_5180,N_1811,N_689);
nand U5181 (N_5181,N_3072,N_590);
nor U5182 (N_5182,N_4128,N_2004);
or U5183 (N_5183,N_1993,N_1562);
nor U5184 (N_5184,N_999,N_2499);
and U5185 (N_5185,N_2921,N_1626);
nand U5186 (N_5186,N_1928,N_1485);
and U5187 (N_5187,N_1555,N_4433);
nand U5188 (N_5188,N_242,N_2183);
nor U5189 (N_5189,N_699,N_4336);
and U5190 (N_5190,N_1417,N_2136);
or U5191 (N_5191,N_3770,N_4302);
or U5192 (N_5192,N_2896,N_4229);
nand U5193 (N_5193,N_3923,N_1733);
nand U5194 (N_5194,N_2261,N_2810);
and U5195 (N_5195,N_307,N_1);
or U5196 (N_5196,N_2974,N_1395);
or U5197 (N_5197,N_3471,N_1493);
or U5198 (N_5198,N_385,N_2080);
nor U5199 (N_5199,N_4789,N_996);
and U5200 (N_5200,N_3480,N_774);
nor U5201 (N_5201,N_420,N_2463);
nor U5202 (N_5202,N_570,N_911);
or U5203 (N_5203,N_1124,N_4694);
nand U5204 (N_5204,N_3586,N_798);
nor U5205 (N_5205,N_4017,N_4163);
or U5206 (N_5206,N_163,N_453);
nand U5207 (N_5207,N_1075,N_2988);
or U5208 (N_5208,N_2096,N_683);
or U5209 (N_5209,N_626,N_1050);
nor U5210 (N_5210,N_1796,N_1096);
or U5211 (N_5211,N_3812,N_2992);
nor U5212 (N_5212,N_1898,N_3769);
nor U5213 (N_5213,N_813,N_3382);
and U5214 (N_5214,N_2012,N_3819);
and U5215 (N_5215,N_1479,N_748);
nand U5216 (N_5216,N_3566,N_2606);
nand U5217 (N_5217,N_1920,N_1290);
nand U5218 (N_5218,N_3517,N_4987);
or U5219 (N_5219,N_4768,N_3763);
nor U5220 (N_5220,N_147,N_3485);
nand U5221 (N_5221,N_2332,N_1267);
or U5222 (N_5222,N_3440,N_1472);
or U5223 (N_5223,N_1825,N_1402);
and U5224 (N_5224,N_1851,N_646);
nand U5225 (N_5225,N_756,N_4822);
and U5226 (N_5226,N_2978,N_3617);
nand U5227 (N_5227,N_3949,N_4125);
and U5228 (N_5228,N_1160,N_4220);
xnor U5229 (N_5229,N_92,N_3924);
and U5230 (N_5230,N_3887,N_901);
and U5231 (N_5231,N_67,N_2184);
or U5232 (N_5232,N_1334,N_1175);
or U5233 (N_5233,N_1540,N_4337);
and U5234 (N_5234,N_2271,N_4540);
nor U5235 (N_5235,N_1584,N_4821);
and U5236 (N_5236,N_1750,N_3389);
nand U5237 (N_5237,N_979,N_4612);
xnor U5238 (N_5238,N_3190,N_3960);
nand U5239 (N_5239,N_3352,N_4711);
nor U5240 (N_5240,N_2418,N_2065);
nand U5241 (N_5241,N_4019,N_3279);
and U5242 (N_5242,N_1454,N_1311);
nor U5243 (N_5243,N_1176,N_2994);
nand U5244 (N_5244,N_2640,N_4388);
and U5245 (N_5245,N_76,N_1403);
or U5246 (N_5246,N_397,N_3902);
nand U5247 (N_5247,N_2132,N_416);
and U5248 (N_5248,N_2809,N_4779);
nand U5249 (N_5249,N_4761,N_305);
or U5250 (N_5250,N_477,N_1600);
nand U5251 (N_5251,N_2531,N_1658);
and U5252 (N_5252,N_4763,N_4572);
nand U5253 (N_5253,N_4552,N_641);
nor U5254 (N_5254,N_1867,N_1242);
or U5255 (N_5255,N_1601,N_35);
nand U5256 (N_5256,N_3800,N_186);
nor U5257 (N_5257,N_4580,N_1392);
or U5258 (N_5258,N_2399,N_797);
nor U5259 (N_5259,N_365,N_3313);
nor U5260 (N_5260,N_1410,N_363);
nand U5261 (N_5261,N_333,N_100);
or U5262 (N_5262,N_906,N_512);
nor U5263 (N_5263,N_963,N_3073);
nand U5264 (N_5264,N_3862,N_1036);
or U5265 (N_5265,N_4780,N_3618);
nor U5266 (N_5266,N_700,N_2516);
nand U5267 (N_5267,N_1878,N_1956);
or U5268 (N_5268,N_2279,N_701);
nor U5269 (N_5269,N_13,N_611);
or U5270 (N_5270,N_450,N_2853);
and U5271 (N_5271,N_2773,N_1725);
nand U5272 (N_5272,N_2411,N_3806);
nand U5273 (N_5273,N_3452,N_4863);
and U5274 (N_5274,N_4501,N_4601);
and U5275 (N_5275,N_1205,N_2006);
nor U5276 (N_5276,N_4293,N_235);
and U5277 (N_5277,N_921,N_1660);
and U5278 (N_5278,N_2017,N_2009);
or U5279 (N_5279,N_3654,N_1130);
nand U5280 (N_5280,N_1844,N_44);
nand U5281 (N_5281,N_3671,N_2804);
nor U5282 (N_5282,N_2240,N_1007);
nor U5283 (N_5283,N_3572,N_1753);
or U5284 (N_5284,N_2700,N_1044);
or U5285 (N_5285,N_2071,N_265);
nand U5286 (N_5286,N_4320,N_1828);
nor U5287 (N_5287,N_2151,N_3776);
nor U5288 (N_5288,N_2633,N_4589);
nand U5289 (N_5289,N_2913,N_615);
nor U5290 (N_5290,N_1365,N_3326);
and U5291 (N_5291,N_2708,N_2511);
nor U5292 (N_5292,N_3738,N_1917);
and U5293 (N_5293,N_313,N_1017);
nor U5294 (N_5294,N_3542,N_1405);
and U5295 (N_5295,N_1827,N_2310);
or U5296 (N_5296,N_3492,N_3076);
and U5297 (N_5297,N_3266,N_4217);
nand U5298 (N_5298,N_4609,N_104);
or U5299 (N_5299,N_787,N_3715);
xor U5300 (N_5300,N_3045,N_2946);
nor U5301 (N_5301,N_595,N_2157);
or U5302 (N_5302,N_1940,N_10);
and U5303 (N_5303,N_3538,N_2687);
nand U5304 (N_5304,N_4375,N_3535);
or U5305 (N_5305,N_3052,N_1673);
and U5306 (N_5306,N_4349,N_3874);
nand U5307 (N_5307,N_1593,N_1462);
and U5308 (N_5308,N_4913,N_2945);
or U5309 (N_5309,N_361,N_3926);
nand U5310 (N_5310,N_3238,N_757);
or U5311 (N_5311,N_4452,N_2167);
xor U5312 (N_5312,N_3412,N_188);
or U5313 (N_5313,N_369,N_2681);
and U5314 (N_5314,N_4448,N_4333);
and U5315 (N_5315,N_3039,N_793);
and U5316 (N_5316,N_2091,N_2843);
nand U5317 (N_5317,N_3780,N_902);
and U5318 (N_5318,N_4211,N_3252);
nand U5319 (N_5319,N_4639,N_845);
nand U5320 (N_5320,N_2095,N_494);
and U5321 (N_5321,N_1172,N_1183);
nand U5322 (N_5322,N_1863,N_1775);
nand U5323 (N_5323,N_1948,N_1275);
and U5324 (N_5324,N_4702,N_636);
and U5325 (N_5325,N_3206,N_3534);
or U5326 (N_5326,N_4746,N_730);
nand U5327 (N_5327,N_4442,N_1052);
nand U5328 (N_5328,N_4940,N_2239);
nor U5329 (N_5329,N_2925,N_3644);
nor U5330 (N_5330,N_2630,N_3130);
nand U5331 (N_5331,N_2369,N_4566);
and U5332 (N_5332,N_3111,N_2032);
nor U5333 (N_5333,N_2287,N_2387);
nor U5334 (N_5334,N_507,N_1815);
nand U5335 (N_5335,N_2003,N_73);
nor U5336 (N_5336,N_4704,N_3463);
nor U5337 (N_5337,N_1374,N_3479);
and U5338 (N_5338,N_891,N_4878);
xor U5339 (N_5339,N_1590,N_488);
nor U5340 (N_5340,N_3977,N_4662);
nand U5341 (N_5341,N_1082,N_2354);
nor U5342 (N_5342,N_2683,N_336);
nand U5343 (N_5343,N_2045,N_165);
nand U5344 (N_5344,N_3131,N_3513);
and U5345 (N_5345,N_1412,N_421);
and U5346 (N_5346,N_3971,N_2748);
or U5347 (N_5347,N_4491,N_211);
nor U5348 (N_5348,N_106,N_665);
nor U5349 (N_5349,N_4826,N_1504);
nor U5350 (N_5350,N_3293,N_3701);
or U5351 (N_5351,N_4446,N_1424);
nand U5352 (N_5352,N_1214,N_111);
nand U5353 (N_5353,N_1615,N_2841);
and U5354 (N_5354,N_2892,N_4595);
or U5355 (N_5355,N_684,N_3999);
or U5356 (N_5356,N_3081,N_3196);
and U5357 (N_5357,N_1713,N_1816);
or U5358 (N_5358,N_4472,N_2826);
nand U5359 (N_5359,N_1734,N_3831);
or U5360 (N_5360,N_2119,N_4428);
nand U5361 (N_5361,N_970,N_4808);
or U5362 (N_5362,N_299,N_1323);
nor U5363 (N_5363,N_1468,N_233);
nand U5364 (N_5364,N_219,N_61);
and U5365 (N_5365,N_3343,N_2777);
or U5366 (N_5366,N_18,N_2850);
xnor U5367 (N_5367,N_1276,N_3970);
nor U5368 (N_5368,N_923,N_718);
nor U5369 (N_5369,N_3105,N_4539);
and U5370 (N_5370,N_3112,N_2251);
or U5371 (N_5371,N_4647,N_2154);
nor U5372 (N_5372,N_4917,N_1469);
and U5373 (N_5373,N_4101,N_2176);
and U5374 (N_5374,N_2528,N_3584);
nor U5375 (N_5375,N_2150,N_2612);
or U5376 (N_5376,N_4565,N_1722);
nand U5377 (N_5377,N_1831,N_705);
and U5378 (N_5378,N_4697,N_1164);
and U5379 (N_5379,N_3891,N_1880);
or U5380 (N_5380,N_4759,N_3386);
and U5381 (N_5381,N_3691,N_998);
nor U5382 (N_5382,N_2789,N_4964);
and U5383 (N_5383,N_680,N_1944);
or U5384 (N_5384,N_2138,N_1874);
xor U5385 (N_5385,N_1683,N_4773);
and U5386 (N_5386,N_1109,N_1671);
or U5387 (N_5387,N_3797,N_120);
nor U5388 (N_5388,N_4383,N_1298);
nor U5389 (N_5389,N_2468,N_43);
nand U5390 (N_5390,N_4576,N_2015);
and U5391 (N_5391,N_3665,N_62);
and U5392 (N_5392,N_3387,N_1024);
or U5393 (N_5393,N_4269,N_2539);
or U5394 (N_5394,N_1791,N_1710);
or U5395 (N_5395,N_4633,N_3065);
nor U5396 (N_5396,N_3402,N_2569);
nand U5397 (N_5397,N_4791,N_2170);
and U5398 (N_5398,N_4689,N_1975);
or U5399 (N_5399,N_1203,N_1581);
or U5400 (N_5400,N_1727,N_4189);
nand U5401 (N_5401,N_4536,N_3486);
or U5402 (N_5402,N_721,N_666);
or U5403 (N_5403,N_1459,N_317);
or U5404 (N_5404,N_1548,N_1264);
and U5405 (N_5405,N_368,N_3690);
nand U5406 (N_5406,N_1197,N_549);
and U5407 (N_5407,N_865,N_1740);
nand U5408 (N_5408,N_1090,N_1642);
nand U5409 (N_5409,N_2967,N_2186);
nor U5410 (N_5410,N_260,N_2023);
nor U5411 (N_5411,N_652,N_565);
nand U5412 (N_5412,N_4827,N_371);
nor U5413 (N_5413,N_1602,N_3242);
or U5414 (N_5414,N_93,N_2815);
or U5415 (N_5415,N_2839,N_1283);
nand U5416 (N_5416,N_1567,N_751);
or U5417 (N_5417,N_3578,N_2028);
or U5418 (N_5418,N_3006,N_1974);
nor U5419 (N_5419,N_1560,N_3025);
nand U5420 (N_5420,N_4551,N_1903);
nor U5421 (N_5421,N_2480,N_4244);
nand U5422 (N_5422,N_4557,N_3121);
nand U5423 (N_5423,N_899,N_659);
nor U5424 (N_5424,N_2158,N_47);
xnor U5425 (N_5425,N_725,N_1107);
and U5426 (N_5426,N_3433,N_1363);
and U5427 (N_5427,N_543,N_4468);
nor U5428 (N_5428,N_3519,N_3254);
nand U5429 (N_5429,N_4951,N_2237);
nand U5430 (N_5430,N_4757,N_3271);
and U5431 (N_5431,N_2784,N_2654);
nand U5432 (N_5432,N_4311,N_4187);
nand U5433 (N_5433,N_897,N_2356);
xnor U5434 (N_5434,N_3673,N_4984);
nor U5435 (N_5435,N_1525,N_1557);
or U5436 (N_5436,N_4667,N_3910);
or U5437 (N_5437,N_2292,N_4143);
or U5438 (N_5438,N_2740,N_2616);
nor U5439 (N_5439,N_1316,N_3468);
and U5440 (N_5440,N_193,N_1565);
and U5441 (N_5441,N_2281,N_1638);
nand U5442 (N_5442,N_3341,N_3685);
nor U5443 (N_5443,N_2282,N_3658);
and U5444 (N_5444,N_4859,N_2047);
nor U5445 (N_5445,N_97,N_1620);
nand U5446 (N_5446,N_298,N_1543);
and U5447 (N_5447,N_3726,N_4018);
or U5448 (N_5448,N_2977,N_1759);
and U5449 (N_5449,N_4876,N_2807);
nand U5450 (N_5450,N_4527,N_1669);
nor U5451 (N_5451,N_4435,N_2731);
and U5452 (N_5452,N_3168,N_28);
and U5453 (N_5453,N_152,N_519);
or U5454 (N_5454,N_2048,N_4983);
nand U5455 (N_5455,N_3706,N_3185);
and U5456 (N_5456,N_29,N_1077);
nand U5457 (N_5457,N_4480,N_2002);
and U5458 (N_5458,N_3116,N_1467);
or U5459 (N_5459,N_3430,N_407);
and U5460 (N_5460,N_4556,N_2653);
or U5461 (N_5461,N_4737,N_3296);
and U5462 (N_5462,N_4563,N_2863);
or U5463 (N_5463,N_827,N_3220);
or U5464 (N_5464,N_3640,N_3421);
or U5465 (N_5465,N_2093,N_714);
or U5466 (N_5466,N_2830,N_4717);
or U5467 (N_5467,N_3151,N_113);
and U5468 (N_5468,N_4581,N_2254);
or U5469 (N_5469,N_1549,N_1058);
and U5470 (N_5470,N_1625,N_388);
nor U5471 (N_5471,N_1604,N_1592);
nand U5472 (N_5472,N_4350,N_1652);
and U5473 (N_5473,N_3441,N_2554);
and U5474 (N_5474,N_167,N_4657);
or U5475 (N_5475,N_4365,N_383);
or U5476 (N_5476,N_4236,N_4039);
and U5477 (N_5477,N_4627,N_2019);
nor U5478 (N_5478,N_513,N_2306);
or U5479 (N_5479,N_3107,N_3314);
and U5480 (N_5480,N_3132,N_2643);
nand U5481 (N_5481,N_178,N_4314);
and U5482 (N_5482,N_3097,N_1110);
nor U5483 (N_5483,N_4832,N_1977);
nand U5484 (N_5484,N_4659,N_2908);
and U5485 (N_5485,N_1150,N_1423);
and U5486 (N_5486,N_2102,N_4867);
nor U5487 (N_5487,N_4230,N_1946);
or U5488 (N_5488,N_3682,N_2835);
xor U5489 (N_5489,N_934,N_4850);
and U5490 (N_5490,N_2694,N_4621);
nor U5491 (N_5491,N_3086,N_3740);
nand U5492 (N_5492,N_2763,N_3509);
or U5493 (N_5493,N_4384,N_2624);
nand U5494 (N_5494,N_2194,N_3457);
nor U5495 (N_5495,N_4200,N_2865);
nor U5496 (N_5496,N_133,N_1301);
and U5497 (N_5497,N_4096,N_3811);
xnor U5498 (N_5498,N_562,N_3307);
or U5499 (N_5499,N_4223,N_3066);
nor U5500 (N_5500,N_3932,N_4914);
and U5501 (N_5501,N_2711,N_4814);
nor U5502 (N_5502,N_2576,N_3024);
or U5503 (N_5503,N_4665,N_4844);
nand U5504 (N_5504,N_985,N_3420);
nor U5505 (N_5505,N_3029,N_3493);
or U5506 (N_5506,N_4394,N_4252);
nor U5507 (N_5507,N_3248,N_3212);
and U5508 (N_5508,N_3843,N_4277);
nor U5509 (N_5509,N_50,N_4459);
and U5510 (N_5510,N_4594,N_3300);
and U5511 (N_5511,N_1125,N_3470);
and U5512 (N_5512,N_3367,N_2542);
nand U5513 (N_5513,N_1979,N_3222);
nand U5514 (N_5514,N_2142,N_1366);
or U5515 (N_5515,N_3051,N_2605);
nor U5516 (N_5516,N_1610,N_1749);
nor U5517 (N_5517,N_2572,N_4824);
nor U5518 (N_5518,N_2721,N_1415);
or U5519 (N_5519,N_837,N_4871);
and U5520 (N_5520,N_3328,N_3545);
nor U5521 (N_5521,N_4107,N_3793);
and U5522 (N_5522,N_400,N_3315);
nand U5523 (N_5523,N_1501,N_857);
nor U5524 (N_5524,N_3992,N_3281);
and U5525 (N_5525,N_4905,N_60);
nor U5526 (N_5526,N_1612,N_2330);
and U5527 (N_5527,N_3550,N_946);
nor U5528 (N_5528,N_1657,N_3573);
nor U5529 (N_5529,N_3070,N_391);
nor U5530 (N_5530,N_2113,N_2806);
and U5531 (N_5531,N_3568,N_2410);
and U5532 (N_5532,N_2018,N_3023);
or U5533 (N_5533,N_1864,N_3366);
and U5534 (N_5534,N_4800,N_3861);
or U5535 (N_5535,N_268,N_1739);
xnor U5536 (N_5536,N_4538,N_1841);
and U5537 (N_5537,N_2313,N_2250);
and U5538 (N_5538,N_3766,N_1375);
and U5539 (N_5539,N_2276,N_4155);
nor U5540 (N_5540,N_3174,N_440);
nor U5541 (N_5541,N_3113,N_4450);
nor U5542 (N_5542,N_1470,N_3953);
and U5543 (N_5543,N_1912,N_4535);
nand U5544 (N_5544,N_2704,N_310);
nor U5545 (N_5545,N_2378,N_1665);
nand U5546 (N_5546,N_4274,N_398);
and U5547 (N_5547,N_2920,N_457);
and U5548 (N_5548,N_2524,N_379);
and U5549 (N_5549,N_988,N_3728);
nor U5550 (N_5550,N_941,N_1456);
or U5551 (N_5551,N_2952,N_3650);
nand U5552 (N_5552,N_541,N_4483);
nor U5553 (N_5553,N_2663,N_2848);
or U5554 (N_5554,N_3466,N_2682);
nand U5555 (N_5555,N_3378,N_184);
or U5556 (N_5556,N_445,N_2690);
nand U5557 (N_5557,N_4179,N_1763);
nand U5558 (N_5558,N_83,N_3009);
or U5559 (N_5559,N_2783,N_1779);
or U5560 (N_5560,N_4849,N_4816);
or U5561 (N_5561,N_807,N_3047);
or U5562 (N_5562,N_191,N_1115);
and U5563 (N_5563,N_0,N_1342);
nor U5564 (N_5564,N_337,N_3158);
nand U5565 (N_5565,N_673,N_1681);
nand U5566 (N_5566,N_4028,N_3592);
or U5567 (N_5567,N_2774,N_3968);
or U5568 (N_5568,N_2350,N_4828);
nand U5569 (N_5569,N_2384,N_297);
and U5570 (N_5570,N_4660,N_3026);
and U5571 (N_5571,N_2595,N_1561);
and U5572 (N_5572,N_1607,N_1534);
or U5573 (N_5573,N_4831,N_1359);
and U5574 (N_5574,N_2600,N_3895);
nor U5575 (N_5575,N_2652,N_4722);
nand U5576 (N_5576,N_1177,N_2227);
and U5577 (N_5577,N_2922,N_1208);
nand U5578 (N_5578,N_2535,N_89);
nor U5579 (N_5579,N_4586,N_245);
and U5580 (N_5580,N_1254,N_1999);
and U5581 (N_5581,N_1270,N_2609);
nand U5582 (N_5582,N_2334,N_2852);
or U5583 (N_5583,N_601,N_1087);
or U5584 (N_5584,N_4895,N_1336);
and U5585 (N_5585,N_278,N_2613);
nand U5586 (N_5586,N_1513,N_964);
and U5587 (N_5587,N_1026,N_3200);
or U5588 (N_5588,N_723,N_3431);
xor U5589 (N_5589,N_800,N_4942);
and U5590 (N_5590,N_3462,N_4505);
and U5591 (N_5591,N_2975,N_4782);
nor U5592 (N_5592,N_122,N_202);
or U5593 (N_5593,N_3312,N_4764);
and U5594 (N_5594,N_4972,N_1074);
or U5595 (N_5595,N_1588,N_3954);
nand U5596 (N_5596,N_2779,N_2217);
and U5597 (N_5597,N_534,N_4058);
nand U5598 (N_5598,N_423,N_4522);
nor U5599 (N_5599,N_3627,N_2526);
nand U5600 (N_5600,N_1335,N_11);
or U5601 (N_5601,N_1324,N_1668);
and U5602 (N_5602,N_1193,N_2760);
nand U5603 (N_5603,N_4324,N_3624);
nor U5604 (N_5604,N_4701,N_2427);
nand U5605 (N_5605,N_4767,N_4212);
and U5606 (N_5606,N_1353,N_2961);
nand U5607 (N_5607,N_54,N_3336);
and U5608 (N_5608,N_2162,N_4806);
and U5609 (N_5609,N_125,N_2808);
nand U5610 (N_5610,N_2838,N_173);
and U5611 (N_5611,N_3942,N_4634);
nor U5612 (N_5612,N_3148,N_3582);
or U5613 (N_5613,N_4514,N_121);
nand U5614 (N_5614,N_4184,N_4771);
and U5615 (N_5615,N_2077,N_1383);
nor U5616 (N_5616,N_16,N_3511);
nand U5617 (N_5617,N_1812,N_4036);
or U5618 (N_5618,N_4997,N_1294);
nand U5619 (N_5619,N_3765,N_2072);
nor U5620 (N_5620,N_1550,N_4465);
and U5621 (N_5621,N_348,N_600);
xnor U5622 (N_5622,N_2385,N_2159);
nor U5623 (N_5623,N_4405,N_2264);
and U5624 (N_5624,N_4399,N_3329);
nand U5625 (N_5625,N_105,N_3890);
nor U5626 (N_5626,N_613,N_4696);
or U5627 (N_5627,N_3962,N_3907);
and U5628 (N_5628,N_2483,N_3409);
or U5629 (N_5629,N_4747,N_592);
nand U5630 (N_5630,N_1049,N_101);
or U5631 (N_5631,N_2164,N_55);
nor U5632 (N_5632,N_1876,N_3127);
or U5633 (N_5633,N_3019,N_406);
nand U5634 (N_5634,N_3080,N_1070);
nor U5635 (N_5635,N_1857,N_784);
nand U5636 (N_5636,N_34,N_311);
or U5637 (N_5637,N_1204,N_304);
and U5638 (N_5638,N_1877,N_4930);
nor U5639 (N_5639,N_953,N_815);
and U5640 (N_5640,N_4321,N_4389);
nor U5641 (N_5641,N_3205,N_3506);
nor U5642 (N_5642,N_2216,N_2347);
xor U5643 (N_5643,N_159,N_2392);
nor U5644 (N_5644,N_2750,N_707);
nand U5645 (N_5645,N_863,N_3423);
and U5646 (N_5646,N_1293,N_1756);
or U5647 (N_5647,N_342,N_3526);
and U5648 (N_5648,N_3795,N_1434);
and U5649 (N_5649,N_210,N_1960);
and U5650 (N_5650,N_1451,N_628);
nor U5651 (N_5651,N_2486,N_3979);
and U5652 (N_5652,N_3711,N_4858);
and U5653 (N_5653,N_3829,N_3904);
nand U5654 (N_5654,N_4635,N_86);
nor U5655 (N_5655,N_3759,N_654);
and U5656 (N_5656,N_4658,N_3491);
nand U5657 (N_5657,N_3651,N_2753);
nor U5658 (N_5658,N_2181,N_761);
nand U5659 (N_5659,N_573,N_1314);
nor U5660 (N_5660,N_4047,N_3866);
and U5661 (N_5661,N_358,N_3369);
nor U5662 (N_5662,N_3555,N_475);
and U5663 (N_5663,N_3267,N_931);
or U5664 (N_5664,N_609,N_3473);
nor U5665 (N_5665,N_1129,N_1698);
xnor U5666 (N_5666,N_3173,N_2379);
nand U5667 (N_5667,N_3695,N_4415);
or U5668 (N_5668,N_2964,N_713);
or U5669 (N_5669,N_2492,N_910);
or U5670 (N_5670,N_1963,N_1411);
and U5671 (N_5671,N_1931,N_4646);
or U5672 (N_5672,N_4453,N_981);
xor U5673 (N_5673,N_1587,N_4315);
nand U5674 (N_5674,N_660,N_2590);
nor U5675 (N_5675,N_1158,N_1191);
or U5676 (N_5676,N_3698,N_1478);
or U5677 (N_5677,N_1766,N_3608);
nand U5678 (N_5678,N_2500,N_2400);
nor U5679 (N_5679,N_3405,N_4386);
or U5680 (N_5680,N_4963,N_4575);
nor U5681 (N_5681,N_3995,N_1330);
and U5682 (N_5682,N_2972,N_4318);
nor U5683 (N_5683,N_2987,N_3656);
nor U5684 (N_5684,N_1596,N_3883);
and U5685 (N_5685,N_2583,N_2213);
or U5686 (N_5686,N_1684,N_2488);
or U5687 (N_5687,N_2327,N_325);
nor U5688 (N_5688,N_3869,N_3149);
nand U5689 (N_5689,N_1289,N_3214);
and U5690 (N_5690,N_1597,N_3083);
and U5691 (N_5691,N_2202,N_3599);
and U5692 (N_5692,N_158,N_3830);
or U5693 (N_5693,N_3037,N_1840);
and U5694 (N_5694,N_4502,N_3364);
and U5695 (N_5695,N_2553,N_1473);
and U5696 (N_5696,N_3437,N_2866);
and U5697 (N_5697,N_102,N_3826);
nand U5698 (N_5698,N_3067,N_547);
nand U5699 (N_5699,N_1859,N_4599);
and U5700 (N_5700,N_1881,N_3804);
and U5701 (N_5701,N_1667,N_3482);
and U5702 (N_5702,N_3408,N_4387);
nor U5703 (N_5703,N_4772,N_3147);
nand U5704 (N_5704,N_324,N_1185);
nand U5705 (N_5705,N_2890,N_2423);
nand U5706 (N_5706,N_1973,N_2730);
nand U5707 (N_5707,N_4931,N_1922);
and U5708 (N_5708,N_3106,N_522);
nor U5709 (N_5709,N_3337,N_732);
and U5710 (N_5710,N_4774,N_4156);
or U5711 (N_5711,N_3102,N_1546);
and U5712 (N_5712,N_3048,N_2917);
and U5713 (N_5713,N_3225,N_1122);
and U5714 (N_5714,N_1510,N_4251);
or U5715 (N_5715,N_1932,N_2618);
nand U5716 (N_5716,N_695,N_821);
nor U5717 (N_5717,N_856,N_1836);
nand U5718 (N_5718,N_4226,N_2041);
and U5719 (N_5719,N_2260,N_1580);
and U5720 (N_5720,N_289,N_1181);
or U5721 (N_5721,N_3501,N_3071);
nand U5722 (N_5722,N_2668,N_3176);
or U5723 (N_5723,N_2893,N_135);
nand U5724 (N_5724,N_2530,N_4588);
and U5725 (N_5725,N_3170,N_1720);
or U5726 (N_5726,N_1955,N_767);
or U5727 (N_5727,N_2556,N_3794);
or U5728 (N_5728,N_2680,N_2274);
or U5729 (N_5729,N_3166,N_2187);
nor U5730 (N_5730,N_1226,N_2883);
nor U5731 (N_5731,N_390,N_2949);
nor U5732 (N_5732,N_1388,N_2658);
and U5733 (N_5733,N_1810,N_1690);
nor U5734 (N_5734,N_668,N_819);
and U5735 (N_5735,N_2795,N_3562);
nand U5736 (N_5736,N_4021,N_2290);
nor U5737 (N_5737,N_130,N_481);
nor U5738 (N_5738,N_1458,N_3342);
nor U5739 (N_5739,N_4174,N_2069);
or U5740 (N_5740,N_1153,N_4529);
and U5741 (N_5741,N_3692,N_1427);
and U5742 (N_5742,N_1179,N_1292);
or U5743 (N_5743,N_2566,N_4493);
nor U5744 (N_5744,N_3935,N_404);
nor U5745 (N_5745,N_3903,N_1888);
nor U5746 (N_5746,N_4611,N_2509);
nor U5747 (N_5747,N_3803,N_2121);
nor U5748 (N_5748,N_3095,N_3813);
and U5749 (N_5749,N_728,N_1120);
or U5750 (N_5750,N_3784,N_1718);
and U5751 (N_5751,N_4776,N_1207);
nor U5752 (N_5752,N_3278,N_3725);
or U5753 (N_5753,N_1095,N_772);
nand U5754 (N_5754,N_1015,N_2421);
nor U5755 (N_5755,N_2174,N_3395);
and U5756 (N_5756,N_1101,N_983);
or U5757 (N_5757,N_3817,N_2501);
or U5758 (N_5758,N_4794,N_2816);
xnor U5759 (N_5759,N_293,N_3322);
or U5760 (N_5760,N_1419,N_1645);
nand U5761 (N_5761,N_3162,N_4231);
nand U5762 (N_5762,N_2756,N_3548);
nor U5763 (N_5763,N_3666,N_2383);
nand U5764 (N_5764,N_4373,N_1742);
and U5765 (N_5765,N_4185,N_4999);
nor U5766 (N_5766,N_974,N_4710);
or U5767 (N_5767,N_4035,N_4626);
and U5768 (N_5768,N_3893,N_1266);
nand U5769 (N_5769,N_4258,N_3483);
nand U5770 (N_5770,N_1261,N_1428);
or U5771 (N_5771,N_478,N_223);
nand U5772 (N_5772,N_1463,N_2705);
or U5773 (N_5773,N_1445,N_4033);
nand U5774 (N_5774,N_3298,N_631);
and U5775 (N_5775,N_2718,N_674);
and U5776 (N_5776,N_2104,N_4778);
and U5777 (N_5777,N_4083,N_2192);
or U5778 (N_5778,N_4154,N_3419);
or U5779 (N_5779,N_3375,N_603);
nand U5780 (N_5780,N_4795,N_1322);
nand U5781 (N_5781,N_3181,N_138);
nor U5782 (N_5782,N_4892,N_2360);
nor U5783 (N_5783,N_893,N_1414);
xor U5784 (N_5784,N_4224,N_883);
nand U5785 (N_5785,N_375,N_2352);
nor U5786 (N_5786,N_2619,N_4503);
and U5787 (N_5787,N_4447,N_3142);
nor U5788 (N_5788,N_790,N_4649);
and U5789 (N_5789,N_2422,N_1755);
nor U5790 (N_5790,N_4600,N_8);
and U5791 (N_5791,N_2199,N_3215);
or U5792 (N_5792,N_2224,N_3853);
and U5793 (N_5793,N_2412,N_2947);
nor U5794 (N_5794,N_1764,N_2791);
nor U5795 (N_5795,N_4119,N_3597);
and U5796 (N_5796,N_4750,N_1906);
nand U5797 (N_5797,N_872,N_2543);
and U5798 (N_5798,N_4618,N_2962);
and U5799 (N_5799,N_2160,N_2924);
xor U5800 (N_5800,N_559,N_1921);
nand U5801 (N_5801,N_3256,N_4515);
and U5802 (N_5802,N_1598,N_4268);
and U5803 (N_5803,N_4048,N_2827);
and U5804 (N_5804,N_4129,N_431);
or U5805 (N_5805,N_2456,N_3964);
or U5806 (N_5806,N_4203,N_3187);
or U5807 (N_5807,N_1004,N_569);
nand U5808 (N_5808,N_2152,N_3934);
nand U5809 (N_5809,N_1585,N_2114);
or U5810 (N_5810,N_825,N_424);
and U5811 (N_5811,N_2116,N_3380);
or U5812 (N_5812,N_3414,N_576);
or U5813 (N_5813,N_3749,N_3598);
and U5814 (N_5814,N_2340,N_3909);
nor U5815 (N_5815,N_3021,N_1799);
or U5816 (N_5816,N_1031,N_194);
nor U5817 (N_5817,N_1224,N_4879);
nor U5818 (N_5818,N_881,N_3521);
or U5819 (N_5819,N_4,N_1219);
or U5820 (N_5820,N_2380,N_1244);
and U5821 (N_5821,N_1659,N_2861);
and U5822 (N_5822,N_4122,N_4995);
nand U5823 (N_5823,N_3594,N_276);
nand U5824 (N_5824,N_3422,N_3616);
nand U5825 (N_5825,N_65,N_1382);
nor U5826 (N_5826,N_491,N_3989);
and U5827 (N_5827,N_3712,N_4392);
and U5828 (N_5828,N_2475,N_1678);
nand U5829 (N_5829,N_4051,N_2177);
nor U5830 (N_5830,N_1892,N_2669);
nand U5831 (N_5831,N_3621,N_3716);
nor U5832 (N_5832,N_1144,N_2241);
and U5833 (N_5833,N_2905,N_236);
and U5834 (N_5834,N_2594,N_1246);
or U5835 (N_5835,N_3317,N_926);
nor U5836 (N_5836,N_4932,N_3103);
or U5837 (N_5837,N_2444,N_3927);
nor U5838 (N_5838,N_4086,N_1202);
nand U5839 (N_5839,N_1834,N_4138);
nor U5840 (N_5840,N_2904,N_4466);
and U5841 (N_5841,N_1056,N_2940);
nand U5842 (N_5842,N_2971,N_2775);
nand U5843 (N_5843,N_977,N_2502);
and U5844 (N_5844,N_4460,N_4356);
nor U5845 (N_5845,N_2879,N_3085);
or U5846 (N_5846,N_677,N_1640);
nand U5847 (N_5847,N_3004,N_593);
or U5848 (N_5848,N_2173,N_2291);
nor U5849 (N_5849,N_415,N_3733);
and U5850 (N_5850,N_706,N_1926);
nand U5851 (N_5851,N_2302,N_2433);
or U5852 (N_5852,N_4059,N_1672);
and U5853 (N_5853,N_244,N_4843);
nand U5854 (N_5854,N_4423,N_3518);
or U5855 (N_5855,N_362,N_3227);
nand U5856 (N_5856,N_3442,N_2587);
nor U5857 (N_5857,N_2425,N_1536);
nand U5858 (N_5858,N_389,N_2859);
or U5859 (N_5859,N_4088,N_1331);
nor U5860 (N_5860,N_2445,N_4164);
and U5861 (N_5861,N_709,N_405);
or U5862 (N_5862,N_264,N_1784);
or U5863 (N_5863,N_1563,N_2932);
nor U5864 (N_5864,N_3438,N_1489);
nor U5865 (N_5865,N_3245,N_4924);
and U5866 (N_5866,N_2470,N_3461);
nand U5867 (N_5867,N_3541,N_568);
or U5868 (N_5868,N_4889,N_1511);
nand U5869 (N_5869,N_869,N_192);
or U5870 (N_5870,N_1890,N_1173);
nand U5871 (N_5871,N_1377,N_1040);
nand U5872 (N_5872,N_170,N_3969);
and U5873 (N_5873,N_621,N_216);
nand U5874 (N_5874,N_3189,N_4921);
or U5875 (N_5875,N_1092,N_3432);
and U5876 (N_5876,N_2442,N_3880);
nand U5877 (N_5877,N_3846,N_3620);
and U5878 (N_5878,N_2075,N_958);
and U5879 (N_5879,N_4492,N_3670);
or U5880 (N_5880,N_4790,N_2074);
or U5881 (N_5881,N_606,N_187);
nand U5882 (N_5882,N_3921,N_1035);
nand U5883 (N_5883,N_4305,N_649);
and U5884 (N_5884,N_4528,N_3469);
or U5885 (N_5885,N_1235,N_98);
nor U5886 (N_5886,N_2766,N_1741);
and U5887 (N_5887,N_3552,N_1808);
nand U5888 (N_5888,N_1263,N_1911);
nand U5889 (N_5889,N_2790,N_736);
or U5890 (N_5890,N_3897,N_4631);
or U5891 (N_5891,N_4473,N_698);
nand U5892 (N_5892,N_3940,N_3850);
nand U5893 (N_5893,N_2702,N_3939);
and U5894 (N_5894,N_3126,N_868);
nor U5895 (N_5895,N_3988,N_3186);
nand U5896 (N_5896,N_808,N_1220);
nand U5897 (N_5897,N_2725,N_1852);
nand U5898 (N_5898,N_1332,N_3889);
or U5899 (N_5899,N_1813,N_1505);
nand U5900 (N_5900,N_156,N_4977);
and U5901 (N_5901,N_687,N_4579);
and U5902 (N_5902,N_3504,N_254);
and U5903 (N_5903,N_1751,N_2611);
nand U5904 (N_5904,N_2212,N_3041);
and U5905 (N_5905,N_422,N_2625);
nand U5906 (N_5906,N_95,N_3397);
and U5907 (N_5907,N_119,N_3495);
or U5908 (N_5908,N_3540,N_1703);
or U5909 (N_5909,N_1041,N_2016);
nor U5910 (N_5910,N_3027,N_2928);
and U5911 (N_5911,N_1884,N_804);
nor U5912 (N_5912,N_4041,N_4313);
or U5913 (N_5913,N_2169,N_3839);
and U5914 (N_5914,N_2094,N_1675);
nand U5915 (N_5915,N_4254,N_1476);
nand U5916 (N_5916,N_456,N_884);
and U5917 (N_5917,N_1195,N_3157);
nand U5918 (N_5918,N_4005,N_117);
nand U5919 (N_5919,N_1889,N_2527);
nand U5920 (N_5920,N_752,N_2950);
nand U5921 (N_5921,N_4919,N_747);
and U5922 (N_5922,N_2382,N_2420);
nand U5923 (N_5923,N_3450,N_4097);
xnor U5924 (N_5924,N_2862,N_4233);
or U5925 (N_5925,N_4304,N_250);
nand U5926 (N_5926,N_3713,N_1738);
xnor U5927 (N_5927,N_3980,N_1736);
nand U5928 (N_5928,N_2046,N_1138);
or U5929 (N_5929,N_330,N_2081);
nand U5930 (N_5930,N_4723,N_4902);
or U5931 (N_5931,N_702,N_2641);
or U5932 (N_5932,N_126,N_12);
nand U5933 (N_5933,N_4933,N_3952);
and U5934 (N_5934,N_266,N_4815);
or U5935 (N_5935,N_269,N_2029);
or U5936 (N_5936,N_4010,N_1258);
nor U5937 (N_5937,N_936,N_2923);
and U5938 (N_5938,N_1312,N_4976);
nor U5939 (N_5939,N_3503,N_1305);
nand U5940 (N_5940,N_1688,N_3202);
nor U5941 (N_5941,N_1680,N_1475);
nand U5942 (N_5942,N_4986,N_1376);
and U5943 (N_5943,N_2373,N_1413);
nand U5944 (N_5944,N_661,N_472);
nor U5945 (N_5945,N_2911,N_1441);
or U5946 (N_5946,N_1777,N_2686);
or U5947 (N_5947,N_3508,N_3082);
and U5948 (N_5948,N_690,N_30);
nand U5949 (N_5949,N_4151,N_3867);
nand U5950 (N_5950,N_3232,N_1033);
and U5951 (N_5951,N_917,N_4298);
and U5952 (N_5952,N_413,N_2636);
nor U5953 (N_5953,N_1576,N_4243);
nor U5954 (N_5954,N_3062,N_3259);
and U5955 (N_5955,N_4671,N_3371);
or U5956 (N_5956,N_2396,N_4829);
and U5957 (N_5957,N_1168,N_2386);
nand U5958 (N_5958,N_1662,N_3017);
nand U5959 (N_5959,N_4199,N_3567);
and U5960 (N_5960,N_1524,N_4731);
and U5961 (N_5961,N_2284,N_4434);
nor U5962 (N_5962,N_3945,N_810);
nor U5963 (N_5963,N_1162,N_938);
and U5964 (N_5964,N_2629,N_3236);
nor U5965 (N_5965,N_3558,N_1079);
and U5966 (N_5966,N_4974,N_2564);
or U5967 (N_5967,N_2579,N_814);
and U5968 (N_5968,N_136,N_3705);
or U5969 (N_5969,N_2437,N_357);
and U5970 (N_5970,N_623,N_779);
nand U5971 (N_5971,N_490,N_227);
nand U5972 (N_5972,N_2837,N_3912);
nand U5973 (N_5973,N_3750,N_572);
and U5974 (N_5974,N_2693,N_3358);
nor U5975 (N_5975,N_2008,N_4715);
or U5976 (N_5976,N_955,N_622);
nand U5977 (N_5977,N_506,N_1532);
xor U5978 (N_5978,N_4684,N_3101);
or U5979 (N_5979,N_2648,N_3340);
and U5980 (N_5980,N_4103,N_786);
and U5981 (N_5981,N_602,N_1104);
or U5982 (N_5982,N_3703,N_2559);
or U5983 (N_5983,N_3565,N_1522);
nand U5984 (N_5984,N_1599,N_3273);
or U5985 (N_5985,N_2638,N_2447);
nor U5986 (N_5986,N_1401,N_1634);
and U5987 (N_5987,N_799,N_118);
nand U5988 (N_5988,N_885,N_81);
or U5989 (N_5989,N_2344,N_1471);
nor U5990 (N_5990,N_2525,N_4864);
or U5991 (N_5991,N_4366,N_2054);
or U5992 (N_5992,N_3120,N_1935);
nor U5993 (N_5993,N_1249,N_3757);
or U5994 (N_5994,N_1145,N_3383);
nand U5995 (N_5995,N_681,N_4418);
or U5996 (N_5996,N_4345,N_2623);
or U5997 (N_5997,N_3782,N_1972);
and U5998 (N_5998,N_877,N_1603);
and U5999 (N_5999,N_2995,N_349);
or U6000 (N_6000,N_741,N_4257);
nor U6001 (N_6001,N_142,N_4003);
xor U6002 (N_6002,N_246,N_720);
or U6003 (N_6003,N_376,N_2719);
xor U6004 (N_6004,N_2389,N_208);
nand U6005 (N_6005,N_1989,N_3129);
nand U6006 (N_6006,N_3801,N_4803);
nand U6007 (N_6007,N_4785,N_3012);
and U6008 (N_6008,N_2889,N_2551);
or U6009 (N_6009,N_3374,N_809);
nand U6010 (N_6010,N_1054,N_2754);
or U6011 (N_6011,N_2401,N_182);
nor U6012 (N_6012,N_2161,N_2953);
and U6013 (N_6013,N_4372,N_3297);
nor U6014 (N_6014,N_1641,N_1632);
and U6015 (N_6015,N_4669,N_4901);
and U6016 (N_6016,N_309,N_2218);
nand U6017 (N_6017,N_734,N_4882);
or U6018 (N_6018,N_2894,N_2051);
nor U6019 (N_6019,N_2745,N_1855);
nor U6020 (N_6020,N_1674,N_1154);
or U6021 (N_6021,N_4422,N_2390);
and U6022 (N_6022,N_2039,N_712);
nand U6023 (N_6023,N_1315,N_2426);
xor U6024 (N_6024,N_4499,N_2549);
nor U6025 (N_6025,N_3610,N_4357);
and U6026 (N_6026,N_3068,N_3384);
nand U6027 (N_6027,N_1357,N_1448);
nand U6028 (N_6028,N_2050,N_4709);
and U6029 (N_6029,N_1512,N_1919);
nand U6030 (N_6030,N_3001,N_777);
xor U6031 (N_6031,N_476,N_2770);
and U6032 (N_6032,N_2312,N_710);
nor U6033 (N_6033,N_530,N_4091);
and U6034 (N_6034,N_2055,N_4441);
nand U6035 (N_6035,N_1517,N_1959);
nand U6036 (N_6036,N_1655,N_3456);
and U6037 (N_6037,N_2823,N_3257);
nand U6038 (N_6038,N_2765,N_4577);
and U6039 (N_6039,N_775,N_4265);
and U6040 (N_6040,N_3454,N_2767);
or U6041 (N_6041,N_3303,N_533);
and U6042 (N_6042,N_1559,N_759);
nor U6043 (N_6043,N_1216,N_2494);
nor U6044 (N_6044,N_2458,N_1466);
and U6045 (N_6045,N_2439,N_2079);
nand U6046 (N_6046,N_24,N_3884);
nor U6047 (N_6047,N_4673,N_2743);
and U6048 (N_6048,N_2521,N_1347);
and U6049 (N_6049,N_711,N_4521);
or U6050 (N_6050,N_107,N_866);
and U6051 (N_6051,N_2258,N_2222);
or U6052 (N_6052,N_1618,N_4954);
xor U6053 (N_6053,N_3474,N_4604);
nor U6054 (N_6054,N_175,N_3152);
xnor U6055 (N_6055,N_1939,N_1080);
nor U6056 (N_6056,N_2298,N_1064);
nor U6057 (N_6057,N_2141,N_1714);
and U6058 (N_6058,N_84,N_1409);
or U6059 (N_6059,N_2308,N_1746);
nand U6060 (N_6060,N_392,N_4628);
and U6061 (N_6061,N_4745,N_1198);
and U6062 (N_6062,N_2578,N_3828);
nand U6063 (N_6063,N_750,N_1279);
nand U6064 (N_6064,N_1446,N_4799);
nand U6065 (N_6065,N_1069,N_3975);
nor U6066 (N_6066,N_341,N_620);
nor U6067 (N_6067,N_203,N_2899);
or U6068 (N_6068,N_3699,N_1901);
nor U6069 (N_6069,N_2498,N_2027);
nor U6070 (N_6070,N_3871,N_2985);
or U6071 (N_6071,N_4113,N_1497);
nand U6072 (N_6072,N_563,N_4839);
or U6073 (N_6073,N_3054,N_3044);
and U6074 (N_6074,N_2958,N_4237);
or U6075 (N_6075,N_4848,N_2296);
nor U6076 (N_6076,N_830,N_2131);
nor U6077 (N_6077,N_1802,N_4896);
or U6078 (N_6078,N_3781,N_1761);
nand U6079 (N_6079,N_1116,N_3428);
or U6080 (N_6080,N_2734,N_2558);
or U6081 (N_6081,N_2269,N_529);
or U6082 (N_6082,N_3602,N_1432);
nor U6083 (N_6083,N_4680,N_2785);
nand U6084 (N_6084,N_4153,N_2140);
or U6085 (N_6085,N_888,N_4168);
or U6086 (N_6086,N_1929,N_2175);
nor U6087 (N_6087,N_920,N_3629);
or U6088 (N_6088,N_3911,N_3569);
and U6089 (N_6089,N_3522,N_2634);
xnor U6090 (N_6090,N_3180,N_2413);
and U6091 (N_6091,N_633,N_38);
or U6092 (N_6092,N_2257,N_4625);
nor U6093 (N_6093,N_1953,N_2471);
nand U6094 (N_6094,N_4193,N_1028);
xnor U6095 (N_6095,N_3709,N_4287);
nor U6096 (N_6096,N_3291,N_3583);
and U6097 (N_6097,N_1481,N_2536);
and U6098 (N_6098,N_3216,N_1988);
and U6099 (N_6099,N_909,N_2870);
nand U6100 (N_6100,N_1542,N_1793);
nand U6101 (N_6101,N_2506,N_1009);
and U6102 (N_6102,N_1695,N_1515);
and U6103 (N_6103,N_2084,N_4173);
nand U6104 (N_6104,N_940,N_59);
nand U6105 (N_6105,N_3609,N_1530);
and U6106 (N_6106,N_727,N_2393);
nand U6107 (N_6107,N_1435,N_3638);
nand U6108 (N_6108,N_2469,N_1754);
and U6109 (N_6109,N_497,N_1821);
nand U6110 (N_6110,N_4340,N_762);
and U6111 (N_6111,N_4754,N_3721);
or U6112 (N_6112,N_2671,N_1086);
nor U6113 (N_6113,N_2956,N_2840);
nor U6114 (N_6114,N_3136,N_2044);
or U6115 (N_6115,N_1983,N_4630);
nor U6116 (N_6116,N_4769,N_3660);
or U6117 (N_6117,N_270,N_3635);
nand U6118 (N_6118,N_1337,N_3104);
or U6119 (N_6119,N_812,N_1328);
nand U6120 (N_6120,N_2226,N_2537);
and U6121 (N_6121,N_3689,N_3011);
nand U6122 (N_6122,N_4877,N_1277);
and U6123 (N_6123,N_2772,N_4368);
nand U6124 (N_6124,N_1904,N_2481);
nand U6125 (N_6125,N_3426,N_3642);
or U6126 (N_6126,N_3734,N_3283);
or U6127 (N_6127,N_1824,N_3007);
nor U6128 (N_6128,N_449,N_1062);
and U6129 (N_6129,N_3477,N_2963);
and U6130 (N_6130,N_1971,N_1707);
nand U6131 (N_6131,N_1072,N_2993);
nand U6132 (N_6132,N_2146,N_3188);
nor U6133 (N_6133,N_1547,N_1151);
nand U6134 (N_6134,N_4406,N_3195);
or U6135 (N_6135,N_2487,N_3877);
or U6136 (N_6136,N_4259,N_3841);
nor U6137 (N_6137,N_4210,N_2803);
and U6138 (N_6138,N_1551,N_3193);
or U6139 (N_6139,N_913,N_1947);
nand U6140 (N_6140,N_2603,N_2872);
nor U6141 (N_6141,N_315,N_2406);
nor U6142 (N_6142,N_2436,N_685);
nor U6143 (N_6143,N_3350,N_3458);
and U6144 (N_6144,N_1393,N_2912);
or U6145 (N_6145,N_2021,N_1910);
nand U6146 (N_6146,N_2513,N_2716);
nor U6147 (N_6147,N_2563,N_2148);
nand U6148 (N_6148,N_2703,N_4756);
nand U6149 (N_6149,N_2515,N_2691);
xor U6150 (N_6150,N_1782,N_3807);
nand U6151 (N_6151,N_1934,N_4040);
or U6152 (N_6152,N_2467,N_4309);
and U6153 (N_6153,N_3141,N_1081);
or U6154 (N_6154,N_3226,N_4727);
nand U6155 (N_6155,N_524,N_1447);
and U6156 (N_6156,N_703,N_544);
nor U6157 (N_6157,N_760,N_3553);
nand U6158 (N_6158,N_3207,N_3652);
and U6159 (N_6159,N_4111,N_4525);
or U6160 (N_6160,N_3346,N_1094);
nand U6161 (N_6161,N_4421,N_1708);
nor U6162 (N_6162,N_2097,N_655);
and U6163 (N_6163,N_3615,N_2980);
and U6164 (N_6164,N_2317,N_3306);
or U6165 (N_6165,N_1474,N_1682);
or U6166 (N_6166,N_986,N_4578);
nor U6167 (N_6167,N_2253,N_4558);
xnor U6168 (N_6168,N_1016,N_4562);
or U6169 (N_6169,N_1941,N_2431);
and U6170 (N_6170,N_1902,N_2395);
nand U6171 (N_6171,N_2455,N_1962);
nor U6172 (N_6172,N_2001,N_3857);
or U6173 (N_6173,N_332,N_3987);
nor U6174 (N_6174,N_1338,N_1321);
nand U6175 (N_6175,N_4523,N_3333);
xnor U6176 (N_6176,N_4682,N_3035);
or U6177 (N_6177,N_295,N_4348);
or U6178 (N_6178,N_1143,N_2931);
nor U6179 (N_6179,N_185,N_2873);
nor U6180 (N_6180,N_441,N_1819);
nor U6181 (N_6181,N_1280,N_2771);
nor U6182 (N_6182,N_1558,N_3686);
and U6183 (N_6183,N_1394,N_735);
nor U6184 (N_6184,N_3718,N_1113);
or U6185 (N_6185,N_943,N_2326);
nand U6186 (N_6186,N_1591,N_2085);
xnor U6187 (N_6187,N_1030,N_3123);
and U6188 (N_6188,N_4400,N_2544);
xor U6189 (N_6189,N_484,N_2155);
nor U6190 (N_6190,N_2983,N_2135);
nand U6191 (N_6191,N_3688,N_4494);
nor U6192 (N_6192,N_2297,N_2429);
nor U6193 (N_6193,N_355,N_1296);
nand U6194 (N_6194,N_785,N_3119);
nand U6195 (N_6195,N_2414,N_1343);
xnor U6196 (N_6196,N_4066,N_439);
xnor U6197 (N_6197,N_2617,N_1344);
nor U6198 (N_6198,N_2293,N_3301);
and U6199 (N_6199,N_3365,N_4075);
or U6200 (N_6200,N_4414,N_6);
nor U6201 (N_6201,N_1918,N_3996);
and U6202 (N_6202,N_1696,N_2205);
nand U6203 (N_6203,N_3741,N_1885);
and U6204 (N_6204,N_2363,N_4167);
or U6205 (N_6205,N_2283,N_3720);
or U6206 (N_6206,N_1046,N_2318);
or U6207 (N_6207,N_3455,N_3972);
or U6208 (N_6208,N_3799,N_4842);
and U6209 (N_6209,N_189,N_3900);
nor U6210 (N_6210,N_373,N_3549);
nand U6211 (N_6211,N_1136,N_197);
or U6212 (N_6212,N_2394,N_4079);
and U6213 (N_6213,N_2377,N_3109);
and U6214 (N_6214,N_4935,N_3858);
and U6215 (N_6215,N_26,N_4509);
or U6216 (N_6216,N_4856,N_1389);
nand U6217 (N_6217,N_2752,N_4194);
nand U6218 (N_6218,N_3637,N_27);
nor U6219 (N_6219,N_4025,N_4261);
and U6220 (N_6220,N_143,N_637);
and U6221 (N_6221,N_308,N_4897);
nand U6222 (N_6222,N_3918,N_2333);
nor U6223 (N_6223,N_2110,N_2111);
nand U6224 (N_6224,N_127,N_222);
nor U6225 (N_6225,N_1286,N_3662);
nor U6226 (N_6226,N_4817,N_2416);
nor U6227 (N_6227,N_4032,N_2076);
and U6228 (N_6228,N_536,N_3014);
and U6229 (N_6229,N_75,N_370);
and U6230 (N_6230,N_4470,N_3361);
nor U6231 (N_6231,N_442,N_2042);
or U6232 (N_6232,N_4147,N_1295);
or U6233 (N_6233,N_2979,N_2792);
nand U6234 (N_6234,N_2738,N_2185);
nor U6235 (N_6235,N_843,N_209);
and U6236 (N_6236,N_1715,N_3028);
nor U6237 (N_6237,N_2747,N_2011);
nor U6238 (N_6238,N_3177,N_3919);
xnor U6239 (N_6239,N_1770,N_3128);
or U6240 (N_6240,N_90,N_4637);
xor U6241 (N_6241,N_4276,N_2825);
or U6242 (N_6242,N_2129,N_2571);
nand U6243 (N_6243,N_239,N_2696);
and U6244 (N_6244,N_4326,N_4729);
nand U6245 (N_6245,N_2272,N_4653);
and U6246 (N_6246,N_2221,N_1986);
and U6247 (N_6247,N_3500,N_4944);
nor U6248 (N_6248,N_1210,N_3792);
or U6249 (N_6249,N_3717,N_3563);
and U6250 (N_6250,N_3219,N_4049);
and U6251 (N_6251,N_3570,N_3018);
nand U6252 (N_6252,N_3873,N_4139);
nor U6253 (N_6253,N_1624,N_2519);
or U6254 (N_6254,N_1265,N_2063);
nor U6255 (N_6255,N_2969,N_1807);
and U6256 (N_6256,N_3385,N_3179);
xnor U6257 (N_6257,N_1872,N_4395);
nand U6258 (N_6258,N_2329,N_1508);
or U6259 (N_6259,N_2919,N_382);
and U6260 (N_6260,N_4196,N_4679);
xnor U6261 (N_6261,N_4923,N_3084);
nor U6262 (N_6262,N_860,N_2153);
and U6263 (N_6263,N_2697,N_3753);
or U6264 (N_6264,N_318,N_402);
nand U6265 (N_6265,N_1084,N_1801);
and U6266 (N_6266,N_4559,N_4734);
or U6267 (N_6267,N_2408,N_1553);
nor U6268 (N_6268,N_3892,N_3512);
nor U6269 (N_6269,N_4275,N_1060);
nor U6270 (N_6270,N_3731,N_2198);
nand U6271 (N_6271,N_1061,N_4885);
and U6272 (N_6272,N_514,N_1837);
nor U6273 (N_6273,N_4288,N_4908);
nor U6274 (N_6274,N_4777,N_499);
nor U6275 (N_6275,N_3681,N_3502);
nand U6276 (N_6276,N_1608,N_840);
and U6277 (N_6277,N_4095,N_724);
nand U6278 (N_6278,N_1399,N_201);
or U6279 (N_6279,N_634,N_4597);
nor U6280 (N_6280,N_2268,N_4110);
nor U6281 (N_6281,N_1896,N_4250);
or U6282 (N_6282,N_2101,N_4956);
and U6283 (N_6283,N_1102,N_3160);
or U6284 (N_6284,N_2038,N_57);
nand U6285 (N_6285,N_1586,N_1571);
or U6286 (N_6286,N_2068,N_4766);
nand U6287 (N_6287,N_3034,N_322);
xnor U6288 (N_6288,N_4114,N_848);
or U6289 (N_6289,N_1037,N_4593);
nand U6290 (N_6290,N_3091,N_3772);
nor U6291 (N_6291,N_754,N_3639);
and U6292 (N_6292,N_4285,N_116);
and U6293 (N_6293,N_1371,N_2066);
nor U6294 (N_6294,N_875,N_2476);
and U6295 (N_6295,N_1726,N_1804);
nand U6296 (N_6296,N_1027,N_688);
nor U6297 (N_6297,N_4246,N_4031);
or U6298 (N_6298,N_4364,N_4181);
or U6299 (N_6299,N_1984,N_3413);
or U6300 (N_6300,N_2876,N_890);
and U6301 (N_6301,N_3856,N_4008);
or U6302 (N_6302,N_738,N_1868);
or U6303 (N_6303,N_664,N_4872);
and U6304 (N_6304,N_4082,N_220);
nor U6305 (N_6305,N_1012,N_69);
and U6306 (N_6306,N_281,N_4805);
or U6307 (N_6307,N_1909,N_112);
or U6308 (N_6308,N_1583,N_2099);
or U6309 (N_6309,N_3122,N_2126);
nand U6310 (N_6310,N_3986,N_2461);
nand U6311 (N_6311,N_4607,N_2645);
and U6312 (N_6312,N_1221,N_2799);
or U6313 (N_6313,N_1149,N_4622);
nor U6314 (N_6314,N_2858,N_1730);
and U6315 (N_6315,N_585,N_3250);
or U6316 (N_6316,N_1250,N_2538);
nand U6317 (N_6317,N_2316,N_2127);
or U6318 (N_6318,N_2289,N_3270);
or U6319 (N_6319,N_1067,N_2902);
and U6320 (N_6320,N_583,N_3997);
nand U6321 (N_6321,N_4713,N_2323);
or U6322 (N_6322,N_366,N_2776);
and U6323 (N_6323,N_4809,N_3619);
and U6324 (N_6324,N_3373,N_4937);
nor U6325 (N_6325,N_3732,N_4692);
nand U6326 (N_6326,N_4728,N_1506);
or U6327 (N_6327,N_1232,N_339);
nand U6328 (N_6328,N_1199,N_4409);
nand U6329 (N_6329,N_3536,N_691);
nand U6330 (N_6330,N_3237,N_485);
nor U6331 (N_6331,N_502,N_4907);
nand U6332 (N_6332,N_4755,N_598);
nand U6333 (N_6333,N_4202,N_2955);
nand U6334 (N_6334,N_33,N_3872);
and U6335 (N_6335,N_3404,N_1010);
nand U6336 (N_6336,N_4454,N_4733);
nor U6337 (N_6337,N_3628,N_3372);
and U6338 (N_6338,N_831,N_1854);
and U6339 (N_6339,N_694,N_2897);
nand U6340 (N_6340,N_4946,N_2546);
and U6341 (N_6341,N_4044,N_218);
nand U6342 (N_6342,N_4560,N_4613);
or U6343 (N_6343,N_2585,N_3668);
or U6344 (N_6344,N_3096,N_1299);
nor U6345 (N_6345,N_3331,N_2368);
and U6346 (N_6346,N_3785,N_282);
and U6347 (N_6347,N_2197,N_3966);
or U6348 (N_6348,N_755,N_2243);
and U6349 (N_6349,N_3821,N_1349);
or U6350 (N_6350,N_4598,N_4118);
and U6351 (N_6351,N_965,N_811);
nand U6352 (N_6352,N_4752,N_4297);
or U6353 (N_6353,N_1579,N_587);
nand U6354 (N_6354,N_2233,N_1131);
nand U6355 (N_6355,N_460,N_859);
and U6356 (N_6356,N_4352,N_2635);
nand U6357 (N_6357,N_669,N_616);
or U6358 (N_6358,N_1247,N_3863);
or U6359 (N_6359,N_198,N_1252);
nand U6360 (N_6360,N_4378,N_4887);
and U6361 (N_6361,N_992,N_4026);
nor U6362 (N_6362,N_2685,N_4141);
nand U6363 (N_6363,N_4346,N_2191);
or U6364 (N_6364,N_2954,N_3013);
nand U6365 (N_6365,N_2211,N_1174);
nor U6366 (N_6366,N_2824,N_2062);
nor U6367 (N_6367,N_380,N_4541);
and U6368 (N_6368,N_1023,N_1211);
nor U6369 (N_6369,N_4532,N_2828);
and U6370 (N_6370,N_231,N_3022);
and U6371 (N_6371,N_3353,N_4419);
nand U6372 (N_6372,N_4743,N_4137);
and U6373 (N_6373,N_4410,N_2812);
or U6374 (N_6374,N_1998,N_817);
nand U6375 (N_6375,N_4353,N_997);
nand U6376 (N_6376,N_1978,N_564);
and U6377 (N_6377,N_2270,N_2464);
nand U6378 (N_6378,N_3150,N_2417);
or U6379 (N_6379,N_2036,N_3557);
and U6380 (N_6380,N_2449,N_464);
or U6381 (N_6381,N_243,N_3933);
and U6382 (N_6382,N_2196,N_1404);
nor U6383 (N_6383,N_4840,N_4688);
nor U6384 (N_6384,N_4605,N_3998);
nor U6385 (N_6385,N_4812,N_3719);
nor U6386 (N_6386,N_39,N_582);
nor U6387 (N_6387,N_32,N_835);
and U6388 (N_6388,N_4993,N_4240);
nand U6389 (N_6389,N_1790,N_4273);
nand U6390 (N_6390,N_2575,N_653);
and U6391 (N_6391,N_704,N_1284);
or U6392 (N_6392,N_1020,N_1656);
or U6393 (N_6393,N_1452,N_3984);
nor U6394 (N_6394,N_1022,N_2262);
and U6395 (N_6395,N_4899,N_3239);
nor U6396 (N_6396,N_2434,N_792);
or U6397 (N_6397,N_4444,N_2733);
xor U6398 (N_6398,N_3309,N_2172);
xnor U6399 (N_6399,N_1196,N_4854);
and U6400 (N_6400,N_1774,N_967);
nor U6401 (N_6401,N_887,N_1420);
nand U6402 (N_6402,N_2802,N_4994);
nor U6403 (N_6403,N_4975,N_3002);
nand U6404 (N_6404,N_466,N_411);
or U6405 (N_6405,N_523,N_1743);
nor U6406 (N_6406,N_987,N_2459);
nand U6407 (N_6407,N_2037,N_2599);
or U6408 (N_6408,N_4567,N_629);
or U6409 (N_6409,N_1731,N_53);
and U6410 (N_6410,N_4762,N_2462);
nand U6411 (N_6411,N_1288,N_3947);
nand U6412 (N_6412,N_4209,N_2631);
nor U6413 (N_6413,N_3399,N_148);
or U6414 (N_6414,N_4076,N_272);
and U6415 (N_6415,N_3677,N_604);
or U6416 (N_6416,N_4726,N_617);
nand U6417 (N_6417,N_3825,N_3117);
nand U6418 (N_6418,N_849,N_3217);
xor U6419 (N_6419,N_2732,N_3265);
and U6420 (N_6420,N_638,N_3476);
nand U6421 (N_6421,N_1001,N_4116);
and U6422 (N_6422,N_1654,N_3646);
or U6423 (N_6423,N_1045,N_4248);
nor U6424 (N_6424,N_2193,N_4099);
nand U6425 (N_6425,N_1206,N_25);
nor U6426 (N_6426,N_1771,N_1066);
and U6427 (N_6427,N_2736,N_3032);
xnor U6428 (N_6428,N_74,N_2496);
or U6429 (N_6429,N_4464,N_1400);
or U6430 (N_6430,N_932,N_1233);
or U6431 (N_6431,N_4884,N_1949);
nand U6432 (N_6432,N_3057,N_1106);
or U6433 (N_6433,N_306,N_4225);
nor U6434 (N_6434,N_259,N_4508);
nand U6435 (N_6435,N_898,N_229);
or U6436 (N_6436,N_3042,N_4482);
nand U6437 (N_6437,N_4674,N_3416);
nand U6438 (N_6438,N_789,N_1653);
and U6439 (N_6439,N_2309,N_2256);
nand U6440 (N_6440,N_4548,N_1537);
nor U6441 (N_6441,N_4695,N_80);
and U6442 (N_6442,N_4981,N_4948);
and U6443 (N_6443,N_3601,N_162);
and U6444 (N_6444,N_2710,N_2746);
nor U6445 (N_6445,N_4520,N_2235);
xor U6446 (N_6446,N_2005,N_995);
nor U6447 (N_6447,N_2353,N_4911);
or U6448 (N_6448,N_3748,N_4796);
and U6449 (N_6449,N_716,N_4063);
nand U6450 (N_6450,N_3211,N_3304);
and U6451 (N_6451,N_1496,N_2723);
or U6452 (N_6452,N_715,N_4862);
xnor U6453 (N_6453,N_3092,N_1927);
xor U6454 (N_6454,N_9,N_4379);
and U6455 (N_6455,N_2741,N_1958);
nor U6456 (N_6456,N_4299,N_1499);
nor U6457 (N_6457,N_4904,N_168);
nand U6458 (N_6458,N_1663,N_4290);
and U6459 (N_6459,N_1735,N_1670);
and U6460 (N_6460,N_4703,N_1355);
or U6461 (N_6461,N_1019,N_2757);
and U6462 (N_6462,N_4705,N_2677);
or U6463 (N_6463,N_975,N_4120);
and U6464 (N_6464,N_2887,N_526);
or U6465 (N_6465,N_2139,N_1135);
nand U6466 (N_6466,N_577,N_443);
nand U6467 (N_6467,N_3767,N_2259);
or U6468 (N_6468,N_1572,N_3488);
and U6469 (N_6469,N_3429,N_3393);
or U6470 (N_6470,N_4926,N_4077);
nand U6471 (N_6471,N_639,N_929);
nand U6472 (N_6472,N_1021,N_2035);
and U6473 (N_6473,N_511,N_3762);
nand U6474 (N_6474,N_4950,N_1528);
nand U6475 (N_6475,N_3707,N_2443);
nor U6476 (N_6476,N_1873,N_4517);
nor U6477 (N_6477,N_2898,N_4797);
nand U6478 (N_6478,N_2577,N_4215);
xnor U6479 (N_6479,N_1938,N_833);
nor U6480 (N_6480,N_3539,N_2252);
or U6481 (N_6481,N_4201,N_521);
nor U6482 (N_6482,N_3576,N_1329);
or U6483 (N_6483,N_2440,N_1773);
nand U6484 (N_6484,N_3319,N_580);
and U6485 (N_6485,N_2604,N_914);
nand U6486 (N_6486,N_731,N_2452);
nor U6487 (N_6487,N_3172,N_4719);
nand U6488 (N_6488,N_2220,N_1218);
and U6489 (N_6489,N_3675,N_430);
nor U6490 (N_6490,N_68,N_2610);
nand U6491 (N_6491,N_1239,N_1187);
nor U6492 (N_6492,N_2497,N_3059);
nor U6493 (N_6493,N_589,N_4641);
or U6494 (N_6494,N_2230,N_302);
and U6495 (N_6495,N_1291,N_4439);
nand U6496 (N_6496,N_489,N_3258);
or U6497 (N_6497,N_428,N_605);
nand U6498 (N_6498,N_2189,N_3403);
nor U6499 (N_6499,N_966,N_103);
or U6500 (N_6500,N_3060,N_4823);
and U6501 (N_6501,N_1350,N_2022);
and U6502 (N_6502,N_1269,N_394);
nand U6503 (N_6503,N_2907,N_2489);
nor U6504 (N_6504,N_842,N_4398);
nand U6505 (N_6505,N_1967,N_1723);
and U6506 (N_6506,N_900,N_458);
nor U6507 (N_6507,N_1617,N_4736);
nand U6508 (N_6508,N_3982,N_4661);
nand U6509 (N_6509,N_99,N_4500);
or U6510 (N_6510,N_4253,N_3661);
nor U6511 (N_6511,N_1482,N_2678);
or U6512 (N_6512,N_4382,N_3379);
or U6513 (N_6513,N_3783,N_2982);
nor U6514 (N_6514,N_4316,N_924);
nand U6515 (N_6515,N_45,N_2597);
nand U6516 (N_6516,N_1744,N_853);
and U6517 (N_6517,N_2875,N_3108);
and U6518 (N_6518,N_1780,N_1169);
nor U6519 (N_6519,N_4030,N_501);
and U6520 (N_6520,N_451,N_1433);
xnor U6521 (N_6521,N_3746,N_1676);
xnor U6522 (N_6522,N_2712,N_3596);
or U6523 (N_6523,N_1354,N_4957);
and U6524 (N_6524,N_2867,N_1712);
nor U6525 (N_6525,N_1241,N_928);
nor U6526 (N_6526,N_2106,N_2495);
xor U6527 (N_6527,N_3579,N_3530);
and U6528 (N_6528,N_3263,N_1798);
or U6529 (N_6529,N_344,N_4263);
or U6530 (N_6530,N_4724,N_889);
nand U6531 (N_6531,N_429,N_327);
and U6532 (N_6532,N_4475,N_4431);
nand U6533 (N_6533,N_2709,N_3814);
nand U6534 (N_6534,N_1908,N_1013);
nand U6535 (N_6535,N_4474,N_292);
nand U6536 (N_6536,N_4104,N_1425);
nor U6537 (N_6537,N_4295,N_4841);
nor U6538 (N_6538,N_1887,N_2620);
and U6539 (N_6539,N_4873,N_4811);
nand U6540 (N_6540,N_2246,N_3038);
or U6541 (N_6541,N_2057,N_546);
xnor U6542 (N_6542,N_1114,N_3898);
or U6543 (N_6543,N_3983,N_4553);
or U6544 (N_6544,N_2991,N_2970);
nand U6545 (N_6545,N_2457,N_553);
and U6546 (N_6546,N_2817,N_2622);
nor U6547 (N_6547,N_2391,N_4793);
and U6548 (N_6548,N_496,N_230);
and U6549 (N_6549,N_294,N_3447);
or U6550 (N_6550,N_279,N_3760);
and U6551 (N_6551,N_4476,N_2209);
and U6552 (N_6552,N_1134,N_4065);
nor U6553 (N_6553,N_3674,N_1648);
or U6554 (N_6554,N_820,N_2547);
nand U6555 (N_6555,N_1063,N_4317);
and U6556 (N_6556,N_1800,N_4685);
or U6557 (N_6557,N_1907,N_2601);
nor U6558 (N_6558,N_1981,N_4218);
and U6559 (N_6559,N_4740,N_4833);
or U6560 (N_6560,N_3040,N_1384);
or U6561 (N_6561,N_2067,N_874);
or U6562 (N_6562,N_2561,N_3859);
nor U6563 (N_6563,N_4328,N_262);
nor U6564 (N_6564,N_776,N_3351);
nor U6565 (N_6565,N_4135,N_3974);
and U6566 (N_6566,N_2149,N_1848);
or U6567 (N_6567,N_670,N_4744);
nand U6568 (N_6568,N_4245,N_1605);
nand U6569 (N_6569,N_2937,N_861);
xor U6570 (N_6570,N_1905,N_2811);
nor U6571 (N_6571,N_3053,N_3554);
or U6572 (N_6572,N_3090,N_2782);
and U6573 (N_6573,N_642,N_1137);
and U6574 (N_6574,N_3055,N_2659);
nor U6575 (N_6575,N_3687,N_1930);
or U6576 (N_6576,N_3845,N_1426);
and U6577 (N_6577,N_3357,N_3820);
nand U6578 (N_6578,N_3327,N_1520);
nor U6579 (N_6579,N_745,N_3906);
nand U6580 (N_6580,N_4687,N_2769);
or U6581 (N_6581,N_2607,N_4362);
nand U6582 (N_6582,N_3901,N_1716);
nand U6583 (N_6583,N_933,N_1362);
or U6584 (N_6584,N_1227,N_2349);
xnor U6585 (N_6585,N_4668,N_4002);
or U6586 (N_6586,N_2238,N_3302);
nor U6587 (N_6587,N_2560,N_3496);
nor U6588 (N_6588,N_3197,N_4330);
xnor U6589 (N_6589,N_2742,N_2375);
nand U6590 (N_6590,N_1272,N_1569);
nand U6591 (N_6591,N_4172,N_1380);
nor U6592 (N_6592,N_3253,N_3808);
and U6593 (N_6593,N_4403,N_452);
nand U6594 (N_6594,N_3171,N_3334);
or U6595 (N_6595,N_3324,N_4818);
nor U6596 (N_6596,N_2248,N_238);
and U6597 (N_6597,N_4192,N_1891);
nand U6598 (N_6598,N_2532,N_4102);
nand U6599 (N_6599,N_3905,N_4610);
xnor U6600 (N_6600,N_1396,N_3046);
or U6601 (N_6601,N_4115,N_3167);
or U6602 (N_6602,N_40,N_3930);
or U6603 (N_6603,N_3937,N_4023);
or U6604 (N_6604,N_1514,N_3262);
xnor U6605 (N_6605,N_4927,N_1772);
nand U6606 (N_6606,N_2909,N_2529);
nand U6607 (N_6607,N_3710,N_4804);
nand U6608 (N_6608,N_2182,N_3497);
or U6609 (N_6609,N_3990,N_4836);
or U6610 (N_6610,N_1368,N_286);
or U6611 (N_6611,N_1171,N_3837);
or U6612 (N_6612,N_1664,N_3355);
nor U6613 (N_6613,N_4319,N_1869);
xor U6614 (N_6614,N_2446,N_4883);
and U6615 (N_6615,N_3100,N_1635);
or U6616 (N_6616,N_4266,N_4970);
nand U6617 (N_6617,N_1406,N_2541);
nor U6618 (N_6618,N_2647,N_647);
or U6619 (N_6619,N_4046,N_2130);
nand U6620 (N_6620,N_1990,N_1055);
nand U6621 (N_6621,N_4510,N_4758);
and U6622 (N_6622,N_1737,N_3835);
and U6623 (N_6623,N_4140,N_4700);
and U6624 (N_6624,N_2343,N_919);
nand U6625 (N_6625,N_4574,N_766);
and U6626 (N_6626,N_4191,N_1783);
nor U6627 (N_6627,N_4894,N_4732);
or U6628 (N_6628,N_2348,N_1966);
and U6629 (N_6629,N_417,N_3546);
and U6630 (N_6630,N_2706,N_1333);
or U6631 (N_6631,N_4301,N_395);
nand U6632 (N_6632,N_4338,N_4960);
nand U6633 (N_6633,N_2087,N_3284);
and U6634 (N_6634,N_520,N_3588);
nor U6635 (N_6635,N_1180,N_314);
or U6636 (N_6636,N_4781,N_2404);
and U6637 (N_6637,N_1341,N_2592);
nand U6638 (N_6638,N_4262,N_190);
nor U6639 (N_6639,N_850,N_3791);
nor U6640 (N_6640,N_2781,N_225);
nor U6641 (N_6641,N_4938,N_3223);
and U6642 (N_6642,N_2856,N_437);
and U6643 (N_6643,N_4401,N_2926);
nor U6644 (N_6644,N_3944,N_3098);
and U6645 (N_6645,N_3514,N_3363);
nor U6646 (N_6646,N_2402,N_4656);
nand U6647 (N_6647,N_1699,N_487);
or U6648 (N_6648,N_3755,N_1059);
nor U6649 (N_6649,N_2424,N_672);
nor U6650 (N_6650,N_839,N_2615);
nor U6651 (N_6651,N_1805,N_4133);
and U6652 (N_6652,N_3064,N_4991);
or U6653 (N_6653,N_1594,N_4869);
or U6654 (N_6654,N_2518,N_948);
or U6655 (N_6655,N_4753,N_4531);
nand U6656 (N_6656,N_4561,N_436);
xnor U6657 (N_6657,N_500,N_1629);
nand U6658 (N_6658,N_2115,N_4011);
nor U6659 (N_6659,N_17,N_3005);
nand U6660 (N_6660,N_78,N_2064);
or U6661 (N_6661,N_2228,N_1461);
or U6662 (N_6662,N_21,N_3079);
xor U6663 (N_6663,N_610,N_3844);
nor U6664 (N_6664,N_4308,N_1595);
or U6665 (N_6665,N_2482,N_2739);
nand U6666 (N_6666,N_2667,N_4408);
or U6667 (N_6667,N_2060,N_1273);
nor U6668 (N_6668,N_3233,N_4979);
nand U6669 (N_6669,N_578,N_882);
or U6670 (N_6670,N_1057,N_2646);
or U6671 (N_6671,N_1146,N_3268);
or U6672 (N_6672,N_4891,N_3963);
nor U6673 (N_6673,N_561,N_4616);
or U6674 (N_6674,N_2581,N_3678);
xor U6675 (N_6675,N_321,N_1643);
nand U6676 (N_6676,N_968,N_2934);
nor U6677 (N_6677,N_4880,N_2362);
and U6678 (N_6678,N_4117,N_4467);
nand U6679 (N_6679,N_114,N_625);
nand U6680 (N_6680,N_249,N_4587);
nand U6681 (N_6681,N_4056,N_1794);
nand U6682 (N_6682,N_558,N_2337);
or U6683 (N_6683,N_4081,N_4939);
nand U6684 (N_6684,N_2300,N_4183);
nand U6685 (N_6685,N_4438,N_1842);
xor U6686 (N_6686,N_2567,N_3833);
or U6687 (N_6687,N_2942,N_4549);
nor U6688 (N_6688,N_1987,N_2717);
nor U6689 (N_6689,N_555,N_4922);
or U6690 (N_6690,N_791,N_4582);
and U6691 (N_6691,N_3946,N_1008);
or U6692 (N_6692,N_4169,N_4256);
and U6693 (N_6693,N_3796,N_2453);
or U6694 (N_6694,N_2304,N_2210);
and U6695 (N_6695,N_4825,N_1644);
nor U6696 (N_6696,N_1111,N_4150);
or U6697 (N_6697,N_2548,N_2366);
nand U6698 (N_6698,N_1870,N_3078);
and U6699 (N_6699,N_2376,N_4424);
and U6700 (N_6700,N_2888,N_4284);
or U6701 (N_6701,N_3537,N_2098);
nor U6702 (N_6702,N_3836,N_4100);
nand U6703 (N_6703,N_2321,N_171);
or U6704 (N_6704,N_4396,N_3295);
and U6705 (N_6705,N_1996,N_643);
nand U6706 (N_6706,N_4706,N_4069);
nor U6707 (N_6707,N_818,N_2764);
and U6708 (N_6708,N_3520,N_2589);
nand U6709 (N_6709,N_1006,N_4526);
and U6710 (N_6710,N_2451,N_42);
and U6711 (N_6711,N_1391,N_1438);
and U6712 (N_6712,N_1933,N_2999);
or U6713 (N_6713,N_624,N_4962);
nand U6714 (N_6714,N_2156,N_3114);
and U6715 (N_6715,N_150,N_2557);
xor U6716 (N_6716,N_410,N_434);
or U6717 (N_6717,N_1623,N_4469);
and U6718 (N_6718,N_1916,N_1850);
xnor U6719 (N_6719,N_4426,N_1611);
nand U6720 (N_6720,N_1507,N_3879);
or U6721 (N_6721,N_651,N_4322);
nor U6722 (N_6722,N_903,N_2805);
nor U6723 (N_6723,N_795,N_4170);
nand U6724 (N_6724,N_3507,N_4875);
and U6725 (N_6725,N_532,N_528);
nand U6726 (N_6726,N_3878,N_2033);
and U6727 (N_6727,N_2078,N_1003);
nor U6728 (N_6728,N_4998,N_708);
nand U6729 (N_6729,N_1494,N_2477);
nand U6730 (N_6730,N_3043,N_4853);
nor U6731 (N_6731,N_937,N_994);
nor U6732 (N_6732,N_4775,N_1190);
and U6733 (N_6733,N_3208,N_345);
or U6734 (N_6734,N_4197,N_3876);
and U6735 (N_6735,N_3183,N_3411);
nor U6736 (N_6736,N_3,N_4242);
nand U6737 (N_6737,N_4936,N_2656);
or U6738 (N_6738,N_2959,N_2180);
and U6739 (N_6739,N_88,N_3745);
nand U6740 (N_6740,N_971,N_2570);
or U6741 (N_6741,N_4371,N_2490);
nand U6742 (N_6742,N_867,N_1051);
or U6743 (N_6743,N_128,N_145);
or U6744 (N_6744,N_3510,N_4504);
nand U6745 (N_6745,N_444,N_2147);
nand U6746 (N_6746,N_4497,N_3774);
xnor U6747 (N_6747,N_2842,N_432);
and U6748 (N_6748,N_3247,N_1088);
and U6749 (N_6749,N_274,N_4078);
xor U6750 (N_6750,N_608,N_2355);
or U6751 (N_6751,N_4061,N_1575);
nor U6752 (N_6752,N_2996,N_1166);
nand U6753 (N_6753,N_3916,N_4134);
nor U6754 (N_6754,N_4693,N_2120);
xor U6755 (N_6755,N_4478,N_782);
nor U6756 (N_6756,N_4542,N_3288);
or U6757 (N_6757,N_20,N_4214);
nor U6758 (N_6758,N_4683,N_4361);
and U6759 (N_6759,N_334,N_301);
or U6760 (N_6760,N_237,N_1636);
nand U6761 (N_6761,N_3135,N_2514);
nor U6762 (N_6762,N_3308,N_2092);
and U6763 (N_6763,N_1108,N_1011);
nor U6764 (N_6764,N_982,N_414);
nand U6765 (N_6765,N_1502,N_109);
and U6766 (N_6766,N_4022,N_548);
or U6767 (N_6767,N_4592,N_2675);
or U6768 (N_6768,N_141,N_85);
nor U6769 (N_6769,N_426,N_635);
or U6770 (N_6770,N_2637,N_4334);
nor U6771 (N_6771,N_2688,N_640);
nor U6772 (N_6772,N_1152,N_4007);
and U6773 (N_6773,N_744,N_2245);
or U6774 (N_6774,N_4080,N_956);
or U6775 (N_6775,N_3163,N_542);
or U6776 (N_6776,N_3571,N_4351);
and U6777 (N_6777,N_2320,N_4020);
nand U6778 (N_6778,N_1378,N_3069);
or U6779 (N_6779,N_3459,N_990);
and U6780 (N_6780,N_3847,N_3928);
and U6781 (N_6781,N_4947,N_255);
nor U6782 (N_6782,N_4286,N_2441);
nor U6783 (N_6783,N_403,N_696);
nand U6784 (N_6784,N_4751,N_1846);
nand U6785 (N_6785,N_846,N_3607);
nor U6786 (N_6786,N_2822,N_1845);
nor U6787 (N_6787,N_2751,N_3590);
and U6788 (N_6788,N_1182,N_4681);
nand U6789 (N_6789,N_139,N_2819);
nand U6790 (N_6790,N_4783,N_2990);
nand U6791 (N_6791,N_2555,N_3636);
or U6792 (N_6792,N_174,N_630);
nand U6793 (N_6793,N_1439,N_498);
nor U6794 (N_6794,N_4620,N_3088);
or U6795 (N_6795,N_4909,N_3204);
nand U6796 (N_6796,N_4360,N_166);
nand U6797 (N_6797,N_4632,N_1381);
nor U6798 (N_6798,N_2698,N_4367);
xnor U6799 (N_6799,N_3915,N_4216);
nand U6800 (N_6800,N_3823,N_2986);
and U6801 (N_6801,N_3559,N_4485);
and U6802 (N_6802,N_2768,N_261);
nor U6803 (N_6803,N_2052,N_2517);
or U6804 (N_6804,N_3490,N_3305);
and U6805 (N_6805,N_2989,N_1132);
and U6806 (N_6806,N_1186,N_3499);
or U6807 (N_6807,N_581,N_4335);
and U6808 (N_6808,N_858,N_717);
nand U6809 (N_6809,N_3282,N_1915);
xor U6810 (N_6810,N_3778,N_1200);
and U6811 (N_6811,N_427,N_591);
and U6812 (N_6812,N_1300,N_3178);
or U6813 (N_6813,N_2178,N_4645);
nor U6814 (N_6814,N_4084,N_4506);
or U6815 (N_6815,N_495,N_2374);
or U6816 (N_6816,N_2311,N_1170);
or U6817 (N_6817,N_4547,N_3036);
nand U6818 (N_6818,N_1309,N_1449);
nand U6819 (N_6819,N_137,N_2628);
nor U6820 (N_6820,N_1970,N_4009);
and U6821 (N_6821,N_1616,N_3231);
nand U6822 (N_6822,N_3580,N_3645);
nand U6823 (N_6823,N_2438,N_224);
xor U6824 (N_6824,N_4057,N_1431);
or U6825 (N_6825,N_3626,N_4436);
and U6826 (N_6826,N_3943,N_4296);
nand U6827 (N_6827,N_3417,N_396);
or U6828 (N_6828,N_2998,N_3957);
nand U6829 (N_6829,N_658,N_729);
and U6830 (N_6830,N_3449,N_2831);
and U6831 (N_6831,N_169,N_1803);
and U6832 (N_6832,N_3547,N_596);
xnor U6833 (N_6833,N_3951,N_918);
nor U6834 (N_6834,N_331,N_4644);
and U6835 (N_6835,N_2465,N_2200);
and U6836 (N_6836,N_4420,N_3528);
or U6837 (N_6837,N_4180,N_4006);
or U6838 (N_6838,N_976,N_768);
nand U6839 (N_6839,N_2794,N_739);
nand U6840 (N_6840,N_2966,N_2013);
and U6841 (N_6841,N_2103,N_2299);
xnor U6842 (N_6842,N_3655,N_2692);
nand U6843 (N_6843,N_4280,N_2325);
nand U6844 (N_6844,N_4255,N_1677);
and U6845 (N_6845,N_1039,N_588);
and U6846 (N_6846,N_3556,N_599);
or U6847 (N_6847,N_329,N_1436);
nor U6848 (N_6848,N_960,N_3516);
or U6849 (N_6849,N_4146,N_864);
or U6850 (N_6850,N_1826,N_1781);
or U6851 (N_6851,N_3427,N_3424);
or U6852 (N_6852,N_1760,N_1518);
nor U6853 (N_6853,N_550,N_2372);
xor U6854 (N_6854,N_3318,N_4358);
nor U6855 (N_6855,N_4232,N_667);
nor U6856 (N_6856,N_4012,N_4015);
nor U6857 (N_6857,N_1443,N_3736);
xnor U6858 (N_6858,N_4227,N_64);
and U6859 (N_6859,N_758,N_3003);
nand U6860 (N_6860,N_2749,N_3985);
and U6861 (N_6861,N_1895,N_4471);
nor U6862 (N_6862,N_802,N_2665);
nor U6863 (N_6863,N_3213,N_3000);
nor U6864 (N_6864,N_2171,N_180);
nand U6865 (N_6865,N_3842,N_2626);
and U6866 (N_6866,N_4742,N_510);
or U6867 (N_6867,N_1234,N_648);
nand U6868 (N_6868,N_2660,N_3978);
nor U6869 (N_6869,N_1271,N_3010);
or U6870 (N_6870,N_3398,N_1440);
and U6871 (N_6871,N_4996,N_1248);
and U6872 (N_6872,N_346,N_4206);
nand U6873 (N_6873,N_3625,N_4810);
nand U6874 (N_6874,N_234,N_1486);
nand U6875 (N_6875,N_468,N_3742);
or U6876 (N_6876,N_378,N_1814);
or U6877 (N_6877,N_4545,N_4292);
nor U6878 (N_6878,N_1706,N_2545);
or U6879 (N_6879,N_2851,N_470);
xor U6880 (N_6880,N_447,N_4903);
nand U6881 (N_6881,N_1105,N_1325);
and U6882 (N_6882,N_3908,N_1320);
and U6883 (N_6883,N_1209,N_3648);
nand U6884 (N_6884,N_4721,N_645);
or U6885 (N_6885,N_796,N_1123);
or U6886 (N_6886,N_2936,N_2342);
nand U6887 (N_6887,N_4429,N_612);
nor U6888 (N_6888,N_2010,N_7);
or U6889 (N_6889,N_1637,N_3338);
nand U6890 (N_6890,N_3377,N_1231);
or U6891 (N_6891,N_3435,N_3191);
or U6892 (N_6892,N_4090,N_1348);
xnor U6893 (N_6893,N_1416,N_70);
and U6894 (N_6894,N_1631,N_1633);
nor U6895 (N_6895,N_2351,N_4000);
nand U6896 (N_6896,N_4437,N_2728);
nor U6897 (N_6897,N_372,N_41);
and U6898 (N_6898,N_3613,N_2460);
nand U6899 (N_6899,N_3400,N_4412);
nor U6900 (N_6900,N_195,N_3543);
or U6901 (N_6901,N_1500,N_3524);
nor U6902 (N_6902,N_1843,N_1076);
or U6903 (N_6903,N_4591,N_880);
and U6904 (N_6904,N_2948,N_4136);
and U6905 (N_6905,N_2914,N_505);
nor U6906 (N_6906,N_4178,N_3848);
and U6907 (N_6907,N_1792,N_3487);
or U6908 (N_6908,N_374,N_2981);
nand U6909 (N_6909,N_1201,N_248);
nand U6910 (N_6910,N_2885,N_1847);
and U6911 (N_6911,N_1184,N_1818);
or U6912 (N_6912,N_984,N_232);
nor U6913 (N_6913,N_2285,N_200);
nand U6914 (N_6914,N_2338,N_2695);
and U6915 (N_6915,N_3827,N_1503);
or U6916 (N_6916,N_4281,N_4691);
and U6917 (N_6917,N_1721,N_3875);
and U6918 (N_6918,N_662,N_3182);
and U6919 (N_6919,N_2505,N_2407);
nor U6920 (N_6920,N_3994,N_1085);
or U6921 (N_6921,N_1582,N_1776);
or U6922 (N_6922,N_4325,N_1351);
or U6923 (N_6923,N_2762,N_1541);
or U6924 (N_6924,N_3381,N_1797);
nor U6925 (N_6925,N_493,N_3443);
or U6926 (N_6926,N_3138,N_4920);
and U6927 (N_6927,N_823,N_1924);
nor U6928 (N_6928,N_4130,N_3464);
xnor U6929 (N_6929,N_3714,N_4407);
and U6930 (N_6930,N_1758,N_2639);
nand U6931 (N_6931,N_1994,N_2208);
nand U6932 (N_6932,N_838,N_3751);
nand U6933 (N_6933,N_801,N_4332);
xnor U6934 (N_6934,N_597,N_2134);
and U6935 (N_6935,N_1327,N_4402);
nor U6936 (N_6936,N_517,N_1883);
and U6937 (N_6937,N_467,N_1032);
or U6938 (N_6938,N_2944,N_3931);
nand U6939 (N_6939,N_4105,N_4533);
nand U6940 (N_6940,N_3606,N_1533);
nor U6941 (N_6941,N_1747,N_3478);
or U6942 (N_6942,N_4786,N_4554);
or U6943 (N_6943,N_2881,N_2214);
nor U6944 (N_6944,N_4004,N_1969);
and U6945 (N_6945,N_4127,N_1408);
nand U6946 (N_6946,N_4819,N_1685);
nand U6947 (N_6947,N_3274,N_3704);
nand U6948 (N_6948,N_36,N_805);
and U6949 (N_6949,N_1089,N_4487);
and U6950 (N_6950,N_2405,N_4555);
nand U6951 (N_6951,N_3630,N_2586);
nor U6952 (N_6952,N_23,N_3604);
or U6953 (N_6953,N_2273,N_961);
and U6954 (N_6954,N_2403,N_4961);
and U6955 (N_6955,N_3603,N_4496);
and U6956 (N_6956,N_2627,N_2031);
nor U6957 (N_6957,N_1387,N_3956);
nor U6958 (N_6958,N_2684,N_4207);
and U6959 (N_6959,N_3822,N_3896);
nand U6960 (N_6960,N_4486,N_1894);
nor U6961 (N_6961,N_4013,N_181);
or U6962 (N_6962,N_2231,N_959);
nand U6963 (N_6963,N_855,N_2735);
and U6964 (N_6964,N_3154,N_110);
nand U6965 (N_6965,N_140,N_4272);
nand U6966 (N_6966,N_4949,N_851);
and U6967 (N_6967,N_3611,N_942);
and U6968 (N_6968,N_656,N_778);
nand U6969 (N_6969,N_1429,N_2124);
nand U6970 (N_6970,N_4865,N_2484);
or U6971 (N_6971,N_614,N_2255);
and U6972 (N_6972,N_2927,N_123);
nand U6973 (N_6973,N_894,N_2878);
and U6974 (N_6974,N_3240,N_1968);
and U6975 (N_6975,N_3752,N_483);
or U6976 (N_6976,N_1490,N_2485);
nor U6977 (N_6977,N_280,N_2301);
nand U6978 (N_6978,N_3391,N_2573);
nor U6979 (N_6979,N_226,N_2089);
nand U6980 (N_6980,N_3722,N_1732);
nor U6981 (N_6981,N_2206,N_1980);
nor U6982 (N_6982,N_4188,N_2984);
or U6983 (N_6983,N_2204,N_2884);
nor U6984 (N_6984,N_149,N_253);
or U6985 (N_6985,N_2263,N_4953);
nand U6986 (N_6986,N_71,N_131);
and U6987 (N_6987,N_1762,N_433);
nor U6988 (N_6988,N_3623,N_1692);
xor U6989 (N_6989,N_1992,N_3310);
and U6990 (N_6990,N_3973,N_2083);
and U6991 (N_6991,N_4344,N_1188);
or U6992 (N_6992,N_2225,N_1127);
and U6993 (N_6993,N_4941,N_1649);
nor U6994 (N_6994,N_743,N_4235);
or U6995 (N_6995,N_4690,N_4916);
nor U6996 (N_6996,N_2357,N_1326);
and U6997 (N_6997,N_3743,N_1048);
nor U6998 (N_6998,N_5,N_1043);
nand U6999 (N_6999,N_4267,N_1858);
nor U7000 (N_7000,N_3354,N_3653);
nand U7001 (N_7001,N_3809,N_176);
and U7002 (N_7002,N_4126,N_408);
nand U7003 (N_7003,N_1230,N_2236);
nor U7004 (N_7004,N_3747,N_4606);
nand U7005 (N_7005,N_4458,N_205);
or U7006 (N_7006,N_196,N_3058);
nand U7007 (N_7007,N_2651,N_993);
and U7008 (N_7008,N_781,N_1385);
nor U7009 (N_7009,N_4516,N_2335);
nor U7010 (N_7010,N_96,N_1464);
nor U7011 (N_7011,N_3448,N_3118);
and U7012 (N_7012,N_3362,N_384);
nand U7013 (N_7013,N_1161,N_1578);
or U7014 (N_7014,N_4038,N_3446);
nor U7015 (N_7015,N_4788,N_3475);
or U7016 (N_7016,N_3575,N_4417);
nor U7017 (N_7017,N_3523,N_1238);
nor U7018 (N_7018,N_4651,N_2662);
nand U7019 (N_7019,N_4686,N_290);
nand U7020 (N_7020,N_3815,N_2288);
or U7021 (N_7021,N_3143,N_2938);
nor U7022 (N_7022,N_4929,N_3049);
and U7023 (N_7023,N_1509,N_824);
or U7024 (N_7024,N_4573,N_619);
and U7025 (N_7025,N_2295,N_291);
nand U7026 (N_7026,N_1430,N_1694);
nor U7027 (N_7027,N_4312,N_2910);
nor U7028 (N_7028,N_3802,N_3229);
or U7029 (N_7029,N_2813,N_2056);
or U7030 (N_7030,N_1498,N_63);
or U7031 (N_7031,N_3885,N_1882);
nor U7032 (N_7032,N_4067,N_678);
and U7033 (N_7033,N_2398,N_4720);
nand U7034 (N_7034,N_4062,N_594);
and U7035 (N_7035,N_52,N_3134);
nor U7036 (N_7036,N_2512,N_82);
nor U7037 (N_7037,N_438,N_480);
or U7038 (N_7038,N_3696,N_3938);
nor U7039 (N_7039,N_1942,N_386);
nand U7040 (N_7040,N_2278,N_4278);
nor U7041 (N_7041,N_1167,N_3676);
nand U7042 (N_7042,N_338,N_3234);
nand U7043 (N_7043,N_1526,N_3489);
or U7044 (N_7044,N_4072,N_847);
and U7045 (N_7045,N_3693,N_2419);
nor U7046 (N_7046,N_1453,N_3824);
nand U7047 (N_7047,N_2713,N_4050);
and U7048 (N_7048,N_571,N_686);
nor U7049 (N_7049,N_4391,N_4241);
or U7050 (N_7050,N_3967,N_3203);
or U7051 (N_7051,N_4098,N_2874);
or U7052 (N_7052,N_1256,N_1422);
or U7053 (N_7053,N_4534,N_2935);
or U7054 (N_7054,N_4886,N_3683);
or U7055 (N_7055,N_3292,N_2588);
or U7056 (N_7056,N_2882,N_2034);
nor U7057 (N_7057,N_3950,N_1752);
nor U7058 (N_7058,N_1465,N_693);
nand U7059 (N_7059,N_2786,N_4239);
nor U7060 (N_7060,N_455,N_77);
or U7061 (N_7061,N_1521,N_1128);
or U7062 (N_7062,N_2796,N_1251);
nor U7063 (N_7063,N_2201,N_4568);
nand U7064 (N_7064,N_4830,N_4219);
nand U7065 (N_7065,N_199,N_3672);
and U7066 (N_7066,N_3564,N_1538);
nand U7067 (N_7067,N_2520,N_4861);
and U7068 (N_7068,N_4784,N_3605);
or U7069 (N_7069,N_3255,N_1189);
nand U7070 (N_7070,N_4377,N_2358);
nand U7071 (N_7071,N_2857,N_2303);
or U7072 (N_7072,N_3194,N_697);
or U7073 (N_7073,N_3260,N_316);
and U7074 (N_7074,N_3560,N_2491);
nand U7075 (N_7075,N_352,N_2903);
and U7076 (N_7076,N_879,N_4698);
nand U7077 (N_7077,N_1820,N_969);
nor U7078 (N_7078,N_3465,N_1833);
nor U7079 (N_7079,N_1483,N_2820);
or U7080 (N_7080,N_3631,N_287);
nor U7081 (N_7081,N_3600,N_4166);
xor U7082 (N_7082,N_448,N_2973);
nor U7083 (N_7083,N_3773,N_3955);
or U7084 (N_7084,N_4966,N_4730);
and U7085 (N_7085,N_2510,N_4385);
and U7086 (N_7086,N_3074,N_351);
nand U7087 (N_7087,N_4374,N_2030);
or U7088 (N_7088,N_3198,N_1523);
or U7089 (N_7089,N_4990,N_1147);
and U7090 (N_7090,N_1442,N_2179);
nand U7091 (N_7091,N_4369,N_3272);
nor U7092 (N_7092,N_2900,N_2328);
or U7093 (N_7093,N_3392,N_4511);
nand U7094 (N_7094,N_1767,N_4073);
and U7095 (N_7095,N_4222,N_4427);
xnor U7096 (N_7096,N_3851,N_3115);
and U7097 (N_7097,N_4851,N_1527);
or U7098 (N_7098,N_1830,N_4890);
nand U7099 (N_7099,N_3669,N_1899);
nand U7100 (N_7100,N_4397,N_4289);
and U7101 (N_7101,N_2324,N_4513);
nor U7102 (N_7102,N_1178,N_3881);
and U7103 (N_7103,N_518,N_2780);
nor U7104 (N_7104,N_2793,N_2108);
nand U7105 (N_7105,N_3261,N_4544);
or U7106 (N_7106,N_1651,N_4489);
nor U7107 (N_7107,N_1719,N_1529);
or U7108 (N_7108,N_474,N_1303);
and U7109 (N_7109,N_4331,N_2968);
or U7110 (N_7110,N_3818,N_4676);
nor U7111 (N_7111,N_4393,N_3805);
nor U7112 (N_7112,N_2043,N_3316);
nor U7113 (N_7113,N_4070,N_2448);
nand U7114 (N_7114,N_206,N_663);
nand U7115 (N_7115,N_3581,N_1613);
and U7116 (N_7116,N_4670,N_4765);
nor U7117 (N_7117,N_783,N_2522);
and U7118 (N_7118,N_1243,N_925);
nor U7119 (N_7119,N_3209,N_2112);
and U7120 (N_7120,N_2534,N_4792);
or U7121 (N_7121,N_2,N_1621);
and U7122 (N_7122,N_2168,N_822);
or U7123 (N_7123,N_4279,N_212);
and U7124 (N_7124,N_4306,N_3133);
and U7125 (N_7125,N_2242,N_4264);
and U7126 (N_7126,N_172,N_1025);
nand U7127 (N_7127,N_2621,N_4910);
or U7128 (N_7128,N_1268,N_4918);
nand U7129 (N_7129,N_876,N_4089);
or U7130 (N_7130,N_425,N_2869);
or U7131 (N_7131,N_3155,N_575);
and U7132 (N_7132,N_66,N_4629);
nor U7133 (N_7133,N_3370,N_354);
xor U7134 (N_7134,N_340,N_1686);
nor U7135 (N_7135,N_1307,N_3077);
nand U7136 (N_7136,N_4760,N_3976);
and U7137 (N_7137,N_1372,N_3634);
nand U7138 (N_7138,N_2133,N_3788);
and U7139 (N_7139,N_277,N_2644);
or U7140 (N_7140,N_3235,N_1240);
nor U7141 (N_7141,N_3595,N_2720);
nor U7142 (N_7142,N_973,N_446);
or U7143 (N_7143,N_1614,N_4260);
or U7144 (N_7144,N_1954,N_4327);
or U7145 (N_7145,N_2860,N_263);
nor U7146 (N_7146,N_1519,N_2568);
and U7147 (N_7147,N_2814,N_4718);
and U7148 (N_7148,N_4969,N_1165);
or U7149 (N_7149,N_2118,N_486);
nor U7150 (N_7150,N_2123,N_3230);
and U7151 (N_7151,N_1029,N_1367);
or U7152 (N_7152,N_4945,N_3694);
nor U7153 (N_7153,N_2122,N_381);
or U7154 (N_7154,N_108,N_1748);
nor U7155 (N_7155,N_3444,N_4071);
and U7156 (N_7156,N_1564,N_3390);
nand U7157 (N_7157,N_1757,N_2540);
nand U7158 (N_7158,N_2331,N_2798);
nand U7159 (N_7159,N_1627,N_4934);
nand U7160 (N_7160,N_3061,N_4570);
nand U7161 (N_7161,N_1795,N_2679);
nor U7162 (N_7162,N_3739,N_3481);
nand U7163 (N_7163,N_2580,N_1038);
nand U7164 (N_7164,N_4204,N_3941);
nand U7165 (N_7165,N_3840,N_4906);
and U7166 (N_7166,N_146,N_2188);
nor U7167 (N_7167,N_3145,N_509);
nand U7168 (N_7168,N_4413,N_49);
nor U7169 (N_7169,N_2758,N_4971);
nand U7170 (N_7170,N_4749,N_829);
or U7171 (N_7171,N_4291,N_4845);
and U7172 (N_7172,N_273,N_2086);
nand U7173 (N_7173,N_535,N_4175);
or U7174 (N_7174,N_4449,N_4837);
nor U7175 (N_7175,N_213,N_353);
or U7176 (N_7176,N_1619,N_3299);
nand U7177 (N_7177,N_2266,N_949);
nand U7178 (N_7178,N_4988,N_2891);
nor U7179 (N_7179,N_4053,N_1853);
nand U7180 (N_7180,N_463,N_4619);
or U7181 (N_7181,N_3647,N_2650);
nor U7182 (N_7182,N_2591,N_4430);
nor U7183 (N_7183,N_1574,N_3094);
nor U7184 (N_7184,N_2797,N_4303);
nand U7185 (N_7185,N_4455,N_1661);
nand U7186 (N_7186,N_3913,N_4602);
nand U7187 (N_7187,N_251,N_3244);
or U7188 (N_7188,N_1835,N_4343);
or U7189 (N_7189,N_1098,N_3708);
nand U7190 (N_7190,N_1100,N_2701);
and U7191 (N_7191,N_2244,N_1701);
and U7192 (N_7192,N_3920,N_4608);
nor U7193 (N_7193,N_1995,N_4060);
nor U7194 (N_7194,N_2834,N_2918);
and U7195 (N_7195,N_2275,N_2707);
nor U7196 (N_7196,N_828,N_1386);
and U7197 (N_7197,N_4381,N_763);
and U7198 (N_7198,N_1705,N_4457);
nand U7199 (N_7199,N_769,N_2049);
nand U7200 (N_7200,N_3697,N_557);
nor U7201 (N_7201,N_4968,N_3798);
or U7202 (N_7202,N_4590,N_94);
xor U7203 (N_7203,N_806,N_4615);
or U7204 (N_7204,N_3633,N_1421);
nor U7205 (N_7205,N_4738,N_2415);
nor U7206 (N_7206,N_1495,N_4672);
nor U7207 (N_7207,N_2397,N_319);
nor U7208 (N_7208,N_3410,N_980);
xor U7209 (N_7209,N_3099,N_742);
nand U7210 (N_7210,N_4866,N_3680);
nand U7211 (N_7211,N_3169,N_1589);
nand U7212 (N_7212,N_4359,N_4870);
and U7213 (N_7213,N_1965,N_1259);
or U7214 (N_7214,N_3415,N_3388);
and U7215 (N_7215,N_4912,N_160);
xor U7216 (N_7216,N_1053,N_1484);
nand U7217 (N_7217,N_4874,N_4238);
xnor U7218 (N_7218,N_3958,N_4411);
nor U7219 (N_7219,N_2674,N_454);
nand U7220 (N_7220,N_51,N_1397);
nor U7221 (N_7221,N_4108,N_1477);
nor U7222 (N_7222,N_2951,N_4888);
and U7223 (N_7223,N_726,N_3332);
nor U7224 (N_7224,N_4087,N_3376);
xnor U7225 (N_7225,N_886,N_3702);
nor U7226 (N_7226,N_1913,N_4221);
and U7227 (N_7227,N_1437,N_3349);
nor U7228 (N_7228,N_56,N_4142);
and U7229 (N_7229,N_2724,N_556);
nand U7230 (N_7230,N_579,N_4640);
nor U7231 (N_7231,N_37,N_2247);
or U7232 (N_7232,N_1943,N_1345);
nor U7233 (N_7233,N_4270,N_2833);
and U7234 (N_7234,N_671,N_1856);
nand U7235 (N_7235,N_1285,N_2800);
and U7236 (N_7236,N_538,N_204);
nand U7237 (N_7237,N_719,N_3667);
nand U7238 (N_7238,N_4654,N_4650);
or U7239 (N_7239,N_3816,N_3089);
nand U7240 (N_7240,N_3775,N_4158);
or U7241 (N_7241,N_1646,N_393);
nor U7242 (N_7242,N_870,N_2314);
xnor U7243 (N_7243,N_3269,N_2215);
and U7244 (N_7244,N_2744,N_4530);
or U7245 (N_7245,N_737,N_3467);
nand U7246 (N_7246,N_3144,N_1068);
nor U7247 (N_7247,N_1647,N_2941);
nor U7248 (N_7248,N_1697,N_1352);
nand U7249 (N_7249,N_771,N_2339);
nor U7250 (N_7250,N_1318,N_4663);
and U7251 (N_7251,N_4699,N_323);
nor U7252 (N_7252,N_3289,N_3243);
and U7253 (N_7253,N_3368,N_749);
nor U7254 (N_7254,N_3744,N_1491);
and U7255 (N_7255,N_2965,N_1487);
or U7256 (N_7256,N_1091,N_1552);
or U7257 (N_7257,N_115,N_2552);
nor U7258 (N_7258,N_4042,N_4678);
nand U7259 (N_7259,N_1666,N_2000);
or U7260 (N_7260,N_794,N_2409);
and U7261 (N_7261,N_1358,N_1018);
or U7262 (N_7262,N_4186,N_3758);
nand U7263 (N_7263,N_3679,N_2190);
nor U7264 (N_7264,N_3591,N_3020);
or U7265 (N_7265,N_4085,N_2836);
nand U7266 (N_7266,N_952,N_2026);
or U7267 (N_7267,N_1455,N_1849);
and U7268 (N_7268,N_3184,N_1709);
nor U7269 (N_7269,N_4852,N_283);
and U7270 (N_7270,N_359,N_540);
or U7271 (N_7271,N_4404,N_4124);
nand U7272 (N_7272,N_3218,N_241);
nor U7273 (N_7273,N_4952,N_3050);
and U7274 (N_7274,N_2125,N_3834);
nor U7275 (N_7275,N_1140,N_1785);
or U7276 (N_7276,N_4355,N_4160);
nand U7277 (N_7277,N_2336,N_4675);
or U7278 (N_7278,N_2930,N_3852);
xor U7279 (N_7279,N_1945,N_228);
and U7280 (N_7280,N_4893,N_1257);
and U7281 (N_7281,N_632,N_2582);
or U7282 (N_7282,N_3228,N_2166);
or U7283 (N_7283,N_1862,N_1339);
nor U7284 (N_7284,N_764,N_1786);
or U7285 (N_7285,N_2818,N_3936);
nor U7286 (N_7286,N_4024,N_2361);
or U7287 (N_7287,N_1005,N_207);
nor U7288 (N_7288,N_4014,N_4342);
and U7289 (N_7289,N_3577,N_803);
nand U7290 (N_7290,N_832,N_1255);
xnor U7291 (N_7291,N_773,N_364);
and U7292 (N_7292,N_2854,N_4205);
nor U7293 (N_7293,N_247,N_296);
or U7294 (N_7294,N_1245,N_2939);
nor U7295 (N_7295,N_2855,N_1554);
xor U7296 (N_7296,N_2117,N_2053);
nor U7297 (N_7297,N_2232,N_3335);
nand U7298 (N_7298,N_4524,N_2165);
nand U7299 (N_7299,N_2943,N_4519);
nor U7300 (N_7300,N_2364,N_1126);
and U7301 (N_7301,N_14,N_303);
nand U7302 (N_7302,N_3870,N_1950);
and U7303 (N_7303,N_473,N_4198);
nor U7304 (N_7304,N_2100,N_904);
nor U7305 (N_7305,N_567,N_2341);
nand U7306 (N_7306,N_4027,N_1789);
or U7307 (N_7307,N_335,N_537);
and U7308 (N_7308,N_4016,N_4376);
nor U7309 (N_7309,N_1711,N_3164);
nor U7310 (N_7310,N_3418,N_3899);
or U7311 (N_7311,N_1745,N_2219);
or U7312 (N_7312,N_4370,N_1531);
nor U7313 (N_7313,N_3277,N_978);
or U7314 (N_7314,N_922,N_4341);
or U7315 (N_7315,N_3161,N_1480);
and U7316 (N_7316,N_4855,N_2821);
and U7317 (N_7317,N_2128,N_2997);
and U7318 (N_7318,N_3344,N_3659);
nand U7319 (N_7319,N_4037,N_4915);
and U7320 (N_7320,N_4161,N_2523);
nor U7321 (N_7321,N_3544,N_753);
nand U7322 (N_7322,N_3727,N_3175);
nand U7323 (N_7323,N_3093,N_4094);
nand U7324 (N_7324,N_3561,N_1728);
and U7325 (N_7325,N_1313,N_907);
and U7326 (N_7326,N_2849,N_1886);
nand U7327 (N_7327,N_2014,N_3641);
and U7328 (N_7328,N_4495,N_4176);
nor U7329 (N_7329,N_161,N_2040);
nor U7330 (N_7330,N_3139,N_4490);
or U7331 (N_7331,N_3264,N_31);
or U7332 (N_7332,N_4985,N_4787);
or U7333 (N_7333,N_4537,N_1982);
nor U7334 (N_7334,N_2203,N_2059);
or U7335 (N_7335,N_780,N_4148);
or U7336 (N_7336,N_1373,N_2787);
and U7337 (N_7337,N_676,N_4943);
and U7338 (N_7338,N_1065,N_1879);
nand U7339 (N_7339,N_72,N_4234);
nor U7340 (N_7340,N_2371,N_4029);
and U7341 (N_7341,N_4144,N_129);
nand U7342 (N_7342,N_2844,N_1360);
and U7343 (N_7343,N_4182,N_3525);
and U7344 (N_7344,N_2163,N_916);
nand U7345 (N_7345,N_2533,N_1097);
nor U7346 (N_7346,N_1103,N_4664);
or U7347 (N_7347,N_1212,N_1302);
or U7348 (N_7348,N_954,N_3110);
and U7349 (N_7349,N_1704,N_4507);
nor U7350 (N_7350,N_3165,N_1861);
or U7351 (N_7351,N_1729,N_1630);
nand U7352 (N_7352,N_367,N_4034);
and U7353 (N_7353,N_4652,N_288);
nand U7354 (N_7354,N_2024,N_3031);
nand U7355 (N_7355,N_2105,N_1297);
or U7356 (N_7356,N_1925,N_844);
or U7357 (N_7357,N_1832,N_1516);
and U7358 (N_7358,N_733,N_4132);
nor U7359 (N_7359,N_124,N_1047);
and U7360 (N_7360,N_1702,N_1139);
or U7361 (N_7361,N_3849,N_1356);
and U7362 (N_7362,N_2234,N_459);
nor U7363 (N_7363,N_4543,N_2673);
and U7364 (N_7364,N_4584,N_3125);
nor U7365 (N_7365,N_4707,N_3075);
and U7366 (N_7366,N_2435,N_945);
and U7367 (N_7367,N_252,N_461);
and U7368 (N_7368,N_409,N_3356);
or U7369 (N_7369,N_895,N_164);
nand U7370 (N_7370,N_1871,N_154);
nand U7371 (N_7371,N_4445,N_1215);
xnor U7372 (N_7372,N_551,N_3632);
xor U7373 (N_7373,N_4451,N_2598);
nand U7374 (N_7374,N_4973,N_4898);
and U7375 (N_7375,N_3287,N_4741);
nand U7376 (N_7376,N_3965,N_3925);
or U7377 (N_7377,N_3159,N_2359);
and U7378 (N_7378,N_1765,N_3724);
or U7379 (N_7379,N_3730,N_2474);
nand U7380 (N_7380,N_3345,N_1133);
nand U7381 (N_7381,N_4159,N_1118);
nand U7382 (N_7382,N_2388,N_2346);
nor U7383 (N_7383,N_4488,N_2428);
or U7384 (N_7384,N_3723,N_1217);
or U7385 (N_7385,N_503,N_3451);
nor U7386 (N_7386,N_3832,N_492);
or U7387 (N_7387,N_4064,N_3737);
nand U7388 (N_7388,N_479,N_2315);
or U7389 (N_7389,N_552,N_4596);
nor U7390 (N_7390,N_2602,N_4638);
or U7391 (N_7391,N_2562,N_2286);
or U7392 (N_7392,N_2207,N_3585);
and U7393 (N_7393,N_1262,N_1159);
nand U7394 (N_7394,N_3394,N_2649);
nor U7395 (N_7395,N_2846,N_300);
or U7396 (N_7396,N_2058,N_2778);
nand U7397 (N_7397,N_3146,N_1287);
nor U7398 (N_7398,N_3663,N_4131);
or U7399 (N_7399,N_4271,N_1609);
or U7400 (N_7400,N_3948,N_2699);
and U7401 (N_7401,N_240,N_3768);
and U7402 (N_7402,N_4860,N_2715);
nor U7403 (N_7403,N_1034,N_4748);
nand U7404 (N_7404,N_275,N_4440);
nand U7405 (N_7405,N_1450,N_873);
nand U7406 (N_7406,N_3156,N_2714);
nor U7407 (N_7407,N_871,N_1806);
or U7408 (N_7408,N_1163,N_4847);
and U7409 (N_7409,N_912,N_4162);
nand U7410 (N_7410,N_3323,N_2365);
nor U7411 (N_7411,N_4569,N_915);
or U7412 (N_7412,N_3406,N_746);
nor U7413 (N_7413,N_320,N_258);
nor U7414 (N_7414,N_471,N_4432);
nand U7415 (N_7415,N_2508,N_3533);
nand U7416 (N_7416,N_826,N_4666);
or U7417 (N_7417,N_2676,N_2466);
and U7418 (N_7418,N_4323,N_3917);
nand U7419 (N_7419,N_1117,N_1639);
or U7420 (N_7420,N_1236,N_3761);
nor U7421 (N_7421,N_3505,N_951);
nand U7422 (N_7422,N_574,N_1817);
nor U7423 (N_7423,N_19,N_3359);
or U7424 (N_7424,N_939,N_2280);
nor U7425 (N_7425,N_2345,N_4068);
nor U7426 (N_7426,N_482,N_1724);
or U7427 (N_7427,N_2020,N_4425);
nand U7428 (N_7428,N_878,N_2503);
nand U7429 (N_7429,N_4835,N_2608);
nor U7430 (N_7430,N_508,N_908);
or U7431 (N_7431,N_836,N_516);
nand U7432 (N_7432,N_2655,N_1961);
nand U7433 (N_7433,N_4282,N_1622);
nand U7434 (N_7434,N_3754,N_1379);
and U7435 (N_7435,N_2801,N_1213);
nor U7436 (N_7436,N_4928,N_1923);
and U7437 (N_7437,N_1539,N_4045);
nand U7438 (N_7438,N_377,N_1976);
and U7439 (N_7439,N_465,N_4770);
nand U7440 (N_7440,N_4617,N_2319);
nor U7441 (N_7441,N_3614,N_3124);
or U7442 (N_7442,N_3241,N_3888);
or U7443 (N_7443,N_4054,N_4152);
nor U7444 (N_7444,N_157,N_3199);
or U7445 (N_7445,N_2367,N_3460);
nand U7446 (N_7446,N_3532,N_2871);
nand U7447 (N_7447,N_2145,N_134);
or U7448 (N_7448,N_4642,N_285);
and U7449 (N_7449,N_1014,N_1141);
nand U7450 (N_7450,N_3786,N_1860);
and U7451 (N_7451,N_722,N_944);
nand U7452 (N_7452,N_1457,N_2267);
nor U7453 (N_7453,N_1346,N_2759);
and U7454 (N_7454,N_387,N_4390);
nand U7455 (N_7455,N_1282,N_3593);
and U7456 (N_7456,N_4802,N_2906);
nor U7457 (N_7457,N_4725,N_4294);
nand U7458 (N_7458,N_3275,N_4477);
and U7459 (N_7459,N_2107,N_1340);
and U7460 (N_7460,N_4798,N_326);
xnor U7461 (N_7461,N_1900,N_765);
nand U7462 (N_7462,N_3201,N_3664);
and U7463 (N_7463,N_1544,N_1310);
and U7464 (N_7464,N_947,N_2061);
or U7465 (N_7465,N_1952,N_3290);
or U7466 (N_7466,N_4043,N_4992);
nor U7467 (N_7467,N_3527,N_221);
nor U7468 (N_7468,N_4603,N_682);
nor U7469 (N_7469,N_4735,N_3657);
nand U7470 (N_7470,N_3498,N_1957);
nor U7471 (N_7471,N_788,N_1361);
nor U7472 (N_7472,N_525,N_1222);
nand U7473 (N_7473,N_1369,N_962);
nand U7474 (N_7474,N_1229,N_2957);
nor U7475 (N_7475,N_4456,N_4708);
nand U7476 (N_7476,N_2880,N_257);
nor U7477 (N_7477,N_4380,N_527);
nand U7478 (N_7478,N_1573,N_4807);
or U7479 (N_7479,N_2877,N_4481);
and U7480 (N_7480,N_46,N_3854);
nor U7481 (N_7481,N_3137,N_2223);
nor U7482 (N_7482,N_4307,N_462);
nor U7483 (N_7483,N_1787,N_4677);
nor U7484 (N_7484,N_3249,N_418);
nor U7485 (N_7485,N_1364,N_1156);
nor U7486 (N_7486,N_2726,N_515);
and U7487 (N_7487,N_2915,N_1407);
nand U7488 (N_7488,N_3865,N_1253);
and U7489 (N_7489,N_896,N_4716);
nand U7490 (N_7490,N_3810,N_179);
xnor U7491 (N_7491,N_4989,N_3280);
nor U7492 (N_7492,N_2381,N_2565);
and U7493 (N_7493,N_2144,N_2929);
nand U7494 (N_7494,N_504,N_4479);
nand U7495 (N_7495,N_256,N_3407);
nand U7496 (N_7496,N_627,N_3643);
nand U7497 (N_7497,N_3321,N_356);
nand U7498 (N_7498,N_3735,N_692);
nand U7499 (N_7499,N_3192,N_3961);
nor U7500 (N_7500,N_3636,N_563);
nand U7501 (N_7501,N_355,N_2300);
nand U7502 (N_7502,N_3361,N_2443);
nand U7503 (N_7503,N_3781,N_4149);
nand U7504 (N_7504,N_2107,N_348);
and U7505 (N_7505,N_488,N_1312);
nor U7506 (N_7506,N_1209,N_1381);
and U7507 (N_7507,N_295,N_4418);
and U7508 (N_7508,N_2475,N_2359);
and U7509 (N_7509,N_2884,N_1839);
and U7510 (N_7510,N_4959,N_4670);
nand U7511 (N_7511,N_4301,N_1935);
nor U7512 (N_7512,N_2731,N_2448);
nor U7513 (N_7513,N_964,N_211);
and U7514 (N_7514,N_2424,N_1521);
nor U7515 (N_7515,N_2411,N_3928);
nor U7516 (N_7516,N_4360,N_3575);
and U7517 (N_7517,N_713,N_2900);
nand U7518 (N_7518,N_4323,N_1800);
nand U7519 (N_7519,N_3081,N_1626);
nand U7520 (N_7520,N_1141,N_1526);
nor U7521 (N_7521,N_4307,N_451);
xor U7522 (N_7522,N_3616,N_4409);
nand U7523 (N_7523,N_189,N_1675);
or U7524 (N_7524,N_3323,N_3934);
nor U7525 (N_7525,N_4371,N_1909);
nor U7526 (N_7526,N_2100,N_4001);
nor U7527 (N_7527,N_114,N_3078);
and U7528 (N_7528,N_941,N_3658);
or U7529 (N_7529,N_4407,N_789);
nand U7530 (N_7530,N_4347,N_3061);
or U7531 (N_7531,N_1220,N_2758);
or U7532 (N_7532,N_1472,N_373);
nand U7533 (N_7533,N_4433,N_915);
nand U7534 (N_7534,N_1865,N_993);
nor U7535 (N_7535,N_2165,N_2601);
or U7536 (N_7536,N_3233,N_2014);
or U7537 (N_7537,N_4507,N_1777);
nor U7538 (N_7538,N_1389,N_1992);
nand U7539 (N_7539,N_4756,N_1083);
nor U7540 (N_7540,N_4616,N_499);
and U7541 (N_7541,N_1792,N_730);
nand U7542 (N_7542,N_4259,N_2000);
or U7543 (N_7543,N_4100,N_79);
nand U7544 (N_7544,N_4124,N_4758);
nand U7545 (N_7545,N_1433,N_3752);
nor U7546 (N_7546,N_3408,N_2804);
or U7547 (N_7547,N_1650,N_292);
and U7548 (N_7548,N_4958,N_2439);
nand U7549 (N_7549,N_3475,N_1415);
or U7550 (N_7550,N_1591,N_1055);
nor U7551 (N_7551,N_490,N_1926);
and U7552 (N_7552,N_1706,N_4530);
or U7553 (N_7553,N_4217,N_4232);
nand U7554 (N_7554,N_386,N_89);
nand U7555 (N_7555,N_1293,N_469);
nand U7556 (N_7556,N_1814,N_3055);
nand U7557 (N_7557,N_4985,N_3499);
or U7558 (N_7558,N_1523,N_882);
and U7559 (N_7559,N_2324,N_3613);
nor U7560 (N_7560,N_4002,N_413);
nand U7561 (N_7561,N_2286,N_3926);
nor U7562 (N_7562,N_2351,N_953);
or U7563 (N_7563,N_3462,N_2372);
or U7564 (N_7564,N_4173,N_2014);
nand U7565 (N_7565,N_3940,N_2528);
nand U7566 (N_7566,N_2729,N_368);
and U7567 (N_7567,N_485,N_3698);
xor U7568 (N_7568,N_3194,N_4987);
nand U7569 (N_7569,N_4039,N_4537);
nand U7570 (N_7570,N_2151,N_1856);
and U7571 (N_7571,N_4137,N_2196);
nor U7572 (N_7572,N_297,N_2547);
and U7573 (N_7573,N_1531,N_4877);
nand U7574 (N_7574,N_4536,N_232);
nor U7575 (N_7575,N_3646,N_2615);
and U7576 (N_7576,N_2895,N_3611);
or U7577 (N_7577,N_2021,N_3865);
or U7578 (N_7578,N_250,N_457);
and U7579 (N_7579,N_1684,N_168);
nand U7580 (N_7580,N_3502,N_1457);
or U7581 (N_7581,N_3067,N_2022);
or U7582 (N_7582,N_293,N_2262);
nand U7583 (N_7583,N_2964,N_2204);
nand U7584 (N_7584,N_3373,N_1952);
or U7585 (N_7585,N_668,N_1281);
nor U7586 (N_7586,N_2799,N_2485);
or U7587 (N_7587,N_99,N_1462);
nor U7588 (N_7588,N_2310,N_3530);
and U7589 (N_7589,N_3455,N_4778);
or U7590 (N_7590,N_1510,N_2574);
and U7591 (N_7591,N_3405,N_1854);
nand U7592 (N_7592,N_2716,N_1906);
nand U7593 (N_7593,N_3767,N_2922);
nand U7594 (N_7594,N_1292,N_2710);
nor U7595 (N_7595,N_2299,N_4446);
or U7596 (N_7596,N_2301,N_4919);
nor U7597 (N_7597,N_2013,N_2984);
xor U7598 (N_7598,N_1382,N_3218);
nor U7599 (N_7599,N_4426,N_1510);
nand U7600 (N_7600,N_4969,N_1067);
or U7601 (N_7601,N_3680,N_487);
nand U7602 (N_7602,N_425,N_1355);
nor U7603 (N_7603,N_0,N_1360);
and U7604 (N_7604,N_4482,N_2366);
nor U7605 (N_7605,N_2547,N_2271);
nor U7606 (N_7606,N_188,N_4985);
and U7607 (N_7607,N_3612,N_4607);
nand U7608 (N_7608,N_1295,N_1054);
nor U7609 (N_7609,N_1930,N_3703);
and U7610 (N_7610,N_2043,N_3800);
xnor U7611 (N_7611,N_646,N_3614);
nand U7612 (N_7612,N_2202,N_3034);
or U7613 (N_7613,N_3297,N_1981);
nand U7614 (N_7614,N_4669,N_2959);
and U7615 (N_7615,N_1324,N_21);
or U7616 (N_7616,N_3842,N_3243);
nand U7617 (N_7617,N_2636,N_1373);
nor U7618 (N_7618,N_3125,N_4492);
or U7619 (N_7619,N_858,N_4771);
and U7620 (N_7620,N_3301,N_712);
xor U7621 (N_7621,N_3392,N_1539);
and U7622 (N_7622,N_849,N_1893);
or U7623 (N_7623,N_369,N_1565);
nand U7624 (N_7624,N_3533,N_4378);
and U7625 (N_7625,N_4397,N_3606);
or U7626 (N_7626,N_2971,N_1661);
and U7627 (N_7627,N_2742,N_1746);
and U7628 (N_7628,N_3474,N_2949);
nor U7629 (N_7629,N_970,N_1692);
and U7630 (N_7630,N_2348,N_2537);
nand U7631 (N_7631,N_241,N_3613);
nand U7632 (N_7632,N_2558,N_1233);
nand U7633 (N_7633,N_4025,N_2346);
nor U7634 (N_7634,N_2746,N_622);
and U7635 (N_7635,N_4994,N_3605);
nand U7636 (N_7636,N_2904,N_839);
and U7637 (N_7637,N_4335,N_2684);
nand U7638 (N_7638,N_4722,N_4930);
and U7639 (N_7639,N_3208,N_2379);
and U7640 (N_7640,N_469,N_4221);
or U7641 (N_7641,N_3329,N_2816);
or U7642 (N_7642,N_2724,N_1670);
or U7643 (N_7643,N_2873,N_1933);
nor U7644 (N_7644,N_4756,N_3658);
nand U7645 (N_7645,N_2275,N_741);
and U7646 (N_7646,N_2137,N_3507);
or U7647 (N_7647,N_1037,N_2240);
nand U7648 (N_7648,N_3575,N_1664);
and U7649 (N_7649,N_58,N_96);
nor U7650 (N_7650,N_4897,N_1203);
nand U7651 (N_7651,N_42,N_2539);
nor U7652 (N_7652,N_1551,N_4405);
or U7653 (N_7653,N_3149,N_2829);
or U7654 (N_7654,N_3630,N_427);
nor U7655 (N_7655,N_3245,N_4514);
or U7656 (N_7656,N_1119,N_691);
nor U7657 (N_7657,N_3225,N_602);
or U7658 (N_7658,N_3026,N_193);
nor U7659 (N_7659,N_3345,N_4727);
nand U7660 (N_7660,N_2575,N_2714);
or U7661 (N_7661,N_2478,N_2679);
nor U7662 (N_7662,N_2972,N_4803);
and U7663 (N_7663,N_2045,N_407);
nand U7664 (N_7664,N_3475,N_3736);
nor U7665 (N_7665,N_3273,N_4189);
nor U7666 (N_7666,N_1166,N_728);
nand U7667 (N_7667,N_97,N_3078);
nor U7668 (N_7668,N_3200,N_722);
or U7669 (N_7669,N_75,N_4312);
or U7670 (N_7670,N_2470,N_74);
and U7671 (N_7671,N_4836,N_2360);
and U7672 (N_7672,N_4372,N_4117);
or U7673 (N_7673,N_3759,N_1690);
or U7674 (N_7674,N_3010,N_2571);
nand U7675 (N_7675,N_623,N_2087);
xnor U7676 (N_7676,N_759,N_266);
and U7677 (N_7677,N_692,N_1759);
nand U7678 (N_7678,N_1859,N_2816);
nand U7679 (N_7679,N_4562,N_1519);
nor U7680 (N_7680,N_4869,N_3994);
and U7681 (N_7681,N_1377,N_2292);
or U7682 (N_7682,N_773,N_580);
nor U7683 (N_7683,N_2190,N_1418);
and U7684 (N_7684,N_2342,N_4446);
nor U7685 (N_7685,N_4741,N_384);
nor U7686 (N_7686,N_1012,N_4889);
and U7687 (N_7687,N_3145,N_592);
or U7688 (N_7688,N_2351,N_3727);
or U7689 (N_7689,N_4992,N_2427);
nand U7690 (N_7690,N_1241,N_3470);
or U7691 (N_7691,N_4267,N_504);
and U7692 (N_7692,N_2434,N_3891);
and U7693 (N_7693,N_3887,N_1036);
nand U7694 (N_7694,N_4848,N_1803);
nor U7695 (N_7695,N_3037,N_2635);
nand U7696 (N_7696,N_2933,N_754);
nand U7697 (N_7697,N_2786,N_3467);
nand U7698 (N_7698,N_1732,N_2767);
or U7699 (N_7699,N_1880,N_3117);
nor U7700 (N_7700,N_3125,N_3584);
and U7701 (N_7701,N_3000,N_4139);
or U7702 (N_7702,N_3774,N_2672);
and U7703 (N_7703,N_2964,N_2776);
xnor U7704 (N_7704,N_4035,N_663);
and U7705 (N_7705,N_2855,N_2408);
nand U7706 (N_7706,N_4588,N_2155);
or U7707 (N_7707,N_3513,N_4774);
nand U7708 (N_7708,N_972,N_1097);
or U7709 (N_7709,N_3959,N_416);
or U7710 (N_7710,N_924,N_3337);
and U7711 (N_7711,N_4361,N_293);
nor U7712 (N_7712,N_2008,N_4596);
and U7713 (N_7713,N_4867,N_1037);
or U7714 (N_7714,N_1095,N_281);
nand U7715 (N_7715,N_3755,N_4029);
nand U7716 (N_7716,N_3552,N_2152);
nand U7717 (N_7717,N_392,N_3352);
or U7718 (N_7718,N_1685,N_1334);
nand U7719 (N_7719,N_3686,N_4598);
and U7720 (N_7720,N_237,N_600);
and U7721 (N_7721,N_3922,N_4947);
nand U7722 (N_7722,N_1101,N_4245);
nand U7723 (N_7723,N_283,N_1907);
nand U7724 (N_7724,N_3318,N_4266);
or U7725 (N_7725,N_5,N_2415);
and U7726 (N_7726,N_4472,N_4649);
nand U7727 (N_7727,N_2744,N_3992);
nor U7728 (N_7728,N_419,N_4410);
nor U7729 (N_7729,N_101,N_3319);
nor U7730 (N_7730,N_4577,N_3824);
or U7731 (N_7731,N_1262,N_4382);
nand U7732 (N_7732,N_4702,N_4611);
nor U7733 (N_7733,N_2787,N_353);
and U7734 (N_7734,N_4059,N_3220);
nand U7735 (N_7735,N_4653,N_963);
xor U7736 (N_7736,N_462,N_2954);
and U7737 (N_7737,N_4873,N_4278);
or U7738 (N_7738,N_722,N_670);
and U7739 (N_7739,N_4287,N_2439);
or U7740 (N_7740,N_3130,N_1225);
nand U7741 (N_7741,N_3003,N_4191);
nand U7742 (N_7742,N_1706,N_4056);
or U7743 (N_7743,N_4669,N_3163);
nand U7744 (N_7744,N_2535,N_515);
nor U7745 (N_7745,N_229,N_590);
and U7746 (N_7746,N_2907,N_2537);
nor U7747 (N_7747,N_3475,N_878);
and U7748 (N_7748,N_2510,N_167);
and U7749 (N_7749,N_1647,N_551);
and U7750 (N_7750,N_1137,N_2222);
nand U7751 (N_7751,N_346,N_1028);
or U7752 (N_7752,N_2925,N_2744);
nor U7753 (N_7753,N_4250,N_4882);
or U7754 (N_7754,N_2836,N_2910);
nand U7755 (N_7755,N_4288,N_3694);
nand U7756 (N_7756,N_581,N_68);
nand U7757 (N_7757,N_2817,N_1966);
nand U7758 (N_7758,N_4798,N_4053);
and U7759 (N_7759,N_2128,N_4639);
nand U7760 (N_7760,N_585,N_998);
or U7761 (N_7761,N_2365,N_1516);
nor U7762 (N_7762,N_4406,N_2480);
or U7763 (N_7763,N_4845,N_663);
xnor U7764 (N_7764,N_2670,N_1989);
or U7765 (N_7765,N_3386,N_4600);
nor U7766 (N_7766,N_2535,N_4039);
or U7767 (N_7767,N_2554,N_2098);
nand U7768 (N_7768,N_1454,N_15);
and U7769 (N_7769,N_3611,N_2222);
or U7770 (N_7770,N_3852,N_1101);
or U7771 (N_7771,N_298,N_1013);
nor U7772 (N_7772,N_4990,N_4869);
nand U7773 (N_7773,N_488,N_1129);
or U7774 (N_7774,N_2892,N_150);
nor U7775 (N_7775,N_4784,N_2623);
nor U7776 (N_7776,N_4168,N_2380);
nand U7777 (N_7777,N_4571,N_60);
nor U7778 (N_7778,N_1704,N_1636);
and U7779 (N_7779,N_4852,N_4630);
nand U7780 (N_7780,N_3822,N_802);
nor U7781 (N_7781,N_4868,N_1841);
nor U7782 (N_7782,N_1040,N_3340);
and U7783 (N_7783,N_2306,N_1656);
nand U7784 (N_7784,N_2545,N_3532);
or U7785 (N_7785,N_2611,N_4714);
nor U7786 (N_7786,N_4227,N_749);
nand U7787 (N_7787,N_3140,N_545);
xnor U7788 (N_7788,N_3396,N_3723);
nor U7789 (N_7789,N_459,N_352);
nand U7790 (N_7790,N_506,N_1447);
nand U7791 (N_7791,N_1055,N_3591);
nand U7792 (N_7792,N_1815,N_718);
or U7793 (N_7793,N_3858,N_160);
and U7794 (N_7794,N_1559,N_4407);
nand U7795 (N_7795,N_2555,N_3978);
nor U7796 (N_7796,N_2215,N_2451);
or U7797 (N_7797,N_4456,N_4315);
and U7798 (N_7798,N_1747,N_2180);
or U7799 (N_7799,N_1264,N_4190);
xnor U7800 (N_7800,N_1882,N_3824);
or U7801 (N_7801,N_4363,N_4101);
and U7802 (N_7802,N_416,N_1128);
nor U7803 (N_7803,N_1633,N_2647);
or U7804 (N_7804,N_1110,N_646);
nand U7805 (N_7805,N_3888,N_3786);
or U7806 (N_7806,N_1273,N_3938);
and U7807 (N_7807,N_980,N_4516);
or U7808 (N_7808,N_3718,N_3939);
and U7809 (N_7809,N_4740,N_2814);
and U7810 (N_7810,N_4222,N_600);
and U7811 (N_7811,N_2706,N_1111);
nand U7812 (N_7812,N_713,N_2682);
or U7813 (N_7813,N_660,N_2048);
nor U7814 (N_7814,N_4215,N_3589);
and U7815 (N_7815,N_4519,N_484);
nor U7816 (N_7816,N_1026,N_2376);
nand U7817 (N_7817,N_4646,N_1832);
or U7818 (N_7818,N_525,N_3866);
nand U7819 (N_7819,N_3400,N_1008);
and U7820 (N_7820,N_4811,N_103);
or U7821 (N_7821,N_4330,N_3072);
nand U7822 (N_7822,N_2296,N_2355);
nor U7823 (N_7823,N_4783,N_4232);
nor U7824 (N_7824,N_4360,N_0);
nor U7825 (N_7825,N_3903,N_2419);
and U7826 (N_7826,N_374,N_4908);
nand U7827 (N_7827,N_2221,N_3165);
nand U7828 (N_7828,N_1684,N_1465);
or U7829 (N_7829,N_4888,N_893);
or U7830 (N_7830,N_4534,N_118);
xnor U7831 (N_7831,N_4148,N_3946);
or U7832 (N_7832,N_1831,N_4782);
and U7833 (N_7833,N_3957,N_4933);
or U7834 (N_7834,N_1969,N_4257);
or U7835 (N_7835,N_2395,N_4634);
and U7836 (N_7836,N_1811,N_4981);
nand U7837 (N_7837,N_734,N_1997);
or U7838 (N_7838,N_1648,N_1735);
nand U7839 (N_7839,N_1984,N_413);
or U7840 (N_7840,N_1086,N_757);
nor U7841 (N_7841,N_3392,N_72);
nor U7842 (N_7842,N_102,N_1767);
nand U7843 (N_7843,N_3297,N_3068);
nand U7844 (N_7844,N_100,N_784);
or U7845 (N_7845,N_4858,N_1434);
or U7846 (N_7846,N_1261,N_4435);
and U7847 (N_7847,N_2180,N_661);
nand U7848 (N_7848,N_297,N_523);
xnor U7849 (N_7849,N_700,N_1557);
nor U7850 (N_7850,N_2354,N_1041);
xor U7851 (N_7851,N_4563,N_310);
xor U7852 (N_7852,N_190,N_2055);
nor U7853 (N_7853,N_2470,N_59);
nand U7854 (N_7854,N_4577,N_53);
and U7855 (N_7855,N_1615,N_748);
nor U7856 (N_7856,N_3514,N_2837);
and U7857 (N_7857,N_1871,N_4696);
nand U7858 (N_7858,N_3892,N_682);
or U7859 (N_7859,N_4204,N_1008);
nand U7860 (N_7860,N_484,N_175);
nor U7861 (N_7861,N_3819,N_2925);
nor U7862 (N_7862,N_4920,N_3482);
nand U7863 (N_7863,N_3903,N_1743);
nand U7864 (N_7864,N_4737,N_2281);
and U7865 (N_7865,N_1082,N_1335);
and U7866 (N_7866,N_4071,N_2754);
nor U7867 (N_7867,N_4770,N_1406);
and U7868 (N_7868,N_4627,N_3258);
nand U7869 (N_7869,N_4884,N_4396);
nor U7870 (N_7870,N_2818,N_3912);
and U7871 (N_7871,N_4381,N_2415);
nand U7872 (N_7872,N_50,N_606);
nand U7873 (N_7873,N_1558,N_2130);
or U7874 (N_7874,N_4675,N_4040);
nand U7875 (N_7875,N_4190,N_2663);
or U7876 (N_7876,N_1362,N_1202);
or U7877 (N_7877,N_4973,N_49);
or U7878 (N_7878,N_155,N_3530);
and U7879 (N_7879,N_1317,N_4190);
and U7880 (N_7880,N_4648,N_277);
or U7881 (N_7881,N_407,N_2870);
or U7882 (N_7882,N_1507,N_348);
nor U7883 (N_7883,N_1381,N_1609);
and U7884 (N_7884,N_1933,N_694);
nor U7885 (N_7885,N_1413,N_2054);
nand U7886 (N_7886,N_1584,N_1054);
and U7887 (N_7887,N_2585,N_1235);
nor U7888 (N_7888,N_1022,N_1401);
or U7889 (N_7889,N_1873,N_1353);
or U7890 (N_7890,N_187,N_3998);
nor U7891 (N_7891,N_663,N_1447);
nand U7892 (N_7892,N_4407,N_2312);
or U7893 (N_7893,N_3635,N_1315);
and U7894 (N_7894,N_4130,N_1592);
nor U7895 (N_7895,N_1277,N_1448);
nand U7896 (N_7896,N_4618,N_749);
or U7897 (N_7897,N_2339,N_4008);
nor U7898 (N_7898,N_4906,N_4962);
xnor U7899 (N_7899,N_598,N_712);
nor U7900 (N_7900,N_3725,N_409);
and U7901 (N_7901,N_4559,N_2764);
or U7902 (N_7902,N_2321,N_3261);
nand U7903 (N_7903,N_1415,N_1518);
nand U7904 (N_7904,N_3908,N_1739);
nor U7905 (N_7905,N_4903,N_1721);
or U7906 (N_7906,N_642,N_734);
or U7907 (N_7907,N_1118,N_3185);
or U7908 (N_7908,N_4287,N_4657);
or U7909 (N_7909,N_2254,N_4091);
and U7910 (N_7910,N_1713,N_3013);
nand U7911 (N_7911,N_4237,N_1116);
nand U7912 (N_7912,N_1220,N_2848);
nand U7913 (N_7913,N_2060,N_1722);
xnor U7914 (N_7914,N_1708,N_489);
nor U7915 (N_7915,N_4974,N_2197);
and U7916 (N_7916,N_4700,N_2796);
or U7917 (N_7917,N_4720,N_2616);
and U7918 (N_7918,N_132,N_2672);
nand U7919 (N_7919,N_4050,N_3341);
nor U7920 (N_7920,N_76,N_2512);
or U7921 (N_7921,N_4463,N_436);
nor U7922 (N_7922,N_4288,N_312);
nand U7923 (N_7923,N_822,N_2056);
nand U7924 (N_7924,N_585,N_4226);
and U7925 (N_7925,N_299,N_1443);
nor U7926 (N_7926,N_1434,N_3933);
and U7927 (N_7927,N_2513,N_405);
nand U7928 (N_7928,N_1076,N_4232);
nand U7929 (N_7929,N_22,N_1586);
nor U7930 (N_7930,N_374,N_2745);
and U7931 (N_7931,N_3328,N_3448);
or U7932 (N_7932,N_3920,N_4587);
nor U7933 (N_7933,N_844,N_364);
or U7934 (N_7934,N_4565,N_4960);
or U7935 (N_7935,N_370,N_2476);
nand U7936 (N_7936,N_4368,N_1536);
nor U7937 (N_7937,N_3146,N_4535);
nor U7938 (N_7938,N_3087,N_781);
and U7939 (N_7939,N_1915,N_4459);
or U7940 (N_7940,N_4331,N_1307);
xor U7941 (N_7941,N_4660,N_208);
nand U7942 (N_7942,N_4863,N_964);
and U7943 (N_7943,N_125,N_3462);
and U7944 (N_7944,N_713,N_4172);
nor U7945 (N_7945,N_513,N_3903);
nand U7946 (N_7946,N_1423,N_3581);
or U7947 (N_7947,N_2231,N_1058);
nor U7948 (N_7948,N_2599,N_1458);
and U7949 (N_7949,N_4844,N_950);
or U7950 (N_7950,N_1606,N_4371);
or U7951 (N_7951,N_2451,N_4402);
and U7952 (N_7952,N_4827,N_1714);
nand U7953 (N_7953,N_4062,N_1355);
or U7954 (N_7954,N_2675,N_93);
or U7955 (N_7955,N_507,N_6);
nor U7956 (N_7956,N_3953,N_2379);
nand U7957 (N_7957,N_3379,N_4006);
nand U7958 (N_7958,N_1657,N_4802);
or U7959 (N_7959,N_4300,N_667);
and U7960 (N_7960,N_3997,N_1952);
nand U7961 (N_7961,N_338,N_2705);
nand U7962 (N_7962,N_1980,N_3328);
nand U7963 (N_7963,N_3288,N_2025);
or U7964 (N_7964,N_2824,N_255);
and U7965 (N_7965,N_3713,N_2785);
nor U7966 (N_7966,N_4097,N_1426);
and U7967 (N_7967,N_1622,N_3704);
nor U7968 (N_7968,N_4579,N_4884);
and U7969 (N_7969,N_1356,N_4652);
or U7970 (N_7970,N_4402,N_291);
nor U7971 (N_7971,N_4257,N_1474);
nand U7972 (N_7972,N_1639,N_4924);
nor U7973 (N_7973,N_4832,N_4346);
nor U7974 (N_7974,N_4777,N_2005);
and U7975 (N_7975,N_3014,N_2873);
nand U7976 (N_7976,N_2905,N_95);
and U7977 (N_7977,N_3088,N_4763);
nand U7978 (N_7978,N_4251,N_3269);
nor U7979 (N_7979,N_2947,N_3312);
or U7980 (N_7980,N_3103,N_3164);
xor U7981 (N_7981,N_1467,N_3077);
and U7982 (N_7982,N_1663,N_3449);
or U7983 (N_7983,N_2508,N_630);
and U7984 (N_7984,N_1543,N_3396);
and U7985 (N_7985,N_3175,N_3921);
nand U7986 (N_7986,N_3319,N_1870);
nor U7987 (N_7987,N_3681,N_2084);
and U7988 (N_7988,N_3504,N_4426);
and U7989 (N_7989,N_4360,N_952);
nor U7990 (N_7990,N_417,N_201);
or U7991 (N_7991,N_4143,N_2024);
or U7992 (N_7992,N_3325,N_3328);
nand U7993 (N_7993,N_4037,N_4317);
nand U7994 (N_7994,N_3204,N_720);
nand U7995 (N_7995,N_967,N_1244);
nor U7996 (N_7996,N_350,N_78);
nand U7997 (N_7997,N_4338,N_4459);
nand U7998 (N_7998,N_354,N_1431);
nor U7999 (N_7999,N_4362,N_2117);
nand U8000 (N_8000,N_2825,N_4933);
nand U8001 (N_8001,N_4101,N_2282);
nand U8002 (N_8002,N_3772,N_2824);
nor U8003 (N_8003,N_2243,N_3635);
nor U8004 (N_8004,N_2959,N_409);
nor U8005 (N_8005,N_351,N_4110);
nand U8006 (N_8006,N_4781,N_3943);
nor U8007 (N_8007,N_4338,N_1662);
nor U8008 (N_8008,N_2325,N_1287);
nand U8009 (N_8009,N_2409,N_4671);
and U8010 (N_8010,N_2976,N_3677);
nand U8011 (N_8011,N_966,N_1201);
nor U8012 (N_8012,N_2225,N_167);
nor U8013 (N_8013,N_1947,N_3555);
and U8014 (N_8014,N_4171,N_1462);
nand U8015 (N_8015,N_812,N_1670);
nand U8016 (N_8016,N_3672,N_2975);
nand U8017 (N_8017,N_3713,N_2146);
or U8018 (N_8018,N_3396,N_3643);
nor U8019 (N_8019,N_3884,N_360);
nand U8020 (N_8020,N_2597,N_4731);
or U8021 (N_8021,N_4737,N_4692);
nor U8022 (N_8022,N_4825,N_3402);
or U8023 (N_8023,N_740,N_3091);
nor U8024 (N_8024,N_2364,N_133);
nor U8025 (N_8025,N_1269,N_402);
nand U8026 (N_8026,N_1058,N_2370);
and U8027 (N_8027,N_2563,N_925);
xnor U8028 (N_8028,N_2587,N_2127);
nor U8029 (N_8029,N_169,N_443);
and U8030 (N_8030,N_1052,N_4369);
nor U8031 (N_8031,N_2336,N_1701);
nor U8032 (N_8032,N_1906,N_4636);
nor U8033 (N_8033,N_4488,N_3901);
or U8034 (N_8034,N_2475,N_4382);
nor U8035 (N_8035,N_4105,N_4354);
nor U8036 (N_8036,N_2944,N_2956);
and U8037 (N_8037,N_12,N_51);
nor U8038 (N_8038,N_3751,N_1988);
nand U8039 (N_8039,N_4911,N_712);
nor U8040 (N_8040,N_4345,N_4107);
or U8041 (N_8041,N_1779,N_2583);
nor U8042 (N_8042,N_810,N_727);
nor U8043 (N_8043,N_983,N_3724);
nand U8044 (N_8044,N_3705,N_2691);
nor U8045 (N_8045,N_3591,N_4290);
and U8046 (N_8046,N_2715,N_4285);
nand U8047 (N_8047,N_2322,N_4999);
or U8048 (N_8048,N_689,N_1532);
xnor U8049 (N_8049,N_5,N_876);
and U8050 (N_8050,N_1395,N_4009);
nand U8051 (N_8051,N_1242,N_3530);
or U8052 (N_8052,N_465,N_833);
and U8053 (N_8053,N_2758,N_394);
nor U8054 (N_8054,N_1665,N_4367);
and U8055 (N_8055,N_164,N_1112);
nand U8056 (N_8056,N_2174,N_268);
and U8057 (N_8057,N_4419,N_2711);
or U8058 (N_8058,N_206,N_300);
and U8059 (N_8059,N_3314,N_2567);
nand U8060 (N_8060,N_3204,N_1011);
nor U8061 (N_8061,N_4296,N_2319);
nor U8062 (N_8062,N_4668,N_4431);
nand U8063 (N_8063,N_694,N_1823);
nand U8064 (N_8064,N_1362,N_1663);
and U8065 (N_8065,N_3460,N_1745);
and U8066 (N_8066,N_978,N_3676);
nand U8067 (N_8067,N_607,N_154);
or U8068 (N_8068,N_1418,N_1891);
nor U8069 (N_8069,N_3543,N_2072);
nand U8070 (N_8070,N_1919,N_2585);
nor U8071 (N_8071,N_562,N_543);
or U8072 (N_8072,N_3850,N_4151);
nor U8073 (N_8073,N_831,N_4272);
nand U8074 (N_8074,N_327,N_3695);
and U8075 (N_8075,N_3332,N_4609);
and U8076 (N_8076,N_212,N_4442);
nand U8077 (N_8077,N_1906,N_4682);
or U8078 (N_8078,N_2608,N_2827);
nor U8079 (N_8079,N_3281,N_1919);
nor U8080 (N_8080,N_465,N_514);
nand U8081 (N_8081,N_3032,N_4245);
nor U8082 (N_8082,N_3764,N_4799);
or U8083 (N_8083,N_4479,N_1589);
nor U8084 (N_8084,N_4804,N_143);
nand U8085 (N_8085,N_4520,N_3928);
or U8086 (N_8086,N_2112,N_3647);
nand U8087 (N_8087,N_3019,N_3537);
nor U8088 (N_8088,N_3577,N_826);
nand U8089 (N_8089,N_4899,N_1778);
nor U8090 (N_8090,N_3706,N_1422);
nor U8091 (N_8091,N_1457,N_542);
or U8092 (N_8092,N_2651,N_1674);
and U8093 (N_8093,N_1733,N_51);
and U8094 (N_8094,N_4446,N_2189);
or U8095 (N_8095,N_1730,N_14);
nand U8096 (N_8096,N_3026,N_707);
or U8097 (N_8097,N_502,N_1156);
or U8098 (N_8098,N_1224,N_3605);
and U8099 (N_8099,N_137,N_1244);
nor U8100 (N_8100,N_4588,N_2553);
and U8101 (N_8101,N_3333,N_1226);
or U8102 (N_8102,N_1654,N_4593);
nor U8103 (N_8103,N_3298,N_2401);
and U8104 (N_8104,N_2901,N_2870);
or U8105 (N_8105,N_995,N_4331);
and U8106 (N_8106,N_4732,N_4750);
and U8107 (N_8107,N_2284,N_3811);
or U8108 (N_8108,N_3311,N_528);
nor U8109 (N_8109,N_1199,N_3984);
nand U8110 (N_8110,N_4197,N_370);
or U8111 (N_8111,N_2203,N_3562);
and U8112 (N_8112,N_4384,N_3289);
nor U8113 (N_8113,N_708,N_142);
nor U8114 (N_8114,N_4786,N_986);
or U8115 (N_8115,N_3518,N_3873);
and U8116 (N_8116,N_4213,N_4785);
nand U8117 (N_8117,N_3226,N_4513);
and U8118 (N_8118,N_96,N_4142);
nand U8119 (N_8119,N_3113,N_1498);
xnor U8120 (N_8120,N_3592,N_334);
and U8121 (N_8121,N_4533,N_3448);
nor U8122 (N_8122,N_3638,N_4403);
nor U8123 (N_8123,N_4573,N_934);
and U8124 (N_8124,N_3454,N_2918);
and U8125 (N_8125,N_4468,N_3022);
nand U8126 (N_8126,N_4902,N_312);
and U8127 (N_8127,N_4307,N_4288);
and U8128 (N_8128,N_1600,N_2320);
nor U8129 (N_8129,N_1075,N_2081);
nor U8130 (N_8130,N_1870,N_4274);
nand U8131 (N_8131,N_4331,N_4971);
nor U8132 (N_8132,N_3343,N_3270);
nand U8133 (N_8133,N_3339,N_2925);
or U8134 (N_8134,N_594,N_4023);
nand U8135 (N_8135,N_3465,N_2567);
nor U8136 (N_8136,N_1213,N_3755);
nor U8137 (N_8137,N_3128,N_1753);
and U8138 (N_8138,N_3944,N_156);
nor U8139 (N_8139,N_539,N_2906);
nor U8140 (N_8140,N_2834,N_4290);
or U8141 (N_8141,N_637,N_3541);
or U8142 (N_8142,N_863,N_3992);
nor U8143 (N_8143,N_1189,N_406);
nand U8144 (N_8144,N_4680,N_1248);
and U8145 (N_8145,N_4691,N_3966);
or U8146 (N_8146,N_3169,N_1767);
and U8147 (N_8147,N_841,N_2943);
nor U8148 (N_8148,N_1668,N_822);
or U8149 (N_8149,N_3957,N_3254);
nand U8150 (N_8150,N_1516,N_2049);
or U8151 (N_8151,N_1877,N_44);
or U8152 (N_8152,N_4734,N_2408);
or U8153 (N_8153,N_1395,N_96);
and U8154 (N_8154,N_2813,N_2962);
or U8155 (N_8155,N_1197,N_4258);
and U8156 (N_8156,N_367,N_2071);
nor U8157 (N_8157,N_2637,N_4961);
or U8158 (N_8158,N_2119,N_1117);
nand U8159 (N_8159,N_4942,N_2016);
nor U8160 (N_8160,N_2580,N_2016);
nand U8161 (N_8161,N_760,N_1321);
and U8162 (N_8162,N_583,N_4779);
nor U8163 (N_8163,N_95,N_107);
nor U8164 (N_8164,N_1185,N_4926);
or U8165 (N_8165,N_1505,N_3895);
or U8166 (N_8166,N_1348,N_2628);
and U8167 (N_8167,N_4069,N_827);
xnor U8168 (N_8168,N_2131,N_4420);
or U8169 (N_8169,N_2139,N_861);
or U8170 (N_8170,N_1780,N_3019);
nand U8171 (N_8171,N_785,N_1318);
nand U8172 (N_8172,N_2345,N_2840);
nand U8173 (N_8173,N_3612,N_4818);
or U8174 (N_8174,N_4417,N_1337);
nor U8175 (N_8175,N_2640,N_4508);
nand U8176 (N_8176,N_2918,N_3332);
nor U8177 (N_8177,N_2638,N_120);
nor U8178 (N_8178,N_4746,N_2264);
nor U8179 (N_8179,N_620,N_2551);
or U8180 (N_8180,N_412,N_1461);
xor U8181 (N_8181,N_2646,N_1742);
nand U8182 (N_8182,N_2585,N_3350);
xnor U8183 (N_8183,N_605,N_3408);
nand U8184 (N_8184,N_3853,N_4582);
nor U8185 (N_8185,N_531,N_1115);
nor U8186 (N_8186,N_4234,N_2916);
or U8187 (N_8187,N_2698,N_1701);
or U8188 (N_8188,N_3957,N_2574);
nand U8189 (N_8189,N_576,N_3331);
or U8190 (N_8190,N_3398,N_3578);
and U8191 (N_8191,N_3239,N_1799);
nand U8192 (N_8192,N_4444,N_3465);
and U8193 (N_8193,N_1866,N_4309);
nand U8194 (N_8194,N_4426,N_4148);
and U8195 (N_8195,N_3892,N_4747);
and U8196 (N_8196,N_2866,N_3952);
and U8197 (N_8197,N_84,N_2449);
nand U8198 (N_8198,N_4596,N_4726);
nand U8199 (N_8199,N_407,N_148);
xnor U8200 (N_8200,N_2216,N_1864);
or U8201 (N_8201,N_3074,N_1199);
and U8202 (N_8202,N_214,N_3348);
or U8203 (N_8203,N_1382,N_580);
nor U8204 (N_8204,N_1866,N_515);
or U8205 (N_8205,N_87,N_4999);
nor U8206 (N_8206,N_3560,N_3973);
nand U8207 (N_8207,N_3689,N_3901);
or U8208 (N_8208,N_3113,N_4811);
xnor U8209 (N_8209,N_162,N_724);
nor U8210 (N_8210,N_1028,N_3463);
nor U8211 (N_8211,N_357,N_4596);
or U8212 (N_8212,N_3598,N_770);
nor U8213 (N_8213,N_860,N_2573);
nor U8214 (N_8214,N_1106,N_1838);
or U8215 (N_8215,N_2101,N_1493);
and U8216 (N_8216,N_1220,N_2770);
nor U8217 (N_8217,N_862,N_2749);
nor U8218 (N_8218,N_4797,N_200);
nand U8219 (N_8219,N_1417,N_2494);
nand U8220 (N_8220,N_4411,N_3337);
nand U8221 (N_8221,N_3956,N_3138);
or U8222 (N_8222,N_2805,N_2215);
nor U8223 (N_8223,N_2518,N_2330);
and U8224 (N_8224,N_1261,N_3948);
and U8225 (N_8225,N_4702,N_2618);
or U8226 (N_8226,N_3596,N_1862);
nand U8227 (N_8227,N_3121,N_3326);
nor U8228 (N_8228,N_1778,N_4586);
and U8229 (N_8229,N_4355,N_4363);
or U8230 (N_8230,N_4149,N_3268);
nor U8231 (N_8231,N_2404,N_3024);
nand U8232 (N_8232,N_1153,N_16);
xor U8233 (N_8233,N_681,N_3036);
and U8234 (N_8234,N_3656,N_3144);
nand U8235 (N_8235,N_1806,N_465);
nand U8236 (N_8236,N_62,N_319);
or U8237 (N_8237,N_3962,N_3925);
and U8238 (N_8238,N_3181,N_3706);
or U8239 (N_8239,N_3874,N_2185);
and U8240 (N_8240,N_110,N_3371);
nand U8241 (N_8241,N_2569,N_2307);
and U8242 (N_8242,N_4128,N_777);
nor U8243 (N_8243,N_4703,N_1747);
nor U8244 (N_8244,N_3071,N_129);
nand U8245 (N_8245,N_1980,N_1846);
or U8246 (N_8246,N_2505,N_4512);
or U8247 (N_8247,N_4827,N_1051);
and U8248 (N_8248,N_4705,N_740);
or U8249 (N_8249,N_3044,N_2360);
nand U8250 (N_8250,N_1502,N_1542);
xor U8251 (N_8251,N_876,N_3616);
nor U8252 (N_8252,N_3856,N_3309);
and U8253 (N_8253,N_1262,N_2065);
or U8254 (N_8254,N_2264,N_2046);
or U8255 (N_8255,N_839,N_1247);
nand U8256 (N_8256,N_4747,N_4028);
nor U8257 (N_8257,N_2919,N_4210);
or U8258 (N_8258,N_4707,N_3604);
nor U8259 (N_8259,N_3830,N_45);
or U8260 (N_8260,N_3478,N_4145);
or U8261 (N_8261,N_2629,N_1170);
nor U8262 (N_8262,N_3623,N_1083);
and U8263 (N_8263,N_4947,N_1876);
xor U8264 (N_8264,N_4673,N_3829);
and U8265 (N_8265,N_492,N_4649);
nor U8266 (N_8266,N_4061,N_2259);
nand U8267 (N_8267,N_4360,N_75);
nor U8268 (N_8268,N_1854,N_2085);
nor U8269 (N_8269,N_958,N_4138);
or U8270 (N_8270,N_2266,N_32);
nor U8271 (N_8271,N_1682,N_3079);
or U8272 (N_8272,N_2716,N_2753);
or U8273 (N_8273,N_4073,N_2108);
nor U8274 (N_8274,N_204,N_474);
and U8275 (N_8275,N_675,N_1851);
and U8276 (N_8276,N_910,N_3742);
nor U8277 (N_8277,N_3322,N_4034);
or U8278 (N_8278,N_3174,N_2236);
and U8279 (N_8279,N_878,N_245);
nor U8280 (N_8280,N_3641,N_2642);
nor U8281 (N_8281,N_1565,N_4688);
nand U8282 (N_8282,N_1327,N_610);
nand U8283 (N_8283,N_2958,N_435);
nor U8284 (N_8284,N_1323,N_3608);
or U8285 (N_8285,N_661,N_374);
nor U8286 (N_8286,N_3417,N_4653);
or U8287 (N_8287,N_3662,N_2879);
or U8288 (N_8288,N_4500,N_4352);
or U8289 (N_8289,N_2194,N_2831);
or U8290 (N_8290,N_4474,N_2938);
and U8291 (N_8291,N_4144,N_1084);
and U8292 (N_8292,N_29,N_1667);
and U8293 (N_8293,N_1888,N_87);
nor U8294 (N_8294,N_2958,N_1347);
nand U8295 (N_8295,N_4221,N_1403);
nor U8296 (N_8296,N_3960,N_2929);
nor U8297 (N_8297,N_3654,N_1361);
xnor U8298 (N_8298,N_387,N_1786);
and U8299 (N_8299,N_2366,N_3527);
nor U8300 (N_8300,N_2248,N_2953);
and U8301 (N_8301,N_1607,N_2193);
and U8302 (N_8302,N_3191,N_2128);
nor U8303 (N_8303,N_4804,N_1654);
nand U8304 (N_8304,N_1227,N_1213);
nor U8305 (N_8305,N_4001,N_4632);
nand U8306 (N_8306,N_2940,N_3788);
nor U8307 (N_8307,N_3073,N_2593);
and U8308 (N_8308,N_420,N_2413);
and U8309 (N_8309,N_967,N_3371);
nand U8310 (N_8310,N_930,N_1191);
nor U8311 (N_8311,N_3572,N_900);
nor U8312 (N_8312,N_618,N_3773);
or U8313 (N_8313,N_2792,N_3084);
nor U8314 (N_8314,N_4471,N_1542);
and U8315 (N_8315,N_895,N_470);
nor U8316 (N_8316,N_3888,N_1446);
and U8317 (N_8317,N_1816,N_1402);
or U8318 (N_8318,N_1877,N_4730);
and U8319 (N_8319,N_1161,N_754);
or U8320 (N_8320,N_47,N_4594);
nor U8321 (N_8321,N_1923,N_1092);
xor U8322 (N_8322,N_1568,N_691);
nor U8323 (N_8323,N_2738,N_741);
nor U8324 (N_8324,N_4947,N_4797);
and U8325 (N_8325,N_3679,N_2076);
or U8326 (N_8326,N_1063,N_4827);
or U8327 (N_8327,N_1928,N_1413);
or U8328 (N_8328,N_2267,N_2643);
or U8329 (N_8329,N_269,N_4846);
or U8330 (N_8330,N_2342,N_3813);
and U8331 (N_8331,N_4506,N_2465);
nor U8332 (N_8332,N_299,N_3492);
and U8333 (N_8333,N_2626,N_4676);
nand U8334 (N_8334,N_4298,N_4142);
nand U8335 (N_8335,N_3229,N_4438);
or U8336 (N_8336,N_297,N_4362);
nand U8337 (N_8337,N_3492,N_1235);
nand U8338 (N_8338,N_1141,N_3792);
and U8339 (N_8339,N_363,N_1168);
and U8340 (N_8340,N_4877,N_829);
nor U8341 (N_8341,N_875,N_1719);
and U8342 (N_8342,N_2629,N_4007);
nor U8343 (N_8343,N_417,N_2906);
nor U8344 (N_8344,N_1810,N_4805);
or U8345 (N_8345,N_4772,N_379);
and U8346 (N_8346,N_669,N_1026);
or U8347 (N_8347,N_717,N_377);
nor U8348 (N_8348,N_3272,N_1536);
or U8349 (N_8349,N_904,N_1844);
and U8350 (N_8350,N_703,N_2759);
nor U8351 (N_8351,N_4604,N_373);
nand U8352 (N_8352,N_468,N_3276);
nor U8353 (N_8353,N_4343,N_1467);
and U8354 (N_8354,N_4572,N_1073);
and U8355 (N_8355,N_1431,N_4177);
and U8356 (N_8356,N_364,N_3892);
nor U8357 (N_8357,N_1845,N_2193);
nand U8358 (N_8358,N_767,N_1489);
and U8359 (N_8359,N_1478,N_3286);
nor U8360 (N_8360,N_4810,N_4047);
nand U8361 (N_8361,N_4490,N_1761);
and U8362 (N_8362,N_3755,N_3118);
and U8363 (N_8363,N_3101,N_3413);
nand U8364 (N_8364,N_4568,N_4777);
or U8365 (N_8365,N_3037,N_4174);
nor U8366 (N_8366,N_117,N_3596);
and U8367 (N_8367,N_4923,N_4472);
xor U8368 (N_8368,N_2408,N_992);
nor U8369 (N_8369,N_4352,N_2092);
nand U8370 (N_8370,N_2671,N_4695);
nor U8371 (N_8371,N_1986,N_980);
nor U8372 (N_8372,N_2175,N_1413);
and U8373 (N_8373,N_2210,N_4441);
and U8374 (N_8374,N_1547,N_4404);
or U8375 (N_8375,N_2955,N_1189);
and U8376 (N_8376,N_1375,N_172);
or U8377 (N_8377,N_3655,N_4545);
nand U8378 (N_8378,N_328,N_1830);
or U8379 (N_8379,N_592,N_2794);
xor U8380 (N_8380,N_1355,N_2240);
xnor U8381 (N_8381,N_1312,N_2717);
nand U8382 (N_8382,N_2270,N_851);
nand U8383 (N_8383,N_1636,N_1181);
and U8384 (N_8384,N_1149,N_3603);
nor U8385 (N_8385,N_2691,N_3216);
and U8386 (N_8386,N_1766,N_1648);
nand U8387 (N_8387,N_1446,N_1343);
and U8388 (N_8388,N_169,N_2929);
and U8389 (N_8389,N_359,N_4948);
or U8390 (N_8390,N_4764,N_3047);
nor U8391 (N_8391,N_1006,N_217);
and U8392 (N_8392,N_47,N_2308);
and U8393 (N_8393,N_1919,N_1249);
nor U8394 (N_8394,N_2953,N_4951);
nor U8395 (N_8395,N_1333,N_3808);
nor U8396 (N_8396,N_3926,N_4387);
nand U8397 (N_8397,N_1725,N_586);
and U8398 (N_8398,N_1097,N_3618);
xnor U8399 (N_8399,N_756,N_931);
nand U8400 (N_8400,N_103,N_2921);
or U8401 (N_8401,N_2353,N_1261);
nor U8402 (N_8402,N_665,N_74);
nor U8403 (N_8403,N_4567,N_2533);
and U8404 (N_8404,N_4843,N_564);
or U8405 (N_8405,N_2032,N_3117);
nor U8406 (N_8406,N_1210,N_836);
or U8407 (N_8407,N_4969,N_1383);
or U8408 (N_8408,N_4483,N_3655);
and U8409 (N_8409,N_2057,N_1043);
nand U8410 (N_8410,N_71,N_2009);
or U8411 (N_8411,N_2162,N_1447);
nand U8412 (N_8412,N_233,N_2253);
and U8413 (N_8413,N_4310,N_2764);
nand U8414 (N_8414,N_4633,N_1368);
or U8415 (N_8415,N_4546,N_3233);
and U8416 (N_8416,N_2369,N_3046);
and U8417 (N_8417,N_4233,N_3778);
xor U8418 (N_8418,N_2033,N_3276);
xor U8419 (N_8419,N_3490,N_4523);
nor U8420 (N_8420,N_4041,N_4595);
or U8421 (N_8421,N_1977,N_2321);
nor U8422 (N_8422,N_2741,N_3190);
and U8423 (N_8423,N_4634,N_662);
nand U8424 (N_8424,N_3719,N_1245);
nand U8425 (N_8425,N_3869,N_3295);
and U8426 (N_8426,N_1774,N_3214);
xnor U8427 (N_8427,N_533,N_3506);
or U8428 (N_8428,N_3136,N_2902);
nand U8429 (N_8429,N_3776,N_2887);
or U8430 (N_8430,N_1433,N_4313);
and U8431 (N_8431,N_1785,N_2017);
nand U8432 (N_8432,N_2337,N_278);
nand U8433 (N_8433,N_4624,N_1915);
nor U8434 (N_8434,N_2739,N_3108);
and U8435 (N_8435,N_4090,N_4868);
xnor U8436 (N_8436,N_10,N_2304);
nor U8437 (N_8437,N_1366,N_1092);
nand U8438 (N_8438,N_2543,N_956);
nand U8439 (N_8439,N_430,N_3121);
nand U8440 (N_8440,N_2439,N_2776);
nand U8441 (N_8441,N_3558,N_2281);
or U8442 (N_8442,N_3443,N_3254);
and U8443 (N_8443,N_1478,N_4875);
and U8444 (N_8444,N_750,N_2049);
and U8445 (N_8445,N_4971,N_3848);
and U8446 (N_8446,N_161,N_3998);
nor U8447 (N_8447,N_677,N_3517);
nor U8448 (N_8448,N_4920,N_959);
or U8449 (N_8449,N_718,N_2748);
and U8450 (N_8450,N_672,N_2289);
or U8451 (N_8451,N_679,N_2393);
nand U8452 (N_8452,N_3892,N_962);
or U8453 (N_8453,N_1431,N_1954);
and U8454 (N_8454,N_4215,N_132);
nand U8455 (N_8455,N_1700,N_1376);
nor U8456 (N_8456,N_3833,N_4256);
nor U8457 (N_8457,N_83,N_2191);
nor U8458 (N_8458,N_4002,N_1772);
and U8459 (N_8459,N_2873,N_2627);
nand U8460 (N_8460,N_3096,N_1234);
xnor U8461 (N_8461,N_3146,N_1200);
or U8462 (N_8462,N_4743,N_4842);
xor U8463 (N_8463,N_2778,N_3015);
nand U8464 (N_8464,N_2094,N_1802);
nor U8465 (N_8465,N_258,N_1324);
and U8466 (N_8466,N_4190,N_642);
or U8467 (N_8467,N_1753,N_4790);
nor U8468 (N_8468,N_270,N_1949);
nand U8469 (N_8469,N_2316,N_1364);
nand U8470 (N_8470,N_4711,N_13);
and U8471 (N_8471,N_345,N_4468);
nor U8472 (N_8472,N_891,N_2656);
and U8473 (N_8473,N_743,N_888);
nor U8474 (N_8474,N_2422,N_875);
and U8475 (N_8475,N_3353,N_4793);
nor U8476 (N_8476,N_204,N_1421);
and U8477 (N_8477,N_2105,N_4583);
or U8478 (N_8478,N_2407,N_1278);
and U8479 (N_8479,N_3966,N_2094);
xor U8480 (N_8480,N_4837,N_276);
nand U8481 (N_8481,N_4242,N_2095);
or U8482 (N_8482,N_3262,N_4124);
nand U8483 (N_8483,N_1221,N_3934);
and U8484 (N_8484,N_1747,N_1150);
nand U8485 (N_8485,N_1151,N_4161);
and U8486 (N_8486,N_659,N_4896);
and U8487 (N_8487,N_331,N_519);
or U8488 (N_8488,N_4580,N_3985);
or U8489 (N_8489,N_2483,N_98);
and U8490 (N_8490,N_2516,N_960);
nand U8491 (N_8491,N_4313,N_4702);
or U8492 (N_8492,N_1982,N_4805);
nand U8493 (N_8493,N_1161,N_2900);
nor U8494 (N_8494,N_485,N_3789);
nor U8495 (N_8495,N_2413,N_2559);
nor U8496 (N_8496,N_3660,N_3685);
nand U8497 (N_8497,N_4813,N_1963);
and U8498 (N_8498,N_646,N_262);
nand U8499 (N_8499,N_1343,N_4622);
xor U8500 (N_8500,N_4533,N_1108);
and U8501 (N_8501,N_3712,N_4735);
nor U8502 (N_8502,N_2253,N_726);
nor U8503 (N_8503,N_1113,N_1758);
or U8504 (N_8504,N_4974,N_3245);
nor U8505 (N_8505,N_4930,N_1582);
and U8506 (N_8506,N_512,N_1885);
and U8507 (N_8507,N_3706,N_3118);
nor U8508 (N_8508,N_3691,N_2646);
and U8509 (N_8509,N_1335,N_389);
and U8510 (N_8510,N_2208,N_664);
and U8511 (N_8511,N_3340,N_1870);
and U8512 (N_8512,N_1429,N_4496);
or U8513 (N_8513,N_3653,N_94);
nor U8514 (N_8514,N_823,N_3454);
xnor U8515 (N_8515,N_3738,N_4737);
or U8516 (N_8516,N_2573,N_4561);
nor U8517 (N_8517,N_1621,N_2641);
or U8518 (N_8518,N_4107,N_4186);
nor U8519 (N_8519,N_1435,N_3707);
nor U8520 (N_8520,N_3595,N_1787);
or U8521 (N_8521,N_4051,N_3050);
nand U8522 (N_8522,N_962,N_2593);
or U8523 (N_8523,N_1388,N_1369);
and U8524 (N_8524,N_4169,N_4178);
and U8525 (N_8525,N_4067,N_3764);
nand U8526 (N_8526,N_1275,N_1729);
nand U8527 (N_8527,N_2036,N_324);
nand U8528 (N_8528,N_2373,N_2081);
nand U8529 (N_8529,N_1845,N_4281);
or U8530 (N_8530,N_4950,N_3489);
nor U8531 (N_8531,N_545,N_966);
and U8532 (N_8532,N_3957,N_1807);
or U8533 (N_8533,N_3443,N_4987);
nand U8534 (N_8534,N_330,N_4369);
and U8535 (N_8535,N_1782,N_255);
and U8536 (N_8536,N_1111,N_3713);
or U8537 (N_8537,N_3351,N_3040);
or U8538 (N_8538,N_2659,N_3476);
and U8539 (N_8539,N_4508,N_975);
or U8540 (N_8540,N_4953,N_1191);
or U8541 (N_8541,N_2089,N_3214);
and U8542 (N_8542,N_2629,N_1658);
nand U8543 (N_8543,N_2223,N_1799);
nor U8544 (N_8544,N_228,N_4645);
or U8545 (N_8545,N_3755,N_4335);
xor U8546 (N_8546,N_3361,N_1076);
and U8547 (N_8547,N_397,N_1141);
nand U8548 (N_8548,N_2582,N_345);
or U8549 (N_8549,N_1962,N_1405);
or U8550 (N_8550,N_4884,N_3546);
or U8551 (N_8551,N_1240,N_4377);
nand U8552 (N_8552,N_3993,N_3912);
nand U8553 (N_8553,N_4824,N_3163);
and U8554 (N_8554,N_2061,N_4274);
nand U8555 (N_8555,N_1346,N_4428);
or U8556 (N_8556,N_4154,N_3049);
and U8557 (N_8557,N_347,N_2150);
and U8558 (N_8558,N_3885,N_4238);
nand U8559 (N_8559,N_2995,N_4571);
or U8560 (N_8560,N_796,N_3951);
and U8561 (N_8561,N_4522,N_3657);
nor U8562 (N_8562,N_4303,N_3689);
and U8563 (N_8563,N_695,N_4658);
and U8564 (N_8564,N_2802,N_1707);
nor U8565 (N_8565,N_1014,N_3428);
or U8566 (N_8566,N_4619,N_4857);
nand U8567 (N_8567,N_167,N_2887);
or U8568 (N_8568,N_3307,N_1218);
or U8569 (N_8569,N_1841,N_1157);
or U8570 (N_8570,N_2201,N_3725);
or U8571 (N_8571,N_4536,N_2969);
nand U8572 (N_8572,N_2118,N_4328);
xnor U8573 (N_8573,N_4544,N_3046);
and U8574 (N_8574,N_2739,N_907);
nor U8575 (N_8575,N_465,N_1825);
nor U8576 (N_8576,N_733,N_2706);
and U8577 (N_8577,N_297,N_1838);
nand U8578 (N_8578,N_27,N_2229);
and U8579 (N_8579,N_4013,N_3532);
or U8580 (N_8580,N_1913,N_3541);
nand U8581 (N_8581,N_502,N_1440);
nand U8582 (N_8582,N_2930,N_3570);
and U8583 (N_8583,N_2560,N_406);
and U8584 (N_8584,N_683,N_4353);
nand U8585 (N_8585,N_2524,N_3673);
nor U8586 (N_8586,N_3249,N_1904);
nand U8587 (N_8587,N_3489,N_4741);
or U8588 (N_8588,N_2486,N_4704);
or U8589 (N_8589,N_579,N_2909);
nand U8590 (N_8590,N_1495,N_593);
nand U8591 (N_8591,N_2756,N_2578);
nand U8592 (N_8592,N_1711,N_1772);
nand U8593 (N_8593,N_1694,N_3676);
nand U8594 (N_8594,N_4897,N_3922);
nor U8595 (N_8595,N_1196,N_2583);
or U8596 (N_8596,N_3080,N_2510);
nor U8597 (N_8597,N_1392,N_4525);
or U8598 (N_8598,N_4485,N_1356);
nor U8599 (N_8599,N_4370,N_4491);
or U8600 (N_8600,N_2236,N_4751);
or U8601 (N_8601,N_4974,N_4306);
or U8602 (N_8602,N_4218,N_4880);
and U8603 (N_8603,N_308,N_4218);
nor U8604 (N_8604,N_941,N_1468);
nand U8605 (N_8605,N_3875,N_4254);
and U8606 (N_8606,N_1130,N_4291);
and U8607 (N_8607,N_374,N_517);
nor U8608 (N_8608,N_4235,N_4366);
nand U8609 (N_8609,N_4437,N_1861);
and U8610 (N_8610,N_2797,N_160);
and U8611 (N_8611,N_789,N_1112);
and U8612 (N_8612,N_2613,N_3402);
nand U8613 (N_8613,N_2866,N_435);
nand U8614 (N_8614,N_139,N_1338);
and U8615 (N_8615,N_4888,N_2083);
nand U8616 (N_8616,N_4712,N_3262);
nand U8617 (N_8617,N_280,N_936);
and U8618 (N_8618,N_1442,N_2802);
and U8619 (N_8619,N_4156,N_4266);
nor U8620 (N_8620,N_2725,N_1570);
nand U8621 (N_8621,N_4252,N_3857);
nor U8622 (N_8622,N_1342,N_2519);
xor U8623 (N_8623,N_1932,N_453);
or U8624 (N_8624,N_3736,N_1088);
or U8625 (N_8625,N_3074,N_837);
and U8626 (N_8626,N_162,N_443);
nor U8627 (N_8627,N_3311,N_3170);
and U8628 (N_8628,N_945,N_2378);
nand U8629 (N_8629,N_3329,N_2339);
and U8630 (N_8630,N_1815,N_4241);
or U8631 (N_8631,N_3081,N_1302);
or U8632 (N_8632,N_3802,N_3197);
nor U8633 (N_8633,N_3731,N_3727);
nor U8634 (N_8634,N_3264,N_3252);
and U8635 (N_8635,N_2449,N_198);
or U8636 (N_8636,N_4396,N_192);
nand U8637 (N_8637,N_342,N_873);
or U8638 (N_8638,N_1862,N_1266);
and U8639 (N_8639,N_2740,N_3435);
nor U8640 (N_8640,N_4534,N_847);
nor U8641 (N_8641,N_3653,N_2159);
or U8642 (N_8642,N_4025,N_4277);
nand U8643 (N_8643,N_4379,N_4387);
nand U8644 (N_8644,N_4881,N_4842);
and U8645 (N_8645,N_4201,N_2356);
or U8646 (N_8646,N_3451,N_480);
nor U8647 (N_8647,N_4022,N_1735);
or U8648 (N_8648,N_204,N_3543);
nand U8649 (N_8649,N_1111,N_3686);
and U8650 (N_8650,N_3031,N_2246);
and U8651 (N_8651,N_2579,N_240);
xnor U8652 (N_8652,N_4164,N_1084);
and U8653 (N_8653,N_3149,N_3424);
or U8654 (N_8654,N_4665,N_4751);
nand U8655 (N_8655,N_3303,N_2850);
and U8656 (N_8656,N_4365,N_521);
and U8657 (N_8657,N_1186,N_3340);
and U8658 (N_8658,N_3104,N_4957);
nor U8659 (N_8659,N_4979,N_4846);
nor U8660 (N_8660,N_227,N_4845);
and U8661 (N_8661,N_2397,N_863);
nand U8662 (N_8662,N_4468,N_849);
or U8663 (N_8663,N_872,N_2411);
nor U8664 (N_8664,N_2401,N_4840);
nand U8665 (N_8665,N_1209,N_2102);
and U8666 (N_8666,N_224,N_3135);
xor U8667 (N_8667,N_4154,N_2000);
and U8668 (N_8668,N_1906,N_2478);
or U8669 (N_8669,N_4482,N_1771);
or U8670 (N_8670,N_4466,N_1232);
nand U8671 (N_8671,N_2247,N_2142);
or U8672 (N_8672,N_1586,N_514);
or U8673 (N_8673,N_1936,N_2793);
or U8674 (N_8674,N_4782,N_4374);
or U8675 (N_8675,N_1437,N_1910);
nand U8676 (N_8676,N_3232,N_3446);
or U8677 (N_8677,N_2632,N_3959);
or U8678 (N_8678,N_3846,N_4510);
or U8679 (N_8679,N_718,N_3257);
nand U8680 (N_8680,N_4807,N_158);
or U8681 (N_8681,N_4434,N_4250);
nand U8682 (N_8682,N_2795,N_3779);
nand U8683 (N_8683,N_3449,N_3023);
or U8684 (N_8684,N_3450,N_4328);
xnor U8685 (N_8685,N_3823,N_4885);
or U8686 (N_8686,N_4666,N_1470);
and U8687 (N_8687,N_62,N_1726);
nor U8688 (N_8688,N_1274,N_2898);
and U8689 (N_8689,N_4185,N_1275);
nor U8690 (N_8690,N_3854,N_309);
or U8691 (N_8691,N_1717,N_236);
or U8692 (N_8692,N_3611,N_2201);
or U8693 (N_8693,N_856,N_2021);
nor U8694 (N_8694,N_1964,N_4850);
nor U8695 (N_8695,N_1108,N_2126);
nor U8696 (N_8696,N_3942,N_4733);
nor U8697 (N_8697,N_4483,N_1601);
and U8698 (N_8698,N_196,N_840);
and U8699 (N_8699,N_1771,N_918);
nor U8700 (N_8700,N_328,N_4759);
nand U8701 (N_8701,N_872,N_418);
or U8702 (N_8702,N_3820,N_2355);
nor U8703 (N_8703,N_3704,N_2372);
nand U8704 (N_8704,N_2655,N_2197);
or U8705 (N_8705,N_4587,N_4295);
or U8706 (N_8706,N_466,N_2527);
and U8707 (N_8707,N_36,N_426);
nor U8708 (N_8708,N_1770,N_886);
nor U8709 (N_8709,N_1442,N_954);
nand U8710 (N_8710,N_2749,N_2001);
and U8711 (N_8711,N_3875,N_1037);
xor U8712 (N_8712,N_4511,N_388);
and U8713 (N_8713,N_2936,N_532);
nand U8714 (N_8714,N_3814,N_941);
nand U8715 (N_8715,N_163,N_1590);
and U8716 (N_8716,N_4238,N_4490);
or U8717 (N_8717,N_1765,N_536);
or U8718 (N_8718,N_4860,N_4519);
or U8719 (N_8719,N_3891,N_1259);
and U8720 (N_8720,N_4706,N_4360);
nor U8721 (N_8721,N_687,N_2016);
nand U8722 (N_8722,N_2748,N_2116);
nand U8723 (N_8723,N_1722,N_2342);
or U8724 (N_8724,N_3519,N_4568);
nor U8725 (N_8725,N_1785,N_2964);
nand U8726 (N_8726,N_4002,N_3660);
nor U8727 (N_8727,N_1021,N_4137);
or U8728 (N_8728,N_2927,N_4602);
nor U8729 (N_8729,N_2392,N_4028);
and U8730 (N_8730,N_2847,N_2253);
and U8731 (N_8731,N_1748,N_1924);
nor U8732 (N_8732,N_1982,N_4371);
and U8733 (N_8733,N_3473,N_3325);
nor U8734 (N_8734,N_2631,N_1910);
and U8735 (N_8735,N_3413,N_1556);
nor U8736 (N_8736,N_1413,N_3783);
and U8737 (N_8737,N_3949,N_4458);
nor U8738 (N_8738,N_4047,N_3874);
or U8739 (N_8739,N_2032,N_4249);
nand U8740 (N_8740,N_2226,N_629);
nand U8741 (N_8741,N_4241,N_226);
and U8742 (N_8742,N_4229,N_3764);
nor U8743 (N_8743,N_1931,N_1273);
or U8744 (N_8744,N_3879,N_1139);
nor U8745 (N_8745,N_3913,N_185);
and U8746 (N_8746,N_423,N_3510);
and U8747 (N_8747,N_1184,N_3434);
nor U8748 (N_8748,N_3531,N_380);
nor U8749 (N_8749,N_602,N_1612);
and U8750 (N_8750,N_171,N_587);
or U8751 (N_8751,N_4212,N_261);
or U8752 (N_8752,N_139,N_2942);
or U8753 (N_8753,N_3995,N_262);
nor U8754 (N_8754,N_3966,N_4771);
nor U8755 (N_8755,N_4024,N_2015);
and U8756 (N_8756,N_952,N_4990);
and U8757 (N_8757,N_2509,N_3394);
nor U8758 (N_8758,N_158,N_2424);
nand U8759 (N_8759,N_967,N_255);
or U8760 (N_8760,N_3356,N_776);
or U8761 (N_8761,N_3980,N_2497);
or U8762 (N_8762,N_501,N_3919);
and U8763 (N_8763,N_1905,N_3780);
or U8764 (N_8764,N_138,N_3149);
and U8765 (N_8765,N_4939,N_4929);
nand U8766 (N_8766,N_1413,N_1796);
nand U8767 (N_8767,N_3564,N_4358);
or U8768 (N_8768,N_2244,N_1378);
and U8769 (N_8769,N_894,N_608);
nand U8770 (N_8770,N_516,N_4091);
and U8771 (N_8771,N_1455,N_3573);
and U8772 (N_8772,N_849,N_916);
nand U8773 (N_8773,N_4151,N_2825);
nor U8774 (N_8774,N_2294,N_1320);
xnor U8775 (N_8775,N_2038,N_832);
nand U8776 (N_8776,N_1613,N_729);
nor U8777 (N_8777,N_4852,N_1554);
and U8778 (N_8778,N_2507,N_1456);
or U8779 (N_8779,N_1611,N_4166);
nand U8780 (N_8780,N_2606,N_29);
nor U8781 (N_8781,N_728,N_2368);
or U8782 (N_8782,N_4048,N_2033);
or U8783 (N_8783,N_3643,N_4299);
and U8784 (N_8784,N_3077,N_263);
or U8785 (N_8785,N_952,N_4925);
and U8786 (N_8786,N_3272,N_3171);
or U8787 (N_8787,N_1592,N_4613);
nand U8788 (N_8788,N_607,N_353);
nand U8789 (N_8789,N_1213,N_2664);
nand U8790 (N_8790,N_1518,N_652);
or U8791 (N_8791,N_254,N_2166);
and U8792 (N_8792,N_2651,N_1263);
nand U8793 (N_8793,N_4439,N_3675);
and U8794 (N_8794,N_1810,N_2963);
nand U8795 (N_8795,N_1135,N_556);
nand U8796 (N_8796,N_1756,N_1746);
nor U8797 (N_8797,N_4040,N_3921);
nor U8798 (N_8798,N_786,N_4041);
and U8799 (N_8799,N_1092,N_4119);
and U8800 (N_8800,N_1462,N_238);
nor U8801 (N_8801,N_3158,N_3204);
or U8802 (N_8802,N_307,N_3979);
and U8803 (N_8803,N_1428,N_3855);
nand U8804 (N_8804,N_1445,N_1783);
or U8805 (N_8805,N_2762,N_1509);
nand U8806 (N_8806,N_3370,N_1942);
nand U8807 (N_8807,N_1277,N_3386);
or U8808 (N_8808,N_4484,N_225);
nand U8809 (N_8809,N_1593,N_4530);
nand U8810 (N_8810,N_3025,N_3152);
or U8811 (N_8811,N_4605,N_2406);
nand U8812 (N_8812,N_1117,N_571);
nor U8813 (N_8813,N_3294,N_2887);
xor U8814 (N_8814,N_3960,N_4197);
nor U8815 (N_8815,N_962,N_3666);
nor U8816 (N_8816,N_3871,N_1626);
xnor U8817 (N_8817,N_309,N_3866);
nor U8818 (N_8818,N_3987,N_3080);
nand U8819 (N_8819,N_1620,N_4049);
nor U8820 (N_8820,N_3571,N_4139);
or U8821 (N_8821,N_2175,N_969);
nand U8822 (N_8822,N_4414,N_2213);
nor U8823 (N_8823,N_4815,N_1303);
or U8824 (N_8824,N_3034,N_2466);
nor U8825 (N_8825,N_2167,N_381);
nor U8826 (N_8826,N_2679,N_4826);
nand U8827 (N_8827,N_4073,N_2411);
nor U8828 (N_8828,N_894,N_3482);
and U8829 (N_8829,N_2369,N_1608);
and U8830 (N_8830,N_3892,N_515);
or U8831 (N_8831,N_2766,N_1060);
and U8832 (N_8832,N_391,N_2489);
and U8833 (N_8833,N_4668,N_3760);
or U8834 (N_8834,N_3883,N_4343);
nor U8835 (N_8835,N_4463,N_1776);
nand U8836 (N_8836,N_1812,N_4642);
nand U8837 (N_8837,N_2074,N_1544);
or U8838 (N_8838,N_2730,N_1086);
nand U8839 (N_8839,N_2079,N_3000);
nor U8840 (N_8840,N_2576,N_1734);
nand U8841 (N_8841,N_1824,N_4956);
nor U8842 (N_8842,N_1617,N_4580);
nand U8843 (N_8843,N_204,N_2569);
or U8844 (N_8844,N_3091,N_4123);
or U8845 (N_8845,N_1184,N_3631);
or U8846 (N_8846,N_2361,N_3224);
and U8847 (N_8847,N_3674,N_241);
or U8848 (N_8848,N_12,N_3057);
nor U8849 (N_8849,N_2706,N_1834);
and U8850 (N_8850,N_2985,N_421);
and U8851 (N_8851,N_152,N_4396);
nor U8852 (N_8852,N_4547,N_3293);
and U8853 (N_8853,N_1930,N_2754);
nor U8854 (N_8854,N_1543,N_3314);
nand U8855 (N_8855,N_2273,N_4844);
or U8856 (N_8856,N_4604,N_1678);
or U8857 (N_8857,N_3598,N_517);
and U8858 (N_8858,N_2218,N_4477);
nor U8859 (N_8859,N_4912,N_3082);
nor U8860 (N_8860,N_845,N_2055);
and U8861 (N_8861,N_4540,N_3169);
nand U8862 (N_8862,N_4012,N_3723);
nor U8863 (N_8863,N_2677,N_1790);
and U8864 (N_8864,N_3004,N_2594);
nand U8865 (N_8865,N_3937,N_2576);
nand U8866 (N_8866,N_4991,N_3891);
nor U8867 (N_8867,N_4553,N_2915);
and U8868 (N_8868,N_666,N_3062);
and U8869 (N_8869,N_2133,N_3880);
or U8870 (N_8870,N_4874,N_4348);
and U8871 (N_8871,N_640,N_720);
nor U8872 (N_8872,N_266,N_2749);
nor U8873 (N_8873,N_1787,N_2111);
and U8874 (N_8874,N_2406,N_1514);
nand U8875 (N_8875,N_282,N_1681);
xor U8876 (N_8876,N_1079,N_231);
and U8877 (N_8877,N_2314,N_1050);
and U8878 (N_8878,N_3561,N_1494);
nand U8879 (N_8879,N_2764,N_4090);
nor U8880 (N_8880,N_2,N_2795);
or U8881 (N_8881,N_2472,N_1841);
nor U8882 (N_8882,N_2283,N_3038);
and U8883 (N_8883,N_2734,N_583);
and U8884 (N_8884,N_1191,N_1323);
nand U8885 (N_8885,N_2788,N_3398);
and U8886 (N_8886,N_745,N_0);
and U8887 (N_8887,N_4250,N_4564);
nand U8888 (N_8888,N_4708,N_1997);
and U8889 (N_8889,N_3948,N_1880);
and U8890 (N_8890,N_4781,N_3746);
nand U8891 (N_8891,N_2543,N_45);
nand U8892 (N_8892,N_221,N_1609);
nand U8893 (N_8893,N_178,N_738);
or U8894 (N_8894,N_1442,N_1794);
xnor U8895 (N_8895,N_2218,N_805);
nand U8896 (N_8896,N_1761,N_1332);
and U8897 (N_8897,N_1036,N_4486);
nor U8898 (N_8898,N_264,N_1003);
nor U8899 (N_8899,N_3906,N_76);
nand U8900 (N_8900,N_4136,N_13);
nor U8901 (N_8901,N_2894,N_2846);
or U8902 (N_8902,N_4024,N_1728);
nor U8903 (N_8903,N_1671,N_2178);
nand U8904 (N_8904,N_4710,N_820);
nor U8905 (N_8905,N_1533,N_4951);
nor U8906 (N_8906,N_679,N_4724);
and U8907 (N_8907,N_4194,N_66);
nor U8908 (N_8908,N_3854,N_2883);
and U8909 (N_8909,N_2468,N_1650);
nand U8910 (N_8910,N_2831,N_56);
nor U8911 (N_8911,N_1857,N_4453);
and U8912 (N_8912,N_4292,N_2463);
nor U8913 (N_8913,N_248,N_2991);
and U8914 (N_8914,N_961,N_2650);
or U8915 (N_8915,N_3751,N_1911);
or U8916 (N_8916,N_377,N_4423);
nand U8917 (N_8917,N_3915,N_783);
nand U8918 (N_8918,N_4383,N_4239);
nand U8919 (N_8919,N_992,N_4663);
and U8920 (N_8920,N_955,N_3115);
nor U8921 (N_8921,N_1567,N_4119);
and U8922 (N_8922,N_3018,N_1224);
nor U8923 (N_8923,N_3905,N_4641);
nand U8924 (N_8924,N_1543,N_2905);
and U8925 (N_8925,N_1325,N_2510);
or U8926 (N_8926,N_1458,N_21);
xor U8927 (N_8927,N_359,N_2261);
nand U8928 (N_8928,N_1698,N_1766);
nor U8929 (N_8929,N_2252,N_4319);
nor U8930 (N_8930,N_4810,N_777);
and U8931 (N_8931,N_4474,N_397);
or U8932 (N_8932,N_4875,N_1651);
and U8933 (N_8933,N_3666,N_4616);
nand U8934 (N_8934,N_1111,N_2477);
or U8935 (N_8935,N_1732,N_3076);
xor U8936 (N_8936,N_3779,N_4144);
nor U8937 (N_8937,N_3129,N_3850);
and U8938 (N_8938,N_1231,N_331);
nand U8939 (N_8939,N_710,N_4517);
nand U8940 (N_8940,N_4673,N_2413);
or U8941 (N_8941,N_2412,N_788);
or U8942 (N_8942,N_3024,N_3637);
and U8943 (N_8943,N_671,N_3306);
and U8944 (N_8944,N_827,N_4158);
or U8945 (N_8945,N_1488,N_66);
and U8946 (N_8946,N_3175,N_4500);
nor U8947 (N_8947,N_4845,N_4119);
nand U8948 (N_8948,N_3508,N_821);
nand U8949 (N_8949,N_20,N_3099);
nand U8950 (N_8950,N_4415,N_2372);
nand U8951 (N_8951,N_204,N_2128);
nor U8952 (N_8952,N_1090,N_3466);
nor U8953 (N_8953,N_2409,N_3570);
nor U8954 (N_8954,N_3314,N_4825);
and U8955 (N_8955,N_3036,N_4699);
nand U8956 (N_8956,N_78,N_3564);
or U8957 (N_8957,N_4264,N_1042);
nand U8958 (N_8958,N_1370,N_2651);
and U8959 (N_8959,N_566,N_2711);
or U8960 (N_8960,N_4237,N_1828);
nand U8961 (N_8961,N_4333,N_4252);
nand U8962 (N_8962,N_2010,N_4760);
or U8963 (N_8963,N_286,N_3538);
and U8964 (N_8964,N_354,N_4122);
or U8965 (N_8965,N_4877,N_4849);
nor U8966 (N_8966,N_3928,N_3346);
nor U8967 (N_8967,N_2412,N_1639);
and U8968 (N_8968,N_3445,N_4988);
nand U8969 (N_8969,N_3314,N_3469);
and U8970 (N_8970,N_2809,N_3613);
or U8971 (N_8971,N_1441,N_4407);
and U8972 (N_8972,N_9,N_3247);
and U8973 (N_8973,N_4424,N_2937);
nand U8974 (N_8974,N_3447,N_4522);
and U8975 (N_8975,N_525,N_3376);
or U8976 (N_8976,N_2598,N_3498);
nor U8977 (N_8977,N_2692,N_2658);
nor U8978 (N_8978,N_4308,N_2634);
xor U8979 (N_8979,N_1288,N_171);
nand U8980 (N_8980,N_4922,N_4148);
or U8981 (N_8981,N_1992,N_4671);
nand U8982 (N_8982,N_304,N_3778);
nand U8983 (N_8983,N_1794,N_1653);
and U8984 (N_8984,N_4547,N_741);
nand U8985 (N_8985,N_3128,N_2066);
or U8986 (N_8986,N_222,N_3901);
nor U8987 (N_8987,N_225,N_3718);
nand U8988 (N_8988,N_929,N_1909);
or U8989 (N_8989,N_4210,N_4279);
or U8990 (N_8990,N_707,N_2033);
or U8991 (N_8991,N_528,N_4375);
or U8992 (N_8992,N_3456,N_4365);
nor U8993 (N_8993,N_3045,N_3973);
and U8994 (N_8994,N_1127,N_1662);
or U8995 (N_8995,N_532,N_1913);
and U8996 (N_8996,N_4516,N_3683);
nand U8997 (N_8997,N_2753,N_3069);
or U8998 (N_8998,N_1830,N_744);
nand U8999 (N_8999,N_161,N_3438);
nor U9000 (N_9000,N_81,N_2267);
and U9001 (N_9001,N_3467,N_577);
nand U9002 (N_9002,N_1265,N_3509);
or U9003 (N_9003,N_7,N_3182);
and U9004 (N_9004,N_1322,N_2928);
and U9005 (N_9005,N_4265,N_3939);
and U9006 (N_9006,N_1842,N_232);
and U9007 (N_9007,N_675,N_2369);
or U9008 (N_9008,N_4862,N_4104);
nand U9009 (N_9009,N_2811,N_904);
or U9010 (N_9010,N_4392,N_3891);
xnor U9011 (N_9011,N_323,N_4434);
and U9012 (N_9012,N_1178,N_4738);
or U9013 (N_9013,N_3837,N_397);
or U9014 (N_9014,N_1595,N_3316);
nor U9015 (N_9015,N_3689,N_66);
xnor U9016 (N_9016,N_977,N_3346);
nor U9017 (N_9017,N_1090,N_2223);
and U9018 (N_9018,N_75,N_1395);
or U9019 (N_9019,N_1128,N_3126);
nand U9020 (N_9020,N_4951,N_2232);
nor U9021 (N_9021,N_4671,N_2778);
nor U9022 (N_9022,N_4504,N_3885);
nor U9023 (N_9023,N_996,N_3028);
nor U9024 (N_9024,N_1365,N_2332);
nor U9025 (N_9025,N_4800,N_4204);
nand U9026 (N_9026,N_481,N_928);
and U9027 (N_9027,N_4317,N_1219);
nand U9028 (N_9028,N_1864,N_1369);
nand U9029 (N_9029,N_868,N_1224);
and U9030 (N_9030,N_1539,N_3218);
nor U9031 (N_9031,N_4407,N_3452);
nor U9032 (N_9032,N_2192,N_1497);
and U9033 (N_9033,N_3636,N_4349);
and U9034 (N_9034,N_1331,N_3865);
and U9035 (N_9035,N_4723,N_972);
and U9036 (N_9036,N_1753,N_1474);
or U9037 (N_9037,N_3112,N_1331);
nand U9038 (N_9038,N_1014,N_3948);
and U9039 (N_9039,N_4677,N_1954);
and U9040 (N_9040,N_1933,N_2572);
or U9041 (N_9041,N_3551,N_291);
nand U9042 (N_9042,N_1675,N_1632);
and U9043 (N_9043,N_819,N_2254);
and U9044 (N_9044,N_405,N_3661);
or U9045 (N_9045,N_0,N_1369);
nor U9046 (N_9046,N_1077,N_2098);
nand U9047 (N_9047,N_802,N_1325);
or U9048 (N_9048,N_279,N_2920);
nand U9049 (N_9049,N_552,N_1004);
nor U9050 (N_9050,N_3326,N_1616);
nand U9051 (N_9051,N_4715,N_603);
and U9052 (N_9052,N_4717,N_508);
and U9053 (N_9053,N_3984,N_3218);
or U9054 (N_9054,N_4931,N_4907);
nand U9055 (N_9055,N_307,N_4856);
nor U9056 (N_9056,N_339,N_3125);
and U9057 (N_9057,N_1906,N_676);
nand U9058 (N_9058,N_3810,N_4755);
and U9059 (N_9059,N_1941,N_4035);
and U9060 (N_9060,N_630,N_1344);
nand U9061 (N_9061,N_1378,N_1909);
nor U9062 (N_9062,N_2964,N_1932);
and U9063 (N_9063,N_2413,N_3354);
xnor U9064 (N_9064,N_1013,N_2481);
xor U9065 (N_9065,N_4134,N_3686);
nand U9066 (N_9066,N_3563,N_2814);
nor U9067 (N_9067,N_2149,N_3899);
nand U9068 (N_9068,N_4797,N_2056);
nand U9069 (N_9069,N_943,N_823);
or U9070 (N_9070,N_2815,N_1972);
nand U9071 (N_9071,N_3904,N_4939);
nor U9072 (N_9072,N_4827,N_3343);
nand U9073 (N_9073,N_4490,N_2239);
xnor U9074 (N_9074,N_2718,N_2988);
nand U9075 (N_9075,N_4558,N_3215);
nor U9076 (N_9076,N_1765,N_4025);
and U9077 (N_9077,N_14,N_2504);
or U9078 (N_9078,N_3020,N_1963);
and U9079 (N_9079,N_3370,N_2256);
nor U9080 (N_9080,N_3276,N_722);
or U9081 (N_9081,N_1668,N_1677);
nor U9082 (N_9082,N_1394,N_1495);
and U9083 (N_9083,N_4255,N_1930);
and U9084 (N_9084,N_540,N_4569);
xor U9085 (N_9085,N_760,N_3449);
nor U9086 (N_9086,N_2513,N_4314);
nand U9087 (N_9087,N_3962,N_4679);
nor U9088 (N_9088,N_4626,N_3110);
nand U9089 (N_9089,N_4282,N_1454);
or U9090 (N_9090,N_1323,N_192);
or U9091 (N_9091,N_740,N_2734);
or U9092 (N_9092,N_396,N_416);
nor U9093 (N_9093,N_2968,N_1718);
nor U9094 (N_9094,N_668,N_3422);
or U9095 (N_9095,N_4391,N_4357);
nor U9096 (N_9096,N_2233,N_148);
or U9097 (N_9097,N_2783,N_3549);
or U9098 (N_9098,N_1705,N_2801);
nor U9099 (N_9099,N_2429,N_1474);
and U9100 (N_9100,N_4161,N_1255);
or U9101 (N_9101,N_1814,N_2715);
or U9102 (N_9102,N_249,N_74);
and U9103 (N_9103,N_27,N_3614);
nand U9104 (N_9104,N_1393,N_448);
nor U9105 (N_9105,N_1890,N_233);
and U9106 (N_9106,N_2637,N_2950);
nand U9107 (N_9107,N_3786,N_130);
and U9108 (N_9108,N_3308,N_953);
and U9109 (N_9109,N_1600,N_4587);
nor U9110 (N_9110,N_3615,N_2554);
nor U9111 (N_9111,N_2901,N_4675);
nor U9112 (N_9112,N_4144,N_2263);
or U9113 (N_9113,N_3068,N_3959);
nand U9114 (N_9114,N_3621,N_4879);
and U9115 (N_9115,N_1211,N_2542);
nand U9116 (N_9116,N_2165,N_1156);
nand U9117 (N_9117,N_3579,N_3017);
or U9118 (N_9118,N_3065,N_2118);
nor U9119 (N_9119,N_875,N_612);
or U9120 (N_9120,N_711,N_102);
or U9121 (N_9121,N_498,N_1994);
xnor U9122 (N_9122,N_4246,N_3050);
nor U9123 (N_9123,N_4336,N_1700);
or U9124 (N_9124,N_4903,N_3914);
or U9125 (N_9125,N_3735,N_4668);
or U9126 (N_9126,N_1753,N_4150);
nand U9127 (N_9127,N_4527,N_3707);
and U9128 (N_9128,N_431,N_371);
or U9129 (N_9129,N_4508,N_1351);
nand U9130 (N_9130,N_4643,N_2835);
nand U9131 (N_9131,N_4449,N_2989);
nor U9132 (N_9132,N_641,N_4754);
nand U9133 (N_9133,N_1359,N_2040);
or U9134 (N_9134,N_2989,N_453);
and U9135 (N_9135,N_1668,N_516);
xnor U9136 (N_9136,N_4429,N_1365);
nor U9137 (N_9137,N_3815,N_1312);
nor U9138 (N_9138,N_3368,N_350);
or U9139 (N_9139,N_876,N_15);
nor U9140 (N_9140,N_992,N_1764);
nand U9141 (N_9141,N_285,N_1612);
nand U9142 (N_9142,N_1276,N_3598);
nand U9143 (N_9143,N_4262,N_4939);
nand U9144 (N_9144,N_3729,N_134);
and U9145 (N_9145,N_3899,N_3640);
nand U9146 (N_9146,N_4946,N_398);
and U9147 (N_9147,N_1031,N_4767);
nand U9148 (N_9148,N_2443,N_2543);
nor U9149 (N_9149,N_237,N_3295);
nand U9150 (N_9150,N_2049,N_854);
nor U9151 (N_9151,N_3194,N_213);
nor U9152 (N_9152,N_2152,N_611);
nor U9153 (N_9153,N_4557,N_1021);
nand U9154 (N_9154,N_3212,N_3701);
and U9155 (N_9155,N_2141,N_3874);
or U9156 (N_9156,N_3979,N_2356);
and U9157 (N_9157,N_4196,N_241);
and U9158 (N_9158,N_4732,N_3841);
nand U9159 (N_9159,N_2060,N_3380);
nand U9160 (N_9160,N_396,N_4139);
xor U9161 (N_9161,N_3825,N_1552);
nand U9162 (N_9162,N_2941,N_519);
nand U9163 (N_9163,N_142,N_1843);
nor U9164 (N_9164,N_265,N_2266);
or U9165 (N_9165,N_3242,N_1386);
or U9166 (N_9166,N_4042,N_1190);
and U9167 (N_9167,N_1120,N_1615);
and U9168 (N_9168,N_3873,N_3896);
nand U9169 (N_9169,N_3223,N_1701);
or U9170 (N_9170,N_3808,N_2721);
or U9171 (N_9171,N_2169,N_3405);
and U9172 (N_9172,N_622,N_1803);
nor U9173 (N_9173,N_2434,N_1798);
nand U9174 (N_9174,N_4004,N_4022);
or U9175 (N_9175,N_2862,N_2941);
xnor U9176 (N_9176,N_1371,N_768);
nand U9177 (N_9177,N_3542,N_3691);
nor U9178 (N_9178,N_3703,N_2180);
nand U9179 (N_9179,N_3056,N_4627);
nand U9180 (N_9180,N_491,N_3432);
nor U9181 (N_9181,N_3644,N_1376);
and U9182 (N_9182,N_2656,N_4961);
and U9183 (N_9183,N_2771,N_2111);
nand U9184 (N_9184,N_4035,N_1574);
or U9185 (N_9185,N_926,N_1584);
nor U9186 (N_9186,N_1573,N_3874);
nor U9187 (N_9187,N_2227,N_124);
nand U9188 (N_9188,N_664,N_3540);
or U9189 (N_9189,N_1580,N_4408);
nor U9190 (N_9190,N_2765,N_947);
nand U9191 (N_9191,N_2889,N_4948);
or U9192 (N_9192,N_767,N_2371);
nor U9193 (N_9193,N_204,N_4322);
nand U9194 (N_9194,N_2852,N_2716);
or U9195 (N_9195,N_797,N_1752);
and U9196 (N_9196,N_924,N_2387);
nand U9197 (N_9197,N_2570,N_4859);
nor U9198 (N_9198,N_2053,N_2006);
or U9199 (N_9199,N_3368,N_300);
nand U9200 (N_9200,N_425,N_2186);
nor U9201 (N_9201,N_3039,N_1861);
nor U9202 (N_9202,N_407,N_3030);
nor U9203 (N_9203,N_3434,N_2191);
nand U9204 (N_9204,N_2801,N_2752);
and U9205 (N_9205,N_49,N_4982);
nand U9206 (N_9206,N_2557,N_1969);
nor U9207 (N_9207,N_1482,N_1156);
or U9208 (N_9208,N_4319,N_481);
or U9209 (N_9209,N_2779,N_3348);
nand U9210 (N_9210,N_2228,N_59);
or U9211 (N_9211,N_2778,N_2488);
nor U9212 (N_9212,N_1971,N_1354);
and U9213 (N_9213,N_3317,N_4568);
and U9214 (N_9214,N_3933,N_4708);
and U9215 (N_9215,N_3415,N_2805);
nor U9216 (N_9216,N_1644,N_136);
and U9217 (N_9217,N_1396,N_559);
or U9218 (N_9218,N_310,N_4638);
nand U9219 (N_9219,N_2182,N_4535);
nand U9220 (N_9220,N_2133,N_4064);
xnor U9221 (N_9221,N_3731,N_547);
nand U9222 (N_9222,N_4192,N_3862);
and U9223 (N_9223,N_1287,N_1317);
and U9224 (N_9224,N_523,N_3877);
and U9225 (N_9225,N_4088,N_2013);
nor U9226 (N_9226,N_883,N_3954);
nor U9227 (N_9227,N_3011,N_4922);
or U9228 (N_9228,N_321,N_287);
and U9229 (N_9229,N_3584,N_1081);
or U9230 (N_9230,N_481,N_2036);
or U9231 (N_9231,N_4942,N_4069);
nand U9232 (N_9232,N_2147,N_4591);
or U9233 (N_9233,N_343,N_1052);
or U9234 (N_9234,N_1852,N_3418);
nor U9235 (N_9235,N_1778,N_2946);
nor U9236 (N_9236,N_1556,N_2638);
and U9237 (N_9237,N_3062,N_1056);
or U9238 (N_9238,N_955,N_2903);
and U9239 (N_9239,N_453,N_870);
nand U9240 (N_9240,N_2921,N_2738);
and U9241 (N_9241,N_4369,N_4882);
and U9242 (N_9242,N_2176,N_4125);
and U9243 (N_9243,N_1891,N_300);
nand U9244 (N_9244,N_106,N_3967);
nand U9245 (N_9245,N_208,N_4944);
nor U9246 (N_9246,N_46,N_3556);
or U9247 (N_9247,N_3164,N_713);
or U9248 (N_9248,N_4578,N_2346);
nor U9249 (N_9249,N_2470,N_4418);
or U9250 (N_9250,N_4634,N_921);
nor U9251 (N_9251,N_2931,N_2956);
or U9252 (N_9252,N_1222,N_2456);
and U9253 (N_9253,N_3549,N_1174);
and U9254 (N_9254,N_2683,N_4969);
or U9255 (N_9255,N_4536,N_1865);
and U9256 (N_9256,N_4082,N_4101);
or U9257 (N_9257,N_788,N_3735);
nand U9258 (N_9258,N_3617,N_2676);
or U9259 (N_9259,N_4224,N_1502);
and U9260 (N_9260,N_2716,N_1723);
nand U9261 (N_9261,N_4052,N_3589);
nand U9262 (N_9262,N_4210,N_2772);
or U9263 (N_9263,N_610,N_1219);
nand U9264 (N_9264,N_2522,N_3618);
and U9265 (N_9265,N_4698,N_2122);
xor U9266 (N_9266,N_2938,N_4145);
nor U9267 (N_9267,N_2650,N_2475);
nand U9268 (N_9268,N_637,N_4238);
nor U9269 (N_9269,N_350,N_2629);
nor U9270 (N_9270,N_4307,N_2552);
nor U9271 (N_9271,N_2483,N_1035);
and U9272 (N_9272,N_4197,N_1330);
and U9273 (N_9273,N_4309,N_1347);
nand U9274 (N_9274,N_2124,N_1737);
or U9275 (N_9275,N_649,N_2770);
nor U9276 (N_9276,N_3512,N_3327);
nand U9277 (N_9277,N_2271,N_584);
nand U9278 (N_9278,N_3510,N_663);
and U9279 (N_9279,N_1869,N_2843);
nor U9280 (N_9280,N_3815,N_3482);
nor U9281 (N_9281,N_233,N_4177);
nand U9282 (N_9282,N_1736,N_1761);
nand U9283 (N_9283,N_3305,N_2196);
or U9284 (N_9284,N_4269,N_28);
nor U9285 (N_9285,N_3667,N_2177);
nor U9286 (N_9286,N_101,N_1292);
nor U9287 (N_9287,N_4541,N_188);
and U9288 (N_9288,N_4133,N_1027);
and U9289 (N_9289,N_1530,N_966);
or U9290 (N_9290,N_4408,N_3819);
and U9291 (N_9291,N_446,N_4523);
or U9292 (N_9292,N_3799,N_2187);
or U9293 (N_9293,N_3923,N_806);
nand U9294 (N_9294,N_432,N_2008);
or U9295 (N_9295,N_4504,N_1779);
xnor U9296 (N_9296,N_3442,N_89);
or U9297 (N_9297,N_3712,N_942);
and U9298 (N_9298,N_3865,N_2);
and U9299 (N_9299,N_1959,N_59);
and U9300 (N_9300,N_3045,N_1245);
nand U9301 (N_9301,N_1704,N_4409);
or U9302 (N_9302,N_2289,N_4735);
nand U9303 (N_9303,N_1598,N_3855);
or U9304 (N_9304,N_3085,N_4099);
nor U9305 (N_9305,N_4429,N_3894);
or U9306 (N_9306,N_3562,N_888);
xor U9307 (N_9307,N_3698,N_2054);
nor U9308 (N_9308,N_4310,N_2927);
and U9309 (N_9309,N_1122,N_1609);
or U9310 (N_9310,N_2274,N_960);
nor U9311 (N_9311,N_2142,N_1899);
or U9312 (N_9312,N_2007,N_1753);
nand U9313 (N_9313,N_4292,N_713);
nor U9314 (N_9314,N_3799,N_1274);
nand U9315 (N_9315,N_2225,N_1662);
or U9316 (N_9316,N_2659,N_88);
nand U9317 (N_9317,N_4647,N_4741);
nand U9318 (N_9318,N_1009,N_3702);
and U9319 (N_9319,N_3477,N_3602);
or U9320 (N_9320,N_4818,N_1438);
and U9321 (N_9321,N_3817,N_2007);
nor U9322 (N_9322,N_2185,N_4523);
or U9323 (N_9323,N_2622,N_4438);
and U9324 (N_9324,N_3581,N_4263);
or U9325 (N_9325,N_2713,N_3054);
or U9326 (N_9326,N_218,N_1522);
or U9327 (N_9327,N_1358,N_585);
nor U9328 (N_9328,N_2211,N_1839);
or U9329 (N_9329,N_2748,N_247);
or U9330 (N_9330,N_3372,N_1399);
and U9331 (N_9331,N_3446,N_3779);
or U9332 (N_9332,N_4908,N_1356);
nor U9333 (N_9333,N_2481,N_3047);
nor U9334 (N_9334,N_4018,N_4986);
and U9335 (N_9335,N_537,N_218);
or U9336 (N_9336,N_3055,N_1753);
nor U9337 (N_9337,N_4921,N_671);
or U9338 (N_9338,N_2960,N_3473);
and U9339 (N_9339,N_4533,N_2352);
or U9340 (N_9340,N_3742,N_1929);
nor U9341 (N_9341,N_2396,N_368);
nand U9342 (N_9342,N_2933,N_4801);
and U9343 (N_9343,N_4251,N_2801);
or U9344 (N_9344,N_4710,N_1637);
or U9345 (N_9345,N_1451,N_4003);
nor U9346 (N_9346,N_2672,N_2479);
and U9347 (N_9347,N_2819,N_4571);
and U9348 (N_9348,N_3623,N_2133);
nor U9349 (N_9349,N_3289,N_1702);
nor U9350 (N_9350,N_16,N_1820);
nand U9351 (N_9351,N_103,N_3810);
nor U9352 (N_9352,N_292,N_2243);
nand U9353 (N_9353,N_3656,N_33);
or U9354 (N_9354,N_3693,N_4009);
nor U9355 (N_9355,N_396,N_1380);
nand U9356 (N_9356,N_806,N_2279);
xnor U9357 (N_9357,N_1870,N_4117);
nand U9358 (N_9358,N_3536,N_2174);
xnor U9359 (N_9359,N_2008,N_2713);
or U9360 (N_9360,N_3211,N_1373);
and U9361 (N_9361,N_4755,N_4517);
nand U9362 (N_9362,N_2868,N_2130);
nand U9363 (N_9363,N_3771,N_1451);
and U9364 (N_9364,N_3026,N_3754);
nand U9365 (N_9365,N_2522,N_4285);
nor U9366 (N_9366,N_2467,N_4727);
nand U9367 (N_9367,N_2095,N_4085);
nand U9368 (N_9368,N_1963,N_288);
xor U9369 (N_9369,N_2617,N_1451);
nor U9370 (N_9370,N_4129,N_3758);
nor U9371 (N_9371,N_2742,N_1395);
or U9372 (N_9372,N_151,N_3407);
and U9373 (N_9373,N_1550,N_4864);
or U9374 (N_9374,N_966,N_4745);
xnor U9375 (N_9375,N_3829,N_1395);
or U9376 (N_9376,N_2678,N_1353);
nand U9377 (N_9377,N_338,N_3761);
nor U9378 (N_9378,N_207,N_3852);
nand U9379 (N_9379,N_4000,N_2249);
nor U9380 (N_9380,N_4295,N_243);
nand U9381 (N_9381,N_4000,N_589);
nand U9382 (N_9382,N_3385,N_4573);
nor U9383 (N_9383,N_2102,N_4345);
xnor U9384 (N_9384,N_4787,N_2450);
nand U9385 (N_9385,N_2281,N_3457);
or U9386 (N_9386,N_701,N_2934);
nor U9387 (N_9387,N_2234,N_1873);
nand U9388 (N_9388,N_2751,N_3850);
or U9389 (N_9389,N_1562,N_3751);
and U9390 (N_9390,N_380,N_262);
or U9391 (N_9391,N_3875,N_4685);
or U9392 (N_9392,N_3846,N_4596);
nor U9393 (N_9393,N_4565,N_1018);
nor U9394 (N_9394,N_1126,N_3989);
nand U9395 (N_9395,N_680,N_4403);
nor U9396 (N_9396,N_4646,N_3781);
nor U9397 (N_9397,N_2308,N_4960);
nor U9398 (N_9398,N_4793,N_1275);
nor U9399 (N_9399,N_4306,N_1616);
nand U9400 (N_9400,N_1821,N_3864);
and U9401 (N_9401,N_259,N_2750);
and U9402 (N_9402,N_3020,N_360);
or U9403 (N_9403,N_4421,N_1545);
or U9404 (N_9404,N_3916,N_1504);
or U9405 (N_9405,N_477,N_4794);
nand U9406 (N_9406,N_4026,N_699);
and U9407 (N_9407,N_1856,N_2078);
and U9408 (N_9408,N_1654,N_4251);
and U9409 (N_9409,N_3321,N_4172);
and U9410 (N_9410,N_1654,N_3670);
or U9411 (N_9411,N_3625,N_967);
nor U9412 (N_9412,N_4356,N_3327);
nand U9413 (N_9413,N_2615,N_1637);
or U9414 (N_9414,N_140,N_1467);
nor U9415 (N_9415,N_271,N_4890);
nand U9416 (N_9416,N_3461,N_3482);
and U9417 (N_9417,N_3036,N_909);
nand U9418 (N_9418,N_4390,N_4705);
nor U9419 (N_9419,N_344,N_3418);
or U9420 (N_9420,N_353,N_1086);
nor U9421 (N_9421,N_715,N_3942);
or U9422 (N_9422,N_4327,N_1943);
nor U9423 (N_9423,N_4871,N_4471);
nor U9424 (N_9424,N_2345,N_61);
nor U9425 (N_9425,N_3091,N_581);
and U9426 (N_9426,N_972,N_92);
nor U9427 (N_9427,N_4584,N_1728);
and U9428 (N_9428,N_4042,N_2260);
nor U9429 (N_9429,N_3085,N_4532);
nor U9430 (N_9430,N_4084,N_4459);
xor U9431 (N_9431,N_2420,N_40);
nor U9432 (N_9432,N_1801,N_2758);
or U9433 (N_9433,N_1437,N_4621);
nor U9434 (N_9434,N_1240,N_2087);
xor U9435 (N_9435,N_1175,N_4485);
nor U9436 (N_9436,N_2218,N_4721);
nand U9437 (N_9437,N_2248,N_1073);
and U9438 (N_9438,N_331,N_4082);
nand U9439 (N_9439,N_4003,N_3194);
xnor U9440 (N_9440,N_3320,N_3787);
or U9441 (N_9441,N_948,N_3951);
nand U9442 (N_9442,N_3645,N_348);
nand U9443 (N_9443,N_4768,N_3465);
and U9444 (N_9444,N_432,N_1987);
nand U9445 (N_9445,N_2759,N_4971);
nor U9446 (N_9446,N_2628,N_2411);
nor U9447 (N_9447,N_3371,N_1549);
nand U9448 (N_9448,N_1294,N_621);
nand U9449 (N_9449,N_4495,N_3425);
xnor U9450 (N_9450,N_658,N_4494);
nor U9451 (N_9451,N_2980,N_1464);
and U9452 (N_9452,N_4034,N_4953);
or U9453 (N_9453,N_2198,N_4936);
nor U9454 (N_9454,N_850,N_4681);
or U9455 (N_9455,N_423,N_2317);
nand U9456 (N_9456,N_1245,N_2247);
nand U9457 (N_9457,N_628,N_3478);
nand U9458 (N_9458,N_1734,N_1325);
nor U9459 (N_9459,N_4976,N_1853);
or U9460 (N_9460,N_1774,N_1671);
or U9461 (N_9461,N_3621,N_1202);
nand U9462 (N_9462,N_4144,N_330);
or U9463 (N_9463,N_1924,N_440);
nor U9464 (N_9464,N_4202,N_1722);
nor U9465 (N_9465,N_4554,N_2378);
or U9466 (N_9466,N_1184,N_4064);
nor U9467 (N_9467,N_3682,N_639);
nor U9468 (N_9468,N_3410,N_1423);
or U9469 (N_9469,N_648,N_4388);
nor U9470 (N_9470,N_2104,N_149);
nand U9471 (N_9471,N_3822,N_2887);
nand U9472 (N_9472,N_1038,N_4516);
and U9473 (N_9473,N_2849,N_4893);
xnor U9474 (N_9474,N_2709,N_4861);
nor U9475 (N_9475,N_2093,N_402);
nand U9476 (N_9476,N_4155,N_1424);
and U9477 (N_9477,N_1514,N_950);
nor U9478 (N_9478,N_2370,N_4122);
and U9479 (N_9479,N_1539,N_1568);
nor U9480 (N_9480,N_1271,N_834);
nor U9481 (N_9481,N_2075,N_2045);
nor U9482 (N_9482,N_4430,N_3548);
nand U9483 (N_9483,N_3493,N_3028);
and U9484 (N_9484,N_3532,N_2930);
nand U9485 (N_9485,N_264,N_2445);
nor U9486 (N_9486,N_2980,N_2380);
nand U9487 (N_9487,N_241,N_695);
nor U9488 (N_9488,N_1597,N_839);
and U9489 (N_9489,N_214,N_1912);
nand U9490 (N_9490,N_2479,N_3781);
and U9491 (N_9491,N_4100,N_4567);
or U9492 (N_9492,N_2265,N_1375);
or U9493 (N_9493,N_4070,N_2463);
or U9494 (N_9494,N_273,N_3344);
nor U9495 (N_9495,N_3275,N_1592);
nand U9496 (N_9496,N_1073,N_1754);
nand U9497 (N_9497,N_740,N_4010);
and U9498 (N_9498,N_676,N_1648);
and U9499 (N_9499,N_2016,N_1970);
and U9500 (N_9500,N_4566,N_4574);
or U9501 (N_9501,N_4576,N_1215);
nor U9502 (N_9502,N_3304,N_1594);
or U9503 (N_9503,N_3432,N_505);
nor U9504 (N_9504,N_642,N_4747);
or U9505 (N_9505,N_4349,N_132);
nand U9506 (N_9506,N_1146,N_4964);
or U9507 (N_9507,N_1868,N_3972);
or U9508 (N_9508,N_1935,N_4215);
nor U9509 (N_9509,N_672,N_3105);
or U9510 (N_9510,N_4155,N_2333);
nor U9511 (N_9511,N_3946,N_3842);
and U9512 (N_9512,N_37,N_430);
nand U9513 (N_9513,N_51,N_4854);
and U9514 (N_9514,N_1165,N_4266);
and U9515 (N_9515,N_481,N_2267);
xnor U9516 (N_9516,N_3905,N_232);
and U9517 (N_9517,N_2849,N_4120);
nor U9518 (N_9518,N_3717,N_4120);
and U9519 (N_9519,N_1646,N_2961);
or U9520 (N_9520,N_3766,N_4199);
nor U9521 (N_9521,N_710,N_2429);
nand U9522 (N_9522,N_1790,N_1895);
or U9523 (N_9523,N_4876,N_68);
nor U9524 (N_9524,N_1043,N_4176);
nand U9525 (N_9525,N_3276,N_4785);
and U9526 (N_9526,N_4526,N_1700);
nand U9527 (N_9527,N_576,N_4586);
nor U9528 (N_9528,N_105,N_4935);
and U9529 (N_9529,N_171,N_2293);
nor U9530 (N_9530,N_2516,N_892);
or U9531 (N_9531,N_1584,N_1627);
or U9532 (N_9532,N_2760,N_3657);
nor U9533 (N_9533,N_4656,N_463);
or U9534 (N_9534,N_1175,N_4155);
nor U9535 (N_9535,N_2947,N_20);
and U9536 (N_9536,N_1291,N_2020);
and U9537 (N_9537,N_3094,N_4162);
or U9538 (N_9538,N_2734,N_163);
or U9539 (N_9539,N_3447,N_1277);
nor U9540 (N_9540,N_519,N_3849);
nor U9541 (N_9541,N_3305,N_1204);
or U9542 (N_9542,N_4427,N_4228);
xor U9543 (N_9543,N_3950,N_4268);
or U9544 (N_9544,N_4638,N_2926);
nor U9545 (N_9545,N_2507,N_3611);
nand U9546 (N_9546,N_1327,N_4790);
or U9547 (N_9547,N_3967,N_3401);
nor U9548 (N_9548,N_2238,N_4264);
and U9549 (N_9549,N_2132,N_2265);
nor U9550 (N_9550,N_1979,N_2781);
nor U9551 (N_9551,N_386,N_4626);
nand U9552 (N_9552,N_337,N_2244);
and U9553 (N_9553,N_862,N_3117);
nand U9554 (N_9554,N_4133,N_3643);
or U9555 (N_9555,N_4320,N_3529);
or U9556 (N_9556,N_2328,N_3619);
or U9557 (N_9557,N_2732,N_3185);
nor U9558 (N_9558,N_1512,N_756);
or U9559 (N_9559,N_2789,N_1921);
nand U9560 (N_9560,N_1258,N_750);
or U9561 (N_9561,N_1063,N_1566);
nand U9562 (N_9562,N_4092,N_327);
nand U9563 (N_9563,N_4770,N_3159);
nand U9564 (N_9564,N_85,N_4675);
or U9565 (N_9565,N_1470,N_1632);
nand U9566 (N_9566,N_2301,N_2689);
nand U9567 (N_9567,N_1132,N_2723);
nor U9568 (N_9568,N_2024,N_695);
and U9569 (N_9569,N_1698,N_2312);
and U9570 (N_9570,N_3930,N_3911);
xnor U9571 (N_9571,N_4487,N_1271);
nand U9572 (N_9572,N_4309,N_963);
nand U9573 (N_9573,N_4426,N_3371);
or U9574 (N_9574,N_4530,N_3568);
nor U9575 (N_9575,N_3962,N_2135);
nor U9576 (N_9576,N_2735,N_3360);
nor U9577 (N_9577,N_1703,N_2925);
or U9578 (N_9578,N_171,N_337);
nand U9579 (N_9579,N_945,N_4127);
and U9580 (N_9580,N_4205,N_2381);
nor U9581 (N_9581,N_4357,N_297);
nor U9582 (N_9582,N_2255,N_2600);
nor U9583 (N_9583,N_755,N_125);
and U9584 (N_9584,N_3513,N_1841);
nand U9585 (N_9585,N_884,N_2688);
or U9586 (N_9586,N_202,N_2885);
nor U9587 (N_9587,N_3451,N_3674);
nor U9588 (N_9588,N_2635,N_67);
and U9589 (N_9589,N_1913,N_4590);
and U9590 (N_9590,N_460,N_619);
and U9591 (N_9591,N_560,N_3479);
xnor U9592 (N_9592,N_1822,N_353);
and U9593 (N_9593,N_3540,N_1669);
nor U9594 (N_9594,N_1401,N_2034);
nand U9595 (N_9595,N_247,N_3630);
nor U9596 (N_9596,N_257,N_3973);
nand U9597 (N_9597,N_3392,N_2745);
or U9598 (N_9598,N_344,N_4010);
or U9599 (N_9599,N_2097,N_1130);
nor U9600 (N_9600,N_1787,N_2642);
and U9601 (N_9601,N_2517,N_1719);
and U9602 (N_9602,N_2687,N_201);
nand U9603 (N_9603,N_1130,N_2557);
nand U9604 (N_9604,N_4822,N_2207);
or U9605 (N_9605,N_1891,N_4913);
or U9606 (N_9606,N_182,N_4993);
nor U9607 (N_9607,N_549,N_4812);
or U9608 (N_9608,N_1380,N_2174);
and U9609 (N_9609,N_4612,N_382);
and U9610 (N_9610,N_3454,N_507);
nand U9611 (N_9611,N_44,N_3597);
nor U9612 (N_9612,N_3441,N_2675);
nor U9613 (N_9613,N_130,N_2307);
and U9614 (N_9614,N_1556,N_1537);
nor U9615 (N_9615,N_2263,N_3364);
or U9616 (N_9616,N_1425,N_1886);
and U9617 (N_9617,N_4611,N_1426);
and U9618 (N_9618,N_2323,N_2084);
nor U9619 (N_9619,N_1696,N_4705);
nand U9620 (N_9620,N_1648,N_447);
nor U9621 (N_9621,N_1881,N_345);
nor U9622 (N_9622,N_337,N_526);
nor U9623 (N_9623,N_534,N_3580);
nand U9624 (N_9624,N_4379,N_3735);
nor U9625 (N_9625,N_1205,N_3349);
or U9626 (N_9626,N_3758,N_203);
or U9627 (N_9627,N_2548,N_3554);
nand U9628 (N_9628,N_3173,N_3956);
and U9629 (N_9629,N_2098,N_3796);
nor U9630 (N_9630,N_223,N_1763);
nor U9631 (N_9631,N_2615,N_1271);
nand U9632 (N_9632,N_1421,N_4933);
and U9633 (N_9633,N_3342,N_2281);
nor U9634 (N_9634,N_144,N_3460);
nand U9635 (N_9635,N_2715,N_3637);
or U9636 (N_9636,N_4805,N_806);
nor U9637 (N_9637,N_1720,N_3165);
and U9638 (N_9638,N_3027,N_72);
nor U9639 (N_9639,N_1587,N_2863);
or U9640 (N_9640,N_135,N_2926);
or U9641 (N_9641,N_2214,N_2749);
or U9642 (N_9642,N_3711,N_2500);
and U9643 (N_9643,N_4932,N_3570);
and U9644 (N_9644,N_70,N_275);
and U9645 (N_9645,N_3492,N_1379);
nand U9646 (N_9646,N_4245,N_1943);
nor U9647 (N_9647,N_123,N_3019);
nand U9648 (N_9648,N_3824,N_217);
nand U9649 (N_9649,N_210,N_2177);
nor U9650 (N_9650,N_3395,N_3055);
and U9651 (N_9651,N_757,N_3197);
or U9652 (N_9652,N_3099,N_3918);
or U9653 (N_9653,N_1352,N_1611);
nand U9654 (N_9654,N_4734,N_870);
or U9655 (N_9655,N_4714,N_727);
nor U9656 (N_9656,N_3020,N_2838);
or U9657 (N_9657,N_1444,N_3193);
and U9658 (N_9658,N_4138,N_1909);
nand U9659 (N_9659,N_4225,N_411);
and U9660 (N_9660,N_3203,N_4123);
and U9661 (N_9661,N_4678,N_1999);
nor U9662 (N_9662,N_3237,N_3928);
nand U9663 (N_9663,N_1692,N_1521);
nor U9664 (N_9664,N_3093,N_3275);
nand U9665 (N_9665,N_828,N_2284);
nor U9666 (N_9666,N_4941,N_4947);
and U9667 (N_9667,N_3398,N_4343);
and U9668 (N_9668,N_1326,N_214);
nand U9669 (N_9669,N_2429,N_88);
nand U9670 (N_9670,N_4949,N_774);
nand U9671 (N_9671,N_3495,N_4003);
and U9672 (N_9672,N_1493,N_684);
nor U9673 (N_9673,N_3852,N_3726);
or U9674 (N_9674,N_1938,N_777);
or U9675 (N_9675,N_1785,N_1392);
nand U9676 (N_9676,N_4707,N_2998);
nand U9677 (N_9677,N_304,N_3549);
or U9678 (N_9678,N_4201,N_185);
or U9679 (N_9679,N_146,N_0);
nand U9680 (N_9680,N_4468,N_3651);
or U9681 (N_9681,N_2262,N_819);
and U9682 (N_9682,N_1320,N_1054);
and U9683 (N_9683,N_1391,N_173);
and U9684 (N_9684,N_4437,N_4302);
nand U9685 (N_9685,N_1363,N_1767);
and U9686 (N_9686,N_65,N_3997);
and U9687 (N_9687,N_2135,N_651);
nand U9688 (N_9688,N_2844,N_3805);
or U9689 (N_9689,N_4759,N_426);
nor U9690 (N_9690,N_1993,N_2995);
and U9691 (N_9691,N_2742,N_4191);
nand U9692 (N_9692,N_117,N_54);
nor U9693 (N_9693,N_3562,N_3481);
and U9694 (N_9694,N_4925,N_4568);
or U9695 (N_9695,N_1082,N_462);
or U9696 (N_9696,N_3377,N_2703);
and U9697 (N_9697,N_877,N_3812);
nor U9698 (N_9698,N_4764,N_2855);
nor U9699 (N_9699,N_1741,N_4833);
or U9700 (N_9700,N_2330,N_2466);
or U9701 (N_9701,N_2960,N_991);
nand U9702 (N_9702,N_2966,N_3783);
nor U9703 (N_9703,N_2355,N_3991);
nand U9704 (N_9704,N_3714,N_805);
or U9705 (N_9705,N_2676,N_1203);
or U9706 (N_9706,N_1418,N_2843);
nor U9707 (N_9707,N_2957,N_1056);
nor U9708 (N_9708,N_3950,N_2115);
nor U9709 (N_9709,N_4812,N_22);
nor U9710 (N_9710,N_4709,N_429);
or U9711 (N_9711,N_3543,N_2188);
nor U9712 (N_9712,N_1733,N_1652);
or U9713 (N_9713,N_3414,N_2592);
and U9714 (N_9714,N_1872,N_3377);
nand U9715 (N_9715,N_1790,N_1777);
and U9716 (N_9716,N_1437,N_627);
nor U9717 (N_9717,N_1,N_3358);
nand U9718 (N_9718,N_3962,N_637);
nand U9719 (N_9719,N_4404,N_2723);
nor U9720 (N_9720,N_3774,N_3993);
nor U9721 (N_9721,N_4775,N_3634);
and U9722 (N_9722,N_4317,N_1505);
nor U9723 (N_9723,N_1159,N_2339);
nor U9724 (N_9724,N_3405,N_3334);
or U9725 (N_9725,N_4688,N_1981);
nor U9726 (N_9726,N_0,N_3349);
nand U9727 (N_9727,N_1899,N_524);
nor U9728 (N_9728,N_2655,N_3395);
nand U9729 (N_9729,N_1606,N_2083);
nor U9730 (N_9730,N_78,N_374);
or U9731 (N_9731,N_4483,N_2533);
nand U9732 (N_9732,N_2408,N_793);
nand U9733 (N_9733,N_4872,N_799);
or U9734 (N_9734,N_4917,N_580);
or U9735 (N_9735,N_4846,N_57);
nor U9736 (N_9736,N_3037,N_1531);
nand U9737 (N_9737,N_3268,N_4357);
or U9738 (N_9738,N_4433,N_3408);
or U9739 (N_9739,N_826,N_3651);
and U9740 (N_9740,N_2908,N_1765);
nand U9741 (N_9741,N_1488,N_989);
or U9742 (N_9742,N_2766,N_879);
nand U9743 (N_9743,N_1967,N_2662);
nor U9744 (N_9744,N_3374,N_3675);
nand U9745 (N_9745,N_1975,N_4562);
or U9746 (N_9746,N_2020,N_1043);
nor U9747 (N_9747,N_3858,N_2951);
and U9748 (N_9748,N_2589,N_2985);
and U9749 (N_9749,N_408,N_4415);
nor U9750 (N_9750,N_3364,N_4101);
or U9751 (N_9751,N_2101,N_4805);
nand U9752 (N_9752,N_4338,N_1116);
or U9753 (N_9753,N_3504,N_3474);
nor U9754 (N_9754,N_862,N_4545);
and U9755 (N_9755,N_2138,N_2161);
nand U9756 (N_9756,N_285,N_2163);
or U9757 (N_9757,N_2564,N_2111);
nand U9758 (N_9758,N_4698,N_3649);
xor U9759 (N_9759,N_3339,N_1769);
or U9760 (N_9760,N_3628,N_4925);
nand U9761 (N_9761,N_2560,N_2175);
or U9762 (N_9762,N_3157,N_4759);
nor U9763 (N_9763,N_477,N_4659);
nand U9764 (N_9764,N_383,N_2613);
nor U9765 (N_9765,N_4206,N_574);
nand U9766 (N_9766,N_4709,N_4369);
or U9767 (N_9767,N_3418,N_1506);
and U9768 (N_9768,N_26,N_2378);
nand U9769 (N_9769,N_3511,N_3532);
or U9770 (N_9770,N_2939,N_4164);
and U9771 (N_9771,N_1214,N_91);
nor U9772 (N_9772,N_1249,N_2023);
and U9773 (N_9773,N_402,N_2732);
nor U9774 (N_9774,N_3051,N_945);
and U9775 (N_9775,N_278,N_924);
and U9776 (N_9776,N_505,N_112);
or U9777 (N_9777,N_4714,N_3094);
and U9778 (N_9778,N_3830,N_3220);
nor U9779 (N_9779,N_2758,N_4474);
nand U9780 (N_9780,N_4716,N_3594);
or U9781 (N_9781,N_2485,N_3836);
or U9782 (N_9782,N_4956,N_1938);
and U9783 (N_9783,N_2862,N_3605);
and U9784 (N_9784,N_2939,N_4423);
or U9785 (N_9785,N_3478,N_3612);
nand U9786 (N_9786,N_4364,N_4111);
and U9787 (N_9787,N_4578,N_4498);
and U9788 (N_9788,N_2850,N_946);
or U9789 (N_9789,N_1269,N_782);
xnor U9790 (N_9790,N_688,N_2667);
and U9791 (N_9791,N_171,N_4345);
xnor U9792 (N_9792,N_1253,N_1265);
or U9793 (N_9793,N_2071,N_1723);
nor U9794 (N_9794,N_1261,N_1103);
or U9795 (N_9795,N_74,N_2033);
nand U9796 (N_9796,N_2432,N_4032);
or U9797 (N_9797,N_3238,N_312);
nand U9798 (N_9798,N_846,N_3526);
nand U9799 (N_9799,N_1480,N_4087);
and U9800 (N_9800,N_4396,N_4126);
xnor U9801 (N_9801,N_3521,N_3770);
or U9802 (N_9802,N_633,N_439);
or U9803 (N_9803,N_3307,N_4257);
nor U9804 (N_9804,N_820,N_2562);
and U9805 (N_9805,N_180,N_1679);
nand U9806 (N_9806,N_3207,N_4706);
nand U9807 (N_9807,N_4572,N_4740);
and U9808 (N_9808,N_1115,N_2201);
and U9809 (N_9809,N_2442,N_3855);
nor U9810 (N_9810,N_1649,N_3510);
and U9811 (N_9811,N_1447,N_306);
and U9812 (N_9812,N_2063,N_2571);
nor U9813 (N_9813,N_2629,N_2677);
or U9814 (N_9814,N_761,N_2903);
nand U9815 (N_9815,N_445,N_3469);
nand U9816 (N_9816,N_4128,N_2299);
nand U9817 (N_9817,N_4265,N_3811);
and U9818 (N_9818,N_2202,N_3054);
nor U9819 (N_9819,N_1536,N_664);
or U9820 (N_9820,N_566,N_4568);
and U9821 (N_9821,N_791,N_2291);
nand U9822 (N_9822,N_4290,N_565);
nor U9823 (N_9823,N_3545,N_4387);
nor U9824 (N_9824,N_2061,N_906);
and U9825 (N_9825,N_1218,N_2793);
xnor U9826 (N_9826,N_2122,N_1444);
nand U9827 (N_9827,N_306,N_2652);
or U9828 (N_9828,N_3342,N_4147);
and U9829 (N_9829,N_2745,N_3074);
or U9830 (N_9830,N_3778,N_4914);
and U9831 (N_9831,N_462,N_343);
and U9832 (N_9832,N_2824,N_4632);
and U9833 (N_9833,N_2619,N_4699);
nor U9834 (N_9834,N_1708,N_2901);
or U9835 (N_9835,N_3659,N_3498);
nand U9836 (N_9836,N_1782,N_3516);
nand U9837 (N_9837,N_1677,N_2222);
and U9838 (N_9838,N_3829,N_4005);
nor U9839 (N_9839,N_103,N_2766);
and U9840 (N_9840,N_3591,N_382);
and U9841 (N_9841,N_3096,N_20);
and U9842 (N_9842,N_3948,N_2464);
and U9843 (N_9843,N_2883,N_773);
and U9844 (N_9844,N_4149,N_1624);
and U9845 (N_9845,N_1926,N_1890);
nor U9846 (N_9846,N_2480,N_798);
nor U9847 (N_9847,N_1288,N_2156);
and U9848 (N_9848,N_2034,N_1388);
nand U9849 (N_9849,N_4649,N_2866);
nor U9850 (N_9850,N_4241,N_2406);
or U9851 (N_9851,N_178,N_1925);
nor U9852 (N_9852,N_3834,N_2663);
nor U9853 (N_9853,N_2209,N_103);
or U9854 (N_9854,N_4695,N_404);
and U9855 (N_9855,N_3699,N_704);
nand U9856 (N_9856,N_4897,N_3832);
nor U9857 (N_9857,N_2956,N_2396);
nor U9858 (N_9858,N_379,N_2977);
or U9859 (N_9859,N_1470,N_4773);
nand U9860 (N_9860,N_1667,N_1931);
or U9861 (N_9861,N_640,N_4260);
nor U9862 (N_9862,N_967,N_530);
nand U9863 (N_9863,N_4011,N_1342);
and U9864 (N_9864,N_899,N_2919);
and U9865 (N_9865,N_2055,N_3657);
and U9866 (N_9866,N_3960,N_4005);
or U9867 (N_9867,N_2390,N_4436);
or U9868 (N_9868,N_1467,N_2991);
and U9869 (N_9869,N_575,N_4678);
nor U9870 (N_9870,N_4475,N_1952);
xnor U9871 (N_9871,N_2572,N_92);
or U9872 (N_9872,N_2305,N_586);
and U9873 (N_9873,N_2837,N_637);
nor U9874 (N_9874,N_3956,N_2492);
nor U9875 (N_9875,N_1700,N_1503);
nand U9876 (N_9876,N_4362,N_1128);
nor U9877 (N_9877,N_532,N_4536);
nor U9878 (N_9878,N_1431,N_4755);
and U9879 (N_9879,N_4892,N_1684);
nand U9880 (N_9880,N_2575,N_997);
and U9881 (N_9881,N_4132,N_709);
nand U9882 (N_9882,N_4152,N_1836);
nor U9883 (N_9883,N_2982,N_4608);
nand U9884 (N_9884,N_4154,N_1669);
nor U9885 (N_9885,N_3028,N_1891);
and U9886 (N_9886,N_2665,N_2083);
and U9887 (N_9887,N_4188,N_4818);
and U9888 (N_9888,N_1045,N_4811);
or U9889 (N_9889,N_4632,N_2276);
nand U9890 (N_9890,N_3438,N_4162);
or U9891 (N_9891,N_1637,N_2738);
nor U9892 (N_9892,N_4621,N_2484);
and U9893 (N_9893,N_2803,N_2574);
nand U9894 (N_9894,N_1605,N_3900);
nand U9895 (N_9895,N_3921,N_2545);
nor U9896 (N_9896,N_4392,N_4261);
nor U9897 (N_9897,N_1750,N_4826);
and U9898 (N_9898,N_2525,N_1611);
and U9899 (N_9899,N_2469,N_2626);
nor U9900 (N_9900,N_2825,N_3635);
nor U9901 (N_9901,N_4926,N_4156);
and U9902 (N_9902,N_2571,N_2031);
or U9903 (N_9903,N_3851,N_595);
nor U9904 (N_9904,N_2672,N_1571);
nor U9905 (N_9905,N_719,N_537);
nand U9906 (N_9906,N_3321,N_3764);
or U9907 (N_9907,N_660,N_1213);
nand U9908 (N_9908,N_2455,N_380);
nand U9909 (N_9909,N_929,N_1034);
or U9910 (N_9910,N_1088,N_1379);
and U9911 (N_9911,N_3918,N_1506);
nor U9912 (N_9912,N_2515,N_2998);
nor U9913 (N_9913,N_1262,N_3500);
nand U9914 (N_9914,N_2256,N_3278);
or U9915 (N_9915,N_753,N_1406);
and U9916 (N_9916,N_126,N_2961);
nor U9917 (N_9917,N_893,N_1702);
and U9918 (N_9918,N_426,N_4726);
or U9919 (N_9919,N_982,N_2400);
or U9920 (N_9920,N_4157,N_2431);
nand U9921 (N_9921,N_666,N_4070);
nand U9922 (N_9922,N_2936,N_147);
or U9923 (N_9923,N_261,N_1200);
xnor U9924 (N_9924,N_4115,N_2199);
nor U9925 (N_9925,N_495,N_603);
and U9926 (N_9926,N_1603,N_2193);
nand U9927 (N_9927,N_3008,N_1393);
nand U9928 (N_9928,N_473,N_918);
or U9929 (N_9929,N_2026,N_3885);
xnor U9930 (N_9930,N_4639,N_1680);
or U9931 (N_9931,N_869,N_1364);
nand U9932 (N_9932,N_691,N_4091);
and U9933 (N_9933,N_2572,N_4311);
nand U9934 (N_9934,N_4139,N_3676);
nand U9935 (N_9935,N_2109,N_3337);
nor U9936 (N_9936,N_1068,N_3569);
or U9937 (N_9937,N_1109,N_4370);
nor U9938 (N_9938,N_2184,N_3962);
nor U9939 (N_9939,N_4647,N_2289);
nor U9940 (N_9940,N_3877,N_1684);
nor U9941 (N_9941,N_1235,N_3612);
nand U9942 (N_9942,N_1177,N_2469);
xnor U9943 (N_9943,N_1260,N_4681);
nand U9944 (N_9944,N_504,N_4533);
nand U9945 (N_9945,N_2125,N_1278);
and U9946 (N_9946,N_2275,N_296);
nand U9947 (N_9947,N_12,N_2440);
xnor U9948 (N_9948,N_19,N_2677);
or U9949 (N_9949,N_3426,N_2199);
nor U9950 (N_9950,N_1729,N_4521);
and U9951 (N_9951,N_3897,N_4410);
or U9952 (N_9952,N_1723,N_890);
nand U9953 (N_9953,N_1651,N_802);
or U9954 (N_9954,N_1983,N_2788);
xor U9955 (N_9955,N_1433,N_1079);
nor U9956 (N_9956,N_1082,N_208);
nand U9957 (N_9957,N_986,N_4567);
nand U9958 (N_9958,N_2708,N_1246);
or U9959 (N_9959,N_4188,N_1796);
or U9960 (N_9960,N_4269,N_47);
or U9961 (N_9961,N_3551,N_307);
xnor U9962 (N_9962,N_4926,N_3362);
nand U9963 (N_9963,N_1796,N_3540);
nor U9964 (N_9964,N_4994,N_4598);
or U9965 (N_9965,N_1801,N_4359);
nor U9966 (N_9966,N_4936,N_1138);
nand U9967 (N_9967,N_2922,N_3821);
nand U9968 (N_9968,N_2506,N_2941);
and U9969 (N_9969,N_3652,N_4959);
nor U9970 (N_9970,N_591,N_1522);
nor U9971 (N_9971,N_1248,N_2424);
or U9972 (N_9972,N_4582,N_2369);
nand U9973 (N_9973,N_3099,N_4099);
or U9974 (N_9974,N_1207,N_2350);
and U9975 (N_9975,N_626,N_1877);
nor U9976 (N_9976,N_2123,N_4877);
or U9977 (N_9977,N_1854,N_1945);
and U9978 (N_9978,N_3903,N_4099);
or U9979 (N_9979,N_4322,N_1542);
nand U9980 (N_9980,N_1985,N_3831);
nor U9981 (N_9981,N_821,N_1775);
and U9982 (N_9982,N_3782,N_645);
nand U9983 (N_9983,N_25,N_3744);
and U9984 (N_9984,N_2736,N_4785);
or U9985 (N_9985,N_4672,N_4095);
nor U9986 (N_9986,N_1214,N_1036);
nand U9987 (N_9987,N_4865,N_2505);
and U9988 (N_9988,N_1893,N_1587);
nand U9989 (N_9989,N_2527,N_720);
and U9990 (N_9990,N_3517,N_4557);
or U9991 (N_9991,N_309,N_3376);
and U9992 (N_9992,N_2373,N_3626);
and U9993 (N_9993,N_4776,N_1136);
nand U9994 (N_9994,N_2461,N_246);
or U9995 (N_9995,N_1634,N_3127);
nor U9996 (N_9996,N_3505,N_846);
and U9997 (N_9997,N_4785,N_3288);
nand U9998 (N_9998,N_4952,N_2661);
or U9999 (N_9999,N_2793,N_1150);
nor U10000 (N_10000,N_6336,N_6186);
nor U10001 (N_10001,N_5463,N_8265);
or U10002 (N_10002,N_6922,N_6899);
nor U10003 (N_10003,N_8157,N_7249);
and U10004 (N_10004,N_9719,N_6198);
nand U10005 (N_10005,N_5424,N_8503);
or U10006 (N_10006,N_6891,N_8842);
nand U10007 (N_10007,N_5117,N_9785);
or U10008 (N_10008,N_5817,N_6791);
nand U10009 (N_10009,N_6923,N_6565);
and U10010 (N_10010,N_9569,N_6196);
and U10011 (N_10011,N_6815,N_8695);
nand U10012 (N_10012,N_9938,N_6517);
and U10013 (N_10013,N_7040,N_6754);
or U10014 (N_10014,N_7625,N_6768);
and U10015 (N_10015,N_8287,N_5605);
and U10016 (N_10016,N_6299,N_5308);
nand U10017 (N_10017,N_6540,N_6395);
nor U10018 (N_10018,N_8596,N_9154);
and U10019 (N_10019,N_8903,N_8873);
and U10020 (N_10020,N_8659,N_7620);
nor U10021 (N_10021,N_6093,N_6499);
and U10022 (N_10022,N_8914,N_9839);
nand U10023 (N_10023,N_8551,N_9511);
or U10024 (N_10024,N_7994,N_8658);
nand U10025 (N_10025,N_9304,N_7489);
or U10026 (N_10026,N_8429,N_5039);
nand U10027 (N_10027,N_7838,N_8812);
and U10028 (N_10028,N_6383,N_6624);
nand U10029 (N_10029,N_7582,N_6012);
xnor U10030 (N_10030,N_8107,N_6570);
nand U10031 (N_10031,N_5724,N_5874);
nor U10032 (N_10032,N_7631,N_6504);
nand U10033 (N_10033,N_7375,N_6458);
and U10034 (N_10034,N_6285,N_7825);
nor U10035 (N_10035,N_6035,N_7422);
or U10036 (N_10036,N_7647,N_8644);
and U10037 (N_10037,N_8719,N_5581);
or U10038 (N_10038,N_7330,N_9484);
or U10039 (N_10039,N_8898,N_6621);
nor U10040 (N_10040,N_7370,N_9611);
or U10041 (N_10041,N_8385,N_6507);
nor U10042 (N_10042,N_7666,N_5657);
xnor U10043 (N_10043,N_8228,N_8422);
nand U10044 (N_10044,N_8282,N_6536);
nor U10045 (N_10045,N_5468,N_7954);
or U10046 (N_10046,N_8307,N_9789);
nand U10047 (N_10047,N_9931,N_7563);
nand U10048 (N_10048,N_8068,N_9197);
nor U10049 (N_10049,N_5661,N_9090);
nor U10050 (N_10050,N_9541,N_5523);
and U10051 (N_10051,N_7983,N_8383);
or U10052 (N_10052,N_9928,N_9645);
nor U10053 (N_10053,N_8703,N_6138);
nand U10054 (N_10054,N_8017,N_7070);
or U10055 (N_10055,N_7674,N_9794);
or U10056 (N_10056,N_6874,N_8798);
and U10057 (N_10057,N_9512,N_9991);
nor U10058 (N_10058,N_9152,N_6075);
or U10059 (N_10059,N_7492,N_9057);
nand U10060 (N_10060,N_8876,N_7786);
or U10061 (N_10061,N_9217,N_8723);
or U10062 (N_10062,N_9535,N_9588);
and U10063 (N_10063,N_7267,N_5006);
nand U10064 (N_10064,N_9817,N_5638);
or U10065 (N_10065,N_5337,N_5350);
nand U10066 (N_10066,N_6257,N_6433);
and U10067 (N_10067,N_8086,N_9486);
and U10068 (N_10068,N_5572,N_6231);
nor U10069 (N_10069,N_8253,N_5241);
or U10070 (N_10070,N_5669,N_7176);
or U10071 (N_10071,N_6320,N_8366);
nand U10072 (N_10072,N_5474,N_7741);
or U10073 (N_10073,N_5680,N_7182);
and U10074 (N_10074,N_5883,N_7399);
nor U10075 (N_10075,N_8747,N_8145);
nand U10076 (N_10076,N_5044,N_5094);
and U10077 (N_10077,N_5888,N_5491);
or U10078 (N_10078,N_7455,N_8928);
or U10079 (N_10079,N_6465,N_8742);
nor U10080 (N_10080,N_7235,N_6003);
or U10081 (N_10081,N_8572,N_9821);
xnor U10082 (N_10082,N_9503,N_9670);
and U10083 (N_10083,N_5076,N_8337);
or U10084 (N_10084,N_6038,N_5989);
xor U10085 (N_10085,N_5443,N_5569);
nor U10086 (N_10086,N_9426,N_6496);
and U10087 (N_10087,N_8395,N_9352);
nand U10088 (N_10088,N_6040,N_5891);
nand U10089 (N_10089,N_6237,N_6324);
and U10090 (N_10090,N_9501,N_8089);
and U10091 (N_10091,N_6284,N_9324);
or U10092 (N_10092,N_9578,N_5882);
nand U10093 (N_10093,N_8188,N_6466);
and U10094 (N_10094,N_6575,N_7774);
nor U10095 (N_10095,N_5890,N_6961);
nand U10096 (N_10096,N_9592,N_5852);
or U10097 (N_10097,N_6409,N_7606);
or U10098 (N_10098,N_9721,N_7279);
and U10099 (N_10099,N_6041,N_5287);
xor U10100 (N_10100,N_9864,N_5920);
nand U10101 (N_10101,N_8257,N_6426);
or U10102 (N_10102,N_7989,N_7123);
or U10103 (N_10103,N_9508,N_8532);
and U10104 (N_10104,N_9002,N_7949);
nand U10105 (N_10105,N_5597,N_9590);
nor U10106 (N_10106,N_8755,N_9895);
nor U10107 (N_10107,N_8748,N_8909);
nor U10108 (N_10108,N_6640,N_8983);
nand U10109 (N_10109,N_5823,N_6490);
nand U10110 (N_10110,N_7209,N_6293);
and U10111 (N_10111,N_8308,N_9335);
and U10112 (N_10112,N_9440,N_6715);
nor U10113 (N_10113,N_6559,N_8635);
and U10114 (N_10114,N_6226,N_5728);
and U10115 (N_10115,N_7591,N_6014);
and U10116 (N_10116,N_8538,N_9058);
nand U10117 (N_10117,N_5098,N_8530);
xor U10118 (N_10118,N_5751,N_5123);
nand U10119 (N_10119,N_9212,N_5666);
nand U10120 (N_10120,N_7392,N_8499);
or U10121 (N_10121,N_6069,N_8069);
and U10122 (N_10122,N_6248,N_5650);
and U10123 (N_10123,N_9402,N_8312);
nor U10124 (N_10124,N_6886,N_6488);
and U10125 (N_10125,N_7614,N_6236);
nor U10126 (N_10126,N_7711,N_8076);
nand U10127 (N_10127,N_9014,N_6592);
nand U10128 (N_10128,N_7733,N_8850);
nand U10129 (N_10129,N_8116,N_5630);
or U10130 (N_10130,N_6515,N_6403);
nor U10131 (N_10131,N_8210,N_5100);
and U10132 (N_10132,N_6586,N_9061);
xor U10133 (N_10133,N_5551,N_6937);
nand U10134 (N_10134,N_7951,N_9963);
and U10135 (N_10135,N_5283,N_9136);
or U10136 (N_10136,N_8881,N_8485);
nand U10137 (N_10137,N_5476,N_6491);
and U10138 (N_10138,N_7452,N_8232);
or U10139 (N_10139,N_7406,N_9914);
nand U10140 (N_10140,N_7996,N_9149);
nand U10141 (N_10141,N_8113,N_8930);
nor U10142 (N_10142,N_6483,N_9393);
nand U10143 (N_10143,N_8368,N_6200);
nor U10144 (N_10144,N_7887,N_5451);
or U10145 (N_10145,N_9722,N_9881);
xor U10146 (N_10146,N_8487,N_5719);
nor U10147 (N_10147,N_6717,N_7790);
nand U10148 (N_10148,N_9325,N_6881);
nor U10149 (N_10149,N_9060,N_5806);
and U10150 (N_10150,N_7942,N_8163);
or U10151 (N_10151,N_7408,N_7086);
and U10152 (N_10152,N_8494,N_8313);
nor U10153 (N_10153,N_7108,N_8333);
nand U10154 (N_10154,N_9676,N_5472);
or U10155 (N_10155,N_8700,N_6702);
nor U10156 (N_10156,N_9565,N_8373);
nor U10157 (N_10157,N_8408,N_8629);
nand U10158 (N_10158,N_7776,N_6927);
nand U10159 (N_10159,N_7331,N_7924);
and U10160 (N_10160,N_8518,N_8254);
and U10161 (N_10161,N_9348,N_9827);
nor U10162 (N_10162,N_6533,N_7119);
nand U10163 (N_10163,N_6027,N_7019);
or U10164 (N_10164,N_5255,N_7819);
nor U10165 (N_10165,N_6314,N_5278);
and U10166 (N_10166,N_6178,N_6520);
nor U10167 (N_10167,N_9870,N_6387);
nor U10168 (N_10168,N_5770,N_9954);
nand U10169 (N_10169,N_5462,N_8998);
nand U10170 (N_10170,N_6745,N_5968);
nand U10171 (N_10171,N_6984,N_8270);
nand U10172 (N_10172,N_5950,N_8979);
nand U10173 (N_10173,N_8272,N_8018);
or U10174 (N_10174,N_9619,N_6099);
nand U10175 (N_10175,N_9280,N_8022);
nor U10176 (N_10176,N_9081,N_7170);
and U10177 (N_10177,N_9457,N_7564);
and U10178 (N_10178,N_5836,N_9295);
or U10179 (N_10179,N_9820,N_8424);
or U10180 (N_10180,N_7476,N_6065);
or U10181 (N_10181,N_9837,N_7839);
nor U10182 (N_10182,N_9939,N_7241);
and U10183 (N_10183,N_9552,N_7527);
and U10184 (N_10184,N_8728,N_6130);
and U10185 (N_10185,N_8939,N_7121);
nor U10186 (N_10186,N_6896,N_8191);
or U10187 (N_10187,N_8513,N_8516);
or U10188 (N_10188,N_5172,N_8033);
nor U10189 (N_10189,N_8846,N_5060);
nand U10190 (N_10190,N_8824,N_9990);
nand U10191 (N_10191,N_5247,N_7254);
nand U10192 (N_10192,N_8460,N_5933);
or U10193 (N_10193,N_5401,N_6825);
nor U10194 (N_10194,N_9211,N_6351);
nand U10195 (N_10195,N_5786,N_9246);
xnor U10196 (N_10196,N_8932,N_7589);
or U10197 (N_10197,N_7622,N_8609);
and U10198 (N_10198,N_8220,N_8016);
nand U10199 (N_10199,N_9048,N_5640);
nand U10200 (N_10200,N_5570,N_5326);
nand U10201 (N_10201,N_5783,N_5410);
nor U10202 (N_10202,N_5613,N_6642);
and U10203 (N_10203,N_7288,N_8687);
xor U10204 (N_10204,N_5186,N_7366);
nand U10205 (N_10205,N_5936,N_5233);
nand U10206 (N_10206,N_8814,N_7383);
nand U10207 (N_10207,N_5899,N_5919);
nand U10208 (N_10208,N_6386,N_6577);
or U10209 (N_10209,N_6061,N_7042);
or U10210 (N_10210,N_5096,N_6232);
or U10211 (N_10211,N_5743,N_9549);
nor U10212 (N_10212,N_7217,N_8866);
nor U10213 (N_10213,N_6921,N_5479);
or U10214 (N_10214,N_5150,N_8779);
and U10215 (N_10215,N_7233,N_5854);
nand U10216 (N_10216,N_9546,N_6235);
and U10217 (N_10217,N_8568,N_5790);
nor U10218 (N_10218,N_9986,N_8843);
or U10219 (N_10219,N_7002,N_8761);
nor U10220 (N_10220,N_8660,N_6736);
and U10221 (N_10221,N_7546,N_5805);
or U10222 (N_10222,N_9347,N_9650);
and U10223 (N_10223,N_7828,N_6853);
and U10224 (N_10224,N_8238,N_7512);
nand U10225 (N_10225,N_6808,N_6141);
or U10226 (N_10226,N_6271,N_7526);
nor U10227 (N_10227,N_6511,N_8054);
or U10228 (N_10228,N_6229,N_9069);
nand U10229 (N_10229,N_9840,N_6510);
and U10230 (N_10230,N_9139,N_8330);
nand U10231 (N_10231,N_7867,N_8533);
nor U10232 (N_10232,N_8486,N_8725);
xnor U10233 (N_10233,N_7573,N_8562);
nor U10234 (N_10234,N_8038,N_7590);
or U10235 (N_10235,N_6078,N_8957);
nor U10236 (N_10236,N_8520,N_7269);
nand U10237 (N_10237,N_6480,N_6476);
or U10238 (N_10238,N_5845,N_5927);
nand U10239 (N_10239,N_9823,N_5238);
and U10240 (N_10240,N_6008,N_8663);
xnor U10241 (N_10241,N_6744,N_8524);
and U10242 (N_10242,N_8787,N_9661);
or U10243 (N_10243,N_8692,N_8620);
nand U10244 (N_10244,N_8139,N_9685);
nand U10245 (N_10245,N_6560,N_9213);
or U10246 (N_10246,N_5069,N_6345);
or U10247 (N_10247,N_5258,N_8565);
or U10248 (N_10248,N_6557,N_7579);
nor U10249 (N_10249,N_7192,N_8441);
nor U10250 (N_10250,N_8137,N_9129);
and U10251 (N_10251,N_9648,N_5007);
nand U10252 (N_10252,N_5125,N_5261);
nor U10253 (N_10253,N_7545,N_9167);
or U10254 (N_10254,N_7745,N_7431);
nand U10255 (N_10255,N_9236,N_7343);
and U10256 (N_10256,N_5140,N_6968);
nor U10257 (N_10257,N_6847,N_6672);
or U10258 (N_10258,N_8488,N_8143);
nand U10259 (N_10259,N_6122,N_7735);
and U10260 (N_10260,N_9615,N_8858);
and U10261 (N_10261,N_6902,N_6172);
nor U10262 (N_10262,N_7253,N_5524);
and U10263 (N_10263,N_5008,N_8744);
nand U10264 (N_10264,N_9413,N_9887);
nand U10265 (N_10265,N_6408,N_7872);
nand U10266 (N_10266,N_6372,N_9239);
nor U10267 (N_10267,N_9193,N_6930);
and U10268 (N_10268,N_5810,N_7138);
nor U10269 (N_10269,N_5302,N_8431);
or U10270 (N_10270,N_9625,N_9664);
nor U10271 (N_10271,N_8216,N_8926);
or U10272 (N_10272,N_5345,N_9117);
or U10273 (N_10273,N_5309,N_6770);
nand U10274 (N_10274,N_8132,N_8314);
xnor U10275 (N_10275,N_5733,N_7039);
and U10276 (N_10276,N_6564,N_6622);
nand U10277 (N_10277,N_6107,N_8675);
nor U10278 (N_10278,N_9669,N_7827);
nand U10279 (N_10279,N_5469,N_7948);
xor U10280 (N_10280,N_8970,N_7821);
and U10281 (N_10281,N_7189,N_5525);
or U10282 (N_10282,N_9783,N_9714);
xnor U10283 (N_10283,N_7200,N_5483);
and U10284 (N_10284,N_6890,N_7760);
and U10285 (N_10285,N_7922,N_7319);
or U10286 (N_10286,N_6331,N_6188);
and U10287 (N_10287,N_9258,N_6174);
nand U10288 (N_10288,N_6365,N_5589);
nor U10289 (N_10289,N_7421,N_9039);
or U10290 (N_10290,N_8340,N_5692);
nand U10291 (N_10291,N_5796,N_6713);
or U10292 (N_10292,N_5236,N_6080);
or U10293 (N_10293,N_7682,N_8212);
nand U10294 (N_10294,N_6435,N_7901);
and U10295 (N_10295,N_6227,N_8569);
nor U10296 (N_10296,N_5380,N_8955);
nand U10297 (N_10297,N_9355,N_6149);
or U10298 (N_10298,N_9753,N_7340);
and U10299 (N_10299,N_7958,N_7640);
nand U10300 (N_10300,N_8831,N_6379);
nand U10301 (N_10301,N_8067,N_9893);
nand U10302 (N_10302,N_8450,N_9663);
nor U10303 (N_10303,N_6725,N_7505);
nand U10304 (N_10304,N_6263,N_6469);
nand U10305 (N_10305,N_7877,N_9107);
and U10306 (N_10306,N_8229,N_6849);
xnor U10307 (N_10307,N_6940,N_7858);
or U10308 (N_10308,N_8258,N_7078);
and U10309 (N_10309,N_6260,N_5161);
xnor U10310 (N_10310,N_8878,N_5934);
nor U10311 (N_10311,N_8531,N_5406);
and U10312 (N_10312,N_7762,N_6604);
and U10313 (N_10313,N_7220,N_7141);
or U10314 (N_10314,N_9718,N_7824);
or U10315 (N_10315,N_5187,N_9679);
nor U10316 (N_10316,N_6451,N_5695);
nand U10317 (N_10317,N_5598,N_7933);
or U10318 (N_10318,N_9302,N_7696);
or U10319 (N_10319,N_7891,N_9805);
and U10320 (N_10320,N_7679,N_5629);
and U10321 (N_10321,N_6848,N_8585);
nor U10322 (N_10322,N_9003,N_7416);
or U10323 (N_10323,N_5996,N_9769);
and U10324 (N_10324,N_7178,N_9027);
nor U10325 (N_10325,N_7283,N_5225);
xnor U10326 (N_10326,N_7243,N_6820);
nor U10327 (N_10327,N_5079,N_9759);
or U10328 (N_10328,N_9475,N_9183);
or U10329 (N_10329,N_5508,N_6784);
nand U10330 (N_10330,N_7829,N_9277);
nor U10331 (N_10331,N_8147,N_6004);
nor U10332 (N_10332,N_6007,N_8050);
nor U10333 (N_10333,N_7908,N_9320);
nor U10334 (N_10334,N_5071,N_9981);
or U10335 (N_10335,N_8203,N_9967);
nand U10336 (N_10336,N_6840,N_6211);
and U10337 (N_10337,N_6264,N_7676);
and U10338 (N_10338,N_6751,N_9017);
nor U10339 (N_10339,N_6571,N_8950);
nand U10340 (N_10340,N_8390,N_7481);
nor U10341 (N_10341,N_8377,N_7895);
nand U10342 (N_10342,N_6824,N_9219);
nor U10343 (N_10343,N_5653,N_8321);
nand U10344 (N_10344,N_5073,N_9741);
or U10345 (N_10345,N_5470,N_6316);
nor U10346 (N_10346,N_6357,N_6760);
nor U10347 (N_10347,N_7362,N_8708);
or U10348 (N_10348,N_6100,N_8665);
nand U10349 (N_10349,N_9897,N_9309);
and U10350 (N_10350,N_9647,N_5399);
and U10351 (N_10351,N_6812,N_8536);
nand U10352 (N_10352,N_8154,N_8769);
or U10353 (N_10353,N_6204,N_9111);
and U10354 (N_10354,N_9982,N_8380);
or U10355 (N_10355,N_9106,N_8410);
nand U10356 (N_10356,N_8246,N_7557);
and U10357 (N_10357,N_7990,N_6615);
and U10358 (N_10358,N_7627,N_9198);
or U10359 (N_10359,N_6865,N_9382);
or U10360 (N_10360,N_7446,N_7817);
and U10361 (N_10361,N_8036,N_8465);
and U10362 (N_10362,N_5562,N_7894);
nor U10363 (N_10363,N_6841,N_6827);
or U10364 (N_10364,N_5361,N_5317);
nor U10365 (N_10365,N_8766,N_7087);
nor U10366 (N_10366,N_9196,N_5700);
or U10367 (N_10367,N_7597,N_5142);
nor U10368 (N_10368,N_9192,N_9510);
nand U10369 (N_10369,N_8586,N_6405);
and U10370 (N_10370,N_6844,N_9879);
and U10371 (N_10371,N_5591,N_8962);
and U10372 (N_10372,N_5394,N_9849);
nor U10373 (N_10373,N_5029,N_8347);
nor U10374 (N_10374,N_8927,N_5028);
or U10375 (N_10375,N_6215,N_9008);
and U10376 (N_10376,N_9960,N_5844);
and U10377 (N_10377,N_7521,N_5343);
xor U10378 (N_10378,N_6421,N_7734);
nor U10379 (N_10379,N_5592,N_8498);
and U10380 (N_10380,N_6101,N_6822);
nor U10381 (N_10381,N_7599,N_7208);
or U10382 (N_10382,N_7298,N_8591);
nand U10383 (N_10383,N_7934,N_7617);
or U10384 (N_10384,N_5516,N_9843);
xor U10385 (N_10385,N_9845,N_5557);
and U10386 (N_10386,N_8561,N_7360);
and U10387 (N_10387,N_8063,N_7124);
nor U10388 (N_10388,N_8448,N_5718);
nand U10389 (N_10389,N_7544,N_6990);
xor U10390 (N_10390,N_7664,N_5875);
and U10391 (N_10391,N_7285,N_9743);
nor U10392 (N_10392,N_7270,N_8495);
or U10393 (N_10393,N_9161,N_8432);
and U10394 (N_10394,N_6733,N_5769);
and U10395 (N_10395,N_6866,N_9121);
nand U10396 (N_10396,N_6005,N_7761);
nor U10397 (N_10397,N_6430,N_8696);
or U10398 (N_10398,N_8793,N_7228);
and U10399 (N_10399,N_9886,N_9370);
nor U10400 (N_10400,N_8535,N_9405);
and U10401 (N_10401,N_9707,N_5437);
nor U10402 (N_10402,N_9563,N_8521);
nand U10403 (N_10403,N_5487,N_5878);
nand U10404 (N_10404,N_6893,N_9976);
or U10405 (N_10405,N_5202,N_8359);
or U10406 (N_10406,N_6350,N_7265);
and U10407 (N_10407,N_8605,N_6718);
nor U10408 (N_10408,N_6197,N_7034);
nand U10409 (N_10409,N_6845,N_7671);
xor U10410 (N_10410,N_5987,N_6422);
and U10411 (N_10411,N_5766,N_6762);
and U10412 (N_10412,N_5847,N_5730);
or U10413 (N_10413,N_8716,N_5024);
and U10414 (N_10414,N_5281,N_6388);
nor U10415 (N_10415,N_8899,N_7278);
or U10416 (N_10416,N_7518,N_6796);
and U10417 (N_10417,N_8006,N_5535);
and U10418 (N_10418,N_5010,N_7258);
or U10419 (N_10419,N_6210,N_9168);
nor U10420 (N_10420,N_5279,N_7353);
or U10421 (N_10421,N_8339,N_6449);
or U10422 (N_10422,N_9275,N_8049);
nand U10423 (N_10423,N_8717,N_6296);
or U10424 (N_10424,N_8686,N_7099);
or U10425 (N_10425,N_8820,N_5955);
nand U10426 (N_10426,N_5252,N_9350);
nand U10427 (N_10427,N_5618,N_7498);
and U10428 (N_10428,N_6993,N_5811);
or U10429 (N_10429,N_6885,N_7067);
nand U10430 (N_10430,N_9918,N_9969);
nand U10431 (N_10431,N_8973,N_5993);
nand U10432 (N_10432,N_5715,N_5198);
nor U10433 (N_10433,N_7104,N_6797);
nand U10434 (N_10434,N_6667,N_5671);
and U10435 (N_10435,N_8822,N_5460);
nand U10436 (N_10436,N_5344,N_6190);
nand U10437 (N_10437,N_5015,N_5956);
or U10438 (N_10438,N_5921,N_8630);
nor U10439 (N_10439,N_5851,N_5564);
or U10440 (N_10440,N_9697,N_6487);
nand U10441 (N_10441,N_6221,N_8466);
and U10442 (N_10442,N_6156,N_7312);
nor U10443 (N_10443,N_7947,N_7484);
or U10444 (N_10444,N_5262,N_7571);
or U10445 (N_10445,N_8219,N_5881);
or U10446 (N_10446,N_5215,N_7555);
nand U10447 (N_10447,N_6276,N_6908);
and U10448 (N_10448,N_9851,N_6707);
or U10449 (N_10449,N_8438,N_8056);
and U10450 (N_10450,N_6817,N_8773);
and U10451 (N_10451,N_6482,N_8632);
nor U10452 (N_10452,N_7763,N_7804);
nor U10453 (N_10453,N_5149,N_6121);
nor U10454 (N_10454,N_8776,N_7356);
or U10455 (N_10455,N_5420,N_5121);
or U10456 (N_10456,N_8934,N_7361);
and U10457 (N_10457,N_9971,N_5082);
or U10458 (N_10458,N_5290,N_7275);
and U10459 (N_10459,N_9736,N_5869);
and U10460 (N_10460,N_5322,N_5405);
and U10461 (N_10461,N_8130,N_7448);
or U10462 (N_10462,N_6044,N_9456);
and U10463 (N_10463,N_5294,N_8890);
xor U10464 (N_10464,N_7751,N_5702);
and U10465 (N_10465,N_8409,N_6897);
nor U10466 (N_10466,N_8999,N_8030);
or U10467 (N_10467,N_6334,N_6023);
and U10468 (N_10468,N_7529,N_6747);
nor U10469 (N_10469,N_6424,N_5639);
nand U10470 (N_10470,N_9720,N_8225);
and U10471 (N_10471,N_7471,N_5174);
nand U10472 (N_10472,N_5944,N_6977);
nand U10473 (N_10473,N_5242,N_9326);
and U10474 (N_10474,N_6134,N_5383);
and U10475 (N_10475,N_6326,N_7859);
nor U10476 (N_10476,N_8305,N_9915);
and U10477 (N_10477,N_8075,N_5590);
or U10478 (N_10478,N_7801,N_8905);
nor U10479 (N_10479,N_9134,N_8767);
nor U10480 (N_10480,N_5030,N_7284);
xnor U10481 (N_10481,N_8548,N_6085);
and U10482 (N_10482,N_6737,N_9717);
or U10483 (N_10483,N_8233,N_6018);
xor U10484 (N_10484,N_7342,N_7088);
nand U10485 (N_10485,N_9169,N_5436);
nor U10486 (N_10486,N_8512,N_8065);
and U10487 (N_10487,N_8628,N_5631);
and U10488 (N_10488,N_9084,N_7112);
nor U10489 (N_10489,N_6111,N_6154);
nand U10490 (N_10490,N_7840,N_6026);
and U10491 (N_10491,N_6399,N_9733);
nand U10492 (N_10492,N_5135,N_6448);
and U10493 (N_10493,N_7061,N_7843);
or U10494 (N_10494,N_9000,N_5027);
or U10495 (N_10495,N_8344,N_9754);
nand U10496 (N_10496,N_6955,N_9380);
and U10497 (N_10497,N_8655,N_9828);
nand U10498 (N_10498,N_7293,N_5683);
and U10499 (N_10499,N_8525,N_6291);
and U10500 (N_10500,N_5327,N_5251);
and U10501 (N_10501,N_6782,N_6834);
and U10502 (N_10502,N_9516,N_9726);
and U10503 (N_10503,N_6690,N_9809);
or U10504 (N_10504,N_7639,N_7681);
nand U10505 (N_10505,N_8560,N_5698);
nor U10506 (N_10506,N_9130,N_9186);
or U10507 (N_10507,N_6495,N_9909);
and U10508 (N_10508,N_9144,N_7878);
or U10509 (N_10509,N_6337,N_5177);
nand U10510 (N_10510,N_8388,N_5457);
and U10511 (N_10511,N_9108,N_6036);
xnor U10512 (N_10512,N_7373,N_7503);
and U10513 (N_10513,N_7569,N_6828);
or U10514 (N_10514,N_7982,N_6224);
or U10515 (N_10515,N_8600,N_6161);
and U10516 (N_10516,N_9816,N_5814);
nand U10517 (N_10517,N_7439,N_6956);
nor U10518 (N_10518,N_9617,N_6428);
and U10519 (N_10519,N_9598,N_5411);
and U10520 (N_10520,N_6904,N_9890);
and U10521 (N_10521,N_9109,N_6531);
and U10522 (N_10522,N_5213,N_5054);
and U10523 (N_10523,N_9228,N_6730);
nand U10524 (N_10524,N_6759,N_6858);
or U10525 (N_10525,N_8025,N_5391);
and U10526 (N_10526,N_5925,N_7004);
and U10527 (N_10527,N_7306,N_6972);
or U10528 (N_10528,N_6567,N_9227);
nand U10529 (N_10529,N_7146,N_6391);
nand U10530 (N_10530,N_5085,N_7913);
or U10531 (N_10531,N_8306,N_6639);
and U10532 (N_10532,N_5422,N_8945);
and U10533 (N_10533,N_9585,N_9674);
nor U10534 (N_10534,N_9016,N_9767);
nand U10535 (N_10535,N_9075,N_8517);
and U10536 (N_10536,N_9416,N_6062);
nor U10537 (N_10537,N_5459,N_7472);
and U10538 (N_10538,N_9341,N_9050);
and U10539 (N_10539,N_5980,N_6059);
nor U10540 (N_10540,N_5554,N_7548);
nor U10541 (N_10541,N_6996,N_6460);
and U10542 (N_10542,N_8019,N_7970);
or U10543 (N_10543,N_8106,N_6318);
nand U10544 (N_10544,N_8712,N_5985);
nand U10545 (N_10545,N_6159,N_9082);
nor U10546 (N_10546,N_9770,N_7635);
and U10547 (N_10547,N_6580,N_6413);
nor U10548 (N_10548,N_6647,N_8126);
and U10549 (N_10549,N_9247,N_5224);
nor U10550 (N_10550,N_8271,N_6063);
nor U10551 (N_10551,N_5295,N_9780);
nor U10552 (N_10552,N_7064,N_6136);
nand U10553 (N_10553,N_7206,N_7987);
or U10554 (N_10554,N_9626,N_7379);
or U10555 (N_10555,N_6474,N_8097);
or U10556 (N_10556,N_8407,N_7705);
or U10557 (N_10557,N_9906,N_6335);
or U10558 (N_10558,N_8985,N_9033);
nor U10559 (N_10559,N_6498,N_8889);
or U10560 (N_10560,N_6677,N_6416);
and U10561 (N_10561,N_6924,N_9904);
and U10562 (N_10562,N_7059,N_6158);
or U10563 (N_10563,N_9737,N_7795);
nand U10564 (N_10564,N_7584,N_7097);
nor U10565 (N_10565,N_7012,N_8165);
or U10566 (N_10566,N_5876,N_6295);
nand U10567 (N_10567,N_9764,N_8949);
and U10568 (N_10568,N_5972,N_8393);
or U10569 (N_10569,N_9468,N_6361);
nor U10570 (N_10570,N_8710,N_5014);
xor U10571 (N_10571,N_6723,N_7651);
nor U10572 (N_10572,N_5196,N_5355);
and U10573 (N_10573,N_5549,N_7609);
nand U10574 (N_10574,N_9666,N_6072);
or U10575 (N_10575,N_7169,N_8496);
nand U10576 (N_10576,N_7063,N_5832);
nand U10577 (N_10577,N_7250,N_5222);
and U10578 (N_10578,N_8433,N_8916);
nor U10579 (N_10579,N_5914,N_7191);
and U10580 (N_10580,N_9284,N_6166);
or U10581 (N_10581,N_8400,N_5379);
and U10582 (N_10582,N_6962,N_9215);
nor U10583 (N_10583,N_6398,N_7787);
nor U10584 (N_10584,N_6452,N_7675);
nor U10585 (N_10585,N_6894,N_7537);
nand U10586 (N_10586,N_9157,N_8077);
and U10587 (N_10587,N_6842,N_8135);
nand U10588 (N_10588,N_8571,N_6073);
nor U10589 (N_10589,N_9363,N_7230);
nand U10590 (N_10590,N_8208,N_6687);
or U10591 (N_10591,N_7559,N_5056);
or U10592 (N_10592,N_9274,N_7873);
xor U10593 (N_10593,N_5812,N_7499);
or U10594 (N_10594,N_7742,N_7107);
and U10595 (N_10595,N_9453,N_8378);
nand U10596 (N_10596,N_9479,N_8341);
nor U10597 (N_10597,N_6218,N_9459);
nor U10598 (N_10598,N_9581,N_7197);
nand U10599 (N_10599,N_9757,N_8758);
and U10600 (N_10600,N_6195,N_5529);
or U10601 (N_10601,N_7558,N_6090);
nand U10602 (N_10602,N_5334,N_8480);
or U10603 (N_10603,N_8953,N_7046);
nor U10604 (N_10604,N_8037,N_9684);
nand U10605 (N_10605,N_5116,N_5374);
nand U10606 (N_10606,N_9076,N_7547);
nand U10607 (N_10607,N_9234,N_6126);
nand U10608 (N_10608,N_9690,N_5226);
nand U10609 (N_10609,N_6382,N_5342);
and U10610 (N_10610,N_9354,N_5720);
nand U10611 (N_10611,N_9349,N_7313);
and U10612 (N_10612,N_8457,N_6205);
or U10613 (N_10613,N_6995,N_8968);
or U10614 (N_10614,N_9729,N_7409);
nand U10615 (N_10615,N_8656,N_9525);
and U10616 (N_10616,N_8468,N_9507);
nor U10617 (N_10617,N_5477,N_6585);
nand U10618 (N_10618,N_5332,N_6583);
xor U10619 (N_10619,N_6392,N_5075);
nor U10620 (N_10620,N_5642,N_6270);
nand U10621 (N_10621,N_6767,N_8546);
and U10622 (N_10622,N_6643,N_7560);
or U10623 (N_10623,N_7417,N_5050);
nor U10624 (N_10624,N_5668,N_9662);
or U10625 (N_10625,N_7964,N_8462);
nor U10626 (N_10626,N_5961,N_6322);
nor U10627 (N_10627,N_7904,N_6106);
nand U10628 (N_10628,N_6514,N_9898);
and U10629 (N_10629,N_9436,N_7334);
nor U10630 (N_10630,N_5108,N_8808);
nor U10631 (N_10631,N_8184,N_5951);
nor U10632 (N_10632,N_9792,N_8131);
or U10633 (N_10633,N_9180,N_6659);
nand U10634 (N_10634,N_6591,N_7369);
or U10635 (N_10635,N_8251,N_5518);
or U10636 (N_10636,N_9892,N_7320);
or U10637 (N_10637,N_8668,N_5645);
and U10638 (N_10638,N_6067,N_8859);
nor U10639 (N_10639,N_7699,N_6199);
nand U10640 (N_10640,N_8989,N_6953);
nor U10641 (N_10641,N_9044,N_9984);
nor U10642 (N_10642,N_6772,N_5741);
or U10643 (N_10643,N_8633,N_6629);
xor U10644 (N_10644,N_5104,N_6509);
nand U10645 (N_10645,N_9964,N_9727);
and U10646 (N_10646,N_7641,N_6143);
and U10647 (N_10647,N_7928,N_5386);
nand U10648 (N_10648,N_7190,N_8900);
or U10649 (N_10649,N_7977,N_5299);
nor U10650 (N_10650,N_8211,N_9911);
nor U10651 (N_10651,N_8595,N_7520);
and U10652 (N_10652,N_8262,N_9047);
nand U10653 (N_10653,N_8396,N_8756);
xnor U10654 (N_10654,N_6952,N_6780);
nor U10655 (N_10655,N_5421,N_8638);
and U10656 (N_10656,N_7953,N_9491);
and U10657 (N_10657,N_9422,N_5298);
or U10658 (N_10658,N_6563,N_7030);
nand U10659 (N_10659,N_9414,N_8919);
or U10660 (N_10660,N_8071,N_7722);
nor U10661 (N_10661,N_5735,N_6459);
nand U10662 (N_10662,N_5975,N_7680);
and U10663 (N_10663,N_9797,N_9437);
nand U10664 (N_10664,N_6117,N_7889);
or U10665 (N_10665,N_6045,N_6758);
nand U10666 (N_10666,N_6776,N_6727);
nor U10667 (N_10667,N_9930,N_6991);
and U10668 (N_10668,N_9242,N_7685);
nor U10669 (N_10669,N_5850,N_6801);
nor U10670 (N_10670,N_7199,N_8974);
and U10671 (N_10671,N_6266,N_5781);
nor U10672 (N_10672,N_6543,N_8138);
nor U10673 (N_10673,N_9866,N_8765);
or U10674 (N_10674,N_6348,N_7568);
nand U10675 (N_10675,N_9997,N_5286);
or U10676 (N_10676,N_5649,N_8014);
nand U10677 (N_10677,N_5235,N_6950);
or U10678 (N_10678,N_9389,N_7968);
and U10679 (N_10679,N_7701,N_6079);
or U10680 (N_10680,N_6209,N_6746);
nor U10681 (N_10681,N_5509,N_8884);
nand U10682 (N_10682,N_5802,N_9237);
nor U10683 (N_10683,N_5091,N_8770);
or U10684 (N_10684,N_6155,N_5667);
nor U10685 (N_10685,N_7516,N_9224);
nand U10686 (N_10686,N_7131,N_8619);
nand U10687 (N_10687,N_5057,N_6976);
or U10688 (N_10688,N_5128,N_8799);
and U10689 (N_10689,N_8862,N_8171);
or U10690 (N_10690,N_6148,N_9693);
or U10691 (N_10691,N_9558,N_6037);
and U10692 (N_10692,N_7427,N_6173);
and U10693 (N_10693,N_9587,N_5148);
xor U10694 (N_10694,N_9022,N_7128);
nor U10695 (N_10695,N_5195,N_6512);
nor U10696 (N_10696,N_8047,N_6010);
and U10697 (N_10697,N_5722,N_5105);
nor U10698 (N_10698,N_9608,N_7195);
nand U10699 (N_10699,N_5456,N_6381);
or U10700 (N_10700,N_6938,N_7136);
or U10701 (N_10701,N_8626,N_8080);
nand U10702 (N_10702,N_9745,N_7980);
and U10703 (N_10703,N_5331,N_5711);
nand U10704 (N_10704,N_9591,N_5369);
nand U10705 (N_10705,N_9353,N_5935);
or U10706 (N_10706,N_6115,N_6919);
nor U10707 (N_10707,N_8834,N_8567);
or U10708 (N_10708,N_9364,N_5497);
and U10709 (N_10709,N_8689,N_7218);
nor U10710 (N_10710,N_9957,N_7363);
and U10711 (N_10711,N_9490,N_9140);
and U10712 (N_10712,N_8372,N_6823);
or U10713 (N_10713,N_6619,N_5423);
and U10714 (N_10714,N_9092,N_7029);
nand U10715 (N_10715,N_8127,N_7247);
and U10716 (N_10716,N_9488,N_8048);
and U10717 (N_10717,N_5390,N_6366);
and U10718 (N_10718,N_6542,N_6104);
nand U10719 (N_10719,N_5620,N_9498);
or U10720 (N_10720,N_8173,N_7359);
and U10721 (N_10721,N_6001,N_7881);
nand U10722 (N_10722,N_7274,N_6553);
or U10723 (N_10723,N_7886,N_8349);
nand U10724 (N_10724,N_6373,N_6606);
nor U10725 (N_10725,N_6501,N_5191);
nor U10726 (N_10726,N_6631,N_5632);
nand U10727 (N_10727,N_7051,N_7598);
and U10728 (N_10728,N_6657,N_5889);
or U10729 (N_10729,N_8887,N_9423);
nor U10730 (N_10730,N_9853,N_7469);
and U10731 (N_10731,N_9774,N_7773);
or U10732 (N_10732,N_6103,N_9632);
or U10733 (N_10733,N_9800,N_9746);
xnor U10734 (N_10734,N_6941,N_7720);
nor U10735 (N_10735,N_9777,N_5958);
nor U10736 (N_10736,N_7602,N_6750);
nor U10737 (N_10737,N_8753,N_5393);
nand U10738 (N_10738,N_7619,N_8778);
nor U10739 (N_10739,N_8160,N_8152);
nand U10740 (N_10740,N_9279,N_8427);
or U10741 (N_10741,N_8583,N_8221);
and U10742 (N_10742,N_9376,N_8379);
nor U10743 (N_10743,N_6957,N_5005);
or U10744 (N_10744,N_7939,N_5819);
or U10745 (N_10745,N_9373,N_5107);
nand U10746 (N_10746,N_9327,N_7198);
nor U10747 (N_10747,N_9787,N_5435);
or U10748 (N_10748,N_9564,N_5759);
and U10749 (N_10749,N_5965,N_7295);
and U10750 (N_10750,N_6742,N_8789);
and U10751 (N_10751,N_5333,N_6676);
nand U10752 (N_10752,N_7084,N_7057);
nand U10753 (N_10753,N_8230,N_8651);
or U10754 (N_10754,N_8681,N_7709);
or U10755 (N_10755,N_7834,N_7515);
and U10756 (N_10756,N_9207,N_7490);
and U10757 (N_10757,N_9978,N_9723);
and U10758 (N_10758,N_7425,N_8389);
nand U10759 (N_10759,N_9649,N_8134);
nor U10760 (N_10760,N_8674,N_9704);
or U10761 (N_10761,N_8837,N_6609);
and U10762 (N_10762,N_9506,N_7350);
nand U10763 (N_10763,N_5885,N_6735);
or U10764 (N_10764,N_6819,N_9473);
nor U10765 (N_10765,N_9297,N_7103);
nand U10766 (N_10766,N_5115,N_6588);
or U10767 (N_10767,N_7926,N_5699);
and U10768 (N_10768,N_6810,N_7744);
nor U10769 (N_10769,N_5559,N_9603);
and U10770 (N_10770,N_9160,N_9807);
nand U10771 (N_10771,N_9291,N_5163);
nand U10772 (N_10772,N_8013,N_9755);
or U10773 (N_10773,N_6980,N_5336);
and U10774 (N_10774,N_8453,N_8099);
or U10775 (N_10775,N_6787,N_6789);
nand U10776 (N_10776,N_5134,N_6786);
nand U10777 (N_10777,N_6638,N_9882);
or U10778 (N_10778,N_7767,N_6646);
and U10779 (N_10779,N_9942,N_9639);
nand U10780 (N_10780,N_7120,N_7337);
nor U10781 (N_10781,N_9379,N_8464);
and U10782 (N_10782,N_5062,N_9202);
and U10783 (N_10783,N_7140,N_5356);
nor U10784 (N_10784,N_7303,N_9962);
and U10785 (N_10785,N_7179,N_7757);
nor U10786 (N_10786,N_7952,N_6298);
or U10787 (N_10787,N_7497,N_8011);
nand U10788 (N_10788,N_9766,N_6308);
nor U10789 (N_10789,N_6120,N_9396);
nor U10790 (N_10790,N_9621,N_9825);
nand U10791 (N_10791,N_7354,N_5126);
nor U10792 (N_10792,N_5721,N_9118);
or U10793 (N_10793,N_6095,N_5145);
xnor U10794 (N_10794,N_9080,N_6616);
and U10795 (N_10795,N_8273,N_9410);
or U10796 (N_10796,N_8729,N_8860);
and U10797 (N_10797,N_7921,N_5930);
and U10798 (N_10798,N_9112,N_9855);
nand U10799 (N_10799,N_7341,N_8227);
or U10800 (N_10800,N_8491,N_7726);
nand U10801 (N_10801,N_6668,N_8997);
nor U10802 (N_10802,N_9966,N_5792);
nand U10803 (N_10803,N_5778,N_8952);
or U10804 (N_10804,N_6029,N_8346);
and U10805 (N_10805,N_5439,N_9034);
nor U10806 (N_10806,N_5614,N_9013);
nand U10807 (N_10807,N_5168,N_8091);
nand U10808 (N_10808,N_5230,N_8133);
nand U10809 (N_10809,N_7060,N_7902);
nand U10810 (N_10810,N_9992,N_8288);
or U10811 (N_10811,N_9170,N_5192);
nand U10812 (N_10812,N_8821,N_8461);
or U10813 (N_10813,N_7377,N_9124);
nor U10814 (N_10814,N_5782,N_9919);
nand U10815 (N_10815,N_8722,N_6741);
xor U10816 (N_10816,N_6673,N_7822);
or U10817 (N_10817,N_6589,N_7624);
or U10818 (N_10818,N_9171,N_9395);
and U10819 (N_10819,N_5677,N_8286);
or U10820 (N_10820,N_7485,N_6411);
and U10821 (N_10821,N_9387,N_6475);
nand U10822 (N_10822,N_5253,N_7662);
or U10823 (N_10823,N_6626,N_7653);
nand U10824 (N_10824,N_9699,N_9368);
nor U10825 (N_10825,N_5872,N_9527);
or U10826 (N_10826,N_8736,N_5627);
nand U10827 (N_10827,N_6347,N_6679);
or U10828 (N_10828,N_9036,N_7022);
nand U10829 (N_10829,N_5528,N_6804);
nor U10830 (N_10830,N_8079,N_5793);
or U10831 (N_10831,N_7324,N_7868);
or U10832 (N_10832,N_5706,N_5166);
or U10833 (N_10833,N_8497,N_5485);
or U10834 (N_10834,N_5540,N_9761);
or U10835 (N_10835,N_7127,N_8268);
nand U10836 (N_10836,N_5795,N_7091);
nand U10837 (N_10837,N_9859,N_8672);
nand U10838 (N_10838,N_8992,N_5033);
and U10839 (N_10839,N_8197,N_6614);
nor U10840 (N_10840,N_6945,N_9605);
or U10841 (N_10841,N_9731,N_6749);
nand U10842 (N_10842,N_6743,N_9344);
nand U10843 (N_10843,N_7261,N_9318);
and U10844 (N_10844,N_8733,N_7799);
or U10845 (N_10845,N_5752,N_6939);
nor U10846 (N_10846,N_9752,N_5498);
and U10847 (N_10847,N_5887,N_9018);
nand U10848 (N_10848,N_5616,N_7412);
and U10849 (N_10849,N_5610,N_5736);
and U10850 (N_10850,N_6213,N_7085);
or U10851 (N_10851,N_9847,N_7973);
nor U10852 (N_10852,N_8563,N_7554);
or U10853 (N_10853,N_8590,N_7562);
and U10854 (N_10854,N_8854,N_8249);
and U10855 (N_10855,N_9985,N_5829);
nand U10856 (N_10856,N_7043,N_9064);
nor U10857 (N_10857,N_9884,N_8259);
or U10858 (N_10858,N_9358,N_8129);
or U10859 (N_10859,N_6884,N_9464);
nor U10860 (N_10860,N_6071,N_8676);
and U10861 (N_10861,N_8796,N_6217);
or U10862 (N_10862,N_5862,N_6305);
nor U10863 (N_10863,N_8593,N_8142);
or U10864 (N_10864,N_7845,N_6022);
and U10865 (N_10865,N_5502,N_5917);
nor U10866 (N_10866,N_7603,N_5587);
nor U10867 (N_10867,N_8501,N_8697);
nor U10868 (N_10868,N_7126,N_5444);
nand U10869 (N_10869,N_6880,N_7038);
nor U10870 (N_10870,N_5074,N_5387);
nand U10871 (N_10871,N_5727,N_7065);
nor U10872 (N_10872,N_5543,N_7115);
nor U10873 (N_10873,N_8613,N_5568);
or U10874 (N_10874,N_6734,N_6843);
nand U10875 (N_10875,N_9249,N_6925);
nor U10876 (N_10876,N_7400,N_8214);
xor U10877 (N_10877,N_5879,N_8519);
nand U10878 (N_10878,N_7344,N_6169);
and U10879 (N_10879,N_5595,N_9653);
nand U10880 (N_10880,N_9889,N_9482);
nor U10881 (N_10881,N_5831,N_9428);
nor U10882 (N_10882,N_5416,N_6635);
nor U10883 (N_10883,N_7892,N_6648);
nor U10884 (N_10884,N_5801,N_9086);
nand U10885 (N_10885,N_6602,N_9319);
xnor U10886 (N_10886,N_7864,N_5478);
and U10887 (N_10887,N_5539,N_7941);
nand U10888 (N_10888,N_6833,N_7044);
nor U10889 (N_10889,N_6597,N_6255);
nand U10890 (N_10890,N_8774,N_6066);
and U10891 (N_10891,N_8631,N_9366);
nor U10892 (N_10892,N_9040,N_8570);
nor U10893 (N_10893,N_9383,N_8327);
or U10894 (N_10894,N_8046,N_7391);
and U10895 (N_10895,N_8698,N_7652);
and U10896 (N_10896,N_9826,N_6457);
nand U10897 (N_10897,N_5335,N_6412);
xor U10898 (N_10898,N_6562,N_5522);
nand U10899 (N_10899,N_6527,N_7114);
and U10900 (N_10900,N_5505,N_5340);
nand U10901 (N_10901,N_5398,N_8290);
nor U10902 (N_10902,N_6319,N_9524);
or U10903 (N_10903,N_8300,N_5271);
or U10904 (N_10904,N_7853,N_9878);
or U10905 (N_10905,N_7937,N_5923);
and U10906 (N_10906,N_6471,N_6798);
nand U10907 (N_10907,N_6954,N_6362);
nand U10908 (N_10908,N_8816,N_5973);
nor U10909 (N_10909,N_7884,N_9658);
and U10910 (N_10910,N_5533,N_7781);
nand U10911 (N_10911,N_8966,N_7862);
and U10912 (N_10912,N_5184,N_6407);
and U10913 (N_10913,N_5245,N_6444);
or U10914 (N_10914,N_6110,N_9912);
nand U10915 (N_10915,N_7991,N_6153);
and U10916 (N_10916,N_5160,N_5450);
or U10917 (N_10917,N_8269,N_6489);
nand U10918 (N_10918,N_7316,N_8090);
or U10919 (N_10919,N_6875,N_7809);
nor U10920 (N_10920,N_9973,N_6076);
or U10921 (N_10921,N_8353,N_7145);
or U10922 (N_10922,N_9595,N_7352);
and U10923 (N_10923,N_6327,N_6959);
and U10924 (N_10924,N_8128,N_9739);
or U10925 (N_10925,N_7028,N_9923);
nand U10926 (N_10926,N_5723,N_8718);
nand U10927 (N_10927,N_8643,N_6070);
and U10928 (N_10928,N_8166,N_8278);
xnor U10929 (N_10929,N_5306,N_5310);
and U10930 (N_10930,N_6272,N_8467);
or U10931 (N_10931,N_9178,N_5583);
nand U10932 (N_10932,N_8164,N_8897);
nand U10933 (N_10933,N_8743,N_7166);
nand U10934 (N_10934,N_9059,N_5349);
nor U10935 (N_10935,N_5896,N_9101);
or U10936 (N_10936,N_7670,N_9863);
nand U10937 (N_10937,N_6763,N_6287);
nor U10938 (N_10938,N_7264,N_9392);
or U10939 (N_10939,N_8029,N_7957);
nand U10940 (N_10940,N_9779,N_9362);
and U10941 (N_10941,N_6310,N_6861);
nand U10942 (N_10942,N_5208,N_9907);
and U10943 (N_10943,N_9751,N_7347);
and U10944 (N_10944,N_7403,N_7703);
or U10945 (N_10945,N_9829,N_8023);
or U10946 (N_10946,N_5373,N_9469);
nor U10947 (N_10947,N_6752,N_8484);
nand U10948 (N_10948,N_6935,N_8034);
nand U10949 (N_10949,N_8584,N_7903);
nor U10950 (N_10950,N_8317,N_6182);
and U10951 (N_10951,N_5628,N_7006);
or U10952 (N_10952,N_7013,N_5078);
xor U10953 (N_10953,N_7623,N_5506);
and U10954 (N_10954,N_5084,N_7310);
and U10955 (N_10955,N_6133,N_8727);
or U10956 (N_10956,N_7567,N_9049);
nor U10957 (N_10957,N_8891,N_6453);
and U10958 (N_10958,N_9273,N_7586);
and U10959 (N_10959,N_8183,N_7089);
nor U10960 (N_10960,N_9860,N_7183);
or U10961 (N_10961,N_8364,N_7222);
and U10962 (N_10962,N_6573,N_6128);
nor U10963 (N_10963,N_7495,N_8709);
nor U10964 (N_10964,N_7348,N_5746);
and U10965 (N_10965,N_7185,N_9660);
nand U10966 (N_10966,N_6164,N_5531);
nor U10967 (N_10967,N_8119,N_5813);
and U10968 (N_10968,N_6966,N_9316);
nand U10969 (N_10969,N_8261,N_8964);
nand U10970 (N_10970,N_7374,N_9494);
nand U10971 (N_10971,N_7814,N_9994);
nand U10972 (N_10972,N_6105,N_5034);
or U10973 (N_10973,N_6030,N_6239);
nand U10974 (N_10974,N_5501,N_5834);
or U10975 (N_10975,N_6601,N_7393);
and U10976 (N_10976,N_8726,N_6329);
or U10977 (N_10977,N_6288,N_7453);
xor U10978 (N_10978,N_7988,N_8870);
nand U10979 (N_10979,N_8582,N_7704);
and U10980 (N_10980,N_8108,N_8328);
nand U10981 (N_10981,N_7765,N_8161);
or U10982 (N_10982,N_7714,N_6028);
and U10983 (N_10983,N_9245,N_8283);
or U10984 (N_10984,N_8840,N_5418);
or U10985 (N_10985,N_6699,N_5527);
nor U10986 (N_10986,N_5219,N_5320);
or U10987 (N_10987,N_9230,N_5892);
and U10988 (N_10988,N_6813,N_5260);
nand U10989 (N_10989,N_5206,N_6986);
nor U10990 (N_10990,N_6584,N_6806);
nand U10991 (N_10991,N_6764,N_5799);
or U10992 (N_10992,N_8412,N_6089);
or U10993 (N_10993,N_7282,N_8136);
and U10994 (N_10994,N_8741,N_5758);
or U10995 (N_10995,N_8425,N_7629);
nand U10996 (N_10996,N_8350,N_8148);
and U10997 (N_10997,N_6805,N_7171);
and U10998 (N_10998,N_9715,N_8362);
nor U10999 (N_10999,N_7224,N_6523);
nand U11000 (N_11000,N_7875,N_6341);
nor U11001 (N_11001,N_7918,N_5169);
nor U11002 (N_11002,N_7542,N_8301);
nor U11003 (N_11003,N_8296,N_8151);
and U11004 (N_11004,N_9266,N_8263);
nor U11005 (N_11005,N_5655,N_7147);
nor U11006 (N_11006,N_6738,N_7216);
nor U11007 (N_11007,N_5825,N_6464);
nand U11008 (N_11008,N_7501,N_7986);
and U11009 (N_11009,N_6525,N_9312);
and U11010 (N_11010,N_5442,N_5388);
or U11011 (N_11011,N_9876,N_9301);
and U11012 (N_11012,N_9712,N_7932);
and U11013 (N_11013,N_5519,N_8081);
or U11014 (N_11014,N_6118,N_5574);
nor U11015 (N_11015,N_9635,N_5982);
xor U11016 (N_11016,N_9339,N_9665);
nand U11017 (N_11017,N_8951,N_7807);
or U11018 (N_11018,N_8677,N_6550);
nor U11019 (N_11019,N_6049,N_7506);
and U11020 (N_11020,N_9902,N_6728);
or U11021 (N_11021,N_7766,N_7721);
and U11022 (N_11022,N_6447,N_7245);
and U11023 (N_11023,N_8701,N_5974);
and U11024 (N_11024,N_9151,N_6982);
nand U11025 (N_11025,N_9599,N_9793);
and U11026 (N_11026,N_6415,N_7999);
nor U11027 (N_11027,N_6102,N_9007);
or U11028 (N_11028,N_5055,N_9365);
or U11029 (N_11029,N_7049,N_7151);
or U11030 (N_11030,N_8052,N_5670);
nand U11031 (N_11031,N_9530,N_7577);
or U11032 (N_11032,N_7710,N_5409);
or U11033 (N_11033,N_8418,N_8740);
and U11034 (N_11034,N_7015,N_9480);
xnor U11035 (N_11035,N_7813,N_9011);
or U11036 (N_11036,N_6963,N_7221);
or U11037 (N_11037,N_6053,N_8640);
or U11038 (N_11038,N_5025,N_6771);
or U11039 (N_11039,N_7387,N_9150);
nand U11040 (N_11040,N_5314,N_7583);
and U11041 (N_11041,N_5353,N_5952);
or U11042 (N_11042,N_7464,N_6055);
nand U11043 (N_11043,N_7188,N_7263);
nor U11044 (N_11044,N_6706,N_9544);
or U11045 (N_11045,N_8476,N_5288);
or U11046 (N_11046,N_7433,N_9848);
nor U11047 (N_11047,N_9688,N_9550);
nand U11048 (N_11048,N_7144,N_6183);
nand U11049 (N_11049,N_6432,N_9830);
nand U11050 (N_11050,N_8661,N_5366);
nand U11051 (N_11051,N_8483,N_8096);
nand U11052 (N_11052,N_5880,N_8436);
nand U11053 (N_11053,N_8202,N_6033);
nor U11054 (N_11054,N_6932,N_8397);
nor U11055 (N_11055,N_5049,N_6669);
or U11056 (N_11056,N_6485,N_6846);
and U11057 (N_11057,N_9394,N_8847);
and U11058 (N_11058,N_8384,N_8092);
and U11059 (N_11059,N_6092,N_7532);
and U11060 (N_11060,N_7226,N_5493);
nand U11061 (N_11061,N_8888,N_5364);
nand U11062 (N_11062,N_7649,N_7098);
and U11063 (N_11063,N_9407,N_5112);
or U11064 (N_11064,N_8456,N_9652);
and U11065 (N_11065,N_8623,N_7397);
nor U11066 (N_11066,N_5646,N_6025);
nor U11067 (N_11067,N_6034,N_5239);
nor U11068 (N_11068,N_5789,N_7096);
nand U11069 (N_11069,N_8669,N_9841);
and U11070 (N_11070,N_5297,N_9651);
and U11071 (N_11071,N_9537,N_5707);
xor U11072 (N_11072,N_5588,N_9765);
or U11073 (N_11073,N_7451,N_7405);
nand U11074 (N_11074,N_7995,N_7536);
nand U11075 (N_11075,N_8430,N_8542);
nand U11076 (N_11076,N_5484,N_5986);
nand U11077 (N_11077,N_6671,N_9357);
and U11078 (N_11078,N_6800,N_5089);
and U11079 (N_11079,N_5714,N_6792);
or U11080 (N_11080,N_6220,N_9289);
and U11081 (N_11081,N_6389,N_9164);
or U11082 (N_11082,N_6694,N_5052);
nor U11083 (N_11083,N_9214,N_6942);
nor U11084 (N_11084,N_9910,N_7326);
xnor U11085 (N_11085,N_6868,N_5313);
and U11086 (N_11086,N_9940,N_5991);
nand U11087 (N_11087,N_7187,N_8274);
or U11088 (N_11088,N_7648,N_9374);
and U11089 (N_11089,N_8956,N_8699);
xor U11090 (N_11090,N_8961,N_7368);
nor U11091 (N_11091,N_7552,N_9703);
xor U11092 (N_11092,N_6729,N_7580);
nand U11093 (N_11093,N_7437,N_8490);
or U11094 (N_11094,N_8602,N_6439);
nor U11095 (N_11095,N_5928,N_5859);
xor U11096 (N_11096,N_9209,N_8045);
nand U11097 (N_11097,N_7610,N_9610);
xor U11098 (N_11098,N_9163,N_7732);
nor U11099 (N_11099,N_9536,N_6185);
nand U11100 (N_11100,N_9071,N_7715);
and U11101 (N_11101,N_9532,N_7255);
nor U11102 (N_11102,N_9520,N_6634);
or U11103 (N_11103,N_9254,N_8207);
xnor U11104 (N_11104,N_6385,N_8421);
and U11105 (N_11105,N_7594,N_6569);
and U11106 (N_11106,N_5087,N_9200);
or U11107 (N_11107,N_5489,N_8549);
and U11108 (N_11108,N_9386,N_5407);
nand U11109 (N_11109,N_9946,N_7837);
nor U11110 (N_11110,N_5705,N_8326);
nand U11111 (N_11111,N_7105,N_9375);
or U11112 (N_11112,N_5648,N_9184);
and U11113 (N_11113,N_7009,N_9472);
nor U11114 (N_11114,N_6613,N_9505);
or U11115 (N_11115,N_8604,N_5229);
and U11116 (N_11116,N_5809,N_6374);
nand U11117 (N_11117,N_6756,N_9980);
and U11118 (N_11118,N_7314,N_6162);
nor U11119 (N_11119,N_7418,N_7962);
nor U11120 (N_11120,N_6630,N_8241);
or U11121 (N_11121,N_5047,N_5697);
nor U11122 (N_11122,N_8140,N_5357);
nor U11123 (N_11123,N_9814,N_7016);
nand U11124 (N_11124,N_8235,N_6704);
or U11125 (N_11125,N_6081,N_5503);
or U11126 (N_11126,N_7698,N_6561);
nor U11127 (N_11127,N_8947,N_8186);
nand U11128 (N_11128,N_9631,N_9175);
nor U11129 (N_11129,N_6020,N_7033);
nand U11130 (N_11130,N_6851,N_6779);
xor U11131 (N_11131,N_6965,N_8871);
or U11132 (N_11132,N_9248,N_8218);
nand U11133 (N_11133,N_9072,N_8627);
and U11134 (N_11134,N_8960,N_9594);
nand U11135 (N_11135,N_6974,N_8320);
or U11136 (N_11136,N_9367,N_7820);
and U11137 (N_11137,N_9026,N_8144);
or U11138 (N_11138,N_5179,N_8304);
nor U11139 (N_11139,N_9888,N_7607);
or U11140 (N_11140,N_9400,N_7678);
or U11141 (N_11141,N_8226,N_5545);
nor U11142 (N_11142,N_6225,N_6587);
nand U11143 (N_11143,N_7690,N_7110);
or U11144 (N_11144,N_8920,N_6644);
nand U11145 (N_11145,N_8612,N_8817);
nor U11146 (N_11146,N_9415,N_8556);
xor U11147 (N_11147,N_8819,N_5275);
and U11148 (N_11148,N_5753,N_8002);
or U11149 (N_11149,N_9614,N_9411);
or U11150 (N_11150,N_7866,N_7443);
nand U11151 (N_11151,N_9322,N_5384);
or U11152 (N_11152,N_7315,N_7857);
nand U11153 (N_11153,N_9159,N_6397);
nand U11154 (N_11154,N_5603,N_9628);
and U11155 (N_11155,N_5434,N_8242);
and U11156 (N_11156,N_7109,N_9749);
and U11157 (N_11157,N_6353,N_5742);
or U11158 (N_11158,N_7321,N_7413);
and U11159 (N_11159,N_5747,N_9190);
nor U11160 (N_11160,N_7553,N_5209);
xnor U11161 (N_11161,N_9880,N_5248);
nor U11162 (N_11162,N_5530,N_8356);
and U11163 (N_11163,N_9656,N_9384);
or U11164 (N_11164,N_6152,N_8392);
nor U11165 (N_11165,N_5894,N_6709);
nand U11166 (N_11166,N_9372,N_9433);
and U11167 (N_11167,N_6177,N_8180);
xnor U11168 (N_11168,N_6912,N_9937);
nor U11169 (N_11169,N_5765,N_9572);
and U11170 (N_11170,N_8666,N_5565);
nand U11171 (N_11171,N_7727,N_8469);
nor U11172 (N_11172,N_9513,N_6364);
or U11173 (N_11173,N_8624,N_5292);
or U11174 (N_11174,N_6024,N_6442);
nor U11175 (N_11175,N_7539,N_9509);
xor U11176 (N_11176,N_8597,N_8293);
and U11177 (N_11177,N_9053,N_5448);
and U11178 (N_11178,N_8239,N_5886);
and U11179 (N_11179,N_5458,N_7764);
nand U11180 (N_11180,N_9560,N_9642);
or U11181 (N_11181,N_6873,N_9310);
and U11182 (N_11182,N_6137,N_5001);
and U11183 (N_11183,N_5032,N_7946);
nand U11184 (N_11184,N_8167,N_6518);
or U11185 (N_11185,N_8452,N_5414);
or U11186 (N_11186,N_8351,N_6719);
nand U11187 (N_11187,N_7860,N_9540);
nand U11188 (N_11188,N_8146,N_6355);
xor U11189 (N_11189,N_5662,N_8750);
nand U11190 (N_11190,N_8150,N_9303);
nor U11191 (N_11191,N_9210,N_7683);
nor U11192 (N_11192,N_6108,N_8185);
and U11193 (N_11193,N_9398,N_6098);
nor U11194 (N_11194,N_7435,N_9775);
nand U11195 (N_11195,N_9035,N_5978);
or U11196 (N_11196,N_8311,N_6666);
nand U11197 (N_11197,N_6689,N_9321);
or U11198 (N_11198,N_9646,N_5482);
nand U11199 (N_11199,N_8885,N_9223);
and U11200 (N_11200,N_9831,N_7630);
or U11201 (N_11201,N_9672,N_5122);
nor U11202 (N_11202,N_8599,N_5954);
nor U11203 (N_11203,N_9531,N_5455);
and U11204 (N_11204,N_9600,N_7286);
nand U11205 (N_11205,N_6920,N_6356);
nand U11206 (N_11206,N_8500,N_7048);
or U11207 (N_11207,N_7338,N_9932);
and U11208 (N_11208,N_9500,N_9216);
nand U11209 (N_11209,N_7707,N_9404);
nand U11210 (N_11210,N_7576,N_5429);
nor U11211 (N_11211,N_5738,N_8544);
nor U11212 (N_11212,N_6440,N_7082);
and U11213 (N_11213,N_9686,N_6829);
nand U11214 (N_11214,N_5454,N_7299);
nand U11215 (N_11215,N_5136,N_7905);
and U11216 (N_11216,N_8552,N_6384);
or U11217 (N_11217,N_7036,N_8095);
nand U11218 (N_11218,N_9263,N_5856);
nand U11219 (N_11219,N_8818,N_6836);
or U11220 (N_11220,N_5623,N_6618);
nand U11221 (N_11221,N_8622,N_9314);
nor U11222 (N_11222,N_5447,N_8731);
and U11223 (N_11223,N_5636,N_8918);
nor U11224 (N_11224,N_7242,N_8963);
or U11225 (N_11225,N_8791,N_6312);
or U11226 (N_11226,N_7142,N_8598);
nand U11227 (N_11227,N_6064,N_6572);
and U11228 (N_11228,N_5984,N_5099);
nor U11229 (N_11229,N_6404,N_9689);
or U11230 (N_11230,N_5201,N_8852);
nor U11231 (N_11231,N_8454,N_9750);
nand U11232 (N_11232,N_8832,N_7430);
nor U11233 (N_11233,N_6219,N_6700);
nand U11234 (N_11234,N_6566,N_7677);
nor U11235 (N_11235,N_8781,N_7724);
or U11236 (N_11236,N_8078,N_8855);
or U11237 (N_11237,N_6050,N_5182);
nor U11238 (N_11238,N_5412,N_7798);
or U11239 (N_11239,N_5971,N_5556);
and U11240 (N_11240,N_5110,N_8688);
and U11241 (N_11241,N_7810,N_8367);
or U11242 (N_11242,N_9205,N_9802);
nand U11243 (N_11243,N_5690,N_7025);
and U11244 (N_11244,N_5061,N_8156);
nand U11245 (N_11245,N_9947,N_5775);
nand U11246 (N_11246,N_9442,N_5635);
or U11247 (N_11247,N_8543,N_6278);
nand U11248 (N_11248,N_5329,N_6262);
or U11249 (N_11249,N_5155,N_9891);
nand U11250 (N_11250,N_5159,N_9811);
nand U11251 (N_11251,N_6286,N_9203);
nor U11252 (N_11252,N_6087,N_5203);
nor U11253 (N_11253,N_9269,N_6486);
nor U11254 (N_11254,N_5515,N_6546);
nor U11255 (N_11255,N_9226,N_6046);
xor U11256 (N_11256,N_9338,N_7355);
nand U11257 (N_11257,N_5905,N_9241);
nand U11258 (N_11258,N_7728,N_6246);
nand U11259 (N_11259,N_9420,N_5983);
or U11260 (N_11260,N_9281,N_8691);
and U11261 (N_11261,N_5761,N_6112);
nand U11262 (N_11262,N_7281,N_9056);
nand U11263 (N_11263,N_5785,N_9673);
or U11264 (N_11264,N_7072,N_5381);
nor U11265 (N_11265,N_7931,N_9445);
and U11266 (N_11266,N_8299,N_9877);
nand U11267 (N_11267,N_9833,N_7204);
nor U11268 (N_11268,N_8083,N_8439);
nand U11269 (N_11269,N_5599,N_6321);
or U11270 (N_11270,N_5841,N_9547);
xnor U11271 (N_11271,N_5609,N_8471);
nor U11272 (N_11272,N_6916,N_8114);
or U11273 (N_11273,N_8442,N_8522);
or U11274 (N_11274,N_7487,N_9872);
or U11275 (N_11275,N_7058,N_7660);
and U11276 (N_11276,N_5146,N_7215);
nor U11277 (N_11277,N_9461,N_9856);
nor U11278 (N_11278,N_5425,N_8024);
nor U11279 (N_11279,N_9243,N_6716);
nand U11280 (N_11280,N_5114,N_6681);
nand U11281 (N_11281,N_6516,N_5534);
nor U11282 (N_11282,N_9462,N_9204);
xor U11283 (N_11283,N_5234,N_8406);
nor U11284 (N_11284,N_8463,N_6660);
nor U11285 (N_11285,N_7936,N_7071);
nand U11286 (N_11286,N_6774,N_6641);
and U11287 (N_11287,N_6113,N_6119);
nand U11288 (N_11288,N_6057,N_9768);
and U11289 (N_11289,N_6251,N_6521);
xor U11290 (N_11290,N_6838,N_5830);
and U11291 (N_11291,N_9128,N_7436);
and U11292 (N_11292,N_8715,N_8473);
xor U11293 (N_11293,N_8345,N_6077);
or U11294 (N_11294,N_7122,N_7010);
nand U11295 (N_11295,N_9125,N_8355);
nor U11296 (N_11296,N_9299,N_6497);
or U11297 (N_11297,N_7693,N_9005);
or U11298 (N_11298,N_9570,N_7538);
or U11299 (N_11299,N_5124,N_5466);
nand U11300 (N_11300,N_9408,N_8671);
nand U11301 (N_11301,N_5617,N_7003);
nor U11302 (N_11302,N_8693,N_9545);
and U11303 (N_11303,N_6088,N_6655);
nand U11304 (N_11304,N_8826,N_5178);
nand U11305 (N_11305,N_7656,N_6835);
or U11306 (N_11306,N_5571,N_8387);
and U11307 (N_11307,N_6610,N_8094);
nor U11308 (N_11308,N_8547,N_5853);
or U11309 (N_11309,N_6443,N_8260);
nor U11310 (N_11310,N_7605,N_9054);
nand U11311 (N_11311,N_5704,N_6150);
and U11312 (N_11312,N_5097,N_8763);
or U11313 (N_11313,N_7793,N_7175);
and U11314 (N_11314,N_8323,N_7201);
nor U11315 (N_11315,N_8169,N_8481);
or U11316 (N_11316,N_8403,N_9538);
nor U11317 (N_11317,N_9194,N_8835);
xor U11318 (N_11318,N_8331,N_6032);
or U11319 (N_11319,N_5264,N_6528);
and U11320 (N_11320,N_5664,N_6901);
nand U11321 (N_11321,N_6590,N_9123);
and U11322 (N_11322,N_5678,N_7459);
and U11323 (N_11323,N_6358,N_7466);
and U11324 (N_11324,N_6094,N_8502);
xor U11325 (N_11325,N_7031,N_8248);
nor U11326 (N_11326,N_5634,N_6282);
and U11327 (N_11327,N_7509,N_8093);
and U11328 (N_11328,N_7351,N_7650);
xor U11329 (N_11329,N_9533,N_9250);
nor U11330 (N_11330,N_8159,N_7632);
nor U11331 (N_11331,N_5371,N_9618);
or U11332 (N_11332,N_6989,N_6757);
and U11333 (N_11333,N_8800,N_5855);
nor U11334 (N_11334,N_9133,N_9261);
nor U11335 (N_11335,N_6803,N_8031);
or U11336 (N_11336,N_9185,N_9842);
or U11337 (N_11337,N_6340,N_9146);
nor U11338 (N_11338,N_5679,N_6368);
nand U11339 (N_11339,N_5739,N_6238);
or U11340 (N_11340,N_8361,N_7523);
or U11341 (N_11341,N_9868,N_6775);
and U11342 (N_11342,N_5641,N_6492);
xnor U11343 (N_11343,N_8401,N_7075);
nor U11344 (N_11344,N_9105,N_8177);
nand U11345 (N_11345,N_7916,N_8318);
nand U11346 (N_11346,N_6731,N_7113);
nand U11347 (N_11347,N_7068,N_6755);
or U11348 (N_11348,N_7129,N_6793);
nor U11349 (N_11349,N_6548,N_9953);
or U11350 (N_11350,N_6948,N_8478);
nor U11351 (N_11351,N_6394,N_8807);
nor U11352 (N_11352,N_5427,N_7802);
or U11353 (N_11353,N_7780,N_5346);
and U11354 (N_11354,N_8886,N_9094);
nand U11355 (N_11355,N_7273,N_9857);
nor U11356 (N_11356,N_5548,N_7888);
or U11357 (N_11357,N_5176,N_9418);
or U11358 (N_11358,N_5431,N_6850);
nand U11359 (N_11359,N_7050,N_8683);
nand U11360 (N_11360,N_8289,N_6652);
or U11361 (N_11361,N_9995,N_5339);
or U11362 (N_11362,N_8786,N_8673);
and U11363 (N_11363,N_7426,N_9702);
or U11364 (N_11364,N_6418,N_6039);
and U11365 (N_11365,N_6253,N_7011);
nand U11366 (N_11366,N_8100,N_9296);
and U11367 (N_11367,N_7687,N_8507);
nand U11368 (N_11368,N_5323,N_8118);
nand U11369 (N_11369,N_9131,N_8573);
and U11370 (N_11370,N_5804,N_8026);
nand U11371 (N_11371,N_7514,N_8754);
xor U11372 (N_11372,N_7234,N_8555);
and U11373 (N_11373,N_9290,N_7783);
and U11374 (N_11374,N_9449,N_7533);
or U11375 (N_11375,N_7959,N_8732);
nor U11376 (N_11376,N_7371,N_7659);
and U11377 (N_11377,N_8845,N_7130);
xnor U11378 (N_11378,N_6695,N_6309);
or U11379 (N_11379,N_7851,N_6047);
or U11380 (N_11380,N_8204,N_6693);
nand U11381 (N_11381,N_8322,N_6907);
and U11382 (N_11382,N_7135,N_8231);
and U11383 (N_11383,N_8381,N_5415);
or U11384 (N_11384,N_7301,N_7510);
nand U11385 (N_11385,N_6675,N_8205);
nor U11386 (N_11386,N_8394,N_9706);
nor U11387 (N_11387,N_5681,N_8564);
nor U11388 (N_11388,N_7979,N_8545);
and U11389 (N_11389,N_6297,N_5833);
or U11390 (N_11390,N_8329,N_5969);
nand U11391 (N_11391,N_6187,N_8324);
nor U11392 (N_11392,N_9999,N_8980);
nand U11393 (N_11393,N_5816,N_9862);
nor U11394 (N_11394,N_6944,N_9908);
or U11395 (N_11395,N_8064,N_9813);
and U11396 (N_11396,N_5827,N_7445);
and U11397 (N_11397,N_6973,N_5165);
and U11398 (N_11398,N_5018,N_9088);
and U11399 (N_11399,N_5093,N_9996);
nor U11400 (N_11400,N_6446,N_9655);
nor U11401 (N_11401,N_9342,N_5656);
and U11402 (N_11402,N_7268,N_7616);
or U11403 (N_11403,N_7719,N_9191);
and U11404 (N_11404,N_8653,N_6233);
xor U11405 (N_11405,N_9253,N_9001);
xor U11406 (N_11406,N_7730,N_8608);
xor U11407 (N_11407,N_6975,N_5228);
or U11408 (N_11408,N_9476,N_8865);
nand U11409 (N_11409,N_8285,N_5576);
nand U11410 (N_11410,N_7482,N_5360);
and U11411 (N_11411,N_6680,N_9694);
and U11412 (N_11412,N_5080,N_7565);
nand U11413 (N_11413,N_9869,N_9235);
nor U11414 (N_11414,N_6878,N_8302);
or U11415 (N_11415,N_5981,N_6593);
nand U11416 (N_11416,N_7461,N_6603);
or U11417 (N_11417,N_5396,N_7748);
and U11418 (N_11418,N_8199,N_8940);
and U11419 (N_11419,N_9066,N_7056);
nor U11420 (N_11420,N_6400,N_5593);
nor U11421 (N_11421,N_7396,N_9346);
and U11422 (N_11422,N_8357,N_8935);
nor U11423 (N_11423,N_5009,N_6724);
nor U11424 (N_11424,N_7723,N_7139);
nand U11425 (N_11425,N_6898,N_8374);
nand U11426 (N_11426,N_7305,N_6867);
nand U11427 (N_11427,N_5270,N_6084);
or U11428 (N_11428,N_6425,N_5237);
or U11429 (N_11429,N_8121,N_5012);
nor U11430 (N_11430,N_7007,N_8804);
or U11431 (N_11431,N_5675,N_7919);
nor U11432 (N_11432,N_5601,N_5188);
nand U11433 (N_11433,N_6140,N_9784);
nor U11434 (N_11434,N_8284,N_8149);
or U11435 (N_11435,N_8342,N_5133);
and U11436 (N_11436,N_8053,N_8880);
nand U11437 (N_11437,N_8087,N_6414);
nand U11438 (N_11438,N_5729,N_8338);
nor U11439 (N_11439,N_8244,N_7702);
or U11440 (N_11440,N_7848,N_6473);
and U11441 (N_11441,N_9905,N_9926);
nor U11442 (N_11442,N_7611,N_6201);
nand U11443 (N_11443,N_5004,N_6250);
nand U11444 (N_11444,N_9287,N_9330);
nor U11445 (N_11445,N_7971,N_7158);
nor U11446 (N_11446,N_9798,N_5573);
or U11447 (N_11447,N_9728,N_8944);
and U11448 (N_11448,N_5250,N_7502);
nor U11449 (N_11449,N_6832,N_9065);
and U11450 (N_11450,N_9791,N_5045);
nand U11451 (N_11451,N_6376,N_9038);
or U11452 (N_11452,N_9238,N_6783);
nand U11453 (N_11453,N_6441,N_8684);
or U11454 (N_11454,N_9502,N_6456);
nand U11455 (N_11455,N_7750,N_6862);
nor U11456 (N_11456,N_6654,N_5619);
and U11457 (N_11457,N_5138,N_5682);
or U11458 (N_11458,N_7081,N_6913);
and U11459 (N_11459,N_6339,N_5776);
nor U11460 (N_11460,N_7642,N_7346);
nand U11461 (N_11461,N_5101,N_6578);
and U11462 (N_11462,N_5268,N_7596);
nand U11463 (N_11463,N_6292,N_7184);
nor U11464 (N_11464,N_5626,N_9921);
or U11465 (N_11465,N_8931,N_9526);
xor U11466 (N_11466,N_7531,N_8906);
nor U11467 (N_11467,N_6852,N_8215);
nand U11468 (N_11468,N_9337,N_7005);
nand U11469 (N_11469,N_5324,N_9559);
nand U11470 (N_11470,N_8245,N_8679);
or U11471 (N_11471,N_9773,N_9206);
nor U11472 (N_11472,N_5818,N_5304);
nor U11473 (N_11473,N_9285,N_9606);
and U11474 (N_11474,N_5162,N_5205);
or U11475 (N_11475,N_7638,N_5561);
and U11476 (N_11476,N_5582,N_6256);
or U11477 (N_11477,N_5694,N_5939);
nand U11478 (N_11478,N_5467,N_8005);
nor U11479 (N_11479,N_9920,N_6328);
or U11480 (N_11480,N_5514,N_5053);
or U11481 (N_11481,N_7035,N_8746);
nand U11482 (N_11482,N_5602,N_7017);
and U11483 (N_11483,N_9553,N_5408);
and U11484 (N_11484,N_7657,N_9493);
nor U11485 (N_11485,N_7420,N_6146);
and U11486 (N_11486,N_6135,N_7841);
nor U11487 (N_11487,N_6258,N_6450);
nor U11488 (N_11488,N_8040,N_8103);
and U11489 (N_11489,N_6985,N_5608);
and U11490 (N_11490,N_8404,N_8508);
or U11491 (N_11491,N_6380,N_8667);
nor U11492 (N_11492,N_8440,N_5560);
and U11493 (N_11493,N_7238,N_8041);
nor U11494 (N_11494,N_8682,N_9725);
or U11495 (N_11495,N_5949,N_7100);
nand U11496 (N_11496,N_5432,N_7308);
nand U11497 (N_11497,N_8706,N_6605);
nand U11498 (N_11498,N_8371,N_8098);
or U11499 (N_11499,N_7398,N_6274);
nand U11500 (N_11500,N_9542,N_7969);
nand U11501 (N_11501,N_8061,N_6809);
or U11502 (N_11502,N_8117,N_7236);
or U11503 (N_11503,N_7955,N_8376);
nand U11504 (N_11504,N_5553,N_9231);
nor U11505 (N_11505,N_6826,N_8986);
or U11506 (N_11506,N_8828,N_8416);
and U11507 (N_11507,N_9029,N_5070);
nor U11508 (N_11508,N_8444,N_5249);
nor U11509 (N_11509,N_7272,N_7927);
and U11510 (N_11510,N_7106,N_9478);
nand U11511 (N_11511,N_6807,N_8780);
and U11512 (N_11512,N_9024,N_9463);
nor U11513 (N_11513,N_8574,N_7214);
and U11514 (N_11514,N_7672,N_7053);
or U11515 (N_11515,N_5063,N_9021);
and U11516 (N_11516,N_6132,N_6558);
nand U11517 (N_11517,N_9158,N_8194);
nand U11518 (N_11518,N_8984,N_9709);
or U11519 (N_11519,N_8735,N_7844);
nor U11520 (N_11520,N_9695,N_8419);
and U11521 (N_11521,N_5691,N_7077);
and U11522 (N_11522,N_8618,N_6463);
xnor U11523 (N_11523,N_8844,N_9305);
or U11524 (N_11524,N_5190,N_6417);
or U11525 (N_11525,N_8912,N_5870);
nor U11526 (N_11526,N_6506,N_5788);
or U11527 (N_11527,N_5154,N_7027);
nor U11528 (N_11528,N_5696,N_7231);
or U11529 (N_11529,N_8295,N_5672);
nand U11530 (N_11530,N_9778,N_8639);
and U11531 (N_11531,N_7404,N_8730);
xor U11532 (N_11532,N_5375,N_7897);
nand U11533 (N_11533,N_5897,N_8559);
nor U11534 (N_11534,N_8652,N_7390);
nor U11535 (N_11535,N_5784,N_9028);
and U11536 (N_11536,N_7297,N_8579);
nor U11537 (N_11537,N_9534,N_8125);
and U11538 (N_11538,N_8649,N_6116);
nor U11539 (N_11539,N_9577,N_8176);
and U11540 (N_11540,N_7885,N_8474);
or U11541 (N_11541,N_8420,N_5216);
nor U11542 (N_11542,N_7384,N_5926);
nand U11543 (N_11543,N_7309,N_8788);
or U11544 (N_11544,N_8833,N_7800);
or U11545 (N_11545,N_8541,N_7349);
and U11546 (N_11546,N_8990,N_9523);
nand U11547 (N_11547,N_6168,N_9037);
nand U11548 (N_11548,N_9276,N_6265);
xor U11549 (N_11549,N_9460,N_9485);
nor U11550 (N_11550,N_7981,N_7593);
nand U11551 (N_11551,N_7854,N_9987);
nor U11552 (N_11552,N_7992,N_7517);
nor U11553 (N_11553,N_9199,N_7001);
nor U11554 (N_11554,N_6096,N_7304);
or U11555 (N_11555,N_9268,N_5948);
nor U11556 (N_11556,N_6222,N_9573);
or U11557 (N_11557,N_9334,N_9288);
and U11558 (N_11558,N_9865,N_5712);
and U11559 (N_11559,N_7148,N_7388);
or U11560 (N_11560,N_7759,N_8848);
nor U11561 (N_11561,N_5330,N_7600);
xnor U11562 (N_11562,N_8690,N_6472);
nand U11563 (N_11563,N_9637,N_8540);
nand U11564 (N_11564,N_9596,N_7300);
xor U11565 (N_11565,N_5037,N_5438);
and U11566 (N_11566,N_9345,N_5495);
nor U11567 (N_11567,N_7914,N_8993);
nand U11568 (N_11568,N_7833,N_5217);
and U11569 (N_11569,N_9113,N_5269);
nand U11570 (N_11570,N_9487,N_7486);
or U11571 (N_11571,N_9602,N_5372);
nor U11572 (N_11572,N_8370,N_7688);
or U11573 (N_11573,N_5762,N_9952);
and U11574 (N_11574,N_6015,N_9257);
or U11575 (N_11575,N_7318,N_5910);
and U11576 (N_11576,N_5492,N_8292);
nand U11577 (N_11577,N_5486,N_5430);
nand U11578 (N_11578,N_8894,N_7442);
nor U11579 (N_11579,N_6423,N_6888);
and U11580 (N_11580,N_7244,N_7083);
nor U11581 (N_11581,N_7271,N_5020);
or U11582 (N_11582,N_8004,N_5658);
nor U11583 (N_11583,N_5904,N_5676);
nor U11584 (N_11584,N_5002,N_9571);
or U11585 (N_11585,N_5036,N_7460);
nor U11586 (N_11586,N_8762,N_9949);
and U11587 (N_11587,N_8771,N_8470);
nand U11588 (N_11588,N_7997,N_6688);
nand U11589 (N_11589,N_6315,N_5596);
nor U11590 (N_11590,N_7522,N_7785);
and U11591 (N_11591,N_7160,N_5307);
nand U11592 (N_11592,N_8112,N_9104);
nand U11593 (N_11593,N_5517,N_8458);
and U11594 (N_11594,N_9091,N_8027);
nor U11595 (N_11595,N_9025,N_8625);
nor U11596 (N_11596,N_9640,N_8240);
nand U11597 (N_11597,N_8455,N_9781);
or U11598 (N_11598,N_7045,N_5452);
or U11599 (N_11599,N_5173,N_8975);
nand U11600 (N_11600,N_9439,N_8252);
xnor U11601 (N_11601,N_9283,N_8012);
and U11602 (N_11602,N_8058,N_5246);
or U11603 (N_11603,N_8402,N_6686);
and U11604 (N_11604,N_7478,N_5130);
nand U11605 (N_11605,N_6633,N_8111);
and U11606 (N_11606,N_7345,N_6277);
nor U11607 (N_11607,N_7974,N_7026);
nor U11608 (N_11608,N_5090,N_5710);
or U11609 (N_11609,N_7743,N_5689);
nor U11610 (N_11610,N_7725,N_9015);
nand U11611 (N_11611,N_6929,N_9331);
or U11612 (N_11612,N_6052,N_7196);
nor U11613 (N_11613,N_8958,N_5600);
or U11614 (N_11614,N_5725,N_8032);
nand U11615 (N_11615,N_6390,N_7945);
nand U11616 (N_11616,N_7252,N_8967);
and U11617 (N_11617,N_8637,N_5959);
nor U11618 (N_11618,N_6781,N_6887);
or U11619 (N_11619,N_9359,N_9356);
or U11620 (N_11620,N_8505,N_5787);
and U11621 (N_11621,N_9574,N_9835);
nand U11622 (N_11622,N_5338,N_9451);
nand U11623 (N_11623,N_8343,N_9917);
or U11624 (N_11624,N_9896,N_6180);
nor U11625 (N_11625,N_7074,N_8200);
nor U11626 (N_11626,N_6917,N_7789);
nand U11627 (N_11627,N_9467,N_5419);
or U11628 (N_11628,N_9317,N_5703);
xnor U11629 (N_11629,N_7280,N_7289);
or U11630 (N_11630,N_7966,N_5953);
or U11631 (N_11631,N_9300,N_7414);
nor U11632 (N_11632,N_5946,N_9378);
nor U11633 (N_11633,N_8255,N_5849);
or U11634 (N_11634,N_6279,N_6011);
and U11635 (N_11635,N_8720,N_9742);
nand U11636 (N_11636,N_8714,N_8994);
nor U11637 (N_11637,N_8482,N_9638);
or U11638 (N_11638,N_7628,N_7364);
or U11639 (N_11639,N_9691,N_8051);
or U11640 (N_11640,N_8415,N_6665);
nand U11641 (N_11641,N_8645,N_7943);
nor U11642 (N_11642,N_5321,N_6216);
or U11643 (N_11643,N_7587,N_9431);
and U11644 (N_11644,N_6802,N_6074);
or U11645 (N_11645,N_6882,N_7232);
or U11646 (N_11646,N_5911,N_5256);
nor U11647 (N_11647,N_5858,N_6097);
nand U11648 (N_11648,N_9483,N_6876);
nand U11649 (N_11649,N_9873,N_8795);
nor U11650 (N_11650,N_7381,N_7419);
nand U11651 (N_11651,N_5755,N_8172);
and U11652 (N_11652,N_6244,N_9127);
and U11653 (N_11653,N_9956,N_9582);
nor U11654 (N_11654,N_6617,N_5924);
or U11655 (N_11655,N_9282,N_7219);
nor U11656 (N_11656,N_5612,N_8610);
nand U11657 (N_11657,N_9073,N_7876);
nor U11658 (N_11658,N_8575,N_6969);
and U11659 (N_11659,N_9955,N_5282);
nor U11660 (N_11660,N_9251,N_6163);
nor U11661 (N_11661,N_5265,N_5768);
nand U11662 (N_11662,N_8195,N_9822);
or U11663 (N_11663,N_7738,N_8515);
or U11664 (N_11664,N_6664,N_9424);
or U11665 (N_11665,N_8335,N_7251);
nand U11666 (N_11666,N_9085,N_5988);
and U11667 (N_11667,N_9259,N_7024);
and U11668 (N_11668,N_8864,N_5038);
nor U11669 (N_11669,N_8539,N_8459);
nor U11670 (N_11670,N_8857,N_9776);
nor U11671 (N_11671,N_7454,N_6872);
nor U11672 (N_11672,N_8553,N_8654);
nor U11673 (N_11673,N_5566,N_5567);
or U11674 (N_11674,N_7883,N_7333);
nor U11675 (N_11675,N_9958,N_5586);
or U11676 (N_11676,N_5821,N_9470);
and U11677 (N_11677,N_6837,N_5504);
and U11678 (N_11678,N_5445,N_8182);
nor U11679 (N_11679,N_6794,N_8941);
nor U11680 (N_11680,N_6830,N_8110);
nor U11681 (N_11681,N_5276,N_9975);
nor U11682 (N_11682,N_8236,N_8749);
nand U11683 (N_11683,N_9786,N_9165);
nand U11684 (N_11684,N_6338,N_5625);
and U11685 (N_11685,N_6579,N_5402);
nand U11686 (N_11686,N_8825,N_8193);
or U11687 (N_11687,N_9361,N_9748);
nand U11688 (N_11688,N_9772,N_5263);
and U11689 (N_11689,N_7322,N_5651);
or U11690 (N_11690,N_5900,N_5500);
nor U11691 (N_11691,N_5749,N_5774);
or U11692 (N_11692,N_9916,N_6193);
nor U11693 (N_11693,N_9122,N_9551);
nand U11694 (N_11694,N_8196,N_6766);
nand U11695 (N_11695,N_6645,N_9528);
and U11696 (N_11696,N_5200,N_7240);
nand U11697 (N_11697,N_5760,N_6243);
nand U11698 (N_11698,N_9782,N_5791);
and U11699 (N_11699,N_8794,N_7550);
and U11700 (N_11700,N_5232,N_5461);
nor U11701 (N_11701,N_9256,N_6502);
nand U11702 (N_11702,N_5395,N_5404);
nor U11703 (N_11703,N_7508,N_9019);
and U11704 (N_11704,N_5922,N_9806);
or U11705 (N_11705,N_8938,N_6997);
nand U11706 (N_11706,N_6739,N_5212);
and U11707 (N_11707,N_9147,N_7772);
and U11708 (N_11708,N_6455,N_9593);
and U11709 (N_11709,N_8405,N_8981);
nor U11710 (N_11710,N_9307,N_9311);
nand U11711 (N_11711,N_5059,N_9201);
nand U11712 (N_11712,N_8933,N_6636);
nor U11713 (N_11713,N_7156,N_8055);
nand U11714 (N_11714,N_9110,N_7874);
nand U11715 (N_11715,N_7618,N_6461);
and U11716 (N_11716,N_5473,N_6494);
nand U11717 (N_11717,N_8868,N_6054);
or U11718 (N_11718,N_5902,N_7815);
or U11719 (N_11719,N_6947,N_7549);
or U11720 (N_11720,N_5909,N_6662);
or U11721 (N_11721,N_9901,N_5803);
nand U11722 (N_11722,N_5686,N_8578);
xor U11723 (N_11723,N_9419,N_7132);
and U11724 (N_11724,N_6595,N_9941);
nor U11725 (N_11725,N_6607,N_9492);
nand U11726 (N_11726,N_7260,N_7054);
and U11727 (N_11727,N_9871,N_6371);
nand U11728 (N_11728,N_8616,N_7092);
nor U11729 (N_11729,N_8363,N_7595);
xnor U11730 (N_11730,N_5243,N_8413);
or U11731 (N_11731,N_5494,N_6259);
nor U11732 (N_11732,N_5318,N_8830);
nor U11733 (N_11733,N_7861,N_6304);
nand U11734 (N_11734,N_8529,N_6056);
nand U11735 (N_11735,N_5916,N_5351);
and U11736 (N_11736,N_6970,N_9004);
nor U11737 (N_11737,N_8446,N_9576);
and U11738 (N_11738,N_9568,N_7637);
or U11739 (N_11739,N_7325,N_7613);
nand U11740 (N_11740,N_9434,N_5048);
nand U11741 (N_11741,N_9900,N_7695);
and U11742 (N_11742,N_7575,N_8001);
nand U11743 (N_11743,N_9945,N_7655);
xnor U11744 (N_11744,N_7307,N_6769);
and U11745 (N_11745,N_8009,N_5688);
nor U11746 (N_11746,N_9409,N_8243);
or U11747 (N_11747,N_7782,N_8015);
xor U11748 (N_11748,N_8021,N_7717);
or U11749 (N_11749,N_9659,N_7329);
and U11750 (N_11750,N_7155,N_5113);
and U11751 (N_11751,N_7920,N_6983);
or U11752 (N_11752,N_8504,N_7479);
nand U11753 (N_11753,N_5210,N_9832);
and U11754 (N_11754,N_7367,N_5717);
or U11755 (N_11755,N_9818,N_9801);
nor U11756 (N_11756,N_7608,N_5120);
and U11757 (N_11757,N_7237,N_5838);
nor U11758 (N_11758,N_6556,N_5426);
and U11759 (N_11759,N_9677,N_7890);
or U11760 (N_11760,N_7998,N_6637);
and U11761 (N_11761,N_8391,N_8910);
nor U11762 (N_11762,N_8423,N_9447);
and U11763 (N_11763,N_6705,N_8636);
and U11764 (N_11764,N_5976,N_6960);
or U11765 (N_11765,N_8428,N_8978);
xnor U11766 (N_11766,N_5022,N_6678);
and U11767 (N_11767,N_5992,N_8634);
nor U11768 (N_11768,N_5624,N_6268);
or U11769 (N_11769,N_7870,N_7842);
nand U11770 (N_11770,N_5031,N_5193);
and U11771 (N_11771,N_8764,N_8434);
nor U11772 (N_11772,N_8802,N_5754);
or U11773 (N_11773,N_7117,N_5453);
nor U11774 (N_11774,N_6043,N_9079);
or U11775 (N_11775,N_6765,N_8072);
nor U11776 (N_11776,N_8102,N_9740);
or U11777 (N_11777,N_7491,N_7803);
and U11778 (N_11778,N_6999,N_7159);
nand U11779 (N_11779,N_8386,N_5962);
nor U11780 (N_11780,N_5218,N_5362);
nor U11781 (N_11781,N_8475,N_6911);
and U11782 (N_11782,N_6785,N_8162);
nor U11783 (N_11783,N_9788,N_9489);
or U11784 (N_11784,N_8936,N_5280);
and U11785 (N_11785,N_5156,N_8901);
and U11786 (N_11786,N_8737,N_6656);
nor U11787 (N_11787,N_8841,N_9220);
nor U11788 (N_11788,N_6696,N_7150);
nand U11789 (N_11789,N_8874,N_7248);
and U11790 (N_11790,N_9474,N_5520);
nor U11791 (N_11791,N_9630,N_8965);
nand U11792 (N_11792,N_7541,N_9968);
nand U11793 (N_11793,N_8174,N_6658);
or U11794 (N_11794,N_8277,N_7339);
nor U11795 (N_11795,N_9336,N_7276);
or U11796 (N_11796,N_9399,N_5868);
nor U11797 (N_11797,N_6068,N_9738);
nor U11798 (N_11798,N_9929,N_8557);
nand U11799 (N_11799,N_5941,N_5465);
nor U11800 (N_11800,N_6576,N_9156);
and U11801 (N_11801,N_5316,N_5143);
nand U11802 (N_11802,N_5931,N_7556);
and U11803 (N_11803,N_9103,N_9682);
nor U11804 (N_11804,N_5757,N_8008);
or U11805 (N_11805,N_9943,N_9450);
and U11806 (N_11806,N_5713,N_8158);
nand U11807 (N_11807,N_9455,N_7706);
nand U11808 (N_11808,N_6290,N_8398);
nor U11809 (N_11809,N_5106,N_8917);
or U11810 (N_11810,N_5131,N_8603);
nand U11811 (N_11811,N_5446,N_8279);
or U11812 (N_11812,N_9173,N_8734);
or U11813 (N_11813,N_8447,N_9070);
nand U11814 (N_11814,N_6839,N_9233);
nand U11815 (N_11815,N_7202,N_6294);
nor U11816 (N_11816,N_6406,N_8369);
nor U11817 (N_11817,N_9616,N_9584);
nor U11818 (N_11818,N_8155,N_9681);
and U11819 (N_11819,N_9096,N_5403);
nor U11820 (N_11820,N_8721,N_9272);
and U11821 (N_11821,N_6454,N_7832);
nand U11822 (N_11822,N_9965,N_7402);
or U11823 (N_11823,N_8000,N_6214);
or U11824 (N_11824,N_7818,N_8120);
nand U11825 (N_11825,N_5824,N_6971);
nand U11826 (N_11826,N_7700,N_6740);
nand U11827 (N_11827,N_5839,N_7173);
or U11828 (N_11828,N_6123,N_9329);
nor U11829 (N_11829,N_6086,N_5144);
nand U11830 (N_11830,N_7149,N_8472);
nand U11831 (N_11831,N_7978,N_8237);
nor U11832 (N_11832,N_9471,N_8566);
nor U11833 (N_11833,N_6167,N_9874);
nor U11834 (N_11834,N_7194,N_5779);
or U11835 (N_11835,N_8670,N_5259);
or U11836 (N_11836,N_9093,N_7669);
and U11837 (N_11837,N_9417,N_7073);
xnor U11838 (N_11838,N_9397,N_6144);
or U11839 (N_11839,N_9539,N_7378);
and U11840 (N_11840,N_6317,N_6632);
nor U11841 (N_11841,N_7327,N_7020);
and U11842 (N_11842,N_7826,N_6083);
nor U11843 (N_11843,N_7395,N_5995);
and U11844 (N_11844,N_8813,N_7737);
nor U11845 (N_11845,N_5127,N_8976);
nor U11846 (N_11846,N_9023,N_7835);
nor U11847 (N_11847,N_8662,N_6753);
and U11848 (N_11848,N_9790,N_5563);
and U11849 (N_11849,N_7907,N_8276);
or U11850 (N_11850,N_6323,N_7740);
or U11851 (N_11851,N_7382,N_7095);
nor U11852 (N_11852,N_7266,N_7561);
nand U11853 (N_11853,N_5397,N_7984);
and U11854 (N_11854,N_7213,N_5737);
nand U11855 (N_11855,N_9225,N_8923);
nor U11856 (N_11856,N_6352,N_7134);
or U11857 (N_11857,N_5019,N_8646);
nor U11858 (N_11858,N_6354,N_5906);
or U11859 (N_11859,N_7909,N_5898);
and U11860 (N_11860,N_5594,N_7462);
and U11861 (N_11861,N_6048,N_9989);
or U11862 (N_11862,N_9177,N_9838);
or U11863 (N_11863,N_8175,N_9589);
nand U11864 (N_11864,N_7806,N_6544);
nand U11865 (N_11865,N_5119,N_9556);
nand U11866 (N_11866,N_9031,N_6206);
nor U11867 (N_11867,N_6539,N_6988);
and U11868 (N_11868,N_9517,N_9586);
and U11869 (N_11869,N_5846,N_8907);
or U11870 (N_11870,N_8883,N_8711);
and U11871 (N_11871,N_5464,N_6191);
nor U11872 (N_11872,N_7500,N_7153);
or U11873 (N_11873,N_7177,N_9052);
nand U11874 (N_11874,N_9294,N_8315);
or U11875 (N_11875,N_9166,N_6189);
or U11876 (N_11876,N_5153,N_6811);
nor U11877 (N_11877,N_8449,N_6234);
nor U11878 (N_11878,N_9043,N_6788);
nor U11879 (N_11879,N_8589,N_7831);
nand U11880 (N_11880,N_5000,N_6360);
and U11881 (N_11881,N_8925,N_7205);
nor U11882 (N_11882,N_5058,N_7440);
or U11883 (N_11883,N_6479,N_8109);
nand U11884 (N_11884,N_8059,N_9711);
nor U11885 (N_11885,N_7654,N_5913);
or U11886 (N_11886,N_7944,N_6964);
xnor U11887 (N_11887,N_8785,N_6179);
or U11888 (N_11888,N_9406,N_5272);
nand U11889 (N_11889,N_5382,N_6951);
or U11890 (N_11890,N_9010,N_9286);
xor U11891 (N_11891,N_7211,N_7863);
and U11892 (N_11892,N_7093,N_5822);
nand U11893 (N_11893,N_6608,N_7985);
nor U11894 (N_11894,N_5341,N_5552);
or U11895 (N_11895,N_7788,N_7494);
and U11896 (N_11896,N_7161,N_7965);
and U11897 (N_11897,N_5575,N_5011);
and U11898 (N_11898,N_9343,N_7372);
nor U11899 (N_11899,N_6582,N_7193);
nor U11900 (N_11900,N_8995,N_7021);
or U11901 (N_11901,N_7673,N_6653);
and U11902 (N_11902,N_7756,N_6176);
nor U11903 (N_11903,N_8352,N_7729);
and U11904 (N_11904,N_5647,N_8319);
nor U11905 (N_11905,N_8805,N_8414);
and U11906 (N_11906,N_6481,N_7746);
and U11907 (N_11907,N_8943,N_8839);
and U11908 (N_11908,N_8863,N_7424);
nor U11909 (N_11909,N_9854,N_7524);
nand U11910 (N_11910,N_5740,N_9006);
or U11911 (N_11911,N_6714,N_9009);
nor U11912 (N_11912,N_8382,N_9222);
nand U11913 (N_11913,N_5507,N_5199);
or U11914 (N_11914,N_8399,N_5385);
nor U11915 (N_11915,N_7102,N_9360);
nand U11916 (N_11916,N_5511,N_8178);
nand U11917 (N_11917,N_6393,N_9087);
nand U11918 (N_11918,N_7925,N_7456);
nor U11919 (N_11919,N_8336,N_6581);
and U11920 (N_11920,N_7450,N_6419);
or U11921 (N_11921,N_7906,N_8554);
nand U11922 (N_11922,N_6230,N_6306);
xnor U11923 (N_11923,N_9575,N_6994);
or U11924 (N_11924,N_7180,N_8375);
nor U11925 (N_11925,N_7816,N_6508);
and U11926 (N_11926,N_5815,N_5907);
nor U11927 (N_11927,N_7758,N_5893);
nor U11928 (N_11928,N_8217,N_5577);
or U11929 (N_11929,N_9885,N_5772);
nand U11930 (N_11930,N_5771,N_9252);
nand U11931 (N_11931,N_6212,N_5764);
or U11932 (N_11932,N_5745,N_6599);
and U11933 (N_11933,N_7871,N_5240);
nand U11934 (N_11934,N_8042,N_5536);
and U11935 (N_11935,N_6300,N_8298);
nor U11936 (N_11936,N_6524,N_7504);
or U11937 (N_11937,N_5546,N_7256);
and U11938 (N_11938,N_8062,N_5042);
or U11939 (N_11939,N_6378,N_9812);
and U11940 (N_11940,N_5615,N_9182);
nand U11941 (N_11941,N_7899,N_9515);
or U11942 (N_11942,N_8911,N_8057);
and U11943 (N_11943,N_9597,N_7210);
nor U11944 (N_11944,N_8836,N_6131);
or U11945 (N_11945,N_8877,N_5512);
nor U11946 (N_11946,N_9824,N_6547);
and U11947 (N_11947,N_6978,N_7287);
xnor U11948 (N_11948,N_6477,N_6701);
nor U11949 (N_11949,N_5303,N_6598);
and U11950 (N_11950,N_9067,N_5828);
or U11951 (N_11951,N_7823,N_9221);
and U11952 (N_11952,N_7910,N_5644);
nor U11953 (N_11953,N_8325,N_5750);
and U11954 (N_11954,N_7239,N_6192);
nand U11955 (N_11955,N_8153,N_9045);
nand U11956 (N_11956,N_5413,N_5673);
nor U11957 (N_11957,N_7684,N_6359);
nor U11958 (N_11958,N_5797,N_8580);
and U11959 (N_11959,N_7152,N_5979);
nand U11960 (N_11960,N_7290,N_7259);
nand U11961 (N_11961,N_9983,N_8074);
and U11962 (N_11962,N_8760,N_8872);
nor U11963 (N_11963,N_6625,N_7697);
nor U11964 (N_11964,N_6002,N_9521);
nor U11965 (N_11965,N_5538,N_6170);
nor U11966 (N_11966,N_5392,N_6254);
nand U11967 (N_11967,N_9271,N_6181);
or U11968 (N_11968,N_8988,N_7432);
and U11969 (N_11969,N_6370,N_9481);
and U11970 (N_11970,N_8206,N_5289);
nand U11971 (N_11971,N_5798,N_7960);
and U11972 (N_11972,N_9042,N_7993);
or U11973 (N_11973,N_9622,N_5932);
or U11974 (N_11974,N_9522,N_5223);
nor U11975 (N_11975,N_7262,N_6325);
and U11976 (N_11976,N_6267,N_8122);
and U11977 (N_11977,N_6568,N_7415);
nand U11978 (N_11978,N_8642,N_7880);
or U11979 (N_11979,N_5687,N_6401);
nor U11980 (N_11980,N_8664,N_6467);
and U11981 (N_11981,N_5967,N_7167);
nor U11982 (N_11982,N_9708,N_8823);
and U11983 (N_11983,N_8588,N_7588);
nand U11984 (N_11984,N_5111,N_7716);
nor U11985 (N_11985,N_6914,N_7796);
or U11986 (N_11986,N_6799,N_8213);
or U11987 (N_11987,N_9032,N_5960);
or U11988 (N_11988,N_9634,N_8806);
xor U11989 (N_11989,N_6943,N_7601);
nor U11990 (N_11990,N_7365,N_7900);
or U11991 (N_11991,N_5867,N_6060);
nand U11992 (N_11992,N_8170,N_8702);
nand U11993 (N_11993,N_9385,N_7865);
nor U11994 (N_11994,N_5937,N_5777);
and U11995 (N_11995,N_5621,N_5693);
nand U11996 (N_11996,N_7438,N_6860);
and U11997 (N_11997,N_5537,N_5660);
and U11998 (N_11998,N_6864,N_8982);
nand U11999 (N_11999,N_7076,N_5526);
and U12000 (N_12000,N_7488,N_7713);
and U12001 (N_12001,N_6245,N_6124);
or U12002 (N_12002,N_7294,N_5046);
or U12003 (N_12003,N_8181,N_7018);
nand U12004 (N_12004,N_5358,N_5794);
nand U12005 (N_12005,N_5637,N_8192);
or U12006 (N_12006,N_5152,N_9441);
nor U12007 (N_12007,N_6242,N_5164);
or U12008 (N_12008,N_5389,N_9390);
or U12009 (N_12009,N_9998,N_5942);
nand U12010 (N_12010,N_7879,N_9583);
or U12011 (N_12011,N_9974,N_5861);
and U12012 (N_12012,N_5026,N_8809);
and U12013 (N_12013,N_6892,N_5139);
nor U12014 (N_12014,N_9858,N_9696);
nor U12015 (N_12015,N_9514,N_9429);
or U12016 (N_12016,N_8922,N_8782);
xor U12017 (N_12017,N_8680,N_7032);
and U12018 (N_12018,N_5041,N_7277);
and U12019 (N_12019,N_5732,N_7291);
or U12020 (N_12020,N_7480,N_9172);
nor U12021 (N_12021,N_8895,N_7407);
or U12022 (N_12022,N_5544,N_8073);
and U12023 (N_12023,N_5929,N_9543);
nor U12024 (N_12024,N_5970,N_8784);
nand U12025 (N_12025,N_5633,N_7755);
nor U12026 (N_12026,N_5267,N_9218);
or U12027 (N_12027,N_9567,N_5998);
nor U12028 (N_12028,N_7661,N_6773);
or U12029 (N_12029,N_6519,N_8971);
or U12030 (N_12030,N_7411,N_7570);
or U12031 (N_12031,N_9683,N_9267);
or U12032 (N_12032,N_6979,N_9333);
nor U12033 (N_12033,N_9654,N_6429);
or U12034 (N_12034,N_6855,N_8280);
nor U12035 (N_12035,N_9579,N_5328);
and U12036 (N_12036,N_8124,N_9181);
or U12037 (N_12037,N_5319,N_8365);
and U12038 (N_12038,N_6333,N_9448);
or U12039 (N_12039,N_7394,N_7643);
or U12040 (N_12040,N_9936,N_9298);
nor U12041 (N_12041,N_9187,N_5475);
nand U12042 (N_12042,N_6906,N_5171);
or U12043 (N_12043,N_5065,N_7836);
or U12044 (N_12044,N_9756,N_8445);
or U12045 (N_12045,N_9819,N_7778);
nand U12046 (N_12046,N_9145,N_7052);
or U12047 (N_12047,N_6207,N_5606);
nor U12048 (N_12048,N_9810,N_6703);
nand U12049 (N_12049,N_5035,N_7663);
nor U12050 (N_12050,N_9315,N_7689);
and U12051 (N_12051,N_7513,N_8310);
and U12052 (N_12052,N_9913,N_8867);
nor U12053 (N_12053,N_9557,N_5773);
and U12054 (N_12054,N_7775,N_7292);
and U12055 (N_12055,N_5665,N_6468);
and U12056 (N_12056,N_8977,N_8601);
and U12057 (N_12057,N_5820,N_8003);
nor U12058 (N_12058,N_8060,N_9403);
and U12059 (N_12059,N_5043,N_6160);
nor U12060 (N_12060,N_9580,N_7458);
nand U12061 (N_12061,N_6532,N_6375);
nor U12062 (N_12062,N_9620,N_8294);
and U12063 (N_12063,N_8493,N_8827);
xnor U12064 (N_12064,N_5848,N_9633);
nor U12065 (N_12065,N_9208,N_5083);
nor U12066 (N_12066,N_9068,N_8451);
and U12067 (N_12067,N_7731,N_5940);
nor U12068 (N_12068,N_8615,N_9732);
or U12069 (N_12069,N_8115,N_8896);
nor U12070 (N_12070,N_5471,N_9401);
and U12071 (N_12071,N_9153,N_9935);
or U12072 (N_12072,N_5301,N_5417);
nand U12073 (N_12073,N_7157,N_9143);
nand U12074 (N_12074,N_8223,N_6926);
nor U12075 (N_12075,N_7898,N_5584);
nor U12076 (N_12076,N_5204,N_7581);
and U12077 (N_12077,N_7143,N_5763);
and U12078 (N_12078,N_9062,N_5947);
nand U12079 (N_12079,N_6612,N_8316);
or U12080 (N_12080,N_7519,N_7604);
and U12081 (N_12081,N_5837,N_6611);
nor U12082 (N_12082,N_7691,N_9950);
nand U12083 (N_12083,N_6682,N_6650);
nand U12084 (N_12084,N_5347,N_7475);
or U12085 (N_12085,N_9836,N_6663);
nor U12086 (N_12086,N_6711,N_9735);
nand U12087 (N_12087,N_8768,N_9504);
nor U12088 (N_12088,N_7585,N_5780);
and U12089 (N_12089,N_9692,N_7457);
nand U12090 (N_12090,N_7972,N_9961);
xor U12091 (N_12091,N_8942,N_5189);
nand U12092 (N_12092,N_5903,N_5312);
or U12093 (N_12093,N_8904,N_9899);
and U12094 (N_12094,N_8594,N_8066);
or U12095 (N_12095,N_5943,N_6541);
and U12096 (N_12096,N_6535,N_8853);
nand U12097 (N_12097,N_6555,N_8678);
nor U12098 (N_12098,N_5908,N_5877);
or U12099 (N_12099,N_7950,N_8492);
nor U12100 (N_12100,N_8509,N_9951);
nor U12101 (N_12101,N_9132,N_9020);
nand U12102 (N_12102,N_5726,N_7172);
nor U12103 (N_12103,N_8921,N_8267);
nand U12104 (N_12104,N_8757,N_5296);
and U12105 (N_12105,N_8685,N_8222);
nor U12106 (N_12106,N_7041,N_5701);
nand U12107 (N_12107,N_5368,N_7511);
or U12108 (N_12108,N_6513,N_7830);
nand U12109 (N_12109,N_7967,N_9499);
nor U12110 (N_12110,N_5744,N_8724);
nor U12111 (N_12111,N_9641,N_6649);
or U12112 (N_12112,N_9427,N_7401);
nand U12113 (N_12113,N_7118,N_9174);
and U12114 (N_12114,N_5578,N_8477);
nor U12115 (N_12115,N_9496,N_9142);
and U12116 (N_12116,N_9804,N_5377);
nand U12117 (N_12117,N_9548,N_6346);
nor U12118 (N_12118,N_7739,N_6698);
and U12119 (N_12119,N_5141,N_5254);
or U12120 (N_12120,N_6031,N_7646);
nor U12121 (N_12121,N_5607,N_9078);
or U12122 (N_12122,N_6934,N_9097);
nand U12123 (N_12123,N_6500,N_8879);
or U12124 (N_12124,N_5957,N_6692);
nor U12125 (N_12125,N_6349,N_6538);
nor U12126 (N_12126,N_7047,N_5441);
nand U12127 (N_12127,N_8537,N_9657);
or U12128 (N_12128,N_8614,N_8489);
and U12129 (N_12129,N_9760,N_6303);
or U12130 (N_12130,N_5137,N_8039);
nand U12131 (N_12131,N_8705,N_7069);
nor U12132 (N_12132,N_8198,N_9762);
and U12133 (N_12133,N_5016,N_9554);
and U12134 (N_12134,N_6879,N_6790);
nor U12135 (N_12135,N_6549,N_9734);
and U12136 (N_12136,N_8510,N_7692);
or U12137 (N_12137,N_7736,N_9232);
nand U12138 (N_12138,N_9604,N_7227);
nand U12139 (N_12139,N_7896,N_8991);
or U12140 (N_12140,N_7332,N_7428);
or U12141 (N_12141,N_8908,N_7165);
and U12142 (N_12142,N_5102,N_7811);
and U12143 (N_12143,N_7525,N_7470);
and U12144 (N_12144,N_6114,N_8082);
and U12145 (N_12145,N_7386,N_5496);
nand U12146 (N_12146,N_9644,N_5277);
nand U12147 (N_12147,N_7911,N_8043);
or U12148 (N_12148,N_6129,N_7621);
nor U12149 (N_12149,N_7207,N_9698);
xnor U12150 (N_12150,N_5158,N_7181);
and U12151 (N_12151,N_5266,N_5214);
nor U12152 (N_12152,N_7223,N_8851);
or U12153 (N_12153,N_5767,N_6710);
and U12154 (N_12154,N_6051,N_7592);
and U12155 (N_12155,N_6869,N_6831);
nand U12156 (N_12156,N_8123,N_6818);
or U12157 (N_12157,N_5541,N_5151);
and U12158 (N_12158,N_7749,N_5748);
nand U12159 (N_12159,N_8234,N_9629);
nor U12160 (N_12160,N_8528,N_6437);
and U12161 (N_12161,N_5183,N_9120);
nor U12162 (N_12162,N_8523,N_5708);
or U12163 (N_12163,N_8954,N_8946);
nand U12164 (N_12164,N_9432,N_7779);
nand U12165 (N_12165,N_5731,N_9796);
or U12166 (N_12166,N_8797,N_5490);
and U12167 (N_12167,N_9934,N_6726);
nor U12168 (N_12168,N_8882,N_5585);
nand U12169 (N_12169,N_8534,N_5359);
nand U12170 (N_12170,N_6208,N_9529);
nor U12171 (N_12171,N_9944,N_5311);
and U12172 (N_12172,N_7869,N_8577);
and U12173 (N_12173,N_6936,N_5866);
nand U12174 (N_12174,N_9609,N_6261);
or U12175 (N_12175,N_8332,N_9555);
or U12176 (N_12176,N_6545,N_7612);
and U12177 (N_12177,N_7125,N_5999);
or U12178 (N_12178,N_6269,N_7686);
and U12179 (N_12179,N_5068,N_9141);
nand U12180 (N_12180,N_8606,N_5843);
and U12181 (N_12181,N_5513,N_9993);
or U12182 (N_12182,N_7441,N_9229);
or U12183 (N_12183,N_5997,N_6967);
nand U12184 (N_12184,N_7791,N_8929);
or U12185 (N_12185,N_7792,N_7929);
or U12186 (N_12186,N_8291,N_5449);
or U12187 (N_12187,N_6900,N_8189);
xor U12188 (N_12188,N_5663,N_9313);
and U12189 (N_12189,N_8190,N_8641);
nand U12190 (N_12190,N_6594,N_7133);
or U12191 (N_12191,N_8281,N_5291);
nand U12192 (N_12192,N_7626,N_5077);
and U12193 (N_12193,N_5895,N_6720);
or U12194 (N_12194,N_8648,N_6301);
or U12195 (N_12195,N_5734,N_8892);
nor U12196 (N_12196,N_7752,N_8792);
or U12197 (N_12197,N_7376,N_9391);
or U12198 (N_12198,N_5095,N_5558);
nor U12199 (N_12199,N_8745,N_7507);
or U12200 (N_12200,N_9668,N_5231);
or U12201 (N_12201,N_9425,N_5547);
nor U12202 (N_12202,N_5221,N_5211);
nor U12203 (N_12203,N_9270,N_8875);
or U12204 (N_12204,N_7771,N_5175);
and U12205 (N_12205,N_5365,N_7090);
nand U12206 (N_12206,N_7956,N_7797);
nand U12207 (N_12207,N_5170,N_8514);
nand U12208 (N_12208,N_7168,N_5994);
nor U12209 (N_12209,N_5147,N_6082);
nor U12210 (N_12210,N_8752,N_7066);
and U12211 (N_12211,N_6016,N_9100);
nor U12212 (N_12212,N_5873,N_9369);
and U12213 (N_12213,N_5643,N_8266);
nor U12214 (N_12214,N_7938,N_9077);
and U12215 (N_12215,N_9497,N_5990);
and U12216 (N_12216,N_5092,N_6281);
nor U12217 (N_12217,N_5807,N_9744);
xor U12218 (N_12218,N_6530,N_7615);
or U12219 (N_12219,N_6684,N_9116);
nand U12220 (N_12220,N_6814,N_9894);
and U12221 (N_12221,N_6445,N_6017);
nand U12222 (N_12222,N_8426,N_7668);
nor U12223 (N_12223,N_6949,N_5129);
nor U12224 (N_12224,N_7658,N_9306);
and U12225 (N_12225,N_9046,N_8354);
nor U12226 (N_12226,N_6330,N_5354);
xor U12227 (N_12227,N_6529,N_8657);
or U12228 (N_12228,N_7493,N_6889);
or U12229 (N_12229,N_6748,N_6596);
nor U12230 (N_12230,N_7850,N_7014);
nand U12231 (N_12231,N_5871,N_7447);
and U12232 (N_12232,N_8479,N_9074);
and U12233 (N_12233,N_5180,N_5013);
or U12234 (N_12234,N_8550,N_5066);
nor U12235 (N_12235,N_6600,N_8141);
nand U12236 (N_12236,N_7317,N_7410);
or U12237 (N_12237,N_8959,N_8168);
and U12238 (N_12238,N_7777,N_7754);
nand U12239 (N_12239,N_6883,N_8587);
nand U12240 (N_12240,N_5064,N_7062);
nor U12241 (N_12241,N_7474,N_7636);
nand U12242 (N_12242,N_5023,N_7465);
nor U12243 (N_12243,N_6275,N_9340);
and U12244 (N_12244,N_8105,N_7449);
nor U12245 (N_12245,N_9262,N_8650);
or U12246 (N_12246,N_7385,N_8581);
nor U12247 (N_12247,N_9179,N_6280);
nand U12248 (N_12248,N_9922,N_6273);
nand U12249 (N_12249,N_6685,N_9875);
or U12250 (N_12250,N_7940,N_8334);
and U12251 (N_12251,N_8913,N_5674);
or U12252 (N_12252,N_5542,N_9435);
and U12253 (N_12253,N_6708,N_8739);
and U12254 (N_12254,N_7473,N_9063);
and U12255 (N_12255,N_6981,N_9446);
xor U12256 (N_12256,N_7530,N_5194);
or U12257 (N_12257,N_6402,N_7257);
or U12258 (N_12258,N_9430,N_7357);
and U12259 (N_12259,N_9561,N_7963);
nor U12260 (N_12260,N_8849,N_7753);
and U12261 (N_12261,N_9624,N_6125);
nand U12262 (N_12262,N_6505,N_7336);
or U12263 (N_12263,N_6905,N_8179);
and U12264 (N_12264,N_6909,N_7667);
or U12265 (N_12265,N_6928,N_7849);
or U12266 (N_12266,N_6691,N_5040);
nand U12267 (N_12267,N_9687,N_6918);
or U12268 (N_12268,N_7543,N_7380);
nor U12269 (N_12269,N_8861,N_6157);
or U12270 (N_12270,N_7633,N_7163);
or U12271 (N_12271,N_5376,N_6434);
or U12272 (N_12272,N_7770,N_6249);
xor U12273 (N_12273,N_6903,N_7535);
nor U12274 (N_12274,N_5315,N_9260);
or U12275 (N_12275,N_9438,N_7768);
or U12276 (N_12276,N_7534,N_6302);
nand U12277 (N_12277,N_6342,N_5285);
and U12278 (N_12278,N_5086,N_5481);
nand U12279 (N_12279,N_7000,N_6857);
or U12280 (N_12280,N_7467,N_6000);
or U12281 (N_12281,N_7358,N_8647);
and U12282 (N_12282,N_7434,N_7164);
nor U12283 (N_12283,N_6165,N_8247);
and U12284 (N_12284,N_9030,N_7477);
nor U12285 (N_12285,N_8007,N_5274);
nand U12286 (N_12286,N_5860,N_5963);
nor U12287 (N_12287,N_8201,N_6697);
and U12288 (N_12288,N_9265,N_9675);
nand U12289 (N_12289,N_8838,N_5109);
nand U12290 (N_12290,N_8969,N_5840);
nand U12291 (N_12291,N_5325,N_9979);
nor U12292 (N_12292,N_6151,N_9351);
and U12293 (N_12293,N_5901,N_6343);
or U12294 (N_12294,N_7694,N_7154);
and U12295 (N_12295,N_8815,N_7463);
nand U12296 (N_12296,N_8511,N_9701);
nor U12297 (N_12297,N_8996,N_8611);
xor U12298 (N_12298,N_8264,N_6470);
and U12299 (N_12299,N_9850,N_6127);
or U12300 (N_12300,N_5284,N_7935);
nor U12301 (N_12301,N_9771,N_5185);
and U12302 (N_12302,N_9948,N_9278);
nor U12303 (N_12303,N_8924,N_7296);
and U12304 (N_12304,N_6307,N_5863);
nor U12305 (N_12305,N_6363,N_7311);
nand U12306 (N_12306,N_9627,N_9977);
nand U12307 (N_12307,N_8759,N_9466);
or U12308 (N_12308,N_8987,N_5157);
nand U12309 (N_12309,N_9834,N_9988);
or U12310 (N_12310,N_7923,N_9115);
nor U12311 (N_12311,N_8790,N_7423);
nand U12312 (N_12312,N_5220,N_9601);
nor U12313 (N_12313,N_8592,N_6778);
nor U12314 (N_12314,N_6396,N_9421);
and U12315 (N_12315,N_8783,N_6367);
nand U12316 (N_12316,N_9308,N_6013);
or U12317 (N_12317,N_9443,N_6761);
or U12318 (N_12318,N_7101,N_9195);
or U12319 (N_12319,N_6933,N_9612);
nand U12320 (N_12320,N_7540,N_5440);
nor U12321 (N_12321,N_9098,N_5842);
nand U12322 (N_12322,N_8707,N_6722);
and U12323 (N_12323,N_9240,N_6628);
nor U12324 (N_12324,N_5305,N_5428);
nor U12325 (N_12325,N_9454,N_7551);
and U12326 (N_12326,N_6427,N_9083);
or U12327 (N_12327,N_8084,N_5550);
or U12328 (N_12328,N_9867,N_6058);
or U12329 (N_12329,N_6410,N_9815);
nand U12330 (N_12330,N_5884,N_9495);
nand U12331 (N_12331,N_5835,N_9458);
nor U12332 (N_12332,N_9970,N_6462);
or U12333 (N_12333,N_7976,N_9452);
nand U12334 (N_12334,N_9114,N_9925);
nor U12335 (N_12335,N_9444,N_9176);
and U12336 (N_12336,N_7784,N_6289);
nor U12337 (N_12337,N_6252,N_7162);
and U12338 (N_12338,N_9138,N_6721);
or U12339 (N_12339,N_9623,N_8437);
nand U12340 (N_12340,N_7328,N_6987);
nand U12341 (N_12341,N_8777,N_6420);
xnor U12342 (N_12342,N_6895,N_6344);
nor U12343 (N_12343,N_9102,N_9041);
nand U12344 (N_12344,N_7912,N_5197);
nand U12345 (N_12345,N_6223,N_6915);
and U12346 (N_12346,N_6551,N_7930);
and U12347 (N_12347,N_7915,N_5857);
nor U12348 (N_12348,N_6431,N_7174);
or U12349 (N_12349,N_5003,N_6992);
and U12350 (N_12350,N_8209,N_5118);
nand U12351 (N_12351,N_7483,N_6503);
nor U12352 (N_12352,N_9758,N_6674);
or U12353 (N_12353,N_6877,N_8250);
and U12354 (N_12354,N_7708,N_7882);
nand U12355 (N_12355,N_7023,N_7566);
or U12356 (N_12356,N_5622,N_9055);
nor U12357 (N_12357,N_9566,N_9162);
nor U12358 (N_12358,N_5088,N_7812);
or U12359 (N_12359,N_6526,N_6777);
or U12360 (N_12360,N_7855,N_7496);
and U12361 (N_12361,N_9095,N_7747);
nand U12362 (N_12362,N_8893,N_6537);
and U12363 (N_12363,N_6042,N_8435);
or U12364 (N_12364,N_5521,N_9713);
nand U12365 (N_12365,N_6202,N_6661);
nor U12366 (N_12366,N_8576,N_9477);
or U12367 (N_12367,N_6795,N_6006);
nand U12368 (N_12368,N_9189,N_7055);
nand U12369 (N_12369,N_8621,N_9051);
nor U12370 (N_12370,N_5167,N_7712);
nor U12371 (N_12371,N_5017,N_9678);
nand U12372 (N_12372,N_5964,N_5207);
nand U12373 (N_12373,N_7572,N_9371);
nand U12374 (N_12374,N_5800,N_7893);
nor U12375 (N_12375,N_9188,N_8309);
and U12376 (N_12376,N_9808,N_5051);
or U12377 (N_12377,N_9846,N_6670);
nor U12378 (N_12378,N_9135,N_5400);
or U12379 (N_12379,N_7665,N_8704);
nor U12380 (N_12380,N_9927,N_8275);
nand U12381 (N_12381,N_5480,N_5378);
or U12382 (N_12382,N_5977,N_7644);
or U12383 (N_12383,N_9099,N_6554);
nor U12384 (N_12384,N_8810,N_9126);
and U12385 (N_12385,N_5756,N_8297);
nand U12386 (N_12386,N_8104,N_7975);
nand U12387 (N_12387,N_8607,N_6241);
nor U12388 (N_12388,N_6522,N_7808);
nand U12389 (N_12389,N_6109,N_8856);
nor U12390 (N_12390,N_8772,N_9844);
or U12391 (N_12391,N_5227,N_8035);
or U12392 (N_12392,N_9388,N_7856);
and U12393 (N_12393,N_6870,N_7574);
nand U12394 (N_12394,N_6856,N_7203);
nand U12395 (N_12395,N_8224,N_5826);
nand U12396 (N_12396,N_9795,N_7429);
xnor U12397 (N_12397,N_5488,N_6194);
nor U12398 (N_12398,N_6283,N_5684);
nand U12399 (N_12399,N_6019,N_9412);
nor U12400 (N_12400,N_7111,N_7847);
nand U12401 (N_12401,N_7335,N_9861);
and U12402 (N_12402,N_5300,N_7528);
nor U12403 (N_12403,N_5555,N_9518);
nor U12404 (N_12404,N_8303,N_7634);
nor U12405 (N_12405,N_6478,N_6574);
or U12406 (N_12406,N_5604,N_9264);
nor U12407 (N_12407,N_6732,N_6240);
nand U12408 (N_12408,N_6139,N_5685);
nand U12409 (N_12409,N_7578,N_5510);
nand U12410 (N_12410,N_9255,N_7225);
and U12411 (N_12411,N_6247,N_6493);
nand U12412 (N_12412,N_5652,N_8751);
nand U12413 (N_12413,N_8811,N_6627);
nor U12414 (N_12414,N_9667,N_8358);
or U12415 (N_12415,N_5966,N_5580);
nor U12416 (N_12416,N_9933,N_6958);
nor U12417 (N_12417,N_5072,N_5273);
and U12418 (N_12418,N_6854,N_7645);
or U12419 (N_12419,N_7302,N_8348);
nand U12420 (N_12420,N_9377,N_9724);
nand U12421 (N_12421,N_5181,N_6552);
nand U12422 (N_12422,N_5499,N_7212);
or U12423 (N_12423,N_9700,N_7186);
and U12424 (N_12424,N_7718,N_8360);
and U12425 (N_12425,N_8617,N_9292);
xor U12426 (N_12426,N_8948,N_7080);
or U12427 (N_12427,N_7008,N_8869);
and U12428 (N_12428,N_6311,N_5912);
and U12429 (N_12429,N_9012,N_9137);
and U12430 (N_12430,N_9852,N_8937);
nand U12431 (N_12431,N_8713,N_8915);
nor U12432 (N_12432,N_6436,N_8972);
or U12433 (N_12433,N_6651,N_7079);
and U12434 (N_12434,N_9763,N_6203);
nor U12435 (N_12435,N_7389,N_8010);
nand U12436 (N_12436,N_7444,N_9730);
or U12437 (N_12437,N_9972,N_8187);
and U12438 (N_12438,N_9607,N_9883);
nor U12439 (N_12439,N_9747,N_6171);
or U12440 (N_12440,N_7846,N_7852);
nand U12441 (N_12441,N_7917,N_7094);
and U12442 (N_12442,N_9323,N_8020);
nor U12443 (N_12443,N_5067,N_8101);
or U12444 (N_12444,N_7323,N_9959);
nand U12445 (N_12445,N_9293,N_8526);
and U12446 (N_12446,N_9903,N_6816);
and U12447 (N_12447,N_6377,N_5348);
and U12448 (N_12448,N_7116,N_8506);
nand U12449 (N_12449,N_8801,N_8088);
nand U12450 (N_12450,N_5433,N_6145);
nor U12451 (N_12451,N_5021,N_6871);
and U12452 (N_12452,N_5709,N_9680);
or U12453 (N_12453,N_5915,N_8070);
and U12454 (N_12454,N_9562,N_6821);
or U12455 (N_12455,N_6175,N_6484);
or U12456 (N_12456,N_5257,N_5864);
nand U12457 (N_12457,N_5945,N_5808);
and U12458 (N_12458,N_6091,N_9519);
or U12459 (N_12459,N_7794,N_6623);
nor U12460 (N_12460,N_8044,N_8694);
nor U12461 (N_12461,N_5918,N_9119);
or U12462 (N_12462,N_6021,N_5579);
or U12463 (N_12463,N_5293,N_5081);
or U12464 (N_12464,N_9799,N_6332);
nand U12465 (N_12465,N_5244,N_6438);
nor U12466 (N_12466,N_8085,N_5352);
nand U12467 (N_12467,N_8527,N_5938);
or U12468 (N_12468,N_6228,N_6910);
nor U12469 (N_12469,N_7805,N_6313);
or U12470 (N_12470,N_5532,N_9465);
nand U12471 (N_12471,N_5659,N_8256);
nor U12472 (N_12472,N_9803,N_6184);
nor U12473 (N_12473,N_9710,N_9613);
or U12474 (N_12474,N_5367,N_5716);
or U12475 (N_12475,N_6683,N_6998);
or U12476 (N_12476,N_8775,N_9332);
and U12477 (N_12477,N_7468,N_5611);
and U12478 (N_12478,N_8411,N_9244);
nor U12479 (N_12479,N_8738,N_7229);
nor U12480 (N_12480,N_7137,N_9716);
nor U12481 (N_12481,N_9705,N_5363);
nor U12482 (N_12482,N_6931,N_6142);
and U12483 (N_12483,N_8902,N_9381);
nand U12484 (N_12484,N_9924,N_7769);
and U12485 (N_12485,N_5865,N_8028);
nand U12486 (N_12486,N_8417,N_6946);
nand U12487 (N_12487,N_5132,N_5103);
and U12488 (N_12488,N_8829,N_6009);
nand U12489 (N_12489,N_6369,N_6620);
nor U12490 (N_12490,N_8803,N_6712);
and U12491 (N_12491,N_6863,N_9155);
nand U12492 (N_12492,N_9148,N_5370);
or U12493 (N_12493,N_8558,N_9636);
nand U12494 (N_12494,N_6859,N_6147);
or U12495 (N_12495,N_7961,N_9328);
or U12496 (N_12496,N_9089,N_6534);
nand U12497 (N_12497,N_7246,N_8443);
or U12498 (N_12498,N_9671,N_5654);
nor U12499 (N_12499,N_9643,N_7037);
nand U12500 (N_12500,N_8153,N_7086);
or U12501 (N_12501,N_5346,N_6632);
or U12502 (N_12502,N_6992,N_8213);
nand U12503 (N_12503,N_6852,N_7062);
nor U12504 (N_12504,N_7031,N_7363);
and U12505 (N_12505,N_9079,N_5476);
nor U12506 (N_12506,N_6107,N_7902);
nand U12507 (N_12507,N_6815,N_8398);
and U12508 (N_12508,N_9314,N_6807);
and U12509 (N_12509,N_7538,N_6064);
xnor U12510 (N_12510,N_8894,N_5460);
or U12511 (N_12511,N_9119,N_5754);
nor U12512 (N_12512,N_6106,N_9769);
nor U12513 (N_12513,N_9702,N_5269);
nor U12514 (N_12514,N_5472,N_9833);
and U12515 (N_12515,N_9319,N_7860);
or U12516 (N_12516,N_8708,N_9224);
or U12517 (N_12517,N_8269,N_7269);
or U12518 (N_12518,N_8730,N_5797);
nor U12519 (N_12519,N_9691,N_7576);
nor U12520 (N_12520,N_6499,N_8362);
and U12521 (N_12521,N_8362,N_7171);
nand U12522 (N_12522,N_5907,N_5461);
nand U12523 (N_12523,N_6494,N_9567);
nor U12524 (N_12524,N_5976,N_6434);
nand U12525 (N_12525,N_6392,N_9210);
nand U12526 (N_12526,N_8547,N_5814);
or U12527 (N_12527,N_5669,N_6619);
nand U12528 (N_12528,N_7362,N_7569);
nand U12529 (N_12529,N_8916,N_7187);
or U12530 (N_12530,N_6061,N_8665);
nand U12531 (N_12531,N_7358,N_8355);
or U12532 (N_12532,N_7789,N_6964);
or U12533 (N_12533,N_6393,N_6881);
nor U12534 (N_12534,N_8693,N_5465);
or U12535 (N_12535,N_5666,N_5111);
nand U12536 (N_12536,N_6212,N_5196);
or U12537 (N_12537,N_6258,N_7727);
nor U12538 (N_12538,N_5711,N_7903);
and U12539 (N_12539,N_9625,N_6536);
and U12540 (N_12540,N_9223,N_6820);
or U12541 (N_12541,N_9877,N_8371);
nand U12542 (N_12542,N_9949,N_7167);
or U12543 (N_12543,N_6267,N_9359);
or U12544 (N_12544,N_7929,N_8385);
nor U12545 (N_12545,N_8926,N_8799);
nand U12546 (N_12546,N_8509,N_7213);
and U12547 (N_12547,N_5067,N_8042);
nor U12548 (N_12548,N_9991,N_6136);
and U12549 (N_12549,N_5823,N_7200);
or U12550 (N_12550,N_7192,N_7153);
xor U12551 (N_12551,N_8369,N_9971);
or U12552 (N_12552,N_5248,N_9940);
nand U12553 (N_12553,N_9367,N_7606);
or U12554 (N_12554,N_5920,N_6943);
nand U12555 (N_12555,N_7631,N_7338);
nor U12556 (N_12556,N_9028,N_9587);
nand U12557 (N_12557,N_5715,N_7878);
nand U12558 (N_12558,N_8306,N_5644);
nor U12559 (N_12559,N_6706,N_7724);
or U12560 (N_12560,N_8222,N_6815);
nor U12561 (N_12561,N_9727,N_7328);
and U12562 (N_12562,N_8973,N_7588);
and U12563 (N_12563,N_8478,N_6528);
or U12564 (N_12564,N_8942,N_8762);
xor U12565 (N_12565,N_7816,N_9977);
nor U12566 (N_12566,N_7827,N_7969);
nand U12567 (N_12567,N_9827,N_8926);
nand U12568 (N_12568,N_6818,N_7203);
nor U12569 (N_12569,N_7637,N_5120);
or U12570 (N_12570,N_7255,N_5631);
and U12571 (N_12571,N_7874,N_8099);
nor U12572 (N_12572,N_6242,N_5161);
or U12573 (N_12573,N_9755,N_6778);
nand U12574 (N_12574,N_5317,N_6341);
or U12575 (N_12575,N_5979,N_5291);
nor U12576 (N_12576,N_6377,N_5667);
nand U12577 (N_12577,N_9661,N_8483);
and U12578 (N_12578,N_9754,N_6652);
nor U12579 (N_12579,N_9728,N_9724);
or U12580 (N_12580,N_6887,N_5530);
nand U12581 (N_12581,N_6187,N_9403);
and U12582 (N_12582,N_7674,N_6945);
nand U12583 (N_12583,N_8244,N_6803);
and U12584 (N_12584,N_7194,N_5672);
and U12585 (N_12585,N_7764,N_9763);
nand U12586 (N_12586,N_9924,N_8708);
or U12587 (N_12587,N_6312,N_7460);
nor U12588 (N_12588,N_5437,N_8417);
or U12589 (N_12589,N_8796,N_7461);
or U12590 (N_12590,N_5172,N_7020);
or U12591 (N_12591,N_7096,N_8763);
nand U12592 (N_12592,N_6027,N_7651);
nor U12593 (N_12593,N_5165,N_7804);
nand U12594 (N_12594,N_7065,N_6685);
nand U12595 (N_12595,N_9632,N_5069);
and U12596 (N_12596,N_8940,N_8772);
nand U12597 (N_12597,N_9507,N_9714);
nor U12598 (N_12598,N_5048,N_9234);
nor U12599 (N_12599,N_5880,N_5129);
and U12600 (N_12600,N_5653,N_6126);
and U12601 (N_12601,N_9614,N_6305);
nor U12602 (N_12602,N_5669,N_5990);
or U12603 (N_12603,N_6132,N_9923);
nor U12604 (N_12604,N_6182,N_8393);
and U12605 (N_12605,N_9997,N_7930);
and U12606 (N_12606,N_9050,N_5297);
nor U12607 (N_12607,N_6682,N_5367);
nor U12608 (N_12608,N_6910,N_8346);
or U12609 (N_12609,N_9311,N_5653);
and U12610 (N_12610,N_8308,N_7664);
or U12611 (N_12611,N_5168,N_6328);
and U12612 (N_12612,N_5138,N_9585);
or U12613 (N_12613,N_7713,N_7013);
and U12614 (N_12614,N_9792,N_9360);
or U12615 (N_12615,N_5394,N_6172);
or U12616 (N_12616,N_6290,N_7840);
or U12617 (N_12617,N_5457,N_5270);
nand U12618 (N_12618,N_5959,N_5593);
nor U12619 (N_12619,N_7074,N_5530);
nand U12620 (N_12620,N_5161,N_8084);
and U12621 (N_12621,N_8754,N_5125);
nand U12622 (N_12622,N_6186,N_5279);
or U12623 (N_12623,N_8042,N_7933);
and U12624 (N_12624,N_9419,N_6534);
and U12625 (N_12625,N_8348,N_6292);
nand U12626 (N_12626,N_6984,N_6110);
and U12627 (N_12627,N_8721,N_6759);
nor U12628 (N_12628,N_5735,N_9505);
and U12629 (N_12629,N_5582,N_9632);
or U12630 (N_12630,N_7115,N_6761);
or U12631 (N_12631,N_5061,N_6758);
and U12632 (N_12632,N_9290,N_8007);
nand U12633 (N_12633,N_8235,N_8302);
xnor U12634 (N_12634,N_5656,N_5977);
and U12635 (N_12635,N_5113,N_7056);
nor U12636 (N_12636,N_5828,N_9578);
and U12637 (N_12637,N_8366,N_9017);
or U12638 (N_12638,N_8759,N_5542);
nand U12639 (N_12639,N_9190,N_5160);
nor U12640 (N_12640,N_5546,N_6679);
and U12641 (N_12641,N_8155,N_8524);
and U12642 (N_12642,N_8885,N_8934);
and U12643 (N_12643,N_8145,N_7958);
nor U12644 (N_12644,N_7555,N_7619);
nor U12645 (N_12645,N_7606,N_6158);
and U12646 (N_12646,N_7962,N_8094);
or U12647 (N_12647,N_8662,N_5042);
nand U12648 (N_12648,N_5934,N_6786);
and U12649 (N_12649,N_6277,N_6259);
and U12650 (N_12650,N_8671,N_8011);
and U12651 (N_12651,N_5337,N_7852);
and U12652 (N_12652,N_5255,N_7487);
nor U12653 (N_12653,N_6950,N_7437);
nor U12654 (N_12654,N_9159,N_8494);
nor U12655 (N_12655,N_5171,N_7324);
nor U12656 (N_12656,N_9336,N_9571);
nor U12657 (N_12657,N_6921,N_9267);
nand U12658 (N_12658,N_6955,N_9803);
and U12659 (N_12659,N_7066,N_7491);
and U12660 (N_12660,N_7962,N_7051);
nor U12661 (N_12661,N_5774,N_8781);
nor U12662 (N_12662,N_9750,N_9122);
or U12663 (N_12663,N_8700,N_5251);
nor U12664 (N_12664,N_9192,N_7515);
or U12665 (N_12665,N_8204,N_6498);
or U12666 (N_12666,N_5126,N_8991);
and U12667 (N_12667,N_9049,N_7067);
or U12668 (N_12668,N_9543,N_7655);
or U12669 (N_12669,N_8614,N_6272);
nand U12670 (N_12670,N_6567,N_6109);
nor U12671 (N_12671,N_6075,N_6720);
nand U12672 (N_12672,N_7255,N_5821);
or U12673 (N_12673,N_5489,N_9251);
nor U12674 (N_12674,N_5351,N_8217);
xor U12675 (N_12675,N_8372,N_5937);
or U12676 (N_12676,N_9556,N_7664);
nor U12677 (N_12677,N_6557,N_6950);
nand U12678 (N_12678,N_7170,N_5469);
and U12679 (N_12679,N_8031,N_8382);
or U12680 (N_12680,N_5729,N_8345);
nor U12681 (N_12681,N_5944,N_8976);
or U12682 (N_12682,N_9822,N_7692);
nor U12683 (N_12683,N_6308,N_6077);
or U12684 (N_12684,N_9681,N_5123);
xnor U12685 (N_12685,N_7755,N_8398);
and U12686 (N_12686,N_9422,N_5141);
and U12687 (N_12687,N_6337,N_8181);
or U12688 (N_12688,N_7841,N_6399);
xor U12689 (N_12689,N_7445,N_9353);
and U12690 (N_12690,N_9569,N_7504);
nand U12691 (N_12691,N_6859,N_7942);
nor U12692 (N_12692,N_6259,N_5960);
nor U12693 (N_12693,N_9917,N_6270);
nand U12694 (N_12694,N_7301,N_7947);
nor U12695 (N_12695,N_9803,N_5394);
or U12696 (N_12696,N_5483,N_6702);
xor U12697 (N_12697,N_7586,N_9977);
and U12698 (N_12698,N_5865,N_5104);
nor U12699 (N_12699,N_8548,N_7769);
and U12700 (N_12700,N_6794,N_9936);
xor U12701 (N_12701,N_6919,N_6786);
nand U12702 (N_12702,N_9702,N_6271);
nor U12703 (N_12703,N_7820,N_8656);
nor U12704 (N_12704,N_6567,N_5300);
nor U12705 (N_12705,N_9333,N_5880);
nand U12706 (N_12706,N_6538,N_7580);
nor U12707 (N_12707,N_8417,N_9645);
and U12708 (N_12708,N_9524,N_5205);
and U12709 (N_12709,N_6889,N_9062);
nand U12710 (N_12710,N_9661,N_8035);
or U12711 (N_12711,N_7887,N_5466);
nand U12712 (N_12712,N_6006,N_7513);
nand U12713 (N_12713,N_9482,N_9020);
and U12714 (N_12714,N_8566,N_8756);
or U12715 (N_12715,N_9222,N_5546);
nor U12716 (N_12716,N_7885,N_8168);
nor U12717 (N_12717,N_6283,N_5807);
or U12718 (N_12718,N_5380,N_7343);
nor U12719 (N_12719,N_5680,N_6438);
or U12720 (N_12720,N_5407,N_9918);
nand U12721 (N_12721,N_6785,N_9939);
nor U12722 (N_12722,N_5288,N_8843);
and U12723 (N_12723,N_9385,N_7376);
nor U12724 (N_12724,N_6124,N_8646);
or U12725 (N_12725,N_9554,N_9847);
or U12726 (N_12726,N_6528,N_8252);
and U12727 (N_12727,N_9368,N_8420);
nor U12728 (N_12728,N_6373,N_6908);
or U12729 (N_12729,N_7159,N_6114);
nand U12730 (N_12730,N_9929,N_7785);
and U12731 (N_12731,N_7664,N_7097);
and U12732 (N_12732,N_8380,N_6192);
nor U12733 (N_12733,N_6549,N_9779);
nand U12734 (N_12734,N_7444,N_9757);
nor U12735 (N_12735,N_6966,N_7247);
or U12736 (N_12736,N_8756,N_5690);
and U12737 (N_12737,N_6545,N_6255);
and U12738 (N_12738,N_5641,N_7686);
nand U12739 (N_12739,N_8786,N_6538);
nand U12740 (N_12740,N_8199,N_8001);
or U12741 (N_12741,N_8556,N_9288);
and U12742 (N_12742,N_9867,N_7262);
nand U12743 (N_12743,N_6032,N_7964);
and U12744 (N_12744,N_7514,N_6442);
nand U12745 (N_12745,N_7675,N_7874);
and U12746 (N_12746,N_8295,N_5988);
or U12747 (N_12747,N_6481,N_7250);
and U12748 (N_12748,N_6554,N_5896);
nor U12749 (N_12749,N_5112,N_7525);
and U12750 (N_12750,N_7091,N_5883);
and U12751 (N_12751,N_9046,N_9150);
nor U12752 (N_12752,N_6911,N_8657);
nand U12753 (N_12753,N_7025,N_8648);
nor U12754 (N_12754,N_6089,N_8154);
nor U12755 (N_12755,N_9662,N_8645);
or U12756 (N_12756,N_5081,N_9880);
and U12757 (N_12757,N_5357,N_8197);
nor U12758 (N_12758,N_6656,N_6985);
or U12759 (N_12759,N_5028,N_6089);
nor U12760 (N_12760,N_6834,N_6908);
nor U12761 (N_12761,N_8029,N_6353);
nor U12762 (N_12762,N_7699,N_5069);
or U12763 (N_12763,N_7158,N_7178);
and U12764 (N_12764,N_6591,N_9309);
nand U12765 (N_12765,N_9050,N_6558);
nand U12766 (N_12766,N_8526,N_6581);
or U12767 (N_12767,N_7622,N_6237);
nor U12768 (N_12768,N_8576,N_6682);
nor U12769 (N_12769,N_5754,N_8852);
nand U12770 (N_12770,N_5329,N_9435);
or U12771 (N_12771,N_7399,N_6986);
nand U12772 (N_12772,N_6776,N_8823);
xor U12773 (N_12773,N_5905,N_5323);
nand U12774 (N_12774,N_7281,N_6264);
nand U12775 (N_12775,N_8732,N_8254);
xor U12776 (N_12776,N_9455,N_8071);
or U12777 (N_12777,N_5145,N_5540);
nor U12778 (N_12778,N_6771,N_7634);
nor U12779 (N_12779,N_9443,N_5669);
and U12780 (N_12780,N_7308,N_9897);
or U12781 (N_12781,N_7341,N_7414);
and U12782 (N_12782,N_7871,N_9191);
nand U12783 (N_12783,N_5705,N_5598);
or U12784 (N_12784,N_8895,N_6510);
and U12785 (N_12785,N_8168,N_9853);
or U12786 (N_12786,N_9545,N_7661);
nand U12787 (N_12787,N_5218,N_8493);
or U12788 (N_12788,N_7384,N_5775);
and U12789 (N_12789,N_7830,N_6041);
or U12790 (N_12790,N_5605,N_8083);
xnor U12791 (N_12791,N_9277,N_9948);
and U12792 (N_12792,N_7502,N_8007);
or U12793 (N_12793,N_5035,N_8881);
and U12794 (N_12794,N_6816,N_9807);
nor U12795 (N_12795,N_5009,N_8529);
nand U12796 (N_12796,N_7332,N_5376);
and U12797 (N_12797,N_8374,N_7947);
and U12798 (N_12798,N_5997,N_9332);
and U12799 (N_12799,N_8579,N_5829);
xnor U12800 (N_12800,N_6162,N_9629);
nor U12801 (N_12801,N_7123,N_6738);
and U12802 (N_12802,N_6893,N_7603);
or U12803 (N_12803,N_8591,N_9101);
or U12804 (N_12804,N_7702,N_8142);
or U12805 (N_12805,N_7488,N_8283);
nand U12806 (N_12806,N_9686,N_8776);
nand U12807 (N_12807,N_6444,N_6252);
nand U12808 (N_12808,N_7288,N_5170);
and U12809 (N_12809,N_9944,N_7613);
nor U12810 (N_12810,N_6998,N_7330);
nor U12811 (N_12811,N_5857,N_5894);
nand U12812 (N_12812,N_6402,N_6633);
or U12813 (N_12813,N_8075,N_9740);
nor U12814 (N_12814,N_5654,N_5728);
nand U12815 (N_12815,N_5416,N_6400);
xor U12816 (N_12816,N_9662,N_7404);
or U12817 (N_12817,N_5180,N_9973);
or U12818 (N_12818,N_5834,N_8537);
or U12819 (N_12819,N_8858,N_5415);
nor U12820 (N_12820,N_7412,N_9737);
and U12821 (N_12821,N_9935,N_5661);
nor U12822 (N_12822,N_7684,N_8273);
nor U12823 (N_12823,N_9513,N_6994);
nand U12824 (N_12824,N_5922,N_6761);
nor U12825 (N_12825,N_7254,N_5940);
nand U12826 (N_12826,N_9154,N_9633);
nor U12827 (N_12827,N_7397,N_8910);
nand U12828 (N_12828,N_9334,N_6685);
and U12829 (N_12829,N_7483,N_7931);
nand U12830 (N_12830,N_9630,N_8836);
nor U12831 (N_12831,N_7797,N_7561);
or U12832 (N_12832,N_5078,N_5452);
and U12833 (N_12833,N_9500,N_9815);
or U12834 (N_12834,N_6732,N_5094);
nand U12835 (N_12835,N_5979,N_7751);
or U12836 (N_12836,N_7670,N_9700);
nor U12837 (N_12837,N_7606,N_7942);
or U12838 (N_12838,N_8606,N_6387);
nand U12839 (N_12839,N_8003,N_7841);
or U12840 (N_12840,N_8472,N_7719);
and U12841 (N_12841,N_6048,N_5052);
nor U12842 (N_12842,N_9379,N_9937);
nand U12843 (N_12843,N_7807,N_6436);
nand U12844 (N_12844,N_9307,N_5170);
and U12845 (N_12845,N_7544,N_7270);
nand U12846 (N_12846,N_6812,N_5387);
nand U12847 (N_12847,N_8878,N_8410);
and U12848 (N_12848,N_8091,N_5397);
nor U12849 (N_12849,N_5138,N_7736);
xor U12850 (N_12850,N_6843,N_9296);
or U12851 (N_12851,N_7460,N_8393);
and U12852 (N_12852,N_7133,N_9070);
and U12853 (N_12853,N_8474,N_8191);
nand U12854 (N_12854,N_7381,N_5358);
or U12855 (N_12855,N_9885,N_5824);
or U12856 (N_12856,N_8355,N_5172);
nand U12857 (N_12857,N_6159,N_7947);
nand U12858 (N_12858,N_8146,N_7332);
and U12859 (N_12859,N_9414,N_6960);
or U12860 (N_12860,N_8070,N_8161);
nor U12861 (N_12861,N_9618,N_7839);
xnor U12862 (N_12862,N_8767,N_5364);
nand U12863 (N_12863,N_9399,N_7268);
and U12864 (N_12864,N_8754,N_5353);
and U12865 (N_12865,N_6126,N_8604);
or U12866 (N_12866,N_7694,N_8619);
and U12867 (N_12867,N_5644,N_7999);
and U12868 (N_12868,N_9633,N_5458);
nor U12869 (N_12869,N_7836,N_8960);
nor U12870 (N_12870,N_6649,N_6619);
or U12871 (N_12871,N_7375,N_9448);
nand U12872 (N_12872,N_8458,N_5482);
nand U12873 (N_12873,N_7739,N_6050);
or U12874 (N_12874,N_6435,N_5907);
xnor U12875 (N_12875,N_6394,N_9466);
nand U12876 (N_12876,N_7887,N_6093);
nor U12877 (N_12877,N_7670,N_5200);
nand U12878 (N_12878,N_6884,N_6702);
xnor U12879 (N_12879,N_8861,N_7914);
nor U12880 (N_12880,N_7787,N_7014);
nand U12881 (N_12881,N_6245,N_6346);
nand U12882 (N_12882,N_6465,N_8277);
or U12883 (N_12883,N_7159,N_9313);
nand U12884 (N_12884,N_8759,N_5453);
or U12885 (N_12885,N_6839,N_8891);
and U12886 (N_12886,N_5779,N_9440);
or U12887 (N_12887,N_5608,N_8206);
nor U12888 (N_12888,N_9901,N_8109);
and U12889 (N_12889,N_9127,N_9938);
or U12890 (N_12890,N_5835,N_5036);
nand U12891 (N_12891,N_7428,N_5512);
nand U12892 (N_12892,N_5865,N_7026);
nor U12893 (N_12893,N_9701,N_7301);
and U12894 (N_12894,N_9391,N_6439);
nand U12895 (N_12895,N_6846,N_7902);
nand U12896 (N_12896,N_8801,N_5698);
or U12897 (N_12897,N_8592,N_6628);
or U12898 (N_12898,N_9038,N_9715);
nand U12899 (N_12899,N_7350,N_9726);
nor U12900 (N_12900,N_6570,N_8357);
nand U12901 (N_12901,N_6436,N_6424);
and U12902 (N_12902,N_6060,N_6301);
or U12903 (N_12903,N_5012,N_9843);
nand U12904 (N_12904,N_8095,N_9900);
and U12905 (N_12905,N_5338,N_8208);
and U12906 (N_12906,N_5251,N_9245);
and U12907 (N_12907,N_6466,N_5623);
and U12908 (N_12908,N_9516,N_8427);
or U12909 (N_12909,N_6537,N_7460);
or U12910 (N_12910,N_9387,N_6292);
nor U12911 (N_12911,N_8630,N_9214);
nand U12912 (N_12912,N_7208,N_8037);
nor U12913 (N_12913,N_5477,N_8158);
nand U12914 (N_12914,N_6065,N_7269);
nand U12915 (N_12915,N_8183,N_5373);
nor U12916 (N_12916,N_6165,N_5772);
and U12917 (N_12917,N_8136,N_5936);
or U12918 (N_12918,N_6311,N_8531);
nor U12919 (N_12919,N_5399,N_7968);
or U12920 (N_12920,N_8928,N_8372);
nand U12921 (N_12921,N_7687,N_5842);
nor U12922 (N_12922,N_7434,N_9365);
and U12923 (N_12923,N_5187,N_5719);
and U12924 (N_12924,N_6728,N_6715);
and U12925 (N_12925,N_7593,N_9634);
nor U12926 (N_12926,N_9456,N_6885);
or U12927 (N_12927,N_6577,N_7706);
nand U12928 (N_12928,N_7358,N_8062);
or U12929 (N_12929,N_6290,N_7222);
xnor U12930 (N_12930,N_9317,N_9598);
nand U12931 (N_12931,N_9307,N_8843);
nor U12932 (N_12932,N_6863,N_7311);
or U12933 (N_12933,N_9323,N_8462);
nand U12934 (N_12934,N_5797,N_6758);
nand U12935 (N_12935,N_6727,N_8962);
or U12936 (N_12936,N_6807,N_5921);
and U12937 (N_12937,N_6339,N_9258);
or U12938 (N_12938,N_9740,N_8788);
nand U12939 (N_12939,N_5432,N_6828);
nor U12940 (N_12940,N_6431,N_6089);
or U12941 (N_12941,N_9496,N_5077);
or U12942 (N_12942,N_9438,N_6056);
and U12943 (N_12943,N_9765,N_8831);
or U12944 (N_12944,N_9850,N_8684);
nand U12945 (N_12945,N_9294,N_9846);
nand U12946 (N_12946,N_8911,N_6660);
nand U12947 (N_12947,N_5452,N_8776);
and U12948 (N_12948,N_6765,N_9456);
nand U12949 (N_12949,N_5878,N_9252);
and U12950 (N_12950,N_5709,N_7843);
nand U12951 (N_12951,N_5755,N_5849);
nor U12952 (N_12952,N_6368,N_9449);
nand U12953 (N_12953,N_9750,N_5103);
or U12954 (N_12954,N_8815,N_8620);
nor U12955 (N_12955,N_7019,N_8334);
nor U12956 (N_12956,N_6416,N_7537);
and U12957 (N_12957,N_8092,N_7203);
or U12958 (N_12958,N_9379,N_8931);
nand U12959 (N_12959,N_8532,N_7409);
nor U12960 (N_12960,N_6181,N_5060);
nand U12961 (N_12961,N_7764,N_8843);
nor U12962 (N_12962,N_7252,N_6581);
and U12963 (N_12963,N_5336,N_9573);
and U12964 (N_12964,N_6351,N_7700);
or U12965 (N_12965,N_8682,N_6932);
and U12966 (N_12966,N_6959,N_5342);
and U12967 (N_12967,N_6128,N_5283);
nand U12968 (N_12968,N_7792,N_6817);
and U12969 (N_12969,N_7475,N_9981);
and U12970 (N_12970,N_8455,N_9275);
or U12971 (N_12971,N_9556,N_8170);
nor U12972 (N_12972,N_5750,N_5013);
nor U12973 (N_12973,N_6283,N_7734);
and U12974 (N_12974,N_7364,N_8618);
nand U12975 (N_12975,N_5278,N_7581);
nand U12976 (N_12976,N_7251,N_9793);
and U12977 (N_12977,N_6934,N_8689);
and U12978 (N_12978,N_7374,N_5169);
xor U12979 (N_12979,N_7372,N_5418);
or U12980 (N_12980,N_5796,N_8188);
and U12981 (N_12981,N_6372,N_8336);
nor U12982 (N_12982,N_6451,N_7357);
and U12983 (N_12983,N_6005,N_8758);
nor U12984 (N_12984,N_5263,N_9907);
and U12985 (N_12985,N_8846,N_7105);
xnor U12986 (N_12986,N_5586,N_7270);
nand U12987 (N_12987,N_9109,N_5073);
or U12988 (N_12988,N_7469,N_8172);
nor U12989 (N_12989,N_5552,N_6609);
or U12990 (N_12990,N_8768,N_8877);
or U12991 (N_12991,N_5147,N_7174);
and U12992 (N_12992,N_6056,N_6583);
or U12993 (N_12993,N_6902,N_8617);
nand U12994 (N_12994,N_8471,N_5295);
nor U12995 (N_12995,N_7711,N_8674);
nand U12996 (N_12996,N_8631,N_6086);
and U12997 (N_12997,N_9511,N_5944);
and U12998 (N_12998,N_8258,N_8267);
nor U12999 (N_12999,N_9246,N_9763);
nand U13000 (N_13000,N_5649,N_8866);
nor U13001 (N_13001,N_8291,N_9178);
xnor U13002 (N_13002,N_9938,N_8862);
nor U13003 (N_13003,N_9768,N_5789);
nor U13004 (N_13004,N_6052,N_9256);
and U13005 (N_13005,N_6709,N_9359);
nand U13006 (N_13006,N_5097,N_5246);
nand U13007 (N_13007,N_7373,N_8621);
and U13008 (N_13008,N_5600,N_9840);
nor U13009 (N_13009,N_8048,N_5198);
and U13010 (N_13010,N_9000,N_5808);
nor U13011 (N_13011,N_8881,N_9701);
nor U13012 (N_13012,N_8861,N_8118);
nand U13013 (N_13013,N_5503,N_8059);
nand U13014 (N_13014,N_7222,N_6609);
or U13015 (N_13015,N_9011,N_6999);
nor U13016 (N_13016,N_8193,N_5475);
and U13017 (N_13017,N_6276,N_8773);
nand U13018 (N_13018,N_5668,N_7746);
or U13019 (N_13019,N_8152,N_5377);
or U13020 (N_13020,N_7269,N_7088);
or U13021 (N_13021,N_5248,N_8688);
and U13022 (N_13022,N_7537,N_9368);
nor U13023 (N_13023,N_5797,N_7158);
nand U13024 (N_13024,N_8577,N_7818);
or U13025 (N_13025,N_8404,N_5369);
nor U13026 (N_13026,N_7420,N_9434);
nand U13027 (N_13027,N_6842,N_6608);
nor U13028 (N_13028,N_6025,N_6671);
nand U13029 (N_13029,N_6620,N_6518);
or U13030 (N_13030,N_7794,N_8978);
nand U13031 (N_13031,N_9984,N_8793);
nand U13032 (N_13032,N_5604,N_6323);
nand U13033 (N_13033,N_5144,N_6053);
nor U13034 (N_13034,N_7382,N_9156);
nand U13035 (N_13035,N_5687,N_9688);
nor U13036 (N_13036,N_9526,N_8275);
nor U13037 (N_13037,N_9640,N_6042);
nor U13038 (N_13038,N_5361,N_8458);
and U13039 (N_13039,N_9843,N_5814);
and U13040 (N_13040,N_5830,N_6211);
nor U13041 (N_13041,N_8170,N_7213);
nor U13042 (N_13042,N_9178,N_7395);
nor U13043 (N_13043,N_5899,N_8539);
nor U13044 (N_13044,N_5554,N_9552);
nand U13045 (N_13045,N_9281,N_9721);
or U13046 (N_13046,N_5483,N_9432);
nor U13047 (N_13047,N_5037,N_7654);
or U13048 (N_13048,N_8221,N_8041);
and U13049 (N_13049,N_7345,N_5644);
nor U13050 (N_13050,N_9213,N_7820);
and U13051 (N_13051,N_7601,N_8895);
and U13052 (N_13052,N_6547,N_8082);
and U13053 (N_13053,N_5082,N_6760);
and U13054 (N_13054,N_6313,N_8611);
or U13055 (N_13055,N_9848,N_9883);
and U13056 (N_13056,N_8169,N_5833);
and U13057 (N_13057,N_5250,N_6346);
or U13058 (N_13058,N_7057,N_6918);
or U13059 (N_13059,N_9868,N_5584);
nand U13060 (N_13060,N_8803,N_7073);
or U13061 (N_13061,N_9951,N_8310);
nand U13062 (N_13062,N_9575,N_8335);
nor U13063 (N_13063,N_9860,N_6616);
and U13064 (N_13064,N_6980,N_8222);
nor U13065 (N_13065,N_7609,N_9850);
nand U13066 (N_13066,N_7833,N_7081);
and U13067 (N_13067,N_7453,N_5561);
nand U13068 (N_13068,N_9124,N_8729);
nor U13069 (N_13069,N_9222,N_6350);
nor U13070 (N_13070,N_5551,N_8379);
and U13071 (N_13071,N_8178,N_5661);
or U13072 (N_13072,N_7325,N_5346);
nor U13073 (N_13073,N_7030,N_8175);
or U13074 (N_13074,N_7880,N_9265);
nor U13075 (N_13075,N_7905,N_7848);
nand U13076 (N_13076,N_9825,N_9458);
or U13077 (N_13077,N_7579,N_8882);
or U13078 (N_13078,N_8756,N_9788);
and U13079 (N_13079,N_7157,N_8700);
nor U13080 (N_13080,N_7789,N_5194);
and U13081 (N_13081,N_9855,N_8433);
and U13082 (N_13082,N_5900,N_8545);
nand U13083 (N_13083,N_9033,N_8269);
or U13084 (N_13084,N_5827,N_5874);
xnor U13085 (N_13085,N_8096,N_5614);
nand U13086 (N_13086,N_8442,N_7120);
nor U13087 (N_13087,N_9321,N_7378);
and U13088 (N_13088,N_5512,N_8302);
or U13089 (N_13089,N_7514,N_5303);
nor U13090 (N_13090,N_9399,N_7118);
and U13091 (N_13091,N_6116,N_5661);
nand U13092 (N_13092,N_6181,N_8849);
and U13093 (N_13093,N_6130,N_5673);
nand U13094 (N_13094,N_8826,N_9451);
nor U13095 (N_13095,N_9611,N_5304);
and U13096 (N_13096,N_7838,N_7074);
or U13097 (N_13097,N_9265,N_5374);
and U13098 (N_13098,N_7897,N_7977);
and U13099 (N_13099,N_9289,N_6251);
and U13100 (N_13100,N_8476,N_5790);
xor U13101 (N_13101,N_8919,N_6342);
or U13102 (N_13102,N_8476,N_6000);
and U13103 (N_13103,N_5785,N_7263);
nor U13104 (N_13104,N_5805,N_9179);
nand U13105 (N_13105,N_6630,N_9843);
nor U13106 (N_13106,N_6099,N_6317);
and U13107 (N_13107,N_9647,N_7295);
and U13108 (N_13108,N_9560,N_5351);
nand U13109 (N_13109,N_6756,N_5733);
nand U13110 (N_13110,N_9515,N_5130);
or U13111 (N_13111,N_5312,N_7829);
or U13112 (N_13112,N_5291,N_5305);
or U13113 (N_13113,N_7842,N_5128);
or U13114 (N_13114,N_5406,N_6751);
and U13115 (N_13115,N_6869,N_7070);
nor U13116 (N_13116,N_8852,N_6696);
nand U13117 (N_13117,N_5166,N_6410);
nor U13118 (N_13118,N_9572,N_6283);
nor U13119 (N_13119,N_9323,N_6486);
or U13120 (N_13120,N_5156,N_7159);
nor U13121 (N_13121,N_6215,N_7568);
and U13122 (N_13122,N_6484,N_8880);
and U13123 (N_13123,N_5562,N_5362);
nor U13124 (N_13124,N_7871,N_6131);
nand U13125 (N_13125,N_9909,N_6357);
nor U13126 (N_13126,N_9398,N_5005);
and U13127 (N_13127,N_5526,N_5747);
and U13128 (N_13128,N_6330,N_9516);
or U13129 (N_13129,N_9139,N_9640);
nand U13130 (N_13130,N_6880,N_6675);
or U13131 (N_13131,N_9474,N_7307);
or U13132 (N_13132,N_6759,N_6527);
or U13133 (N_13133,N_6420,N_6694);
nor U13134 (N_13134,N_9024,N_7951);
or U13135 (N_13135,N_9097,N_6705);
nor U13136 (N_13136,N_6331,N_5127);
nand U13137 (N_13137,N_8922,N_9111);
nand U13138 (N_13138,N_9660,N_6569);
or U13139 (N_13139,N_5383,N_5049);
or U13140 (N_13140,N_7620,N_8132);
or U13141 (N_13141,N_5751,N_6046);
nor U13142 (N_13142,N_8224,N_9439);
nand U13143 (N_13143,N_7647,N_5367);
and U13144 (N_13144,N_8874,N_7772);
or U13145 (N_13145,N_9018,N_5793);
nor U13146 (N_13146,N_7583,N_8199);
and U13147 (N_13147,N_8465,N_9162);
and U13148 (N_13148,N_9353,N_7788);
and U13149 (N_13149,N_8910,N_5003);
and U13150 (N_13150,N_9789,N_6199);
nor U13151 (N_13151,N_6650,N_7316);
and U13152 (N_13152,N_5028,N_8537);
or U13153 (N_13153,N_8045,N_6763);
or U13154 (N_13154,N_7754,N_6436);
xnor U13155 (N_13155,N_5126,N_5893);
nand U13156 (N_13156,N_7014,N_8570);
nand U13157 (N_13157,N_8743,N_9692);
and U13158 (N_13158,N_7289,N_8937);
nor U13159 (N_13159,N_8252,N_9195);
and U13160 (N_13160,N_6661,N_7310);
nor U13161 (N_13161,N_9837,N_7025);
and U13162 (N_13162,N_9361,N_9033);
nand U13163 (N_13163,N_6970,N_9333);
nand U13164 (N_13164,N_8874,N_8581);
nor U13165 (N_13165,N_8176,N_5925);
or U13166 (N_13166,N_7923,N_5114);
and U13167 (N_13167,N_7460,N_7491);
nand U13168 (N_13168,N_5369,N_6418);
nand U13169 (N_13169,N_6255,N_5721);
nand U13170 (N_13170,N_6429,N_6722);
and U13171 (N_13171,N_6188,N_6298);
and U13172 (N_13172,N_5344,N_9081);
nand U13173 (N_13173,N_8527,N_9089);
nand U13174 (N_13174,N_9814,N_7038);
or U13175 (N_13175,N_9650,N_8863);
or U13176 (N_13176,N_6457,N_5473);
nand U13177 (N_13177,N_9877,N_9873);
nor U13178 (N_13178,N_8158,N_5432);
nor U13179 (N_13179,N_7212,N_7349);
nor U13180 (N_13180,N_6785,N_5374);
nand U13181 (N_13181,N_5934,N_9407);
and U13182 (N_13182,N_6852,N_9113);
nand U13183 (N_13183,N_6280,N_7596);
and U13184 (N_13184,N_9216,N_8920);
nor U13185 (N_13185,N_8927,N_5768);
nand U13186 (N_13186,N_5924,N_5843);
or U13187 (N_13187,N_6001,N_9016);
or U13188 (N_13188,N_7747,N_9648);
or U13189 (N_13189,N_7083,N_9840);
nand U13190 (N_13190,N_7164,N_8810);
or U13191 (N_13191,N_9757,N_9106);
nand U13192 (N_13192,N_9357,N_9367);
xor U13193 (N_13193,N_8470,N_8512);
and U13194 (N_13194,N_5805,N_7169);
nand U13195 (N_13195,N_9851,N_9514);
nand U13196 (N_13196,N_7109,N_9626);
and U13197 (N_13197,N_5195,N_7931);
nand U13198 (N_13198,N_9390,N_5435);
nand U13199 (N_13199,N_8343,N_7658);
or U13200 (N_13200,N_6158,N_6275);
or U13201 (N_13201,N_7786,N_5141);
and U13202 (N_13202,N_6934,N_5095);
or U13203 (N_13203,N_5841,N_9961);
xor U13204 (N_13204,N_9115,N_8439);
and U13205 (N_13205,N_6251,N_5102);
nand U13206 (N_13206,N_7462,N_5813);
or U13207 (N_13207,N_9798,N_7151);
or U13208 (N_13208,N_5322,N_5465);
nor U13209 (N_13209,N_5792,N_7660);
nand U13210 (N_13210,N_9174,N_9871);
nand U13211 (N_13211,N_8156,N_8028);
nand U13212 (N_13212,N_9872,N_5892);
nor U13213 (N_13213,N_6883,N_6721);
nor U13214 (N_13214,N_7873,N_9082);
or U13215 (N_13215,N_5235,N_9149);
nor U13216 (N_13216,N_8958,N_9245);
or U13217 (N_13217,N_6815,N_8807);
nand U13218 (N_13218,N_7658,N_9463);
nand U13219 (N_13219,N_6750,N_5376);
or U13220 (N_13220,N_9490,N_5360);
xor U13221 (N_13221,N_7140,N_8570);
or U13222 (N_13222,N_5918,N_8046);
or U13223 (N_13223,N_5493,N_7616);
nor U13224 (N_13224,N_5677,N_6591);
nand U13225 (N_13225,N_5195,N_9693);
nor U13226 (N_13226,N_6997,N_5749);
nand U13227 (N_13227,N_7448,N_8424);
nand U13228 (N_13228,N_7644,N_5686);
and U13229 (N_13229,N_7871,N_8265);
and U13230 (N_13230,N_5399,N_5390);
and U13231 (N_13231,N_6903,N_8935);
nand U13232 (N_13232,N_9149,N_5983);
nor U13233 (N_13233,N_5429,N_5527);
nand U13234 (N_13234,N_7838,N_8802);
and U13235 (N_13235,N_8139,N_5396);
nor U13236 (N_13236,N_8237,N_7100);
nor U13237 (N_13237,N_9737,N_5757);
nand U13238 (N_13238,N_8653,N_8513);
or U13239 (N_13239,N_6470,N_5212);
and U13240 (N_13240,N_8616,N_6422);
or U13241 (N_13241,N_8623,N_9689);
nand U13242 (N_13242,N_7632,N_9364);
nand U13243 (N_13243,N_7573,N_9842);
nand U13244 (N_13244,N_6593,N_7421);
and U13245 (N_13245,N_5612,N_9390);
nor U13246 (N_13246,N_8082,N_9974);
or U13247 (N_13247,N_7882,N_6012);
or U13248 (N_13248,N_6051,N_5741);
nor U13249 (N_13249,N_9969,N_6287);
and U13250 (N_13250,N_5420,N_8300);
and U13251 (N_13251,N_6129,N_5251);
or U13252 (N_13252,N_7432,N_9447);
nor U13253 (N_13253,N_7732,N_7201);
or U13254 (N_13254,N_6761,N_7501);
nor U13255 (N_13255,N_5694,N_5710);
or U13256 (N_13256,N_6861,N_9982);
and U13257 (N_13257,N_8960,N_6425);
nand U13258 (N_13258,N_9007,N_8948);
or U13259 (N_13259,N_8851,N_9196);
nor U13260 (N_13260,N_6146,N_7990);
and U13261 (N_13261,N_7443,N_5735);
or U13262 (N_13262,N_7342,N_8595);
and U13263 (N_13263,N_5377,N_7386);
nand U13264 (N_13264,N_6245,N_6762);
or U13265 (N_13265,N_7055,N_7728);
and U13266 (N_13266,N_6996,N_9177);
nand U13267 (N_13267,N_8360,N_6290);
nor U13268 (N_13268,N_6215,N_8792);
or U13269 (N_13269,N_6927,N_9110);
nor U13270 (N_13270,N_9043,N_7411);
nand U13271 (N_13271,N_9086,N_5203);
or U13272 (N_13272,N_8993,N_7918);
or U13273 (N_13273,N_7066,N_6277);
nand U13274 (N_13274,N_9706,N_8276);
nor U13275 (N_13275,N_8711,N_8310);
and U13276 (N_13276,N_5354,N_5966);
nand U13277 (N_13277,N_9478,N_5804);
or U13278 (N_13278,N_6447,N_6108);
nor U13279 (N_13279,N_9634,N_9705);
nor U13280 (N_13280,N_6935,N_7783);
or U13281 (N_13281,N_9008,N_7682);
nand U13282 (N_13282,N_5004,N_9876);
and U13283 (N_13283,N_5811,N_8225);
or U13284 (N_13284,N_6752,N_7243);
nor U13285 (N_13285,N_8002,N_6339);
nor U13286 (N_13286,N_7734,N_7711);
nand U13287 (N_13287,N_5823,N_8620);
nand U13288 (N_13288,N_5458,N_7962);
nor U13289 (N_13289,N_9481,N_9422);
xor U13290 (N_13290,N_8560,N_8248);
and U13291 (N_13291,N_8053,N_7506);
or U13292 (N_13292,N_9261,N_9894);
xor U13293 (N_13293,N_7355,N_8216);
nor U13294 (N_13294,N_7455,N_8282);
or U13295 (N_13295,N_5729,N_8536);
nand U13296 (N_13296,N_6884,N_5630);
or U13297 (N_13297,N_7020,N_6865);
and U13298 (N_13298,N_7366,N_9504);
nand U13299 (N_13299,N_6512,N_9031);
xnor U13300 (N_13300,N_9412,N_5371);
and U13301 (N_13301,N_9995,N_9341);
and U13302 (N_13302,N_7277,N_6541);
nand U13303 (N_13303,N_7007,N_7921);
nand U13304 (N_13304,N_9668,N_5907);
or U13305 (N_13305,N_5583,N_5021);
or U13306 (N_13306,N_9148,N_9212);
nand U13307 (N_13307,N_7785,N_6649);
nor U13308 (N_13308,N_7860,N_9999);
and U13309 (N_13309,N_7603,N_6564);
nand U13310 (N_13310,N_7227,N_8974);
nor U13311 (N_13311,N_8740,N_8864);
nand U13312 (N_13312,N_7537,N_6967);
nand U13313 (N_13313,N_8547,N_9932);
and U13314 (N_13314,N_9022,N_7897);
or U13315 (N_13315,N_9869,N_6337);
or U13316 (N_13316,N_9533,N_8310);
or U13317 (N_13317,N_5532,N_6463);
nand U13318 (N_13318,N_7548,N_5708);
nand U13319 (N_13319,N_7331,N_6523);
and U13320 (N_13320,N_8434,N_6613);
nor U13321 (N_13321,N_7142,N_8402);
nand U13322 (N_13322,N_7340,N_8332);
nand U13323 (N_13323,N_5281,N_6598);
nor U13324 (N_13324,N_5043,N_9219);
and U13325 (N_13325,N_5768,N_7454);
nand U13326 (N_13326,N_6678,N_8522);
or U13327 (N_13327,N_7946,N_9468);
nand U13328 (N_13328,N_8144,N_8279);
and U13329 (N_13329,N_9051,N_7563);
or U13330 (N_13330,N_5589,N_6508);
nand U13331 (N_13331,N_7679,N_6733);
nor U13332 (N_13332,N_9341,N_6203);
nor U13333 (N_13333,N_7146,N_6449);
or U13334 (N_13334,N_6182,N_5055);
or U13335 (N_13335,N_8330,N_7854);
or U13336 (N_13336,N_8507,N_8815);
nand U13337 (N_13337,N_5913,N_7834);
nand U13338 (N_13338,N_8404,N_9428);
and U13339 (N_13339,N_8328,N_5544);
nand U13340 (N_13340,N_5579,N_9267);
nand U13341 (N_13341,N_9362,N_6110);
nand U13342 (N_13342,N_7595,N_5633);
nor U13343 (N_13343,N_7695,N_8832);
and U13344 (N_13344,N_9925,N_9910);
nand U13345 (N_13345,N_5480,N_9306);
nor U13346 (N_13346,N_6025,N_5498);
nand U13347 (N_13347,N_6117,N_7753);
and U13348 (N_13348,N_5060,N_7295);
nand U13349 (N_13349,N_7648,N_6373);
and U13350 (N_13350,N_8458,N_9941);
or U13351 (N_13351,N_5533,N_7428);
nand U13352 (N_13352,N_7300,N_7871);
nor U13353 (N_13353,N_9046,N_7486);
nand U13354 (N_13354,N_8566,N_7641);
nor U13355 (N_13355,N_6009,N_9967);
or U13356 (N_13356,N_6044,N_9730);
or U13357 (N_13357,N_7151,N_8571);
or U13358 (N_13358,N_5717,N_5578);
or U13359 (N_13359,N_8676,N_9172);
and U13360 (N_13360,N_6580,N_9330);
or U13361 (N_13361,N_5423,N_7146);
or U13362 (N_13362,N_6991,N_8736);
or U13363 (N_13363,N_6670,N_7027);
nand U13364 (N_13364,N_8843,N_5032);
nand U13365 (N_13365,N_8859,N_8928);
and U13366 (N_13366,N_8215,N_6791);
nor U13367 (N_13367,N_7114,N_6557);
or U13368 (N_13368,N_8921,N_9458);
and U13369 (N_13369,N_6507,N_7003);
or U13370 (N_13370,N_8948,N_7654);
nor U13371 (N_13371,N_8367,N_7388);
and U13372 (N_13372,N_5122,N_5988);
and U13373 (N_13373,N_6466,N_6354);
nor U13374 (N_13374,N_8832,N_7410);
and U13375 (N_13375,N_6626,N_5670);
nor U13376 (N_13376,N_9789,N_5729);
nor U13377 (N_13377,N_6978,N_9634);
or U13378 (N_13378,N_5557,N_5771);
nand U13379 (N_13379,N_8862,N_7427);
nand U13380 (N_13380,N_8956,N_9068);
nor U13381 (N_13381,N_5581,N_5381);
or U13382 (N_13382,N_8372,N_6516);
nor U13383 (N_13383,N_9347,N_5824);
nor U13384 (N_13384,N_7268,N_6959);
or U13385 (N_13385,N_6602,N_6300);
nor U13386 (N_13386,N_8175,N_7020);
nand U13387 (N_13387,N_7130,N_8390);
nand U13388 (N_13388,N_5666,N_6545);
nor U13389 (N_13389,N_9345,N_8467);
or U13390 (N_13390,N_7118,N_6310);
xor U13391 (N_13391,N_6416,N_8570);
nand U13392 (N_13392,N_5336,N_5432);
nor U13393 (N_13393,N_7311,N_6786);
nand U13394 (N_13394,N_6120,N_5312);
nand U13395 (N_13395,N_9983,N_5994);
nand U13396 (N_13396,N_6410,N_9245);
and U13397 (N_13397,N_6282,N_6521);
nand U13398 (N_13398,N_9658,N_9870);
or U13399 (N_13399,N_9593,N_5452);
nand U13400 (N_13400,N_7998,N_7594);
nor U13401 (N_13401,N_9456,N_5406);
and U13402 (N_13402,N_8398,N_6653);
nand U13403 (N_13403,N_9882,N_8081);
and U13404 (N_13404,N_8504,N_7346);
nor U13405 (N_13405,N_6098,N_6389);
nor U13406 (N_13406,N_9064,N_7778);
nor U13407 (N_13407,N_8499,N_8135);
or U13408 (N_13408,N_9231,N_7793);
and U13409 (N_13409,N_7490,N_9109);
or U13410 (N_13410,N_7886,N_9851);
or U13411 (N_13411,N_6181,N_8452);
nor U13412 (N_13412,N_9536,N_7085);
or U13413 (N_13413,N_6529,N_7120);
nor U13414 (N_13414,N_8541,N_5854);
or U13415 (N_13415,N_5917,N_7279);
or U13416 (N_13416,N_8788,N_8656);
and U13417 (N_13417,N_8014,N_8629);
nand U13418 (N_13418,N_5669,N_8582);
nor U13419 (N_13419,N_9340,N_8846);
nor U13420 (N_13420,N_6002,N_6527);
and U13421 (N_13421,N_7091,N_8226);
nand U13422 (N_13422,N_5010,N_7686);
and U13423 (N_13423,N_9208,N_9738);
or U13424 (N_13424,N_5743,N_6890);
nor U13425 (N_13425,N_8548,N_6311);
or U13426 (N_13426,N_7298,N_5764);
nand U13427 (N_13427,N_9694,N_7315);
or U13428 (N_13428,N_8996,N_8907);
nand U13429 (N_13429,N_7124,N_5249);
nor U13430 (N_13430,N_9468,N_5362);
and U13431 (N_13431,N_6317,N_7784);
or U13432 (N_13432,N_8620,N_7084);
or U13433 (N_13433,N_7453,N_6847);
or U13434 (N_13434,N_9989,N_6435);
or U13435 (N_13435,N_8988,N_7946);
nand U13436 (N_13436,N_9769,N_5389);
nor U13437 (N_13437,N_7790,N_6917);
or U13438 (N_13438,N_9469,N_5266);
and U13439 (N_13439,N_5378,N_6890);
and U13440 (N_13440,N_5482,N_9886);
nor U13441 (N_13441,N_8985,N_5145);
xor U13442 (N_13442,N_8508,N_7962);
nand U13443 (N_13443,N_5686,N_8087);
and U13444 (N_13444,N_6120,N_8138);
or U13445 (N_13445,N_6882,N_5795);
and U13446 (N_13446,N_5316,N_6479);
or U13447 (N_13447,N_9138,N_8953);
nand U13448 (N_13448,N_5755,N_7009);
or U13449 (N_13449,N_9400,N_9773);
nand U13450 (N_13450,N_6908,N_7656);
nor U13451 (N_13451,N_8962,N_6893);
or U13452 (N_13452,N_8276,N_8267);
nand U13453 (N_13453,N_5720,N_8781);
nand U13454 (N_13454,N_8244,N_5085);
nor U13455 (N_13455,N_6799,N_5347);
or U13456 (N_13456,N_7803,N_9278);
nor U13457 (N_13457,N_7455,N_9415);
nand U13458 (N_13458,N_8041,N_9646);
and U13459 (N_13459,N_5581,N_9743);
or U13460 (N_13460,N_6841,N_5832);
and U13461 (N_13461,N_5996,N_5527);
nor U13462 (N_13462,N_9391,N_9818);
and U13463 (N_13463,N_9865,N_7196);
nor U13464 (N_13464,N_5995,N_7296);
nand U13465 (N_13465,N_8253,N_8993);
xnor U13466 (N_13466,N_5487,N_5106);
and U13467 (N_13467,N_9522,N_9066);
and U13468 (N_13468,N_9289,N_7453);
nand U13469 (N_13469,N_6441,N_6163);
and U13470 (N_13470,N_6332,N_5464);
or U13471 (N_13471,N_9653,N_8260);
nor U13472 (N_13472,N_9627,N_7023);
and U13473 (N_13473,N_7687,N_5555);
nand U13474 (N_13474,N_9780,N_9398);
or U13475 (N_13475,N_8146,N_5926);
and U13476 (N_13476,N_7162,N_5146);
nand U13477 (N_13477,N_9248,N_9402);
nand U13478 (N_13478,N_6854,N_9570);
or U13479 (N_13479,N_8439,N_6202);
nor U13480 (N_13480,N_8688,N_8915);
and U13481 (N_13481,N_9144,N_6044);
nand U13482 (N_13482,N_5873,N_9163);
nor U13483 (N_13483,N_8394,N_7049);
and U13484 (N_13484,N_9952,N_6823);
nand U13485 (N_13485,N_8998,N_9737);
nor U13486 (N_13486,N_5512,N_7486);
nor U13487 (N_13487,N_9033,N_7122);
or U13488 (N_13488,N_8212,N_6086);
and U13489 (N_13489,N_6987,N_7768);
or U13490 (N_13490,N_8837,N_8967);
nand U13491 (N_13491,N_6308,N_7943);
nand U13492 (N_13492,N_8590,N_8105);
nor U13493 (N_13493,N_9994,N_5554);
nor U13494 (N_13494,N_7620,N_6894);
or U13495 (N_13495,N_6316,N_7744);
nand U13496 (N_13496,N_5661,N_8247);
nand U13497 (N_13497,N_8189,N_7651);
and U13498 (N_13498,N_9980,N_8076);
nand U13499 (N_13499,N_7081,N_9275);
and U13500 (N_13500,N_6807,N_9464);
nand U13501 (N_13501,N_7919,N_6324);
nor U13502 (N_13502,N_8733,N_6763);
or U13503 (N_13503,N_9521,N_6491);
and U13504 (N_13504,N_5760,N_5795);
nand U13505 (N_13505,N_7409,N_6687);
and U13506 (N_13506,N_7129,N_8377);
and U13507 (N_13507,N_7508,N_5321);
or U13508 (N_13508,N_8317,N_9634);
xor U13509 (N_13509,N_8203,N_7405);
and U13510 (N_13510,N_8758,N_5242);
and U13511 (N_13511,N_5608,N_9396);
and U13512 (N_13512,N_7342,N_5201);
nor U13513 (N_13513,N_6571,N_9977);
or U13514 (N_13514,N_8519,N_7371);
and U13515 (N_13515,N_9523,N_8845);
or U13516 (N_13516,N_9720,N_5241);
and U13517 (N_13517,N_7536,N_5912);
or U13518 (N_13518,N_8203,N_6989);
nand U13519 (N_13519,N_8520,N_5011);
or U13520 (N_13520,N_8083,N_5858);
or U13521 (N_13521,N_8607,N_6996);
and U13522 (N_13522,N_9015,N_7244);
nor U13523 (N_13523,N_7428,N_6310);
or U13524 (N_13524,N_7963,N_7266);
and U13525 (N_13525,N_8130,N_5433);
xnor U13526 (N_13526,N_6175,N_7398);
nand U13527 (N_13527,N_7873,N_8679);
nand U13528 (N_13528,N_6105,N_5783);
nand U13529 (N_13529,N_6811,N_5008);
nor U13530 (N_13530,N_7814,N_7345);
and U13531 (N_13531,N_7426,N_7417);
nand U13532 (N_13532,N_5049,N_5720);
nor U13533 (N_13533,N_9184,N_9657);
nor U13534 (N_13534,N_9998,N_8676);
and U13535 (N_13535,N_6559,N_5200);
or U13536 (N_13536,N_5828,N_7415);
nor U13537 (N_13537,N_8407,N_8632);
and U13538 (N_13538,N_5794,N_7433);
or U13539 (N_13539,N_7961,N_7683);
xor U13540 (N_13540,N_9266,N_7838);
xnor U13541 (N_13541,N_8416,N_5953);
nand U13542 (N_13542,N_8085,N_7496);
nand U13543 (N_13543,N_9680,N_6217);
or U13544 (N_13544,N_5892,N_8012);
xor U13545 (N_13545,N_6088,N_8234);
nand U13546 (N_13546,N_5163,N_8589);
and U13547 (N_13547,N_7384,N_6400);
nand U13548 (N_13548,N_8443,N_5771);
nand U13549 (N_13549,N_5517,N_8633);
and U13550 (N_13550,N_6162,N_9816);
or U13551 (N_13551,N_8868,N_8181);
or U13552 (N_13552,N_5839,N_6251);
and U13553 (N_13553,N_8033,N_8626);
nand U13554 (N_13554,N_6626,N_9931);
nand U13555 (N_13555,N_5358,N_5484);
nand U13556 (N_13556,N_9774,N_9514);
nand U13557 (N_13557,N_8477,N_5392);
nand U13558 (N_13558,N_5574,N_6104);
or U13559 (N_13559,N_7484,N_7928);
xor U13560 (N_13560,N_9269,N_7906);
nand U13561 (N_13561,N_9365,N_7042);
and U13562 (N_13562,N_5246,N_7601);
and U13563 (N_13563,N_8757,N_5678);
nand U13564 (N_13564,N_5948,N_6397);
xnor U13565 (N_13565,N_5372,N_9589);
nor U13566 (N_13566,N_6656,N_8994);
and U13567 (N_13567,N_9393,N_6807);
and U13568 (N_13568,N_8028,N_9584);
or U13569 (N_13569,N_7489,N_8760);
xnor U13570 (N_13570,N_6968,N_5732);
or U13571 (N_13571,N_8081,N_5698);
nor U13572 (N_13572,N_9947,N_9114);
and U13573 (N_13573,N_7348,N_6822);
nand U13574 (N_13574,N_9715,N_8102);
nand U13575 (N_13575,N_5188,N_7479);
nand U13576 (N_13576,N_7185,N_5239);
nor U13577 (N_13577,N_8465,N_7350);
nand U13578 (N_13578,N_6850,N_8493);
nand U13579 (N_13579,N_6180,N_6203);
and U13580 (N_13580,N_5396,N_7039);
nor U13581 (N_13581,N_5295,N_6411);
and U13582 (N_13582,N_9910,N_7870);
nand U13583 (N_13583,N_6412,N_6678);
nor U13584 (N_13584,N_5279,N_5318);
nor U13585 (N_13585,N_5286,N_8457);
and U13586 (N_13586,N_9265,N_8974);
and U13587 (N_13587,N_9435,N_7812);
nand U13588 (N_13588,N_7740,N_7362);
or U13589 (N_13589,N_9841,N_5001);
and U13590 (N_13590,N_6519,N_7160);
nor U13591 (N_13591,N_6873,N_6492);
nand U13592 (N_13592,N_7660,N_5263);
and U13593 (N_13593,N_9889,N_7927);
nand U13594 (N_13594,N_8301,N_7140);
nor U13595 (N_13595,N_8683,N_7324);
or U13596 (N_13596,N_5436,N_7183);
nor U13597 (N_13597,N_9588,N_8842);
nand U13598 (N_13598,N_7796,N_7216);
and U13599 (N_13599,N_9013,N_7377);
and U13600 (N_13600,N_7146,N_7167);
and U13601 (N_13601,N_8174,N_9940);
nor U13602 (N_13602,N_6161,N_7770);
nand U13603 (N_13603,N_8209,N_9646);
nor U13604 (N_13604,N_5308,N_7790);
nand U13605 (N_13605,N_9240,N_9342);
or U13606 (N_13606,N_5924,N_9770);
or U13607 (N_13607,N_5296,N_5587);
nand U13608 (N_13608,N_9746,N_5370);
and U13609 (N_13609,N_5611,N_5292);
and U13610 (N_13610,N_8284,N_5028);
or U13611 (N_13611,N_5729,N_7729);
or U13612 (N_13612,N_9038,N_6285);
nand U13613 (N_13613,N_6034,N_6088);
nor U13614 (N_13614,N_9974,N_7792);
and U13615 (N_13615,N_5229,N_6069);
and U13616 (N_13616,N_5369,N_6985);
nor U13617 (N_13617,N_8408,N_8067);
and U13618 (N_13618,N_9879,N_7248);
or U13619 (N_13619,N_7649,N_8141);
and U13620 (N_13620,N_7618,N_9081);
nor U13621 (N_13621,N_7223,N_7435);
or U13622 (N_13622,N_5639,N_5995);
nand U13623 (N_13623,N_5840,N_7929);
nand U13624 (N_13624,N_7918,N_7195);
or U13625 (N_13625,N_5609,N_5597);
nand U13626 (N_13626,N_9478,N_9645);
nor U13627 (N_13627,N_6286,N_8234);
nor U13628 (N_13628,N_9464,N_5719);
nor U13629 (N_13629,N_7952,N_7185);
nor U13630 (N_13630,N_9363,N_7244);
nand U13631 (N_13631,N_8961,N_5916);
nor U13632 (N_13632,N_7887,N_7013);
nor U13633 (N_13633,N_7598,N_7145);
and U13634 (N_13634,N_9697,N_5368);
nor U13635 (N_13635,N_8974,N_6082);
nand U13636 (N_13636,N_7994,N_8544);
nand U13637 (N_13637,N_6270,N_7900);
and U13638 (N_13638,N_6575,N_9330);
nor U13639 (N_13639,N_5942,N_9214);
nand U13640 (N_13640,N_9155,N_5261);
nor U13641 (N_13641,N_7900,N_8553);
and U13642 (N_13642,N_9051,N_7601);
and U13643 (N_13643,N_6300,N_6288);
nor U13644 (N_13644,N_5450,N_5433);
xor U13645 (N_13645,N_8764,N_5958);
nor U13646 (N_13646,N_9384,N_5598);
nand U13647 (N_13647,N_5201,N_5613);
nand U13648 (N_13648,N_7372,N_9398);
or U13649 (N_13649,N_5150,N_7515);
and U13650 (N_13650,N_8772,N_8655);
or U13651 (N_13651,N_8882,N_9130);
and U13652 (N_13652,N_9708,N_6969);
and U13653 (N_13653,N_5337,N_5808);
or U13654 (N_13654,N_6124,N_5663);
nor U13655 (N_13655,N_5507,N_6334);
or U13656 (N_13656,N_7486,N_5844);
and U13657 (N_13657,N_8747,N_8961);
or U13658 (N_13658,N_8379,N_8380);
or U13659 (N_13659,N_6247,N_5567);
or U13660 (N_13660,N_7694,N_7238);
and U13661 (N_13661,N_8614,N_6022);
nor U13662 (N_13662,N_5745,N_8993);
or U13663 (N_13663,N_7474,N_6960);
and U13664 (N_13664,N_5384,N_5252);
or U13665 (N_13665,N_6567,N_5318);
and U13666 (N_13666,N_7060,N_9001);
nor U13667 (N_13667,N_7538,N_9590);
or U13668 (N_13668,N_9605,N_5429);
and U13669 (N_13669,N_9024,N_6375);
nand U13670 (N_13670,N_7187,N_5478);
or U13671 (N_13671,N_8138,N_7538);
and U13672 (N_13672,N_7773,N_5022);
and U13673 (N_13673,N_7787,N_7117);
nor U13674 (N_13674,N_6890,N_8650);
or U13675 (N_13675,N_7015,N_8613);
and U13676 (N_13676,N_8629,N_8885);
or U13677 (N_13677,N_9933,N_6574);
nand U13678 (N_13678,N_7869,N_6270);
and U13679 (N_13679,N_5440,N_8092);
nand U13680 (N_13680,N_7147,N_7874);
and U13681 (N_13681,N_7940,N_9654);
nand U13682 (N_13682,N_5679,N_8861);
xnor U13683 (N_13683,N_8464,N_9862);
and U13684 (N_13684,N_5436,N_9400);
and U13685 (N_13685,N_9715,N_6784);
or U13686 (N_13686,N_8624,N_6136);
or U13687 (N_13687,N_6168,N_9542);
or U13688 (N_13688,N_7248,N_6422);
or U13689 (N_13689,N_8524,N_5845);
nor U13690 (N_13690,N_5167,N_5131);
and U13691 (N_13691,N_6521,N_5162);
and U13692 (N_13692,N_5434,N_5074);
and U13693 (N_13693,N_8217,N_7117);
nor U13694 (N_13694,N_9848,N_6232);
and U13695 (N_13695,N_5907,N_5680);
nor U13696 (N_13696,N_6329,N_7504);
nor U13697 (N_13697,N_5903,N_5365);
nor U13698 (N_13698,N_6339,N_8589);
nand U13699 (N_13699,N_5998,N_7612);
or U13700 (N_13700,N_9752,N_5063);
or U13701 (N_13701,N_8345,N_5351);
nand U13702 (N_13702,N_7152,N_7426);
nand U13703 (N_13703,N_5239,N_5442);
or U13704 (N_13704,N_6610,N_5471);
and U13705 (N_13705,N_6898,N_9219);
nand U13706 (N_13706,N_9549,N_6645);
xnor U13707 (N_13707,N_5150,N_7218);
nand U13708 (N_13708,N_9005,N_8532);
nand U13709 (N_13709,N_8232,N_7172);
or U13710 (N_13710,N_5389,N_6043);
and U13711 (N_13711,N_6193,N_8998);
nor U13712 (N_13712,N_9396,N_7165);
or U13713 (N_13713,N_9045,N_9807);
nor U13714 (N_13714,N_9881,N_5494);
or U13715 (N_13715,N_7871,N_8933);
nand U13716 (N_13716,N_8525,N_8857);
and U13717 (N_13717,N_8856,N_9914);
nor U13718 (N_13718,N_6278,N_8022);
or U13719 (N_13719,N_9046,N_8135);
and U13720 (N_13720,N_9762,N_6335);
and U13721 (N_13721,N_9049,N_9527);
or U13722 (N_13722,N_6419,N_5169);
and U13723 (N_13723,N_7666,N_8144);
and U13724 (N_13724,N_9766,N_6806);
or U13725 (N_13725,N_8318,N_6435);
or U13726 (N_13726,N_5890,N_5234);
nor U13727 (N_13727,N_8326,N_7904);
nand U13728 (N_13728,N_8374,N_8528);
nand U13729 (N_13729,N_5308,N_7075);
nor U13730 (N_13730,N_8117,N_5601);
nand U13731 (N_13731,N_5472,N_9992);
nand U13732 (N_13732,N_9178,N_5455);
nor U13733 (N_13733,N_9276,N_5340);
nor U13734 (N_13734,N_7676,N_7267);
or U13735 (N_13735,N_6923,N_8247);
or U13736 (N_13736,N_8265,N_7140);
xor U13737 (N_13737,N_9536,N_7059);
or U13738 (N_13738,N_6706,N_7502);
xor U13739 (N_13739,N_5087,N_5132);
and U13740 (N_13740,N_6995,N_6818);
nand U13741 (N_13741,N_7455,N_7850);
xor U13742 (N_13742,N_9851,N_7827);
nand U13743 (N_13743,N_8527,N_9352);
nor U13744 (N_13744,N_5018,N_8654);
or U13745 (N_13745,N_5261,N_8981);
nor U13746 (N_13746,N_9363,N_8867);
nor U13747 (N_13747,N_7091,N_6834);
and U13748 (N_13748,N_6525,N_9415);
and U13749 (N_13749,N_8261,N_7965);
and U13750 (N_13750,N_7565,N_8077);
nor U13751 (N_13751,N_6560,N_9810);
or U13752 (N_13752,N_6868,N_6878);
and U13753 (N_13753,N_6907,N_9336);
nor U13754 (N_13754,N_6905,N_7059);
or U13755 (N_13755,N_5890,N_8333);
and U13756 (N_13756,N_5573,N_5405);
or U13757 (N_13757,N_9124,N_9108);
nand U13758 (N_13758,N_9185,N_7343);
nand U13759 (N_13759,N_6552,N_8562);
and U13760 (N_13760,N_7554,N_8962);
or U13761 (N_13761,N_7329,N_8919);
nor U13762 (N_13762,N_7688,N_9927);
or U13763 (N_13763,N_6519,N_8229);
nand U13764 (N_13764,N_9013,N_9813);
nor U13765 (N_13765,N_8985,N_6524);
xor U13766 (N_13766,N_7325,N_9739);
and U13767 (N_13767,N_8461,N_9190);
nand U13768 (N_13768,N_5608,N_6353);
or U13769 (N_13769,N_6739,N_8248);
and U13770 (N_13770,N_5642,N_9436);
nor U13771 (N_13771,N_7398,N_9735);
and U13772 (N_13772,N_7245,N_5635);
or U13773 (N_13773,N_7179,N_5194);
and U13774 (N_13774,N_5131,N_8835);
nand U13775 (N_13775,N_9845,N_9599);
and U13776 (N_13776,N_5318,N_9206);
or U13777 (N_13777,N_7600,N_8977);
or U13778 (N_13778,N_9935,N_5091);
nand U13779 (N_13779,N_7964,N_5648);
or U13780 (N_13780,N_6106,N_9263);
nor U13781 (N_13781,N_6636,N_9374);
nor U13782 (N_13782,N_5771,N_7494);
nor U13783 (N_13783,N_7585,N_8047);
xor U13784 (N_13784,N_6396,N_7424);
nand U13785 (N_13785,N_9014,N_5451);
xor U13786 (N_13786,N_8359,N_5266);
and U13787 (N_13787,N_8292,N_6362);
nand U13788 (N_13788,N_6233,N_6205);
nand U13789 (N_13789,N_5519,N_7185);
and U13790 (N_13790,N_6516,N_6988);
nor U13791 (N_13791,N_8782,N_9920);
nand U13792 (N_13792,N_8765,N_7472);
or U13793 (N_13793,N_8295,N_9525);
xor U13794 (N_13794,N_7548,N_8840);
nor U13795 (N_13795,N_6166,N_5114);
and U13796 (N_13796,N_8461,N_8584);
and U13797 (N_13797,N_7757,N_9536);
or U13798 (N_13798,N_9562,N_6118);
or U13799 (N_13799,N_6921,N_5661);
nand U13800 (N_13800,N_8713,N_6079);
or U13801 (N_13801,N_9049,N_5380);
and U13802 (N_13802,N_9239,N_9491);
or U13803 (N_13803,N_7463,N_9381);
nor U13804 (N_13804,N_9105,N_8705);
nand U13805 (N_13805,N_7585,N_7136);
nor U13806 (N_13806,N_9668,N_9491);
nor U13807 (N_13807,N_5107,N_6549);
nand U13808 (N_13808,N_9927,N_5737);
nand U13809 (N_13809,N_8120,N_6044);
nand U13810 (N_13810,N_7084,N_6311);
and U13811 (N_13811,N_9818,N_9777);
and U13812 (N_13812,N_8906,N_9395);
and U13813 (N_13813,N_5932,N_7775);
and U13814 (N_13814,N_8057,N_6829);
nand U13815 (N_13815,N_7984,N_6318);
nor U13816 (N_13816,N_9213,N_9359);
and U13817 (N_13817,N_8422,N_6261);
or U13818 (N_13818,N_5568,N_7124);
nor U13819 (N_13819,N_7861,N_8243);
or U13820 (N_13820,N_6079,N_9308);
and U13821 (N_13821,N_5790,N_9824);
nor U13822 (N_13822,N_6875,N_7829);
nand U13823 (N_13823,N_8074,N_7342);
nor U13824 (N_13824,N_5179,N_9989);
nor U13825 (N_13825,N_7216,N_7837);
nand U13826 (N_13826,N_9337,N_6878);
and U13827 (N_13827,N_7677,N_7495);
and U13828 (N_13828,N_5620,N_6808);
or U13829 (N_13829,N_8961,N_7091);
xor U13830 (N_13830,N_7492,N_9958);
nand U13831 (N_13831,N_5324,N_8316);
or U13832 (N_13832,N_9279,N_5671);
xnor U13833 (N_13833,N_6976,N_7526);
or U13834 (N_13834,N_5795,N_7955);
and U13835 (N_13835,N_5270,N_6711);
nand U13836 (N_13836,N_9422,N_9434);
nand U13837 (N_13837,N_7029,N_5354);
nand U13838 (N_13838,N_6888,N_9671);
nand U13839 (N_13839,N_8847,N_8030);
and U13840 (N_13840,N_7926,N_8976);
and U13841 (N_13841,N_5417,N_7878);
nor U13842 (N_13842,N_7720,N_8679);
nor U13843 (N_13843,N_7237,N_6177);
or U13844 (N_13844,N_7624,N_6563);
nor U13845 (N_13845,N_7377,N_8142);
or U13846 (N_13846,N_5635,N_5517);
nor U13847 (N_13847,N_5298,N_9793);
and U13848 (N_13848,N_9960,N_6114);
nor U13849 (N_13849,N_5290,N_6477);
nor U13850 (N_13850,N_6145,N_6356);
nor U13851 (N_13851,N_6930,N_9016);
nand U13852 (N_13852,N_5324,N_5157);
and U13853 (N_13853,N_9028,N_8279);
nor U13854 (N_13854,N_7898,N_7110);
nand U13855 (N_13855,N_9558,N_7392);
nand U13856 (N_13856,N_5194,N_8312);
and U13857 (N_13857,N_7626,N_8143);
and U13858 (N_13858,N_7384,N_5750);
nor U13859 (N_13859,N_9468,N_8719);
and U13860 (N_13860,N_7781,N_6653);
and U13861 (N_13861,N_9431,N_7857);
nand U13862 (N_13862,N_6234,N_7340);
and U13863 (N_13863,N_9688,N_5061);
and U13864 (N_13864,N_6697,N_9927);
nor U13865 (N_13865,N_5805,N_6199);
nor U13866 (N_13866,N_7768,N_5270);
nor U13867 (N_13867,N_6831,N_9857);
nor U13868 (N_13868,N_9190,N_9750);
and U13869 (N_13869,N_8143,N_8675);
nand U13870 (N_13870,N_7206,N_6935);
and U13871 (N_13871,N_7546,N_7556);
or U13872 (N_13872,N_8214,N_9171);
and U13873 (N_13873,N_9746,N_6289);
and U13874 (N_13874,N_5530,N_7148);
nand U13875 (N_13875,N_7947,N_7438);
nor U13876 (N_13876,N_6125,N_9706);
nor U13877 (N_13877,N_7022,N_8343);
or U13878 (N_13878,N_6896,N_6383);
and U13879 (N_13879,N_8878,N_8483);
nand U13880 (N_13880,N_5513,N_9305);
nand U13881 (N_13881,N_7770,N_9063);
and U13882 (N_13882,N_9575,N_5447);
or U13883 (N_13883,N_9516,N_5136);
or U13884 (N_13884,N_8782,N_9149);
or U13885 (N_13885,N_8997,N_8625);
nor U13886 (N_13886,N_9395,N_7367);
nand U13887 (N_13887,N_8118,N_9860);
and U13888 (N_13888,N_8794,N_5608);
nor U13889 (N_13889,N_9101,N_6153);
and U13890 (N_13890,N_7479,N_5582);
nor U13891 (N_13891,N_5881,N_5299);
or U13892 (N_13892,N_8497,N_5514);
and U13893 (N_13893,N_7422,N_8278);
nand U13894 (N_13894,N_9592,N_6050);
xnor U13895 (N_13895,N_6291,N_6194);
nor U13896 (N_13896,N_9446,N_8504);
and U13897 (N_13897,N_8388,N_7054);
or U13898 (N_13898,N_8773,N_6452);
nor U13899 (N_13899,N_5353,N_9816);
or U13900 (N_13900,N_6469,N_6363);
nand U13901 (N_13901,N_6396,N_5486);
nor U13902 (N_13902,N_5268,N_5154);
nand U13903 (N_13903,N_7606,N_8008);
and U13904 (N_13904,N_7095,N_5343);
or U13905 (N_13905,N_9211,N_7191);
and U13906 (N_13906,N_9842,N_9082);
or U13907 (N_13907,N_8353,N_7048);
nor U13908 (N_13908,N_5878,N_9806);
xor U13909 (N_13909,N_9071,N_5130);
and U13910 (N_13910,N_5933,N_6341);
or U13911 (N_13911,N_9274,N_9884);
xor U13912 (N_13912,N_9707,N_8503);
and U13913 (N_13913,N_8253,N_9354);
nor U13914 (N_13914,N_5039,N_8771);
nor U13915 (N_13915,N_7569,N_7804);
nor U13916 (N_13916,N_6755,N_6715);
or U13917 (N_13917,N_6695,N_6493);
and U13918 (N_13918,N_8246,N_9721);
nor U13919 (N_13919,N_6908,N_8712);
or U13920 (N_13920,N_5155,N_8268);
nor U13921 (N_13921,N_8112,N_9690);
nor U13922 (N_13922,N_5166,N_8840);
and U13923 (N_13923,N_7267,N_7355);
nor U13924 (N_13924,N_6047,N_5578);
nor U13925 (N_13925,N_8780,N_8274);
or U13926 (N_13926,N_5733,N_8457);
nand U13927 (N_13927,N_9503,N_6846);
nand U13928 (N_13928,N_9483,N_5890);
and U13929 (N_13929,N_6285,N_6249);
nand U13930 (N_13930,N_6351,N_8648);
nor U13931 (N_13931,N_8887,N_7766);
nor U13932 (N_13932,N_6540,N_9394);
nand U13933 (N_13933,N_8831,N_5565);
and U13934 (N_13934,N_8108,N_7336);
nor U13935 (N_13935,N_9564,N_6522);
and U13936 (N_13936,N_7919,N_9017);
nor U13937 (N_13937,N_7778,N_5438);
and U13938 (N_13938,N_8938,N_8182);
nand U13939 (N_13939,N_8148,N_5714);
nand U13940 (N_13940,N_6476,N_8954);
nor U13941 (N_13941,N_9111,N_5062);
and U13942 (N_13942,N_8190,N_8152);
nor U13943 (N_13943,N_5053,N_6365);
or U13944 (N_13944,N_8456,N_7587);
nand U13945 (N_13945,N_9027,N_5598);
and U13946 (N_13946,N_8617,N_7535);
and U13947 (N_13947,N_8720,N_8582);
nand U13948 (N_13948,N_7554,N_9187);
and U13949 (N_13949,N_5098,N_8242);
and U13950 (N_13950,N_7458,N_7479);
or U13951 (N_13951,N_5503,N_8302);
nand U13952 (N_13952,N_8028,N_9525);
nor U13953 (N_13953,N_9375,N_7053);
or U13954 (N_13954,N_8770,N_8057);
or U13955 (N_13955,N_6681,N_6719);
nand U13956 (N_13956,N_9441,N_8901);
nor U13957 (N_13957,N_8381,N_6936);
nor U13958 (N_13958,N_9024,N_6606);
nand U13959 (N_13959,N_7455,N_7156);
or U13960 (N_13960,N_6419,N_5205);
and U13961 (N_13961,N_5986,N_5068);
and U13962 (N_13962,N_6595,N_9939);
or U13963 (N_13963,N_6047,N_8135);
nor U13964 (N_13964,N_5172,N_6651);
nand U13965 (N_13965,N_6306,N_8223);
and U13966 (N_13966,N_7039,N_5515);
or U13967 (N_13967,N_5644,N_5913);
and U13968 (N_13968,N_9177,N_7404);
or U13969 (N_13969,N_8819,N_5891);
nor U13970 (N_13970,N_9452,N_6280);
or U13971 (N_13971,N_5988,N_6854);
nor U13972 (N_13972,N_9158,N_9213);
nor U13973 (N_13973,N_6324,N_9517);
nor U13974 (N_13974,N_8255,N_8834);
or U13975 (N_13975,N_7015,N_5267);
nor U13976 (N_13976,N_8665,N_8729);
nand U13977 (N_13977,N_7411,N_8007);
nor U13978 (N_13978,N_5043,N_7562);
nor U13979 (N_13979,N_9141,N_5711);
and U13980 (N_13980,N_5994,N_7117);
and U13981 (N_13981,N_6072,N_7198);
nor U13982 (N_13982,N_9181,N_9969);
and U13983 (N_13983,N_6389,N_6715);
nand U13984 (N_13984,N_7991,N_5806);
xnor U13985 (N_13985,N_7012,N_8129);
nor U13986 (N_13986,N_8595,N_8487);
or U13987 (N_13987,N_9611,N_9652);
nand U13988 (N_13988,N_9485,N_5506);
xnor U13989 (N_13989,N_6816,N_8800);
nor U13990 (N_13990,N_6691,N_5014);
nor U13991 (N_13991,N_7082,N_8644);
nor U13992 (N_13992,N_6663,N_9891);
and U13993 (N_13993,N_8287,N_9711);
nand U13994 (N_13994,N_6473,N_6855);
and U13995 (N_13995,N_8423,N_9276);
nand U13996 (N_13996,N_5305,N_7193);
and U13997 (N_13997,N_7978,N_6693);
nand U13998 (N_13998,N_5013,N_9075);
nor U13999 (N_13999,N_8891,N_9681);
or U14000 (N_14000,N_5204,N_7748);
and U14001 (N_14001,N_8871,N_5000);
nor U14002 (N_14002,N_5727,N_6241);
or U14003 (N_14003,N_5318,N_7120);
nor U14004 (N_14004,N_8197,N_8234);
nand U14005 (N_14005,N_6607,N_8501);
nand U14006 (N_14006,N_8497,N_8162);
and U14007 (N_14007,N_8648,N_6930);
nor U14008 (N_14008,N_8288,N_9789);
or U14009 (N_14009,N_6128,N_6631);
nand U14010 (N_14010,N_8431,N_6731);
nand U14011 (N_14011,N_9391,N_5054);
nor U14012 (N_14012,N_9106,N_6047);
nand U14013 (N_14013,N_7489,N_9404);
nand U14014 (N_14014,N_6346,N_9233);
nand U14015 (N_14015,N_8048,N_8892);
nor U14016 (N_14016,N_5948,N_5081);
nor U14017 (N_14017,N_7387,N_5085);
or U14018 (N_14018,N_6110,N_6010);
and U14019 (N_14019,N_7988,N_7829);
nor U14020 (N_14020,N_8466,N_8883);
nor U14021 (N_14021,N_8012,N_9925);
nand U14022 (N_14022,N_5511,N_8486);
nor U14023 (N_14023,N_7619,N_6156);
and U14024 (N_14024,N_7198,N_5097);
and U14025 (N_14025,N_7948,N_8530);
or U14026 (N_14026,N_7332,N_8994);
nand U14027 (N_14027,N_5461,N_6628);
nand U14028 (N_14028,N_8793,N_6606);
nor U14029 (N_14029,N_6268,N_6984);
nand U14030 (N_14030,N_7248,N_9606);
nor U14031 (N_14031,N_6405,N_7166);
nand U14032 (N_14032,N_6007,N_6913);
and U14033 (N_14033,N_5879,N_7663);
or U14034 (N_14034,N_5988,N_9473);
or U14035 (N_14035,N_7278,N_5250);
or U14036 (N_14036,N_5674,N_9098);
or U14037 (N_14037,N_9441,N_8287);
or U14038 (N_14038,N_7844,N_9102);
nor U14039 (N_14039,N_7845,N_9505);
and U14040 (N_14040,N_5657,N_5623);
nor U14041 (N_14041,N_5638,N_9307);
or U14042 (N_14042,N_7638,N_6558);
nand U14043 (N_14043,N_5223,N_9010);
or U14044 (N_14044,N_5810,N_5050);
xor U14045 (N_14045,N_7070,N_8554);
nor U14046 (N_14046,N_6799,N_6132);
nor U14047 (N_14047,N_9937,N_5041);
or U14048 (N_14048,N_8309,N_6225);
xor U14049 (N_14049,N_8475,N_9231);
nand U14050 (N_14050,N_5649,N_8164);
nand U14051 (N_14051,N_9983,N_6175);
nor U14052 (N_14052,N_8663,N_9595);
or U14053 (N_14053,N_8140,N_7313);
nand U14054 (N_14054,N_5659,N_9833);
or U14055 (N_14055,N_9393,N_9704);
nand U14056 (N_14056,N_5245,N_5234);
nor U14057 (N_14057,N_7277,N_8006);
and U14058 (N_14058,N_6787,N_7505);
nand U14059 (N_14059,N_7037,N_8984);
nand U14060 (N_14060,N_9178,N_5407);
or U14061 (N_14061,N_5378,N_6473);
nor U14062 (N_14062,N_5151,N_7162);
nand U14063 (N_14063,N_7817,N_6333);
nor U14064 (N_14064,N_6842,N_6585);
and U14065 (N_14065,N_9601,N_9577);
or U14066 (N_14066,N_8617,N_5226);
nand U14067 (N_14067,N_5520,N_9493);
or U14068 (N_14068,N_9095,N_7964);
nor U14069 (N_14069,N_7201,N_7239);
and U14070 (N_14070,N_6567,N_5649);
and U14071 (N_14071,N_5655,N_6305);
and U14072 (N_14072,N_7828,N_6120);
nor U14073 (N_14073,N_5396,N_7016);
nor U14074 (N_14074,N_8439,N_5392);
and U14075 (N_14075,N_6301,N_5641);
nand U14076 (N_14076,N_7632,N_8696);
nor U14077 (N_14077,N_8249,N_8609);
and U14078 (N_14078,N_5066,N_5087);
or U14079 (N_14079,N_7590,N_6907);
or U14080 (N_14080,N_5720,N_7373);
or U14081 (N_14081,N_7068,N_9386);
or U14082 (N_14082,N_6227,N_6476);
nor U14083 (N_14083,N_6947,N_5427);
nor U14084 (N_14084,N_7408,N_8798);
nand U14085 (N_14085,N_8809,N_7539);
and U14086 (N_14086,N_9833,N_9260);
and U14087 (N_14087,N_6235,N_6117);
or U14088 (N_14088,N_5349,N_9394);
nor U14089 (N_14089,N_8949,N_8341);
or U14090 (N_14090,N_6358,N_6901);
xnor U14091 (N_14091,N_6815,N_5332);
nand U14092 (N_14092,N_7992,N_9740);
nor U14093 (N_14093,N_6050,N_7612);
nand U14094 (N_14094,N_8467,N_7151);
nand U14095 (N_14095,N_8898,N_7644);
or U14096 (N_14096,N_7636,N_6701);
or U14097 (N_14097,N_7353,N_6677);
or U14098 (N_14098,N_9177,N_8793);
nor U14099 (N_14099,N_8365,N_5140);
or U14100 (N_14100,N_7000,N_5754);
and U14101 (N_14101,N_7179,N_8577);
nand U14102 (N_14102,N_9305,N_8900);
and U14103 (N_14103,N_8888,N_7676);
nand U14104 (N_14104,N_7338,N_9756);
and U14105 (N_14105,N_9137,N_8738);
and U14106 (N_14106,N_7304,N_7778);
or U14107 (N_14107,N_7524,N_9327);
or U14108 (N_14108,N_5424,N_6249);
or U14109 (N_14109,N_5096,N_5172);
and U14110 (N_14110,N_5943,N_6593);
or U14111 (N_14111,N_8416,N_5128);
or U14112 (N_14112,N_8333,N_7812);
or U14113 (N_14113,N_7616,N_8467);
and U14114 (N_14114,N_6413,N_7592);
or U14115 (N_14115,N_8751,N_5351);
nor U14116 (N_14116,N_6715,N_9632);
or U14117 (N_14117,N_8511,N_7793);
nor U14118 (N_14118,N_5102,N_7665);
nand U14119 (N_14119,N_9720,N_5901);
nor U14120 (N_14120,N_6535,N_5525);
and U14121 (N_14121,N_9711,N_7072);
or U14122 (N_14122,N_6409,N_7876);
nor U14123 (N_14123,N_9734,N_6345);
nand U14124 (N_14124,N_5864,N_5069);
nand U14125 (N_14125,N_7624,N_6209);
xnor U14126 (N_14126,N_6096,N_5049);
nor U14127 (N_14127,N_9205,N_9766);
or U14128 (N_14128,N_9009,N_8648);
nand U14129 (N_14129,N_6630,N_8554);
and U14130 (N_14130,N_5666,N_6011);
or U14131 (N_14131,N_9071,N_8101);
or U14132 (N_14132,N_8210,N_7942);
nor U14133 (N_14133,N_5346,N_9502);
nand U14134 (N_14134,N_6526,N_6822);
or U14135 (N_14135,N_7481,N_7714);
or U14136 (N_14136,N_5228,N_8765);
nor U14137 (N_14137,N_8289,N_5013);
and U14138 (N_14138,N_9720,N_8349);
nand U14139 (N_14139,N_5021,N_9092);
nor U14140 (N_14140,N_7825,N_9175);
nor U14141 (N_14141,N_6969,N_9794);
and U14142 (N_14142,N_5839,N_5860);
nor U14143 (N_14143,N_7809,N_9587);
nand U14144 (N_14144,N_5376,N_5206);
nor U14145 (N_14145,N_6406,N_6671);
or U14146 (N_14146,N_5933,N_8929);
or U14147 (N_14147,N_7206,N_5661);
and U14148 (N_14148,N_8440,N_9866);
and U14149 (N_14149,N_6943,N_5425);
nor U14150 (N_14150,N_5150,N_6442);
or U14151 (N_14151,N_9348,N_8851);
and U14152 (N_14152,N_5058,N_7935);
and U14153 (N_14153,N_9842,N_9694);
or U14154 (N_14154,N_6626,N_9545);
and U14155 (N_14155,N_8781,N_8297);
nor U14156 (N_14156,N_9584,N_9381);
or U14157 (N_14157,N_7608,N_8148);
or U14158 (N_14158,N_8612,N_5028);
or U14159 (N_14159,N_6745,N_9881);
or U14160 (N_14160,N_7484,N_6519);
nand U14161 (N_14161,N_6406,N_9384);
nand U14162 (N_14162,N_6834,N_7961);
xor U14163 (N_14163,N_7930,N_8059);
and U14164 (N_14164,N_8379,N_8212);
and U14165 (N_14165,N_6778,N_7636);
nand U14166 (N_14166,N_9194,N_9056);
or U14167 (N_14167,N_5046,N_6465);
nor U14168 (N_14168,N_8252,N_6655);
and U14169 (N_14169,N_5753,N_7702);
nand U14170 (N_14170,N_9526,N_9233);
and U14171 (N_14171,N_8911,N_7167);
or U14172 (N_14172,N_5403,N_9086);
nand U14173 (N_14173,N_8899,N_5525);
and U14174 (N_14174,N_9427,N_6699);
and U14175 (N_14175,N_8701,N_5363);
nand U14176 (N_14176,N_5239,N_9746);
nor U14177 (N_14177,N_5926,N_6011);
nand U14178 (N_14178,N_9953,N_7273);
or U14179 (N_14179,N_5558,N_7616);
nor U14180 (N_14180,N_6310,N_7219);
and U14181 (N_14181,N_9281,N_7981);
nor U14182 (N_14182,N_7719,N_6816);
nor U14183 (N_14183,N_9283,N_5221);
nand U14184 (N_14184,N_8769,N_5870);
nor U14185 (N_14185,N_7607,N_5741);
or U14186 (N_14186,N_7460,N_7826);
or U14187 (N_14187,N_9081,N_8729);
or U14188 (N_14188,N_5290,N_8856);
and U14189 (N_14189,N_6511,N_5553);
and U14190 (N_14190,N_6661,N_9214);
and U14191 (N_14191,N_9326,N_7428);
and U14192 (N_14192,N_6612,N_8543);
nand U14193 (N_14193,N_7518,N_8529);
nand U14194 (N_14194,N_7104,N_8928);
nor U14195 (N_14195,N_5782,N_8683);
nand U14196 (N_14196,N_7216,N_6415);
nand U14197 (N_14197,N_9915,N_5489);
and U14198 (N_14198,N_6257,N_5168);
or U14199 (N_14199,N_6147,N_7921);
and U14200 (N_14200,N_5543,N_6355);
nand U14201 (N_14201,N_5821,N_5586);
and U14202 (N_14202,N_9545,N_9686);
and U14203 (N_14203,N_8085,N_8641);
nand U14204 (N_14204,N_9219,N_5287);
nand U14205 (N_14205,N_7434,N_7760);
and U14206 (N_14206,N_9070,N_5104);
or U14207 (N_14207,N_7974,N_6201);
nand U14208 (N_14208,N_9458,N_7041);
nor U14209 (N_14209,N_6511,N_5152);
and U14210 (N_14210,N_5159,N_5581);
nand U14211 (N_14211,N_6913,N_7984);
or U14212 (N_14212,N_9531,N_5081);
and U14213 (N_14213,N_8632,N_8192);
and U14214 (N_14214,N_8695,N_9840);
xnor U14215 (N_14215,N_8801,N_8218);
nand U14216 (N_14216,N_5265,N_8666);
and U14217 (N_14217,N_6421,N_7332);
nor U14218 (N_14218,N_6223,N_5475);
or U14219 (N_14219,N_5991,N_5039);
and U14220 (N_14220,N_7550,N_9668);
nor U14221 (N_14221,N_6598,N_5347);
or U14222 (N_14222,N_9211,N_8433);
nand U14223 (N_14223,N_7912,N_7643);
and U14224 (N_14224,N_6855,N_9550);
nor U14225 (N_14225,N_7461,N_9856);
nand U14226 (N_14226,N_5674,N_7048);
or U14227 (N_14227,N_5177,N_8911);
xor U14228 (N_14228,N_7370,N_8917);
and U14229 (N_14229,N_6188,N_9670);
or U14230 (N_14230,N_7669,N_8270);
nand U14231 (N_14231,N_6013,N_9467);
nand U14232 (N_14232,N_5035,N_6944);
xnor U14233 (N_14233,N_5496,N_5546);
nand U14234 (N_14234,N_7603,N_6672);
nand U14235 (N_14235,N_9852,N_6605);
nand U14236 (N_14236,N_6743,N_5766);
xnor U14237 (N_14237,N_5847,N_5385);
or U14238 (N_14238,N_8636,N_5298);
or U14239 (N_14239,N_8464,N_5537);
nor U14240 (N_14240,N_8778,N_9567);
or U14241 (N_14241,N_5313,N_7611);
nor U14242 (N_14242,N_9884,N_7286);
and U14243 (N_14243,N_8760,N_5140);
nor U14244 (N_14244,N_5987,N_7398);
nor U14245 (N_14245,N_8184,N_8748);
nand U14246 (N_14246,N_7920,N_8822);
nor U14247 (N_14247,N_6003,N_7498);
or U14248 (N_14248,N_6743,N_5429);
or U14249 (N_14249,N_8805,N_7066);
nor U14250 (N_14250,N_7028,N_7011);
nor U14251 (N_14251,N_6387,N_9392);
nand U14252 (N_14252,N_6886,N_6892);
nand U14253 (N_14253,N_9893,N_8961);
xnor U14254 (N_14254,N_7541,N_6613);
and U14255 (N_14255,N_6230,N_7147);
nor U14256 (N_14256,N_6490,N_9270);
and U14257 (N_14257,N_9269,N_5866);
and U14258 (N_14258,N_5821,N_8404);
and U14259 (N_14259,N_7679,N_6858);
nor U14260 (N_14260,N_5262,N_6691);
or U14261 (N_14261,N_9838,N_6609);
or U14262 (N_14262,N_5856,N_9074);
nand U14263 (N_14263,N_5331,N_6134);
or U14264 (N_14264,N_7191,N_8712);
nor U14265 (N_14265,N_6203,N_7886);
or U14266 (N_14266,N_9342,N_7023);
nand U14267 (N_14267,N_8399,N_5599);
and U14268 (N_14268,N_5367,N_8401);
nor U14269 (N_14269,N_6272,N_9183);
and U14270 (N_14270,N_5883,N_9266);
nand U14271 (N_14271,N_5702,N_6172);
nand U14272 (N_14272,N_9635,N_8342);
nor U14273 (N_14273,N_7967,N_7221);
or U14274 (N_14274,N_5318,N_6005);
and U14275 (N_14275,N_8715,N_5225);
nor U14276 (N_14276,N_8715,N_9882);
nand U14277 (N_14277,N_8761,N_8717);
and U14278 (N_14278,N_6335,N_5847);
nor U14279 (N_14279,N_5816,N_8545);
nand U14280 (N_14280,N_9270,N_7757);
or U14281 (N_14281,N_5869,N_5921);
nor U14282 (N_14282,N_5497,N_7081);
nor U14283 (N_14283,N_8241,N_7193);
nand U14284 (N_14284,N_6662,N_7115);
or U14285 (N_14285,N_6263,N_7503);
nand U14286 (N_14286,N_5053,N_9532);
nor U14287 (N_14287,N_5107,N_5060);
or U14288 (N_14288,N_8041,N_6978);
xor U14289 (N_14289,N_9843,N_6528);
nor U14290 (N_14290,N_6674,N_7624);
nor U14291 (N_14291,N_8386,N_7374);
nor U14292 (N_14292,N_7267,N_9652);
and U14293 (N_14293,N_6983,N_6678);
nor U14294 (N_14294,N_6203,N_5274);
nor U14295 (N_14295,N_9512,N_6298);
nor U14296 (N_14296,N_8153,N_7056);
nor U14297 (N_14297,N_8108,N_8312);
and U14298 (N_14298,N_5255,N_9031);
or U14299 (N_14299,N_5658,N_5267);
and U14300 (N_14300,N_5274,N_8852);
nor U14301 (N_14301,N_5035,N_8256);
and U14302 (N_14302,N_8211,N_9344);
and U14303 (N_14303,N_8694,N_9592);
or U14304 (N_14304,N_7587,N_7986);
nor U14305 (N_14305,N_7987,N_5019);
or U14306 (N_14306,N_9855,N_9078);
nand U14307 (N_14307,N_5454,N_6059);
nand U14308 (N_14308,N_9425,N_9864);
and U14309 (N_14309,N_8737,N_9413);
nand U14310 (N_14310,N_6473,N_6708);
or U14311 (N_14311,N_6074,N_9798);
nand U14312 (N_14312,N_7325,N_8576);
nand U14313 (N_14313,N_9279,N_5476);
or U14314 (N_14314,N_7811,N_5569);
or U14315 (N_14315,N_6902,N_9829);
nand U14316 (N_14316,N_5777,N_7444);
nor U14317 (N_14317,N_5312,N_5912);
and U14318 (N_14318,N_8256,N_8156);
nor U14319 (N_14319,N_8356,N_9438);
nand U14320 (N_14320,N_5419,N_5374);
nand U14321 (N_14321,N_7844,N_9508);
and U14322 (N_14322,N_9236,N_9168);
or U14323 (N_14323,N_6619,N_5062);
nor U14324 (N_14324,N_6574,N_7224);
and U14325 (N_14325,N_6145,N_7464);
nor U14326 (N_14326,N_8773,N_7969);
or U14327 (N_14327,N_8127,N_8032);
and U14328 (N_14328,N_8861,N_5150);
or U14329 (N_14329,N_7038,N_7151);
nor U14330 (N_14330,N_8433,N_6502);
nand U14331 (N_14331,N_6200,N_9675);
nand U14332 (N_14332,N_6983,N_9204);
nor U14333 (N_14333,N_5547,N_8933);
nand U14334 (N_14334,N_8029,N_5862);
and U14335 (N_14335,N_7145,N_9778);
nor U14336 (N_14336,N_8568,N_9401);
and U14337 (N_14337,N_7387,N_9906);
or U14338 (N_14338,N_9287,N_8606);
or U14339 (N_14339,N_5605,N_6977);
nor U14340 (N_14340,N_8189,N_5114);
and U14341 (N_14341,N_7379,N_8804);
and U14342 (N_14342,N_5186,N_5110);
nor U14343 (N_14343,N_5213,N_7458);
nor U14344 (N_14344,N_9231,N_6136);
and U14345 (N_14345,N_7962,N_6916);
or U14346 (N_14346,N_6372,N_5967);
nand U14347 (N_14347,N_8738,N_6705);
nor U14348 (N_14348,N_7513,N_8318);
nor U14349 (N_14349,N_8250,N_6666);
nand U14350 (N_14350,N_6700,N_6286);
or U14351 (N_14351,N_5536,N_5227);
or U14352 (N_14352,N_5596,N_5634);
and U14353 (N_14353,N_9939,N_7361);
nor U14354 (N_14354,N_9908,N_9520);
nor U14355 (N_14355,N_7831,N_9246);
nor U14356 (N_14356,N_5094,N_6194);
and U14357 (N_14357,N_9536,N_8735);
or U14358 (N_14358,N_7222,N_9132);
or U14359 (N_14359,N_6499,N_7783);
or U14360 (N_14360,N_8302,N_5631);
and U14361 (N_14361,N_9663,N_6502);
and U14362 (N_14362,N_8424,N_8455);
and U14363 (N_14363,N_5289,N_7811);
nor U14364 (N_14364,N_9422,N_6342);
or U14365 (N_14365,N_6605,N_9047);
nand U14366 (N_14366,N_7831,N_6929);
nand U14367 (N_14367,N_7284,N_5238);
or U14368 (N_14368,N_8811,N_6764);
and U14369 (N_14369,N_9232,N_6027);
or U14370 (N_14370,N_6192,N_6155);
nor U14371 (N_14371,N_5877,N_8989);
nor U14372 (N_14372,N_8040,N_8626);
nor U14373 (N_14373,N_5099,N_5038);
or U14374 (N_14374,N_5008,N_8236);
or U14375 (N_14375,N_8683,N_9826);
nand U14376 (N_14376,N_5176,N_6592);
nor U14377 (N_14377,N_8880,N_7423);
and U14378 (N_14378,N_8844,N_8899);
nor U14379 (N_14379,N_7427,N_7662);
or U14380 (N_14380,N_8463,N_8607);
nor U14381 (N_14381,N_5265,N_9864);
nand U14382 (N_14382,N_7526,N_8928);
nand U14383 (N_14383,N_5298,N_9613);
xnor U14384 (N_14384,N_7836,N_6273);
or U14385 (N_14385,N_5214,N_6494);
nor U14386 (N_14386,N_8305,N_5709);
and U14387 (N_14387,N_9257,N_6798);
nand U14388 (N_14388,N_8676,N_9040);
and U14389 (N_14389,N_7300,N_9778);
and U14390 (N_14390,N_7082,N_5171);
and U14391 (N_14391,N_9956,N_6731);
or U14392 (N_14392,N_5354,N_7975);
nor U14393 (N_14393,N_7056,N_8274);
or U14394 (N_14394,N_5369,N_9548);
or U14395 (N_14395,N_7705,N_5281);
or U14396 (N_14396,N_7830,N_7993);
or U14397 (N_14397,N_7190,N_6262);
nand U14398 (N_14398,N_6331,N_5196);
or U14399 (N_14399,N_8499,N_5164);
and U14400 (N_14400,N_8155,N_9931);
nor U14401 (N_14401,N_8112,N_5689);
or U14402 (N_14402,N_5201,N_9486);
or U14403 (N_14403,N_9149,N_5925);
nand U14404 (N_14404,N_5962,N_8203);
nor U14405 (N_14405,N_6313,N_9733);
nor U14406 (N_14406,N_6090,N_9924);
nor U14407 (N_14407,N_6477,N_9102);
nor U14408 (N_14408,N_5807,N_5543);
nor U14409 (N_14409,N_6322,N_6736);
and U14410 (N_14410,N_6513,N_9166);
nor U14411 (N_14411,N_5507,N_9913);
and U14412 (N_14412,N_9815,N_8826);
and U14413 (N_14413,N_7009,N_6450);
and U14414 (N_14414,N_9523,N_7261);
xor U14415 (N_14415,N_7840,N_7189);
xnor U14416 (N_14416,N_5607,N_6671);
nand U14417 (N_14417,N_7687,N_7563);
nor U14418 (N_14418,N_7112,N_7830);
nor U14419 (N_14419,N_8879,N_5485);
nor U14420 (N_14420,N_8931,N_8862);
or U14421 (N_14421,N_8389,N_6227);
or U14422 (N_14422,N_8647,N_7068);
nand U14423 (N_14423,N_7075,N_9889);
or U14424 (N_14424,N_8482,N_6057);
nor U14425 (N_14425,N_5450,N_5400);
and U14426 (N_14426,N_5567,N_7947);
nor U14427 (N_14427,N_6295,N_9038);
nand U14428 (N_14428,N_6166,N_6768);
nor U14429 (N_14429,N_8460,N_8560);
nand U14430 (N_14430,N_7218,N_8268);
and U14431 (N_14431,N_5560,N_7673);
and U14432 (N_14432,N_6282,N_5512);
and U14433 (N_14433,N_7714,N_6978);
nor U14434 (N_14434,N_9310,N_7244);
nand U14435 (N_14435,N_8643,N_9184);
nand U14436 (N_14436,N_7590,N_9047);
nor U14437 (N_14437,N_7893,N_9402);
nor U14438 (N_14438,N_8884,N_7356);
nand U14439 (N_14439,N_6325,N_9742);
nand U14440 (N_14440,N_6842,N_5424);
xnor U14441 (N_14441,N_7292,N_7327);
nand U14442 (N_14442,N_8891,N_7588);
nor U14443 (N_14443,N_6627,N_6534);
or U14444 (N_14444,N_6368,N_7775);
or U14445 (N_14445,N_9876,N_5814);
or U14446 (N_14446,N_9070,N_7777);
or U14447 (N_14447,N_5055,N_9564);
nor U14448 (N_14448,N_7051,N_7127);
and U14449 (N_14449,N_6341,N_7231);
and U14450 (N_14450,N_8897,N_5003);
and U14451 (N_14451,N_5445,N_7248);
nor U14452 (N_14452,N_6074,N_7258);
nand U14453 (N_14453,N_5310,N_8402);
and U14454 (N_14454,N_9689,N_5568);
nor U14455 (N_14455,N_7550,N_7151);
and U14456 (N_14456,N_8683,N_8714);
nand U14457 (N_14457,N_9857,N_8971);
and U14458 (N_14458,N_9241,N_5196);
or U14459 (N_14459,N_6000,N_6543);
nor U14460 (N_14460,N_6899,N_7617);
or U14461 (N_14461,N_5581,N_5846);
nand U14462 (N_14462,N_9263,N_5737);
and U14463 (N_14463,N_7800,N_6354);
nand U14464 (N_14464,N_5850,N_7631);
nand U14465 (N_14465,N_9877,N_5698);
nor U14466 (N_14466,N_7772,N_5879);
nor U14467 (N_14467,N_6321,N_5578);
nand U14468 (N_14468,N_5102,N_8403);
nor U14469 (N_14469,N_6505,N_7576);
nand U14470 (N_14470,N_8822,N_7195);
and U14471 (N_14471,N_7826,N_5328);
or U14472 (N_14472,N_7321,N_7533);
nand U14473 (N_14473,N_9897,N_6641);
nor U14474 (N_14474,N_8234,N_5946);
or U14475 (N_14475,N_7125,N_7233);
xor U14476 (N_14476,N_7225,N_5356);
nand U14477 (N_14477,N_8785,N_8879);
nor U14478 (N_14478,N_5375,N_6322);
nor U14479 (N_14479,N_9082,N_8218);
or U14480 (N_14480,N_7876,N_5167);
and U14481 (N_14481,N_5595,N_8096);
nand U14482 (N_14482,N_9650,N_7654);
or U14483 (N_14483,N_5425,N_6433);
and U14484 (N_14484,N_6560,N_6811);
nor U14485 (N_14485,N_5455,N_9429);
or U14486 (N_14486,N_7255,N_5246);
and U14487 (N_14487,N_5429,N_9608);
nor U14488 (N_14488,N_7019,N_6669);
nand U14489 (N_14489,N_9398,N_6230);
nand U14490 (N_14490,N_6623,N_9162);
and U14491 (N_14491,N_9955,N_8753);
and U14492 (N_14492,N_8301,N_5574);
nor U14493 (N_14493,N_9338,N_7286);
nand U14494 (N_14494,N_5154,N_8104);
or U14495 (N_14495,N_6711,N_9478);
and U14496 (N_14496,N_5597,N_8810);
and U14497 (N_14497,N_9069,N_8899);
nor U14498 (N_14498,N_5493,N_5774);
and U14499 (N_14499,N_7295,N_6328);
or U14500 (N_14500,N_8172,N_6601);
or U14501 (N_14501,N_8572,N_6660);
nor U14502 (N_14502,N_5392,N_5039);
nand U14503 (N_14503,N_5586,N_6626);
and U14504 (N_14504,N_9987,N_8357);
nor U14505 (N_14505,N_7590,N_5978);
nor U14506 (N_14506,N_8046,N_7789);
nand U14507 (N_14507,N_9959,N_5710);
or U14508 (N_14508,N_5120,N_5344);
nand U14509 (N_14509,N_6158,N_7203);
or U14510 (N_14510,N_7159,N_6403);
and U14511 (N_14511,N_5001,N_5625);
nor U14512 (N_14512,N_5951,N_5236);
and U14513 (N_14513,N_6960,N_8108);
nor U14514 (N_14514,N_8286,N_7812);
nand U14515 (N_14515,N_9668,N_9344);
or U14516 (N_14516,N_8458,N_5848);
nor U14517 (N_14517,N_6717,N_5698);
nor U14518 (N_14518,N_9207,N_5855);
and U14519 (N_14519,N_6351,N_6209);
xor U14520 (N_14520,N_9571,N_7838);
nand U14521 (N_14521,N_8046,N_5447);
nand U14522 (N_14522,N_6170,N_5870);
nand U14523 (N_14523,N_5650,N_5938);
and U14524 (N_14524,N_7009,N_7850);
nand U14525 (N_14525,N_8030,N_9326);
and U14526 (N_14526,N_7178,N_5001);
nand U14527 (N_14527,N_5807,N_8660);
nor U14528 (N_14528,N_9811,N_5148);
and U14529 (N_14529,N_7971,N_5677);
nand U14530 (N_14530,N_5031,N_9832);
xnor U14531 (N_14531,N_8964,N_6663);
and U14532 (N_14532,N_9692,N_5087);
or U14533 (N_14533,N_7910,N_5131);
nor U14534 (N_14534,N_6312,N_8846);
and U14535 (N_14535,N_5272,N_7688);
or U14536 (N_14536,N_8264,N_9154);
or U14537 (N_14537,N_9998,N_9349);
nand U14538 (N_14538,N_6159,N_7645);
and U14539 (N_14539,N_8150,N_5344);
and U14540 (N_14540,N_5482,N_7253);
and U14541 (N_14541,N_5282,N_7083);
or U14542 (N_14542,N_8056,N_5591);
nand U14543 (N_14543,N_7293,N_9181);
nor U14544 (N_14544,N_6862,N_9935);
and U14545 (N_14545,N_9705,N_5834);
and U14546 (N_14546,N_5001,N_7877);
nand U14547 (N_14547,N_7255,N_9264);
and U14548 (N_14548,N_9167,N_8132);
nor U14549 (N_14549,N_6210,N_7298);
nand U14550 (N_14550,N_8174,N_5123);
or U14551 (N_14551,N_7212,N_7133);
or U14552 (N_14552,N_9648,N_8375);
nor U14553 (N_14553,N_7055,N_9713);
and U14554 (N_14554,N_9052,N_7660);
or U14555 (N_14555,N_6539,N_7415);
or U14556 (N_14556,N_7978,N_6723);
and U14557 (N_14557,N_7537,N_5608);
or U14558 (N_14558,N_5937,N_9896);
nand U14559 (N_14559,N_9655,N_6326);
nand U14560 (N_14560,N_7113,N_9210);
or U14561 (N_14561,N_8077,N_5858);
nor U14562 (N_14562,N_5284,N_7923);
nor U14563 (N_14563,N_7968,N_7436);
and U14564 (N_14564,N_9918,N_7631);
or U14565 (N_14565,N_7269,N_9945);
nor U14566 (N_14566,N_8636,N_5376);
nand U14567 (N_14567,N_9288,N_9160);
or U14568 (N_14568,N_8198,N_5998);
or U14569 (N_14569,N_9400,N_6226);
and U14570 (N_14570,N_7086,N_5912);
nor U14571 (N_14571,N_7839,N_6962);
nor U14572 (N_14572,N_5002,N_8116);
and U14573 (N_14573,N_5835,N_9138);
or U14574 (N_14574,N_6595,N_9711);
and U14575 (N_14575,N_9548,N_6064);
nand U14576 (N_14576,N_5559,N_5827);
nor U14577 (N_14577,N_6285,N_5719);
nor U14578 (N_14578,N_5828,N_8708);
and U14579 (N_14579,N_5744,N_6968);
and U14580 (N_14580,N_7731,N_6077);
or U14581 (N_14581,N_8897,N_7705);
or U14582 (N_14582,N_6640,N_6217);
nor U14583 (N_14583,N_9493,N_7984);
or U14584 (N_14584,N_6014,N_8790);
nand U14585 (N_14585,N_5000,N_6848);
and U14586 (N_14586,N_5573,N_5159);
or U14587 (N_14587,N_6750,N_9657);
and U14588 (N_14588,N_7006,N_9280);
xnor U14589 (N_14589,N_7596,N_8439);
nor U14590 (N_14590,N_5489,N_8518);
nand U14591 (N_14591,N_8261,N_6247);
nor U14592 (N_14592,N_6739,N_6731);
and U14593 (N_14593,N_5826,N_9601);
and U14594 (N_14594,N_9653,N_5791);
and U14595 (N_14595,N_6621,N_5323);
and U14596 (N_14596,N_5608,N_8024);
or U14597 (N_14597,N_6981,N_9159);
nand U14598 (N_14598,N_9429,N_9592);
nand U14599 (N_14599,N_6739,N_9683);
and U14600 (N_14600,N_8969,N_6786);
nand U14601 (N_14601,N_9292,N_9778);
nor U14602 (N_14602,N_6243,N_9397);
or U14603 (N_14603,N_8180,N_8282);
nor U14604 (N_14604,N_5635,N_6487);
or U14605 (N_14605,N_6467,N_5914);
nor U14606 (N_14606,N_9964,N_8439);
and U14607 (N_14607,N_9416,N_8458);
nand U14608 (N_14608,N_9624,N_5985);
and U14609 (N_14609,N_6113,N_9020);
or U14610 (N_14610,N_6701,N_7670);
nand U14611 (N_14611,N_8786,N_6211);
nand U14612 (N_14612,N_5364,N_6175);
nand U14613 (N_14613,N_8465,N_7724);
or U14614 (N_14614,N_6943,N_5977);
and U14615 (N_14615,N_6385,N_6080);
nand U14616 (N_14616,N_9090,N_6169);
nand U14617 (N_14617,N_5976,N_7966);
xnor U14618 (N_14618,N_6832,N_6847);
or U14619 (N_14619,N_9870,N_8286);
nand U14620 (N_14620,N_5446,N_8376);
or U14621 (N_14621,N_9501,N_9178);
or U14622 (N_14622,N_9822,N_6524);
nand U14623 (N_14623,N_6782,N_9994);
and U14624 (N_14624,N_8499,N_6499);
nand U14625 (N_14625,N_6840,N_6242);
nand U14626 (N_14626,N_6940,N_9077);
nor U14627 (N_14627,N_7772,N_8102);
nor U14628 (N_14628,N_8701,N_6581);
nor U14629 (N_14629,N_7478,N_8443);
or U14630 (N_14630,N_6106,N_6702);
or U14631 (N_14631,N_7801,N_5194);
or U14632 (N_14632,N_7890,N_5128);
or U14633 (N_14633,N_5799,N_6015);
and U14634 (N_14634,N_9452,N_8452);
nor U14635 (N_14635,N_6273,N_8122);
nand U14636 (N_14636,N_8173,N_6353);
nor U14637 (N_14637,N_8866,N_8332);
and U14638 (N_14638,N_5821,N_8429);
nor U14639 (N_14639,N_9133,N_8652);
nand U14640 (N_14640,N_5823,N_5118);
nor U14641 (N_14641,N_6933,N_5721);
nor U14642 (N_14642,N_7625,N_7451);
nor U14643 (N_14643,N_7767,N_9008);
nand U14644 (N_14644,N_5496,N_8044);
or U14645 (N_14645,N_8583,N_5663);
or U14646 (N_14646,N_7021,N_7531);
nor U14647 (N_14647,N_8262,N_6408);
and U14648 (N_14648,N_5749,N_9084);
nor U14649 (N_14649,N_6994,N_7319);
or U14650 (N_14650,N_8155,N_7750);
or U14651 (N_14651,N_7846,N_5245);
nor U14652 (N_14652,N_8554,N_6717);
or U14653 (N_14653,N_5466,N_9033);
xnor U14654 (N_14654,N_8994,N_9984);
nand U14655 (N_14655,N_9974,N_5639);
and U14656 (N_14656,N_9967,N_6637);
nand U14657 (N_14657,N_6320,N_5100);
and U14658 (N_14658,N_7167,N_5632);
or U14659 (N_14659,N_8775,N_8894);
nor U14660 (N_14660,N_5764,N_6237);
nand U14661 (N_14661,N_7334,N_7180);
and U14662 (N_14662,N_5196,N_6018);
nand U14663 (N_14663,N_8522,N_7249);
nor U14664 (N_14664,N_9571,N_8192);
nor U14665 (N_14665,N_9873,N_6949);
and U14666 (N_14666,N_9621,N_5434);
nor U14667 (N_14667,N_5981,N_5534);
or U14668 (N_14668,N_6743,N_9709);
nor U14669 (N_14669,N_6650,N_8809);
or U14670 (N_14670,N_7723,N_9544);
or U14671 (N_14671,N_6706,N_7323);
nor U14672 (N_14672,N_7487,N_5093);
nor U14673 (N_14673,N_8845,N_7636);
or U14674 (N_14674,N_8390,N_7946);
xnor U14675 (N_14675,N_5000,N_9737);
nand U14676 (N_14676,N_5969,N_7698);
nor U14677 (N_14677,N_8468,N_9174);
and U14678 (N_14678,N_5684,N_6900);
and U14679 (N_14679,N_8439,N_8637);
nand U14680 (N_14680,N_8154,N_6789);
nand U14681 (N_14681,N_8930,N_9568);
and U14682 (N_14682,N_5442,N_6005);
nand U14683 (N_14683,N_7691,N_7590);
nand U14684 (N_14684,N_7926,N_5445);
nor U14685 (N_14685,N_9060,N_7966);
nand U14686 (N_14686,N_6981,N_5275);
or U14687 (N_14687,N_5489,N_6657);
nor U14688 (N_14688,N_7673,N_7183);
nor U14689 (N_14689,N_6385,N_6652);
and U14690 (N_14690,N_8492,N_8787);
and U14691 (N_14691,N_7417,N_9212);
and U14692 (N_14692,N_9700,N_5784);
or U14693 (N_14693,N_8926,N_5924);
and U14694 (N_14694,N_5815,N_6427);
or U14695 (N_14695,N_9165,N_8118);
nor U14696 (N_14696,N_9462,N_9893);
or U14697 (N_14697,N_9729,N_8710);
and U14698 (N_14698,N_9845,N_6242);
or U14699 (N_14699,N_6937,N_5217);
nor U14700 (N_14700,N_9660,N_5768);
nand U14701 (N_14701,N_5374,N_9326);
and U14702 (N_14702,N_8914,N_6433);
and U14703 (N_14703,N_9486,N_6511);
nor U14704 (N_14704,N_8284,N_9291);
nand U14705 (N_14705,N_6510,N_9935);
or U14706 (N_14706,N_8757,N_8693);
or U14707 (N_14707,N_7474,N_6947);
or U14708 (N_14708,N_6676,N_9494);
and U14709 (N_14709,N_6852,N_6408);
xor U14710 (N_14710,N_8602,N_8732);
or U14711 (N_14711,N_5255,N_7370);
nand U14712 (N_14712,N_5764,N_6321);
nand U14713 (N_14713,N_9616,N_8512);
nor U14714 (N_14714,N_9265,N_5138);
and U14715 (N_14715,N_9673,N_9584);
and U14716 (N_14716,N_8214,N_7552);
and U14717 (N_14717,N_9937,N_5845);
or U14718 (N_14718,N_8550,N_5384);
or U14719 (N_14719,N_7310,N_6360);
and U14720 (N_14720,N_6240,N_9630);
nand U14721 (N_14721,N_5198,N_6690);
or U14722 (N_14722,N_6762,N_5109);
nor U14723 (N_14723,N_8716,N_9852);
xnor U14724 (N_14724,N_5531,N_5910);
nand U14725 (N_14725,N_9234,N_6964);
or U14726 (N_14726,N_9619,N_5266);
nor U14727 (N_14727,N_8544,N_8412);
or U14728 (N_14728,N_6976,N_6337);
and U14729 (N_14729,N_7638,N_9985);
or U14730 (N_14730,N_6202,N_7169);
or U14731 (N_14731,N_8952,N_6839);
nor U14732 (N_14732,N_9298,N_6686);
nand U14733 (N_14733,N_5582,N_9014);
nor U14734 (N_14734,N_6521,N_5909);
or U14735 (N_14735,N_5753,N_7001);
or U14736 (N_14736,N_5245,N_9520);
or U14737 (N_14737,N_9247,N_9962);
nand U14738 (N_14738,N_8721,N_9039);
or U14739 (N_14739,N_7380,N_9817);
and U14740 (N_14740,N_5637,N_5060);
nor U14741 (N_14741,N_9213,N_6249);
or U14742 (N_14742,N_8093,N_7243);
nand U14743 (N_14743,N_8157,N_7591);
or U14744 (N_14744,N_7947,N_6288);
and U14745 (N_14745,N_8948,N_9882);
or U14746 (N_14746,N_6287,N_8000);
nand U14747 (N_14747,N_7165,N_6346);
nor U14748 (N_14748,N_7285,N_6702);
nor U14749 (N_14749,N_7011,N_6204);
or U14750 (N_14750,N_7245,N_7122);
and U14751 (N_14751,N_5042,N_8728);
nand U14752 (N_14752,N_7852,N_7101);
or U14753 (N_14753,N_8075,N_7973);
nor U14754 (N_14754,N_9181,N_8550);
and U14755 (N_14755,N_5804,N_9708);
and U14756 (N_14756,N_6434,N_8805);
nor U14757 (N_14757,N_6656,N_8032);
and U14758 (N_14758,N_6796,N_8558);
or U14759 (N_14759,N_8677,N_5991);
and U14760 (N_14760,N_9323,N_7451);
and U14761 (N_14761,N_9365,N_5592);
nor U14762 (N_14762,N_8745,N_8095);
and U14763 (N_14763,N_8461,N_9947);
and U14764 (N_14764,N_8154,N_9528);
xor U14765 (N_14765,N_7781,N_9542);
and U14766 (N_14766,N_8334,N_7067);
nor U14767 (N_14767,N_9437,N_7956);
and U14768 (N_14768,N_9206,N_6188);
and U14769 (N_14769,N_9933,N_9069);
or U14770 (N_14770,N_5153,N_8177);
nand U14771 (N_14771,N_7043,N_7080);
or U14772 (N_14772,N_9908,N_7879);
and U14773 (N_14773,N_9612,N_5904);
or U14774 (N_14774,N_8653,N_6502);
and U14775 (N_14775,N_8782,N_8527);
or U14776 (N_14776,N_7497,N_6771);
nand U14777 (N_14777,N_7572,N_7792);
xnor U14778 (N_14778,N_6842,N_9132);
nor U14779 (N_14779,N_9622,N_8163);
and U14780 (N_14780,N_8631,N_7609);
nand U14781 (N_14781,N_8874,N_7446);
nand U14782 (N_14782,N_7702,N_6089);
nor U14783 (N_14783,N_7484,N_8483);
nor U14784 (N_14784,N_7853,N_5616);
nand U14785 (N_14785,N_8190,N_6391);
nand U14786 (N_14786,N_6477,N_7946);
or U14787 (N_14787,N_6462,N_7563);
nand U14788 (N_14788,N_6865,N_5454);
and U14789 (N_14789,N_6128,N_7396);
and U14790 (N_14790,N_5637,N_8069);
nand U14791 (N_14791,N_5834,N_7520);
nand U14792 (N_14792,N_6999,N_9978);
nand U14793 (N_14793,N_8641,N_7373);
xnor U14794 (N_14794,N_7314,N_8749);
nor U14795 (N_14795,N_8461,N_7588);
xnor U14796 (N_14796,N_6501,N_8538);
xor U14797 (N_14797,N_8044,N_8637);
or U14798 (N_14798,N_8105,N_8372);
nor U14799 (N_14799,N_5444,N_6193);
xor U14800 (N_14800,N_5609,N_9345);
nand U14801 (N_14801,N_8628,N_6259);
xor U14802 (N_14802,N_7439,N_5827);
nand U14803 (N_14803,N_6797,N_7508);
nand U14804 (N_14804,N_7157,N_6232);
nor U14805 (N_14805,N_8201,N_7480);
nand U14806 (N_14806,N_5125,N_6060);
nand U14807 (N_14807,N_5508,N_5624);
nor U14808 (N_14808,N_7448,N_7166);
nand U14809 (N_14809,N_7402,N_6615);
or U14810 (N_14810,N_8457,N_6120);
nand U14811 (N_14811,N_9746,N_8508);
nor U14812 (N_14812,N_5221,N_8595);
and U14813 (N_14813,N_9888,N_8997);
nor U14814 (N_14814,N_8079,N_8185);
nand U14815 (N_14815,N_7280,N_5430);
or U14816 (N_14816,N_9131,N_6339);
nor U14817 (N_14817,N_8812,N_5040);
and U14818 (N_14818,N_6747,N_5815);
nor U14819 (N_14819,N_8237,N_9790);
nand U14820 (N_14820,N_9486,N_9565);
and U14821 (N_14821,N_6255,N_7407);
or U14822 (N_14822,N_5695,N_8233);
or U14823 (N_14823,N_7886,N_8310);
and U14824 (N_14824,N_9729,N_7872);
nand U14825 (N_14825,N_6661,N_7349);
nand U14826 (N_14826,N_5521,N_9868);
nor U14827 (N_14827,N_9805,N_6050);
xnor U14828 (N_14828,N_5054,N_8214);
or U14829 (N_14829,N_8120,N_8546);
nor U14830 (N_14830,N_8186,N_8454);
nand U14831 (N_14831,N_5861,N_8779);
and U14832 (N_14832,N_5370,N_8368);
nand U14833 (N_14833,N_9084,N_6609);
or U14834 (N_14834,N_6657,N_7874);
or U14835 (N_14835,N_8043,N_6764);
and U14836 (N_14836,N_8858,N_8800);
nor U14837 (N_14837,N_6392,N_5872);
and U14838 (N_14838,N_5345,N_6943);
nand U14839 (N_14839,N_9524,N_9710);
or U14840 (N_14840,N_8691,N_6284);
nand U14841 (N_14841,N_8685,N_7058);
nand U14842 (N_14842,N_5957,N_5305);
nand U14843 (N_14843,N_5448,N_9344);
nand U14844 (N_14844,N_9197,N_5434);
or U14845 (N_14845,N_6647,N_9237);
nor U14846 (N_14846,N_5898,N_5120);
nand U14847 (N_14847,N_9107,N_7184);
xor U14848 (N_14848,N_9296,N_6328);
xor U14849 (N_14849,N_6322,N_5435);
nand U14850 (N_14850,N_7863,N_8879);
xnor U14851 (N_14851,N_5466,N_7981);
nand U14852 (N_14852,N_6152,N_8275);
and U14853 (N_14853,N_8256,N_7681);
nand U14854 (N_14854,N_5661,N_8400);
and U14855 (N_14855,N_9549,N_9155);
or U14856 (N_14856,N_7499,N_5739);
or U14857 (N_14857,N_6397,N_8642);
or U14858 (N_14858,N_7395,N_7062);
nor U14859 (N_14859,N_7578,N_6992);
and U14860 (N_14860,N_5067,N_8666);
or U14861 (N_14861,N_9065,N_5484);
nor U14862 (N_14862,N_9059,N_7103);
nor U14863 (N_14863,N_7866,N_8862);
or U14864 (N_14864,N_5575,N_6501);
nor U14865 (N_14865,N_5403,N_9175);
nor U14866 (N_14866,N_6424,N_5568);
and U14867 (N_14867,N_9669,N_7607);
or U14868 (N_14868,N_5243,N_6978);
nor U14869 (N_14869,N_7623,N_5779);
nor U14870 (N_14870,N_9399,N_9936);
nand U14871 (N_14871,N_8461,N_5936);
nand U14872 (N_14872,N_5975,N_5398);
or U14873 (N_14873,N_7086,N_7619);
or U14874 (N_14874,N_5366,N_6918);
nor U14875 (N_14875,N_5981,N_8836);
nand U14876 (N_14876,N_6248,N_5785);
nand U14877 (N_14877,N_7018,N_9615);
nor U14878 (N_14878,N_7776,N_7958);
xor U14879 (N_14879,N_5870,N_9914);
nor U14880 (N_14880,N_7495,N_8991);
and U14881 (N_14881,N_7644,N_5725);
and U14882 (N_14882,N_6677,N_8447);
and U14883 (N_14883,N_6668,N_9835);
nor U14884 (N_14884,N_9706,N_6168);
nor U14885 (N_14885,N_7009,N_8492);
xor U14886 (N_14886,N_9215,N_5870);
and U14887 (N_14887,N_5806,N_7432);
nand U14888 (N_14888,N_9283,N_8905);
nor U14889 (N_14889,N_9559,N_7594);
nor U14890 (N_14890,N_9590,N_6636);
nor U14891 (N_14891,N_8900,N_9860);
nor U14892 (N_14892,N_6367,N_7793);
and U14893 (N_14893,N_9732,N_5934);
or U14894 (N_14894,N_6732,N_7563);
nor U14895 (N_14895,N_5212,N_5274);
and U14896 (N_14896,N_6905,N_5914);
nand U14897 (N_14897,N_6994,N_6901);
and U14898 (N_14898,N_8947,N_5286);
nor U14899 (N_14899,N_9174,N_8610);
nand U14900 (N_14900,N_5198,N_9438);
nor U14901 (N_14901,N_9350,N_7733);
nor U14902 (N_14902,N_7906,N_9200);
nor U14903 (N_14903,N_9694,N_6283);
and U14904 (N_14904,N_8676,N_8953);
nand U14905 (N_14905,N_6543,N_9124);
xor U14906 (N_14906,N_8155,N_7994);
nand U14907 (N_14907,N_6450,N_7958);
or U14908 (N_14908,N_7675,N_5356);
or U14909 (N_14909,N_5015,N_6372);
or U14910 (N_14910,N_5386,N_8493);
or U14911 (N_14911,N_9048,N_8491);
nand U14912 (N_14912,N_5092,N_6721);
nor U14913 (N_14913,N_9961,N_8367);
and U14914 (N_14914,N_5638,N_9724);
nor U14915 (N_14915,N_9065,N_8032);
and U14916 (N_14916,N_6602,N_9499);
nor U14917 (N_14917,N_5531,N_6823);
and U14918 (N_14918,N_9395,N_8304);
and U14919 (N_14919,N_9528,N_6183);
nand U14920 (N_14920,N_6496,N_9741);
nand U14921 (N_14921,N_5265,N_5316);
nor U14922 (N_14922,N_7640,N_8470);
and U14923 (N_14923,N_8889,N_8784);
xnor U14924 (N_14924,N_6750,N_7306);
or U14925 (N_14925,N_9077,N_6357);
nor U14926 (N_14926,N_6831,N_8478);
nand U14927 (N_14927,N_9860,N_6398);
nand U14928 (N_14928,N_9412,N_8818);
nand U14929 (N_14929,N_7342,N_6961);
or U14930 (N_14930,N_8266,N_5714);
and U14931 (N_14931,N_6239,N_8160);
nand U14932 (N_14932,N_5972,N_7407);
or U14933 (N_14933,N_9781,N_9837);
and U14934 (N_14934,N_6683,N_6456);
nand U14935 (N_14935,N_8845,N_9482);
and U14936 (N_14936,N_7304,N_9380);
and U14937 (N_14937,N_5856,N_6240);
or U14938 (N_14938,N_7627,N_5473);
nand U14939 (N_14939,N_9360,N_7756);
and U14940 (N_14940,N_8070,N_6994);
nand U14941 (N_14941,N_5244,N_9036);
nor U14942 (N_14942,N_5876,N_8067);
or U14943 (N_14943,N_5879,N_8009);
and U14944 (N_14944,N_7016,N_5949);
nor U14945 (N_14945,N_6524,N_9721);
and U14946 (N_14946,N_8155,N_6687);
and U14947 (N_14947,N_9359,N_7696);
and U14948 (N_14948,N_9672,N_6754);
nor U14949 (N_14949,N_7335,N_7677);
nand U14950 (N_14950,N_5177,N_6872);
or U14951 (N_14951,N_8102,N_8506);
nor U14952 (N_14952,N_7949,N_8505);
nand U14953 (N_14953,N_9047,N_6731);
xor U14954 (N_14954,N_6566,N_9922);
nand U14955 (N_14955,N_7514,N_9635);
nand U14956 (N_14956,N_5146,N_5575);
nor U14957 (N_14957,N_9427,N_9627);
nor U14958 (N_14958,N_6588,N_8946);
xnor U14959 (N_14959,N_8660,N_8565);
and U14960 (N_14960,N_5961,N_7178);
nor U14961 (N_14961,N_9506,N_9932);
nor U14962 (N_14962,N_9335,N_5870);
nand U14963 (N_14963,N_9824,N_7942);
or U14964 (N_14964,N_5605,N_8412);
and U14965 (N_14965,N_7297,N_6817);
nand U14966 (N_14966,N_9679,N_9445);
nand U14967 (N_14967,N_8259,N_7775);
or U14968 (N_14968,N_5406,N_6907);
or U14969 (N_14969,N_7258,N_8736);
nor U14970 (N_14970,N_5639,N_5434);
and U14971 (N_14971,N_7932,N_9240);
nand U14972 (N_14972,N_7584,N_7965);
nand U14973 (N_14973,N_8296,N_5494);
nand U14974 (N_14974,N_7740,N_5865);
or U14975 (N_14975,N_7966,N_8721);
nand U14976 (N_14976,N_5219,N_8193);
or U14977 (N_14977,N_7083,N_8694);
and U14978 (N_14978,N_7619,N_7582);
nor U14979 (N_14979,N_6060,N_6658);
or U14980 (N_14980,N_7242,N_7910);
nor U14981 (N_14981,N_9798,N_7263);
and U14982 (N_14982,N_8410,N_8423);
or U14983 (N_14983,N_8837,N_6569);
nor U14984 (N_14984,N_9315,N_5133);
nand U14985 (N_14985,N_5239,N_7539);
nand U14986 (N_14986,N_5229,N_7538);
nor U14987 (N_14987,N_9469,N_5375);
and U14988 (N_14988,N_9420,N_8934);
and U14989 (N_14989,N_5425,N_6443);
and U14990 (N_14990,N_9474,N_9197);
and U14991 (N_14991,N_6139,N_5627);
or U14992 (N_14992,N_8008,N_9385);
or U14993 (N_14993,N_8796,N_6441);
or U14994 (N_14994,N_7287,N_6919);
nand U14995 (N_14995,N_9419,N_6576);
nand U14996 (N_14996,N_5984,N_7521);
nor U14997 (N_14997,N_7444,N_9303);
and U14998 (N_14998,N_9556,N_5266);
nor U14999 (N_14999,N_9392,N_7955);
nand UO_0 (O_0,N_12585,N_11124);
and UO_1 (O_1,N_13955,N_11338);
nand UO_2 (O_2,N_12000,N_13388);
nand UO_3 (O_3,N_14622,N_12477);
nand UO_4 (O_4,N_11034,N_12047);
or UO_5 (O_5,N_11846,N_11234);
and UO_6 (O_6,N_11159,N_11170);
nor UO_7 (O_7,N_12395,N_11558);
and UO_8 (O_8,N_10164,N_11378);
and UO_9 (O_9,N_10741,N_13016);
nor UO_10 (O_10,N_13007,N_11887);
or UO_11 (O_11,N_11021,N_13817);
or UO_12 (O_12,N_13069,N_11551);
or UO_13 (O_13,N_11516,N_14303);
or UO_14 (O_14,N_10757,N_14386);
nor UO_15 (O_15,N_11067,N_10719);
nand UO_16 (O_16,N_13249,N_10252);
or UO_17 (O_17,N_11235,N_14959);
or UO_18 (O_18,N_10834,N_11517);
nor UO_19 (O_19,N_14063,N_13229);
or UO_20 (O_20,N_14084,N_14343);
and UO_21 (O_21,N_13285,N_14742);
nor UO_22 (O_22,N_10400,N_10798);
nor UO_23 (O_23,N_14675,N_13088);
and UO_24 (O_24,N_12162,N_12236);
or UO_25 (O_25,N_13198,N_14526);
nor UO_26 (O_26,N_12911,N_13361);
or UO_27 (O_27,N_12074,N_12837);
or UO_28 (O_28,N_11582,N_10549);
and UO_29 (O_29,N_11876,N_13337);
and UO_30 (O_30,N_10978,N_13423);
nor UO_31 (O_31,N_11443,N_10825);
and UO_32 (O_32,N_11926,N_14522);
nand UO_33 (O_33,N_12091,N_10368);
nor UO_34 (O_34,N_12145,N_13497);
nor UO_35 (O_35,N_14064,N_12918);
nor UO_36 (O_36,N_12922,N_14460);
nor UO_37 (O_37,N_10673,N_14909);
and UO_38 (O_38,N_12247,N_12470);
and UO_39 (O_39,N_10904,N_10930);
nand UO_40 (O_40,N_10344,N_11025);
nor UO_41 (O_41,N_11527,N_12723);
nor UO_42 (O_42,N_12989,N_13605);
or UO_43 (O_43,N_13734,N_12063);
nor UO_44 (O_44,N_11473,N_10081);
nor UO_45 (O_45,N_13597,N_11142);
nor UO_46 (O_46,N_13414,N_11705);
or UO_47 (O_47,N_12773,N_11716);
and UO_48 (O_48,N_12133,N_10919);
and UO_49 (O_49,N_14430,N_10781);
and UO_50 (O_50,N_12886,N_13091);
and UO_51 (O_51,N_13496,N_10106);
or UO_52 (O_52,N_14586,N_14336);
and UO_53 (O_53,N_12718,N_12439);
or UO_54 (O_54,N_14022,N_14344);
nand UO_55 (O_55,N_12956,N_10233);
and UO_56 (O_56,N_12045,N_12154);
or UO_57 (O_57,N_11864,N_11560);
nand UO_58 (O_58,N_12218,N_12969);
or UO_59 (O_59,N_13818,N_12607);
and UO_60 (O_60,N_13868,N_12110);
or UO_61 (O_61,N_12589,N_10989);
nor UO_62 (O_62,N_11015,N_12117);
or UO_63 (O_63,N_10500,N_14059);
nor UO_64 (O_64,N_12840,N_10955);
or UO_65 (O_65,N_14703,N_14677);
nor UO_66 (O_66,N_11192,N_11083);
or UO_67 (O_67,N_11950,N_14974);
nor UO_68 (O_68,N_11165,N_10687);
nor UO_69 (O_69,N_12704,N_14918);
or UO_70 (O_70,N_10382,N_11737);
and UO_71 (O_71,N_13537,N_11735);
or UO_72 (O_72,N_10421,N_11964);
nand UO_73 (O_73,N_10685,N_10112);
nand UO_74 (O_74,N_13363,N_10574);
nor UO_75 (O_75,N_10702,N_11143);
or UO_76 (O_76,N_13051,N_11260);
nand UO_77 (O_77,N_14815,N_12243);
or UO_78 (O_78,N_10912,N_10176);
nor UO_79 (O_79,N_10950,N_11005);
and UO_80 (O_80,N_10525,N_10486);
or UO_81 (O_81,N_11168,N_13312);
and UO_82 (O_82,N_12590,N_12284);
and UO_83 (O_83,N_14783,N_14953);
nor UO_84 (O_84,N_11559,N_13023);
and UO_85 (O_85,N_13653,N_10315);
and UO_86 (O_86,N_11528,N_13167);
and UO_87 (O_87,N_11684,N_12643);
or UO_88 (O_88,N_10841,N_13146);
nor UO_89 (O_89,N_12090,N_11413);
nand UO_90 (O_90,N_11689,N_14427);
nor UO_91 (O_91,N_11725,N_12797);
or UO_92 (O_92,N_13438,N_12616);
and UO_93 (O_93,N_13319,N_13060);
nand UO_94 (O_94,N_10823,N_14501);
nand UO_95 (O_95,N_14672,N_10737);
and UO_96 (O_96,N_11388,N_13222);
nor UO_97 (O_97,N_12546,N_11662);
and UO_98 (O_98,N_11721,N_13972);
or UO_99 (O_99,N_11878,N_14168);
nand UO_100 (O_100,N_13988,N_12936);
nor UO_101 (O_101,N_11982,N_12142);
and UO_102 (O_102,N_12564,N_14905);
and UO_103 (O_103,N_12229,N_14973);
and UO_104 (O_104,N_11714,N_13459);
nand UO_105 (O_105,N_13122,N_11387);
nand UO_106 (O_106,N_10513,N_12424);
and UO_107 (O_107,N_14512,N_13776);
nor UO_108 (O_108,N_10839,N_12124);
nand UO_109 (O_109,N_12135,N_13384);
nand UO_110 (O_110,N_12964,N_11902);
nand UO_111 (O_111,N_12664,N_10494);
or UO_112 (O_112,N_11284,N_13846);
or UO_113 (O_113,N_11773,N_12605);
and UO_114 (O_114,N_10546,N_11127);
xnor UO_115 (O_115,N_10680,N_10416);
nand UO_116 (O_116,N_10872,N_11693);
or UO_117 (O_117,N_10042,N_13819);
nand UO_118 (O_118,N_11750,N_10111);
or UO_119 (O_119,N_13159,N_14514);
nand UO_120 (O_120,N_13834,N_12908);
and UO_121 (O_121,N_13591,N_14319);
or UO_122 (O_122,N_13108,N_12088);
or UO_123 (O_123,N_11374,N_10257);
or UO_124 (O_124,N_13386,N_13073);
nor UO_125 (O_125,N_13473,N_13435);
or UO_126 (O_126,N_12128,N_14813);
or UO_127 (O_127,N_13969,N_14618);
or UO_128 (O_128,N_12534,N_11213);
nand UO_129 (O_129,N_10827,N_12623);
nand UO_130 (O_130,N_11086,N_10538);
or UO_131 (O_131,N_13329,N_12639);
or UO_132 (O_132,N_13499,N_11101);
nor UO_133 (O_133,N_10490,N_10566);
and UO_134 (O_134,N_14454,N_13451);
nor UO_135 (O_135,N_12671,N_11660);
and UO_136 (O_136,N_14060,N_14692);
and UO_137 (O_137,N_11727,N_12998);
nor UO_138 (O_138,N_10796,N_12249);
and UO_139 (O_139,N_12370,N_12848);
nand UO_140 (O_140,N_13560,N_13567);
xnor UO_141 (O_141,N_11783,N_12137);
xnor UO_142 (O_142,N_14264,N_14024);
or UO_143 (O_143,N_12121,N_13749);
nand UO_144 (O_144,N_10529,N_13411);
nand UO_145 (O_145,N_12985,N_13291);
nor UO_146 (O_146,N_13658,N_10711);
nor UO_147 (O_147,N_11497,N_10761);
nor UO_148 (O_148,N_11202,N_11011);
or UO_149 (O_149,N_12944,N_13804);
nand UO_150 (O_150,N_10283,N_12600);
and UO_151 (O_151,N_14612,N_11477);
nand UO_152 (O_152,N_10888,N_14708);
or UO_153 (O_153,N_12553,N_12581);
nand UO_154 (O_154,N_10752,N_12914);
and UO_155 (O_155,N_10663,N_12877);
or UO_156 (O_156,N_10578,N_10943);
nand UO_157 (O_157,N_10646,N_12673);
and UO_158 (O_158,N_11007,N_13533);
nor UO_159 (O_159,N_13068,N_11571);
nand UO_160 (O_160,N_10868,N_14626);
or UO_161 (O_161,N_10173,N_14422);
nor UO_162 (O_162,N_12920,N_10146);
or UO_163 (O_163,N_12267,N_13121);
nand UO_164 (O_164,N_10745,N_14090);
nor UO_165 (O_165,N_10581,N_11405);
or UO_166 (O_166,N_11091,N_10805);
nor UO_167 (O_167,N_10947,N_13678);
and UO_168 (O_168,N_12160,N_14348);
nor UO_169 (O_169,N_10028,N_11930);
nand UO_170 (O_170,N_10776,N_13688);
nand UO_171 (O_171,N_10148,N_14238);
nor UO_172 (O_172,N_10532,N_14653);
nor UO_173 (O_173,N_12663,N_10429);
nand UO_174 (O_174,N_10598,N_12491);
and UO_175 (O_175,N_10223,N_14435);
nand UO_176 (O_176,N_13092,N_14868);
and UO_177 (O_177,N_11460,N_12732);
or UO_178 (O_178,N_13349,N_10411);
or UO_179 (O_179,N_14505,N_12120);
or UO_180 (O_180,N_10863,N_10672);
nand UO_181 (O_181,N_13015,N_11045);
or UO_182 (O_182,N_13794,N_11332);
nand UO_183 (O_183,N_11096,N_11752);
nor UO_184 (O_184,N_10976,N_11164);
nand UO_185 (O_185,N_11184,N_12881);
and UO_186 (O_186,N_12510,N_13885);
and UO_187 (O_187,N_14880,N_13244);
nand UO_188 (O_188,N_10445,N_12321);
nor UO_189 (O_189,N_12651,N_13266);
nor UO_190 (O_190,N_11268,N_11478);
and UO_191 (O_191,N_13067,N_13735);
or UO_192 (O_192,N_13293,N_14242);
or UO_193 (O_193,N_11825,N_10481);
nand UO_194 (O_194,N_13071,N_13436);
and UO_195 (O_195,N_12994,N_10789);
and UO_196 (O_196,N_13135,N_13783);
nor UO_197 (O_197,N_11506,N_12924);
nor UO_198 (O_198,N_10640,N_11932);
nor UO_199 (O_199,N_13324,N_13295);
and UO_200 (O_200,N_12237,N_12131);
nor UO_201 (O_201,N_12661,N_10985);
nor UO_202 (O_202,N_10509,N_11061);
and UO_203 (O_203,N_14822,N_10265);
or UO_204 (O_204,N_11563,N_12845);
or UO_205 (O_205,N_14236,N_12305);
nand UO_206 (O_206,N_11562,N_13635);
and UO_207 (O_207,N_11016,N_12084);
and UO_208 (O_208,N_10448,N_14785);
nand UO_209 (O_209,N_13033,N_13975);
nor UO_210 (O_210,N_10077,N_10883);
and UO_211 (O_211,N_13536,N_13509);
or UO_212 (O_212,N_14132,N_13990);
nor UO_213 (O_213,N_10683,N_11505);
and UO_214 (O_214,N_14010,N_12948);
nor UO_215 (O_215,N_14334,N_13055);
nand UO_216 (O_216,N_10234,N_10703);
and UO_217 (O_217,N_12642,N_13265);
nand UO_218 (O_218,N_10221,N_14478);
nor UO_219 (O_219,N_14362,N_14206);
and UO_220 (O_220,N_12155,N_12447);
or UO_221 (O_221,N_11272,N_13401);
nand UO_222 (O_222,N_12980,N_12547);
nand UO_223 (O_223,N_13609,N_13276);
nor UO_224 (O_224,N_12233,N_14706);
nand UO_225 (O_225,N_14342,N_11906);
and UO_226 (O_226,N_13449,N_11112);
nand UO_227 (O_227,N_13883,N_12052);
nor UO_228 (O_228,N_12729,N_14472);
nor UO_229 (O_229,N_10551,N_13627);
nor UO_230 (O_230,N_13516,N_12649);
nand UO_231 (O_231,N_14922,N_10918);
or UO_232 (O_232,N_11905,N_12039);
nand UO_233 (O_233,N_13484,N_13177);
nor UO_234 (O_234,N_12612,N_11126);
nand UO_235 (O_235,N_14580,N_13194);
nor UO_236 (O_236,N_11316,N_13645);
or UO_237 (O_237,N_14183,N_11307);
nand UO_238 (O_238,N_10542,N_11400);
or UO_239 (O_239,N_10437,N_10634);
nor UO_240 (O_240,N_10025,N_12053);
and UO_241 (O_241,N_10960,N_13781);
or UO_242 (O_242,N_10853,N_10880);
and UO_243 (O_243,N_14149,N_11257);
xnor UO_244 (O_244,N_14109,N_11232);
nor UO_245 (O_245,N_11064,N_10425);
and UO_246 (O_246,N_13080,N_14452);
nand UO_247 (O_247,N_13682,N_14419);
nor UO_248 (O_248,N_11057,N_11765);
nor UO_249 (O_249,N_12101,N_12753);
nand UO_250 (O_250,N_11448,N_10763);
or UO_251 (O_251,N_12380,N_14124);
nor UO_252 (O_252,N_11815,N_14667);
and UO_253 (O_253,N_14438,N_11771);
nand UO_254 (O_254,N_13157,N_14794);
nor UO_255 (O_255,N_13942,N_10260);
nor UO_256 (O_256,N_12250,N_14338);
or UO_257 (O_257,N_10651,N_14963);
or UO_258 (O_258,N_14004,N_11366);
or UO_259 (O_259,N_14701,N_11324);
xor UO_260 (O_260,N_13862,N_13274);
and UO_261 (O_261,N_12792,N_10463);
or UO_262 (O_262,N_10365,N_13570);
xor UO_263 (O_263,N_10984,N_10621);
or UO_264 (O_264,N_12786,N_11784);
nand UO_265 (O_265,N_12670,N_13544);
nor UO_266 (O_266,N_10231,N_12388);
or UO_267 (O_267,N_14572,N_12206);
xnor UO_268 (O_268,N_14499,N_13982);
nor UO_269 (O_269,N_10877,N_10996);
or UO_270 (O_270,N_12310,N_13822);
nor UO_271 (O_271,N_13145,N_14251);
nor UO_272 (O_272,N_10705,N_10386);
nor UO_273 (O_273,N_10632,N_14987);
and UO_274 (O_274,N_12488,N_10945);
nor UO_275 (O_275,N_14574,N_11245);
nand UO_276 (O_276,N_14786,N_13926);
or UO_277 (O_277,N_10762,N_13503);
and UO_278 (O_278,N_10108,N_14417);
and UO_279 (O_279,N_13815,N_14535);
and UO_280 (O_280,N_12733,N_10491);
and UO_281 (O_281,N_12355,N_10890);
or UO_282 (O_282,N_14763,N_11146);
and UO_283 (O_283,N_13890,N_11301);
nor UO_284 (O_284,N_12941,N_10414);
nand UO_285 (O_285,N_13501,N_12288);
nor UO_286 (O_286,N_10684,N_11909);
nand UO_287 (O_287,N_14494,N_10541);
and UO_288 (O_288,N_10301,N_11363);
and UO_289 (O_289,N_14518,N_13486);
or UO_290 (O_290,N_14223,N_13928);
nor UO_291 (O_291,N_12629,N_11487);
nand UO_292 (O_292,N_10389,N_10946);
and UO_293 (O_293,N_12529,N_10855);
or UO_294 (O_294,N_10436,N_11147);
and UO_295 (O_295,N_10917,N_12660);
and UO_296 (O_296,N_13392,N_10939);
and UO_297 (O_297,N_12608,N_14732);
nor UO_298 (O_298,N_11241,N_12909);
and UO_299 (O_299,N_12526,N_13922);
nor UO_300 (O_300,N_11479,N_11075);
nand UO_301 (O_301,N_12406,N_11258);
nor UO_302 (O_302,N_13076,N_13661);
nor UO_303 (O_303,N_11854,N_13947);
or UO_304 (O_304,N_13753,N_13095);
nor UO_305 (O_305,N_14311,N_11029);
and UO_306 (O_306,N_12967,N_13318);
nand UO_307 (O_307,N_12330,N_11039);
and UO_308 (O_308,N_11440,N_13756);
and UO_309 (O_309,N_13886,N_14545);
nor UO_310 (O_310,N_11701,N_10248);
nor UO_311 (O_311,N_14830,N_14284);
and UO_312 (O_312,N_14766,N_14772);
nand UO_313 (O_313,N_14248,N_11669);
and UO_314 (O_314,N_11218,N_12173);
nand UO_315 (O_315,N_10602,N_12319);
nor UO_316 (O_316,N_13750,N_14051);
or UO_317 (O_317,N_12610,N_13864);
nand UO_318 (O_318,N_10354,N_12828);
nor UO_319 (O_319,N_10279,N_13037);
and UO_320 (O_320,N_11646,N_11754);
and UO_321 (O_321,N_10992,N_13877);
nand UO_322 (O_322,N_10132,N_12582);
nor UO_323 (O_323,N_12680,N_11566);
nor UO_324 (O_324,N_14517,N_11942);
nor UO_325 (O_325,N_11238,N_10179);
nand UO_326 (O_326,N_14134,N_12397);
xor UO_327 (O_327,N_10070,N_11970);
or UO_328 (O_328,N_10076,N_10772);
or UO_329 (O_329,N_14804,N_10390);
xnor UO_330 (O_330,N_12460,N_13660);
nand UO_331 (O_331,N_12092,N_11461);
or UO_332 (O_332,N_12022,N_13830);
and UO_333 (O_333,N_14698,N_10607);
nor UO_334 (O_334,N_14935,N_11874);
and UO_335 (O_335,N_12528,N_14628);
nor UO_336 (O_336,N_13136,N_13385);
nor UO_337 (O_337,N_12505,N_12502);
nor UO_338 (O_338,N_13831,N_11077);
nor UO_339 (O_339,N_12569,N_11785);
and UO_340 (O_340,N_14523,N_12595);
or UO_341 (O_341,N_10840,N_12175);
nand UO_342 (O_342,N_14116,N_11863);
or UO_343 (O_343,N_10330,N_12975);
xnor UO_344 (O_344,N_11177,N_13649);
or UO_345 (O_345,N_13614,N_10338);
nor UO_346 (O_346,N_13299,N_10066);
and UO_347 (O_347,N_13872,N_10172);
nand UO_348 (O_348,N_12153,N_13467);
and UO_349 (O_349,N_10851,N_11099);
xor UO_350 (O_350,N_12344,N_10932);
nand UO_351 (O_351,N_13107,N_12365);
or UO_352 (O_352,N_10953,N_12401);
and UO_353 (O_353,N_14182,N_10180);
and UO_354 (O_354,N_12573,N_10540);
nand UO_355 (O_355,N_14533,N_14927);
xor UO_356 (O_356,N_10505,N_10573);
or UO_357 (O_357,N_11627,N_14043);
xnor UO_358 (O_358,N_13995,N_12521);
or UO_359 (O_359,N_14374,N_14884);
nor UO_360 (O_360,N_14012,N_11610);
or UO_361 (O_361,N_14819,N_13072);
or UO_362 (O_362,N_10163,N_14743);
nand UO_363 (O_363,N_12820,N_11462);
and UO_364 (O_364,N_11327,N_14158);
and UO_365 (O_365,N_14107,N_12774);
nand UO_366 (O_366,N_10061,N_10369);
and UO_367 (O_367,N_14122,N_10474);
nor UO_368 (O_368,N_14713,N_11012);
or UO_369 (O_369,N_14846,N_11090);
and UO_370 (O_370,N_14805,N_10082);
or UO_371 (O_371,N_11002,N_14562);
nor UO_372 (O_372,N_10456,N_10304);
nor UO_373 (O_373,N_13722,N_12437);
or UO_374 (O_374,N_11833,N_13469);
nand UO_375 (O_375,N_10620,N_14137);
nor UO_376 (O_376,N_13383,N_13683);
and UO_377 (O_377,N_14656,N_10667);
and UO_378 (O_378,N_11222,N_14421);
and UO_379 (O_379,N_11872,N_13706);
and UO_380 (O_380,N_12915,N_13863);
or UO_381 (O_381,N_12869,N_10069);
nand UO_382 (O_382,N_11160,N_11131);
nand UO_383 (O_383,N_14226,N_14077);
nor UO_384 (O_384,N_10157,N_12042);
or UO_385 (O_385,N_12109,N_10749);
nor UO_386 (O_386,N_13226,N_13745);
nor UO_387 (O_387,N_10251,N_14507);
nand UO_388 (O_388,N_13320,N_11990);
nor UO_389 (O_389,N_11348,N_11987);
and UO_390 (O_390,N_13182,N_14916);
or UO_391 (O_391,N_13607,N_13719);
and UO_392 (O_392,N_10181,N_10318);
nor UO_393 (O_393,N_11577,N_10794);
nor UO_394 (O_394,N_12412,N_12385);
or UO_395 (O_395,N_10117,N_11006);
or UO_396 (O_396,N_10935,N_13790);
or UO_397 (O_397,N_13366,N_12937);
nor UO_398 (O_398,N_14117,N_10842);
and UO_399 (O_399,N_14468,N_13825);
nand UO_400 (O_400,N_10256,N_13720);
nand UO_401 (O_401,N_10879,N_12178);
nor UO_402 (O_402,N_13715,N_10766);
or UO_403 (O_403,N_14221,N_12801);
and UO_404 (O_404,N_12276,N_12880);
nand UO_405 (O_405,N_12228,N_12266);
nand UO_406 (O_406,N_13691,N_12668);
or UO_407 (O_407,N_10864,N_14657);
or UO_408 (O_408,N_10099,N_14824);
and UO_409 (O_409,N_12254,N_13882);
or UO_410 (O_410,N_12245,N_14693);
nor UO_411 (O_411,N_11054,N_13773);
nor UO_412 (O_412,N_13490,N_11549);
nand UO_413 (O_413,N_10149,N_12691);
or UO_414 (O_414,N_11897,N_11634);
and UO_415 (O_415,N_13984,N_11561);
or UO_416 (O_416,N_13871,N_13281);
nor UO_417 (O_417,N_10432,N_14309);
or UO_418 (O_418,N_10972,N_14633);
or UO_419 (O_419,N_11992,N_13236);
nor UO_420 (O_420,N_14497,N_11550);
and UO_421 (O_421,N_10596,N_13221);
or UO_422 (O_422,N_12032,N_14461);
or UO_423 (O_423,N_13454,N_14073);
and UO_424 (O_424,N_14899,N_13606);
and UO_425 (O_425,N_11078,N_11967);
nand UO_426 (O_426,N_11601,N_14714);
or UO_427 (O_427,N_14131,N_12294);
nand UO_428 (O_428,N_10334,N_12504);
or UO_429 (O_429,N_13889,N_11792);
nand UO_430 (O_430,N_14385,N_11641);
and UO_431 (O_431,N_13224,N_12679);
and UO_432 (O_432,N_14071,N_14254);
or UO_433 (O_433,N_13010,N_14013);
and UO_434 (O_434,N_12552,N_10802);
or UO_435 (O_435,N_12050,N_10593);
and UO_436 (O_436,N_14997,N_13478);
and UO_437 (O_437,N_11896,N_11704);
nor UO_438 (O_438,N_10502,N_14908);
nand UO_439 (O_439,N_13322,N_14210);
nand UO_440 (O_440,N_11507,N_12809);
nand UO_441 (O_441,N_12626,N_12832);
nor UO_442 (O_442,N_13402,N_12478);
nor UO_443 (O_443,N_11486,N_13233);
nand UO_444 (O_444,N_13415,N_11824);
or UO_445 (O_445,N_10485,N_13553);
nand UO_446 (O_446,N_12361,N_10022);
and UO_447 (O_447,N_10130,N_14198);
nor UO_448 (O_448,N_10966,N_12688);
or UO_449 (O_449,N_13911,N_13041);
nand UO_450 (O_450,N_13271,N_13666);
or UO_451 (O_451,N_12693,N_10898);
nand UO_452 (O_452,N_10536,N_14532);
and UO_453 (O_453,N_10190,N_14752);
nand UO_454 (O_454,N_10046,N_13357);
nand UO_455 (O_455,N_10122,N_14173);
nor UO_456 (O_456,N_11821,N_12147);
nand UO_457 (O_457,N_10743,N_14389);
nand UO_458 (O_458,N_11826,N_14711);
nand UO_459 (O_459,N_12093,N_12019);
and UO_460 (O_460,N_12325,N_10940);
or UO_461 (O_461,N_13945,N_12686);
and UO_462 (O_462,N_14350,N_14647);
xor UO_463 (O_463,N_14923,N_11535);
or UO_464 (O_464,N_13949,N_11789);
nor UO_465 (O_465,N_14106,N_14269);
nor UO_466 (O_466,N_13382,N_14006);
nor UO_467 (O_467,N_11432,N_12632);
nand UO_468 (O_468,N_11913,N_10013);
nand UO_469 (O_469,N_11584,N_13724);
or UO_470 (O_470,N_14929,N_10662);
and UO_471 (O_471,N_11637,N_12844);
or UO_472 (O_472,N_11575,N_13180);
nor UO_473 (O_473,N_11526,N_14885);
nand UO_474 (O_474,N_14531,N_10071);
nor UO_475 (O_475,N_10928,N_14863);
nand UO_476 (O_476,N_12788,N_12739);
and UO_477 (O_477,N_14759,N_13613);
or UO_478 (O_478,N_12705,N_13770);
nor UO_479 (O_479,N_11943,N_10367);
nand UO_480 (O_480,N_13256,N_10212);
nand UO_481 (O_481,N_13842,N_10314);
and UO_482 (O_482,N_11553,N_12903);
and UO_483 (O_483,N_12394,N_12973);
and UO_484 (O_484,N_11071,N_10508);
or UO_485 (O_485,N_14047,N_14347);
or UO_486 (O_486,N_14636,N_12104);
nor UO_487 (O_487,N_10771,N_11877);
nand UO_488 (O_488,N_10833,N_11195);
and UO_489 (O_489,N_11624,N_14806);
or UO_490 (O_490,N_10087,N_13596);
nor UO_491 (O_491,N_12953,N_13812);
and UO_492 (O_492,N_13317,N_11998);
or UO_493 (O_493,N_13848,N_11554);
and UO_494 (O_494,N_13138,N_12010);
nor UO_495 (O_495,N_13580,N_12351);
or UO_496 (O_496,N_14428,N_10889);
nor UO_497 (O_497,N_12687,N_13421);
nand UO_498 (O_498,N_13489,N_12240);
nand UO_499 (O_499,N_14289,N_10374);
nand UO_500 (O_500,N_11940,N_10821);
nand UO_501 (O_501,N_11278,N_13154);
and UO_502 (O_502,N_14201,N_13424);
nor UO_503 (O_503,N_12163,N_11630);
nand UO_504 (O_504,N_13339,N_10608);
nor UO_505 (O_505,N_12111,N_14617);
nand UO_506 (O_506,N_13594,N_12354);
or UO_507 (O_507,N_10100,N_10583);
and UO_508 (O_508,N_12296,N_14891);
or UO_509 (O_509,N_13493,N_12619);
or UO_510 (O_510,N_13852,N_14143);
nor UO_511 (O_511,N_14089,N_10910);
nor UO_512 (O_512,N_10388,N_13711);
nand UO_513 (O_513,N_12230,N_12721);
or UO_514 (O_514,N_12858,N_10732);
or UO_515 (O_515,N_11121,N_12404);
or UO_516 (O_516,N_13737,N_11230);
nor UO_517 (O_517,N_14651,N_13568);
and UO_518 (O_518,N_12747,N_12625);
or UO_519 (O_519,N_10322,N_14977);
nor UO_520 (O_520,N_13488,N_11428);
nand UO_521 (O_521,N_12896,N_10878);
nor UO_522 (O_522,N_10056,N_12885);
nand UO_523 (O_523,N_10769,N_10218);
nand UO_524 (O_524,N_13462,N_13482);
xnor UO_525 (O_525,N_14735,N_14103);
and UO_526 (O_526,N_14816,N_14687);
or UO_527 (O_527,N_11774,N_13908);
nand UO_528 (O_528,N_11066,N_12764);
and UO_529 (O_529,N_10913,N_10199);
and UO_530 (O_530,N_10591,N_10981);
or UO_531 (O_531,N_10577,N_10707);
or UO_532 (O_532,N_10993,N_12041);
or UO_533 (O_533,N_14156,N_10193);
nor UO_534 (O_534,N_14575,N_14560);
nor UO_535 (O_535,N_13575,N_13900);
nor UO_536 (O_536,N_11315,N_11059);
nor UO_537 (O_537,N_10349,N_11154);
or UO_538 (O_538,N_14998,N_14469);
or UO_539 (O_539,N_11620,N_11888);
or UO_540 (O_540,N_13029,N_13270);
nand UO_541 (O_541,N_11088,N_10226);
xnor UO_542 (O_542,N_12622,N_12060);
nor UO_543 (O_543,N_11677,N_10503);
or UO_544 (O_544,N_11251,N_13054);
and UO_545 (O_545,N_12805,N_11608);
nand UO_546 (O_546,N_11139,N_13565);
nor UO_547 (O_547,N_11076,N_10306);
nor UO_548 (O_548,N_14605,N_11794);
nand UO_549 (O_549,N_10088,N_10874);
and UO_550 (O_550,N_13806,N_12728);
and UO_551 (O_551,N_14642,N_13986);
nor UO_552 (O_552,N_14758,N_13555);
nor UO_553 (O_553,N_13861,N_12631);
or UO_554 (O_554,N_11611,N_10290);
nor UO_555 (O_555,N_12555,N_11927);
and UO_556 (O_556,N_13480,N_12018);
nand UO_557 (O_557,N_14473,N_12199);
or UO_558 (O_558,N_13083,N_14061);
nor UO_559 (O_559,N_11808,N_13134);
and UO_560 (O_560,N_13081,N_11707);
and UO_561 (O_561,N_12857,N_12715);
nor UO_562 (O_562,N_14381,N_11410);
or UO_563 (O_563,N_11838,N_13954);
xnor UO_564 (O_564,N_13056,N_13332);
nor UO_565 (O_565,N_12040,N_14465);
nand UO_566 (O_566,N_11081,N_13631);
and UO_567 (O_567,N_13426,N_12796);
or UO_568 (O_568,N_12299,N_11380);
or UO_569 (O_569,N_12690,N_12246);
nor UO_570 (O_570,N_10731,N_14433);
nand UO_571 (O_571,N_14050,N_12780);
or UO_572 (O_572,N_11968,N_10381);
and UO_573 (O_573,N_12278,N_12692);
nand UO_574 (O_574,N_11632,N_13838);
nor UO_575 (O_575,N_11687,N_12672);
nor UO_576 (O_576,N_10387,N_10113);
nor UO_577 (O_577,N_11313,N_13340);
nand UO_578 (O_578,N_13875,N_12291);
and UO_579 (O_579,N_12152,N_12122);
nand UO_580 (O_580,N_11654,N_11211);
nor UO_581 (O_581,N_13085,N_14205);
nand UO_582 (O_582,N_12737,N_10885);
and UO_583 (O_583,N_14695,N_12298);
nor UO_584 (O_584,N_10054,N_10024);
or UO_585 (O_585,N_11581,N_11895);
nand UO_586 (O_586,N_12697,N_14390);
and UO_587 (O_587,N_11053,N_12223);
nor UO_588 (O_588,N_13637,N_14730);
xnor UO_589 (O_589,N_11595,N_14224);
or UO_590 (O_590,N_14645,N_13049);
and UO_591 (O_591,N_10938,N_13771);
xnor UO_592 (O_592,N_14485,N_12306);
and UO_593 (O_593,N_10351,N_10384);
and UO_594 (O_594,N_10039,N_13168);
nor UO_595 (O_595,N_11276,N_14558);
or UO_596 (O_596,N_10498,N_14776);
nand UO_597 (O_597,N_13021,N_13303);
and UO_598 (O_598,N_13718,N_14875);
nor UO_599 (O_599,N_10983,N_10739);
nand UO_600 (O_600,N_11882,N_12641);
nor UO_601 (O_601,N_10990,N_11105);
and UO_602 (O_602,N_13269,N_12549);
and UO_603 (O_603,N_10133,N_11008);
xor UO_604 (O_604,N_12719,N_10435);
or UO_605 (O_605,N_11357,N_13185);
nor UO_606 (O_606,N_13429,N_10353);
nor UO_607 (O_607,N_14190,N_14400);
nand UO_608 (O_608,N_14471,N_14958);
nor UO_609 (O_609,N_11894,N_11556);
nand UO_610 (O_610,N_11267,N_12749);
nand UO_611 (O_611,N_13245,N_14278);
nor UO_612 (O_612,N_11080,N_10142);
and UO_613 (O_613,N_13677,N_10266);
and UO_614 (O_614,N_11344,N_13460);
and UO_615 (O_615,N_14644,N_14496);
nor UO_616 (O_616,N_14466,N_14585);
nor UO_617 (O_617,N_12905,N_12479);
or UO_618 (O_618,N_12509,N_11648);
or UO_619 (O_619,N_13934,N_14429);
nand UO_620 (O_620,N_14108,N_14133);
and UO_621 (O_621,N_13618,N_13187);
nand UO_622 (O_622,N_11084,N_13215);
nand UO_623 (O_623,N_13498,N_10728);
or UO_624 (O_624,N_11722,N_13638);
or UO_625 (O_625,N_10473,N_13662);
and UO_626 (O_626,N_13811,N_13858);
and UO_627 (O_627,N_13470,N_12432);
nor UO_628 (O_628,N_14397,N_14394);
and UO_629 (O_629,N_14148,N_11856);
nor UO_630 (O_630,N_14065,N_14890);
nor UO_631 (O_631,N_11706,N_12997);
nor UO_632 (O_632,N_10926,N_10614);
or UO_633 (O_633,N_12362,N_10929);
nand UO_634 (O_634,N_11341,N_10264);
and UO_635 (O_635,N_14281,N_11997);
or UO_636 (O_636,N_13869,N_10994);
nor UO_637 (O_637,N_12961,N_12965);
nand UO_638 (O_638,N_10419,N_11529);
nor UO_639 (O_639,N_14002,N_13116);
nand UO_640 (O_640,N_12059,N_13115);
and UO_641 (O_641,N_12750,N_13802);
or UO_642 (O_642,N_10927,N_10921);
nand UO_643 (O_643,N_11585,N_10923);
and UO_644 (O_644,N_13255,N_12211);
or UO_645 (O_645,N_11188,N_11130);
or UO_646 (O_646,N_12444,N_11424);
and UO_647 (O_647,N_13369,N_10859);
and UO_648 (O_648,N_13242,N_10019);
nor UO_649 (O_649,N_14709,N_12894);
xor UO_650 (O_650,N_12224,N_13479);
nor UO_651 (O_651,N_11097,N_14257);
nor UO_652 (O_652,N_11475,N_13152);
nor UO_653 (O_653,N_13374,N_14506);
nor UO_654 (O_654,N_10895,N_12119);
nand UO_655 (O_655,N_10258,N_13465);
and UO_656 (O_656,N_12003,N_12188);
or UO_657 (O_657,N_13933,N_11830);
nor UO_658 (O_658,N_14227,N_14955);
nor UO_659 (O_659,N_12675,N_11587);
nor UO_660 (O_660,N_14392,N_14455);
nor UO_661 (O_661,N_10555,N_11718);
nor UO_662 (O_662,N_10469,N_12293);
and UO_663 (O_663,N_13624,N_13087);
nor UO_664 (O_664,N_10829,N_12900);
xnor UO_665 (O_665,N_11730,N_11450);
nor UO_666 (O_666,N_12850,N_14016);
and UO_667 (O_667,N_10489,N_12352);
nand UO_668 (O_668,N_11988,N_13938);
nand UO_669 (O_669,N_10422,N_11829);
nor UO_670 (O_670,N_12930,N_10340);
nand UO_671 (O_671,N_14262,N_13985);
or UO_672 (O_672,N_12182,N_13195);
or UO_673 (O_673,N_13744,N_11638);
and UO_674 (O_674,N_11346,N_12094);
and UO_675 (O_675,N_12203,N_11918);
and UO_676 (O_676,N_11702,N_10359);
and UO_677 (O_677,N_14773,N_11120);
and UO_678 (O_678,N_11254,N_13093);
and UO_679 (O_679,N_14356,N_12817);
and UO_680 (O_680,N_14482,N_12096);
nor UO_681 (O_681,N_10706,N_10043);
and UO_682 (O_682,N_12058,N_13632);
nor UO_683 (O_683,N_10162,N_14439);
nand UO_684 (O_684,N_12226,N_14611);
nand UO_685 (O_685,N_10143,N_10975);
or UO_686 (O_686,N_13169,N_10712);
or UO_687 (O_687,N_11819,N_13630);
nand UO_688 (O_688,N_13727,N_10623);
nand UO_689 (O_689,N_12991,N_12048);
or UO_690 (O_690,N_13859,N_11901);
xnor UO_691 (O_691,N_10005,N_14808);
and UO_692 (O_692,N_10724,N_10693);
and UO_693 (O_693,N_10843,N_10616);
nand UO_694 (O_694,N_12483,N_14383);
xor UO_695 (O_695,N_10084,N_12511);
nor UO_696 (O_696,N_13381,N_13651);
nor UO_697 (O_697,N_14627,N_10599);
or UO_698 (O_698,N_10204,N_13671);
nor UO_699 (O_699,N_12139,N_13562);
or UO_700 (O_700,N_14689,N_13079);
nor UO_701 (O_701,N_13696,N_12279);
nand UO_702 (O_702,N_11471,N_11282);
or UO_703 (O_703,N_14780,N_12902);
nor UO_704 (O_704,N_12127,N_12043);
nor UO_705 (O_705,N_10664,N_10145);
and UO_706 (O_706,N_12945,N_12669);
nand UO_707 (O_707,N_12455,N_13902);
nand UO_708 (O_708,N_10067,N_13994);
nand UO_709 (O_709,N_11263,N_14181);
and UO_710 (O_710,N_10109,N_12417);
and UO_711 (O_711,N_10654,N_12855);
and UO_712 (O_712,N_11360,N_10615);
or UO_713 (O_713,N_10775,N_10465);
nand UO_714 (O_714,N_12320,N_10227);
nor UO_715 (O_715,N_12978,N_11488);
and UO_716 (O_716,N_12984,N_11144);
and UO_717 (O_717,N_12384,N_13201);
and UO_718 (O_718,N_12766,N_14099);
or UO_719 (O_719,N_11215,N_13389);
nand UO_720 (O_720,N_14299,N_14716);
xnor UO_721 (O_721,N_14462,N_12037);
xnor UO_722 (O_722,N_13220,N_10803);
nor UO_723 (O_723,N_13006,N_14749);
or UO_724 (O_724,N_12508,N_10735);
nor UO_725 (O_725,N_11135,N_14321);
nor UO_726 (O_726,N_12758,N_13809);
and UO_727 (O_727,N_13784,N_14279);
xor UO_728 (O_728,N_14094,N_13111);
nor UO_729 (O_729,N_10458,N_11757);
nor UO_730 (O_730,N_12403,N_14539);
xor UO_731 (O_731,N_12186,N_11564);
nor UO_732 (O_732,N_13504,N_14352);
nor UO_733 (O_733,N_14513,N_12210);
or UO_734 (O_734,N_11599,N_12020);
nor UO_735 (O_735,N_12185,N_10175);
nor UO_736 (O_736,N_13901,N_10755);
or UO_737 (O_737,N_11724,N_13629);
and UO_738 (O_738,N_10671,N_10240);
nor UO_739 (O_739,N_10727,N_11482);
nor UO_740 (O_740,N_10361,N_12292);
or UO_741 (O_741,N_14423,N_11598);
or UO_742 (O_742,N_10822,N_11555);
and UO_743 (O_743,N_13420,N_12440);
and UO_744 (O_744,N_12443,N_14258);
nand UO_745 (O_745,N_10278,N_10198);
nand UO_746 (O_746,N_12714,N_11666);
nand UO_747 (O_747,N_14722,N_10116);
or UO_748 (O_748,N_11732,N_11062);
nand UO_749 (O_749,N_11676,N_14267);
nor UO_750 (O_750,N_13512,N_10303);
nor UO_751 (O_751,N_13432,N_12169);
and UO_752 (O_752,N_10128,N_11444);
nor UO_753 (O_753,N_14796,N_10187);
nor UO_754 (O_754,N_10764,N_12016);
nor UO_755 (O_755,N_11393,N_11855);
nor UO_756 (O_756,N_14993,N_10965);
or UO_757 (O_757,N_10431,N_10207);
nor UO_758 (O_758,N_13059,N_11936);
or UO_759 (O_759,N_10000,N_11814);
or UO_760 (O_760,N_14854,N_13212);
nand UO_761 (O_761,N_12570,N_13523);
nor UO_762 (O_762,N_10339,N_11300);
or UO_763 (O_763,N_10969,N_14793);
and UO_764 (O_764,N_11051,N_12200);
nor UO_765 (O_765,N_14547,N_12027);
nor UO_766 (O_766,N_11166,N_13268);
or UO_767 (O_767,N_12372,N_14030);
xnor UO_768 (O_768,N_10900,N_14318);
nand UO_769 (O_769,N_12895,N_13321);
or UO_770 (O_770,N_13595,N_14220);
and UO_771 (O_771,N_11586,N_10734);
nand UO_772 (O_772,N_14615,N_14364);
and UO_773 (O_773,N_12834,N_11781);
or UO_774 (O_774,N_13893,N_14525);
or UO_775 (O_775,N_13761,N_10557);
nand UO_776 (O_776,N_14972,N_11502);
and UO_777 (O_777,N_10861,N_14865);
and UO_778 (O_778,N_10454,N_10127);
and UO_779 (O_779,N_11381,N_11416);
nor UO_780 (O_780,N_13350,N_14204);
nor UO_781 (O_781,N_12332,N_13345);
nand UO_782 (O_782,N_11285,N_13702);
and UO_783 (O_783,N_10427,N_14164);
or UO_784 (O_784,N_14136,N_14791);
or UO_785 (O_785,N_12793,N_14212);
nand UO_786 (O_786,N_10140,N_11474);
and UO_787 (O_787,N_11772,N_11437);
xor UO_788 (O_788,N_12428,N_13044);
and UO_789 (O_789,N_10302,N_12559);
nor UO_790 (O_790,N_14017,N_13050);
nand UO_791 (O_791,N_11612,N_14192);
and UO_792 (O_792,N_14682,N_13726);
nand UO_793 (O_793,N_12017,N_10564);
nor UO_794 (O_794,N_11796,N_13681);
nand UO_795 (O_795,N_14045,N_12252);
and UO_796 (O_796,N_10401,N_10483);
or UO_797 (O_797,N_12255,N_11760);
and UO_798 (O_798,N_13936,N_14982);
nor UO_799 (O_799,N_12057,N_11858);
nor UO_800 (O_800,N_12086,N_12685);
or UO_801 (O_801,N_14437,N_10356);
nor UO_802 (O_802,N_14736,N_10725);
nand UO_803 (O_803,N_12898,N_13119);
nand UO_804 (O_804,N_13826,N_14330);
nand UO_805 (O_805,N_13398,N_10200);
nor UO_806 (O_806,N_10478,N_13450);
or UO_807 (O_807,N_13485,N_10971);
and UO_808 (O_808,N_10259,N_13937);
or UO_809 (O_809,N_11343,N_11273);
or UO_810 (O_810,N_11606,N_13202);
or UO_811 (O_811,N_12363,N_10466);
nor UO_812 (O_812,N_12722,N_10665);
nand UO_813 (O_813,N_11185,N_14936);
and UO_814 (O_814,N_12892,N_12441);
or UO_815 (O_815,N_14576,N_12818);
nor UO_816 (O_816,N_13914,N_12421);
and UO_817 (O_817,N_14588,N_14306);
nand UO_818 (O_818,N_13063,N_10471);
and UO_819 (O_819,N_10123,N_14680);
and UO_820 (O_820,N_12067,N_12258);
and UO_821 (O_821,N_10377,N_11775);
nor UO_822 (O_822,N_11132,N_12525);
or UO_823 (O_823,N_14066,N_13316);
or UO_824 (O_824,N_11311,N_13648);
nand UO_825 (O_825,N_10792,N_12174);
nor UO_826 (O_826,N_12410,N_13150);
nand UO_827 (O_827,N_11212,N_13471);
nor UO_828 (O_828,N_13315,N_12578);
or UO_829 (O_829,N_13599,N_13918);
or UO_830 (O_830,N_11682,N_14503);
and UO_831 (O_831,N_10915,N_13541);
nor UO_832 (O_832,N_10692,N_13639);
nor UO_833 (O_833,N_14603,N_12453);
nor UO_834 (O_834,N_14620,N_12280);
nor UO_835 (O_835,N_13058,N_14731);
nor UO_836 (O_836,N_14011,N_11973);
xor UO_837 (O_837,N_10297,N_10053);
xnor UO_838 (O_838,N_13556,N_10778);
nor UO_839 (O_839,N_14755,N_10094);
xor UO_840 (O_840,N_11411,N_13500);
nor UO_841 (O_841,N_10428,N_10810);
or UO_842 (O_842,N_12532,N_13854);
and UO_843 (O_843,N_12489,N_12974);
and UO_844 (O_844,N_13304,N_13008);
and UO_845 (O_845,N_11199,N_14609);
or UO_846 (O_846,N_14515,N_12634);
nand UO_847 (O_847,N_14632,N_14845);
nand UO_848 (O_848,N_11023,N_13697);
xor UO_849 (O_849,N_14444,N_12202);
nor UO_850 (O_850,N_13685,N_10048);
nor UO_851 (O_851,N_13833,N_13675);
nand UO_852 (O_852,N_13277,N_10413);
or UO_853 (O_853,N_10595,N_11800);
nand UO_854 (O_854,N_10211,N_13153);
and UO_855 (O_855,N_10051,N_13030);
and UO_856 (O_856,N_14582,N_11221);
nand UO_857 (O_857,N_11947,N_11141);
and UO_858 (O_858,N_10410,N_14327);
nand UO_859 (O_859,N_13839,N_12338);
xnor UO_860 (O_860,N_13231,N_11664);
or UO_861 (O_861,N_14096,N_13785);
or UO_862 (O_862,N_14896,N_13729);
and UO_863 (O_863,N_13957,N_13679);
or UO_864 (O_864,N_14762,N_10824);
or UO_865 (O_865,N_11111,N_12681);
and UO_866 (O_866,N_13966,N_13647);
or UO_867 (O_867,N_11074,N_11787);
nand UO_868 (O_868,N_13376,N_11622);
nor UO_869 (O_869,N_14767,N_10561);
and UO_870 (O_870,N_12879,N_12527);
nor UO_871 (O_871,N_14876,N_12846);
nand UO_872 (O_872,N_11459,N_13354);
nor UO_873 (O_873,N_13434,N_13730);
nor UO_874 (O_874,N_11093,N_10908);
or UO_875 (O_875,N_10903,N_13701);
or UO_876 (O_876,N_11873,N_12999);
or UO_877 (O_877,N_14683,N_12301);
or UO_878 (O_878,N_11532,N_12803);
or UO_879 (O_879,N_13019,N_10780);
xor UO_880 (O_880,N_14484,N_14159);
nand UO_881 (O_881,N_10345,N_13557);
nor UO_882 (O_882,N_12860,N_12854);
and UO_883 (O_883,N_12544,N_14754);
or UO_884 (O_884,N_13944,N_11513);
nor UO_885 (O_885,N_12498,N_13131);
nor UO_886 (O_886,N_13228,N_14193);
nor UO_887 (O_887,N_14274,N_11201);
nand UO_888 (O_888,N_10487,N_14768);
nand UO_889 (O_889,N_11588,N_10030);
or UO_890 (O_890,N_11339,N_13887);
or UO_891 (O_891,N_11740,N_14697);
and UO_892 (O_892,N_11415,N_10565);
and UO_893 (O_893,N_14288,N_13690);
or UO_894 (O_894,N_10495,N_11158);
and UO_895 (O_895,N_10569,N_13173);
or UO_896 (O_896,N_12405,N_11840);
nor UO_897 (O_897,N_13284,N_14740);
nand UO_898 (O_898,N_10224,N_10787);
nand UO_899 (O_899,N_11489,N_12684);
xor UO_900 (O_900,N_13476,N_11196);
and UO_901 (O_901,N_10205,N_14459);
or UO_902 (O_902,N_11880,N_13207);
or UO_903 (O_903,N_14033,N_11578);
or UO_904 (O_904,N_11209,N_10228);
nand UO_905 (O_905,N_12315,N_13664);
nor UO_906 (O_906,N_12724,N_13517);
or UO_907 (O_907,N_11296,N_14571);
and UO_908 (O_908,N_13400,N_10420);
nand UO_909 (O_909,N_13952,N_13760);
and UO_910 (O_910,N_10378,N_11019);
nand UO_911 (O_911,N_11048,N_14634);
or UO_912 (O_912,N_12099,N_14665);
or UO_913 (O_913,N_10329,N_12804);
nor UO_914 (O_914,N_14831,N_12138);
nand UO_915 (O_915,N_13130,N_14395);
or UO_916 (O_916,N_12463,N_13686);
nor UO_917 (O_917,N_10441,N_14502);
and UO_918 (O_918,N_13456,N_11745);
and UO_919 (O_919,N_11652,N_10403);
or UO_920 (O_920,N_13644,N_10570);
nor UO_921 (O_921,N_14995,N_13634);
or UO_922 (O_922,N_10399,N_14602);
nand UO_923 (O_923,N_13147,N_13909);
nor UO_924 (O_924,N_14255,N_14631);
or UO_925 (O_925,N_12089,N_12698);
nor UO_926 (O_926,N_14895,N_12767);
and UO_927 (O_927,N_12007,N_10366);
nor UO_928 (O_928,N_11376,N_13204);
or UO_929 (O_929,N_11694,N_10690);
nor UO_930 (O_930,N_14639,N_14969);
nor UO_931 (O_931,N_10836,N_12227);
nand UO_932 (O_932,N_11436,N_13530);
or UO_933 (O_933,N_12656,N_10660);
nor UO_934 (O_934,N_10430,N_10479);
and UO_935 (O_935,N_13290,N_12906);
or UO_936 (O_936,N_13915,N_11651);
nor UO_937 (O_937,N_10085,N_12342);
or UO_938 (O_938,N_13045,N_14354);
and UO_939 (O_939,N_12942,N_12442);
and UO_940 (O_940,N_10768,N_11068);
and UO_941 (O_941,N_12928,N_11458);
or UO_942 (O_942,N_11567,N_13405);
and UO_943 (O_943,N_10214,N_11481);
or UO_944 (O_944,N_10288,N_11713);
nand UO_945 (O_945,N_10974,N_12464);
nand UO_946 (O_946,N_14296,N_12515);
nand UO_947 (O_947,N_14524,N_13279);
nor UO_948 (O_948,N_13208,N_10423);
and UO_949 (O_949,N_11835,N_14119);
nand UO_950 (O_950,N_10718,N_14950);
and UO_951 (O_951,N_13881,N_10447);
nand UO_952 (O_952,N_13891,N_12378);
or UO_953 (O_953,N_11503,N_12015);
and UO_954 (O_954,N_14285,N_12604);
nor UO_955 (O_955,N_11429,N_12731);
or UO_956 (O_956,N_11552,N_11056);
nor UO_957 (O_957,N_12710,N_11644);
nor UO_958 (O_958,N_13813,N_11665);
or UO_959 (O_959,N_14710,N_10375);
xor UO_960 (O_960,N_11969,N_10342);
and UO_961 (O_961,N_12467,N_10958);
and UO_962 (O_962,N_11249,N_11469);
nor UO_963 (O_963,N_12103,N_12674);
and UO_964 (O_964,N_14834,N_14844);
or UO_965 (O_965,N_14062,N_13109);
nand UO_966 (O_966,N_10865,N_10701);
nand UO_967 (O_967,N_12474,N_10372);
or UO_968 (O_968,N_12275,N_11152);
or UO_969 (O_969,N_14250,N_11910);
and UO_970 (O_970,N_10216,N_10037);
or UO_971 (O_971,N_13211,N_14500);
and UO_972 (O_972,N_13355,N_13663);
or UO_973 (O_973,N_14590,N_12377);
and UO_974 (O_974,N_12825,N_10544);
nand UO_975 (O_975,N_10450,N_10622);
nor UO_976 (O_976,N_11698,N_14607);
or UO_977 (O_977,N_11514,N_11744);
nor UO_978 (O_978,N_14699,N_11426);
and UO_979 (O_979,N_13592,N_14619);
nand UO_980 (O_980,N_10870,N_13547);
and UO_981 (O_981,N_12125,N_12348);
and UO_982 (O_982,N_13218,N_10587);
nor UO_983 (O_983,N_10782,N_13808);
and UO_984 (O_984,N_14938,N_14996);
nor UO_985 (O_985,N_12986,N_12494);
xor UO_986 (O_986,N_13425,N_10681);
and UO_987 (O_987,N_14733,N_11836);
nand UO_988 (O_988,N_12189,N_11001);
nand UO_989 (O_989,N_14856,N_13053);
and UO_990 (O_990,N_11442,N_10936);
or UO_991 (O_991,N_11013,N_11631);
or UO_992 (O_992,N_14150,N_11903);
nor UO_993 (O_993,N_10675,N_13767);
nor UO_994 (O_994,N_12996,N_11377);
or UO_995 (O_995,N_11671,N_13175);
and UO_996 (O_996,N_13065,N_10507);
or UO_997 (O_997,N_13943,N_10759);
nand UO_998 (O_998,N_12070,N_10605);
and UO_999 (O_999,N_11999,N_14165);
or UO_1000 (O_1000,N_13920,N_12530);
nor UO_1001 (O_1001,N_12346,N_12072);
or UO_1002 (O_1002,N_12083,N_14493);
or UO_1003 (O_1003,N_10995,N_11959);
xor UO_1004 (O_1004,N_10814,N_11495);
nand UO_1005 (O_1005,N_11384,N_14037);
and UO_1006 (O_1006,N_14869,N_11948);
or UO_1007 (O_1007,N_12537,N_13919);
nand UO_1008 (O_1008,N_14189,N_13930);
or UO_1009 (O_1009,N_10488,N_11464);
nor UO_1010 (O_1010,N_13197,N_14897);
and UO_1011 (O_1011,N_11843,N_10397);
and UO_1012 (O_1012,N_10131,N_11129);
nor UO_1013 (O_1013,N_10272,N_14237);
and UO_1014 (O_1014,N_10552,N_12934);
or UO_1015 (O_1015,N_13948,N_13235);
and UO_1016 (O_1016,N_14329,N_14216);
and UO_1017 (O_1017,N_11394,N_12654);
nand UO_1018 (O_1018,N_12333,N_14375);
and UO_1019 (O_1019,N_10136,N_10134);
nor UO_1020 (O_1020,N_12821,N_12887);
nor UO_1021 (O_1021,N_10060,N_13528);
and UO_1022 (O_1022,N_11512,N_13074);
nor UO_1023 (O_1023,N_12655,N_14534);
nand UO_1024 (O_1024,N_13330,N_13126);
nor UO_1025 (O_1025,N_14921,N_14067);
and UO_1026 (O_1026,N_11996,N_11100);
nand UO_1027 (O_1027,N_14346,N_10751);
nor UO_1028 (O_1028,N_11033,N_10906);
nor UO_1029 (O_1029,N_13200,N_10527);
nand UO_1030 (O_1030,N_14900,N_12636);
nand UO_1031 (O_1031,N_10520,N_10846);
nand UO_1032 (O_1032,N_12768,N_11089);
xor UO_1033 (O_1033,N_14187,N_14966);
or UO_1034 (O_1034,N_14557,N_10852);
nand UO_1035 (O_1035,N_13779,N_11193);
and UO_1036 (O_1036,N_13896,N_14111);
or UO_1037 (O_1037,N_13612,N_13416);
nand UO_1038 (O_1038,N_14217,N_10689);
nor UO_1039 (O_1039,N_14432,N_13625);
and UO_1040 (O_1040,N_14178,N_14425);
xnor UO_1041 (O_1041,N_14601,N_14883);
or UO_1042 (O_1042,N_14643,N_11491);
and UO_1043 (O_1043,N_11922,N_13668);
nand UO_1044 (O_1044,N_10160,N_14898);
or UO_1045 (O_1045,N_14451,N_14125);
nor UO_1046 (O_1046,N_10580,N_14162);
and UO_1047 (O_1047,N_11573,N_11225);
and UO_1048 (O_1048,N_13587,N_10186);
or UO_1049 (O_1049,N_11688,N_14146);
nor UO_1050 (O_1050,N_13510,N_11180);
and UO_1051 (O_1051,N_12695,N_12112);
and UO_1052 (O_1052,N_14630,N_12044);
nand UO_1053 (O_1053,N_14795,N_10635);
or UO_1054 (O_1054,N_11626,N_10371);
nand UO_1055 (O_1055,N_10610,N_14747);
nand UO_1056 (O_1056,N_13288,N_13259);
or UO_1057 (O_1057,N_10786,N_14076);
nor UO_1058 (O_1058,N_10875,N_11137);
and UO_1059 (O_1059,N_11372,N_12779);
nand UO_1060 (O_1060,N_13193,N_13965);
nand UO_1061 (O_1061,N_12562,N_11308);
nor UO_1062 (O_1062,N_11041,N_10120);
nor UO_1063 (O_1063,N_11945,N_11465);
nor UO_1064 (O_1064,N_12480,N_10462);
or UO_1065 (O_1065,N_11040,N_13333);
nand UO_1066 (O_1066,N_10010,N_11949);
nor UO_1067 (O_1067,N_11044,N_14847);
nor UO_1068 (O_1068,N_12126,N_14244);
or UO_1069 (O_1069,N_10177,N_10412);
or UO_1070 (O_1070,N_11741,N_11993);
nand UO_1071 (O_1071,N_12157,N_11223);
nor UO_1072 (O_1072,N_11224,N_12653);
nor UO_1073 (O_1073,N_11073,N_10592);
and UO_1074 (O_1074,N_12734,N_14388);
and UO_1075 (O_1075,N_11125,N_14301);
or UO_1076 (O_1076,N_10791,N_13532);
and UO_1077 (O_1077,N_14504,N_14313);
nor UO_1078 (O_1078,N_11816,N_13821);
nor UO_1079 (O_1079,N_13137,N_12742);
and UO_1080 (O_1080,N_12976,N_14823);
or UO_1081 (O_1081,N_10284,N_11297);
nand UO_1082 (O_1082,N_12778,N_11788);
or UO_1083 (O_1083,N_11767,N_13247);
or UO_1084 (O_1084,N_14676,N_14928);
and UO_1085 (O_1085,N_13549,N_14937);
or UO_1086 (O_1086,N_11367,N_11500);
nand UO_1087 (O_1087,N_12248,N_14556);
nand UO_1088 (O_1088,N_12130,N_11525);
or UO_1089 (O_1089,N_14637,N_12150);
xnor UO_1090 (O_1090,N_11456,N_11548);
nand UO_1091 (O_1091,N_10230,N_13652);
nand UO_1092 (O_1092,N_14491,N_10155);
nor UO_1093 (O_1093,N_11962,N_13250);
or UO_1094 (O_1094,N_13566,N_12164);
nor UO_1095 (O_1095,N_11419,N_14679);
nor UO_1096 (O_1096,N_12862,N_12727);
or UO_1097 (O_1097,N_12784,N_10871);
nand UO_1098 (O_1098,N_14404,N_10467);
nor UO_1099 (O_1099,N_10192,N_11305);
nor UO_1100 (O_1100,N_14177,N_14573);
nand UO_1101 (O_1101,N_11149,N_14666);
nand UO_1102 (O_1102,N_14925,N_13884);
nor UO_1103 (O_1103,N_13757,N_13874);
nor UO_1104 (O_1104,N_11349,N_10700);
nor UO_1105 (O_1105,N_12702,N_10804);
nor UO_1106 (O_1106,N_13325,N_12677);
nand UO_1107 (O_1107,N_11270,N_13487);
or UO_1108 (O_1108,N_10942,N_12161);
nand UO_1109 (O_1109,N_10310,N_12966);
or UO_1110 (O_1110,N_13656,N_13124);
and UO_1111 (O_1111,N_13976,N_13585);
nand UO_1112 (O_1112,N_13552,N_11253);
and UO_1113 (O_1113,N_11498,N_11667);
and UO_1114 (O_1114,N_11134,N_12628);
and UO_1115 (O_1115,N_10695,N_14508);
nor UO_1116 (O_1116,N_11145,N_14829);
and UO_1117 (O_1117,N_13052,N_12743);
and UO_1118 (O_1118,N_14594,N_13028);
nand UO_1119 (O_1119,N_13959,N_13778);
nor UO_1120 (O_1120,N_10235,N_13143);
and UO_1121 (O_1121,N_11435,N_10894);
nor UO_1122 (O_1122,N_12875,N_13125);
nand UO_1123 (O_1123,N_12958,N_14587);
and UO_1124 (O_1124,N_13951,N_12216);
or UO_1125 (O_1125,N_14486,N_13998);
and UO_1126 (O_1126,N_11163,N_12364);
and UO_1127 (O_1127,N_10254,N_14797);
nor UO_1128 (O_1128,N_12235,N_14145);
nand UO_1129 (O_1129,N_13328,N_12550);
and UO_1130 (O_1130,N_11438,N_11764);
and UO_1131 (O_1131,N_10601,N_10406);
and UO_1132 (O_1132,N_11886,N_14787);
nor UO_1133 (O_1133,N_12523,N_14082);
and UO_1134 (O_1134,N_14986,N_10121);
and UO_1135 (O_1135,N_11680,N_10044);
nor UO_1136 (O_1136,N_12775,N_13003);
xnor UO_1137 (O_1137,N_14858,N_13980);
or UO_1138 (O_1138,N_13139,N_14369);
nand UO_1139 (O_1139,N_10604,N_14368);
nor UO_1140 (O_1140,N_14351,N_11010);
or UO_1141 (O_1141,N_14790,N_13346);
and UO_1142 (O_1142,N_14985,N_13766);
and UO_1143 (O_1143,N_10287,N_11236);
nand UO_1144 (O_1144,N_14873,N_11590);
and UO_1145 (O_1145,N_13163,N_10091);
and UO_1146 (O_1146,N_12277,N_11593);
and UO_1147 (O_1147,N_12148,N_14968);
xor UO_1148 (O_1148,N_12241,N_11944);
or UO_1149 (O_1149,N_14947,N_13004);
or UO_1150 (O_1150,N_11262,N_10518);
nand UO_1151 (O_1151,N_14020,N_11079);
and UO_1152 (O_1152,N_11038,N_14650);
nor UO_1153 (O_1153,N_11271,N_10434);
nand UO_1154 (O_1154,N_14144,N_14638);
and UO_1155 (O_1155,N_10512,N_14894);
xnor UO_1156 (O_1156,N_12466,N_11108);
nand UO_1157 (O_1157,N_12253,N_12624);
or UO_1158 (O_1158,N_12375,N_14161);
nor UO_1159 (O_1159,N_11522,N_11404);
nor UO_1160 (O_1160,N_13593,N_10409);
nor UO_1161 (O_1161,N_11361,N_12452);
nand UO_1162 (O_1162,N_11373,N_14414);
nand UO_1163 (O_1163,N_10715,N_13309);
nor UO_1164 (O_1164,N_12213,N_12398);
and UO_1165 (O_1165,N_14153,N_10720);
or UO_1166 (O_1166,N_14337,N_12456);
nor UO_1167 (O_1167,N_14310,N_14054);
and UO_1168 (O_1168,N_12567,N_11369);
nand UO_1169 (O_1169,N_14720,N_12950);
or UO_1170 (O_1170,N_10335,N_14287);
or UO_1171 (O_1171,N_12113,N_13518);
nor UO_1172 (O_1172,N_11246,N_13075);
nor UO_1173 (O_1173,N_13742,N_12335);
or UO_1174 (O_1174,N_10275,N_10464);
or UO_1175 (O_1175,N_12085,N_13531);
or UO_1176 (O_1176,N_14138,N_10537);
or UO_1177 (O_1177,N_12535,N_11484);
nor UO_1178 (O_1178,N_10815,N_13404);
and UO_1179 (O_1179,N_10736,N_11293);
and UO_1180 (O_1180,N_11233,N_13455);
or UO_1181 (O_1181,N_13999,N_12772);
nor UO_1182 (O_1182,N_14277,N_11848);
xnor UO_1183 (O_1183,N_13367,N_11329);
and UO_1184 (O_1184,N_13582,N_12904);
and UO_1185 (O_1185,N_14314,N_13160);
and UO_1186 (O_1186,N_10449,N_13311);
nand UO_1187 (O_1187,N_10102,N_12481);
nand UO_1188 (O_1188,N_10808,N_12268);
and UO_1189 (O_1189,N_11837,N_10790);
and UO_1190 (O_1190,N_13310,N_10336);
or UO_1191 (O_1191,N_10713,N_12951);
nor UO_1192 (O_1192,N_11813,N_14353);
nor UO_1193 (O_1193,N_14241,N_14914);
and UO_1194 (O_1194,N_13443,N_14910);
nand UO_1195 (O_1195,N_11037,N_10332);
nand UO_1196 (O_1196,N_14800,N_14331);
nand UO_1197 (O_1197,N_13110,N_14726);
or UO_1198 (O_1198,N_14775,N_11889);
or UO_1199 (O_1199,N_10576,N_11807);
and UO_1200 (O_1200,N_14616,N_14234);
or UO_1201 (O_1201,N_10753,N_10178);
or UO_1202 (O_1202,N_14546,N_14447);
nor UO_1203 (O_1203,N_10470,N_12191);
nor UO_1204 (O_1204,N_12031,N_13619);
nand UO_1205 (O_1205,N_12492,N_10443);
nand UO_1206 (O_1206,N_12339,N_10586);
and UO_1207 (O_1207,N_13046,N_13468);
or UO_1208 (O_1208,N_14932,N_14685);
xnor UO_1209 (O_1209,N_14492,N_14120);
and UO_1210 (O_1210,N_11020,N_14112);
nor UO_1211 (O_1211,N_10896,N_12069);
nand UO_1212 (O_1212,N_13238,N_11931);
and UO_1213 (O_1213,N_11709,N_14606);
or UO_1214 (O_1214,N_12689,N_13301);
or UO_1215 (O_1215,N_11492,N_10522);
and UO_1216 (O_1216,N_12465,N_10261);
or UO_1217 (O_1217,N_10560,N_12938);
or UO_1218 (O_1218,N_14554,N_11085);
or UO_1219 (O_1219,N_13406,N_11445);
nor UO_1220 (O_1220,N_12617,N_13378);
nand UO_1221 (O_1221,N_11200,N_12597);
and UO_1222 (O_1222,N_14083,N_11717);
or UO_1223 (O_1223,N_10360,N_10876);
and UO_1224 (O_1224,N_12580,N_14592);
nor UO_1225 (O_1225,N_12449,N_14579);
and UO_1226 (O_1226,N_12744,N_13788);
nor UO_1227 (O_1227,N_12730,N_10065);
and UO_1228 (O_1228,N_13129,N_14222);
nor UO_1229 (O_1229,N_11453,N_10161);
and UO_1230 (O_1230,N_10034,N_11457);
nor UO_1231 (O_1231,N_14038,N_12972);
nor UO_1232 (O_1232,N_14479,N_12572);
nand UO_1233 (O_1233,N_14157,N_11427);
nand UO_1234 (O_1234,N_14266,N_10656);
nand UO_1235 (O_1235,N_10831,N_12822);
nor UO_1236 (O_1236,N_13031,N_13186);
xor UO_1237 (O_1237,N_11977,N_13005);
nand UO_1238 (O_1238,N_11541,N_12849);
nand UO_1239 (O_1239,N_11295,N_11421);
and UO_1240 (O_1240,N_12579,N_13022);
nor UO_1241 (O_1241,N_11642,N_12014);
nor UO_1242 (O_1242,N_13253,N_13375);
xnor UO_1243 (O_1243,N_14931,N_12613);
and UO_1244 (O_1244,N_14213,N_11000);
or UO_1245 (O_1245,N_10661,N_11657);
nand UO_1246 (O_1246,N_11510,N_11565);
nand UO_1247 (O_1247,N_14249,N_14920);
or UO_1248 (O_1248,N_11831,N_13754);
or UO_1249 (O_1249,N_11956,N_11032);
or UO_1250 (O_1250,N_14176,N_13796);
nand UO_1251 (O_1251,N_14335,N_14549);
or UO_1252 (O_1252,N_11853,N_11592);
and UO_1253 (O_1253,N_13261,N_14233);
and UO_1254 (O_1254,N_11028,N_13352);
and UO_1255 (O_1255,N_13857,N_11058);
nand UO_1256 (O_1256,N_12806,N_13086);
or UO_1257 (O_1257,N_11519,N_14135);
and UO_1258 (O_1258,N_13042,N_13924);
nand UO_1259 (O_1259,N_12098,N_12399);
or UO_1260 (O_1260,N_14719,N_10104);
nor UO_1261 (O_1261,N_10337,N_13441);
or UO_1262 (O_1262,N_14961,N_14140);
and UO_1263 (O_1263,N_10819,N_14035);
or UO_1264 (O_1264,N_14801,N_14610);
nor UO_1265 (O_1265,N_14007,N_10438);
and UO_1266 (O_1266,N_13464,N_11220);
and UO_1267 (O_1267,N_14652,N_13096);
or UO_1268 (O_1268,N_11370,N_12038);
or UO_1269 (O_1269,N_12923,N_12082);
or UO_1270 (O_1270,N_13968,N_10862);
or UO_1271 (O_1271,N_11570,N_11981);
and UO_1272 (O_1272,N_14690,N_10944);
or UO_1273 (O_1273,N_12507,N_10045);
nor UO_1274 (O_1274,N_13725,N_11534);
nor UO_1275 (O_1275,N_11187,N_13775);
nand UO_1276 (O_1276,N_11065,N_14911);
nor UO_1277 (O_1277,N_13397,N_12414);
nor UO_1278 (O_1278,N_12259,N_10818);
or UO_1279 (O_1279,N_14139,N_13561);
nor UO_1280 (O_1280,N_12771,N_13241);
nor UO_1281 (O_1281,N_13932,N_13314);
nand UO_1282 (O_1282,N_14068,N_11365);
or UO_1283 (O_1283,N_11470,N_14405);
and UO_1284 (O_1284,N_12172,N_13752);
nor UO_1285 (O_1285,N_11917,N_13287);
xnor UO_1286 (O_1286,N_12080,N_11321);
or UO_1287 (O_1287,N_13640,N_12242);
and UO_1288 (O_1288,N_14886,N_13192);
nand UO_1289 (O_1289,N_13258,N_14537);
nand UO_1290 (O_1290,N_14812,N_12563);
nor UO_1291 (O_1291,N_14169,N_11904);
nor UO_1292 (O_1292,N_13856,N_14668);
nor UO_1293 (O_1293,N_12273,N_10630);
and UO_1294 (O_1294,N_14608,N_14326);
or UO_1295 (O_1295,N_14595,N_13844);
or UO_1296 (O_1296,N_14686,N_12791);
and UO_1297 (O_1297,N_14942,N_14912);
or UO_1298 (O_1298,N_13801,N_14203);
and UO_1299 (O_1299,N_10642,N_14565);
and UO_1300 (O_1300,N_14861,N_10887);
nand UO_1301 (O_1301,N_13394,N_11615);
or UO_1302 (O_1302,N_11804,N_11494);
or UO_1303 (O_1303,N_11389,N_12781);
nor UO_1304 (O_1304,N_12376,N_10460);
and UO_1305 (O_1305,N_13800,N_10147);
xor UO_1306 (O_1306,N_14377,N_10281);
nand UO_1307 (O_1307,N_10517,N_12475);
nand UO_1308 (O_1308,N_14253,N_11423);
nand UO_1309 (O_1309,N_13929,N_12931);
or UO_1310 (O_1310,N_14848,N_12304);
nand UO_1311 (O_1311,N_10062,N_11914);
nor UO_1312 (O_1312,N_10726,N_10957);
or UO_1313 (O_1313,N_13440,N_13206);
nand UO_1314 (O_1314,N_11991,N_11983);
nand UO_1315 (O_1315,N_13743,N_10119);
nand UO_1316 (O_1316,N_11989,N_10124);
or UO_1317 (O_1317,N_13522,N_11893);
or UO_1318 (O_1318,N_13219,N_10609);
and UO_1319 (O_1319,N_12446,N_10003);
and UO_1320 (O_1320,N_14317,N_12574);
nand UO_1321 (O_1321,N_10676,N_10138);
nand UO_1322 (O_1322,N_12637,N_14229);
nor UO_1323 (O_1323,N_13100,N_12143);
nand UO_1324 (O_1324,N_11336,N_14378);
nor UO_1325 (O_1325,N_11653,N_13112);
and UO_1326 (O_1326,N_11279,N_11971);
nand UO_1327 (O_1327,N_11371,N_13396);
or UO_1328 (O_1328,N_13867,N_10866);
nor UO_1329 (O_1329,N_13077,N_13002);
xnor UO_1330 (O_1330,N_12322,N_14069);
or UO_1331 (O_1331,N_12036,N_12949);
nor UO_1332 (O_1332,N_12251,N_13447);
and UO_1333 (O_1333,N_12725,N_14339);
and UO_1334 (O_1334,N_14705,N_10925);
or UO_1335 (O_1335,N_10424,N_12584);
nand UO_1336 (O_1336,N_14371,N_12851);
nand UO_1337 (O_1337,N_13967,N_10243);
nand UO_1338 (O_1338,N_12012,N_13899);
nand UO_1339 (O_1339,N_11449,N_13789);
xor UO_1340 (O_1340,N_12717,N_10647);
nor UO_1341 (O_1341,N_14600,N_12707);
or UO_1342 (O_1342,N_14563,N_11237);
nand UO_1343 (O_1343,N_10613,N_10550);
nand UO_1344 (O_1344,N_12891,N_12350);
xor UO_1345 (O_1345,N_14589,N_13987);
and UO_1346 (O_1346,N_14239,N_12221);
nor UO_1347 (O_1347,N_14214,N_12457);
nand UO_1348 (O_1348,N_14744,N_14097);
nand UO_1349 (O_1349,N_12004,N_14115);
nand UO_1350 (O_1350,N_10154,N_13359);
and UO_1351 (O_1351,N_12317,N_11198);
nor UO_1352 (O_1352,N_10844,N_10393);
and UO_1353 (O_1353,N_10040,N_12988);
or UO_1354 (O_1354,N_14481,N_14408);
and UO_1355 (O_1355,N_12551,N_10029);
and UO_1356 (O_1356,N_10461,N_14304);
nor UO_1357 (O_1357,N_12852,N_10571);
nand UO_1358 (O_1358,N_14919,N_12473);
nand UO_1359 (O_1359,N_11715,N_11434);
or UO_1360 (O_1360,N_13820,N_14933);
or UO_1361 (O_1361,N_10232,N_12932);
or UO_1362 (O_1362,N_12308,N_11433);
or UO_1363 (O_1363,N_10504,N_11602);
or UO_1364 (O_1364,N_13971,N_12826);
nand UO_1365 (O_1365,N_14151,N_14260);
and UO_1366 (O_1366,N_13978,N_10217);
and UO_1367 (O_1367,N_14208,N_13188);
nand UO_1368 (O_1368,N_14458,N_13564);
or UO_1369 (O_1369,N_11823,N_11818);
and UO_1370 (O_1370,N_10708,N_10152);
nor UO_1371 (O_1371,N_10242,N_10832);
and UO_1372 (O_1372,N_11368,N_13132);
or UO_1373 (O_1373,N_14694,N_13997);
nand UO_1374 (O_1374,N_11524,N_11847);
and UO_1375 (O_1375,N_13659,N_11810);
or UO_1376 (O_1376,N_10168,N_12878);
or UO_1377 (O_1377,N_13765,N_10493);
or UO_1378 (O_1378,N_13343,N_11504);
or UO_1379 (O_1379,N_12302,N_14184);
or UO_1380 (O_1380,N_14757,N_11004);
and UO_1381 (O_1381,N_10558,N_10869);
or UO_1382 (O_1382,N_13227,N_11203);
nand UO_1383 (O_1383,N_13084,N_10886);
xnor UO_1384 (O_1384,N_11546,N_10305);
nand UO_1385 (O_1385,N_10007,N_13141);
and UO_1386 (O_1386,N_11777,N_12274);
nand UO_1387 (O_1387,N_11892,N_12586);
or UO_1388 (O_1388,N_10158,N_14833);
and UO_1389 (O_1389,N_13832,N_13860);
nand UO_1390 (O_1390,N_14751,N_13149);
or UO_1391 (O_1391,N_13641,N_10323);
and UO_1392 (O_1392,N_10860,N_11523);
and UO_1393 (O_1393,N_14292,N_10417);
and UO_1394 (O_1394,N_14091,N_11496);
nor UO_1395 (O_1395,N_14949,N_12283);
nand UO_1396 (O_1396,N_14821,N_13576);
or UO_1397 (O_1397,N_12013,N_10236);
or UO_1398 (O_1398,N_11616,N_11625);
nand UO_1399 (O_1399,N_11244,N_13507);
and UO_1400 (O_1400,N_13161,N_13026);
and UO_1401 (O_1401,N_11743,N_13407);
nand UO_1402 (O_1402,N_12369,N_10110);
or UO_1403 (O_1403,N_13853,N_11264);
nor UO_1404 (O_1404,N_11544,N_10276);
nor UO_1405 (O_1405,N_11695,N_14312);
and UO_1406 (O_1406,N_13090,N_14570);
or UO_1407 (O_1407,N_14970,N_14741);
and UO_1408 (O_1408,N_14688,N_14197);
or UO_1409 (O_1409,N_13408,N_13989);
nor UO_1410 (O_1410,N_13731,N_13946);
and UO_1411 (O_1411,N_12712,N_14027);
and UO_1412 (O_1412,N_10244,N_12863);
or UO_1413 (O_1413,N_13545,N_10901);
or UO_1414 (O_1414,N_14774,N_11603);
nand UO_1415 (O_1415,N_10639,N_10210);
or UO_1416 (O_1416,N_12238,N_10291);
or UO_1417 (O_1417,N_13393,N_12149);
or UO_1418 (O_1418,N_13981,N_14147);
nand UO_1419 (O_1419,N_12751,N_12921);
nand UO_1420 (O_1420,N_13294,N_12916);
nand UO_1421 (O_1421,N_13171,N_14413);
and UO_1422 (O_1422,N_11350,N_13123);
and UO_1423 (O_1423,N_11974,N_13009);
or UO_1424 (O_1424,N_12287,N_10617);
nand UO_1425 (O_1425,N_12652,N_12151);
nor UO_1426 (O_1426,N_13148,N_13466);
nand UO_1427 (O_1427,N_14945,N_11509);
nor UO_1428 (O_1428,N_14446,N_10625);
nor UO_1429 (O_1429,N_12217,N_13836);
or UO_1430 (O_1430,N_11414,N_10459);
nand UO_1431 (O_1431,N_10669,N_14658);
nor UO_1432 (O_1432,N_12843,N_11568);
or UO_1433 (O_1433,N_12601,N_11072);
nand UO_1434 (O_1434,N_11579,N_12516);
nor UO_1435 (O_1435,N_13539,N_13921);
nor UO_1436 (O_1436,N_13027,N_12484);
and UO_1437 (O_1437,N_10657,N_14976);
nand UO_1438 (O_1438,N_10774,N_13057);
nor UO_1439 (O_1439,N_11916,N_13603);
nor UO_1440 (O_1440,N_12602,N_11953);
and UO_1441 (O_1441,N_10440,N_14357);
or UO_1442 (O_1442,N_10285,N_10882);
nor UO_1443 (O_1443,N_11155,N_10296);
and UO_1444 (O_1444,N_13740,N_12713);
and UO_1445 (O_1445,N_10838,N_10093);
nand UO_1446 (O_1446,N_10107,N_11984);
or UO_1447 (O_1447,N_13769,N_11972);
nor UO_1448 (O_1448,N_11026,N_10668);
nor UO_1449 (O_1449,N_12367,N_14345);
and UO_1450 (O_1450,N_14273,N_13483);
and UO_1451 (O_1451,N_10499,N_13621);
nand UO_1452 (O_1452,N_10820,N_12081);
xnor UO_1453 (O_1453,N_14946,N_11396);
nand UO_1454 (O_1454,N_13758,N_14186);
nor UO_1455 (O_1455,N_14366,N_14980);
and UO_1456 (O_1456,N_11645,N_11098);
nand UO_1457 (O_1457,N_13841,N_14788);
and UO_1458 (O_1458,N_10799,N_12028);
nor UO_1459 (O_1459,N_10267,N_11406);
nor UO_1460 (O_1460,N_13559,N_11589);
nor UO_1461 (O_1461,N_14835,N_12979);
nand UO_1462 (O_1462,N_10072,N_12087);
nand UO_1463 (O_1463,N_12208,N_10597);
nand UO_1464 (O_1464,N_14498,N_10092);
nand UO_1465 (O_1465,N_12402,N_14596);
nand UO_1466 (O_1466,N_14849,N_11476);
nand UO_1467 (O_1467,N_13305,N_10933);
nor UO_1468 (O_1468,N_13799,N_14127);
nor UO_1469 (O_1469,N_11161,N_12343);
and UO_1470 (O_1470,N_10426,N_13888);
nand UO_1471 (O_1471,N_11242,N_11294);
or UO_1472 (O_1472,N_11619,N_12272);
and UO_1473 (O_1473,N_10073,N_12141);
or UO_1474 (O_1474,N_14559,N_13535);
nor UO_1475 (O_1475,N_11851,N_10679);
and UO_1476 (O_1476,N_14811,N_14333);
nand UO_1477 (O_1477,N_11803,N_10058);
nor UO_1478 (O_1478,N_13505,N_13463);
and UO_1479 (O_1479,N_14081,N_14202);
nand UO_1480 (O_1480,N_10826,N_14036);
nand UO_1481 (O_1481,N_14000,N_12129);
nand UO_1482 (O_1482,N_12281,N_14530);
nor UO_1483 (O_1483,N_14660,N_11326);
and UO_1484 (O_1484,N_14355,N_13521);
and UO_1485 (O_1485,N_14055,N_11951);
or UO_1486 (O_1486,N_11306,N_14906);
nand UO_1487 (O_1487,N_13390,N_11621);
nand UO_1488 (O_1488,N_14975,N_11793);
and UO_1489 (O_1489,N_12379,N_13903);
or UO_1490 (O_1490,N_12575,N_13203);
nor UO_1491 (O_1491,N_12583,N_14056);
or UO_1492 (O_1492,N_11925,N_14828);
or UO_1493 (O_1493,N_11629,N_14130);
nor UO_1494 (O_1494,N_11786,N_13446);
xnor UO_1495 (O_1495,N_10026,N_13654);
nor UO_1496 (O_1496,N_14291,N_12513);
nor UO_1497 (O_1497,N_13917,N_14944);
or UO_1498 (O_1498,N_13243,N_12560);
nor UO_1499 (O_1499,N_14365,N_10255);
and UO_1500 (O_1500,N_10856,N_12049);
xnor UO_1501 (O_1501,N_12893,N_14725);
nor UO_1502 (O_1502,N_14991,N_11114);
or UO_1503 (O_1503,N_11985,N_10321);
nor UO_1504 (O_1504,N_12156,N_12873);
or UO_1505 (O_1505,N_12962,N_14101);
nor UO_1506 (O_1506,N_10327,N_10041);
nor UO_1507 (O_1507,N_12368,N_14624);
or UO_1508 (O_1508,N_14814,N_12897);
nand UO_1509 (O_1509,N_13427,N_13906);
and UO_1510 (O_1510,N_10362,N_11446);
or UO_1511 (O_1511,N_14155,N_10588);
and UO_1512 (O_1512,N_11148,N_13963);
or UO_1513 (O_1513,N_11266,N_13172);
nor UO_1514 (O_1514,N_13120,N_10484);
or UO_1515 (O_1515,N_10312,N_11934);
nor UO_1516 (O_1516,N_12503,N_13230);
nand UO_1517 (O_1517,N_13755,N_10744);
nand UO_1518 (O_1518,N_14443,N_10137);
or UO_1519 (O_1519,N_14964,N_11686);
nor UO_1520 (O_1520,N_10830,N_10023);
nor UO_1521 (O_1521,N_11407,N_11480);
nand UO_1522 (O_1522,N_13380,N_12309);
nor UO_1523 (O_1523,N_14855,N_12181);
and UO_1524 (O_1524,N_13979,N_10612);
nand UO_1525 (O_1525,N_13209,N_14298);
and UO_1526 (O_1526,N_12520,N_12180);
nor UO_1527 (O_1527,N_12556,N_10688);
nand UO_1528 (O_1528,N_12497,N_11122);
nand UO_1529 (O_1529,N_14662,N_10086);
xnor UO_1530 (O_1530,N_12426,N_14199);
nand UO_1531 (O_1531,N_11070,N_10407);
nor UO_1532 (O_1532,N_12620,N_10979);
or UO_1533 (O_1533,N_11650,N_14028);
and UO_1534 (O_1534,N_11182,N_12239);
nand UO_1535 (O_1535,N_12389,N_11605);
and UO_1536 (O_1536,N_11281,N_11719);
nand UO_1537 (O_1537,N_13272,N_11451);
nand UO_1538 (O_1538,N_10948,N_12459);
nor UO_1539 (O_1539,N_11762,N_14764);
xor UO_1540 (O_1540,N_14648,N_12260);
or UO_1541 (O_1541,N_11292,N_14174);
and UO_1542 (O_1542,N_12490,N_11303);
or UO_1543 (O_1543,N_14852,N_14818);
nand UO_1544 (O_1544,N_13646,N_10166);
nor UO_1545 (O_1545,N_14172,N_11859);
nor UO_1546 (O_1546,N_11302,N_11290);
nand UO_1547 (O_1547,N_10433,N_13260);
nor UO_1548 (O_1548,N_12146,N_12313);
nor UO_1549 (O_1549,N_13038,N_10008);
nand UO_1550 (O_1550,N_11866,N_14207);
and UO_1551 (O_1551,N_11420,N_14086);
nand UO_1552 (O_1552,N_11390,N_14449);
and UO_1553 (O_1553,N_14511,N_10170);
or UO_1554 (O_1554,N_14440,N_13372);
or UO_1555 (O_1555,N_10373,N_14225);
or UO_1556 (O_1556,N_12374,N_12271);
nor UO_1557 (O_1557,N_11243,N_13205);
nor UO_1558 (O_1558,N_10857,N_12647);
and UO_1559 (O_1559,N_10519,N_13520);
and UO_1560 (O_1560,N_10582,N_13011);
nand UO_1561 (O_1561,N_14031,N_13542);
and UO_1562 (O_1562,N_14359,N_12312);
and UO_1563 (O_1563,N_12219,N_10059);
nand UO_1564 (O_1564,N_12171,N_12977);
nor UO_1565 (O_1565,N_10047,N_13732);
nand UO_1566 (O_1566,N_13248,N_12957);
nand UO_1567 (O_1567,N_11769,N_11941);
and UO_1568 (O_1568,N_12847,N_13403);
or UO_1569 (O_1569,N_14087,N_11966);
nand UO_1570 (O_1570,N_14302,N_10723);
nor UO_1571 (O_1571,N_12034,N_13714);
nor UO_1572 (O_1572,N_10202,N_13964);
and UO_1573 (O_1573,N_12001,N_10032);
nand UO_1574 (O_1574,N_11027,N_11175);
nor UO_1575 (O_1575,N_14092,N_10987);
nor UO_1576 (O_1576,N_11617,N_14057);
or UO_1577 (O_1577,N_14049,N_14209);
nand UO_1578 (O_1578,N_13728,N_10916);
nand UO_1579 (O_1579,N_12757,N_14320);
nor UO_1580 (O_1580,N_10973,N_12445);
and UO_1581 (O_1581,N_12183,N_10348);
and UO_1582 (O_1582,N_11828,N_14142);
nand UO_1583 (O_1583,N_14072,N_12448);
or UO_1584 (O_1584,N_10001,N_10309);
nand UO_1585 (O_1585,N_13307,N_13240);
and UO_1586 (O_1586,N_14488,N_14376);
nand UO_1587 (O_1587,N_13155,N_13956);
or UO_1588 (O_1588,N_10590,N_14809);
nor UO_1589 (O_1589,N_13586,N_14519);
and UO_1590 (O_1590,N_10816,N_12360);
nand UO_1591 (O_1591,N_13712,N_14235);
or UO_1592 (O_1592,N_11362,N_14555);
nand UO_1593 (O_1593,N_13970,N_13341);
or UO_1594 (O_1594,N_12311,N_12910);
and UO_1595 (O_1595,N_12167,N_13166);
and UO_1596 (O_1596,N_11780,N_14727);
or UO_1597 (O_1597,N_14940,N_10931);
nor UO_1598 (O_1598,N_10398,N_13292);
nor UO_1599 (O_1599,N_11703,N_13334);
or UO_1600 (O_1600,N_14954,N_11907);
nor UO_1601 (O_1601,N_12678,N_11286);
nand UO_1602 (O_1602,N_14231,N_11063);
nor UO_1603 (O_1603,N_12011,N_11017);
and UO_1604 (O_1604,N_10767,N_14541);
nand UO_1605 (O_1605,N_11102,N_12140);
nand UO_1606 (O_1606,N_14128,N_11995);
nand UO_1607 (O_1607,N_10033,N_13492);
nor UO_1608 (O_1608,N_12963,N_11499);
nor UO_1609 (O_1609,N_10225,N_14553);
nor UO_1610 (O_1610,N_11455,N_10129);
nand UO_1611 (O_1611,N_13941,N_12021);
xor UO_1612 (O_1612,N_10991,N_14048);
nor UO_1613 (O_1613,N_11539,N_10893);
nor UO_1614 (O_1614,N_13097,N_14951);
nor UO_1615 (O_1615,N_11255,N_11335);
nor UO_1616 (O_1616,N_13223,N_12300);
nand UO_1617 (O_1617,N_11980,N_11128);
or UO_1618 (O_1618,N_11649,N_14282);
nand UO_1619 (O_1619,N_14654,N_10189);
and UO_1620 (O_1620,N_10355,N_14965);
nand UO_1621 (O_1621,N_10986,N_14219);
and UO_1622 (O_1622,N_12409,N_10952);
and UO_1623 (O_1623,N_12499,N_14581);
nand UO_1624 (O_1624,N_11094,N_12419);
or UO_1625 (O_1625,N_14529,N_14276);
and UO_1626 (O_1626,N_14259,N_14009);
nand UO_1627 (O_1627,N_12621,N_13748);
and UO_1628 (O_1628,N_13014,N_14584);
and UO_1629 (O_1629,N_10777,N_14979);
or UO_1630 (O_1630,N_10553,N_14561);
nor UO_1631 (O_1631,N_14761,N_12829);
and UO_1632 (O_1632,N_14171,N_14121);
or UO_1633 (O_1633,N_11696,N_13590);
or UO_1634 (O_1634,N_10095,N_11656);
or UO_1635 (O_1635,N_14888,N_14543);
nor UO_1636 (O_1636,N_12889,N_12983);
nand UO_1637 (O_1637,N_10144,N_13513);
nand UO_1638 (O_1638,N_12002,N_11022);
xor UO_1639 (O_1639,N_12076,N_12783);
or UO_1640 (O_1640,N_14989,N_14406);
or UO_1641 (O_1641,N_11042,N_11939);
and UO_1642 (O_1642,N_14014,N_12472);
or UO_1643 (O_1643,N_13643,N_10269);
or UO_1644 (O_1644,N_10643,N_12204);
nor UO_1645 (O_1645,N_10150,N_14678);
xor UO_1646 (O_1646,N_13577,N_11683);
nor UO_1647 (O_1647,N_12813,N_12097);
nor UO_1648 (O_1648,N_10268,N_11355);
nand UO_1649 (O_1649,N_14340,N_12917);
nor UO_1650 (O_1650,N_12741,N_13673);
nor UO_1651 (O_1651,N_11672,N_12868);
nand UO_1652 (O_1652,N_12699,N_10299);
and UO_1653 (O_1653,N_13448,N_13190);
or UO_1654 (O_1654,N_13035,N_13894);
or UO_1655 (O_1655,N_14075,N_12468);
nand UO_1656 (O_1656,N_11256,N_11770);
or UO_1657 (O_1657,N_10213,N_10035);
nand UO_1658 (O_1658,N_11340,N_11812);
xnor UO_1659 (O_1659,N_12077,N_14477);
and UO_1660 (O_1660,N_10611,N_13845);
nor UO_1661 (O_1661,N_13843,N_10222);
or UO_1662 (O_1662,N_14704,N_13814);
and UO_1663 (O_1663,N_11392,N_11153);
or UO_1664 (O_1664,N_14962,N_12776);
or UO_1665 (O_1665,N_13519,N_13140);
and UO_1666 (O_1666,N_13713,N_12830);
xor UO_1667 (O_1667,N_12487,N_11533);
or UO_1668 (O_1668,N_14325,N_11174);
nand UO_1669 (O_1669,N_14475,N_13387);
nand UO_1670 (O_1670,N_11118,N_10967);
nor UO_1671 (O_1671,N_14129,N_14810);
nor UO_1672 (O_1672,N_11508,N_14838);
nand UO_1673 (O_1673,N_14293,N_14872);
and UO_1674 (O_1674,N_10418,N_14409);
nor UO_1675 (O_1675,N_13040,N_11317);
or UO_1676 (O_1676,N_12485,N_12222);
and UO_1677 (O_1677,N_14211,N_13695);
nand UO_1678 (O_1678,N_12328,N_14372);
or UO_1679 (O_1679,N_10694,N_10250);
nor UO_1680 (O_1680,N_11345,N_14907);
nand UO_1681 (O_1681,N_12396,N_14684);
xor UO_1682 (O_1682,N_12676,N_13105);
nor UO_1683 (O_1683,N_11511,N_11868);
or UO_1684 (O_1684,N_12872,N_13278);
nand UO_1685 (O_1685,N_10828,N_12524);
or UO_1686 (O_1686,N_14228,N_11607);
nor UO_1687 (O_1687,N_11176,N_11207);
and UO_1688 (O_1688,N_14180,N_14396);
and UO_1689 (O_1689,N_10637,N_14510);
nor UO_1690 (O_1690,N_14874,N_10274);
nor UO_1691 (O_1691,N_10277,N_10760);
or UO_1692 (O_1692,N_13538,N_14926);
or UO_1693 (O_1693,N_12752,N_12533);
nand UO_1694 (O_1694,N_14939,N_12633);
nor UO_1695 (O_1695,N_14591,N_12939);
nor UO_1696 (O_1696,N_13262,N_11515);
or UO_1697 (O_1697,N_12356,N_11318);
nand UO_1698 (O_1698,N_12888,N_13927);
or UO_1699 (O_1699,N_10331,N_13113);
or UO_1700 (O_1700,N_13151,N_10009);
nor UO_1701 (O_1701,N_14154,N_14230);
and UO_1702 (O_1702,N_13283,N_13433);
nor UO_1703 (O_1703,N_10677,N_12907);
or UO_1704 (O_1704,N_11899,N_14930);
or UO_1705 (O_1705,N_10914,N_14840);
nand UO_1706 (O_1706,N_13300,N_10195);
and UO_1707 (O_1707,N_12420,N_12358);
nor UO_1708 (O_1708,N_14832,N_12864);
or UO_1709 (O_1709,N_13866,N_10219);
nand UO_1710 (O_1710,N_11104,N_10245);
nor UO_1711 (O_1711,N_13472,N_11673);
xor UO_1712 (O_1712,N_12763,N_10346);
nor UO_1713 (O_1713,N_14160,N_13362);
nand UO_1714 (O_1714,N_11655,N_14080);
nor UO_1715 (O_1715,N_13025,N_13960);
xor UO_1716 (O_1716,N_11309,N_10899);
or UO_1717 (O_1717,N_11247,N_13667);
and UO_1718 (O_1718,N_13551,N_11046);
or UO_1719 (O_1719,N_12476,N_11751);
xnor UO_1720 (O_1720,N_13239,N_14542);
and UO_1721 (O_1721,N_10729,N_13589);
xnor UO_1722 (O_1722,N_14401,N_13020);
nand UO_1723 (O_1723,N_13331,N_12486);
or UO_1724 (O_1724,N_14882,N_12833);
and UO_1725 (O_1725,N_10881,N_13013);
nand UO_1726 (O_1726,N_10716,N_12381);
nand UO_1727 (O_1727,N_10027,N_13365);
nand UO_1728 (O_1728,N_14696,N_11385);
and UO_1729 (O_1729,N_14817,N_11043);
nand UO_1730 (O_1730,N_13665,N_10396);
nand UO_1731 (O_1731,N_12548,N_14550);
and UO_1732 (O_1732,N_10962,N_12458);
nor UO_1733 (O_1733,N_12648,N_14820);
nor UO_1734 (O_1734,N_14509,N_13066);
or UO_1735 (O_1735,N_14540,N_12194);
nor UO_1736 (O_1736,N_10920,N_11060);
nand UO_1737 (O_1737,N_10905,N_13704);
nand UO_1738 (O_1738,N_12353,N_11337);
nand UO_1739 (O_1739,N_14957,N_11342);
nand UO_1740 (O_1740,N_11178,N_13344);
and UO_1741 (O_1741,N_14967,N_10629);
or UO_1742 (O_1742,N_12536,N_12760);
or UO_1743 (O_1743,N_10999,N_14841);
nand UO_1744 (O_1744,N_12382,N_12740);
or UO_1745 (O_1745,N_10439,N_12785);
or UO_1746 (O_1746,N_11790,N_10858);
and UO_1747 (O_1747,N_13082,N_13506);
nor UO_1748 (O_1748,N_12811,N_11138);
nor UO_1749 (O_1749,N_10849,N_11857);
or UO_1750 (O_1750,N_12196,N_14879);
or UO_1751 (O_1751,N_12025,N_13633);
xnor UO_1752 (O_1752,N_14416,N_13870);
nand UO_1753 (O_1753,N_10742,N_10185);
and UO_1754 (O_1754,N_12073,N_11181);
nand UO_1755 (O_1755,N_14434,N_13370);
and UO_1756 (O_1756,N_12195,N_14826);
and UO_1757 (O_1757,N_10171,N_14655);
and UO_1758 (O_1758,N_14297,N_10579);
and UO_1759 (O_1759,N_11490,N_13189);
nand UO_1760 (O_1760,N_11197,N_11658);
nand UO_1761 (O_1761,N_10686,N_14100);
nand UO_1762 (O_1762,N_13610,N_10196);
xor UO_1763 (O_1763,N_11685,N_10208);
nand UO_1764 (O_1764,N_13707,N_12683);
xnor UO_1765 (O_1765,N_13534,N_14407);
and UO_1766 (O_1766,N_12159,N_11545);
and UO_1767 (O_1767,N_11412,N_14280);
and UO_1768 (O_1768,N_11150,N_14163);
or UO_1769 (O_1769,N_13214,N_10229);
nor UO_1770 (O_1770,N_14712,N_12500);
nand UO_1771 (O_1771,N_12522,N_12318);
nand UO_1772 (O_1772,N_12264,N_10575);
and UO_1773 (O_1773,N_11742,N_13935);
or UO_1774 (O_1774,N_13550,N_11191);
nand UO_1775 (O_1775,N_11186,N_11867);
nor UO_1776 (O_1776,N_14960,N_10103);
and UO_1777 (O_1777,N_14825,N_11259);
xor UO_1778 (O_1778,N_10263,N_13689);
nand UO_1779 (O_1779,N_10444,N_12594);
nand UO_1780 (O_1780,N_11119,N_12874);
and UO_1781 (O_1781,N_11663,N_13176);
nor UO_1782 (O_1782,N_11623,N_11425);
or UO_1783 (O_1783,N_12471,N_11173);
nand UO_1784 (O_1784,N_13940,N_13974);
or UO_1785 (O_1785,N_13313,N_12853);
or UO_1786 (O_1786,N_12115,N_13216);
or UO_1787 (O_1787,N_12800,N_11136);
nor UO_1788 (O_1788,N_10080,N_11386);
and UO_1789 (O_1789,N_11205,N_11674);
nor UO_1790 (O_1790,N_13234,N_13412);
xnor UO_1791 (O_1791,N_10959,N_14256);
nand UO_1792 (O_1792,N_11881,N_12738);
nand UO_1793 (O_1793,N_12329,N_11879);
nor UO_1794 (O_1794,N_11976,N_12450);
and UO_1795 (O_1795,N_13584,N_13824);
and UO_1796 (O_1796,N_12762,N_10159);
nand UO_1797 (O_1797,N_10699,N_11334);
nand UO_1798 (O_1798,N_11299,N_13588);
and UO_1799 (O_1799,N_11975,N_12798);
and UO_1800 (O_1800,N_12416,N_12425);
or UO_1801 (O_1801,N_14681,N_12925);
and UO_1802 (O_1802,N_11547,N_13751);
and UO_1803 (O_1803,N_11208,N_13524);
and UO_1804 (O_1804,N_10090,N_13526);
and UO_1805 (O_1805,N_13196,N_11409);
or UO_1806 (O_1806,N_12646,N_12232);
or UO_1807 (O_1807,N_12824,N_11755);
or UO_1808 (O_1808,N_12066,N_13892);
nand UO_1809 (O_1809,N_13763,N_14948);
nand UO_1810 (O_1810,N_11240,N_10797);
nor UO_1811 (O_1811,N_11842,N_12841);
nor UO_1812 (O_1812,N_12105,N_12261);
nand UO_1813 (O_1813,N_12592,N_10514);
nand UO_1814 (O_1814,N_13368,N_14032);
or UO_1815 (O_1815,N_14717,N_14803);
and UO_1816 (O_1816,N_10325,N_14843);
nand UO_1817 (O_1817,N_12635,N_13502);
nand UO_1818 (O_1818,N_14901,N_13477);
and UO_1819 (O_1819,N_13018,N_11024);
or UO_1820 (O_1820,N_10696,N_10125);
nand UO_1821 (O_1821,N_13353,N_13128);
and UO_1822 (O_1822,N_14728,N_11194);
or UO_1823 (O_1823,N_10770,N_14418);
nand UO_1824 (O_1824,N_10891,N_12899);
or UO_1825 (O_1825,N_10114,N_11801);
or UO_1826 (O_1826,N_11708,N_10717);
and UO_1827 (O_1827,N_12913,N_10795);
and UO_1828 (O_1828,N_13939,N_13993);
or UO_1829 (O_1829,N_14026,N_12838);
nand UO_1830 (O_1830,N_10653,N_13430);
nor UO_1831 (O_1831,N_11618,N_10358);
or UO_1832 (O_1832,N_13579,N_12960);
and UO_1833 (O_1833,N_14489,N_11609);
or UO_1834 (O_1834,N_13458,N_11395);
and UO_1835 (O_1835,N_14521,N_10101);
xor UO_1836 (O_1836,N_14476,N_11113);
or UO_1837 (O_1837,N_13481,N_14669);
nand UO_1838 (O_1838,N_11422,N_10941);
and UO_1839 (O_1839,N_11123,N_14341);
nor UO_1840 (O_1840,N_14023,N_10295);
nor UO_1841 (O_1841,N_13275,N_11679);
or UO_1842 (O_1842,N_11289,N_13650);
nor UO_1843 (O_1843,N_12051,N_11003);
or UO_1844 (O_1844,N_12024,N_12543);
xnor UO_1845 (O_1845,N_12599,N_11869);
or UO_1846 (O_1846,N_13849,N_13905);
nand UO_1847 (O_1847,N_12720,N_13457);
xnor UO_1848 (O_1848,N_14750,N_12469);
nor UO_1849 (O_1849,N_13364,N_13578);
nor UO_1850 (O_1850,N_13326,N_10455);
nand UO_1851 (O_1851,N_11747,N_10526);
nor UO_1852 (O_1852,N_11994,N_14426);
nand UO_1853 (O_1853,N_11955,N_11352);
nand UO_1854 (O_1854,N_11883,N_14467);
nor UO_1855 (O_1855,N_11322,N_10884);
or UO_1856 (O_1856,N_13162,N_12334);
or UO_1857 (O_1857,N_14200,N_10453);
nor UO_1858 (O_1858,N_11580,N_13371);
nor UO_1859 (O_1859,N_14807,N_10606);
or UO_1860 (O_1860,N_11946,N_13774);
nand UO_1861 (O_1861,N_14739,N_13910);
and UO_1862 (O_1862,N_11675,N_11162);
nand UO_1863 (O_1863,N_10068,N_10655);
or UO_1864 (O_1864,N_14934,N_14599);
and UO_1865 (O_1865,N_14034,N_10253);
and UO_1866 (O_1866,N_10636,N_13237);
and UO_1867 (O_1867,N_12436,N_13827);
or UO_1868 (O_1868,N_13991,N_11639);
and UO_1869 (O_1869,N_12807,N_14232);
and UO_1870 (O_1870,N_13805,N_10562);
or UO_1871 (O_1871,N_13642,N_14246);
nand UO_1872 (O_1872,N_13183,N_11151);
nor UO_1873 (O_1873,N_12859,N_11472);
nand UO_1874 (O_1874,N_10313,N_14673);
and UO_1875 (O_1875,N_13573,N_12207);
nor UO_1876 (O_1876,N_14604,N_13508);
or UO_1877 (O_1877,N_10141,N_12407);
and UO_1878 (O_1878,N_10638,N_12357);
and UO_1879 (O_1879,N_12618,N_10352);
or UO_1880 (O_1880,N_13444,N_13062);
nand UO_1881 (O_1881,N_13494,N_13399);
or UO_1882 (O_1882,N_13217,N_14456);
nand UO_1883 (O_1883,N_10835,N_10730);
or UO_1884 (O_1884,N_13708,N_14889);
or UO_1885 (O_1885,N_12870,N_13983);
and UO_1886 (O_1886,N_12866,N_14691);
and UO_1887 (O_1887,N_14008,N_14862);
nor UO_1888 (O_1888,N_12061,N_13012);
nor UO_1889 (O_1889,N_11319,N_12644);
nor UO_1890 (O_1890,N_12970,N_14748);
nor UO_1891 (O_1891,N_10982,N_10600);
nand UO_1892 (O_1892,N_14756,N_14598);
nor UO_1893 (O_1893,N_14019,N_12716);
and UO_1894 (O_1894,N_10031,N_14635);
nor UO_1895 (O_1895,N_10911,N_12748);
and UO_1896 (O_1896,N_13428,N_11353);
or UO_1897 (O_1897,N_13064,N_13296);
and UO_1898 (O_1898,N_13569,N_10873);
xnor UO_1899 (O_1899,N_12179,N_13527);
nor UO_1900 (O_1900,N_13923,N_13895);
and UO_1901 (O_1901,N_13099,N_13780);
nor UO_1902 (O_1902,N_11723,N_11797);
nand UO_1903 (O_1903,N_11483,N_13795);
or UO_1904 (O_1904,N_13442,N_14271);
nor UO_1905 (O_1905,N_13101,N_11439);
or UO_1906 (O_1906,N_10678,N_14941);
or UO_1907 (O_1907,N_12802,N_14990);
or UO_1908 (O_1908,N_13181,N_14323);
nor UO_1909 (O_1909,N_12095,N_14663);
nor UO_1910 (O_1910,N_11965,N_11776);
nand UO_1911 (O_1911,N_14102,N_10215);
nand UO_1912 (O_1912,N_12046,N_11738);
nand UO_1913 (O_1913,N_12390,N_10539);
nor UO_1914 (O_1914,N_10385,N_13474);
and UO_1915 (O_1915,N_10165,N_13762);
and UO_1916 (O_1916,N_10548,N_10294);
or UO_1917 (O_1917,N_12696,N_14373);
and UO_1918 (O_1918,N_13699,N_11574);
or UO_1919 (O_1919,N_12215,N_12429);
nor UO_1920 (O_1920,N_14290,N_14702);
nor UO_1921 (O_1921,N_10788,N_13257);
or UO_1922 (O_1922,N_14307,N_10151);
nor UO_1923 (O_1923,N_14025,N_11613);
nor UO_1924 (O_1924,N_12166,N_10954);
and UO_1925 (O_1925,N_11697,N_12435);
or UO_1926 (O_1926,N_10201,N_12611);
nor UO_1927 (O_1927,N_12777,N_10238);
or UO_1928 (O_1928,N_10182,N_11358);
nor UO_1929 (O_1929,N_11640,N_12954);
xnor UO_1930 (O_1930,N_12078,N_12982);
or UO_1931 (O_1931,N_14715,N_12192);
and UO_1932 (O_1932,N_13347,N_13114);
or UO_1933 (O_1933,N_12114,N_14837);
nor UO_1934 (O_1934,N_14799,N_13873);
nand UO_1935 (O_1935,N_14420,N_12810);
and UO_1936 (O_1936,N_14367,N_13179);
nor UO_1937 (O_1937,N_10247,N_10050);
and UO_1938 (O_1938,N_13571,N_12542);
and UO_1939 (O_1939,N_14729,N_10006);
nand UO_1940 (O_1940,N_11226,N_11690);
xnor UO_1941 (O_1941,N_11431,N_14544);
and UO_1942 (O_1942,N_12427,N_10311);
xor UO_1943 (O_1943,N_11978,N_14286);
and UO_1944 (O_1944,N_13717,N_10015);
nand UO_1945 (O_1945,N_12493,N_12746);
or UO_1946 (O_1946,N_11169,N_13089);
nand UO_1947 (O_1947,N_12630,N_11572);
nor UO_1948 (O_1948,N_10018,N_10897);
nand UO_1949 (O_1949,N_10038,N_10594);
or UO_1950 (O_1950,N_11351,N_11921);
and UO_1951 (O_1951,N_12009,N_13840);
nor UO_1952 (O_1952,N_11862,N_12598);
nand UO_1953 (O_1953,N_14379,N_10183);
or UO_1954 (O_1954,N_12769,N_14548);
nor UO_1955 (O_1955,N_11958,N_11463);
and UO_1956 (O_1956,N_13232,N_10482);
or UO_1957 (O_1957,N_14272,N_11018);
xor UO_1958 (O_1958,N_14516,N_14866);
nor UO_1959 (O_1959,N_10452,N_14723);
and UO_1960 (O_1960,N_10153,N_13847);
or UO_1961 (O_1961,N_12132,N_10115);
or UO_1962 (O_1962,N_12134,N_11219);
nand UO_1963 (O_1963,N_13422,N_12799);
and UO_1964 (O_1964,N_11047,N_13684);
nor UO_1965 (O_1965,N_14621,N_12244);
and UO_1966 (O_1966,N_12366,N_11782);
or UO_1967 (O_1967,N_10659,N_13563);
or UO_1968 (O_1968,N_14528,N_10682);
or UO_1969 (O_1969,N_11809,N_13144);
nand UO_1970 (O_1970,N_14393,N_14263);
nor UO_1971 (O_1971,N_11600,N_10098);
and UO_1972 (O_1972,N_10206,N_11849);
nand UO_1973 (O_1973,N_10572,N_13772);
and UO_1974 (O_1974,N_13118,N_11227);
nand UO_1975 (O_1975,N_14270,N_11543);
and UO_1976 (O_1976,N_14983,N_13733);
and UO_1977 (O_1977,N_12971,N_10547);
and UO_1978 (O_1978,N_13254,N_12257);
nand UO_1979 (O_1979,N_14569,N_10765);
or UO_1980 (O_1980,N_12694,N_10892);
nand UO_1981 (O_1981,N_12106,N_13977);
or UO_1982 (O_1982,N_12512,N_12307);
and UO_1983 (O_1983,N_14044,N_11092);
nand UO_1984 (O_1984,N_10650,N_11520);
and UO_1985 (O_1985,N_10515,N_12606);
or UO_1986 (O_1986,N_12100,N_10194);
nor UO_1987 (O_1987,N_13142,N_10812);
or UO_1988 (O_1988,N_12591,N_14623);
nand UO_1989 (O_1989,N_12225,N_14483);
nand UO_1990 (O_1990,N_10241,N_11157);
or UO_1991 (O_1991,N_10079,N_11106);
or UO_1992 (O_1992,N_10126,N_11291);
and UO_1993 (O_1993,N_12168,N_14984);
and UO_1994 (O_1994,N_11891,N_12812);
and UO_1995 (O_1995,N_13703,N_10089);
xnor UO_1996 (O_1996,N_11283,N_11729);
or UO_1997 (O_1997,N_14463,N_10934);
nand UO_1998 (O_1998,N_10477,N_11720);
or UO_1999 (O_1999,N_14771,N_14114);
endmodule