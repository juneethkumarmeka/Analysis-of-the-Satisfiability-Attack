module basic_500_3000_500_15_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_471,In_496);
nor U1 (N_1,In_61,In_402);
nor U2 (N_2,In_164,In_484);
nor U3 (N_3,In_111,In_428);
nand U4 (N_4,In_250,In_150);
nand U5 (N_5,In_218,In_482);
and U6 (N_6,In_406,In_327);
or U7 (N_7,In_110,In_84);
nor U8 (N_8,In_200,In_384);
nor U9 (N_9,In_261,In_314);
nor U10 (N_10,In_331,In_215);
nor U11 (N_11,In_232,In_497);
nor U12 (N_12,In_297,In_400);
or U13 (N_13,In_442,In_429);
xnor U14 (N_14,In_452,In_199);
nor U15 (N_15,In_301,In_25);
and U16 (N_16,In_489,In_268);
xnor U17 (N_17,In_125,In_324);
nand U18 (N_18,In_222,In_330);
nor U19 (N_19,In_131,In_269);
and U20 (N_20,In_485,In_385);
or U21 (N_21,In_210,In_226);
or U22 (N_22,In_239,In_202);
and U23 (N_23,In_145,In_85);
or U24 (N_24,In_291,In_329);
nand U25 (N_25,In_244,In_168);
nand U26 (N_26,In_336,In_368);
or U27 (N_27,In_24,In_286);
nand U28 (N_28,In_183,In_119);
and U29 (N_29,In_68,In_127);
or U30 (N_30,In_77,In_151);
or U31 (N_31,In_326,In_63);
and U32 (N_32,In_399,In_405);
nand U33 (N_33,In_86,In_108);
xor U34 (N_34,In_389,In_133);
nor U35 (N_35,In_416,In_432);
nor U36 (N_36,In_352,In_375);
and U37 (N_37,In_453,In_97);
and U38 (N_38,In_190,In_309);
nor U39 (N_39,In_284,In_444);
and U40 (N_40,In_454,In_191);
nand U41 (N_41,In_19,In_498);
xor U42 (N_42,In_251,In_342);
xnor U43 (N_43,In_130,In_383);
and U44 (N_44,In_12,In_414);
or U45 (N_45,In_185,In_128);
and U46 (N_46,In_358,In_413);
or U47 (N_47,In_209,In_134);
or U48 (N_48,In_212,In_236);
nand U49 (N_49,In_466,In_14);
nor U50 (N_50,In_163,In_319);
nand U51 (N_51,In_347,In_462);
and U52 (N_52,In_0,In_499);
or U53 (N_53,In_182,In_493);
and U54 (N_54,In_231,In_121);
nor U55 (N_55,In_270,In_247);
nor U56 (N_56,In_157,In_6);
and U57 (N_57,In_170,In_470);
or U58 (N_58,In_95,In_274);
xor U59 (N_59,In_227,In_278);
or U60 (N_60,In_320,In_92);
or U61 (N_61,In_66,In_17);
or U62 (N_62,In_192,In_287);
or U63 (N_63,In_217,In_390);
nand U64 (N_64,In_197,In_420);
and U65 (N_65,In_44,In_457);
nand U66 (N_66,In_27,In_280);
or U67 (N_67,In_488,In_79);
nand U68 (N_68,In_43,In_203);
nor U69 (N_69,In_441,In_245);
or U70 (N_70,In_15,In_120);
xnor U71 (N_71,In_80,In_418);
and U72 (N_72,In_123,In_117);
nand U73 (N_73,In_308,In_57);
xnor U74 (N_74,In_208,In_118);
nor U75 (N_75,In_253,In_22);
nor U76 (N_76,In_341,In_29);
nor U77 (N_77,In_282,In_285);
nand U78 (N_78,In_101,In_40);
or U79 (N_79,In_310,In_303);
nor U80 (N_80,In_337,In_49);
nor U81 (N_81,In_373,In_275);
nand U82 (N_82,In_51,In_221);
nand U83 (N_83,In_211,In_76);
nand U84 (N_84,In_483,In_255);
and U85 (N_85,In_315,In_60);
and U86 (N_86,In_381,In_196);
or U87 (N_87,In_494,In_173);
nor U88 (N_88,In_451,In_394);
and U89 (N_89,In_423,In_379);
and U90 (N_90,In_403,In_219);
nor U91 (N_91,In_139,In_370);
nor U92 (N_92,In_20,In_38);
xnor U93 (N_93,In_431,In_82);
xnor U94 (N_94,In_272,In_45);
nor U95 (N_95,In_81,In_129);
nor U96 (N_96,In_9,In_407);
nor U97 (N_97,In_276,In_289);
nand U98 (N_98,In_333,In_178);
nand U99 (N_99,In_96,In_249);
or U100 (N_100,In_321,In_435);
and U101 (N_101,In_140,In_88);
or U102 (N_102,In_75,In_165);
nor U103 (N_103,In_56,In_214);
nor U104 (N_104,In_317,In_467);
nand U105 (N_105,In_447,In_106);
nor U106 (N_106,In_446,In_356);
xnor U107 (N_107,In_355,In_476);
xor U108 (N_108,In_136,In_230);
xnor U109 (N_109,In_419,In_229);
nand U110 (N_110,In_122,In_186);
or U111 (N_111,In_34,In_152);
nand U112 (N_112,In_380,In_137);
and U113 (N_113,In_455,In_223);
nand U114 (N_114,In_141,In_475);
nand U115 (N_115,In_322,In_158);
nor U116 (N_116,In_39,In_436);
nand U117 (N_117,In_166,In_69);
nor U118 (N_118,In_89,In_159);
nand U119 (N_119,In_126,In_401);
and U120 (N_120,In_148,In_338);
xnor U121 (N_121,In_26,In_490);
nor U122 (N_122,In_65,In_464);
nand U123 (N_123,In_33,In_194);
or U124 (N_124,In_264,In_67);
nor U125 (N_125,In_187,In_382);
and U126 (N_126,In_257,In_458);
nor U127 (N_127,In_31,In_228);
nor U128 (N_128,In_486,In_288);
nor U129 (N_129,In_100,In_91);
or U130 (N_130,In_213,In_115);
nand U131 (N_131,In_47,In_369);
nand U132 (N_132,In_357,In_396);
xnor U133 (N_133,In_201,In_367);
nand U134 (N_134,In_225,In_204);
or U135 (N_135,In_293,In_36);
or U136 (N_136,In_411,In_160);
nor U137 (N_137,In_397,In_359);
or U138 (N_138,In_42,In_99);
and U139 (N_139,In_28,In_70);
xor U140 (N_140,In_35,In_50);
or U141 (N_141,In_109,In_177);
xor U142 (N_142,In_410,In_393);
and U143 (N_143,In_283,In_216);
or U144 (N_144,In_325,In_262);
and U145 (N_145,In_180,In_374);
or U146 (N_146,In_37,In_332);
xnor U147 (N_147,In_426,In_468);
nor U148 (N_148,In_449,In_237);
or U149 (N_149,In_434,In_238);
nor U150 (N_150,In_354,In_344);
xor U151 (N_151,In_93,In_450);
nand U152 (N_152,In_167,In_312);
or U153 (N_153,In_13,In_445);
and U154 (N_154,In_235,In_343);
and U155 (N_155,In_113,In_459);
nand U156 (N_156,In_353,In_59);
xnor U157 (N_157,In_90,In_437);
and U158 (N_158,In_348,In_71);
nor U159 (N_159,In_304,In_30);
nor U160 (N_160,In_292,In_491);
or U161 (N_161,In_345,In_64);
nor U162 (N_162,In_103,In_181);
xor U163 (N_163,In_105,In_16);
and U164 (N_164,In_439,In_266);
nor U165 (N_165,In_339,In_480);
nand U166 (N_166,In_302,In_346);
and U167 (N_167,In_477,In_4);
nor U168 (N_168,In_277,In_472);
nand U169 (N_169,In_72,In_386);
and U170 (N_170,In_74,In_273);
or U171 (N_171,In_184,In_162);
nor U172 (N_172,In_252,In_300);
and U173 (N_173,In_5,In_169);
and U174 (N_174,In_335,In_398);
nand U175 (N_175,In_243,In_328);
nand U176 (N_176,In_424,In_154);
xnor U177 (N_177,In_112,In_478);
nor U178 (N_178,In_408,In_156);
and U179 (N_179,In_421,In_104);
or U180 (N_180,In_487,In_363);
or U181 (N_181,In_364,In_461);
or U182 (N_182,In_21,In_149);
nor U183 (N_183,In_299,In_195);
nand U184 (N_184,In_233,In_412);
xnor U185 (N_185,In_58,In_438);
or U186 (N_186,In_404,In_495);
nand U187 (N_187,In_469,In_298);
and U188 (N_188,In_189,In_430);
nand U189 (N_189,In_98,In_271);
and U190 (N_190,In_143,In_433);
nor U191 (N_191,In_360,In_425);
nor U192 (N_192,In_371,In_366);
or U193 (N_193,In_87,In_54);
nand U194 (N_194,In_440,In_175);
or U195 (N_195,In_174,In_395);
and U196 (N_196,In_18,In_296);
nand U197 (N_197,In_155,In_172);
nand U198 (N_198,In_207,In_267);
nand U199 (N_199,In_142,In_107);
nor U200 (N_200,In_1,In_307);
nand U201 (N_201,N_129,N_87);
nor U202 (N_202,In_2,N_196);
and U203 (N_203,N_144,N_104);
nor U204 (N_204,In_281,N_50);
nor U205 (N_205,N_70,In_417);
nor U206 (N_206,N_121,In_448);
nor U207 (N_207,N_59,N_26);
and U208 (N_208,N_36,N_157);
and U209 (N_209,N_147,N_187);
nand U210 (N_210,In_362,N_34);
or U211 (N_211,N_130,N_38);
and U212 (N_212,N_43,N_161);
and U213 (N_213,N_162,N_137);
nand U214 (N_214,N_6,N_178);
nor U215 (N_215,N_169,In_3);
and U216 (N_216,In_188,N_167);
nor U217 (N_217,In_443,In_11);
or U218 (N_218,In_316,N_84);
or U219 (N_219,In_176,N_106);
or U220 (N_220,N_71,In_147);
nand U221 (N_221,N_37,N_9);
nand U222 (N_222,N_95,In_32);
or U223 (N_223,N_25,In_460);
nand U224 (N_224,N_41,In_193);
xor U225 (N_225,N_176,In_258);
or U226 (N_226,N_81,N_64);
nor U227 (N_227,N_153,N_175);
nand U228 (N_228,In_479,N_16);
nor U229 (N_229,N_126,N_125);
nor U230 (N_230,In_124,N_116);
and U231 (N_231,In_422,N_15);
nand U232 (N_232,In_351,N_94);
xnor U233 (N_233,In_427,N_140);
and U234 (N_234,In_94,N_1);
xor U235 (N_235,N_57,N_63);
nor U236 (N_236,In_305,N_148);
and U237 (N_237,N_164,In_290);
nand U238 (N_238,In_391,N_99);
nor U239 (N_239,In_388,In_392);
or U240 (N_240,In_224,N_73);
nand U241 (N_241,N_188,N_173);
nor U242 (N_242,N_139,N_168);
or U243 (N_243,N_75,N_105);
nor U244 (N_244,N_24,N_96);
or U245 (N_245,N_183,N_2);
nor U246 (N_246,N_151,N_179);
and U247 (N_247,N_160,In_350);
nand U248 (N_248,In_206,N_150);
nor U249 (N_249,N_80,N_155);
and U250 (N_250,N_159,In_78);
nor U251 (N_251,In_114,N_45);
nor U252 (N_252,N_66,N_65);
nand U253 (N_253,N_127,In_179);
or U254 (N_254,In_73,N_93);
and U255 (N_255,N_193,In_306);
and U256 (N_256,In_265,N_10);
nand U257 (N_257,N_107,N_29);
nor U258 (N_258,N_54,N_101);
nand U259 (N_259,In_340,In_294);
nor U260 (N_260,N_182,N_194);
or U261 (N_261,N_18,N_119);
xor U262 (N_262,N_112,N_171);
and U263 (N_263,In_474,N_172);
nand U264 (N_264,N_11,N_100);
and U265 (N_265,N_78,N_74);
or U266 (N_266,N_32,In_146);
and U267 (N_267,N_102,N_86);
nand U268 (N_268,N_28,In_334);
or U269 (N_269,In_256,N_103);
nand U270 (N_270,N_141,N_166);
nor U271 (N_271,In_8,In_349);
or U272 (N_272,N_3,N_198);
nand U273 (N_273,In_144,N_67);
nor U274 (N_274,N_118,N_8);
and U275 (N_275,N_4,N_55);
and U276 (N_276,N_195,N_138);
and U277 (N_277,N_149,N_7);
nand U278 (N_278,In_53,N_180);
or U279 (N_279,N_77,N_35);
and U280 (N_280,N_135,In_473);
nand U281 (N_281,In_135,N_111);
nor U282 (N_282,In_248,N_115);
nor U283 (N_283,In_171,N_48);
nor U284 (N_284,N_82,N_117);
and U285 (N_285,N_184,In_279);
or U286 (N_286,N_190,In_387);
nor U287 (N_287,N_13,N_185);
nand U288 (N_288,N_56,N_49);
xnor U289 (N_289,In_132,N_145);
and U290 (N_290,In_83,N_83);
or U291 (N_291,N_97,N_47);
or U292 (N_292,N_61,N_154);
nor U293 (N_293,In_465,N_33);
nor U294 (N_294,In_138,N_136);
or U295 (N_295,In_242,N_199);
and U296 (N_296,In_48,In_318);
nand U297 (N_297,N_158,N_52);
and U298 (N_298,N_156,N_0);
or U299 (N_299,In_55,N_146);
nor U300 (N_300,In_41,N_123);
and U301 (N_301,N_143,N_170);
nand U302 (N_302,N_114,In_241);
and U303 (N_303,N_5,N_98);
nand U304 (N_304,In_409,N_60);
nor U305 (N_305,N_31,In_254);
and U306 (N_306,In_376,N_191);
nor U307 (N_307,In_246,In_220);
or U308 (N_308,N_79,N_69);
nand U309 (N_309,N_197,In_198);
and U310 (N_310,N_189,In_365);
nand U311 (N_311,In_260,In_161);
nand U312 (N_312,In_311,In_52);
or U313 (N_313,N_40,N_27);
or U314 (N_314,N_22,N_30);
and U315 (N_315,N_89,N_14);
nor U316 (N_316,In_46,N_142);
nand U317 (N_317,N_51,N_12);
xor U318 (N_318,N_44,In_102);
and U319 (N_319,N_92,In_240);
nand U320 (N_320,N_113,N_174);
and U321 (N_321,In_378,In_116);
or U322 (N_322,N_85,In_313);
nand U323 (N_323,N_21,In_323);
nor U324 (N_324,N_165,In_481);
or U325 (N_325,N_128,N_186);
and U326 (N_326,In_263,N_131);
nor U327 (N_327,N_110,N_134);
and U328 (N_328,N_23,N_68);
and U329 (N_329,N_177,N_19);
nor U330 (N_330,N_53,In_62);
and U331 (N_331,In_377,In_10);
xnor U332 (N_332,N_62,N_152);
nand U333 (N_333,N_72,In_463);
and U334 (N_334,N_46,N_132);
nand U335 (N_335,In_492,N_108);
nand U336 (N_336,N_120,N_39);
and U337 (N_337,N_192,In_361);
nor U338 (N_338,N_20,N_122);
xnor U339 (N_339,In_295,N_91);
or U340 (N_340,In_415,N_109);
or U341 (N_341,In_372,N_90);
and U342 (N_342,In_205,N_163);
nor U343 (N_343,In_23,N_42);
nand U344 (N_344,In_259,In_234);
nor U345 (N_345,N_76,N_124);
and U346 (N_346,In_456,In_153);
nand U347 (N_347,N_58,N_88);
nand U348 (N_348,N_181,In_7);
and U349 (N_349,N_17,N_133);
nand U350 (N_350,N_34,N_147);
and U351 (N_351,N_9,N_80);
nor U352 (N_352,N_184,In_10);
and U353 (N_353,N_134,N_50);
nand U354 (N_354,In_260,N_95);
nand U355 (N_355,In_46,In_176);
or U356 (N_356,In_83,In_193);
and U357 (N_357,In_306,N_101);
nand U358 (N_358,N_113,N_2);
nor U359 (N_359,N_160,N_144);
nor U360 (N_360,N_50,N_71);
or U361 (N_361,N_47,N_119);
or U362 (N_362,N_155,N_166);
nor U363 (N_363,In_290,In_377);
or U364 (N_364,In_492,N_157);
nand U365 (N_365,N_136,N_173);
nand U366 (N_366,N_10,In_193);
nor U367 (N_367,N_173,N_138);
and U368 (N_368,In_161,N_106);
nor U369 (N_369,In_281,N_42);
and U370 (N_370,N_55,In_171);
nand U371 (N_371,N_73,In_62);
xnor U372 (N_372,N_127,In_248);
nand U373 (N_373,N_84,In_116);
nand U374 (N_374,N_181,N_124);
nand U375 (N_375,N_133,N_81);
nor U376 (N_376,In_473,In_263);
nand U377 (N_377,In_281,N_28);
nor U378 (N_378,N_94,N_196);
xor U379 (N_379,In_365,N_11);
nand U380 (N_380,N_47,N_192);
nand U381 (N_381,N_125,N_3);
xnor U382 (N_382,In_259,N_197);
or U383 (N_383,N_104,In_365);
and U384 (N_384,N_123,N_131);
and U385 (N_385,N_46,N_59);
nor U386 (N_386,N_50,N_126);
xnor U387 (N_387,In_311,N_49);
and U388 (N_388,In_114,N_134);
nand U389 (N_389,N_57,N_176);
nor U390 (N_390,In_147,N_94);
and U391 (N_391,In_188,In_179);
nor U392 (N_392,N_168,N_95);
nor U393 (N_393,N_122,In_246);
xnor U394 (N_394,N_10,N_173);
and U395 (N_395,In_474,N_49);
nand U396 (N_396,N_35,N_69);
nand U397 (N_397,In_263,N_9);
nand U398 (N_398,N_71,In_409);
nand U399 (N_399,In_260,N_104);
or U400 (N_400,N_296,N_377);
and U401 (N_401,N_203,N_213);
nand U402 (N_402,N_276,N_343);
nor U403 (N_403,N_378,N_304);
and U404 (N_404,N_201,N_389);
nand U405 (N_405,N_279,N_216);
or U406 (N_406,N_372,N_281);
nor U407 (N_407,N_282,N_251);
and U408 (N_408,N_268,N_208);
and U409 (N_409,N_395,N_374);
nor U410 (N_410,N_223,N_301);
and U411 (N_411,N_326,N_212);
nand U412 (N_412,N_332,N_253);
or U413 (N_413,N_250,N_324);
nor U414 (N_414,N_278,N_215);
or U415 (N_415,N_323,N_340);
nor U416 (N_416,N_351,N_328);
and U417 (N_417,N_355,N_202);
nor U418 (N_418,N_360,N_295);
or U419 (N_419,N_273,N_393);
and U420 (N_420,N_277,N_322);
nor U421 (N_421,N_225,N_342);
xor U422 (N_422,N_238,N_298);
and U423 (N_423,N_233,N_263);
nor U424 (N_424,N_347,N_361);
or U425 (N_425,N_362,N_310);
nand U426 (N_426,N_200,N_205);
and U427 (N_427,N_339,N_218);
xnor U428 (N_428,N_386,N_232);
nor U429 (N_429,N_337,N_290);
and U430 (N_430,N_221,N_266);
or U431 (N_431,N_239,N_317);
or U432 (N_432,N_248,N_262);
or U433 (N_433,N_204,N_283);
nor U434 (N_434,N_256,N_396);
and U435 (N_435,N_359,N_388);
nor U436 (N_436,N_382,N_379);
nand U437 (N_437,N_292,N_207);
or U438 (N_438,N_274,N_289);
nor U439 (N_439,N_210,N_315);
nor U440 (N_440,N_391,N_269);
nor U441 (N_441,N_270,N_261);
or U442 (N_442,N_217,N_333);
nand U443 (N_443,N_222,N_398);
or U444 (N_444,N_257,N_285);
xnor U445 (N_445,N_275,N_329);
nand U446 (N_446,N_381,N_231);
nand U447 (N_447,N_272,N_319);
and U448 (N_448,N_247,N_363);
and U449 (N_449,N_211,N_244);
nor U450 (N_450,N_305,N_299);
or U451 (N_451,N_380,N_294);
nor U452 (N_452,N_330,N_373);
nand U453 (N_453,N_255,N_287);
nand U454 (N_454,N_271,N_227);
nand U455 (N_455,N_311,N_334);
and U456 (N_456,N_242,N_325);
and U457 (N_457,N_387,N_376);
and U458 (N_458,N_397,N_369);
nor U459 (N_459,N_288,N_349);
nor U460 (N_460,N_254,N_246);
and U461 (N_461,N_224,N_314);
and U462 (N_462,N_243,N_300);
or U463 (N_463,N_209,N_241);
and U464 (N_464,N_371,N_370);
and U465 (N_465,N_358,N_367);
nand U466 (N_466,N_214,N_291);
nand U467 (N_467,N_318,N_338);
nor U468 (N_468,N_308,N_364);
or U469 (N_469,N_228,N_356);
and U470 (N_470,N_365,N_302);
nand U471 (N_471,N_220,N_354);
or U472 (N_472,N_249,N_252);
xor U473 (N_473,N_341,N_344);
nand U474 (N_474,N_384,N_335);
nor U475 (N_475,N_316,N_206);
and U476 (N_476,N_394,N_280);
nand U477 (N_477,N_237,N_235);
xnor U478 (N_478,N_368,N_345);
nand U479 (N_479,N_383,N_353);
nor U480 (N_480,N_284,N_321);
or U481 (N_481,N_390,N_348);
and U482 (N_482,N_240,N_327);
nor U483 (N_483,N_357,N_350);
nand U484 (N_484,N_307,N_346);
nand U485 (N_485,N_259,N_306);
nand U486 (N_486,N_297,N_392);
and U487 (N_487,N_336,N_258);
nor U488 (N_488,N_331,N_264);
or U489 (N_489,N_375,N_230);
or U490 (N_490,N_385,N_245);
nand U491 (N_491,N_309,N_234);
or U492 (N_492,N_219,N_265);
or U493 (N_493,N_313,N_320);
xor U494 (N_494,N_229,N_312);
nor U495 (N_495,N_293,N_352);
and U496 (N_496,N_260,N_267);
or U497 (N_497,N_399,N_303);
nor U498 (N_498,N_226,N_236);
nand U499 (N_499,N_366,N_286);
and U500 (N_500,N_394,N_296);
nor U501 (N_501,N_231,N_252);
nor U502 (N_502,N_350,N_250);
nor U503 (N_503,N_350,N_262);
nand U504 (N_504,N_341,N_252);
nand U505 (N_505,N_234,N_210);
and U506 (N_506,N_205,N_392);
nor U507 (N_507,N_382,N_357);
nand U508 (N_508,N_397,N_264);
xor U509 (N_509,N_213,N_369);
or U510 (N_510,N_335,N_332);
nand U511 (N_511,N_381,N_228);
or U512 (N_512,N_313,N_390);
nand U513 (N_513,N_231,N_294);
nand U514 (N_514,N_359,N_314);
nand U515 (N_515,N_376,N_379);
or U516 (N_516,N_383,N_321);
or U517 (N_517,N_326,N_324);
nor U518 (N_518,N_336,N_344);
and U519 (N_519,N_294,N_252);
xor U520 (N_520,N_222,N_390);
nor U521 (N_521,N_338,N_395);
nor U522 (N_522,N_356,N_304);
and U523 (N_523,N_362,N_206);
xnor U524 (N_524,N_331,N_267);
or U525 (N_525,N_217,N_345);
nor U526 (N_526,N_383,N_333);
and U527 (N_527,N_333,N_331);
and U528 (N_528,N_299,N_312);
nand U529 (N_529,N_275,N_216);
nor U530 (N_530,N_367,N_330);
nand U531 (N_531,N_299,N_260);
or U532 (N_532,N_339,N_247);
or U533 (N_533,N_320,N_264);
nor U534 (N_534,N_392,N_359);
and U535 (N_535,N_224,N_395);
and U536 (N_536,N_247,N_233);
or U537 (N_537,N_334,N_227);
nand U538 (N_538,N_211,N_208);
nor U539 (N_539,N_389,N_326);
or U540 (N_540,N_214,N_391);
and U541 (N_541,N_333,N_274);
nand U542 (N_542,N_392,N_282);
nand U543 (N_543,N_346,N_375);
nor U544 (N_544,N_355,N_338);
and U545 (N_545,N_225,N_273);
nor U546 (N_546,N_305,N_223);
nand U547 (N_547,N_254,N_212);
or U548 (N_548,N_281,N_338);
nor U549 (N_549,N_205,N_287);
nand U550 (N_550,N_205,N_288);
nor U551 (N_551,N_284,N_316);
nand U552 (N_552,N_209,N_306);
and U553 (N_553,N_268,N_261);
nor U554 (N_554,N_330,N_345);
or U555 (N_555,N_278,N_259);
and U556 (N_556,N_335,N_245);
or U557 (N_557,N_302,N_355);
nand U558 (N_558,N_211,N_225);
or U559 (N_559,N_355,N_342);
nor U560 (N_560,N_337,N_286);
or U561 (N_561,N_324,N_390);
nor U562 (N_562,N_251,N_272);
and U563 (N_563,N_237,N_256);
nand U564 (N_564,N_306,N_372);
and U565 (N_565,N_328,N_336);
nor U566 (N_566,N_321,N_310);
and U567 (N_567,N_328,N_246);
nand U568 (N_568,N_306,N_283);
nor U569 (N_569,N_294,N_264);
xnor U570 (N_570,N_395,N_202);
xnor U571 (N_571,N_357,N_338);
and U572 (N_572,N_214,N_213);
nor U573 (N_573,N_277,N_236);
nand U574 (N_574,N_233,N_258);
nor U575 (N_575,N_261,N_254);
or U576 (N_576,N_260,N_325);
nand U577 (N_577,N_320,N_279);
and U578 (N_578,N_220,N_329);
nor U579 (N_579,N_238,N_310);
nand U580 (N_580,N_254,N_252);
nand U581 (N_581,N_285,N_352);
or U582 (N_582,N_305,N_254);
xnor U583 (N_583,N_289,N_376);
nor U584 (N_584,N_354,N_323);
and U585 (N_585,N_395,N_216);
nor U586 (N_586,N_269,N_222);
nand U587 (N_587,N_330,N_281);
nor U588 (N_588,N_221,N_244);
or U589 (N_589,N_257,N_329);
and U590 (N_590,N_248,N_364);
or U591 (N_591,N_388,N_318);
or U592 (N_592,N_231,N_276);
nand U593 (N_593,N_320,N_352);
and U594 (N_594,N_351,N_382);
and U595 (N_595,N_370,N_347);
nor U596 (N_596,N_246,N_251);
nor U597 (N_597,N_260,N_275);
or U598 (N_598,N_337,N_328);
nor U599 (N_599,N_337,N_329);
nand U600 (N_600,N_521,N_417);
or U601 (N_601,N_524,N_549);
and U602 (N_602,N_447,N_473);
nand U603 (N_603,N_481,N_562);
nand U604 (N_604,N_418,N_449);
or U605 (N_605,N_464,N_500);
nand U606 (N_606,N_561,N_408);
or U607 (N_607,N_434,N_499);
nand U608 (N_608,N_593,N_427);
xor U609 (N_609,N_528,N_520);
or U610 (N_610,N_595,N_517);
and U611 (N_611,N_444,N_410);
nand U612 (N_612,N_443,N_547);
nand U613 (N_613,N_483,N_507);
nand U614 (N_614,N_510,N_541);
nor U615 (N_615,N_453,N_498);
nor U616 (N_616,N_576,N_506);
or U617 (N_617,N_597,N_514);
nor U618 (N_618,N_455,N_589);
nor U619 (N_619,N_565,N_594);
nand U620 (N_620,N_573,N_470);
and U621 (N_621,N_530,N_463);
xor U622 (N_622,N_478,N_582);
nor U623 (N_623,N_441,N_508);
or U624 (N_624,N_446,N_414);
nand U625 (N_625,N_495,N_445);
and U626 (N_626,N_590,N_402);
nand U627 (N_627,N_407,N_485);
or U628 (N_628,N_522,N_502);
and U629 (N_629,N_525,N_489);
and U630 (N_630,N_543,N_542);
and U631 (N_631,N_511,N_580);
and U632 (N_632,N_513,N_527);
and U633 (N_633,N_454,N_532);
or U634 (N_634,N_574,N_544);
nor U635 (N_635,N_493,N_588);
xnor U636 (N_636,N_433,N_519);
nor U637 (N_637,N_570,N_459);
nand U638 (N_638,N_404,N_421);
nand U639 (N_639,N_428,N_553);
nand U640 (N_640,N_509,N_581);
nand U641 (N_641,N_531,N_467);
and U642 (N_642,N_462,N_585);
or U643 (N_643,N_490,N_450);
or U644 (N_644,N_476,N_523);
and U645 (N_645,N_496,N_566);
nand U646 (N_646,N_458,N_461);
nor U647 (N_647,N_409,N_599);
xnor U648 (N_648,N_480,N_424);
and U649 (N_649,N_457,N_540);
or U650 (N_650,N_555,N_534);
nor U651 (N_651,N_429,N_487);
nor U652 (N_652,N_503,N_557);
or U653 (N_653,N_563,N_430);
nor U654 (N_654,N_515,N_419);
nand U655 (N_655,N_479,N_415);
nor U656 (N_656,N_488,N_413);
nor U657 (N_657,N_596,N_504);
and U658 (N_658,N_539,N_516);
or U659 (N_659,N_512,N_583);
nor U660 (N_660,N_571,N_431);
nand U661 (N_661,N_405,N_587);
nor U662 (N_662,N_411,N_578);
nand U663 (N_663,N_400,N_559);
and U664 (N_664,N_469,N_468);
nor U665 (N_665,N_475,N_586);
or U666 (N_666,N_577,N_472);
nor U667 (N_667,N_422,N_505);
nand U668 (N_668,N_437,N_584);
nand U669 (N_669,N_567,N_451);
nand U670 (N_670,N_448,N_435);
nor U671 (N_671,N_403,N_484);
nand U672 (N_672,N_533,N_569);
nor U673 (N_673,N_406,N_526);
or U674 (N_674,N_564,N_416);
or U675 (N_675,N_466,N_420);
nand U676 (N_676,N_438,N_529);
nor U677 (N_677,N_538,N_572);
xnor U678 (N_678,N_497,N_494);
or U679 (N_679,N_545,N_432);
nor U680 (N_680,N_554,N_551);
nand U681 (N_681,N_536,N_560);
nor U682 (N_682,N_492,N_401);
nand U683 (N_683,N_477,N_423);
xnor U684 (N_684,N_592,N_579);
and U685 (N_685,N_442,N_568);
xnor U686 (N_686,N_546,N_591);
or U687 (N_687,N_537,N_425);
or U688 (N_688,N_518,N_491);
or U689 (N_689,N_482,N_440);
xor U690 (N_690,N_452,N_486);
nor U691 (N_691,N_575,N_474);
and U692 (N_692,N_439,N_598);
nand U693 (N_693,N_550,N_535);
xor U694 (N_694,N_465,N_558);
nand U695 (N_695,N_501,N_556);
or U696 (N_696,N_426,N_436);
nor U697 (N_697,N_456,N_460);
nand U698 (N_698,N_552,N_412);
or U699 (N_699,N_548,N_471);
nand U700 (N_700,N_587,N_470);
xor U701 (N_701,N_504,N_430);
or U702 (N_702,N_483,N_562);
xor U703 (N_703,N_546,N_417);
nor U704 (N_704,N_539,N_520);
and U705 (N_705,N_405,N_459);
nor U706 (N_706,N_464,N_470);
nor U707 (N_707,N_551,N_576);
nor U708 (N_708,N_503,N_494);
or U709 (N_709,N_504,N_410);
nor U710 (N_710,N_507,N_458);
or U711 (N_711,N_525,N_428);
or U712 (N_712,N_555,N_564);
or U713 (N_713,N_533,N_577);
and U714 (N_714,N_566,N_492);
nor U715 (N_715,N_437,N_445);
nor U716 (N_716,N_572,N_540);
xnor U717 (N_717,N_561,N_478);
xor U718 (N_718,N_463,N_483);
nor U719 (N_719,N_598,N_558);
or U720 (N_720,N_504,N_592);
nand U721 (N_721,N_406,N_466);
and U722 (N_722,N_454,N_424);
and U723 (N_723,N_592,N_419);
and U724 (N_724,N_519,N_450);
and U725 (N_725,N_485,N_537);
xor U726 (N_726,N_483,N_431);
nand U727 (N_727,N_478,N_509);
xor U728 (N_728,N_423,N_439);
and U729 (N_729,N_423,N_406);
nor U730 (N_730,N_565,N_499);
xnor U731 (N_731,N_546,N_599);
nand U732 (N_732,N_519,N_590);
nand U733 (N_733,N_460,N_429);
nor U734 (N_734,N_446,N_482);
nand U735 (N_735,N_535,N_553);
or U736 (N_736,N_577,N_548);
or U737 (N_737,N_515,N_516);
nand U738 (N_738,N_532,N_442);
nor U739 (N_739,N_410,N_574);
nor U740 (N_740,N_525,N_567);
and U741 (N_741,N_528,N_580);
or U742 (N_742,N_429,N_497);
xnor U743 (N_743,N_506,N_549);
or U744 (N_744,N_508,N_547);
xor U745 (N_745,N_484,N_534);
nor U746 (N_746,N_536,N_423);
nand U747 (N_747,N_555,N_586);
or U748 (N_748,N_569,N_495);
and U749 (N_749,N_418,N_537);
nor U750 (N_750,N_407,N_443);
or U751 (N_751,N_523,N_473);
xnor U752 (N_752,N_597,N_455);
xor U753 (N_753,N_589,N_580);
nor U754 (N_754,N_456,N_465);
nand U755 (N_755,N_564,N_418);
nor U756 (N_756,N_440,N_596);
or U757 (N_757,N_580,N_488);
or U758 (N_758,N_493,N_440);
and U759 (N_759,N_432,N_491);
nor U760 (N_760,N_463,N_419);
nor U761 (N_761,N_467,N_426);
or U762 (N_762,N_525,N_444);
or U763 (N_763,N_510,N_433);
nor U764 (N_764,N_417,N_480);
nor U765 (N_765,N_478,N_475);
nand U766 (N_766,N_492,N_576);
and U767 (N_767,N_428,N_474);
nor U768 (N_768,N_479,N_446);
and U769 (N_769,N_520,N_434);
and U770 (N_770,N_490,N_588);
and U771 (N_771,N_428,N_511);
nor U772 (N_772,N_431,N_416);
nor U773 (N_773,N_405,N_540);
nor U774 (N_774,N_598,N_497);
nand U775 (N_775,N_561,N_467);
xor U776 (N_776,N_404,N_457);
or U777 (N_777,N_491,N_479);
nand U778 (N_778,N_492,N_467);
and U779 (N_779,N_424,N_422);
or U780 (N_780,N_561,N_587);
or U781 (N_781,N_450,N_500);
and U782 (N_782,N_526,N_440);
nor U783 (N_783,N_541,N_547);
or U784 (N_784,N_557,N_516);
nand U785 (N_785,N_448,N_510);
and U786 (N_786,N_487,N_459);
nor U787 (N_787,N_414,N_443);
or U788 (N_788,N_514,N_571);
or U789 (N_789,N_577,N_494);
or U790 (N_790,N_537,N_558);
nand U791 (N_791,N_449,N_577);
xor U792 (N_792,N_539,N_499);
nor U793 (N_793,N_584,N_591);
and U794 (N_794,N_569,N_412);
and U795 (N_795,N_412,N_578);
and U796 (N_796,N_489,N_482);
nor U797 (N_797,N_493,N_451);
and U798 (N_798,N_540,N_496);
xnor U799 (N_799,N_427,N_453);
and U800 (N_800,N_770,N_678);
nand U801 (N_801,N_662,N_723);
nor U802 (N_802,N_722,N_633);
nor U803 (N_803,N_734,N_666);
and U804 (N_804,N_772,N_744);
nand U805 (N_805,N_602,N_753);
and U806 (N_806,N_785,N_653);
or U807 (N_807,N_671,N_726);
nand U808 (N_808,N_679,N_790);
and U809 (N_809,N_637,N_645);
or U810 (N_810,N_618,N_698);
nor U811 (N_811,N_616,N_787);
nand U812 (N_812,N_651,N_783);
and U813 (N_813,N_699,N_688);
nor U814 (N_814,N_605,N_740);
nor U815 (N_815,N_642,N_631);
and U816 (N_816,N_617,N_661);
xnor U817 (N_817,N_696,N_748);
xor U818 (N_818,N_650,N_792);
or U819 (N_819,N_768,N_669);
and U820 (N_820,N_766,N_708);
nor U821 (N_821,N_784,N_691);
and U822 (N_822,N_647,N_683);
or U823 (N_823,N_771,N_764);
nand U824 (N_824,N_632,N_627);
and U825 (N_825,N_675,N_603);
nor U826 (N_826,N_735,N_635);
nor U827 (N_827,N_695,N_686);
or U828 (N_828,N_614,N_724);
and U829 (N_829,N_659,N_737);
and U830 (N_830,N_681,N_777);
nand U831 (N_831,N_743,N_611);
xnor U832 (N_832,N_747,N_796);
nand U833 (N_833,N_621,N_622);
nand U834 (N_834,N_758,N_655);
nor U835 (N_835,N_711,N_652);
or U836 (N_836,N_721,N_729);
nand U837 (N_837,N_780,N_640);
and U838 (N_838,N_791,N_638);
and U839 (N_839,N_776,N_730);
and U840 (N_840,N_755,N_704);
nor U841 (N_841,N_738,N_763);
and U842 (N_842,N_630,N_687);
and U843 (N_843,N_667,N_767);
nand U844 (N_844,N_705,N_750);
nand U845 (N_845,N_676,N_778);
nor U846 (N_846,N_794,N_749);
and U847 (N_847,N_690,N_693);
nand U848 (N_848,N_646,N_754);
nor U849 (N_849,N_761,N_673);
or U850 (N_850,N_782,N_709);
or U851 (N_851,N_786,N_628);
or U852 (N_852,N_774,N_719);
and U853 (N_853,N_615,N_702);
and U854 (N_854,N_643,N_689);
nor U855 (N_855,N_715,N_619);
xor U856 (N_856,N_793,N_757);
nand U857 (N_857,N_641,N_625);
and U858 (N_858,N_692,N_649);
or U859 (N_859,N_733,N_701);
and U860 (N_860,N_684,N_680);
and U861 (N_861,N_613,N_658);
or U862 (N_862,N_656,N_798);
and U863 (N_863,N_665,N_685);
and U864 (N_864,N_736,N_712);
or U865 (N_865,N_677,N_670);
or U866 (N_866,N_718,N_720);
or U867 (N_867,N_788,N_795);
nand U868 (N_868,N_752,N_639);
or U869 (N_869,N_773,N_604);
and U870 (N_870,N_725,N_600);
nor U871 (N_871,N_742,N_716);
nor U872 (N_872,N_769,N_739);
nor U873 (N_873,N_657,N_797);
nor U874 (N_874,N_612,N_608);
nor U875 (N_875,N_756,N_674);
nand U876 (N_876,N_745,N_728);
nand U877 (N_877,N_765,N_707);
nor U878 (N_878,N_606,N_746);
nor U879 (N_879,N_751,N_775);
or U880 (N_880,N_629,N_713);
or U881 (N_881,N_636,N_732);
and U882 (N_882,N_700,N_623);
and U883 (N_883,N_731,N_703);
nand U884 (N_884,N_660,N_609);
nand U885 (N_885,N_634,N_672);
nor U886 (N_886,N_610,N_644);
xor U887 (N_887,N_779,N_668);
nand U888 (N_888,N_663,N_620);
nand U889 (N_889,N_601,N_781);
or U890 (N_890,N_710,N_624);
nor U891 (N_891,N_706,N_694);
nand U892 (N_892,N_648,N_799);
nor U893 (N_893,N_607,N_760);
and U894 (N_894,N_626,N_664);
and U895 (N_895,N_714,N_727);
and U896 (N_896,N_759,N_654);
or U897 (N_897,N_762,N_682);
nor U898 (N_898,N_717,N_741);
nor U899 (N_899,N_789,N_697);
and U900 (N_900,N_743,N_632);
nor U901 (N_901,N_645,N_757);
or U902 (N_902,N_746,N_732);
and U903 (N_903,N_766,N_624);
xor U904 (N_904,N_779,N_667);
and U905 (N_905,N_627,N_658);
and U906 (N_906,N_749,N_637);
and U907 (N_907,N_658,N_750);
nor U908 (N_908,N_606,N_747);
xor U909 (N_909,N_603,N_654);
xor U910 (N_910,N_712,N_765);
or U911 (N_911,N_697,N_709);
and U912 (N_912,N_740,N_699);
and U913 (N_913,N_698,N_794);
and U914 (N_914,N_629,N_738);
nor U915 (N_915,N_746,N_799);
and U916 (N_916,N_608,N_753);
or U917 (N_917,N_792,N_606);
nand U918 (N_918,N_782,N_610);
xnor U919 (N_919,N_606,N_646);
nand U920 (N_920,N_674,N_788);
nand U921 (N_921,N_658,N_684);
and U922 (N_922,N_622,N_793);
nor U923 (N_923,N_792,N_705);
nor U924 (N_924,N_721,N_672);
or U925 (N_925,N_644,N_780);
and U926 (N_926,N_613,N_684);
or U927 (N_927,N_731,N_660);
nand U928 (N_928,N_665,N_719);
nor U929 (N_929,N_663,N_609);
and U930 (N_930,N_681,N_792);
or U931 (N_931,N_681,N_729);
xnor U932 (N_932,N_795,N_675);
nor U933 (N_933,N_749,N_761);
xor U934 (N_934,N_723,N_706);
nor U935 (N_935,N_647,N_658);
nor U936 (N_936,N_704,N_780);
xor U937 (N_937,N_691,N_717);
xnor U938 (N_938,N_677,N_700);
nand U939 (N_939,N_778,N_653);
nor U940 (N_940,N_608,N_768);
nor U941 (N_941,N_600,N_687);
or U942 (N_942,N_613,N_676);
nor U943 (N_943,N_684,N_645);
nand U944 (N_944,N_761,N_745);
nor U945 (N_945,N_621,N_616);
nor U946 (N_946,N_715,N_609);
or U947 (N_947,N_691,N_618);
or U948 (N_948,N_609,N_639);
nor U949 (N_949,N_790,N_647);
or U950 (N_950,N_638,N_786);
and U951 (N_951,N_625,N_732);
nor U952 (N_952,N_624,N_687);
and U953 (N_953,N_619,N_762);
nand U954 (N_954,N_679,N_743);
nor U955 (N_955,N_750,N_674);
nand U956 (N_956,N_734,N_799);
xnor U957 (N_957,N_700,N_717);
or U958 (N_958,N_797,N_765);
or U959 (N_959,N_670,N_694);
nor U960 (N_960,N_642,N_601);
or U961 (N_961,N_639,N_712);
nor U962 (N_962,N_784,N_766);
or U963 (N_963,N_720,N_630);
or U964 (N_964,N_751,N_758);
nand U965 (N_965,N_634,N_771);
and U966 (N_966,N_654,N_782);
or U967 (N_967,N_618,N_714);
and U968 (N_968,N_613,N_705);
or U969 (N_969,N_656,N_786);
nor U970 (N_970,N_659,N_792);
or U971 (N_971,N_718,N_776);
xnor U972 (N_972,N_610,N_608);
xor U973 (N_973,N_609,N_749);
nor U974 (N_974,N_783,N_667);
nand U975 (N_975,N_728,N_644);
nand U976 (N_976,N_791,N_654);
or U977 (N_977,N_797,N_603);
nor U978 (N_978,N_602,N_689);
and U979 (N_979,N_752,N_676);
nor U980 (N_980,N_702,N_667);
or U981 (N_981,N_621,N_699);
or U982 (N_982,N_606,N_787);
nor U983 (N_983,N_723,N_635);
or U984 (N_984,N_678,N_797);
nand U985 (N_985,N_758,N_785);
and U986 (N_986,N_601,N_794);
xor U987 (N_987,N_686,N_652);
nand U988 (N_988,N_660,N_702);
nor U989 (N_989,N_762,N_644);
nand U990 (N_990,N_648,N_655);
and U991 (N_991,N_710,N_740);
nor U992 (N_992,N_751,N_760);
and U993 (N_993,N_696,N_677);
and U994 (N_994,N_708,N_726);
or U995 (N_995,N_652,N_660);
nand U996 (N_996,N_784,N_603);
or U997 (N_997,N_602,N_783);
nor U998 (N_998,N_615,N_787);
nor U999 (N_999,N_737,N_783);
nor U1000 (N_1000,N_819,N_898);
nor U1001 (N_1001,N_902,N_877);
and U1002 (N_1002,N_936,N_944);
or U1003 (N_1003,N_829,N_891);
or U1004 (N_1004,N_809,N_913);
and U1005 (N_1005,N_850,N_835);
nand U1006 (N_1006,N_893,N_808);
nor U1007 (N_1007,N_978,N_943);
nor U1008 (N_1008,N_910,N_836);
and U1009 (N_1009,N_875,N_803);
or U1010 (N_1010,N_823,N_991);
nand U1011 (N_1011,N_916,N_952);
or U1012 (N_1012,N_818,N_820);
nor U1013 (N_1013,N_919,N_946);
nor U1014 (N_1014,N_889,N_921);
nand U1015 (N_1015,N_970,N_924);
nand U1016 (N_1016,N_870,N_934);
and U1017 (N_1017,N_873,N_942);
nor U1018 (N_1018,N_865,N_941);
and U1019 (N_1019,N_988,N_949);
nand U1020 (N_1020,N_805,N_989);
nor U1021 (N_1021,N_860,N_918);
and U1022 (N_1022,N_849,N_866);
nand U1023 (N_1023,N_811,N_925);
xor U1024 (N_1024,N_998,N_983);
nor U1025 (N_1025,N_857,N_892);
nand U1026 (N_1026,N_985,N_960);
and U1027 (N_1027,N_801,N_879);
nor U1028 (N_1028,N_954,N_948);
and U1029 (N_1029,N_828,N_999);
nor U1030 (N_1030,N_896,N_871);
xnor U1031 (N_1031,N_982,N_832);
or U1032 (N_1032,N_996,N_872);
nor U1033 (N_1033,N_880,N_861);
nand U1034 (N_1034,N_881,N_974);
nand U1035 (N_1035,N_951,N_812);
nor U1036 (N_1036,N_980,N_838);
or U1037 (N_1037,N_917,N_800);
nor U1038 (N_1038,N_802,N_817);
nor U1039 (N_1039,N_862,N_926);
or U1040 (N_1040,N_968,N_844);
nor U1041 (N_1041,N_940,N_986);
and U1042 (N_1042,N_956,N_953);
or U1043 (N_1043,N_923,N_945);
nor U1044 (N_1044,N_930,N_843);
nand U1045 (N_1045,N_962,N_971);
or U1046 (N_1046,N_937,N_947);
nor U1047 (N_1047,N_905,N_842);
nand U1048 (N_1048,N_906,N_863);
nand U1049 (N_1049,N_884,N_848);
or U1050 (N_1050,N_839,N_987);
nor U1051 (N_1051,N_885,N_890);
nand U1052 (N_1052,N_837,N_966);
nand U1053 (N_1053,N_964,N_959);
nand U1054 (N_1054,N_977,N_826);
nand U1055 (N_1055,N_907,N_810);
and U1056 (N_1056,N_876,N_914);
or U1057 (N_1057,N_992,N_806);
and U1058 (N_1058,N_824,N_932);
nor U1059 (N_1059,N_858,N_864);
or U1060 (N_1060,N_928,N_939);
or U1061 (N_1061,N_869,N_868);
xor U1062 (N_1062,N_967,N_990);
or U1063 (N_1063,N_965,N_852);
or U1064 (N_1064,N_840,N_938);
nand U1065 (N_1065,N_899,N_845);
nor U1066 (N_1066,N_815,N_993);
nand U1067 (N_1067,N_894,N_908);
or U1068 (N_1068,N_927,N_833);
xor U1069 (N_1069,N_935,N_895);
nor U1070 (N_1070,N_855,N_958);
nor U1071 (N_1071,N_979,N_950);
nor U1072 (N_1072,N_909,N_834);
and U1073 (N_1073,N_981,N_851);
nand U1074 (N_1074,N_900,N_897);
nand U1075 (N_1075,N_911,N_874);
or U1076 (N_1076,N_867,N_901);
and U1077 (N_1077,N_882,N_853);
or U1078 (N_1078,N_846,N_878);
nor U1079 (N_1079,N_963,N_957);
nor U1080 (N_1080,N_929,N_822);
or U1081 (N_1081,N_827,N_969);
nand U1082 (N_1082,N_816,N_975);
nand U1083 (N_1083,N_994,N_831);
nor U1084 (N_1084,N_807,N_922);
and U1085 (N_1085,N_915,N_804);
xor U1086 (N_1086,N_886,N_972);
and U1087 (N_1087,N_888,N_931);
xor U1088 (N_1088,N_984,N_883);
or U1089 (N_1089,N_854,N_821);
nand U1090 (N_1090,N_997,N_903);
nand U1091 (N_1091,N_995,N_887);
nor U1092 (N_1092,N_904,N_973);
and U1093 (N_1093,N_856,N_847);
and U1094 (N_1094,N_961,N_933);
or U1095 (N_1095,N_920,N_825);
nand U1096 (N_1096,N_955,N_830);
nor U1097 (N_1097,N_912,N_813);
nor U1098 (N_1098,N_976,N_814);
or U1099 (N_1099,N_841,N_859);
nor U1100 (N_1100,N_844,N_949);
and U1101 (N_1101,N_869,N_877);
or U1102 (N_1102,N_965,N_842);
nor U1103 (N_1103,N_865,N_855);
nand U1104 (N_1104,N_825,N_979);
or U1105 (N_1105,N_917,N_965);
or U1106 (N_1106,N_837,N_983);
nor U1107 (N_1107,N_963,N_811);
and U1108 (N_1108,N_911,N_906);
nor U1109 (N_1109,N_819,N_890);
nor U1110 (N_1110,N_867,N_913);
and U1111 (N_1111,N_930,N_984);
nand U1112 (N_1112,N_815,N_838);
and U1113 (N_1113,N_981,N_832);
or U1114 (N_1114,N_998,N_839);
xnor U1115 (N_1115,N_816,N_847);
or U1116 (N_1116,N_819,N_973);
nor U1117 (N_1117,N_977,N_831);
or U1118 (N_1118,N_930,N_817);
or U1119 (N_1119,N_996,N_805);
nand U1120 (N_1120,N_831,N_845);
nand U1121 (N_1121,N_876,N_882);
and U1122 (N_1122,N_974,N_931);
or U1123 (N_1123,N_882,N_958);
and U1124 (N_1124,N_838,N_949);
nand U1125 (N_1125,N_826,N_833);
or U1126 (N_1126,N_806,N_960);
nand U1127 (N_1127,N_970,N_847);
and U1128 (N_1128,N_922,N_884);
and U1129 (N_1129,N_973,N_845);
nor U1130 (N_1130,N_959,N_895);
nor U1131 (N_1131,N_829,N_897);
and U1132 (N_1132,N_819,N_853);
nand U1133 (N_1133,N_862,N_982);
nor U1134 (N_1134,N_859,N_912);
and U1135 (N_1135,N_943,N_853);
nor U1136 (N_1136,N_876,N_965);
xor U1137 (N_1137,N_914,N_992);
nor U1138 (N_1138,N_996,N_987);
nand U1139 (N_1139,N_824,N_985);
or U1140 (N_1140,N_824,N_803);
nand U1141 (N_1141,N_918,N_915);
nor U1142 (N_1142,N_926,N_840);
or U1143 (N_1143,N_849,N_828);
nor U1144 (N_1144,N_827,N_814);
and U1145 (N_1145,N_810,N_804);
nand U1146 (N_1146,N_833,N_943);
nor U1147 (N_1147,N_818,N_926);
nor U1148 (N_1148,N_810,N_927);
nand U1149 (N_1149,N_967,N_858);
nor U1150 (N_1150,N_875,N_929);
or U1151 (N_1151,N_818,N_942);
xnor U1152 (N_1152,N_995,N_992);
nor U1153 (N_1153,N_919,N_881);
and U1154 (N_1154,N_989,N_802);
xnor U1155 (N_1155,N_897,N_957);
nor U1156 (N_1156,N_923,N_893);
or U1157 (N_1157,N_977,N_860);
nor U1158 (N_1158,N_908,N_817);
nor U1159 (N_1159,N_980,N_891);
nor U1160 (N_1160,N_804,N_969);
xnor U1161 (N_1161,N_882,N_972);
xor U1162 (N_1162,N_855,N_861);
or U1163 (N_1163,N_838,N_917);
xnor U1164 (N_1164,N_854,N_835);
and U1165 (N_1165,N_854,N_896);
and U1166 (N_1166,N_885,N_948);
xor U1167 (N_1167,N_872,N_808);
or U1168 (N_1168,N_849,N_874);
nand U1169 (N_1169,N_931,N_926);
nor U1170 (N_1170,N_900,N_886);
or U1171 (N_1171,N_860,N_829);
and U1172 (N_1172,N_883,N_845);
nand U1173 (N_1173,N_885,N_935);
nor U1174 (N_1174,N_896,N_997);
or U1175 (N_1175,N_910,N_949);
and U1176 (N_1176,N_953,N_835);
and U1177 (N_1177,N_933,N_993);
and U1178 (N_1178,N_945,N_982);
nand U1179 (N_1179,N_881,N_966);
and U1180 (N_1180,N_878,N_828);
nand U1181 (N_1181,N_986,N_840);
nor U1182 (N_1182,N_938,N_876);
nor U1183 (N_1183,N_873,N_917);
and U1184 (N_1184,N_818,N_940);
and U1185 (N_1185,N_822,N_937);
and U1186 (N_1186,N_821,N_988);
or U1187 (N_1187,N_872,N_970);
or U1188 (N_1188,N_948,N_985);
nor U1189 (N_1189,N_861,N_844);
and U1190 (N_1190,N_807,N_925);
nor U1191 (N_1191,N_938,N_862);
or U1192 (N_1192,N_908,N_890);
nor U1193 (N_1193,N_860,N_839);
or U1194 (N_1194,N_992,N_921);
or U1195 (N_1195,N_894,N_958);
nand U1196 (N_1196,N_870,N_929);
nor U1197 (N_1197,N_938,N_843);
nand U1198 (N_1198,N_961,N_870);
nand U1199 (N_1199,N_826,N_868);
nor U1200 (N_1200,N_1150,N_1072);
or U1201 (N_1201,N_1125,N_1083);
and U1202 (N_1202,N_1086,N_1011);
nor U1203 (N_1203,N_1053,N_1103);
and U1204 (N_1204,N_1171,N_1050);
and U1205 (N_1205,N_1193,N_1074);
and U1206 (N_1206,N_1000,N_1029);
nand U1207 (N_1207,N_1005,N_1087);
nand U1208 (N_1208,N_1049,N_1035);
nor U1209 (N_1209,N_1160,N_1131);
nor U1210 (N_1210,N_1180,N_1059);
and U1211 (N_1211,N_1143,N_1190);
xnor U1212 (N_1212,N_1196,N_1023);
xnor U1213 (N_1213,N_1199,N_1033);
xor U1214 (N_1214,N_1166,N_1060);
and U1215 (N_1215,N_1128,N_1032);
nand U1216 (N_1216,N_1172,N_1069);
and U1217 (N_1217,N_1066,N_1079);
nand U1218 (N_1218,N_1122,N_1198);
nand U1219 (N_1219,N_1110,N_1040);
or U1220 (N_1220,N_1186,N_1139);
and U1221 (N_1221,N_1115,N_1098);
or U1222 (N_1222,N_1149,N_1068);
and U1223 (N_1223,N_1124,N_1152);
nand U1224 (N_1224,N_1088,N_1127);
and U1225 (N_1225,N_1022,N_1157);
nand U1226 (N_1226,N_1082,N_1016);
nand U1227 (N_1227,N_1075,N_1030);
or U1228 (N_1228,N_1001,N_1179);
nor U1229 (N_1229,N_1104,N_1020);
nand U1230 (N_1230,N_1126,N_1167);
or U1231 (N_1231,N_1107,N_1177);
nand U1232 (N_1232,N_1043,N_1188);
nor U1233 (N_1233,N_1147,N_1056);
nor U1234 (N_1234,N_1194,N_1070);
or U1235 (N_1235,N_1117,N_1112);
nor U1236 (N_1236,N_1197,N_1006);
and U1237 (N_1237,N_1123,N_1034);
nand U1238 (N_1238,N_1192,N_1090);
nand U1239 (N_1239,N_1021,N_1114);
or U1240 (N_1240,N_1003,N_1091);
and U1241 (N_1241,N_1015,N_1010);
and U1242 (N_1242,N_1101,N_1159);
nor U1243 (N_1243,N_1044,N_1158);
and U1244 (N_1244,N_1061,N_1116);
nor U1245 (N_1245,N_1064,N_1054);
nand U1246 (N_1246,N_1067,N_1132);
xor U1247 (N_1247,N_1096,N_1118);
nor U1248 (N_1248,N_1014,N_1146);
xnor U1249 (N_1249,N_1076,N_1028);
and U1250 (N_1250,N_1012,N_1121);
or U1251 (N_1251,N_1169,N_1111);
xor U1252 (N_1252,N_1130,N_1153);
nand U1253 (N_1253,N_1073,N_1140);
xor U1254 (N_1254,N_1134,N_1183);
or U1255 (N_1255,N_1155,N_1185);
or U1256 (N_1256,N_1105,N_1120);
xor U1257 (N_1257,N_1008,N_1195);
and U1258 (N_1258,N_1093,N_1163);
nand U1259 (N_1259,N_1106,N_1065);
nor U1260 (N_1260,N_1164,N_1099);
nand U1261 (N_1261,N_1063,N_1038);
nand U1262 (N_1262,N_1048,N_1089);
or U1263 (N_1263,N_1162,N_1100);
or U1264 (N_1264,N_1189,N_1097);
and U1265 (N_1265,N_1046,N_1081);
and U1266 (N_1266,N_1113,N_1154);
nand U1267 (N_1267,N_1170,N_1168);
nand U1268 (N_1268,N_1027,N_1133);
nand U1269 (N_1269,N_1142,N_1129);
nor U1270 (N_1270,N_1095,N_1148);
and U1271 (N_1271,N_1119,N_1151);
or U1272 (N_1272,N_1025,N_1004);
or U1273 (N_1273,N_1047,N_1058);
nor U1274 (N_1274,N_1084,N_1055);
nand U1275 (N_1275,N_1135,N_1085);
nand U1276 (N_1276,N_1108,N_1007);
nor U1277 (N_1277,N_1102,N_1042);
nand U1278 (N_1278,N_1031,N_1175);
or U1279 (N_1279,N_1045,N_1002);
or U1280 (N_1280,N_1156,N_1009);
and U1281 (N_1281,N_1165,N_1018);
nor U1282 (N_1282,N_1041,N_1019);
xnor U1283 (N_1283,N_1184,N_1178);
and U1284 (N_1284,N_1094,N_1182);
nand U1285 (N_1285,N_1145,N_1024);
nor U1286 (N_1286,N_1137,N_1052);
nor U1287 (N_1287,N_1062,N_1176);
or U1288 (N_1288,N_1191,N_1174);
nor U1289 (N_1289,N_1161,N_1080);
or U1290 (N_1290,N_1173,N_1181);
nand U1291 (N_1291,N_1036,N_1109);
nor U1292 (N_1292,N_1013,N_1071);
nor U1293 (N_1293,N_1141,N_1187);
nor U1294 (N_1294,N_1136,N_1138);
nor U1295 (N_1295,N_1078,N_1144);
nand U1296 (N_1296,N_1026,N_1057);
nor U1297 (N_1297,N_1077,N_1092);
nor U1298 (N_1298,N_1051,N_1037);
nor U1299 (N_1299,N_1017,N_1039);
or U1300 (N_1300,N_1076,N_1037);
nand U1301 (N_1301,N_1061,N_1044);
and U1302 (N_1302,N_1024,N_1048);
nor U1303 (N_1303,N_1034,N_1048);
nor U1304 (N_1304,N_1033,N_1171);
and U1305 (N_1305,N_1142,N_1037);
or U1306 (N_1306,N_1027,N_1134);
nand U1307 (N_1307,N_1150,N_1049);
and U1308 (N_1308,N_1111,N_1070);
nand U1309 (N_1309,N_1189,N_1109);
xor U1310 (N_1310,N_1095,N_1017);
and U1311 (N_1311,N_1125,N_1178);
or U1312 (N_1312,N_1198,N_1147);
xor U1313 (N_1313,N_1173,N_1004);
nand U1314 (N_1314,N_1096,N_1106);
or U1315 (N_1315,N_1059,N_1132);
xnor U1316 (N_1316,N_1197,N_1079);
or U1317 (N_1317,N_1037,N_1001);
nand U1318 (N_1318,N_1138,N_1132);
and U1319 (N_1319,N_1073,N_1119);
nor U1320 (N_1320,N_1176,N_1087);
xor U1321 (N_1321,N_1197,N_1053);
nand U1322 (N_1322,N_1047,N_1053);
and U1323 (N_1323,N_1017,N_1076);
nand U1324 (N_1324,N_1082,N_1158);
or U1325 (N_1325,N_1032,N_1195);
nand U1326 (N_1326,N_1158,N_1118);
nand U1327 (N_1327,N_1060,N_1159);
and U1328 (N_1328,N_1116,N_1161);
xnor U1329 (N_1329,N_1063,N_1197);
or U1330 (N_1330,N_1051,N_1054);
or U1331 (N_1331,N_1173,N_1084);
nand U1332 (N_1332,N_1059,N_1146);
or U1333 (N_1333,N_1109,N_1081);
and U1334 (N_1334,N_1190,N_1178);
or U1335 (N_1335,N_1154,N_1020);
nand U1336 (N_1336,N_1176,N_1179);
nand U1337 (N_1337,N_1141,N_1135);
xnor U1338 (N_1338,N_1190,N_1033);
or U1339 (N_1339,N_1166,N_1183);
nand U1340 (N_1340,N_1115,N_1021);
or U1341 (N_1341,N_1119,N_1120);
or U1342 (N_1342,N_1179,N_1008);
nand U1343 (N_1343,N_1045,N_1173);
nor U1344 (N_1344,N_1119,N_1042);
nand U1345 (N_1345,N_1065,N_1159);
nand U1346 (N_1346,N_1155,N_1053);
xor U1347 (N_1347,N_1003,N_1102);
and U1348 (N_1348,N_1190,N_1130);
xor U1349 (N_1349,N_1174,N_1082);
and U1350 (N_1350,N_1183,N_1180);
nand U1351 (N_1351,N_1141,N_1007);
nand U1352 (N_1352,N_1050,N_1069);
and U1353 (N_1353,N_1151,N_1086);
nand U1354 (N_1354,N_1134,N_1169);
nand U1355 (N_1355,N_1051,N_1160);
and U1356 (N_1356,N_1130,N_1141);
nand U1357 (N_1357,N_1059,N_1081);
and U1358 (N_1358,N_1064,N_1055);
nand U1359 (N_1359,N_1032,N_1089);
and U1360 (N_1360,N_1097,N_1067);
nor U1361 (N_1361,N_1144,N_1069);
nand U1362 (N_1362,N_1048,N_1056);
nor U1363 (N_1363,N_1160,N_1110);
nand U1364 (N_1364,N_1106,N_1177);
and U1365 (N_1365,N_1041,N_1131);
nand U1366 (N_1366,N_1050,N_1093);
nor U1367 (N_1367,N_1041,N_1126);
nand U1368 (N_1368,N_1189,N_1131);
nand U1369 (N_1369,N_1002,N_1026);
and U1370 (N_1370,N_1127,N_1160);
and U1371 (N_1371,N_1095,N_1061);
xnor U1372 (N_1372,N_1038,N_1127);
or U1373 (N_1373,N_1045,N_1180);
xnor U1374 (N_1374,N_1069,N_1128);
nor U1375 (N_1375,N_1063,N_1163);
nand U1376 (N_1376,N_1072,N_1006);
xor U1377 (N_1377,N_1138,N_1188);
or U1378 (N_1378,N_1176,N_1112);
nor U1379 (N_1379,N_1148,N_1108);
xnor U1380 (N_1380,N_1172,N_1083);
or U1381 (N_1381,N_1080,N_1033);
and U1382 (N_1382,N_1082,N_1138);
or U1383 (N_1383,N_1161,N_1053);
or U1384 (N_1384,N_1178,N_1016);
nand U1385 (N_1385,N_1023,N_1024);
or U1386 (N_1386,N_1180,N_1039);
or U1387 (N_1387,N_1122,N_1192);
and U1388 (N_1388,N_1040,N_1076);
nand U1389 (N_1389,N_1164,N_1015);
xor U1390 (N_1390,N_1055,N_1151);
and U1391 (N_1391,N_1124,N_1051);
nor U1392 (N_1392,N_1175,N_1169);
and U1393 (N_1393,N_1142,N_1145);
or U1394 (N_1394,N_1084,N_1024);
nand U1395 (N_1395,N_1198,N_1035);
nor U1396 (N_1396,N_1097,N_1047);
nor U1397 (N_1397,N_1075,N_1107);
or U1398 (N_1398,N_1047,N_1070);
nand U1399 (N_1399,N_1084,N_1109);
nor U1400 (N_1400,N_1284,N_1393);
and U1401 (N_1401,N_1330,N_1278);
or U1402 (N_1402,N_1362,N_1229);
or U1403 (N_1403,N_1342,N_1212);
nand U1404 (N_1404,N_1301,N_1371);
or U1405 (N_1405,N_1219,N_1213);
and U1406 (N_1406,N_1261,N_1260);
or U1407 (N_1407,N_1345,N_1272);
and U1408 (N_1408,N_1200,N_1235);
or U1409 (N_1409,N_1254,N_1273);
nand U1410 (N_1410,N_1205,N_1243);
xnor U1411 (N_1411,N_1232,N_1341);
or U1412 (N_1412,N_1311,N_1337);
xor U1413 (N_1413,N_1265,N_1258);
nor U1414 (N_1414,N_1269,N_1281);
nor U1415 (N_1415,N_1223,N_1293);
nand U1416 (N_1416,N_1207,N_1359);
xnor U1417 (N_1417,N_1392,N_1233);
and U1418 (N_1418,N_1230,N_1394);
or U1419 (N_1419,N_1334,N_1307);
nand U1420 (N_1420,N_1364,N_1326);
and U1421 (N_1421,N_1288,N_1202);
or U1422 (N_1422,N_1343,N_1249);
nand U1423 (N_1423,N_1331,N_1287);
nand U1424 (N_1424,N_1375,N_1339);
nor U1425 (N_1425,N_1312,N_1216);
nand U1426 (N_1426,N_1239,N_1310);
and U1427 (N_1427,N_1351,N_1338);
or U1428 (N_1428,N_1355,N_1380);
or U1429 (N_1429,N_1237,N_1313);
or U1430 (N_1430,N_1365,N_1257);
and U1431 (N_1431,N_1327,N_1224);
xor U1432 (N_1432,N_1289,N_1305);
xor U1433 (N_1433,N_1335,N_1373);
nor U1434 (N_1434,N_1347,N_1250);
nand U1435 (N_1435,N_1302,N_1384);
xnor U1436 (N_1436,N_1298,N_1391);
or U1437 (N_1437,N_1321,N_1306);
nor U1438 (N_1438,N_1374,N_1317);
nand U1439 (N_1439,N_1352,N_1316);
and U1440 (N_1440,N_1280,N_1336);
and U1441 (N_1441,N_1304,N_1206);
or U1442 (N_1442,N_1376,N_1366);
nand U1443 (N_1443,N_1228,N_1214);
or U1444 (N_1444,N_1270,N_1299);
and U1445 (N_1445,N_1396,N_1291);
and U1446 (N_1446,N_1218,N_1294);
or U1447 (N_1447,N_1350,N_1292);
or U1448 (N_1448,N_1263,N_1262);
and U1449 (N_1449,N_1322,N_1377);
and U1450 (N_1450,N_1353,N_1357);
nor U1451 (N_1451,N_1369,N_1340);
nand U1452 (N_1452,N_1279,N_1363);
nand U1453 (N_1453,N_1325,N_1385);
or U1454 (N_1454,N_1348,N_1276);
or U1455 (N_1455,N_1389,N_1323);
and U1456 (N_1456,N_1244,N_1253);
nand U1457 (N_1457,N_1388,N_1215);
nor U1458 (N_1458,N_1381,N_1264);
nor U1459 (N_1459,N_1309,N_1277);
and U1460 (N_1460,N_1209,N_1300);
nor U1461 (N_1461,N_1295,N_1274);
nand U1462 (N_1462,N_1226,N_1259);
or U1463 (N_1463,N_1217,N_1319);
nor U1464 (N_1464,N_1231,N_1203);
and U1465 (N_1465,N_1344,N_1399);
and U1466 (N_1466,N_1296,N_1286);
nor U1467 (N_1467,N_1251,N_1329);
and U1468 (N_1468,N_1320,N_1383);
xnor U1469 (N_1469,N_1245,N_1266);
nand U1470 (N_1470,N_1246,N_1358);
nand U1471 (N_1471,N_1354,N_1248);
and U1472 (N_1472,N_1382,N_1318);
or U1473 (N_1473,N_1220,N_1387);
and U1474 (N_1474,N_1255,N_1204);
or U1475 (N_1475,N_1379,N_1314);
nand U1476 (N_1476,N_1349,N_1256);
and U1477 (N_1477,N_1290,N_1275);
nand U1478 (N_1478,N_1201,N_1395);
xnor U1479 (N_1479,N_1271,N_1333);
nor U1480 (N_1480,N_1221,N_1378);
xnor U1481 (N_1481,N_1315,N_1238);
and U1482 (N_1482,N_1283,N_1390);
or U1483 (N_1483,N_1234,N_1368);
nand U1484 (N_1484,N_1346,N_1360);
nand U1485 (N_1485,N_1208,N_1328);
nor U1486 (N_1486,N_1297,N_1247);
or U1487 (N_1487,N_1332,N_1397);
or U1488 (N_1488,N_1241,N_1225);
nor U1489 (N_1489,N_1370,N_1211);
nor U1490 (N_1490,N_1361,N_1285);
or U1491 (N_1491,N_1227,N_1386);
nor U1492 (N_1492,N_1398,N_1303);
or U1493 (N_1493,N_1252,N_1282);
nand U1494 (N_1494,N_1210,N_1240);
and U1495 (N_1495,N_1367,N_1308);
nor U1496 (N_1496,N_1268,N_1236);
or U1497 (N_1497,N_1242,N_1372);
nor U1498 (N_1498,N_1222,N_1324);
and U1499 (N_1499,N_1356,N_1267);
nor U1500 (N_1500,N_1215,N_1205);
or U1501 (N_1501,N_1344,N_1372);
or U1502 (N_1502,N_1349,N_1334);
nor U1503 (N_1503,N_1239,N_1247);
nand U1504 (N_1504,N_1338,N_1226);
nor U1505 (N_1505,N_1206,N_1381);
nand U1506 (N_1506,N_1363,N_1203);
nor U1507 (N_1507,N_1229,N_1313);
or U1508 (N_1508,N_1281,N_1237);
and U1509 (N_1509,N_1258,N_1313);
nand U1510 (N_1510,N_1224,N_1263);
or U1511 (N_1511,N_1334,N_1207);
nand U1512 (N_1512,N_1251,N_1233);
nand U1513 (N_1513,N_1322,N_1249);
nor U1514 (N_1514,N_1262,N_1221);
and U1515 (N_1515,N_1369,N_1378);
nand U1516 (N_1516,N_1301,N_1267);
and U1517 (N_1517,N_1362,N_1389);
and U1518 (N_1518,N_1389,N_1344);
and U1519 (N_1519,N_1255,N_1331);
or U1520 (N_1520,N_1395,N_1355);
nand U1521 (N_1521,N_1290,N_1243);
xnor U1522 (N_1522,N_1256,N_1278);
nor U1523 (N_1523,N_1372,N_1225);
and U1524 (N_1524,N_1288,N_1251);
nand U1525 (N_1525,N_1214,N_1371);
and U1526 (N_1526,N_1200,N_1257);
or U1527 (N_1527,N_1348,N_1377);
or U1528 (N_1528,N_1214,N_1249);
nor U1529 (N_1529,N_1305,N_1228);
nand U1530 (N_1530,N_1375,N_1228);
and U1531 (N_1531,N_1386,N_1262);
and U1532 (N_1532,N_1279,N_1340);
or U1533 (N_1533,N_1200,N_1333);
nor U1534 (N_1534,N_1324,N_1220);
or U1535 (N_1535,N_1381,N_1319);
or U1536 (N_1536,N_1365,N_1286);
and U1537 (N_1537,N_1202,N_1261);
nor U1538 (N_1538,N_1209,N_1386);
nor U1539 (N_1539,N_1243,N_1395);
nor U1540 (N_1540,N_1331,N_1397);
and U1541 (N_1541,N_1239,N_1227);
nand U1542 (N_1542,N_1290,N_1225);
nand U1543 (N_1543,N_1356,N_1374);
nand U1544 (N_1544,N_1330,N_1282);
and U1545 (N_1545,N_1295,N_1384);
nor U1546 (N_1546,N_1215,N_1234);
nor U1547 (N_1547,N_1351,N_1274);
xnor U1548 (N_1548,N_1326,N_1356);
or U1549 (N_1549,N_1305,N_1283);
nand U1550 (N_1550,N_1360,N_1285);
and U1551 (N_1551,N_1215,N_1222);
nand U1552 (N_1552,N_1270,N_1265);
or U1553 (N_1553,N_1322,N_1394);
or U1554 (N_1554,N_1237,N_1390);
and U1555 (N_1555,N_1216,N_1360);
nand U1556 (N_1556,N_1222,N_1335);
nand U1557 (N_1557,N_1300,N_1266);
or U1558 (N_1558,N_1391,N_1372);
nand U1559 (N_1559,N_1380,N_1229);
or U1560 (N_1560,N_1344,N_1313);
and U1561 (N_1561,N_1300,N_1230);
nand U1562 (N_1562,N_1243,N_1300);
xnor U1563 (N_1563,N_1263,N_1357);
and U1564 (N_1564,N_1243,N_1271);
and U1565 (N_1565,N_1237,N_1288);
or U1566 (N_1566,N_1259,N_1244);
and U1567 (N_1567,N_1243,N_1394);
nor U1568 (N_1568,N_1300,N_1320);
nand U1569 (N_1569,N_1204,N_1289);
or U1570 (N_1570,N_1346,N_1312);
nand U1571 (N_1571,N_1325,N_1262);
nor U1572 (N_1572,N_1287,N_1262);
nand U1573 (N_1573,N_1236,N_1332);
or U1574 (N_1574,N_1308,N_1240);
and U1575 (N_1575,N_1380,N_1266);
or U1576 (N_1576,N_1364,N_1362);
or U1577 (N_1577,N_1342,N_1229);
or U1578 (N_1578,N_1276,N_1308);
nand U1579 (N_1579,N_1219,N_1371);
nand U1580 (N_1580,N_1265,N_1282);
and U1581 (N_1581,N_1211,N_1337);
and U1582 (N_1582,N_1355,N_1242);
nand U1583 (N_1583,N_1342,N_1331);
nor U1584 (N_1584,N_1342,N_1287);
and U1585 (N_1585,N_1360,N_1281);
nand U1586 (N_1586,N_1236,N_1374);
xor U1587 (N_1587,N_1243,N_1227);
and U1588 (N_1588,N_1316,N_1219);
and U1589 (N_1589,N_1201,N_1210);
nand U1590 (N_1590,N_1254,N_1399);
nand U1591 (N_1591,N_1238,N_1380);
and U1592 (N_1592,N_1273,N_1256);
and U1593 (N_1593,N_1341,N_1278);
nand U1594 (N_1594,N_1270,N_1210);
xnor U1595 (N_1595,N_1293,N_1326);
and U1596 (N_1596,N_1218,N_1259);
nor U1597 (N_1597,N_1338,N_1289);
nand U1598 (N_1598,N_1247,N_1230);
and U1599 (N_1599,N_1256,N_1341);
xnor U1600 (N_1600,N_1415,N_1566);
nand U1601 (N_1601,N_1448,N_1581);
or U1602 (N_1602,N_1521,N_1432);
nor U1603 (N_1603,N_1598,N_1403);
or U1604 (N_1604,N_1429,N_1585);
nand U1605 (N_1605,N_1577,N_1594);
and U1606 (N_1606,N_1578,N_1492);
nand U1607 (N_1607,N_1590,N_1494);
and U1608 (N_1608,N_1536,N_1453);
nor U1609 (N_1609,N_1472,N_1505);
nor U1610 (N_1610,N_1484,N_1479);
or U1611 (N_1611,N_1567,N_1593);
nor U1612 (N_1612,N_1475,N_1428);
xor U1613 (N_1613,N_1512,N_1540);
nor U1614 (N_1614,N_1467,N_1431);
nand U1615 (N_1615,N_1478,N_1547);
nor U1616 (N_1616,N_1524,N_1446);
nand U1617 (N_1617,N_1460,N_1551);
nor U1618 (N_1618,N_1421,N_1586);
nor U1619 (N_1619,N_1569,N_1412);
nor U1620 (N_1620,N_1571,N_1424);
and U1621 (N_1621,N_1481,N_1499);
nand U1622 (N_1622,N_1506,N_1595);
or U1623 (N_1623,N_1400,N_1596);
nor U1624 (N_1624,N_1516,N_1497);
and U1625 (N_1625,N_1447,N_1407);
nand U1626 (N_1626,N_1565,N_1573);
nand U1627 (N_1627,N_1525,N_1477);
nand U1628 (N_1628,N_1452,N_1483);
nand U1629 (N_1629,N_1410,N_1416);
or U1630 (N_1630,N_1461,N_1473);
nand U1631 (N_1631,N_1574,N_1509);
xor U1632 (N_1632,N_1480,N_1556);
nand U1633 (N_1633,N_1425,N_1535);
nand U1634 (N_1634,N_1588,N_1559);
or U1635 (N_1635,N_1599,N_1465);
nand U1636 (N_1636,N_1557,N_1562);
nor U1637 (N_1637,N_1462,N_1463);
nand U1638 (N_1638,N_1564,N_1541);
and U1639 (N_1639,N_1532,N_1510);
nor U1640 (N_1640,N_1401,N_1458);
and U1641 (N_1641,N_1413,N_1560);
nor U1642 (N_1642,N_1518,N_1455);
or U1643 (N_1643,N_1515,N_1549);
xnor U1644 (N_1644,N_1597,N_1470);
and U1645 (N_1645,N_1522,N_1466);
xor U1646 (N_1646,N_1563,N_1539);
or U1647 (N_1647,N_1527,N_1439);
nor U1648 (N_1648,N_1482,N_1427);
and U1649 (N_1649,N_1488,N_1528);
or U1650 (N_1650,N_1406,N_1568);
nor U1651 (N_1651,N_1500,N_1529);
or U1652 (N_1652,N_1583,N_1553);
xor U1653 (N_1653,N_1434,N_1514);
or U1654 (N_1654,N_1579,N_1417);
and U1655 (N_1655,N_1454,N_1450);
nand U1656 (N_1656,N_1449,N_1423);
nand U1657 (N_1657,N_1501,N_1422);
nor U1658 (N_1658,N_1513,N_1438);
nand U1659 (N_1659,N_1493,N_1584);
and U1660 (N_1660,N_1476,N_1485);
and U1661 (N_1661,N_1420,N_1457);
nand U1662 (N_1662,N_1404,N_1440);
nand U1663 (N_1663,N_1519,N_1526);
nor U1664 (N_1664,N_1542,N_1495);
nor U1665 (N_1665,N_1570,N_1508);
or U1666 (N_1666,N_1503,N_1436);
and U1667 (N_1667,N_1437,N_1572);
nand U1668 (N_1668,N_1441,N_1402);
or U1669 (N_1669,N_1414,N_1418);
nor U1670 (N_1670,N_1486,N_1411);
nor U1671 (N_1671,N_1561,N_1546);
or U1672 (N_1672,N_1582,N_1405);
nor U1673 (N_1673,N_1534,N_1538);
or U1674 (N_1674,N_1544,N_1530);
or U1675 (N_1675,N_1443,N_1537);
nand U1676 (N_1676,N_1487,N_1444);
and U1677 (N_1677,N_1552,N_1592);
nand U1678 (N_1678,N_1451,N_1419);
or U1679 (N_1679,N_1456,N_1517);
nor U1680 (N_1680,N_1533,N_1543);
xor U1681 (N_1681,N_1511,N_1531);
nand U1682 (N_1682,N_1426,N_1445);
nor U1683 (N_1683,N_1554,N_1496);
or U1684 (N_1684,N_1468,N_1591);
nor U1685 (N_1685,N_1555,N_1489);
xor U1686 (N_1686,N_1490,N_1504);
and U1687 (N_1687,N_1575,N_1548);
and U1688 (N_1688,N_1464,N_1442);
or U1689 (N_1689,N_1545,N_1408);
or U1690 (N_1690,N_1507,N_1498);
or U1691 (N_1691,N_1502,N_1523);
nor U1692 (N_1692,N_1471,N_1469);
nor U1693 (N_1693,N_1430,N_1491);
nor U1694 (N_1694,N_1576,N_1550);
nor U1695 (N_1695,N_1520,N_1474);
nand U1696 (N_1696,N_1587,N_1409);
and U1697 (N_1697,N_1459,N_1558);
nor U1698 (N_1698,N_1580,N_1589);
or U1699 (N_1699,N_1433,N_1435);
xnor U1700 (N_1700,N_1430,N_1508);
or U1701 (N_1701,N_1598,N_1561);
xor U1702 (N_1702,N_1461,N_1553);
and U1703 (N_1703,N_1521,N_1463);
nand U1704 (N_1704,N_1555,N_1472);
nor U1705 (N_1705,N_1583,N_1595);
or U1706 (N_1706,N_1425,N_1544);
nor U1707 (N_1707,N_1426,N_1401);
or U1708 (N_1708,N_1481,N_1567);
nor U1709 (N_1709,N_1465,N_1495);
nand U1710 (N_1710,N_1532,N_1517);
or U1711 (N_1711,N_1510,N_1434);
nor U1712 (N_1712,N_1504,N_1484);
nor U1713 (N_1713,N_1492,N_1556);
nand U1714 (N_1714,N_1535,N_1507);
xnor U1715 (N_1715,N_1474,N_1442);
xor U1716 (N_1716,N_1405,N_1522);
and U1717 (N_1717,N_1466,N_1488);
nor U1718 (N_1718,N_1520,N_1551);
or U1719 (N_1719,N_1518,N_1406);
or U1720 (N_1720,N_1573,N_1523);
nand U1721 (N_1721,N_1403,N_1415);
and U1722 (N_1722,N_1508,N_1411);
or U1723 (N_1723,N_1408,N_1548);
nand U1724 (N_1724,N_1414,N_1426);
xnor U1725 (N_1725,N_1506,N_1412);
or U1726 (N_1726,N_1571,N_1583);
and U1727 (N_1727,N_1410,N_1544);
or U1728 (N_1728,N_1586,N_1557);
nand U1729 (N_1729,N_1540,N_1562);
or U1730 (N_1730,N_1560,N_1513);
nor U1731 (N_1731,N_1522,N_1592);
nor U1732 (N_1732,N_1482,N_1410);
nand U1733 (N_1733,N_1467,N_1419);
or U1734 (N_1734,N_1544,N_1523);
and U1735 (N_1735,N_1432,N_1590);
nand U1736 (N_1736,N_1426,N_1591);
nor U1737 (N_1737,N_1544,N_1568);
xor U1738 (N_1738,N_1447,N_1571);
and U1739 (N_1739,N_1462,N_1539);
nor U1740 (N_1740,N_1560,N_1519);
nor U1741 (N_1741,N_1434,N_1579);
nor U1742 (N_1742,N_1480,N_1579);
or U1743 (N_1743,N_1599,N_1536);
nor U1744 (N_1744,N_1436,N_1407);
and U1745 (N_1745,N_1475,N_1427);
and U1746 (N_1746,N_1522,N_1444);
nand U1747 (N_1747,N_1500,N_1469);
nand U1748 (N_1748,N_1560,N_1497);
xnor U1749 (N_1749,N_1513,N_1476);
and U1750 (N_1750,N_1546,N_1505);
or U1751 (N_1751,N_1471,N_1520);
nor U1752 (N_1752,N_1493,N_1596);
nor U1753 (N_1753,N_1590,N_1569);
or U1754 (N_1754,N_1594,N_1581);
nand U1755 (N_1755,N_1449,N_1427);
or U1756 (N_1756,N_1503,N_1425);
xnor U1757 (N_1757,N_1423,N_1420);
or U1758 (N_1758,N_1556,N_1456);
nor U1759 (N_1759,N_1568,N_1545);
or U1760 (N_1760,N_1400,N_1567);
or U1761 (N_1761,N_1475,N_1599);
and U1762 (N_1762,N_1424,N_1407);
nand U1763 (N_1763,N_1539,N_1416);
nor U1764 (N_1764,N_1536,N_1445);
and U1765 (N_1765,N_1473,N_1493);
nand U1766 (N_1766,N_1584,N_1503);
or U1767 (N_1767,N_1431,N_1416);
and U1768 (N_1768,N_1424,N_1455);
nor U1769 (N_1769,N_1426,N_1406);
nand U1770 (N_1770,N_1549,N_1583);
and U1771 (N_1771,N_1584,N_1408);
nand U1772 (N_1772,N_1504,N_1411);
nor U1773 (N_1773,N_1540,N_1584);
or U1774 (N_1774,N_1503,N_1489);
and U1775 (N_1775,N_1409,N_1453);
or U1776 (N_1776,N_1465,N_1502);
nand U1777 (N_1777,N_1593,N_1455);
and U1778 (N_1778,N_1582,N_1565);
nand U1779 (N_1779,N_1436,N_1505);
and U1780 (N_1780,N_1417,N_1581);
nand U1781 (N_1781,N_1488,N_1575);
nand U1782 (N_1782,N_1473,N_1537);
and U1783 (N_1783,N_1402,N_1482);
nor U1784 (N_1784,N_1583,N_1470);
nor U1785 (N_1785,N_1459,N_1417);
nand U1786 (N_1786,N_1577,N_1539);
nand U1787 (N_1787,N_1457,N_1427);
nand U1788 (N_1788,N_1514,N_1468);
or U1789 (N_1789,N_1452,N_1500);
xor U1790 (N_1790,N_1541,N_1452);
and U1791 (N_1791,N_1434,N_1580);
xor U1792 (N_1792,N_1510,N_1410);
nor U1793 (N_1793,N_1545,N_1506);
nand U1794 (N_1794,N_1470,N_1512);
or U1795 (N_1795,N_1584,N_1591);
xor U1796 (N_1796,N_1571,N_1486);
nor U1797 (N_1797,N_1457,N_1417);
nor U1798 (N_1798,N_1446,N_1409);
nand U1799 (N_1799,N_1529,N_1538);
nor U1800 (N_1800,N_1636,N_1615);
nand U1801 (N_1801,N_1698,N_1730);
xnor U1802 (N_1802,N_1640,N_1750);
or U1803 (N_1803,N_1658,N_1774);
and U1804 (N_1804,N_1650,N_1798);
nand U1805 (N_1805,N_1669,N_1675);
nor U1806 (N_1806,N_1646,N_1627);
and U1807 (N_1807,N_1696,N_1619);
xor U1808 (N_1808,N_1768,N_1771);
or U1809 (N_1809,N_1729,N_1746);
nor U1810 (N_1810,N_1783,N_1604);
and U1811 (N_1811,N_1652,N_1797);
or U1812 (N_1812,N_1602,N_1731);
and U1813 (N_1813,N_1717,N_1739);
nor U1814 (N_1814,N_1688,N_1668);
nand U1815 (N_1815,N_1787,N_1689);
and U1816 (N_1816,N_1641,N_1722);
xor U1817 (N_1817,N_1605,N_1654);
or U1818 (N_1818,N_1794,N_1721);
nand U1819 (N_1819,N_1753,N_1789);
nand U1820 (N_1820,N_1744,N_1666);
or U1821 (N_1821,N_1706,N_1611);
or U1822 (N_1822,N_1647,N_1740);
nand U1823 (N_1823,N_1610,N_1607);
nand U1824 (N_1824,N_1703,N_1694);
and U1825 (N_1825,N_1763,N_1714);
nand U1826 (N_1826,N_1649,N_1770);
nor U1827 (N_1827,N_1792,N_1758);
nand U1828 (N_1828,N_1709,N_1724);
or U1829 (N_1829,N_1712,N_1671);
nand U1830 (N_1830,N_1653,N_1651);
and U1831 (N_1831,N_1680,N_1733);
or U1832 (N_1832,N_1681,N_1795);
and U1833 (N_1833,N_1687,N_1663);
nor U1834 (N_1834,N_1626,N_1628);
xor U1835 (N_1835,N_1690,N_1677);
nand U1836 (N_1836,N_1643,N_1664);
and U1837 (N_1837,N_1685,N_1735);
or U1838 (N_1838,N_1693,N_1767);
nand U1839 (N_1839,N_1629,N_1762);
and U1840 (N_1840,N_1727,N_1618);
xor U1841 (N_1841,N_1701,N_1738);
or U1842 (N_1842,N_1655,N_1785);
or U1843 (N_1843,N_1662,N_1700);
nand U1844 (N_1844,N_1796,N_1606);
nand U1845 (N_1845,N_1632,N_1773);
nor U1846 (N_1846,N_1786,N_1782);
nand U1847 (N_1847,N_1755,N_1648);
nor U1848 (N_1848,N_1639,N_1743);
or U1849 (N_1849,N_1745,N_1665);
nand U1850 (N_1850,N_1683,N_1778);
xnor U1851 (N_1851,N_1737,N_1793);
or U1852 (N_1852,N_1631,N_1682);
nor U1853 (N_1853,N_1708,N_1761);
nand U1854 (N_1854,N_1635,N_1711);
and U1855 (N_1855,N_1766,N_1644);
nor U1856 (N_1856,N_1757,N_1634);
or U1857 (N_1857,N_1725,N_1776);
nand U1858 (N_1858,N_1678,N_1747);
nor U1859 (N_1859,N_1660,N_1601);
and U1860 (N_1860,N_1715,N_1760);
xnor U1861 (N_1861,N_1670,N_1790);
nor U1862 (N_1862,N_1764,N_1720);
or U1863 (N_1863,N_1705,N_1697);
and U1864 (N_1864,N_1719,N_1781);
nor U1865 (N_1865,N_1661,N_1765);
nor U1866 (N_1866,N_1679,N_1754);
and U1867 (N_1867,N_1630,N_1673);
or U1868 (N_1868,N_1726,N_1633);
and U1869 (N_1869,N_1617,N_1759);
and U1870 (N_1870,N_1614,N_1710);
nand U1871 (N_1871,N_1672,N_1624);
nor U1872 (N_1872,N_1613,N_1692);
or U1873 (N_1873,N_1788,N_1749);
nand U1874 (N_1874,N_1609,N_1695);
xnor U1875 (N_1875,N_1642,N_1772);
nor U1876 (N_1876,N_1718,N_1612);
and U1877 (N_1877,N_1691,N_1704);
nand U1878 (N_1878,N_1645,N_1623);
nor U1879 (N_1879,N_1622,N_1656);
and U1880 (N_1880,N_1723,N_1637);
or U1881 (N_1881,N_1676,N_1784);
nand U1882 (N_1882,N_1777,N_1752);
xnor U1883 (N_1883,N_1732,N_1608);
nor U1884 (N_1884,N_1741,N_1699);
xnor U1885 (N_1885,N_1621,N_1742);
nor U1886 (N_1886,N_1734,N_1620);
nand U1887 (N_1887,N_1603,N_1667);
nor U1888 (N_1888,N_1659,N_1799);
nand U1889 (N_1889,N_1625,N_1702);
or U1890 (N_1890,N_1716,N_1713);
nand U1891 (N_1891,N_1791,N_1779);
and U1892 (N_1892,N_1756,N_1775);
and U1893 (N_1893,N_1674,N_1686);
nand U1894 (N_1894,N_1751,N_1748);
xor U1895 (N_1895,N_1657,N_1684);
nand U1896 (N_1896,N_1638,N_1707);
xor U1897 (N_1897,N_1780,N_1769);
nor U1898 (N_1898,N_1600,N_1736);
nand U1899 (N_1899,N_1728,N_1616);
or U1900 (N_1900,N_1665,N_1644);
nand U1901 (N_1901,N_1645,N_1718);
and U1902 (N_1902,N_1626,N_1798);
nand U1903 (N_1903,N_1759,N_1697);
nand U1904 (N_1904,N_1682,N_1620);
or U1905 (N_1905,N_1734,N_1732);
nand U1906 (N_1906,N_1791,N_1710);
and U1907 (N_1907,N_1774,N_1635);
and U1908 (N_1908,N_1740,N_1790);
nand U1909 (N_1909,N_1691,N_1706);
or U1910 (N_1910,N_1712,N_1615);
nand U1911 (N_1911,N_1671,N_1686);
or U1912 (N_1912,N_1641,N_1613);
or U1913 (N_1913,N_1610,N_1677);
xor U1914 (N_1914,N_1695,N_1754);
or U1915 (N_1915,N_1673,N_1664);
and U1916 (N_1916,N_1685,N_1603);
or U1917 (N_1917,N_1715,N_1719);
nand U1918 (N_1918,N_1753,N_1738);
and U1919 (N_1919,N_1788,N_1692);
nor U1920 (N_1920,N_1602,N_1610);
nor U1921 (N_1921,N_1762,N_1747);
nor U1922 (N_1922,N_1745,N_1731);
nand U1923 (N_1923,N_1711,N_1691);
nand U1924 (N_1924,N_1744,N_1636);
nand U1925 (N_1925,N_1727,N_1785);
or U1926 (N_1926,N_1631,N_1622);
or U1927 (N_1927,N_1644,N_1648);
nor U1928 (N_1928,N_1735,N_1686);
nand U1929 (N_1929,N_1780,N_1788);
nor U1930 (N_1930,N_1794,N_1709);
or U1931 (N_1931,N_1627,N_1611);
xnor U1932 (N_1932,N_1716,N_1714);
and U1933 (N_1933,N_1733,N_1724);
nor U1934 (N_1934,N_1789,N_1710);
or U1935 (N_1935,N_1669,N_1768);
or U1936 (N_1936,N_1649,N_1641);
or U1937 (N_1937,N_1752,N_1734);
nor U1938 (N_1938,N_1625,N_1784);
xnor U1939 (N_1939,N_1704,N_1621);
nor U1940 (N_1940,N_1679,N_1734);
nand U1941 (N_1941,N_1765,N_1689);
nor U1942 (N_1942,N_1630,N_1666);
or U1943 (N_1943,N_1732,N_1621);
or U1944 (N_1944,N_1610,N_1749);
xor U1945 (N_1945,N_1738,N_1767);
nor U1946 (N_1946,N_1654,N_1609);
nor U1947 (N_1947,N_1751,N_1628);
nand U1948 (N_1948,N_1735,N_1683);
nand U1949 (N_1949,N_1705,N_1702);
nand U1950 (N_1950,N_1696,N_1793);
and U1951 (N_1951,N_1640,N_1732);
nor U1952 (N_1952,N_1668,N_1764);
xor U1953 (N_1953,N_1682,N_1689);
or U1954 (N_1954,N_1784,N_1603);
or U1955 (N_1955,N_1737,N_1684);
nand U1956 (N_1956,N_1647,N_1785);
or U1957 (N_1957,N_1730,N_1647);
and U1958 (N_1958,N_1602,N_1649);
nand U1959 (N_1959,N_1739,N_1649);
nand U1960 (N_1960,N_1669,N_1718);
xor U1961 (N_1961,N_1798,N_1743);
nor U1962 (N_1962,N_1798,N_1767);
nor U1963 (N_1963,N_1785,N_1742);
and U1964 (N_1964,N_1701,N_1730);
nor U1965 (N_1965,N_1609,N_1747);
and U1966 (N_1966,N_1732,N_1760);
or U1967 (N_1967,N_1731,N_1659);
nand U1968 (N_1968,N_1600,N_1631);
or U1969 (N_1969,N_1610,N_1628);
nor U1970 (N_1970,N_1660,N_1722);
and U1971 (N_1971,N_1755,N_1742);
nor U1972 (N_1972,N_1612,N_1621);
and U1973 (N_1973,N_1690,N_1691);
xnor U1974 (N_1974,N_1660,N_1717);
and U1975 (N_1975,N_1789,N_1762);
and U1976 (N_1976,N_1693,N_1722);
nor U1977 (N_1977,N_1777,N_1703);
xor U1978 (N_1978,N_1757,N_1734);
and U1979 (N_1979,N_1730,N_1642);
and U1980 (N_1980,N_1704,N_1719);
or U1981 (N_1981,N_1776,N_1688);
nor U1982 (N_1982,N_1700,N_1650);
and U1983 (N_1983,N_1704,N_1778);
or U1984 (N_1984,N_1674,N_1695);
nor U1985 (N_1985,N_1793,N_1678);
and U1986 (N_1986,N_1722,N_1745);
nor U1987 (N_1987,N_1725,N_1705);
nand U1988 (N_1988,N_1704,N_1684);
nor U1989 (N_1989,N_1725,N_1641);
nand U1990 (N_1990,N_1786,N_1617);
or U1991 (N_1991,N_1645,N_1717);
xnor U1992 (N_1992,N_1764,N_1644);
and U1993 (N_1993,N_1678,N_1712);
xnor U1994 (N_1994,N_1725,N_1727);
xnor U1995 (N_1995,N_1775,N_1729);
nor U1996 (N_1996,N_1602,N_1646);
and U1997 (N_1997,N_1696,N_1640);
nand U1998 (N_1998,N_1724,N_1671);
xor U1999 (N_1999,N_1790,N_1673);
xor U2000 (N_2000,N_1892,N_1891);
or U2001 (N_2001,N_1864,N_1986);
or U2002 (N_2002,N_1823,N_1981);
nand U2003 (N_2003,N_1984,N_1894);
nand U2004 (N_2004,N_1959,N_1839);
nand U2005 (N_2005,N_1968,N_1855);
xnor U2006 (N_2006,N_1869,N_1901);
and U2007 (N_2007,N_1873,N_1857);
and U2008 (N_2008,N_1938,N_1859);
or U2009 (N_2009,N_1808,N_1918);
or U2010 (N_2010,N_1896,N_1847);
nand U2011 (N_2011,N_1890,N_1899);
and U2012 (N_2012,N_1805,N_1877);
and U2013 (N_2013,N_1881,N_1867);
nand U2014 (N_2014,N_1957,N_1951);
xnor U2015 (N_2015,N_1974,N_1827);
nand U2016 (N_2016,N_1856,N_1926);
nand U2017 (N_2017,N_1841,N_1860);
nand U2018 (N_2018,N_1818,N_1935);
and U2019 (N_2019,N_1963,N_1848);
xor U2020 (N_2020,N_1943,N_1842);
nand U2021 (N_2021,N_1954,N_1939);
nor U2022 (N_2022,N_1833,N_1915);
and U2023 (N_2023,N_1948,N_1977);
and U2024 (N_2024,N_1865,N_1975);
nor U2025 (N_2025,N_1967,N_1846);
and U2026 (N_2026,N_1844,N_1940);
or U2027 (N_2027,N_1987,N_1911);
nor U2028 (N_2028,N_1962,N_1834);
or U2029 (N_2029,N_1863,N_1964);
nor U2030 (N_2030,N_1982,N_1817);
nor U2031 (N_2031,N_1988,N_1931);
and U2032 (N_2032,N_1908,N_1868);
nand U2033 (N_2033,N_1913,N_1870);
and U2034 (N_2034,N_1871,N_1999);
nand U2035 (N_2035,N_1893,N_1830);
and U2036 (N_2036,N_1858,N_1919);
or U2037 (N_2037,N_1904,N_1993);
nor U2038 (N_2038,N_1972,N_1971);
and U2039 (N_2039,N_1809,N_1946);
and U2040 (N_2040,N_1813,N_1806);
and U2041 (N_2041,N_1861,N_1875);
nand U2042 (N_2042,N_1850,N_1804);
or U2043 (N_2043,N_1980,N_1933);
xnor U2044 (N_2044,N_1945,N_1801);
nand U2045 (N_2045,N_1888,N_1955);
nor U2046 (N_2046,N_1979,N_1889);
nand U2047 (N_2047,N_1832,N_1929);
or U2048 (N_2048,N_1998,N_1900);
and U2049 (N_2049,N_1831,N_1995);
or U2050 (N_2050,N_1862,N_1851);
nand U2051 (N_2051,N_1953,N_1944);
xnor U2052 (N_2052,N_1887,N_1837);
xor U2053 (N_2053,N_1985,N_1976);
nor U2054 (N_2054,N_1897,N_1878);
and U2055 (N_2055,N_1879,N_1880);
nor U2056 (N_2056,N_1825,N_1910);
or U2057 (N_2057,N_1824,N_1973);
and U2058 (N_2058,N_1950,N_1952);
and U2059 (N_2059,N_1916,N_1895);
or U2060 (N_2060,N_1942,N_1990);
or U2061 (N_2061,N_1934,N_1958);
nor U2062 (N_2062,N_1905,N_1812);
or U2063 (N_2063,N_1961,N_1994);
nand U2064 (N_2064,N_1937,N_1883);
and U2065 (N_2065,N_1800,N_1989);
and U2066 (N_2066,N_1826,N_1969);
or U2067 (N_2067,N_1807,N_1902);
and U2068 (N_2068,N_1885,N_1996);
and U2069 (N_2069,N_1836,N_1811);
and U2070 (N_2070,N_1923,N_1936);
and U2071 (N_2071,N_1997,N_1835);
and U2072 (N_2072,N_1882,N_1909);
nand U2073 (N_2073,N_1922,N_1840);
or U2074 (N_2074,N_1898,N_1920);
nand U2075 (N_2075,N_1917,N_1843);
and U2076 (N_2076,N_1956,N_1924);
nor U2077 (N_2077,N_1970,N_1810);
and U2078 (N_2078,N_1903,N_1928);
and U2079 (N_2079,N_1838,N_1966);
or U2080 (N_2080,N_1991,N_1978);
nand U2081 (N_2081,N_1828,N_1925);
and U2082 (N_2082,N_1866,N_1907);
xnor U2083 (N_2083,N_1819,N_1965);
or U2084 (N_2084,N_1853,N_1820);
xor U2085 (N_2085,N_1992,N_1872);
nor U2086 (N_2086,N_1960,N_1884);
or U2087 (N_2087,N_1947,N_1816);
nand U2088 (N_2088,N_1921,N_1854);
nor U2089 (N_2089,N_1821,N_1932);
or U2090 (N_2090,N_1829,N_1849);
and U2091 (N_2091,N_1927,N_1802);
xor U2092 (N_2092,N_1941,N_1876);
or U2093 (N_2093,N_1930,N_1949);
nand U2094 (N_2094,N_1906,N_1914);
or U2095 (N_2095,N_1815,N_1845);
nand U2096 (N_2096,N_1886,N_1983);
and U2097 (N_2097,N_1822,N_1852);
and U2098 (N_2098,N_1803,N_1814);
nand U2099 (N_2099,N_1874,N_1912);
xor U2100 (N_2100,N_1847,N_1974);
nor U2101 (N_2101,N_1922,N_1955);
nand U2102 (N_2102,N_1890,N_1916);
and U2103 (N_2103,N_1839,N_1951);
nand U2104 (N_2104,N_1839,N_1828);
or U2105 (N_2105,N_1938,N_1856);
nand U2106 (N_2106,N_1898,N_1876);
or U2107 (N_2107,N_1963,N_1913);
or U2108 (N_2108,N_1909,N_1944);
nor U2109 (N_2109,N_1864,N_1943);
and U2110 (N_2110,N_1996,N_1918);
and U2111 (N_2111,N_1995,N_1815);
or U2112 (N_2112,N_1828,N_1998);
nor U2113 (N_2113,N_1848,N_1870);
xor U2114 (N_2114,N_1866,N_1947);
nand U2115 (N_2115,N_1958,N_1904);
or U2116 (N_2116,N_1837,N_1903);
nand U2117 (N_2117,N_1812,N_1981);
xor U2118 (N_2118,N_1834,N_1976);
nor U2119 (N_2119,N_1838,N_1926);
or U2120 (N_2120,N_1888,N_1861);
or U2121 (N_2121,N_1864,N_1958);
and U2122 (N_2122,N_1909,N_1884);
or U2123 (N_2123,N_1899,N_1915);
xor U2124 (N_2124,N_1908,N_1861);
nand U2125 (N_2125,N_1925,N_1889);
or U2126 (N_2126,N_1820,N_1999);
or U2127 (N_2127,N_1973,N_1858);
nor U2128 (N_2128,N_1885,N_1868);
or U2129 (N_2129,N_1979,N_1996);
or U2130 (N_2130,N_1825,N_1960);
nor U2131 (N_2131,N_1980,N_1948);
nand U2132 (N_2132,N_1800,N_1841);
nor U2133 (N_2133,N_1992,N_1837);
nor U2134 (N_2134,N_1862,N_1896);
nand U2135 (N_2135,N_1935,N_1888);
nor U2136 (N_2136,N_1884,N_1875);
or U2137 (N_2137,N_1855,N_1905);
nand U2138 (N_2138,N_1910,N_1962);
nor U2139 (N_2139,N_1967,N_1886);
nor U2140 (N_2140,N_1905,N_1955);
and U2141 (N_2141,N_1860,N_1975);
nor U2142 (N_2142,N_1902,N_1899);
or U2143 (N_2143,N_1830,N_1983);
nand U2144 (N_2144,N_1874,N_1867);
and U2145 (N_2145,N_1898,N_1932);
xor U2146 (N_2146,N_1844,N_1961);
nor U2147 (N_2147,N_1802,N_1877);
nor U2148 (N_2148,N_1875,N_1822);
nand U2149 (N_2149,N_1846,N_1916);
nor U2150 (N_2150,N_1875,N_1831);
and U2151 (N_2151,N_1944,N_1880);
nor U2152 (N_2152,N_1900,N_1971);
nor U2153 (N_2153,N_1847,N_1841);
nor U2154 (N_2154,N_1961,N_1900);
nor U2155 (N_2155,N_1989,N_1889);
and U2156 (N_2156,N_1933,N_1916);
or U2157 (N_2157,N_1981,N_1845);
or U2158 (N_2158,N_1878,N_1970);
xnor U2159 (N_2159,N_1919,N_1812);
nor U2160 (N_2160,N_1875,N_1956);
and U2161 (N_2161,N_1851,N_1938);
and U2162 (N_2162,N_1952,N_1858);
or U2163 (N_2163,N_1974,N_1888);
or U2164 (N_2164,N_1911,N_1812);
or U2165 (N_2165,N_1988,N_1930);
nand U2166 (N_2166,N_1815,N_1890);
nor U2167 (N_2167,N_1870,N_1861);
nor U2168 (N_2168,N_1841,N_1975);
xor U2169 (N_2169,N_1825,N_1913);
nand U2170 (N_2170,N_1867,N_1824);
nand U2171 (N_2171,N_1984,N_1862);
nand U2172 (N_2172,N_1960,N_1942);
or U2173 (N_2173,N_1952,N_1879);
nor U2174 (N_2174,N_1906,N_1922);
nor U2175 (N_2175,N_1879,N_1956);
or U2176 (N_2176,N_1822,N_1906);
or U2177 (N_2177,N_1814,N_1950);
and U2178 (N_2178,N_1815,N_1941);
nor U2179 (N_2179,N_1880,N_1923);
xor U2180 (N_2180,N_1972,N_1880);
nor U2181 (N_2181,N_1892,N_1831);
or U2182 (N_2182,N_1820,N_1921);
or U2183 (N_2183,N_1834,N_1961);
xor U2184 (N_2184,N_1971,N_1922);
nor U2185 (N_2185,N_1968,N_1865);
xor U2186 (N_2186,N_1806,N_1868);
nor U2187 (N_2187,N_1838,N_1882);
or U2188 (N_2188,N_1919,N_1962);
or U2189 (N_2189,N_1864,N_1920);
xnor U2190 (N_2190,N_1865,N_1801);
or U2191 (N_2191,N_1828,N_1898);
and U2192 (N_2192,N_1951,N_1845);
nor U2193 (N_2193,N_1865,N_1870);
nand U2194 (N_2194,N_1934,N_1863);
and U2195 (N_2195,N_1903,N_1888);
nor U2196 (N_2196,N_1813,N_1814);
nand U2197 (N_2197,N_1886,N_1966);
xnor U2198 (N_2198,N_1828,N_1819);
nand U2199 (N_2199,N_1898,N_1979);
xor U2200 (N_2200,N_2111,N_2020);
nand U2201 (N_2201,N_2096,N_2191);
nor U2202 (N_2202,N_2144,N_2147);
and U2203 (N_2203,N_2161,N_2124);
or U2204 (N_2204,N_2092,N_2066);
nor U2205 (N_2205,N_2070,N_2118);
or U2206 (N_2206,N_2018,N_2047);
nand U2207 (N_2207,N_2159,N_2175);
nand U2208 (N_2208,N_2028,N_2164);
nor U2209 (N_2209,N_2157,N_2193);
nor U2210 (N_2210,N_2142,N_2171);
nor U2211 (N_2211,N_2100,N_2052);
xnor U2212 (N_2212,N_2044,N_2071);
or U2213 (N_2213,N_2005,N_2058);
nor U2214 (N_2214,N_2065,N_2141);
nand U2215 (N_2215,N_2126,N_2059);
nand U2216 (N_2216,N_2021,N_2120);
and U2217 (N_2217,N_2080,N_2112);
nand U2218 (N_2218,N_2033,N_2117);
or U2219 (N_2219,N_2133,N_2131);
xnor U2220 (N_2220,N_2069,N_2031);
and U2221 (N_2221,N_2034,N_2169);
nand U2222 (N_2222,N_2048,N_2087);
or U2223 (N_2223,N_2167,N_2097);
xor U2224 (N_2224,N_2160,N_2003);
or U2225 (N_2225,N_2168,N_2061);
nor U2226 (N_2226,N_2158,N_2057);
nand U2227 (N_2227,N_2180,N_2105);
xnor U2228 (N_2228,N_2125,N_2053);
xor U2229 (N_2229,N_2068,N_2104);
xnor U2230 (N_2230,N_2074,N_2001);
and U2231 (N_2231,N_2049,N_2063);
or U2232 (N_2232,N_2054,N_2011);
nand U2233 (N_2233,N_2146,N_2010);
xnor U2234 (N_2234,N_2132,N_2006);
or U2235 (N_2235,N_2002,N_2121);
or U2236 (N_2236,N_2152,N_2185);
nor U2237 (N_2237,N_2076,N_2007);
nor U2238 (N_2238,N_2036,N_2148);
xor U2239 (N_2239,N_2172,N_2198);
or U2240 (N_2240,N_2176,N_2182);
nor U2241 (N_2241,N_2122,N_2025);
or U2242 (N_2242,N_2149,N_2012);
nand U2243 (N_2243,N_2064,N_2109);
nor U2244 (N_2244,N_2199,N_2127);
and U2245 (N_2245,N_2027,N_2186);
nor U2246 (N_2246,N_2178,N_2195);
or U2247 (N_2247,N_2155,N_2107);
and U2248 (N_2248,N_2079,N_2123);
xnor U2249 (N_2249,N_2009,N_2136);
xnor U2250 (N_2250,N_2140,N_2017);
nand U2251 (N_2251,N_2015,N_2154);
xor U2252 (N_2252,N_2040,N_2098);
or U2253 (N_2253,N_2077,N_2162);
and U2254 (N_2254,N_2137,N_2099);
and U2255 (N_2255,N_2151,N_2103);
xor U2256 (N_2256,N_2037,N_2114);
and U2257 (N_2257,N_2170,N_2026);
nor U2258 (N_2258,N_2073,N_2110);
xor U2259 (N_2259,N_2188,N_2115);
and U2260 (N_2260,N_2039,N_2116);
and U2261 (N_2261,N_2041,N_2085);
and U2262 (N_2262,N_2135,N_2050);
and U2263 (N_2263,N_2067,N_2043);
or U2264 (N_2264,N_2177,N_2045);
xnor U2265 (N_2265,N_2084,N_2106);
and U2266 (N_2266,N_2101,N_2143);
and U2267 (N_2267,N_2089,N_2090);
nand U2268 (N_2268,N_2163,N_2086);
and U2269 (N_2269,N_2187,N_2094);
nor U2270 (N_2270,N_2016,N_2183);
nor U2271 (N_2271,N_2023,N_2032);
nand U2272 (N_2272,N_2189,N_2075);
nor U2273 (N_2273,N_2156,N_2093);
and U2274 (N_2274,N_2165,N_2000);
nor U2275 (N_2275,N_2130,N_2102);
nand U2276 (N_2276,N_2129,N_2174);
nor U2277 (N_2277,N_2197,N_2072);
and U2278 (N_2278,N_2091,N_2056);
nor U2279 (N_2279,N_2166,N_2008);
nor U2280 (N_2280,N_2095,N_2153);
or U2281 (N_2281,N_2030,N_2194);
or U2282 (N_2282,N_2024,N_2035);
or U2283 (N_2283,N_2108,N_2150);
or U2284 (N_2284,N_2134,N_2013);
or U2285 (N_2285,N_2029,N_2062);
and U2286 (N_2286,N_2055,N_2060);
or U2287 (N_2287,N_2083,N_2192);
or U2288 (N_2288,N_2004,N_2138);
and U2289 (N_2289,N_2081,N_2088);
or U2290 (N_2290,N_2139,N_2022);
and U2291 (N_2291,N_2113,N_2046);
or U2292 (N_2292,N_2014,N_2051);
and U2293 (N_2293,N_2082,N_2019);
nand U2294 (N_2294,N_2042,N_2184);
nor U2295 (N_2295,N_2119,N_2078);
or U2296 (N_2296,N_2190,N_2173);
nor U2297 (N_2297,N_2038,N_2181);
nor U2298 (N_2298,N_2196,N_2128);
or U2299 (N_2299,N_2179,N_2145);
nand U2300 (N_2300,N_2097,N_2129);
nor U2301 (N_2301,N_2180,N_2032);
nor U2302 (N_2302,N_2028,N_2085);
nor U2303 (N_2303,N_2191,N_2098);
and U2304 (N_2304,N_2043,N_2127);
and U2305 (N_2305,N_2170,N_2081);
xnor U2306 (N_2306,N_2037,N_2029);
and U2307 (N_2307,N_2091,N_2173);
nor U2308 (N_2308,N_2113,N_2021);
and U2309 (N_2309,N_2183,N_2118);
and U2310 (N_2310,N_2101,N_2104);
and U2311 (N_2311,N_2162,N_2025);
or U2312 (N_2312,N_2010,N_2074);
nand U2313 (N_2313,N_2117,N_2140);
or U2314 (N_2314,N_2013,N_2067);
nand U2315 (N_2315,N_2114,N_2143);
nor U2316 (N_2316,N_2020,N_2078);
nor U2317 (N_2317,N_2110,N_2039);
and U2318 (N_2318,N_2148,N_2129);
and U2319 (N_2319,N_2000,N_2176);
nand U2320 (N_2320,N_2117,N_2162);
or U2321 (N_2321,N_2142,N_2114);
or U2322 (N_2322,N_2005,N_2167);
nand U2323 (N_2323,N_2033,N_2066);
and U2324 (N_2324,N_2166,N_2061);
and U2325 (N_2325,N_2112,N_2142);
nand U2326 (N_2326,N_2069,N_2147);
or U2327 (N_2327,N_2006,N_2119);
nor U2328 (N_2328,N_2082,N_2124);
nor U2329 (N_2329,N_2118,N_2150);
or U2330 (N_2330,N_2054,N_2052);
or U2331 (N_2331,N_2105,N_2163);
xor U2332 (N_2332,N_2014,N_2137);
nor U2333 (N_2333,N_2152,N_2024);
xnor U2334 (N_2334,N_2162,N_2002);
nand U2335 (N_2335,N_2108,N_2104);
and U2336 (N_2336,N_2178,N_2061);
nor U2337 (N_2337,N_2076,N_2017);
nand U2338 (N_2338,N_2098,N_2065);
xor U2339 (N_2339,N_2164,N_2034);
nor U2340 (N_2340,N_2016,N_2123);
nor U2341 (N_2341,N_2169,N_2029);
xnor U2342 (N_2342,N_2027,N_2070);
nor U2343 (N_2343,N_2185,N_2170);
and U2344 (N_2344,N_2105,N_2123);
nor U2345 (N_2345,N_2097,N_2073);
and U2346 (N_2346,N_2101,N_2005);
nor U2347 (N_2347,N_2048,N_2160);
xor U2348 (N_2348,N_2170,N_2028);
nand U2349 (N_2349,N_2161,N_2018);
or U2350 (N_2350,N_2004,N_2016);
xor U2351 (N_2351,N_2086,N_2074);
and U2352 (N_2352,N_2017,N_2130);
nand U2353 (N_2353,N_2082,N_2003);
and U2354 (N_2354,N_2051,N_2019);
and U2355 (N_2355,N_2020,N_2192);
nand U2356 (N_2356,N_2015,N_2080);
nor U2357 (N_2357,N_2048,N_2190);
or U2358 (N_2358,N_2001,N_2014);
nand U2359 (N_2359,N_2154,N_2125);
or U2360 (N_2360,N_2066,N_2071);
nor U2361 (N_2361,N_2040,N_2049);
xnor U2362 (N_2362,N_2018,N_2088);
xnor U2363 (N_2363,N_2051,N_2122);
nor U2364 (N_2364,N_2049,N_2095);
and U2365 (N_2365,N_2029,N_2110);
nor U2366 (N_2366,N_2093,N_2110);
xnor U2367 (N_2367,N_2108,N_2014);
nor U2368 (N_2368,N_2130,N_2103);
and U2369 (N_2369,N_2199,N_2075);
or U2370 (N_2370,N_2167,N_2028);
or U2371 (N_2371,N_2097,N_2104);
nor U2372 (N_2372,N_2056,N_2075);
and U2373 (N_2373,N_2159,N_2099);
xnor U2374 (N_2374,N_2134,N_2077);
nand U2375 (N_2375,N_2073,N_2185);
or U2376 (N_2376,N_2195,N_2086);
or U2377 (N_2377,N_2051,N_2054);
xor U2378 (N_2378,N_2152,N_2097);
nor U2379 (N_2379,N_2142,N_2199);
nand U2380 (N_2380,N_2040,N_2001);
nor U2381 (N_2381,N_2159,N_2084);
and U2382 (N_2382,N_2110,N_2143);
or U2383 (N_2383,N_2062,N_2184);
nor U2384 (N_2384,N_2019,N_2040);
and U2385 (N_2385,N_2034,N_2041);
and U2386 (N_2386,N_2132,N_2070);
nand U2387 (N_2387,N_2175,N_2097);
nand U2388 (N_2388,N_2003,N_2072);
xnor U2389 (N_2389,N_2101,N_2096);
nor U2390 (N_2390,N_2023,N_2148);
or U2391 (N_2391,N_2141,N_2187);
xor U2392 (N_2392,N_2033,N_2195);
and U2393 (N_2393,N_2143,N_2009);
and U2394 (N_2394,N_2161,N_2055);
nand U2395 (N_2395,N_2023,N_2104);
and U2396 (N_2396,N_2084,N_2104);
and U2397 (N_2397,N_2143,N_2058);
xor U2398 (N_2398,N_2102,N_2007);
or U2399 (N_2399,N_2058,N_2029);
xor U2400 (N_2400,N_2335,N_2386);
and U2401 (N_2401,N_2297,N_2204);
or U2402 (N_2402,N_2242,N_2228);
nand U2403 (N_2403,N_2232,N_2203);
or U2404 (N_2404,N_2276,N_2226);
and U2405 (N_2405,N_2362,N_2284);
nor U2406 (N_2406,N_2272,N_2270);
xor U2407 (N_2407,N_2225,N_2283);
or U2408 (N_2408,N_2248,N_2239);
or U2409 (N_2409,N_2332,N_2217);
xnor U2410 (N_2410,N_2287,N_2398);
nand U2411 (N_2411,N_2372,N_2329);
nand U2412 (N_2412,N_2383,N_2392);
nand U2413 (N_2413,N_2236,N_2300);
or U2414 (N_2414,N_2299,N_2359);
nand U2415 (N_2415,N_2351,N_2364);
nand U2416 (N_2416,N_2349,N_2258);
and U2417 (N_2417,N_2315,N_2215);
nand U2418 (N_2418,N_2245,N_2288);
nor U2419 (N_2419,N_2353,N_2265);
or U2420 (N_2420,N_2330,N_2393);
and U2421 (N_2421,N_2388,N_2323);
and U2422 (N_2422,N_2354,N_2379);
nor U2423 (N_2423,N_2210,N_2326);
nor U2424 (N_2424,N_2396,N_2333);
and U2425 (N_2425,N_2279,N_2244);
xor U2426 (N_2426,N_2376,N_2338);
nand U2427 (N_2427,N_2325,N_2294);
nor U2428 (N_2428,N_2373,N_2307);
and U2429 (N_2429,N_2221,N_2316);
and U2430 (N_2430,N_2317,N_2296);
and U2431 (N_2431,N_2319,N_2394);
nand U2432 (N_2432,N_2247,N_2304);
or U2433 (N_2433,N_2237,N_2397);
nor U2434 (N_2434,N_2200,N_2266);
nor U2435 (N_2435,N_2292,N_2262);
nor U2436 (N_2436,N_2229,N_2365);
and U2437 (N_2437,N_2253,N_2213);
nand U2438 (N_2438,N_2259,N_2395);
or U2439 (N_2439,N_2233,N_2309);
or U2440 (N_2440,N_2336,N_2263);
nand U2441 (N_2441,N_2337,N_2235);
nand U2442 (N_2442,N_2243,N_2305);
nor U2443 (N_2443,N_2391,N_2231);
nor U2444 (N_2444,N_2306,N_2381);
nand U2445 (N_2445,N_2352,N_2238);
and U2446 (N_2446,N_2252,N_2343);
nand U2447 (N_2447,N_2342,N_2251);
xor U2448 (N_2448,N_2312,N_2291);
nor U2449 (N_2449,N_2360,N_2254);
and U2450 (N_2450,N_2348,N_2334);
nor U2451 (N_2451,N_2216,N_2261);
or U2452 (N_2452,N_2240,N_2387);
and U2453 (N_2453,N_2267,N_2209);
nand U2454 (N_2454,N_2370,N_2285);
nor U2455 (N_2455,N_2281,N_2399);
nand U2456 (N_2456,N_2246,N_2212);
nand U2457 (N_2457,N_2314,N_2311);
and U2458 (N_2458,N_2382,N_2369);
or U2459 (N_2459,N_2222,N_2277);
xnor U2460 (N_2460,N_2289,N_2389);
and U2461 (N_2461,N_2385,N_2241);
and U2462 (N_2462,N_2218,N_2282);
and U2463 (N_2463,N_2271,N_2341);
or U2464 (N_2464,N_2380,N_2250);
nor U2465 (N_2465,N_2224,N_2278);
nor U2466 (N_2466,N_2350,N_2327);
nand U2467 (N_2467,N_2206,N_2374);
or U2468 (N_2468,N_2301,N_2331);
xor U2469 (N_2469,N_2205,N_2310);
or U2470 (N_2470,N_2269,N_2275);
xnor U2471 (N_2471,N_2356,N_2303);
nor U2472 (N_2472,N_2290,N_2227);
nand U2473 (N_2473,N_2346,N_2207);
or U2474 (N_2474,N_2390,N_2220);
or U2475 (N_2475,N_2286,N_2321);
and U2476 (N_2476,N_2223,N_2367);
nand U2477 (N_2477,N_2230,N_2320);
nand U2478 (N_2478,N_2219,N_2366);
and U2479 (N_2479,N_2249,N_2308);
nor U2480 (N_2480,N_2344,N_2322);
and U2481 (N_2481,N_2328,N_2256);
and U2482 (N_2482,N_2313,N_2280);
xor U2483 (N_2483,N_2201,N_2273);
nor U2484 (N_2484,N_2260,N_2255);
xnor U2485 (N_2485,N_2264,N_2345);
nor U2486 (N_2486,N_2324,N_2268);
xnor U2487 (N_2487,N_2368,N_2384);
nor U2488 (N_2488,N_2340,N_2363);
and U2489 (N_2489,N_2318,N_2361);
nor U2490 (N_2490,N_2234,N_2357);
and U2491 (N_2491,N_2371,N_2375);
nor U2492 (N_2492,N_2358,N_2211);
nor U2493 (N_2493,N_2208,N_2202);
or U2494 (N_2494,N_2274,N_2295);
nand U2495 (N_2495,N_2302,N_2339);
and U2496 (N_2496,N_2355,N_2257);
nor U2497 (N_2497,N_2214,N_2293);
xnor U2498 (N_2498,N_2378,N_2347);
nor U2499 (N_2499,N_2298,N_2377);
and U2500 (N_2500,N_2293,N_2291);
and U2501 (N_2501,N_2219,N_2213);
nor U2502 (N_2502,N_2205,N_2254);
and U2503 (N_2503,N_2262,N_2388);
xor U2504 (N_2504,N_2368,N_2238);
or U2505 (N_2505,N_2324,N_2206);
xnor U2506 (N_2506,N_2213,N_2209);
or U2507 (N_2507,N_2397,N_2384);
or U2508 (N_2508,N_2384,N_2381);
or U2509 (N_2509,N_2310,N_2234);
nor U2510 (N_2510,N_2222,N_2200);
nor U2511 (N_2511,N_2336,N_2201);
or U2512 (N_2512,N_2222,N_2284);
xnor U2513 (N_2513,N_2215,N_2382);
nand U2514 (N_2514,N_2389,N_2255);
or U2515 (N_2515,N_2391,N_2344);
nor U2516 (N_2516,N_2273,N_2277);
and U2517 (N_2517,N_2230,N_2378);
and U2518 (N_2518,N_2245,N_2231);
or U2519 (N_2519,N_2241,N_2376);
nor U2520 (N_2520,N_2331,N_2232);
nand U2521 (N_2521,N_2254,N_2346);
or U2522 (N_2522,N_2312,N_2263);
or U2523 (N_2523,N_2353,N_2234);
or U2524 (N_2524,N_2253,N_2216);
or U2525 (N_2525,N_2298,N_2371);
and U2526 (N_2526,N_2302,N_2353);
nor U2527 (N_2527,N_2231,N_2368);
nand U2528 (N_2528,N_2322,N_2279);
xnor U2529 (N_2529,N_2204,N_2246);
nor U2530 (N_2530,N_2222,N_2308);
nand U2531 (N_2531,N_2230,N_2392);
or U2532 (N_2532,N_2304,N_2290);
nand U2533 (N_2533,N_2226,N_2321);
nand U2534 (N_2534,N_2204,N_2260);
nor U2535 (N_2535,N_2333,N_2253);
or U2536 (N_2536,N_2374,N_2373);
nor U2537 (N_2537,N_2281,N_2355);
nand U2538 (N_2538,N_2291,N_2204);
nand U2539 (N_2539,N_2226,N_2328);
and U2540 (N_2540,N_2293,N_2346);
and U2541 (N_2541,N_2202,N_2266);
or U2542 (N_2542,N_2243,N_2379);
or U2543 (N_2543,N_2298,N_2287);
nor U2544 (N_2544,N_2235,N_2206);
and U2545 (N_2545,N_2253,N_2222);
or U2546 (N_2546,N_2393,N_2378);
nor U2547 (N_2547,N_2228,N_2269);
or U2548 (N_2548,N_2361,N_2236);
xor U2549 (N_2549,N_2306,N_2347);
nand U2550 (N_2550,N_2378,N_2308);
and U2551 (N_2551,N_2324,N_2211);
and U2552 (N_2552,N_2395,N_2231);
and U2553 (N_2553,N_2219,N_2301);
or U2554 (N_2554,N_2360,N_2363);
nand U2555 (N_2555,N_2291,N_2250);
or U2556 (N_2556,N_2347,N_2248);
nor U2557 (N_2557,N_2212,N_2201);
and U2558 (N_2558,N_2322,N_2352);
or U2559 (N_2559,N_2208,N_2365);
nor U2560 (N_2560,N_2370,N_2353);
nand U2561 (N_2561,N_2345,N_2214);
nand U2562 (N_2562,N_2228,N_2258);
nand U2563 (N_2563,N_2329,N_2360);
nor U2564 (N_2564,N_2311,N_2392);
or U2565 (N_2565,N_2334,N_2257);
and U2566 (N_2566,N_2221,N_2398);
nand U2567 (N_2567,N_2393,N_2284);
and U2568 (N_2568,N_2348,N_2270);
nand U2569 (N_2569,N_2306,N_2271);
nand U2570 (N_2570,N_2343,N_2242);
nand U2571 (N_2571,N_2253,N_2311);
and U2572 (N_2572,N_2330,N_2357);
nor U2573 (N_2573,N_2353,N_2352);
and U2574 (N_2574,N_2269,N_2285);
nor U2575 (N_2575,N_2396,N_2324);
xor U2576 (N_2576,N_2373,N_2277);
nor U2577 (N_2577,N_2319,N_2284);
xor U2578 (N_2578,N_2255,N_2354);
nor U2579 (N_2579,N_2229,N_2210);
nor U2580 (N_2580,N_2311,N_2324);
and U2581 (N_2581,N_2374,N_2377);
and U2582 (N_2582,N_2278,N_2389);
or U2583 (N_2583,N_2370,N_2343);
or U2584 (N_2584,N_2247,N_2220);
xor U2585 (N_2585,N_2249,N_2299);
nor U2586 (N_2586,N_2312,N_2389);
or U2587 (N_2587,N_2366,N_2308);
and U2588 (N_2588,N_2308,N_2332);
and U2589 (N_2589,N_2376,N_2213);
or U2590 (N_2590,N_2399,N_2218);
xor U2591 (N_2591,N_2379,N_2302);
xor U2592 (N_2592,N_2246,N_2399);
nor U2593 (N_2593,N_2383,N_2342);
nand U2594 (N_2594,N_2370,N_2388);
and U2595 (N_2595,N_2301,N_2385);
nor U2596 (N_2596,N_2257,N_2396);
and U2597 (N_2597,N_2247,N_2319);
and U2598 (N_2598,N_2216,N_2316);
nor U2599 (N_2599,N_2271,N_2244);
nand U2600 (N_2600,N_2426,N_2477);
xor U2601 (N_2601,N_2468,N_2476);
nand U2602 (N_2602,N_2566,N_2595);
nand U2603 (N_2603,N_2444,N_2584);
and U2604 (N_2604,N_2434,N_2545);
nand U2605 (N_2605,N_2553,N_2464);
or U2606 (N_2606,N_2417,N_2556);
or U2607 (N_2607,N_2461,N_2500);
or U2608 (N_2608,N_2586,N_2403);
and U2609 (N_2609,N_2501,N_2537);
nand U2610 (N_2610,N_2546,N_2448);
nor U2611 (N_2611,N_2587,N_2543);
xnor U2612 (N_2612,N_2446,N_2588);
or U2613 (N_2613,N_2466,N_2410);
xor U2614 (N_2614,N_2591,N_2491);
nor U2615 (N_2615,N_2521,N_2436);
and U2616 (N_2616,N_2408,N_2452);
and U2617 (N_2617,N_2506,N_2547);
xor U2618 (N_2618,N_2516,N_2442);
or U2619 (N_2619,N_2401,N_2526);
xnor U2620 (N_2620,N_2599,N_2480);
nand U2621 (N_2621,N_2593,N_2435);
or U2622 (N_2622,N_2421,N_2441);
and U2623 (N_2623,N_2459,N_2525);
and U2624 (N_2624,N_2535,N_2503);
and U2625 (N_2625,N_2419,N_2530);
or U2626 (N_2626,N_2457,N_2504);
nand U2627 (N_2627,N_2469,N_2576);
nor U2628 (N_2628,N_2559,N_2416);
and U2629 (N_2629,N_2458,N_2578);
nor U2630 (N_2630,N_2497,N_2422);
xor U2631 (N_2631,N_2524,N_2598);
and U2632 (N_2632,N_2437,N_2523);
nor U2633 (N_2633,N_2567,N_2470);
nor U2634 (N_2634,N_2423,N_2445);
and U2635 (N_2635,N_2509,N_2471);
or U2636 (N_2636,N_2558,N_2564);
nor U2637 (N_2637,N_2433,N_2590);
nor U2638 (N_2638,N_2571,N_2494);
or U2639 (N_2639,N_2549,N_2453);
nor U2640 (N_2640,N_2573,N_2498);
and U2641 (N_2641,N_2431,N_2438);
and U2642 (N_2642,N_2511,N_2552);
nor U2643 (N_2643,N_2542,N_2551);
and U2644 (N_2644,N_2577,N_2548);
or U2645 (N_2645,N_2574,N_2518);
nor U2646 (N_2646,N_2589,N_2413);
nor U2647 (N_2647,N_2505,N_2414);
or U2648 (N_2648,N_2429,N_2432);
or U2649 (N_2649,N_2405,N_2527);
nor U2650 (N_2650,N_2463,N_2534);
or U2651 (N_2651,N_2490,N_2406);
xnor U2652 (N_2652,N_2579,N_2596);
nor U2653 (N_2653,N_2541,N_2404);
nor U2654 (N_2654,N_2424,N_2447);
xnor U2655 (N_2655,N_2495,N_2594);
or U2656 (N_2656,N_2455,N_2568);
nand U2657 (N_2657,N_2532,N_2473);
nand U2658 (N_2658,N_2415,N_2462);
and U2659 (N_2659,N_2488,N_2507);
nor U2660 (N_2660,N_2440,N_2485);
or U2661 (N_2661,N_2557,N_2533);
nor U2662 (N_2662,N_2544,N_2418);
and U2663 (N_2663,N_2560,N_2474);
and U2664 (N_2664,N_2597,N_2402);
or U2665 (N_2665,N_2478,N_2540);
nor U2666 (N_2666,N_2420,N_2565);
and U2667 (N_2667,N_2483,N_2430);
nor U2668 (N_2668,N_2427,N_2450);
nor U2669 (N_2669,N_2492,N_2502);
or U2670 (N_2670,N_2515,N_2467);
and U2671 (N_2671,N_2449,N_2465);
nand U2672 (N_2672,N_2569,N_2531);
and U2673 (N_2673,N_2489,N_2487);
or U2674 (N_2674,N_2400,N_2513);
nand U2675 (N_2675,N_2562,N_2451);
and U2676 (N_2676,N_2561,N_2512);
and U2677 (N_2677,N_2536,N_2425);
nor U2678 (N_2678,N_2570,N_2580);
or U2679 (N_2679,N_2412,N_2479);
nor U2680 (N_2680,N_2439,N_2575);
and U2681 (N_2681,N_2428,N_2529);
nand U2682 (N_2682,N_2517,N_2550);
xor U2683 (N_2683,N_2522,N_2481);
xor U2684 (N_2684,N_2499,N_2592);
nand U2685 (N_2685,N_2409,N_2475);
nand U2686 (N_2686,N_2496,N_2538);
nand U2687 (N_2687,N_2407,N_2555);
and U2688 (N_2688,N_2472,N_2484);
nor U2689 (N_2689,N_2508,N_2482);
and U2690 (N_2690,N_2528,N_2510);
nand U2691 (N_2691,N_2581,N_2454);
nand U2692 (N_2692,N_2520,N_2554);
and U2693 (N_2693,N_2460,N_2539);
or U2694 (N_2694,N_2585,N_2486);
and U2695 (N_2695,N_2582,N_2563);
and U2696 (N_2696,N_2456,N_2572);
and U2697 (N_2697,N_2583,N_2493);
nor U2698 (N_2698,N_2514,N_2519);
or U2699 (N_2699,N_2443,N_2411);
nor U2700 (N_2700,N_2558,N_2576);
nor U2701 (N_2701,N_2428,N_2473);
nand U2702 (N_2702,N_2487,N_2571);
nor U2703 (N_2703,N_2558,N_2579);
xor U2704 (N_2704,N_2520,N_2532);
or U2705 (N_2705,N_2580,N_2520);
and U2706 (N_2706,N_2464,N_2425);
and U2707 (N_2707,N_2522,N_2447);
nor U2708 (N_2708,N_2407,N_2496);
or U2709 (N_2709,N_2517,N_2443);
and U2710 (N_2710,N_2514,N_2536);
nand U2711 (N_2711,N_2552,N_2591);
nor U2712 (N_2712,N_2420,N_2417);
and U2713 (N_2713,N_2546,N_2592);
and U2714 (N_2714,N_2499,N_2522);
and U2715 (N_2715,N_2506,N_2443);
xor U2716 (N_2716,N_2515,N_2541);
nor U2717 (N_2717,N_2425,N_2549);
nand U2718 (N_2718,N_2430,N_2522);
and U2719 (N_2719,N_2494,N_2411);
nand U2720 (N_2720,N_2430,N_2472);
and U2721 (N_2721,N_2474,N_2489);
or U2722 (N_2722,N_2439,N_2527);
nand U2723 (N_2723,N_2476,N_2477);
and U2724 (N_2724,N_2424,N_2453);
nand U2725 (N_2725,N_2453,N_2586);
nand U2726 (N_2726,N_2466,N_2486);
xor U2727 (N_2727,N_2412,N_2583);
or U2728 (N_2728,N_2451,N_2526);
or U2729 (N_2729,N_2410,N_2571);
or U2730 (N_2730,N_2506,N_2402);
or U2731 (N_2731,N_2553,N_2416);
or U2732 (N_2732,N_2456,N_2483);
xor U2733 (N_2733,N_2449,N_2567);
and U2734 (N_2734,N_2580,N_2485);
and U2735 (N_2735,N_2545,N_2440);
or U2736 (N_2736,N_2509,N_2513);
nand U2737 (N_2737,N_2470,N_2408);
nand U2738 (N_2738,N_2569,N_2507);
nand U2739 (N_2739,N_2511,N_2595);
xnor U2740 (N_2740,N_2581,N_2456);
nor U2741 (N_2741,N_2519,N_2577);
nor U2742 (N_2742,N_2413,N_2437);
or U2743 (N_2743,N_2520,N_2522);
nand U2744 (N_2744,N_2446,N_2414);
nor U2745 (N_2745,N_2477,N_2594);
nor U2746 (N_2746,N_2500,N_2483);
xnor U2747 (N_2747,N_2493,N_2425);
and U2748 (N_2748,N_2485,N_2470);
and U2749 (N_2749,N_2541,N_2510);
and U2750 (N_2750,N_2489,N_2499);
nand U2751 (N_2751,N_2484,N_2570);
and U2752 (N_2752,N_2536,N_2482);
or U2753 (N_2753,N_2400,N_2403);
and U2754 (N_2754,N_2440,N_2506);
and U2755 (N_2755,N_2505,N_2574);
nand U2756 (N_2756,N_2490,N_2551);
nand U2757 (N_2757,N_2584,N_2481);
or U2758 (N_2758,N_2482,N_2500);
or U2759 (N_2759,N_2406,N_2402);
nand U2760 (N_2760,N_2548,N_2594);
and U2761 (N_2761,N_2589,N_2471);
nand U2762 (N_2762,N_2463,N_2481);
nor U2763 (N_2763,N_2508,N_2577);
and U2764 (N_2764,N_2502,N_2559);
or U2765 (N_2765,N_2406,N_2492);
and U2766 (N_2766,N_2423,N_2552);
xor U2767 (N_2767,N_2565,N_2534);
xor U2768 (N_2768,N_2513,N_2444);
or U2769 (N_2769,N_2565,N_2457);
or U2770 (N_2770,N_2501,N_2475);
nand U2771 (N_2771,N_2521,N_2547);
or U2772 (N_2772,N_2458,N_2569);
or U2773 (N_2773,N_2585,N_2535);
and U2774 (N_2774,N_2501,N_2441);
and U2775 (N_2775,N_2448,N_2505);
nor U2776 (N_2776,N_2432,N_2463);
nor U2777 (N_2777,N_2504,N_2527);
nand U2778 (N_2778,N_2422,N_2527);
nand U2779 (N_2779,N_2452,N_2577);
nor U2780 (N_2780,N_2466,N_2500);
and U2781 (N_2781,N_2570,N_2509);
xor U2782 (N_2782,N_2476,N_2478);
nand U2783 (N_2783,N_2439,N_2487);
and U2784 (N_2784,N_2538,N_2505);
or U2785 (N_2785,N_2518,N_2599);
and U2786 (N_2786,N_2412,N_2448);
or U2787 (N_2787,N_2485,N_2433);
or U2788 (N_2788,N_2491,N_2507);
nor U2789 (N_2789,N_2436,N_2539);
and U2790 (N_2790,N_2428,N_2546);
and U2791 (N_2791,N_2497,N_2549);
xor U2792 (N_2792,N_2550,N_2521);
nor U2793 (N_2793,N_2401,N_2490);
or U2794 (N_2794,N_2430,N_2415);
and U2795 (N_2795,N_2535,N_2406);
nor U2796 (N_2796,N_2531,N_2454);
and U2797 (N_2797,N_2407,N_2467);
nor U2798 (N_2798,N_2497,N_2532);
nand U2799 (N_2799,N_2542,N_2521);
and U2800 (N_2800,N_2795,N_2783);
nor U2801 (N_2801,N_2677,N_2780);
xor U2802 (N_2802,N_2738,N_2704);
or U2803 (N_2803,N_2778,N_2727);
or U2804 (N_2804,N_2753,N_2664);
or U2805 (N_2805,N_2633,N_2752);
xor U2806 (N_2806,N_2608,N_2690);
and U2807 (N_2807,N_2676,N_2659);
or U2808 (N_2808,N_2697,N_2731);
xor U2809 (N_2809,N_2632,N_2730);
nor U2810 (N_2810,N_2662,N_2779);
xor U2811 (N_2811,N_2788,N_2652);
or U2812 (N_2812,N_2735,N_2777);
nor U2813 (N_2813,N_2737,N_2725);
nand U2814 (N_2814,N_2767,N_2768);
nand U2815 (N_2815,N_2713,N_2673);
and U2816 (N_2816,N_2774,N_2723);
nand U2817 (N_2817,N_2683,N_2601);
or U2818 (N_2818,N_2605,N_2651);
nand U2819 (N_2819,N_2760,N_2756);
nand U2820 (N_2820,N_2631,N_2609);
nand U2821 (N_2821,N_2695,N_2791);
or U2822 (N_2822,N_2610,N_2669);
nor U2823 (N_2823,N_2642,N_2649);
nand U2824 (N_2824,N_2734,N_2688);
nand U2825 (N_2825,N_2686,N_2627);
and U2826 (N_2826,N_2786,N_2739);
xnor U2827 (N_2827,N_2623,N_2702);
and U2828 (N_2828,N_2653,N_2660);
nand U2829 (N_2829,N_2687,N_2724);
or U2830 (N_2830,N_2674,N_2720);
nand U2831 (N_2831,N_2692,N_2604);
and U2832 (N_2832,N_2665,N_2773);
and U2833 (N_2833,N_2626,N_2717);
nor U2834 (N_2834,N_2728,N_2635);
or U2835 (N_2835,N_2707,N_2769);
nand U2836 (N_2836,N_2751,N_2775);
xor U2837 (N_2837,N_2616,N_2763);
xnor U2838 (N_2838,N_2696,N_2667);
or U2839 (N_2839,N_2655,N_2622);
nor U2840 (N_2840,N_2640,N_2625);
nor U2841 (N_2841,N_2785,N_2705);
nand U2842 (N_2842,N_2758,N_2617);
and U2843 (N_2843,N_2711,N_2666);
or U2844 (N_2844,N_2618,N_2663);
xnor U2845 (N_2845,N_2733,N_2634);
or U2846 (N_2846,N_2754,N_2603);
nand U2847 (N_2847,N_2797,N_2790);
nor U2848 (N_2848,N_2619,N_2643);
and U2849 (N_2849,N_2799,N_2680);
or U2850 (N_2850,N_2722,N_2787);
and U2851 (N_2851,N_2743,N_2691);
or U2852 (N_2852,N_2796,N_2689);
xnor U2853 (N_2853,N_2636,N_2670);
nor U2854 (N_2854,N_2793,N_2709);
and U2855 (N_2855,N_2715,N_2607);
and U2856 (N_2856,N_2710,N_2654);
and U2857 (N_2857,N_2766,N_2741);
nand U2858 (N_2858,N_2721,N_2650);
nor U2859 (N_2859,N_2745,N_2716);
and U2860 (N_2860,N_2776,N_2638);
and U2861 (N_2861,N_2679,N_2606);
or U2862 (N_2862,N_2755,N_2684);
and U2863 (N_2863,N_2742,N_2613);
and U2864 (N_2864,N_2628,N_2759);
nor U2865 (N_2865,N_2600,N_2614);
or U2866 (N_2866,N_2789,N_2764);
xnor U2867 (N_2867,N_2668,N_2639);
and U2868 (N_2868,N_2732,N_2749);
nand U2869 (N_2869,N_2646,N_2693);
and U2870 (N_2870,N_2784,N_2637);
or U2871 (N_2871,N_2656,N_2761);
and U2872 (N_2872,N_2748,N_2700);
and U2873 (N_2873,N_2706,N_2672);
and U2874 (N_2874,N_2611,N_2681);
nand U2875 (N_2875,N_2729,N_2675);
nor U2876 (N_2876,N_2740,N_2624);
nor U2877 (N_2877,N_2644,N_2602);
nor U2878 (N_2878,N_2762,N_2736);
nand U2879 (N_2879,N_2694,N_2621);
nand U2880 (N_2880,N_2657,N_2661);
nand U2881 (N_2881,N_2718,N_2703);
nor U2882 (N_2882,N_2772,N_2792);
xor U2883 (N_2883,N_2771,N_2648);
nand U2884 (N_2884,N_2658,N_2781);
and U2885 (N_2885,N_2615,N_2712);
or U2886 (N_2886,N_2629,N_2770);
nand U2887 (N_2887,N_2612,N_2641);
xor U2888 (N_2888,N_2794,N_2744);
or U2889 (N_2889,N_2698,N_2782);
nand U2890 (N_2890,N_2647,N_2701);
or U2891 (N_2891,N_2765,N_2708);
nand U2892 (N_2892,N_2671,N_2798);
nand U2893 (N_2893,N_2719,N_2757);
or U2894 (N_2894,N_2678,N_2685);
or U2895 (N_2895,N_2630,N_2750);
or U2896 (N_2896,N_2714,N_2726);
or U2897 (N_2897,N_2747,N_2746);
or U2898 (N_2898,N_2699,N_2645);
nor U2899 (N_2899,N_2682,N_2620);
nor U2900 (N_2900,N_2722,N_2766);
nand U2901 (N_2901,N_2654,N_2736);
xor U2902 (N_2902,N_2793,N_2780);
xor U2903 (N_2903,N_2682,N_2616);
nor U2904 (N_2904,N_2646,N_2747);
or U2905 (N_2905,N_2631,N_2672);
and U2906 (N_2906,N_2635,N_2679);
nand U2907 (N_2907,N_2642,N_2799);
or U2908 (N_2908,N_2641,N_2758);
nand U2909 (N_2909,N_2790,N_2744);
nand U2910 (N_2910,N_2752,N_2603);
or U2911 (N_2911,N_2621,N_2778);
nand U2912 (N_2912,N_2694,N_2730);
xnor U2913 (N_2913,N_2745,N_2691);
or U2914 (N_2914,N_2603,N_2635);
xnor U2915 (N_2915,N_2677,N_2632);
or U2916 (N_2916,N_2778,N_2655);
and U2917 (N_2917,N_2774,N_2705);
nor U2918 (N_2918,N_2749,N_2664);
or U2919 (N_2919,N_2657,N_2761);
or U2920 (N_2920,N_2670,N_2754);
or U2921 (N_2921,N_2609,N_2649);
nor U2922 (N_2922,N_2732,N_2621);
or U2923 (N_2923,N_2754,N_2655);
or U2924 (N_2924,N_2671,N_2751);
or U2925 (N_2925,N_2603,N_2788);
or U2926 (N_2926,N_2754,N_2796);
and U2927 (N_2927,N_2643,N_2783);
nand U2928 (N_2928,N_2621,N_2776);
xor U2929 (N_2929,N_2649,N_2739);
or U2930 (N_2930,N_2791,N_2767);
or U2931 (N_2931,N_2714,N_2664);
nor U2932 (N_2932,N_2704,N_2688);
nor U2933 (N_2933,N_2632,N_2670);
xnor U2934 (N_2934,N_2616,N_2799);
nand U2935 (N_2935,N_2687,N_2627);
or U2936 (N_2936,N_2600,N_2790);
and U2937 (N_2937,N_2781,N_2728);
or U2938 (N_2938,N_2782,N_2696);
and U2939 (N_2939,N_2778,N_2669);
nand U2940 (N_2940,N_2742,N_2645);
and U2941 (N_2941,N_2715,N_2685);
and U2942 (N_2942,N_2669,N_2635);
and U2943 (N_2943,N_2757,N_2763);
nor U2944 (N_2944,N_2774,N_2778);
or U2945 (N_2945,N_2725,N_2773);
nand U2946 (N_2946,N_2750,N_2691);
xor U2947 (N_2947,N_2640,N_2642);
and U2948 (N_2948,N_2753,N_2640);
and U2949 (N_2949,N_2710,N_2749);
or U2950 (N_2950,N_2662,N_2673);
xnor U2951 (N_2951,N_2691,N_2682);
nand U2952 (N_2952,N_2709,N_2671);
and U2953 (N_2953,N_2669,N_2603);
and U2954 (N_2954,N_2699,N_2623);
nor U2955 (N_2955,N_2792,N_2646);
or U2956 (N_2956,N_2719,N_2793);
nand U2957 (N_2957,N_2660,N_2666);
and U2958 (N_2958,N_2621,N_2604);
nor U2959 (N_2959,N_2621,N_2710);
nand U2960 (N_2960,N_2610,N_2674);
xnor U2961 (N_2961,N_2628,N_2647);
nand U2962 (N_2962,N_2642,N_2728);
and U2963 (N_2963,N_2694,N_2686);
nand U2964 (N_2964,N_2764,N_2737);
nor U2965 (N_2965,N_2678,N_2688);
or U2966 (N_2966,N_2674,N_2606);
xnor U2967 (N_2967,N_2614,N_2611);
xor U2968 (N_2968,N_2698,N_2625);
or U2969 (N_2969,N_2773,N_2639);
nand U2970 (N_2970,N_2655,N_2725);
and U2971 (N_2971,N_2657,N_2635);
or U2972 (N_2972,N_2738,N_2615);
nand U2973 (N_2973,N_2651,N_2775);
and U2974 (N_2974,N_2792,N_2734);
nor U2975 (N_2975,N_2795,N_2737);
nand U2976 (N_2976,N_2603,N_2643);
xor U2977 (N_2977,N_2618,N_2651);
and U2978 (N_2978,N_2675,N_2616);
and U2979 (N_2979,N_2779,N_2658);
nor U2980 (N_2980,N_2617,N_2715);
nand U2981 (N_2981,N_2762,N_2643);
nor U2982 (N_2982,N_2781,N_2607);
or U2983 (N_2983,N_2729,N_2746);
or U2984 (N_2984,N_2687,N_2754);
or U2985 (N_2985,N_2696,N_2741);
and U2986 (N_2986,N_2716,N_2749);
nor U2987 (N_2987,N_2766,N_2668);
and U2988 (N_2988,N_2714,N_2619);
nor U2989 (N_2989,N_2784,N_2690);
or U2990 (N_2990,N_2644,N_2605);
nand U2991 (N_2991,N_2664,N_2614);
nand U2992 (N_2992,N_2734,N_2673);
nor U2993 (N_2993,N_2695,N_2737);
or U2994 (N_2994,N_2766,N_2638);
and U2995 (N_2995,N_2690,N_2665);
or U2996 (N_2996,N_2735,N_2687);
nand U2997 (N_2997,N_2790,N_2623);
and U2998 (N_2998,N_2657,N_2765);
or U2999 (N_2999,N_2613,N_2638);
nand UO_0 (O_0,N_2866,N_2860);
nor UO_1 (O_1,N_2804,N_2997);
and UO_2 (O_2,N_2824,N_2940);
and UO_3 (O_3,N_2835,N_2894);
or UO_4 (O_4,N_2851,N_2806);
and UO_5 (O_5,N_2996,N_2810);
nor UO_6 (O_6,N_2879,N_2842);
and UO_7 (O_7,N_2950,N_2888);
nand UO_8 (O_8,N_2926,N_2920);
and UO_9 (O_9,N_2915,N_2838);
xor UO_10 (O_10,N_2887,N_2972);
nor UO_11 (O_11,N_2977,N_2832);
nor UO_12 (O_12,N_2812,N_2858);
nor UO_13 (O_13,N_2949,N_2979);
and UO_14 (O_14,N_2957,N_2992);
or UO_15 (O_15,N_2864,N_2813);
or UO_16 (O_16,N_2811,N_2966);
nand UO_17 (O_17,N_2924,N_2880);
nor UO_18 (O_18,N_2905,N_2937);
or UO_19 (O_19,N_2857,N_2931);
or UO_20 (O_20,N_2827,N_2981);
xor UO_21 (O_21,N_2897,N_2876);
nand UO_22 (O_22,N_2985,N_2934);
or UO_23 (O_23,N_2840,N_2906);
nor UO_24 (O_24,N_2903,N_2984);
or UO_25 (O_25,N_2976,N_2823);
and UO_26 (O_26,N_2862,N_2890);
and UO_27 (O_27,N_2875,N_2961);
and UO_28 (O_28,N_2891,N_2834);
nor UO_29 (O_29,N_2816,N_2861);
nand UO_30 (O_30,N_2854,N_2807);
xor UO_31 (O_31,N_2973,N_2913);
and UO_32 (O_32,N_2874,N_2809);
or UO_33 (O_33,N_2922,N_2872);
nor UO_34 (O_34,N_2945,N_2941);
nor UO_35 (O_35,N_2983,N_2871);
nor UO_36 (O_36,N_2898,N_2955);
and UO_37 (O_37,N_2882,N_2946);
and UO_38 (O_38,N_2819,N_2930);
xor UO_39 (O_39,N_2933,N_2829);
nor UO_40 (O_40,N_2837,N_2974);
nor UO_41 (O_41,N_2918,N_2938);
or UO_42 (O_42,N_2896,N_2952);
nand UO_43 (O_43,N_2849,N_2803);
nand UO_44 (O_44,N_2883,N_2867);
or UO_45 (O_45,N_2942,N_2911);
nand UO_46 (O_46,N_2947,N_2999);
or UO_47 (O_47,N_2841,N_2919);
and UO_48 (O_48,N_2873,N_2828);
or UO_49 (O_49,N_2923,N_2969);
or UO_50 (O_50,N_2989,N_2825);
and UO_51 (O_51,N_2865,N_2956);
nand UO_52 (O_52,N_2970,N_2801);
or UO_53 (O_53,N_2893,N_2948);
nor UO_54 (O_54,N_2800,N_2988);
and UO_55 (O_55,N_2987,N_2939);
or UO_56 (O_56,N_2892,N_2993);
or UO_57 (O_57,N_2895,N_2845);
nand UO_58 (O_58,N_2843,N_2982);
nand UO_59 (O_59,N_2986,N_2953);
and UO_60 (O_60,N_2971,N_2967);
nor UO_61 (O_61,N_2991,N_2826);
nand UO_62 (O_62,N_2932,N_2886);
nor UO_63 (O_63,N_2877,N_2912);
or UO_64 (O_64,N_2889,N_2910);
or UO_65 (O_65,N_2960,N_2869);
nor UO_66 (O_66,N_2847,N_2990);
nand UO_67 (O_67,N_2808,N_2878);
nand UO_68 (O_68,N_2975,N_2954);
xor UO_69 (O_69,N_2850,N_2968);
nand UO_70 (O_70,N_2901,N_2815);
nor UO_71 (O_71,N_2929,N_2814);
xnor UO_72 (O_72,N_2936,N_2964);
or UO_73 (O_73,N_2963,N_2925);
nor UO_74 (O_74,N_2881,N_2818);
nand UO_75 (O_75,N_2909,N_2943);
xnor UO_76 (O_76,N_2994,N_2836);
and UO_77 (O_77,N_2853,N_2908);
nand UO_78 (O_78,N_2852,N_2927);
xor UO_79 (O_79,N_2907,N_2805);
and UO_80 (O_80,N_2928,N_2830);
or UO_81 (O_81,N_2856,N_2914);
or UO_82 (O_82,N_2916,N_2833);
nand UO_83 (O_83,N_2917,N_2821);
nand UO_84 (O_84,N_2802,N_2859);
and UO_85 (O_85,N_2839,N_2900);
nand UO_86 (O_86,N_2855,N_2935);
or UO_87 (O_87,N_2958,N_2959);
nand UO_88 (O_88,N_2884,N_2868);
xor UO_89 (O_89,N_2844,N_2995);
and UO_90 (O_90,N_2978,N_2822);
xnor UO_91 (O_91,N_2870,N_2921);
nand UO_92 (O_92,N_2831,N_2820);
nor UO_93 (O_93,N_2962,N_2998);
and UO_94 (O_94,N_2944,N_2902);
nand UO_95 (O_95,N_2980,N_2846);
or UO_96 (O_96,N_2904,N_2817);
and UO_97 (O_97,N_2848,N_2951);
nand UO_98 (O_98,N_2965,N_2899);
nor UO_99 (O_99,N_2885,N_2863);
xnor UO_100 (O_100,N_2855,N_2967);
and UO_101 (O_101,N_2813,N_2947);
nand UO_102 (O_102,N_2878,N_2995);
or UO_103 (O_103,N_2832,N_2838);
xnor UO_104 (O_104,N_2992,N_2976);
and UO_105 (O_105,N_2820,N_2812);
xor UO_106 (O_106,N_2879,N_2832);
nor UO_107 (O_107,N_2811,N_2947);
xnor UO_108 (O_108,N_2814,N_2926);
or UO_109 (O_109,N_2924,N_2905);
and UO_110 (O_110,N_2949,N_2859);
nor UO_111 (O_111,N_2913,N_2974);
or UO_112 (O_112,N_2974,N_2894);
or UO_113 (O_113,N_2904,N_2886);
or UO_114 (O_114,N_2995,N_2837);
or UO_115 (O_115,N_2993,N_2845);
nand UO_116 (O_116,N_2822,N_2995);
or UO_117 (O_117,N_2923,N_2961);
and UO_118 (O_118,N_2893,N_2973);
or UO_119 (O_119,N_2984,N_2921);
and UO_120 (O_120,N_2977,N_2863);
or UO_121 (O_121,N_2910,N_2993);
nor UO_122 (O_122,N_2857,N_2956);
nand UO_123 (O_123,N_2973,N_2816);
xnor UO_124 (O_124,N_2826,N_2949);
or UO_125 (O_125,N_2862,N_2924);
nand UO_126 (O_126,N_2812,N_2829);
nor UO_127 (O_127,N_2930,N_2989);
nand UO_128 (O_128,N_2954,N_2948);
nand UO_129 (O_129,N_2880,N_2963);
and UO_130 (O_130,N_2875,N_2940);
nand UO_131 (O_131,N_2873,N_2935);
nor UO_132 (O_132,N_2857,N_2806);
nand UO_133 (O_133,N_2900,N_2897);
nor UO_134 (O_134,N_2811,N_2929);
nor UO_135 (O_135,N_2868,N_2963);
nor UO_136 (O_136,N_2854,N_2850);
or UO_137 (O_137,N_2986,N_2868);
nand UO_138 (O_138,N_2941,N_2924);
nand UO_139 (O_139,N_2964,N_2997);
and UO_140 (O_140,N_2876,N_2887);
and UO_141 (O_141,N_2851,N_2929);
and UO_142 (O_142,N_2867,N_2932);
xnor UO_143 (O_143,N_2980,N_2919);
nand UO_144 (O_144,N_2990,N_2917);
nand UO_145 (O_145,N_2986,N_2963);
or UO_146 (O_146,N_2890,N_2845);
and UO_147 (O_147,N_2985,N_2999);
and UO_148 (O_148,N_2904,N_2854);
nor UO_149 (O_149,N_2887,N_2985);
or UO_150 (O_150,N_2918,N_2874);
or UO_151 (O_151,N_2962,N_2836);
and UO_152 (O_152,N_2862,N_2922);
or UO_153 (O_153,N_2900,N_2986);
nand UO_154 (O_154,N_2960,N_2935);
nor UO_155 (O_155,N_2843,N_2959);
and UO_156 (O_156,N_2804,N_2852);
nand UO_157 (O_157,N_2808,N_2907);
xnor UO_158 (O_158,N_2971,N_2928);
or UO_159 (O_159,N_2868,N_2952);
nor UO_160 (O_160,N_2840,N_2948);
nand UO_161 (O_161,N_2832,N_2894);
and UO_162 (O_162,N_2837,N_2858);
and UO_163 (O_163,N_2983,N_2959);
nor UO_164 (O_164,N_2936,N_2878);
xnor UO_165 (O_165,N_2874,N_2988);
and UO_166 (O_166,N_2925,N_2832);
and UO_167 (O_167,N_2876,N_2808);
nor UO_168 (O_168,N_2904,N_2835);
or UO_169 (O_169,N_2883,N_2918);
nand UO_170 (O_170,N_2851,N_2927);
or UO_171 (O_171,N_2979,N_2891);
nand UO_172 (O_172,N_2813,N_2844);
or UO_173 (O_173,N_2949,N_2966);
xor UO_174 (O_174,N_2850,N_2878);
nor UO_175 (O_175,N_2992,N_2889);
and UO_176 (O_176,N_2950,N_2850);
or UO_177 (O_177,N_2909,N_2814);
nand UO_178 (O_178,N_2892,N_2947);
nand UO_179 (O_179,N_2911,N_2987);
and UO_180 (O_180,N_2987,N_2905);
nand UO_181 (O_181,N_2824,N_2890);
or UO_182 (O_182,N_2835,N_2821);
nand UO_183 (O_183,N_2855,N_2925);
or UO_184 (O_184,N_2942,N_2893);
nor UO_185 (O_185,N_2946,N_2870);
or UO_186 (O_186,N_2874,N_2987);
nand UO_187 (O_187,N_2887,N_2838);
or UO_188 (O_188,N_2899,N_2816);
nand UO_189 (O_189,N_2965,N_2846);
and UO_190 (O_190,N_2850,N_2947);
nand UO_191 (O_191,N_2895,N_2901);
nand UO_192 (O_192,N_2827,N_2985);
nor UO_193 (O_193,N_2878,N_2866);
nor UO_194 (O_194,N_2866,N_2899);
xor UO_195 (O_195,N_2867,N_2961);
nand UO_196 (O_196,N_2976,N_2989);
and UO_197 (O_197,N_2854,N_2813);
nand UO_198 (O_198,N_2825,N_2870);
nor UO_199 (O_199,N_2992,N_2935);
nor UO_200 (O_200,N_2872,N_2921);
or UO_201 (O_201,N_2952,N_2856);
or UO_202 (O_202,N_2958,N_2866);
and UO_203 (O_203,N_2991,N_2830);
or UO_204 (O_204,N_2895,N_2832);
xor UO_205 (O_205,N_2897,N_2888);
nor UO_206 (O_206,N_2981,N_2965);
and UO_207 (O_207,N_2904,N_2961);
nand UO_208 (O_208,N_2897,N_2986);
or UO_209 (O_209,N_2981,N_2808);
nor UO_210 (O_210,N_2887,N_2895);
nor UO_211 (O_211,N_2932,N_2929);
nor UO_212 (O_212,N_2984,N_2842);
xnor UO_213 (O_213,N_2828,N_2838);
or UO_214 (O_214,N_2931,N_2966);
nand UO_215 (O_215,N_2840,N_2914);
nor UO_216 (O_216,N_2873,N_2899);
nand UO_217 (O_217,N_2913,N_2986);
nor UO_218 (O_218,N_2829,N_2823);
nor UO_219 (O_219,N_2969,N_2863);
nor UO_220 (O_220,N_2974,N_2985);
or UO_221 (O_221,N_2889,N_2931);
or UO_222 (O_222,N_2916,N_2838);
nor UO_223 (O_223,N_2964,N_2863);
xor UO_224 (O_224,N_2962,N_2858);
nor UO_225 (O_225,N_2930,N_2948);
or UO_226 (O_226,N_2876,N_2804);
xnor UO_227 (O_227,N_2972,N_2936);
nor UO_228 (O_228,N_2935,N_2829);
nor UO_229 (O_229,N_2821,N_2973);
nor UO_230 (O_230,N_2819,N_2988);
nor UO_231 (O_231,N_2979,N_2965);
or UO_232 (O_232,N_2884,N_2990);
nand UO_233 (O_233,N_2801,N_2819);
and UO_234 (O_234,N_2957,N_2852);
nand UO_235 (O_235,N_2867,N_2832);
and UO_236 (O_236,N_2881,N_2967);
nand UO_237 (O_237,N_2956,N_2908);
and UO_238 (O_238,N_2834,N_2979);
nand UO_239 (O_239,N_2974,N_2917);
and UO_240 (O_240,N_2841,N_2955);
or UO_241 (O_241,N_2837,N_2920);
nor UO_242 (O_242,N_2901,N_2991);
nand UO_243 (O_243,N_2958,N_2817);
and UO_244 (O_244,N_2807,N_2989);
or UO_245 (O_245,N_2863,N_2904);
xnor UO_246 (O_246,N_2888,N_2813);
nand UO_247 (O_247,N_2883,N_2999);
nor UO_248 (O_248,N_2833,N_2947);
xor UO_249 (O_249,N_2890,N_2967);
xor UO_250 (O_250,N_2954,N_2891);
nor UO_251 (O_251,N_2985,N_2982);
or UO_252 (O_252,N_2994,N_2943);
nor UO_253 (O_253,N_2991,N_2995);
nand UO_254 (O_254,N_2838,N_2864);
nand UO_255 (O_255,N_2923,N_2850);
nor UO_256 (O_256,N_2858,N_2807);
nand UO_257 (O_257,N_2924,N_2949);
and UO_258 (O_258,N_2822,N_2897);
or UO_259 (O_259,N_2812,N_2873);
or UO_260 (O_260,N_2951,N_2906);
nor UO_261 (O_261,N_2812,N_2836);
nand UO_262 (O_262,N_2977,N_2916);
and UO_263 (O_263,N_2941,N_2949);
nand UO_264 (O_264,N_2900,N_2808);
nor UO_265 (O_265,N_2868,N_2874);
nor UO_266 (O_266,N_2825,N_2929);
and UO_267 (O_267,N_2814,N_2935);
nand UO_268 (O_268,N_2818,N_2843);
xnor UO_269 (O_269,N_2873,N_2843);
or UO_270 (O_270,N_2904,N_2814);
or UO_271 (O_271,N_2850,N_2915);
nor UO_272 (O_272,N_2930,N_2910);
nand UO_273 (O_273,N_2809,N_2944);
nor UO_274 (O_274,N_2863,N_2922);
nor UO_275 (O_275,N_2889,N_2810);
and UO_276 (O_276,N_2958,N_2973);
and UO_277 (O_277,N_2894,N_2827);
or UO_278 (O_278,N_2928,N_2983);
nand UO_279 (O_279,N_2939,N_2811);
nor UO_280 (O_280,N_2802,N_2803);
and UO_281 (O_281,N_2961,N_2821);
nor UO_282 (O_282,N_2866,N_2869);
nand UO_283 (O_283,N_2801,N_2981);
or UO_284 (O_284,N_2843,N_2917);
or UO_285 (O_285,N_2867,N_2865);
xor UO_286 (O_286,N_2890,N_2989);
nand UO_287 (O_287,N_2859,N_2980);
xnor UO_288 (O_288,N_2951,N_2946);
or UO_289 (O_289,N_2815,N_2914);
and UO_290 (O_290,N_2922,N_2954);
or UO_291 (O_291,N_2912,N_2918);
nor UO_292 (O_292,N_2882,N_2889);
and UO_293 (O_293,N_2801,N_2897);
or UO_294 (O_294,N_2987,N_2805);
nor UO_295 (O_295,N_2956,N_2909);
nand UO_296 (O_296,N_2970,N_2819);
nand UO_297 (O_297,N_2964,N_2862);
nand UO_298 (O_298,N_2911,N_2849);
nor UO_299 (O_299,N_2805,N_2816);
and UO_300 (O_300,N_2968,N_2986);
xnor UO_301 (O_301,N_2957,N_2808);
nand UO_302 (O_302,N_2953,N_2855);
and UO_303 (O_303,N_2912,N_2887);
nor UO_304 (O_304,N_2837,N_2822);
nand UO_305 (O_305,N_2946,N_2868);
nand UO_306 (O_306,N_2843,N_2973);
nor UO_307 (O_307,N_2963,N_2896);
xnor UO_308 (O_308,N_2988,N_2853);
nand UO_309 (O_309,N_2985,N_2950);
or UO_310 (O_310,N_2861,N_2813);
nand UO_311 (O_311,N_2828,N_2814);
xor UO_312 (O_312,N_2919,N_2987);
xnor UO_313 (O_313,N_2862,N_2945);
nor UO_314 (O_314,N_2962,N_2911);
nor UO_315 (O_315,N_2919,N_2891);
nor UO_316 (O_316,N_2992,N_2987);
nor UO_317 (O_317,N_2997,N_2974);
or UO_318 (O_318,N_2824,N_2808);
xnor UO_319 (O_319,N_2942,N_2800);
and UO_320 (O_320,N_2970,N_2929);
nand UO_321 (O_321,N_2905,N_2991);
or UO_322 (O_322,N_2900,N_2823);
nand UO_323 (O_323,N_2833,N_2998);
nor UO_324 (O_324,N_2912,N_2852);
or UO_325 (O_325,N_2872,N_2887);
nand UO_326 (O_326,N_2829,N_2958);
or UO_327 (O_327,N_2995,N_2972);
or UO_328 (O_328,N_2945,N_2993);
nor UO_329 (O_329,N_2831,N_2823);
nor UO_330 (O_330,N_2830,N_2945);
xor UO_331 (O_331,N_2920,N_2884);
and UO_332 (O_332,N_2868,N_2918);
and UO_333 (O_333,N_2838,N_2928);
nor UO_334 (O_334,N_2826,N_2831);
nor UO_335 (O_335,N_2814,N_2915);
nand UO_336 (O_336,N_2844,N_2873);
or UO_337 (O_337,N_2800,N_2900);
nand UO_338 (O_338,N_2861,N_2884);
nand UO_339 (O_339,N_2950,N_2803);
nand UO_340 (O_340,N_2918,N_2872);
and UO_341 (O_341,N_2905,N_2807);
nand UO_342 (O_342,N_2834,N_2900);
nand UO_343 (O_343,N_2973,N_2910);
or UO_344 (O_344,N_2843,N_2831);
or UO_345 (O_345,N_2937,N_2883);
xor UO_346 (O_346,N_2975,N_2826);
nor UO_347 (O_347,N_2963,N_2940);
or UO_348 (O_348,N_2984,N_2849);
nand UO_349 (O_349,N_2910,N_2966);
or UO_350 (O_350,N_2813,N_2843);
or UO_351 (O_351,N_2829,N_2984);
nor UO_352 (O_352,N_2831,N_2911);
and UO_353 (O_353,N_2923,N_2976);
nand UO_354 (O_354,N_2987,N_2922);
nor UO_355 (O_355,N_2945,N_2854);
or UO_356 (O_356,N_2890,N_2806);
or UO_357 (O_357,N_2978,N_2949);
nor UO_358 (O_358,N_2928,N_2985);
nor UO_359 (O_359,N_2839,N_2952);
nor UO_360 (O_360,N_2831,N_2937);
nor UO_361 (O_361,N_2839,N_2975);
and UO_362 (O_362,N_2845,N_2837);
xnor UO_363 (O_363,N_2892,N_2972);
nand UO_364 (O_364,N_2980,N_2884);
nor UO_365 (O_365,N_2892,N_2849);
xor UO_366 (O_366,N_2939,N_2838);
nand UO_367 (O_367,N_2824,N_2835);
nand UO_368 (O_368,N_2965,N_2916);
or UO_369 (O_369,N_2827,N_2954);
and UO_370 (O_370,N_2976,N_2908);
and UO_371 (O_371,N_2966,N_2851);
or UO_372 (O_372,N_2803,N_2893);
or UO_373 (O_373,N_2810,N_2906);
nor UO_374 (O_374,N_2981,N_2822);
xnor UO_375 (O_375,N_2816,N_2877);
and UO_376 (O_376,N_2886,N_2990);
nand UO_377 (O_377,N_2894,N_2903);
nand UO_378 (O_378,N_2920,N_2959);
xnor UO_379 (O_379,N_2908,N_2933);
nand UO_380 (O_380,N_2918,N_2865);
nand UO_381 (O_381,N_2852,N_2975);
nor UO_382 (O_382,N_2985,N_2879);
nor UO_383 (O_383,N_2944,N_2901);
nor UO_384 (O_384,N_2908,N_2841);
nand UO_385 (O_385,N_2897,N_2804);
nand UO_386 (O_386,N_2941,N_2873);
and UO_387 (O_387,N_2963,N_2802);
and UO_388 (O_388,N_2820,N_2853);
nand UO_389 (O_389,N_2893,N_2830);
nor UO_390 (O_390,N_2853,N_2831);
nand UO_391 (O_391,N_2803,N_2919);
nor UO_392 (O_392,N_2965,N_2957);
xnor UO_393 (O_393,N_2839,N_2830);
or UO_394 (O_394,N_2969,N_2986);
or UO_395 (O_395,N_2872,N_2857);
or UO_396 (O_396,N_2879,N_2851);
and UO_397 (O_397,N_2874,N_2820);
nand UO_398 (O_398,N_2990,N_2965);
nand UO_399 (O_399,N_2890,N_2966);
nor UO_400 (O_400,N_2923,N_2941);
and UO_401 (O_401,N_2881,N_2945);
and UO_402 (O_402,N_2912,N_2999);
nand UO_403 (O_403,N_2981,N_2852);
xnor UO_404 (O_404,N_2872,N_2808);
nand UO_405 (O_405,N_2831,N_2879);
or UO_406 (O_406,N_2839,N_2849);
nor UO_407 (O_407,N_2878,N_2800);
or UO_408 (O_408,N_2889,N_2835);
nand UO_409 (O_409,N_2996,N_2958);
and UO_410 (O_410,N_2812,N_2854);
nor UO_411 (O_411,N_2854,N_2855);
nand UO_412 (O_412,N_2836,N_2840);
nand UO_413 (O_413,N_2958,N_2889);
or UO_414 (O_414,N_2835,N_2895);
nor UO_415 (O_415,N_2970,N_2950);
xnor UO_416 (O_416,N_2942,N_2803);
xnor UO_417 (O_417,N_2811,N_2961);
nor UO_418 (O_418,N_2851,N_2987);
nand UO_419 (O_419,N_2855,N_2923);
nor UO_420 (O_420,N_2947,N_2984);
xnor UO_421 (O_421,N_2994,N_2810);
and UO_422 (O_422,N_2996,N_2914);
nor UO_423 (O_423,N_2821,N_2853);
or UO_424 (O_424,N_2948,N_2855);
nand UO_425 (O_425,N_2852,N_2817);
nor UO_426 (O_426,N_2865,N_2911);
nand UO_427 (O_427,N_2973,N_2878);
nor UO_428 (O_428,N_2983,N_2839);
and UO_429 (O_429,N_2844,N_2820);
nand UO_430 (O_430,N_2985,N_2913);
xnor UO_431 (O_431,N_2963,N_2897);
nor UO_432 (O_432,N_2802,N_2999);
nor UO_433 (O_433,N_2938,N_2969);
nor UO_434 (O_434,N_2994,N_2885);
nand UO_435 (O_435,N_2839,N_2841);
nor UO_436 (O_436,N_2845,N_2852);
or UO_437 (O_437,N_2977,N_2823);
and UO_438 (O_438,N_2904,N_2820);
nand UO_439 (O_439,N_2935,N_2816);
and UO_440 (O_440,N_2808,N_2870);
or UO_441 (O_441,N_2931,N_2820);
nand UO_442 (O_442,N_2931,N_2828);
nor UO_443 (O_443,N_2874,N_2957);
and UO_444 (O_444,N_2862,N_2844);
or UO_445 (O_445,N_2935,N_2968);
nor UO_446 (O_446,N_2982,N_2888);
nand UO_447 (O_447,N_2938,N_2949);
xor UO_448 (O_448,N_2919,N_2929);
nand UO_449 (O_449,N_2993,N_2954);
and UO_450 (O_450,N_2857,N_2913);
or UO_451 (O_451,N_2810,N_2921);
or UO_452 (O_452,N_2947,N_2917);
xnor UO_453 (O_453,N_2939,N_2823);
xor UO_454 (O_454,N_2838,N_2873);
nand UO_455 (O_455,N_2976,N_2816);
or UO_456 (O_456,N_2915,N_2929);
or UO_457 (O_457,N_2972,N_2827);
nand UO_458 (O_458,N_2843,N_2985);
nor UO_459 (O_459,N_2916,N_2868);
and UO_460 (O_460,N_2901,N_2805);
nor UO_461 (O_461,N_2959,N_2806);
or UO_462 (O_462,N_2929,N_2897);
and UO_463 (O_463,N_2961,N_2967);
nor UO_464 (O_464,N_2885,N_2912);
and UO_465 (O_465,N_2864,N_2957);
xnor UO_466 (O_466,N_2884,N_2934);
nand UO_467 (O_467,N_2816,N_2852);
and UO_468 (O_468,N_2926,N_2931);
nor UO_469 (O_469,N_2823,N_2811);
nand UO_470 (O_470,N_2972,N_2836);
nor UO_471 (O_471,N_2976,N_2855);
or UO_472 (O_472,N_2860,N_2917);
and UO_473 (O_473,N_2836,N_2864);
nor UO_474 (O_474,N_2852,N_2878);
nor UO_475 (O_475,N_2938,N_2906);
xor UO_476 (O_476,N_2845,N_2916);
xor UO_477 (O_477,N_2851,N_2823);
and UO_478 (O_478,N_2947,N_2849);
or UO_479 (O_479,N_2826,N_2955);
and UO_480 (O_480,N_2962,N_2942);
xnor UO_481 (O_481,N_2850,N_2919);
nor UO_482 (O_482,N_2879,N_2995);
nor UO_483 (O_483,N_2913,N_2950);
nor UO_484 (O_484,N_2823,N_2962);
nand UO_485 (O_485,N_2901,N_2833);
nand UO_486 (O_486,N_2896,N_2847);
and UO_487 (O_487,N_2996,N_2880);
and UO_488 (O_488,N_2888,N_2953);
nor UO_489 (O_489,N_2899,N_2811);
and UO_490 (O_490,N_2933,N_2800);
or UO_491 (O_491,N_2927,N_2937);
xor UO_492 (O_492,N_2941,N_2915);
or UO_493 (O_493,N_2817,N_2871);
or UO_494 (O_494,N_2888,N_2981);
nor UO_495 (O_495,N_2988,N_2805);
nand UO_496 (O_496,N_2941,N_2928);
nor UO_497 (O_497,N_2835,N_2905);
nand UO_498 (O_498,N_2843,N_2800);
nand UO_499 (O_499,N_2871,N_2870);
endmodule