module basic_750_5000_1000_5_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_257,In_358);
nand U1 (N_1,In_535,In_360);
and U2 (N_2,In_318,In_136);
nor U3 (N_3,In_573,In_471);
or U4 (N_4,In_221,In_339);
and U5 (N_5,In_348,In_73);
nand U6 (N_6,In_186,In_503);
and U7 (N_7,In_4,In_292);
or U8 (N_8,In_351,In_240);
or U9 (N_9,In_95,In_706);
and U10 (N_10,In_261,In_116);
or U11 (N_11,In_330,In_671);
nor U12 (N_12,In_310,In_316);
and U13 (N_13,In_622,In_396);
or U14 (N_14,In_599,In_420);
and U15 (N_15,In_490,In_407);
or U16 (N_16,In_170,In_556);
nor U17 (N_17,In_506,In_476);
or U18 (N_18,In_75,In_642);
or U19 (N_19,In_434,In_14);
nand U20 (N_20,In_25,In_362);
nor U21 (N_21,In_593,In_250);
and U22 (N_22,In_210,In_206);
and U23 (N_23,In_495,In_524);
or U24 (N_24,In_543,In_349);
and U25 (N_25,In_686,In_595);
nor U26 (N_26,In_284,In_588);
and U27 (N_27,In_294,In_20);
and U28 (N_28,In_201,In_224);
nor U29 (N_29,In_167,In_392);
and U30 (N_30,In_322,In_522);
or U31 (N_31,In_426,In_67);
and U32 (N_32,In_165,In_118);
or U33 (N_33,In_679,In_600);
or U34 (N_34,In_323,In_291);
or U35 (N_35,In_277,In_460);
nor U36 (N_36,In_16,In_333);
nor U37 (N_37,In_24,In_41);
and U38 (N_38,In_602,In_704);
or U39 (N_39,In_367,In_590);
and U40 (N_40,In_43,In_244);
nand U41 (N_41,In_158,In_681);
nand U42 (N_42,In_701,In_619);
and U43 (N_43,In_492,In_368);
nor U44 (N_44,In_587,In_419);
nand U45 (N_45,In_189,In_427);
and U46 (N_46,In_370,In_161);
nor U47 (N_47,In_327,In_440);
or U48 (N_48,In_612,In_585);
or U49 (N_49,In_733,In_516);
nor U50 (N_50,In_504,In_26);
and U51 (N_51,In_262,In_698);
nand U52 (N_52,In_449,In_29);
and U53 (N_53,In_744,In_636);
or U54 (N_54,In_480,In_107);
and U55 (N_55,In_93,In_450);
nand U56 (N_56,In_313,In_32);
or U57 (N_57,In_695,In_68);
nor U58 (N_58,In_501,In_238);
nor U59 (N_59,In_552,In_463);
nand U60 (N_60,In_731,In_63);
nor U61 (N_61,In_547,In_180);
and U62 (N_62,In_464,In_306);
or U63 (N_63,In_336,In_727);
and U64 (N_64,In_70,In_468);
and U65 (N_65,In_168,In_28);
and U66 (N_66,In_272,In_138);
and U67 (N_67,In_613,In_246);
or U68 (N_68,In_565,In_641);
nand U69 (N_69,In_705,In_694);
and U70 (N_70,In_36,In_536);
nand U71 (N_71,In_363,In_69);
and U72 (N_72,In_187,In_149);
nor U73 (N_73,In_532,In_27);
nor U74 (N_74,In_5,In_675);
nor U75 (N_75,In_15,In_541);
nand U76 (N_76,In_331,In_231);
nor U77 (N_77,In_605,In_634);
or U78 (N_78,In_620,In_345);
nand U79 (N_79,In_53,In_315);
nand U80 (N_80,In_376,In_472);
or U81 (N_81,In_281,In_720);
nand U82 (N_82,In_126,In_309);
or U83 (N_83,In_483,In_544);
and U84 (N_84,In_559,In_373);
nor U85 (N_85,In_269,In_160);
or U86 (N_86,In_117,In_743);
nand U87 (N_87,In_132,In_729);
or U88 (N_88,In_576,In_498);
nor U89 (N_89,In_656,In_438);
or U90 (N_90,In_655,In_665);
nor U91 (N_91,In_410,In_652);
nand U92 (N_92,In_44,In_623);
nor U93 (N_93,In_216,In_539);
and U94 (N_94,In_265,In_23);
or U95 (N_95,In_403,In_562);
nor U96 (N_96,In_494,In_79);
nand U97 (N_97,In_629,In_283);
or U98 (N_98,In_305,In_597);
or U99 (N_99,In_399,In_275);
nor U100 (N_100,In_65,In_371);
nor U101 (N_101,In_430,In_418);
or U102 (N_102,In_437,In_372);
nand U103 (N_103,In_156,In_645);
nor U104 (N_104,In_726,In_582);
nand U105 (N_105,In_337,In_550);
nor U106 (N_106,In_81,In_62);
and U107 (N_107,In_435,In_299);
nor U108 (N_108,In_431,In_596);
and U109 (N_109,In_130,In_215);
nor U110 (N_110,In_626,In_542);
or U111 (N_111,In_135,In_718);
nand U112 (N_112,In_604,In_3);
nand U113 (N_113,In_97,In_555);
or U114 (N_114,In_445,In_157);
or U115 (N_115,In_179,In_611);
or U116 (N_116,In_683,In_572);
or U117 (N_117,In_98,In_297);
nor U118 (N_118,In_200,In_659);
nor U119 (N_119,In_227,In_346);
nand U120 (N_120,In_690,In_329);
and U121 (N_121,In_499,In_377);
nor U122 (N_122,In_394,In_223);
nand U123 (N_123,In_577,In_512);
nand U124 (N_124,In_405,In_293);
or U125 (N_125,In_57,In_134);
or U126 (N_126,In_379,In_112);
and U127 (N_127,In_575,In_166);
or U128 (N_128,In_198,In_458);
and U129 (N_129,In_260,In_228);
and U130 (N_130,In_99,In_508);
nor U131 (N_131,In_343,In_52);
or U132 (N_132,In_510,In_74);
nor U133 (N_133,In_666,In_314);
nand U134 (N_134,In_670,In_267);
or U135 (N_135,In_185,In_728);
and U136 (N_136,In_13,In_563);
and U137 (N_137,In_312,In_719);
and U138 (N_138,In_153,In_355);
and U139 (N_139,In_553,In_571);
nand U140 (N_140,In_411,In_442);
or U141 (N_141,In_457,In_129);
nor U142 (N_142,In_621,In_569);
nor U143 (N_143,In_661,In_644);
and U144 (N_144,In_658,In_513);
and U145 (N_145,In_252,In_321);
or U146 (N_146,In_567,In_692);
nor U147 (N_147,In_342,In_691);
and U148 (N_148,In_366,In_338);
and U149 (N_149,In_748,In_183);
nor U150 (N_150,In_341,In_48);
and U151 (N_151,In_255,In_326);
nand U152 (N_152,In_359,In_745);
nor U153 (N_153,In_172,In_459);
nand U154 (N_154,In_609,In_101);
and U155 (N_155,In_296,In_311);
and U156 (N_156,In_266,In_251);
nor U157 (N_157,In_664,In_702);
nor U158 (N_158,In_689,In_643);
nor U159 (N_159,In_102,In_398);
nand U160 (N_160,In_710,In_334);
and U161 (N_161,In_663,In_518);
nand U162 (N_162,In_628,In_159);
nand U163 (N_163,In_625,In_415);
and U164 (N_164,In_213,In_236);
or U165 (N_165,In_182,In_328);
or U166 (N_166,In_162,In_303);
nor U167 (N_167,In_466,In_638);
or U168 (N_168,In_12,In_648);
nand U169 (N_169,In_127,In_601);
nand U170 (N_170,In_493,In_249);
nand U171 (N_171,In_523,In_538);
nand U172 (N_172,In_64,In_491);
and U173 (N_173,In_361,In_150);
nor U174 (N_174,In_667,In_416);
nor U175 (N_175,In_340,In_531);
nor U176 (N_176,In_365,In_247);
and U177 (N_177,In_10,In_594);
or U178 (N_178,In_274,In_732);
nand U179 (N_179,In_549,In_651);
or U180 (N_180,In_712,In_222);
nand U181 (N_181,In_196,In_708);
nand U182 (N_182,In_724,In_421);
nor U183 (N_183,In_711,In_17);
nand U184 (N_184,In_395,In_288);
nand U185 (N_185,In_402,In_46);
nand U186 (N_186,In_557,In_680);
nor U187 (N_187,In_143,In_624);
and U188 (N_188,In_540,In_233);
or U189 (N_189,In_214,In_39);
nand U190 (N_190,In_615,In_649);
nand U191 (N_191,In_717,In_389);
and U192 (N_192,In_703,In_470);
and U193 (N_193,In_509,In_635);
nand U194 (N_194,In_113,In_232);
and U195 (N_195,In_248,In_465);
nand U196 (N_196,In_114,In_614);
and U197 (N_197,In_105,In_104);
nor U198 (N_198,In_7,In_738);
nor U199 (N_199,In_59,In_413);
and U200 (N_200,In_86,In_482);
and U201 (N_201,In_80,In_696);
nor U202 (N_202,In_324,In_525);
and U203 (N_203,In_357,In_401);
or U204 (N_204,In_146,In_447);
nor U205 (N_205,In_374,In_320);
and U206 (N_206,In_546,In_106);
and U207 (N_207,In_171,In_137);
or U208 (N_208,In_739,In_78);
nand U209 (N_209,In_647,In_253);
or U210 (N_210,In_287,In_583);
or U211 (N_211,In_0,In_519);
nand U212 (N_212,In_205,In_742);
nand U213 (N_213,In_1,In_264);
nor U214 (N_214,In_534,In_225);
and U215 (N_215,In_486,In_259);
and U216 (N_216,In_424,In_388);
nor U217 (N_217,In_479,In_607);
and U218 (N_218,In_242,In_528);
nand U219 (N_219,In_497,In_674);
nor U220 (N_220,In_409,In_688);
nand U221 (N_221,In_735,In_347);
nand U222 (N_222,In_85,In_352);
nor U223 (N_223,In_489,In_737);
nor U224 (N_224,In_488,In_481);
or U225 (N_225,In_131,In_527);
or U226 (N_226,In_397,In_746);
nor U227 (N_227,In_515,In_617);
and U228 (N_228,In_496,In_278);
and U229 (N_229,In_404,In_382);
nor U230 (N_230,In_685,In_715);
nand U231 (N_231,In_124,In_428);
nor U232 (N_232,In_653,In_684);
or U233 (N_233,In_22,In_608);
nor U234 (N_234,In_241,In_422);
nor U235 (N_235,In_574,In_190);
nor U236 (N_236,In_660,In_406);
or U237 (N_237,In_592,In_34);
and U238 (N_238,In_254,In_603);
and U239 (N_239,In_687,In_475);
or U240 (N_240,In_256,In_61);
nand U241 (N_241,In_42,In_672);
and U242 (N_242,In_484,In_175);
nor U243 (N_243,In_616,In_469);
nand U244 (N_244,In_386,In_290);
nand U245 (N_245,In_178,In_375);
or U246 (N_246,In_353,In_91);
and U247 (N_247,In_474,In_521);
nand U248 (N_248,In_417,In_123);
and U249 (N_249,In_207,In_530);
and U250 (N_250,In_217,In_630);
nand U251 (N_251,In_699,In_286);
nor U252 (N_252,In_195,In_258);
nand U253 (N_253,In_66,In_237);
or U254 (N_254,In_441,In_443);
and U255 (N_255,In_700,In_586);
and U256 (N_256,In_133,In_45);
nor U257 (N_257,In_268,In_707);
nor U258 (N_258,In_220,In_94);
nand U259 (N_259,In_736,In_35);
nand U260 (N_260,In_335,In_282);
nand U261 (N_261,In_298,In_747);
and U262 (N_262,In_423,In_439);
and U263 (N_263,In_354,In_657);
or U264 (N_264,In_204,In_451);
nand U265 (N_265,In_177,In_721);
or U266 (N_266,In_208,In_304);
nand U267 (N_267,In_148,In_212);
or U268 (N_268,In_56,In_164);
nand U269 (N_269,In_570,In_425);
nor U270 (N_270,In_199,In_125);
nand U271 (N_271,In_332,In_285);
and U272 (N_272,In_115,In_414);
nor U273 (N_273,In_151,In_722);
nand U274 (N_274,In_239,In_72);
nand U275 (N_275,In_30,In_551);
or U276 (N_276,In_84,In_245);
nand U277 (N_277,In_307,In_144);
or U278 (N_278,In_537,In_561);
xnor U279 (N_279,In_589,In_381);
and U280 (N_280,In_194,In_693);
and U281 (N_281,In_507,In_502);
or U282 (N_282,In_673,In_369);
or U283 (N_283,In_76,In_90);
nand U284 (N_284,In_654,In_77);
or U285 (N_285,In_325,In_723);
or U286 (N_286,In_568,In_174);
nor U287 (N_287,In_122,In_218);
and U288 (N_288,In_610,In_640);
or U289 (N_289,In_432,In_669);
nand U290 (N_290,In_209,In_446);
or U291 (N_291,In_477,In_140);
nand U292 (N_292,In_92,In_109);
nor U293 (N_293,In_120,In_50);
or U294 (N_294,In_580,In_100);
or U295 (N_295,In_230,In_142);
and U296 (N_296,In_716,In_154);
nand U297 (N_297,In_485,In_678);
nand U298 (N_298,In_234,In_300);
or U299 (N_299,In_37,In_197);
nor U300 (N_300,In_581,In_383);
and U301 (N_301,In_713,In_749);
and U302 (N_302,In_55,In_147);
or U303 (N_303,In_203,In_83);
nor U304 (N_304,In_520,In_650);
nor U305 (N_305,In_181,In_219);
xnor U306 (N_306,In_380,In_356);
nand U307 (N_307,In_89,In_505);
nor U308 (N_308,In_364,In_633);
nand U309 (N_309,In_47,In_54);
or U310 (N_310,In_40,In_243);
nand U311 (N_311,In_631,In_58);
or U312 (N_312,In_526,In_514);
or U313 (N_313,In_176,In_71);
or U314 (N_314,In_578,In_591);
nand U315 (N_315,In_725,In_662);
and U316 (N_316,In_682,In_229);
nand U317 (N_317,In_226,In_408);
xnor U318 (N_318,In_145,In_139);
and U319 (N_319,In_271,In_155);
or U320 (N_320,In_734,In_487);
nand U321 (N_321,In_19,In_280);
and U322 (N_322,In_344,In_308);
nor U323 (N_323,In_128,In_51);
nor U324 (N_324,In_639,In_202);
or U325 (N_325,In_319,In_632);
or U326 (N_326,In_211,In_387);
and U327 (N_327,In_270,In_730);
nor U328 (N_328,In_677,In_276);
or U329 (N_329,In_21,In_235);
nand U330 (N_330,In_49,In_385);
nand U331 (N_331,In_558,In_455);
or U332 (N_332,In_301,In_714);
nand U333 (N_333,In_152,In_412);
nand U334 (N_334,In_317,In_709);
or U335 (N_335,In_478,In_88);
nor U336 (N_336,In_627,In_31);
nor U337 (N_337,In_646,In_511);
nor U338 (N_338,In_545,In_9);
and U339 (N_339,In_393,In_668);
nand U340 (N_340,In_6,In_110);
or U341 (N_341,In_429,In_467);
nand U342 (N_342,In_163,In_584);
or U343 (N_343,In_384,In_350);
nor U344 (N_344,In_8,In_448);
and U345 (N_345,In_579,In_141);
or U346 (N_346,In_444,In_566);
nand U347 (N_347,In_289,In_184);
nand U348 (N_348,In_87,In_391);
and U349 (N_349,In_188,In_454);
or U350 (N_350,In_462,In_529);
nand U351 (N_351,In_18,In_461);
nand U352 (N_352,In_740,In_554);
and U353 (N_353,In_169,In_598);
nor U354 (N_354,In_606,In_191);
nor U355 (N_355,In_453,In_697);
nand U356 (N_356,In_436,In_96);
and U357 (N_357,In_302,In_618);
and U358 (N_358,In_533,In_279);
and U359 (N_359,In_548,In_517);
nand U360 (N_360,In_108,In_173);
and U361 (N_361,In_192,In_111);
and U362 (N_362,In_400,In_38);
nand U363 (N_363,In_456,In_560);
or U364 (N_364,In_741,In_263);
nor U365 (N_365,In_390,In_273);
or U366 (N_366,In_82,In_452);
and U367 (N_367,In_637,In_60);
or U368 (N_368,In_11,In_564);
and U369 (N_369,In_119,In_500);
nor U370 (N_370,In_433,In_295);
nand U371 (N_371,In_103,In_676);
nand U372 (N_372,In_473,In_2);
nand U373 (N_373,In_378,In_33);
nor U374 (N_374,In_193,In_121);
or U375 (N_375,In_331,In_473);
and U376 (N_376,In_389,In_289);
and U377 (N_377,In_599,In_167);
and U378 (N_378,In_321,In_225);
and U379 (N_379,In_188,In_30);
or U380 (N_380,In_181,In_460);
nand U381 (N_381,In_409,In_202);
and U382 (N_382,In_92,In_622);
and U383 (N_383,In_497,In_344);
nand U384 (N_384,In_348,In_744);
and U385 (N_385,In_277,In_598);
nor U386 (N_386,In_590,In_20);
or U387 (N_387,In_208,In_211);
nor U388 (N_388,In_736,In_462);
and U389 (N_389,In_507,In_632);
xnor U390 (N_390,In_248,In_121);
and U391 (N_391,In_83,In_701);
and U392 (N_392,In_536,In_353);
nor U393 (N_393,In_60,In_28);
nor U394 (N_394,In_548,In_98);
nand U395 (N_395,In_17,In_237);
and U396 (N_396,In_661,In_626);
nor U397 (N_397,In_210,In_279);
nand U398 (N_398,In_471,In_738);
and U399 (N_399,In_627,In_292);
or U400 (N_400,In_677,In_584);
nor U401 (N_401,In_212,In_242);
and U402 (N_402,In_17,In_314);
nor U403 (N_403,In_110,In_568);
or U404 (N_404,In_230,In_389);
nor U405 (N_405,In_638,In_526);
nor U406 (N_406,In_154,In_354);
or U407 (N_407,In_745,In_387);
nor U408 (N_408,In_664,In_676);
and U409 (N_409,In_225,In_560);
nand U410 (N_410,In_540,In_732);
nor U411 (N_411,In_47,In_616);
and U412 (N_412,In_585,In_305);
nor U413 (N_413,In_403,In_647);
nor U414 (N_414,In_553,In_315);
and U415 (N_415,In_276,In_274);
nor U416 (N_416,In_701,In_133);
nor U417 (N_417,In_340,In_302);
and U418 (N_418,In_253,In_387);
nand U419 (N_419,In_422,In_543);
and U420 (N_420,In_542,In_83);
nand U421 (N_421,In_130,In_691);
or U422 (N_422,In_626,In_372);
nor U423 (N_423,In_583,In_75);
nand U424 (N_424,In_487,In_193);
nor U425 (N_425,In_741,In_710);
and U426 (N_426,In_205,In_741);
and U427 (N_427,In_337,In_503);
nor U428 (N_428,In_286,In_108);
nor U429 (N_429,In_229,In_596);
and U430 (N_430,In_359,In_519);
or U431 (N_431,In_312,In_482);
and U432 (N_432,In_7,In_222);
or U433 (N_433,In_725,In_261);
and U434 (N_434,In_466,In_133);
nor U435 (N_435,In_39,In_267);
or U436 (N_436,In_413,In_150);
nor U437 (N_437,In_443,In_170);
and U438 (N_438,In_415,In_512);
and U439 (N_439,In_500,In_81);
or U440 (N_440,In_251,In_241);
nand U441 (N_441,In_345,In_214);
nand U442 (N_442,In_487,In_522);
nor U443 (N_443,In_189,In_27);
nand U444 (N_444,In_373,In_148);
or U445 (N_445,In_489,In_668);
nand U446 (N_446,In_296,In_116);
or U447 (N_447,In_213,In_510);
and U448 (N_448,In_148,In_223);
and U449 (N_449,In_626,In_91);
and U450 (N_450,In_171,In_262);
and U451 (N_451,In_344,In_116);
nor U452 (N_452,In_492,In_241);
and U453 (N_453,In_230,In_160);
nor U454 (N_454,In_11,In_648);
nand U455 (N_455,In_89,In_321);
or U456 (N_456,In_158,In_293);
and U457 (N_457,In_690,In_98);
and U458 (N_458,In_571,In_306);
and U459 (N_459,In_683,In_193);
and U460 (N_460,In_117,In_680);
or U461 (N_461,In_211,In_657);
nor U462 (N_462,In_495,In_533);
or U463 (N_463,In_92,In_170);
or U464 (N_464,In_145,In_244);
nor U465 (N_465,In_578,In_590);
and U466 (N_466,In_70,In_449);
nor U467 (N_467,In_559,In_699);
nand U468 (N_468,In_204,In_523);
nand U469 (N_469,In_707,In_340);
nand U470 (N_470,In_107,In_242);
and U471 (N_471,In_591,In_289);
or U472 (N_472,In_262,In_172);
nor U473 (N_473,In_556,In_719);
nand U474 (N_474,In_4,In_201);
or U475 (N_475,In_351,In_574);
nor U476 (N_476,In_434,In_613);
or U477 (N_477,In_261,In_744);
nand U478 (N_478,In_102,In_213);
or U479 (N_479,In_190,In_172);
nand U480 (N_480,In_530,In_200);
and U481 (N_481,In_461,In_21);
nand U482 (N_482,In_431,In_740);
and U483 (N_483,In_211,In_396);
or U484 (N_484,In_615,In_285);
or U485 (N_485,In_542,In_513);
nand U486 (N_486,In_183,In_53);
or U487 (N_487,In_349,In_59);
and U488 (N_488,In_624,In_374);
nor U489 (N_489,In_357,In_250);
nor U490 (N_490,In_71,In_570);
or U491 (N_491,In_610,In_537);
nand U492 (N_492,In_213,In_306);
nand U493 (N_493,In_728,In_146);
nand U494 (N_494,In_356,In_53);
xnor U495 (N_495,In_580,In_488);
and U496 (N_496,In_559,In_730);
nand U497 (N_497,In_725,In_139);
and U498 (N_498,In_631,In_257);
nand U499 (N_499,In_402,In_569);
or U500 (N_500,In_689,In_369);
and U501 (N_501,In_310,In_581);
nor U502 (N_502,In_589,In_610);
nand U503 (N_503,In_284,In_206);
nor U504 (N_504,In_36,In_704);
nor U505 (N_505,In_45,In_717);
nor U506 (N_506,In_530,In_633);
nor U507 (N_507,In_83,In_347);
nand U508 (N_508,In_22,In_130);
or U509 (N_509,In_199,In_325);
or U510 (N_510,In_444,In_154);
and U511 (N_511,In_106,In_256);
nor U512 (N_512,In_239,In_705);
and U513 (N_513,In_670,In_526);
or U514 (N_514,In_500,In_573);
nand U515 (N_515,In_320,In_184);
or U516 (N_516,In_242,In_552);
and U517 (N_517,In_375,In_72);
nand U518 (N_518,In_292,In_563);
or U519 (N_519,In_580,In_621);
or U520 (N_520,In_388,In_576);
or U521 (N_521,In_672,In_727);
nand U522 (N_522,In_413,In_741);
nor U523 (N_523,In_309,In_429);
nor U524 (N_524,In_629,In_351);
nand U525 (N_525,In_373,In_80);
or U526 (N_526,In_294,In_67);
and U527 (N_527,In_231,In_425);
nand U528 (N_528,In_149,In_686);
nor U529 (N_529,In_498,In_495);
nand U530 (N_530,In_641,In_232);
nor U531 (N_531,In_708,In_435);
or U532 (N_532,In_97,In_618);
nor U533 (N_533,In_680,In_71);
nand U534 (N_534,In_37,In_320);
or U535 (N_535,In_221,In_63);
nand U536 (N_536,In_478,In_266);
nor U537 (N_537,In_532,In_352);
and U538 (N_538,In_340,In_404);
xnor U539 (N_539,In_114,In_403);
nand U540 (N_540,In_515,In_618);
and U541 (N_541,In_286,In_476);
xor U542 (N_542,In_651,In_131);
or U543 (N_543,In_157,In_438);
nor U544 (N_544,In_659,In_612);
nand U545 (N_545,In_193,In_280);
nand U546 (N_546,In_122,In_615);
or U547 (N_547,In_110,In_270);
and U548 (N_548,In_60,In_479);
nand U549 (N_549,In_671,In_284);
or U550 (N_550,In_446,In_481);
and U551 (N_551,In_630,In_20);
nor U552 (N_552,In_233,In_142);
or U553 (N_553,In_738,In_478);
and U554 (N_554,In_82,In_259);
or U555 (N_555,In_447,In_73);
nor U556 (N_556,In_74,In_120);
nand U557 (N_557,In_18,In_451);
or U558 (N_558,In_705,In_586);
nor U559 (N_559,In_719,In_178);
or U560 (N_560,In_744,In_223);
nand U561 (N_561,In_384,In_428);
or U562 (N_562,In_245,In_316);
nand U563 (N_563,In_196,In_305);
and U564 (N_564,In_33,In_556);
xor U565 (N_565,In_456,In_473);
nand U566 (N_566,In_272,In_63);
nand U567 (N_567,In_280,In_179);
or U568 (N_568,In_642,In_46);
or U569 (N_569,In_298,In_729);
nor U570 (N_570,In_189,In_522);
and U571 (N_571,In_343,In_717);
nor U572 (N_572,In_105,In_342);
or U573 (N_573,In_611,In_431);
nor U574 (N_574,In_309,In_561);
or U575 (N_575,In_108,In_185);
nor U576 (N_576,In_503,In_433);
nor U577 (N_577,In_0,In_323);
nand U578 (N_578,In_570,In_703);
nor U579 (N_579,In_735,In_208);
xor U580 (N_580,In_89,In_563);
and U581 (N_581,In_457,In_742);
nand U582 (N_582,In_317,In_123);
nand U583 (N_583,In_578,In_141);
nand U584 (N_584,In_22,In_579);
nor U585 (N_585,In_427,In_530);
nor U586 (N_586,In_196,In_303);
and U587 (N_587,In_546,In_349);
and U588 (N_588,In_252,In_52);
nor U589 (N_589,In_15,In_625);
and U590 (N_590,In_661,In_723);
or U591 (N_591,In_415,In_361);
nor U592 (N_592,In_638,In_113);
and U593 (N_593,In_288,In_2);
and U594 (N_594,In_131,In_318);
nand U595 (N_595,In_692,In_472);
nand U596 (N_596,In_7,In_107);
and U597 (N_597,In_719,In_138);
and U598 (N_598,In_236,In_691);
and U599 (N_599,In_1,In_386);
and U600 (N_600,In_181,In_21);
nand U601 (N_601,In_12,In_140);
or U602 (N_602,In_166,In_597);
nor U603 (N_603,In_390,In_582);
nand U604 (N_604,In_700,In_150);
nor U605 (N_605,In_0,In_531);
and U606 (N_606,In_217,In_185);
nand U607 (N_607,In_506,In_565);
or U608 (N_608,In_262,In_98);
nor U609 (N_609,In_644,In_281);
and U610 (N_610,In_290,In_219);
nand U611 (N_611,In_644,In_714);
and U612 (N_612,In_491,In_699);
and U613 (N_613,In_351,In_608);
or U614 (N_614,In_102,In_588);
or U615 (N_615,In_539,In_601);
or U616 (N_616,In_67,In_490);
nor U617 (N_617,In_354,In_99);
or U618 (N_618,In_485,In_44);
nor U619 (N_619,In_39,In_126);
nor U620 (N_620,In_731,In_275);
or U621 (N_621,In_109,In_626);
xor U622 (N_622,In_666,In_147);
nor U623 (N_623,In_127,In_106);
or U624 (N_624,In_706,In_52);
nand U625 (N_625,In_459,In_247);
and U626 (N_626,In_222,In_308);
nand U627 (N_627,In_563,In_363);
nand U628 (N_628,In_705,In_134);
nand U629 (N_629,In_749,In_22);
and U630 (N_630,In_206,In_29);
and U631 (N_631,In_297,In_727);
nor U632 (N_632,In_481,In_484);
and U633 (N_633,In_193,In_742);
nor U634 (N_634,In_365,In_576);
nor U635 (N_635,In_194,In_477);
and U636 (N_636,In_290,In_465);
nand U637 (N_637,In_602,In_570);
and U638 (N_638,In_258,In_178);
nand U639 (N_639,In_305,In_547);
nor U640 (N_640,In_459,In_701);
nand U641 (N_641,In_410,In_343);
nor U642 (N_642,In_75,In_677);
or U643 (N_643,In_730,In_369);
or U644 (N_644,In_324,In_214);
xor U645 (N_645,In_260,In_547);
and U646 (N_646,In_573,In_306);
and U647 (N_647,In_41,In_467);
or U648 (N_648,In_246,In_137);
nand U649 (N_649,In_420,In_12);
and U650 (N_650,In_546,In_332);
or U651 (N_651,In_552,In_231);
and U652 (N_652,In_287,In_615);
or U653 (N_653,In_467,In_485);
and U654 (N_654,In_7,In_339);
or U655 (N_655,In_189,In_418);
and U656 (N_656,In_637,In_523);
and U657 (N_657,In_124,In_714);
and U658 (N_658,In_528,In_195);
or U659 (N_659,In_93,In_665);
or U660 (N_660,In_696,In_221);
nor U661 (N_661,In_236,In_210);
or U662 (N_662,In_214,In_43);
or U663 (N_663,In_248,In_419);
and U664 (N_664,In_319,In_364);
nor U665 (N_665,In_430,In_325);
nand U666 (N_666,In_727,In_558);
and U667 (N_667,In_19,In_558);
nor U668 (N_668,In_722,In_645);
nand U669 (N_669,In_314,In_325);
and U670 (N_670,In_13,In_258);
or U671 (N_671,In_442,In_338);
and U672 (N_672,In_413,In_360);
nand U673 (N_673,In_171,In_119);
nor U674 (N_674,In_44,In_64);
nand U675 (N_675,In_500,In_209);
and U676 (N_676,In_452,In_388);
nand U677 (N_677,In_523,In_453);
nor U678 (N_678,In_366,In_232);
nor U679 (N_679,In_353,In_295);
and U680 (N_680,In_505,In_345);
and U681 (N_681,In_120,In_90);
nand U682 (N_682,In_82,In_45);
and U683 (N_683,In_436,In_219);
and U684 (N_684,In_243,In_11);
nand U685 (N_685,In_655,In_305);
nor U686 (N_686,In_423,In_455);
and U687 (N_687,In_341,In_262);
and U688 (N_688,In_420,In_494);
nand U689 (N_689,In_425,In_470);
nor U690 (N_690,In_86,In_528);
and U691 (N_691,In_167,In_36);
nand U692 (N_692,In_86,In_594);
nor U693 (N_693,In_412,In_28);
nor U694 (N_694,In_520,In_140);
or U695 (N_695,In_606,In_57);
nor U696 (N_696,In_204,In_713);
nor U697 (N_697,In_241,In_580);
and U698 (N_698,In_643,In_329);
nor U699 (N_699,In_466,In_254);
nor U700 (N_700,In_451,In_393);
xnor U701 (N_701,In_202,In_401);
nand U702 (N_702,In_265,In_395);
and U703 (N_703,In_540,In_537);
nor U704 (N_704,In_732,In_488);
and U705 (N_705,In_447,In_416);
nand U706 (N_706,In_314,In_726);
or U707 (N_707,In_596,In_612);
nand U708 (N_708,In_679,In_394);
nor U709 (N_709,In_275,In_620);
and U710 (N_710,In_179,In_500);
and U711 (N_711,In_462,In_463);
or U712 (N_712,In_249,In_252);
and U713 (N_713,In_479,In_297);
and U714 (N_714,In_302,In_626);
or U715 (N_715,In_644,In_575);
nand U716 (N_716,In_196,In_397);
nand U717 (N_717,In_62,In_477);
and U718 (N_718,In_301,In_428);
nand U719 (N_719,In_155,In_33);
nor U720 (N_720,In_226,In_686);
and U721 (N_721,In_562,In_19);
and U722 (N_722,In_479,In_433);
nand U723 (N_723,In_51,In_687);
nor U724 (N_724,In_156,In_340);
nor U725 (N_725,In_588,In_27);
or U726 (N_726,In_416,In_549);
nand U727 (N_727,In_106,In_510);
nor U728 (N_728,In_359,In_174);
nor U729 (N_729,In_612,In_554);
nor U730 (N_730,In_13,In_463);
nand U731 (N_731,In_236,In_67);
or U732 (N_732,In_178,In_449);
nand U733 (N_733,In_352,In_64);
or U734 (N_734,In_498,In_146);
or U735 (N_735,In_447,In_410);
and U736 (N_736,In_519,In_529);
and U737 (N_737,In_87,In_108);
nand U738 (N_738,In_556,In_264);
and U739 (N_739,In_182,In_661);
and U740 (N_740,In_370,In_693);
nand U741 (N_741,In_21,In_613);
and U742 (N_742,In_436,In_207);
nor U743 (N_743,In_577,In_432);
and U744 (N_744,In_197,In_586);
nor U745 (N_745,In_223,In_291);
and U746 (N_746,In_749,In_630);
and U747 (N_747,In_161,In_314);
or U748 (N_748,In_563,In_234);
or U749 (N_749,In_728,In_166);
and U750 (N_750,In_216,In_469);
and U751 (N_751,In_41,In_617);
or U752 (N_752,In_16,In_749);
or U753 (N_753,In_444,In_59);
nand U754 (N_754,In_242,In_740);
nor U755 (N_755,In_680,In_251);
nor U756 (N_756,In_512,In_348);
and U757 (N_757,In_572,In_89);
nand U758 (N_758,In_496,In_138);
nand U759 (N_759,In_489,In_676);
nor U760 (N_760,In_599,In_574);
nand U761 (N_761,In_698,In_91);
nand U762 (N_762,In_181,In_537);
nor U763 (N_763,In_197,In_236);
or U764 (N_764,In_249,In_455);
nor U765 (N_765,In_717,In_48);
or U766 (N_766,In_281,In_542);
or U767 (N_767,In_159,In_47);
nand U768 (N_768,In_642,In_245);
and U769 (N_769,In_129,In_249);
nor U770 (N_770,In_36,In_307);
nor U771 (N_771,In_654,In_95);
or U772 (N_772,In_4,In_28);
or U773 (N_773,In_477,In_391);
nor U774 (N_774,In_233,In_709);
nand U775 (N_775,In_369,In_129);
and U776 (N_776,In_104,In_143);
nand U777 (N_777,In_406,In_71);
nand U778 (N_778,In_668,In_74);
nand U779 (N_779,In_50,In_399);
nand U780 (N_780,In_653,In_391);
nor U781 (N_781,In_197,In_720);
nand U782 (N_782,In_45,In_528);
or U783 (N_783,In_127,In_555);
nor U784 (N_784,In_24,In_370);
or U785 (N_785,In_486,In_269);
nor U786 (N_786,In_30,In_212);
nand U787 (N_787,In_628,In_406);
or U788 (N_788,In_241,In_379);
nor U789 (N_789,In_256,In_622);
nand U790 (N_790,In_179,In_478);
and U791 (N_791,In_401,In_308);
and U792 (N_792,In_469,In_313);
and U793 (N_793,In_712,In_613);
nand U794 (N_794,In_162,In_723);
or U795 (N_795,In_538,In_378);
and U796 (N_796,In_642,In_673);
or U797 (N_797,In_484,In_210);
nand U798 (N_798,In_567,In_661);
nor U799 (N_799,In_491,In_473);
or U800 (N_800,In_411,In_371);
nand U801 (N_801,In_539,In_262);
and U802 (N_802,In_497,In_535);
or U803 (N_803,In_649,In_696);
or U804 (N_804,In_488,In_518);
and U805 (N_805,In_672,In_30);
nand U806 (N_806,In_167,In_331);
or U807 (N_807,In_661,In_472);
nor U808 (N_808,In_299,In_104);
nand U809 (N_809,In_734,In_700);
nand U810 (N_810,In_112,In_685);
and U811 (N_811,In_175,In_673);
or U812 (N_812,In_209,In_155);
and U813 (N_813,In_294,In_202);
and U814 (N_814,In_150,In_149);
nand U815 (N_815,In_147,In_590);
and U816 (N_816,In_336,In_419);
and U817 (N_817,In_599,In_673);
and U818 (N_818,In_348,In_469);
nand U819 (N_819,In_465,In_196);
nand U820 (N_820,In_251,In_720);
nand U821 (N_821,In_534,In_586);
nand U822 (N_822,In_407,In_377);
and U823 (N_823,In_116,In_323);
nor U824 (N_824,In_219,In_681);
and U825 (N_825,In_62,In_426);
or U826 (N_826,In_477,In_571);
or U827 (N_827,In_203,In_722);
nor U828 (N_828,In_191,In_342);
nor U829 (N_829,In_401,In_23);
nand U830 (N_830,In_130,In_475);
nand U831 (N_831,In_447,In_681);
or U832 (N_832,In_382,In_93);
and U833 (N_833,In_227,In_292);
xnor U834 (N_834,In_121,In_353);
nor U835 (N_835,In_448,In_198);
and U836 (N_836,In_401,In_348);
and U837 (N_837,In_191,In_525);
and U838 (N_838,In_337,In_214);
and U839 (N_839,In_7,In_423);
nor U840 (N_840,In_124,In_748);
and U841 (N_841,In_137,In_668);
nor U842 (N_842,In_267,In_311);
or U843 (N_843,In_643,In_430);
nand U844 (N_844,In_742,In_580);
nand U845 (N_845,In_107,In_96);
and U846 (N_846,In_314,In_308);
or U847 (N_847,In_253,In_631);
or U848 (N_848,In_600,In_531);
or U849 (N_849,In_651,In_331);
and U850 (N_850,In_234,In_286);
and U851 (N_851,In_162,In_481);
nand U852 (N_852,In_30,In_239);
or U853 (N_853,In_746,In_524);
nor U854 (N_854,In_401,In_522);
and U855 (N_855,In_62,In_215);
nand U856 (N_856,In_609,In_261);
and U857 (N_857,In_50,In_211);
nor U858 (N_858,In_247,In_226);
nor U859 (N_859,In_174,In_159);
nand U860 (N_860,In_42,In_218);
or U861 (N_861,In_464,In_253);
nor U862 (N_862,In_694,In_382);
or U863 (N_863,In_258,In_539);
nand U864 (N_864,In_445,In_143);
or U865 (N_865,In_44,In_718);
nand U866 (N_866,In_237,In_652);
or U867 (N_867,In_279,In_283);
nand U868 (N_868,In_168,In_119);
and U869 (N_869,In_303,In_80);
xor U870 (N_870,In_104,In_313);
nand U871 (N_871,In_302,In_571);
or U872 (N_872,In_9,In_434);
and U873 (N_873,In_540,In_490);
nand U874 (N_874,In_582,In_240);
nor U875 (N_875,In_597,In_304);
and U876 (N_876,In_419,In_13);
and U877 (N_877,In_566,In_308);
and U878 (N_878,In_405,In_231);
xnor U879 (N_879,In_482,In_182);
or U880 (N_880,In_678,In_467);
nor U881 (N_881,In_94,In_77);
or U882 (N_882,In_728,In_165);
nand U883 (N_883,In_310,In_92);
and U884 (N_884,In_366,In_173);
nor U885 (N_885,In_682,In_733);
and U886 (N_886,In_319,In_276);
nor U887 (N_887,In_129,In_436);
nand U888 (N_888,In_397,In_388);
nor U889 (N_889,In_676,In_46);
or U890 (N_890,In_381,In_107);
nor U891 (N_891,In_212,In_469);
nor U892 (N_892,In_207,In_567);
nor U893 (N_893,In_625,In_150);
or U894 (N_894,In_374,In_286);
and U895 (N_895,In_432,In_302);
or U896 (N_896,In_668,In_634);
nor U897 (N_897,In_367,In_53);
or U898 (N_898,In_637,In_543);
and U899 (N_899,In_522,In_127);
nand U900 (N_900,In_691,In_526);
nor U901 (N_901,In_375,In_486);
or U902 (N_902,In_609,In_661);
nand U903 (N_903,In_296,In_176);
or U904 (N_904,In_91,In_517);
or U905 (N_905,In_371,In_710);
nor U906 (N_906,In_711,In_329);
nand U907 (N_907,In_537,In_22);
and U908 (N_908,In_93,In_290);
and U909 (N_909,In_696,In_531);
and U910 (N_910,In_518,In_497);
nor U911 (N_911,In_83,In_547);
and U912 (N_912,In_589,In_272);
nand U913 (N_913,In_270,In_599);
nand U914 (N_914,In_350,In_35);
nor U915 (N_915,In_617,In_388);
nor U916 (N_916,In_471,In_599);
nand U917 (N_917,In_82,In_631);
and U918 (N_918,In_533,In_525);
nand U919 (N_919,In_130,In_234);
nand U920 (N_920,In_207,In_179);
or U921 (N_921,In_599,In_238);
nor U922 (N_922,In_123,In_505);
nand U923 (N_923,In_364,In_342);
nand U924 (N_924,In_200,In_362);
nand U925 (N_925,In_408,In_319);
and U926 (N_926,In_191,In_225);
and U927 (N_927,In_641,In_414);
and U928 (N_928,In_365,In_747);
nor U929 (N_929,In_186,In_75);
and U930 (N_930,In_731,In_461);
nor U931 (N_931,In_539,In_33);
or U932 (N_932,In_699,In_553);
or U933 (N_933,In_732,In_265);
or U934 (N_934,In_147,In_655);
nor U935 (N_935,In_730,In_38);
or U936 (N_936,In_594,In_63);
nand U937 (N_937,In_621,In_556);
nor U938 (N_938,In_55,In_563);
nor U939 (N_939,In_458,In_354);
nand U940 (N_940,In_527,In_115);
or U941 (N_941,In_101,In_312);
and U942 (N_942,In_558,In_132);
nor U943 (N_943,In_348,In_710);
nor U944 (N_944,In_603,In_93);
nand U945 (N_945,In_594,In_324);
nand U946 (N_946,In_287,In_594);
and U947 (N_947,In_506,In_343);
and U948 (N_948,In_376,In_188);
nor U949 (N_949,In_476,In_133);
or U950 (N_950,In_141,In_477);
and U951 (N_951,In_681,In_239);
nor U952 (N_952,In_137,In_312);
nor U953 (N_953,In_470,In_207);
or U954 (N_954,In_373,In_724);
nor U955 (N_955,In_205,In_334);
nand U956 (N_956,In_679,In_61);
nand U957 (N_957,In_586,In_435);
or U958 (N_958,In_417,In_591);
nor U959 (N_959,In_518,In_120);
nor U960 (N_960,In_492,In_169);
or U961 (N_961,In_127,In_440);
and U962 (N_962,In_142,In_128);
and U963 (N_963,In_177,In_64);
and U964 (N_964,In_78,In_667);
or U965 (N_965,In_701,In_237);
nor U966 (N_966,In_344,In_634);
nor U967 (N_967,In_337,In_114);
nor U968 (N_968,In_522,In_532);
nor U969 (N_969,In_402,In_489);
nor U970 (N_970,In_690,In_362);
and U971 (N_971,In_142,In_655);
nand U972 (N_972,In_379,In_93);
nor U973 (N_973,In_442,In_503);
or U974 (N_974,In_544,In_740);
or U975 (N_975,In_121,In_127);
and U976 (N_976,In_147,In_445);
nor U977 (N_977,In_95,In_637);
nand U978 (N_978,In_133,In_749);
nand U979 (N_979,In_269,In_290);
and U980 (N_980,In_611,In_217);
and U981 (N_981,In_682,In_216);
nand U982 (N_982,In_667,In_680);
and U983 (N_983,In_297,In_113);
nor U984 (N_984,In_104,In_321);
and U985 (N_985,In_416,In_25);
and U986 (N_986,In_72,In_259);
and U987 (N_987,In_130,In_575);
nor U988 (N_988,In_593,In_529);
nand U989 (N_989,In_104,In_630);
nand U990 (N_990,In_137,In_12);
nor U991 (N_991,In_453,In_288);
and U992 (N_992,In_112,In_665);
or U993 (N_993,In_268,In_285);
nor U994 (N_994,In_698,In_143);
nand U995 (N_995,In_607,In_218);
nand U996 (N_996,In_419,In_406);
xnor U997 (N_997,In_694,In_325);
or U998 (N_998,In_494,In_510);
nand U999 (N_999,In_661,In_517);
and U1000 (N_1000,N_691,N_296);
or U1001 (N_1001,N_736,N_857);
nand U1002 (N_1002,N_954,N_340);
and U1003 (N_1003,N_336,N_256);
or U1004 (N_1004,N_908,N_990);
nor U1005 (N_1005,N_612,N_593);
and U1006 (N_1006,N_155,N_659);
or U1007 (N_1007,N_871,N_700);
nor U1008 (N_1008,N_530,N_166);
nor U1009 (N_1009,N_280,N_828);
and U1010 (N_1010,N_348,N_709);
or U1011 (N_1011,N_764,N_727);
nor U1012 (N_1012,N_360,N_257);
or U1013 (N_1013,N_672,N_290);
nand U1014 (N_1014,N_670,N_345);
nand U1015 (N_1015,N_852,N_146);
nand U1016 (N_1016,N_886,N_883);
or U1017 (N_1017,N_416,N_689);
or U1018 (N_1018,N_29,N_654);
and U1019 (N_1019,N_497,N_765);
or U1020 (N_1020,N_832,N_442);
nor U1021 (N_1021,N_59,N_71);
and U1022 (N_1022,N_374,N_815);
or U1023 (N_1023,N_353,N_979);
and U1024 (N_1024,N_65,N_434);
and U1025 (N_1025,N_826,N_321);
or U1026 (N_1026,N_669,N_112);
and U1027 (N_1027,N_568,N_113);
and U1028 (N_1028,N_77,N_724);
nor U1029 (N_1029,N_680,N_238);
or U1030 (N_1030,N_314,N_437);
and U1031 (N_1031,N_362,N_817);
nand U1032 (N_1032,N_732,N_159);
or U1033 (N_1033,N_465,N_474);
nor U1034 (N_1034,N_897,N_705);
and U1035 (N_1035,N_236,N_748);
and U1036 (N_1036,N_911,N_658);
nor U1037 (N_1037,N_754,N_295);
nand U1038 (N_1038,N_119,N_310);
nor U1039 (N_1039,N_60,N_17);
nand U1040 (N_1040,N_190,N_618);
and U1041 (N_1041,N_508,N_140);
xnor U1042 (N_1042,N_68,N_169);
and U1043 (N_1043,N_436,N_781);
nand U1044 (N_1044,N_377,N_453);
and U1045 (N_1045,N_116,N_164);
nand U1046 (N_1046,N_821,N_619);
nor U1047 (N_1047,N_745,N_307);
or U1048 (N_1048,N_933,N_779);
and U1049 (N_1049,N_10,N_513);
or U1050 (N_1050,N_484,N_992);
or U1051 (N_1051,N_70,N_837);
or U1052 (N_1052,N_585,N_414);
and U1053 (N_1053,N_786,N_952);
nor U1054 (N_1054,N_961,N_565);
or U1055 (N_1055,N_291,N_981);
or U1056 (N_1056,N_989,N_167);
nand U1057 (N_1057,N_872,N_531);
and U1058 (N_1058,N_186,N_99);
and U1059 (N_1059,N_664,N_389);
nor U1060 (N_1060,N_865,N_249);
nand U1061 (N_1061,N_46,N_48);
or U1062 (N_1062,N_413,N_40);
and U1063 (N_1063,N_163,N_793);
nor U1064 (N_1064,N_873,N_608);
and U1065 (N_1065,N_763,N_673);
nand U1066 (N_1066,N_197,N_762);
and U1067 (N_1067,N_639,N_769);
nand U1068 (N_1068,N_429,N_556);
nor U1069 (N_1069,N_827,N_583);
or U1070 (N_1070,N_239,N_549);
or U1071 (N_1071,N_675,N_785);
nor U1072 (N_1072,N_546,N_797);
or U1073 (N_1073,N_304,N_8);
nand U1074 (N_1074,N_835,N_807);
and U1075 (N_1075,N_199,N_423);
and U1076 (N_1076,N_7,N_312);
or U1077 (N_1077,N_2,N_853);
or U1078 (N_1078,N_634,N_635);
nor U1079 (N_1079,N_20,N_172);
or U1080 (N_1080,N_25,N_544);
nand U1081 (N_1081,N_35,N_766);
nor U1082 (N_1082,N_175,N_253);
nand U1083 (N_1083,N_373,N_428);
and U1084 (N_1084,N_333,N_346);
nor U1085 (N_1085,N_461,N_581);
nor U1086 (N_1086,N_882,N_927);
or U1087 (N_1087,N_126,N_720);
or U1088 (N_1088,N_219,N_301);
nor U1089 (N_1089,N_616,N_161);
nor U1090 (N_1090,N_445,N_722);
nand U1091 (N_1091,N_569,N_642);
or U1092 (N_1092,N_144,N_114);
and U1093 (N_1093,N_36,N_802);
nand U1094 (N_1094,N_127,N_212);
nand U1095 (N_1095,N_452,N_316);
or U1096 (N_1096,N_468,N_196);
nand U1097 (N_1097,N_884,N_814);
nand U1098 (N_1098,N_214,N_137);
or U1099 (N_1099,N_305,N_363);
nor U1100 (N_1100,N_129,N_912);
or U1101 (N_1101,N_647,N_730);
or U1102 (N_1102,N_154,N_225);
or U1103 (N_1103,N_274,N_630);
and U1104 (N_1104,N_498,N_610);
or U1105 (N_1105,N_187,N_838);
nand U1106 (N_1106,N_152,N_517);
nand U1107 (N_1107,N_412,N_607);
nand U1108 (N_1108,N_715,N_139);
and U1109 (N_1109,N_939,N_157);
and U1110 (N_1110,N_868,N_455);
or U1111 (N_1111,N_731,N_209);
nor U1112 (N_1112,N_261,N_358);
and U1113 (N_1113,N_796,N_105);
or U1114 (N_1114,N_276,N_767);
nor U1115 (N_1115,N_877,N_458);
nor U1116 (N_1116,N_601,N_859);
or U1117 (N_1117,N_842,N_170);
nor U1118 (N_1118,N_171,N_582);
xnor U1119 (N_1119,N_231,N_875);
nor U1120 (N_1120,N_79,N_904);
nand U1121 (N_1121,N_539,N_75);
nand U1122 (N_1122,N_491,N_393);
and U1123 (N_1123,N_486,N_289);
and U1124 (N_1124,N_52,N_138);
or U1125 (N_1125,N_650,N_192);
and U1126 (N_1126,N_536,N_425);
nor U1127 (N_1127,N_967,N_726);
nand U1128 (N_1128,N_391,N_831);
nor U1129 (N_1129,N_141,N_419);
or U1130 (N_1130,N_299,N_602);
or U1131 (N_1131,N_410,N_198);
or U1132 (N_1132,N_194,N_6);
or U1133 (N_1133,N_179,N_281);
nand U1134 (N_1134,N_712,N_746);
nand U1135 (N_1135,N_801,N_921);
nor U1136 (N_1136,N_646,N_782);
nor U1137 (N_1137,N_266,N_790);
nor U1138 (N_1138,N_120,N_302);
and U1139 (N_1139,N_205,N_522);
nor U1140 (N_1140,N_799,N_101);
nand U1141 (N_1141,N_660,N_328);
and U1142 (N_1142,N_207,N_394);
nand U1143 (N_1143,N_621,N_791);
nor U1144 (N_1144,N_311,N_824);
or U1145 (N_1145,N_996,N_264);
or U1146 (N_1146,N_400,N_469);
or U1147 (N_1147,N_697,N_991);
nor U1148 (N_1148,N_218,N_858);
nand U1149 (N_1149,N_938,N_822);
nor U1150 (N_1150,N_507,N_648);
or U1151 (N_1151,N_645,N_665);
nand U1152 (N_1152,N_854,N_788);
nand U1153 (N_1153,N_655,N_994);
nand U1154 (N_1154,N_11,N_719);
and U1155 (N_1155,N_232,N_477);
nor U1156 (N_1156,N_624,N_255);
nor U1157 (N_1157,N_955,N_269);
and U1158 (N_1158,N_1,N_623);
nand U1159 (N_1159,N_337,N_37);
or U1160 (N_1160,N_287,N_846);
nor U1161 (N_1161,N_331,N_13);
nor U1162 (N_1162,N_43,N_923);
nand U1163 (N_1163,N_576,N_64);
and U1164 (N_1164,N_557,N_999);
and U1165 (N_1165,N_87,N_133);
or U1166 (N_1166,N_118,N_433);
nand U1167 (N_1167,N_690,N_751);
or U1168 (N_1168,N_258,N_243);
or U1169 (N_1169,N_351,N_446);
or U1170 (N_1170,N_149,N_956);
and U1171 (N_1171,N_512,N_403);
nand U1172 (N_1172,N_158,N_472);
nand U1173 (N_1173,N_386,N_834);
or U1174 (N_1174,N_267,N_696);
nand U1175 (N_1175,N_251,N_860);
and U1176 (N_1176,N_605,N_866);
nor U1177 (N_1177,N_756,N_338);
nand U1178 (N_1178,N_183,N_739);
or U1179 (N_1179,N_698,N_687);
nor U1180 (N_1180,N_679,N_57);
nand U1181 (N_1181,N_203,N_117);
nor U1182 (N_1182,N_734,N_851);
nor U1183 (N_1183,N_339,N_550);
nor U1184 (N_1184,N_496,N_711);
and U1185 (N_1185,N_561,N_298);
nand U1186 (N_1186,N_24,N_368);
or U1187 (N_1187,N_109,N_747);
or U1188 (N_1188,N_110,N_547);
nand U1189 (N_1189,N_622,N_843);
nand U1190 (N_1190,N_957,N_663);
or U1191 (N_1191,N_81,N_603);
or U1192 (N_1192,N_111,N_326);
nor U1193 (N_1193,N_702,N_356);
or U1194 (N_1194,N_986,N_833);
nor U1195 (N_1195,N_44,N_916);
or U1196 (N_1196,N_143,N_88);
nor U1197 (N_1197,N_968,N_153);
and U1198 (N_1198,N_392,N_935);
nand U1199 (N_1199,N_626,N_604);
or U1200 (N_1200,N_589,N_228);
nor U1201 (N_1201,N_847,N_534);
or U1202 (N_1202,N_580,N_27);
and U1203 (N_1203,N_692,N_643);
or U1204 (N_1204,N_819,N_401);
nand U1205 (N_1205,N_188,N_708);
and U1206 (N_1206,N_804,N_347);
or U1207 (N_1207,N_502,N_638);
nand U1208 (N_1208,N_735,N_733);
and U1209 (N_1209,N_685,N_949);
and U1210 (N_1210,N_9,N_876);
nor U1211 (N_1211,N_361,N_716);
nor U1212 (N_1212,N_49,N_103);
and U1213 (N_1213,N_315,N_424);
nor U1214 (N_1214,N_760,N_202);
or U1215 (N_1215,N_344,N_93);
and U1216 (N_1216,N_84,N_910);
or U1217 (N_1217,N_511,N_600);
nand U1218 (N_1218,N_591,N_850);
or U1219 (N_1219,N_867,N_409);
and U1220 (N_1220,N_844,N_62);
nor U1221 (N_1221,N_275,N_753);
or U1222 (N_1222,N_382,N_805);
nand U1223 (N_1223,N_572,N_430);
or U1224 (N_1224,N_743,N_30);
nor U1225 (N_1225,N_217,N_879);
or U1226 (N_1226,N_470,N_278);
or U1227 (N_1227,N_548,N_984);
and U1228 (N_1228,N_324,N_222);
or U1229 (N_1229,N_926,N_123);
and U1230 (N_1230,N_946,N_463);
and U1231 (N_1231,N_271,N_542);
or U1232 (N_1232,N_628,N_95);
nor U1233 (N_1233,N_620,N_718);
nand U1234 (N_1234,N_778,N_893);
or U1235 (N_1235,N_3,N_829);
or U1236 (N_1236,N_150,N_878);
nand U1237 (N_1237,N_662,N_66);
nand U1238 (N_1238,N_651,N_862);
and U1239 (N_1239,N_951,N_447);
and U1240 (N_1240,N_761,N_206);
nor U1241 (N_1241,N_554,N_282);
or U1242 (N_1242,N_487,N_880);
nor U1243 (N_1243,N_941,N_841);
and U1244 (N_1244,N_334,N_518);
or U1245 (N_1245,N_286,N_263);
nor U1246 (N_1246,N_869,N_519);
and U1247 (N_1247,N_0,N_555);
nand U1248 (N_1248,N_825,N_595);
nor U1249 (N_1249,N_122,N_124);
or U1250 (N_1250,N_38,N_421);
or U1251 (N_1251,N_320,N_365);
nand U1252 (N_1252,N_96,N_988);
nor U1253 (N_1253,N_76,N_578);
nand U1254 (N_1254,N_980,N_586);
or U1255 (N_1255,N_323,N_970);
and U1256 (N_1256,N_641,N_388);
or U1257 (N_1257,N_740,N_381);
nand U1258 (N_1258,N_744,N_372);
nand U1259 (N_1259,N_693,N_390);
and U1260 (N_1260,N_246,N_840);
nor U1261 (N_1261,N_224,N_142);
nand U1262 (N_1262,N_737,N_772);
nor U1263 (N_1263,N_537,N_467);
nand U1264 (N_1264,N_184,N_631);
nor U1265 (N_1265,N_770,N_349);
or U1266 (N_1266,N_915,N_579);
nand U1267 (N_1267,N_242,N_402);
nand U1268 (N_1268,N_783,N_115);
nand U1269 (N_1269,N_245,N_566);
or U1270 (N_1270,N_73,N_83);
nor U1271 (N_1271,N_695,N_703);
nor U1272 (N_1272,N_63,N_803);
nor U1273 (N_1273,N_776,N_350);
nor U1274 (N_1274,N_473,N_792);
nand U1275 (N_1275,N_758,N_335);
and U1276 (N_1276,N_962,N_478);
nor U1277 (N_1277,N_969,N_535);
nor U1278 (N_1278,N_812,N_454);
nand U1279 (N_1279,N_451,N_584);
nor U1280 (N_1280,N_395,N_864);
nand U1281 (N_1281,N_406,N_268);
nor U1282 (N_1282,N_293,N_900);
and U1283 (N_1283,N_592,N_182);
or U1284 (N_1284,N_247,N_431);
xor U1285 (N_1285,N_42,N_676);
nand U1286 (N_1286,N_924,N_890);
nand U1287 (N_1287,N_449,N_914);
and U1288 (N_1288,N_714,N_47);
or U1289 (N_1289,N_919,N_490);
or U1290 (N_1290,N_818,N_270);
and U1291 (N_1291,N_907,N_525);
xnor U1292 (N_1292,N_930,N_456);
or U1293 (N_1293,N_493,N_12);
and U1294 (N_1294,N_283,N_387);
or U1295 (N_1295,N_252,N_235);
xnor U1296 (N_1296,N_541,N_435);
nor U1297 (N_1297,N_977,N_678);
and U1298 (N_1298,N_19,N_272);
and U1299 (N_1299,N_504,N_148);
or U1300 (N_1300,N_376,N_396);
or U1301 (N_1301,N_789,N_427);
and U1302 (N_1302,N_317,N_925);
xor U1303 (N_1303,N_405,N_173);
or U1304 (N_1304,N_599,N_855);
xor U1305 (N_1305,N_520,N_983);
nand U1306 (N_1306,N_699,N_755);
and U1307 (N_1307,N_237,N_902);
nor U1308 (N_1308,N_78,N_964);
nand U1309 (N_1309,N_404,N_516);
nand U1310 (N_1310,N_160,N_614);
or U1311 (N_1311,N_909,N_810);
and U1312 (N_1312,N_514,N_459);
or U1313 (N_1313,N_370,N_521);
nand U1314 (N_1314,N_553,N_21);
nor U1315 (N_1315,N_637,N_944);
and U1316 (N_1316,N_495,N_411);
nand U1317 (N_1317,N_313,N_891);
nor U1318 (N_1318,N_885,N_359);
and U1319 (N_1319,N_809,N_178);
nor U1320 (N_1320,N_422,N_971);
nor U1321 (N_1321,N_613,N_342);
nor U1322 (N_1322,N_378,N_54);
nor U1323 (N_1323,N_899,N_777);
or U1324 (N_1324,N_426,N_707);
or U1325 (N_1325,N_575,N_125);
or U1326 (N_1326,N_993,N_713);
nor U1327 (N_1327,N_367,N_108);
nand U1328 (N_1328,N_471,N_527);
nand U1329 (N_1329,N_505,N_509);
and U1330 (N_1330,N_438,N_784);
and U1331 (N_1331,N_227,N_440);
or U1332 (N_1332,N_757,N_917);
and U1333 (N_1333,N_901,N_32);
and U1334 (N_1334,N_398,N_50);
and U1335 (N_1335,N_657,N_67);
or U1336 (N_1336,N_895,N_92);
nor U1337 (N_1337,N_51,N_482);
nand U1338 (N_1338,N_611,N_545);
nor U1339 (N_1339,N_723,N_432);
and U1340 (N_1340,N_987,N_501);
nand U1341 (N_1341,N_942,N_627);
and U1342 (N_1342,N_538,N_98);
nor U1343 (N_1343,N_168,N_318);
xor U1344 (N_1344,N_948,N_773);
nand U1345 (N_1345,N_4,N_573);
nor U1346 (N_1346,N_997,N_976);
or U1347 (N_1347,N_800,N_259);
or U1348 (N_1348,N_649,N_947);
nor U1349 (N_1349,N_288,N_982);
and U1350 (N_1350,N_375,N_384);
nor U1351 (N_1351,N_870,N_364);
nand U1352 (N_1352,N_823,N_151);
xnor U1353 (N_1353,N_450,N_798);
nor U1354 (N_1354,N_352,N_226);
nand U1355 (N_1355,N_552,N_479);
and U1356 (N_1356,N_683,N_540);
and U1357 (N_1357,N_500,N_606);
and U1358 (N_1358,N_932,N_510);
or U1359 (N_1359,N_667,N_366);
nor U1360 (N_1360,N_972,N_562);
or U1361 (N_1361,N_806,N_617);
nor U1362 (N_1362,N_906,N_262);
nor U1363 (N_1363,N_371,N_418);
and U1364 (N_1364,N_845,N_330);
and U1365 (N_1365,N_597,N_343);
and U1366 (N_1366,N_567,N_889);
and U1367 (N_1367,N_574,N_185);
or U1368 (N_1368,N_128,N_441);
and U1369 (N_1369,N_5,N_380);
and U1370 (N_1370,N_590,N_529);
and U1371 (N_1371,N_250,N_85);
nor U1372 (N_1372,N_913,N_480);
or U1373 (N_1373,N_811,N_201);
or U1374 (N_1374,N_145,N_922);
nand U1375 (N_1375,N_625,N_265);
nand U1376 (N_1376,N_355,N_640);
and U1377 (N_1377,N_559,N_959);
or U1378 (N_1378,N_230,N_849);
nor U1379 (N_1379,N_56,N_920);
or U1380 (N_1380,N_39,N_26);
or U1381 (N_1381,N_45,N_162);
and U1382 (N_1382,N_515,N_684);
and U1383 (N_1383,N_407,N_41);
nor U1384 (N_1384,N_577,N_725);
nor U1385 (N_1385,N_974,N_180);
nor U1386 (N_1386,N_80,N_874);
or U1387 (N_1387,N_457,N_200);
and U1388 (N_1388,N_966,N_89);
nor U1389 (N_1389,N_379,N_503);
and U1390 (N_1390,N_945,N_587);
nand U1391 (N_1391,N_998,N_466);
and U1392 (N_1392,N_958,N_571);
or U1393 (N_1393,N_18,N_694);
nor U1394 (N_1394,N_813,N_195);
nand U1395 (N_1395,N_551,N_830);
nand U1396 (N_1396,N_905,N_294);
or U1397 (N_1397,N_357,N_385);
and U1398 (N_1398,N_488,N_856);
nor U1399 (N_1399,N_609,N_934);
nor U1400 (N_1400,N_420,N_681);
nand U1401 (N_1401,N_327,N_615);
and U1402 (N_1402,N_668,N_74);
or U1403 (N_1403,N_448,N_848);
nor U1404 (N_1404,N_808,N_863);
nand U1405 (N_1405,N_960,N_701);
or U1406 (N_1406,N_91,N_965);
or U1407 (N_1407,N_894,N_896);
and U1408 (N_1408,N_729,N_963);
nor U1409 (N_1409,N_55,N_629);
and U1410 (N_1410,N_706,N_444);
or U1411 (N_1411,N_686,N_943);
nand U1412 (N_1412,N_929,N_306);
nand U1413 (N_1413,N_973,N_774);
nand U1414 (N_1414,N_775,N_653);
nand U1415 (N_1415,N_903,N_644);
nor U1416 (N_1416,N_309,N_558);
nor U1417 (N_1417,N_666,N_97);
nor U1418 (N_1418,N_260,N_53);
xor U1419 (N_1419,N_759,N_292);
or U1420 (N_1420,N_107,N_594);
nor U1421 (N_1421,N_526,N_717);
or U1422 (N_1422,N_887,N_369);
and U1423 (N_1423,N_134,N_28);
nor U1424 (N_1424,N_241,N_652);
nand U1425 (N_1425,N_839,N_329);
nand U1426 (N_1426,N_240,N_216);
and U1427 (N_1427,N_147,N_995);
nand U1428 (N_1428,N_978,N_499);
and U1429 (N_1429,N_279,N_90);
or U1430 (N_1430,N_688,N_397);
or U1431 (N_1431,N_254,N_898);
nand U1432 (N_1432,N_485,N_588);
nand U1433 (N_1433,N_383,N_165);
nor U1434 (N_1434,N_728,N_415);
nor U1435 (N_1435,N_322,N_234);
nor U1436 (N_1436,N_481,N_524);
or U1437 (N_1437,N_771,N_928);
or U1438 (N_1438,N_58,N_297);
and U1439 (N_1439,N_677,N_130);
and U1440 (N_1440,N_86,N_749);
and U1441 (N_1441,N_795,N_104);
and U1442 (N_1442,N_94,N_439);
or U1443 (N_1443,N_506,N_303);
and U1444 (N_1444,N_121,N_23);
nor U1445 (N_1445,N_223,N_768);
nor U1446 (N_1446,N_888,N_950);
nor U1447 (N_1447,N_752,N_273);
or U1448 (N_1448,N_820,N_636);
or U1449 (N_1449,N_156,N_931);
nor U1450 (N_1450,N_210,N_953);
and U1451 (N_1451,N_523,N_710);
nor U1452 (N_1452,N_215,N_570);
or U1453 (N_1453,N_189,N_213);
nor U1454 (N_1454,N_132,N_598);
nor U1455 (N_1455,N_674,N_31);
nor U1456 (N_1456,N_492,N_325);
and U1457 (N_1457,N_82,N_936);
nor U1458 (N_1458,N_563,N_102);
nand U1459 (N_1459,N_174,N_285);
and U1460 (N_1460,N_72,N_787);
and U1461 (N_1461,N_277,N_861);
nor U1462 (N_1462,N_354,N_671);
and U1463 (N_1463,N_16,N_308);
nor U1464 (N_1464,N_918,N_136);
and U1465 (N_1465,N_284,N_181);
nand U1466 (N_1466,N_69,N_61);
and U1467 (N_1467,N_937,N_229);
and U1468 (N_1468,N_475,N_208);
nand U1469 (N_1469,N_476,N_816);
nand U1470 (N_1470,N_221,N_443);
nand U1471 (N_1471,N_177,N_248);
or U1472 (N_1472,N_135,N_417);
nand U1473 (N_1473,N_489,N_176);
or U1474 (N_1474,N_204,N_34);
nor U1475 (N_1475,N_564,N_780);
nor U1476 (N_1476,N_211,N_191);
or U1477 (N_1477,N_682,N_483);
xor U1478 (N_1478,N_131,N_332);
or U1479 (N_1479,N_533,N_738);
nor U1480 (N_1480,N_633,N_233);
or U1481 (N_1481,N_892,N_15);
nand U1482 (N_1482,N_532,N_656);
nand U1483 (N_1483,N_106,N_14);
nor U1484 (N_1484,N_244,N_220);
nor U1485 (N_1485,N_596,N_975);
nand U1486 (N_1486,N_193,N_836);
or U1487 (N_1487,N_794,N_408);
nand U1488 (N_1488,N_462,N_528);
or U1489 (N_1489,N_881,N_742);
nand U1490 (N_1490,N_985,N_399);
or U1491 (N_1491,N_464,N_741);
nand U1492 (N_1492,N_33,N_460);
nand U1493 (N_1493,N_300,N_341);
or U1494 (N_1494,N_704,N_543);
nand U1495 (N_1495,N_661,N_319);
nand U1496 (N_1496,N_494,N_100);
and U1497 (N_1497,N_750,N_22);
or U1498 (N_1498,N_940,N_632);
and U1499 (N_1499,N_560,N_721);
and U1500 (N_1500,N_696,N_343);
and U1501 (N_1501,N_661,N_739);
and U1502 (N_1502,N_341,N_364);
nand U1503 (N_1503,N_430,N_394);
or U1504 (N_1504,N_953,N_464);
and U1505 (N_1505,N_78,N_634);
nand U1506 (N_1506,N_422,N_646);
nor U1507 (N_1507,N_201,N_700);
and U1508 (N_1508,N_483,N_589);
or U1509 (N_1509,N_56,N_441);
and U1510 (N_1510,N_940,N_447);
and U1511 (N_1511,N_992,N_309);
nor U1512 (N_1512,N_498,N_147);
and U1513 (N_1513,N_603,N_200);
nor U1514 (N_1514,N_268,N_255);
nor U1515 (N_1515,N_944,N_591);
nand U1516 (N_1516,N_87,N_263);
or U1517 (N_1517,N_870,N_234);
nor U1518 (N_1518,N_993,N_222);
or U1519 (N_1519,N_804,N_518);
nor U1520 (N_1520,N_402,N_309);
nand U1521 (N_1521,N_212,N_458);
nor U1522 (N_1522,N_181,N_601);
nand U1523 (N_1523,N_894,N_547);
and U1524 (N_1524,N_257,N_982);
nand U1525 (N_1525,N_68,N_209);
nor U1526 (N_1526,N_55,N_129);
and U1527 (N_1527,N_76,N_146);
nor U1528 (N_1528,N_980,N_607);
xor U1529 (N_1529,N_428,N_721);
or U1530 (N_1530,N_520,N_421);
nor U1531 (N_1531,N_974,N_949);
nand U1532 (N_1532,N_284,N_530);
nor U1533 (N_1533,N_882,N_687);
nand U1534 (N_1534,N_318,N_396);
nand U1535 (N_1535,N_961,N_665);
nand U1536 (N_1536,N_822,N_199);
and U1537 (N_1537,N_204,N_385);
and U1538 (N_1538,N_879,N_488);
nor U1539 (N_1539,N_330,N_65);
nor U1540 (N_1540,N_886,N_643);
nor U1541 (N_1541,N_577,N_72);
nor U1542 (N_1542,N_130,N_162);
and U1543 (N_1543,N_711,N_411);
nor U1544 (N_1544,N_472,N_402);
or U1545 (N_1545,N_218,N_805);
and U1546 (N_1546,N_699,N_570);
and U1547 (N_1547,N_65,N_172);
and U1548 (N_1548,N_252,N_788);
or U1549 (N_1549,N_696,N_446);
or U1550 (N_1550,N_150,N_303);
or U1551 (N_1551,N_584,N_974);
nor U1552 (N_1552,N_555,N_746);
nand U1553 (N_1553,N_512,N_151);
or U1554 (N_1554,N_325,N_731);
or U1555 (N_1555,N_86,N_106);
and U1556 (N_1556,N_517,N_275);
nor U1557 (N_1557,N_36,N_271);
nand U1558 (N_1558,N_146,N_889);
nand U1559 (N_1559,N_746,N_871);
nor U1560 (N_1560,N_604,N_245);
or U1561 (N_1561,N_951,N_390);
and U1562 (N_1562,N_892,N_735);
and U1563 (N_1563,N_199,N_591);
nor U1564 (N_1564,N_30,N_225);
and U1565 (N_1565,N_95,N_265);
nor U1566 (N_1566,N_81,N_279);
nor U1567 (N_1567,N_431,N_893);
and U1568 (N_1568,N_774,N_939);
or U1569 (N_1569,N_756,N_43);
nand U1570 (N_1570,N_304,N_695);
or U1571 (N_1571,N_824,N_722);
or U1572 (N_1572,N_221,N_985);
nand U1573 (N_1573,N_743,N_77);
and U1574 (N_1574,N_244,N_468);
and U1575 (N_1575,N_529,N_526);
nor U1576 (N_1576,N_315,N_556);
and U1577 (N_1577,N_467,N_560);
or U1578 (N_1578,N_275,N_547);
nand U1579 (N_1579,N_981,N_36);
and U1580 (N_1580,N_190,N_144);
or U1581 (N_1581,N_635,N_16);
or U1582 (N_1582,N_535,N_86);
and U1583 (N_1583,N_661,N_567);
or U1584 (N_1584,N_758,N_647);
or U1585 (N_1585,N_425,N_712);
or U1586 (N_1586,N_470,N_435);
nand U1587 (N_1587,N_616,N_456);
nand U1588 (N_1588,N_456,N_924);
nand U1589 (N_1589,N_656,N_510);
nor U1590 (N_1590,N_612,N_960);
or U1591 (N_1591,N_695,N_891);
nor U1592 (N_1592,N_803,N_810);
nor U1593 (N_1593,N_159,N_550);
or U1594 (N_1594,N_396,N_505);
nor U1595 (N_1595,N_963,N_215);
and U1596 (N_1596,N_306,N_372);
and U1597 (N_1597,N_627,N_326);
and U1598 (N_1598,N_376,N_57);
and U1599 (N_1599,N_284,N_429);
and U1600 (N_1600,N_175,N_842);
nor U1601 (N_1601,N_395,N_504);
or U1602 (N_1602,N_56,N_178);
nand U1603 (N_1603,N_365,N_256);
nor U1604 (N_1604,N_532,N_3);
and U1605 (N_1605,N_934,N_265);
nand U1606 (N_1606,N_724,N_366);
and U1607 (N_1607,N_949,N_130);
and U1608 (N_1608,N_325,N_526);
and U1609 (N_1609,N_178,N_618);
xnor U1610 (N_1610,N_79,N_762);
nor U1611 (N_1611,N_67,N_176);
or U1612 (N_1612,N_338,N_532);
nor U1613 (N_1613,N_307,N_80);
nor U1614 (N_1614,N_398,N_712);
and U1615 (N_1615,N_79,N_191);
nor U1616 (N_1616,N_680,N_794);
and U1617 (N_1617,N_570,N_939);
nand U1618 (N_1618,N_977,N_553);
or U1619 (N_1619,N_643,N_459);
nand U1620 (N_1620,N_181,N_226);
nand U1621 (N_1621,N_613,N_467);
nor U1622 (N_1622,N_251,N_718);
and U1623 (N_1623,N_957,N_283);
nor U1624 (N_1624,N_293,N_97);
and U1625 (N_1625,N_667,N_503);
nor U1626 (N_1626,N_170,N_934);
nand U1627 (N_1627,N_845,N_656);
or U1628 (N_1628,N_839,N_958);
nand U1629 (N_1629,N_855,N_46);
and U1630 (N_1630,N_687,N_223);
and U1631 (N_1631,N_531,N_647);
or U1632 (N_1632,N_81,N_46);
or U1633 (N_1633,N_825,N_728);
nand U1634 (N_1634,N_755,N_299);
or U1635 (N_1635,N_117,N_369);
nand U1636 (N_1636,N_624,N_23);
or U1637 (N_1637,N_106,N_547);
or U1638 (N_1638,N_21,N_540);
or U1639 (N_1639,N_859,N_519);
nor U1640 (N_1640,N_356,N_958);
nor U1641 (N_1641,N_795,N_53);
and U1642 (N_1642,N_710,N_992);
nor U1643 (N_1643,N_480,N_291);
nand U1644 (N_1644,N_524,N_683);
and U1645 (N_1645,N_488,N_105);
nor U1646 (N_1646,N_558,N_927);
and U1647 (N_1647,N_293,N_477);
nand U1648 (N_1648,N_619,N_891);
nand U1649 (N_1649,N_527,N_360);
nor U1650 (N_1650,N_50,N_176);
and U1651 (N_1651,N_863,N_739);
nor U1652 (N_1652,N_568,N_414);
nor U1653 (N_1653,N_927,N_401);
or U1654 (N_1654,N_173,N_705);
or U1655 (N_1655,N_172,N_215);
nor U1656 (N_1656,N_290,N_441);
and U1657 (N_1657,N_225,N_720);
nor U1658 (N_1658,N_651,N_691);
nor U1659 (N_1659,N_838,N_80);
nand U1660 (N_1660,N_848,N_598);
nor U1661 (N_1661,N_441,N_421);
or U1662 (N_1662,N_116,N_641);
nor U1663 (N_1663,N_407,N_860);
or U1664 (N_1664,N_840,N_713);
or U1665 (N_1665,N_277,N_700);
or U1666 (N_1666,N_640,N_233);
nand U1667 (N_1667,N_465,N_577);
or U1668 (N_1668,N_498,N_388);
and U1669 (N_1669,N_597,N_15);
or U1670 (N_1670,N_637,N_23);
nor U1671 (N_1671,N_740,N_345);
and U1672 (N_1672,N_10,N_586);
nor U1673 (N_1673,N_184,N_967);
and U1674 (N_1674,N_22,N_68);
nand U1675 (N_1675,N_790,N_472);
nand U1676 (N_1676,N_309,N_990);
or U1677 (N_1677,N_929,N_397);
nor U1678 (N_1678,N_118,N_925);
nand U1679 (N_1679,N_270,N_382);
or U1680 (N_1680,N_734,N_892);
nor U1681 (N_1681,N_550,N_43);
nor U1682 (N_1682,N_827,N_792);
and U1683 (N_1683,N_995,N_62);
or U1684 (N_1684,N_49,N_642);
or U1685 (N_1685,N_293,N_994);
or U1686 (N_1686,N_782,N_665);
nor U1687 (N_1687,N_640,N_538);
or U1688 (N_1688,N_147,N_520);
or U1689 (N_1689,N_689,N_548);
nor U1690 (N_1690,N_570,N_634);
and U1691 (N_1691,N_601,N_459);
nand U1692 (N_1692,N_465,N_618);
nor U1693 (N_1693,N_31,N_225);
and U1694 (N_1694,N_713,N_851);
nor U1695 (N_1695,N_435,N_368);
nor U1696 (N_1696,N_411,N_187);
nand U1697 (N_1697,N_217,N_986);
or U1698 (N_1698,N_757,N_906);
nor U1699 (N_1699,N_235,N_780);
or U1700 (N_1700,N_260,N_551);
nor U1701 (N_1701,N_395,N_207);
nor U1702 (N_1702,N_982,N_486);
and U1703 (N_1703,N_271,N_831);
or U1704 (N_1704,N_423,N_583);
nand U1705 (N_1705,N_299,N_495);
nand U1706 (N_1706,N_583,N_189);
nand U1707 (N_1707,N_128,N_423);
and U1708 (N_1708,N_655,N_786);
nor U1709 (N_1709,N_935,N_696);
and U1710 (N_1710,N_822,N_352);
nor U1711 (N_1711,N_877,N_923);
nand U1712 (N_1712,N_518,N_406);
or U1713 (N_1713,N_112,N_524);
nand U1714 (N_1714,N_131,N_413);
or U1715 (N_1715,N_891,N_83);
nand U1716 (N_1716,N_457,N_786);
nand U1717 (N_1717,N_68,N_435);
or U1718 (N_1718,N_0,N_373);
and U1719 (N_1719,N_829,N_715);
or U1720 (N_1720,N_204,N_81);
and U1721 (N_1721,N_608,N_557);
and U1722 (N_1722,N_242,N_601);
xor U1723 (N_1723,N_645,N_406);
or U1724 (N_1724,N_995,N_322);
or U1725 (N_1725,N_641,N_838);
and U1726 (N_1726,N_814,N_23);
or U1727 (N_1727,N_462,N_724);
nand U1728 (N_1728,N_133,N_319);
and U1729 (N_1729,N_667,N_229);
and U1730 (N_1730,N_825,N_379);
and U1731 (N_1731,N_876,N_70);
nor U1732 (N_1732,N_205,N_548);
nor U1733 (N_1733,N_529,N_492);
and U1734 (N_1734,N_714,N_453);
nand U1735 (N_1735,N_133,N_458);
or U1736 (N_1736,N_518,N_499);
nor U1737 (N_1737,N_111,N_122);
nor U1738 (N_1738,N_694,N_913);
or U1739 (N_1739,N_921,N_415);
nand U1740 (N_1740,N_641,N_5);
nand U1741 (N_1741,N_216,N_832);
nor U1742 (N_1742,N_40,N_396);
nand U1743 (N_1743,N_905,N_228);
or U1744 (N_1744,N_708,N_812);
or U1745 (N_1745,N_166,N_118);
nor U1746 (N_1746,N_854,N_566);
nand U1747 (N_1747,N_577,N_986);
nor U1748 (N_1748,N_371,N_795);
or U1749 (N_1749,N_805,N_821);
or U1750 (N_1750,N_736,N_206);
or U1751 (N_1751,N_509,N_257);
nor U1752 (N_1752,N_268,N_202);
and U1753 (N_1753,N_100,N_936);
nor U1754 (N_1754,N_164,N_404);
or U1755 (N_1755,N_851,N_698);
nor U1756 (N_1756,N_141,N_104);
nand U1757 (N_1757,N_207,N_844);
or U1758 (N_1758,N_565,N_20);
and U1759 (N_1759,N_764,N_162);
and U1760 (N_1760,N_150,N_672);
or U1761 (N_1761,N_103,N_153);
and U1762 (N_1762,N_902,N_669);
nand U1763 (N_1763,N_585,N_962);
nand U1764 (N_1764,N_91,N_594);
nor U1765 (N_1765,N_545,N_36);
nand U1766 (N_1766,N_156,N_568);
or U1767 (N_1767,N_724,N_509);
or U1768 (N_1768,N_631,N_173);
and U1769 (N_1769,N_758,N_612);
nor U1770 (N_1770,N_199,N_90);
and U1771 (N_1771,N_131,N_716);
nand U1772 (N_1772,N_269,N_759);
and U1773 (N_1773,N_882,N_761);
and U1774 (N_1774,N_649,N_228);
nand U1775 (N_1775,N_864,N_325);
nor U1776 (N_1776,N_969,N_863);
nor U1777 (N_1777,N_793,N_338);
nand U1778 (N_1778,N_807,N_648);
and U1779 (N_1779,N_197,N_152);
and U1780 (N_1780,N_858,N_245);
nand U1781 (N_1781,N_459,N_597);
or U1782 (N_1782,N_470,N_379);
and U1783 (N_1783,N_373,N_662);
nand U1784 (N_1784,N_131,N_494);
nand U1785 (N_1785,N_829,N_77);
nor U1786 (N_1786,N_177,N_984);
or U1787 (N_1787,N_922,N_499);
or U1788 (N_1788,N_152,N_507);
nor U1789 (N_1789,N_545,N_47);
nand U1790 (N_1790,N_789,N_324);
and U1791 (N_1791,N_560,N_670);
or U1792 (N_1792,N_408,N_353);
or U1793 (N_1793,N_80,N_359);
nand U1794 (N_1794,N_315,N_583);
or U1795 (N_1795,N_665,N_71);
nor U1796 (N_1796,N_733,N_906);
or U1797 (N_1797,N_346,N_665);
or U1798 (N_1798,N_229,N_711);
and U1799 (N_1799,N_99,N_15);
or U1800 (N_1800,N_955,N_268);
or U1801 (N_1801,N_987,N_334);
or U1802 (N_1802,N_995,N_749);
nand U1803 (N_1803,N_396,N_450);
nand U1804 (N_1804,N_853,N_326);
and U1805 (N_1805,N_667,N_457);
xor U1806 (N_1806,N_420,N_482);
or U1807 (N_1807,N_584,N_131);
nor U1808 (N_1808,N_123,N_245);
or U1809 (N_1809,N_769,N_733);
or U1810 (N_1810,N_511,N_975);
and U1811 (N_1811,N_378,N_290);
nor U1812 (N_1812,N_224,N_97);
nand U1813 (N_1813,N_976,N_873);
nand U1814 (N_1814,N_198,N_88);
and U1815 (N_1815,N_678,N_796);
nor U1816 (N_1816,N_255,N_108);
or U1817 (N_1817,N_753,N_879);
nor U1818 (N_1818,N_118,N_155);
xnor U1819 (N_1819,N_510,N_998);
nor U1820 (N_1820,N_608,N_135);
or U1821 (N_1821,N_826,N_212);
and U1822 (N_1822,N_949,N_250);
nor U1823 (N_1823,N_546,N_24);
nand U1824 (N_1824,N_213,N_208);
nand U1825 (N_1825,N_986,N_331);
or U1826 (N_1826,N_794,N_264);
nor U1827 (N_1827,N_477,N_785);
nor U1828 (N_1828,N_971,N_121);
nor U1829 (N_1829,N_936,N_219);
nor U1830 (N_1830,N_418,N_771);
or U1831 (N_1831,N_847,N_615);
or U1832 (N_1832,N_472,N_295);
nand U1833 (N_1833,N_679,N_245);
nand U1834 (N_1834,N_234,N_752);
nand U1835 (N_1835,N_176,N_919);
nor U1836 (N_1836,N_707,N_209);
nor U1837 (N_1837,N_743,N_943);
nand U1838 (N_1838,N_971,N_608);
nand U1839 (N_1839,N_461,N_829);
nand U1840 (N_1840,N_894,N_159);
or U1841 (N_1841,N_459,N_267);
nor U1842 (N_1842,N_311,N_68);
nor U1843 (N_1843,N_906,N_316);
nor U1844 (N_1844,N_827,N_787);
nor U1845 (N_1845,N_397,N_180);
and U1846 (N_1846,N_872,N_173);
nand U1847 (N_1847,N_211,N_791);
nor U1848 (N_1848,N_270,N_315);
and U1849 (N_1849,N_567,N_326);
and U1850 (N_1850,N_800,N_167);
nor U1851 (N_1851,N_889,N_791);
nand U1852 (N_1852,N_606,N_816);
or U1853 (N_1853,N_63,N_989);
nor U1854 (N_1854,N_627,N_394);
or U1855 (N_1855,N_997,N_304);
nor U1856 (N_1856,N_310,N_649);
or U1857 (N_1857,N_251,N_998);
or U1858 (N_1858,N_211,N_718);
nand U1859 (N_1859,N_24,N_752);
and U1860 (N_1860,N_711,N_731);
nand U1861 (N_1861,N_93,N_684);
nand U1862 (N_1862,N_214,N_903);
nor U1863 (N_1863,N_787,N_604);
and U1864 (N_1864,N_206,N_103);
and U1865 (N_1865,N_666,N_17);
nor U1866 (N_1866,N_326,N_66);
nand U1867 (N_1867,N_278,N_737);
nand U1868 (N_1868,N_216,N_826);
or U1869 (N_1869,N_21,N_732);
and U1870 (N_1870,N_702,N_273);
nor U1871 (N_1871,N_446,N_429);
nor U1872 (N_1872,N_25,N_652);
nand U1873 (N_1873,N_143,N_68);
and U1874 (N_1874,N_122,N_501);
or U1875 (N_1875,N_327,N_570);
nand U1876 (N_1876,N_643,N_479);
nor U1877 (N_1877,N_396,N_401);
nand U1878 (N_1878,N_646,N_141);
and U1879 (N_1879,N_716,N_804);
and U1880 (N_1880,N_713,N_808);
and U1881 (N_1881,N_117,N_907);
nor U1882 (N_1882,N_947,N_445);
or U1883 (N_1883,N_868,N_36);
nor U1884 (N_1884,N_572,N_17);
nor U1885 (N_1885,N_407,N_40);
nand U1886 (N_1886,N_856,N_41);
nand U1887 (N_1887,N_17,N_728);
or U1888 (N_1888,N_875,N_609);
and U1889 (N_1889,N_461,N_788);
or U1890 (N_1890,N_485,N_286);
nor U1891 (N_1891,N_909,N_578);
or U1892 (N_1892,N_495,N_360);
nor U1893 (N_1893,N_151,N_475);
and U1894 (N_1894,N_557,N_245);
or U1895 (N_1895,N_973,N_445);
or U1896 (N_1896,N_348,N_183);
nand U1897 (N_1897,N_865,N_591);
nor U1898 (N_1898,N_602,N_669);
nor U1899 (N_1899,N_517,N_41);
nand U1900 (N_1900,N_921,N_292);
nor U1901 (N_1901,N_207,N_324);
nand U1902 (N_1902,N_319,N_713);
nand U1903 (N_1903,N_309,N_161);
or U1904 (N_1904,N_153,N_809);
or U1905 (N_1905,N_699,N_134);
nor U1906 (N_1906,N_946,N_762);
and U1907 (N_1907,N_722,N_805);
nand U1908 (N_1908,N_268,N_234);
or U1909 (N_1909,N_314,N_391);
and U1910 (N_1910,N_479,N_182);
and U1911 (N_1911,N_181,N_406);
or U1912 (N_1912,N_302,N_132);
and U1913 (N_1913,N_880,N_1);
xor U1914 (N_1914,N_620,N_181);
and U1915 (N_1915,N_890,N_619);
and U1916 (N_1916,N_899,N_45);
and U1917 (N_1917,N_934,N_742);
nor U1918 (N_1918,N_195,N_156);
nand U1919 (N_1919,N_817,N_737);
and U1920 (N_1920,N_479,N_383);
nand U1921 (N_1921,N_882,N_747);
or U1922 (N_1922,N_777,N_129);
nor U1923 (N_1923,N_337,N_51);
nor U1924 (N_1924,N_535,N_338);
and U1925 (N_1925,N_931,N_419);
nand U1926 (N_1926,N_900,N_950);
or U1927 (N_1927,N_256,N_899);
or U1928 (N_1928,N_950,N_578);
nand U1929 (N_1929,N_835,N_423);
or U1930 (N_1930,N_173,N_850);
nor U1931 (N_1931,N_331,N_805);
or U1932 (N_1932,N_890,N_187);
nand U1933 (N_1933,N_430,N_369);
nand U1934 (N_1934,N_866,N_333);
and U1935 (N_1935,N_881,N_464);
nand U1936 (N_1936,N_650,N_788);
or U1937 (N_1937,N_39,N_975);
or U1938 (N_1938,N_293,N_723);
nand U1939 (N_1939,N_2,N_322);
nand U1940 (N_1940,N_522,N_824);
and U1941 (N_1941,N_610,N_329);
nand U1942 (N_1942,N_569,N_791);
or U1943 (N_1943,N_22,N_305);
and U1944 (N_1944,N_281,N_788);
and U1945 (N_1945,N_67,N_755);
nand U1946 (N_1946,N_234,N_819);
nor U1947 (N_1947,N_788,N_435);
and U1948 (N_1948,N_863,N_790);
nand U1949 (N_1949,N_581,N_97);
and U1950 (N_1950,N_51,N_225);
or U1951 (N_1951,N_650,N_560);
nor U1952 (N_1952,N_222,N_10);
nor U1953 (N_1953,N_708,N_866);
and U1954 (N_1954,N_571,N_924);
nor U1955 (N_1955,N_59,N_633);
and U1956 (N_1956,N_627,N_915);
nand U1957 (N_1957,N_674,N_874);
nor U1958 (N_1958,N_24,N_81);
nor U1959 (N_1959,N_219,N_356);
nand U1960 (N_1960,N_223,N_751);
nand U1961 (N_1961,N_497,N_145);
or U1962 (N_1962,N_127,N_579);
and U1963 (N_1963,N_262,N_549);
or U1964 (N_1964,N_728,N_620);
and U1965 (N_1965,N_42,N_64);
and U1966 (N_1966,N_358,N_341);
and U1967 (N_1967,N_364,N_840);
nor U1968 (N_1968,N_998,N_398);
or U1969 (N_1969,N_182,N_53);
nand U1970 (N_1970,N_947,N_247);
nand U1971 (N_1971,N_632,N_894);
or U1972 (N_1972,N_891,N_645);
and U1973 (N_1973,N_311,N_200);
or U1974 (N_1974,N_635,N_614);
nor U1975 (N_1975,N_745,N_62);
nand U1976 (N_1976,N_624,N_253);
nand U1977 (N_1977,N_645,N_29);
nand U1978 (N_1978,N_530,N_77);
nand U1979 (N_1979,N_632,N_526);
or U1980 (N_1980,N_341,N_216);
nor U1981 (N_1981,N_588,N_419);
nor U1982 (N_1982,N_23,N_673);
or U1983 (N_1983,N_709,N_414);
nor U1984 (N_1984,N_171,N_237);
and U1985 (N_1985,N_388,N_292);
xor U1986 (N_1986,N_387,N_377);
or U1987 (N_1987,N_760,N_166);
nand U1988 (N_1988,N_849,N_896);
nand U1989 (N_1989,N_588,N_762);
and U1990 (N_1990,N_607,N_173);
or U1991 (N_1991,N_157,N_336);
and U1992 (N_1992,N_426,N_287);
or U1993 (N_1993,N_0,N_501);
nand U1994 (N_1994,N_802,N_0);
nor U1995 (N_1995,N_736,N_350);
nand U1996 (N_1996,N_270,N_309);
or U1997 (N_1997,N_87,N_322);
and U1998 (N_1998,N_458,N_145);
nor U1999 (N_1999,N_762,N_358);
nor U2000 (N_2000,N_1849,N_1259);
nor U2001 (N_2001,N_1710,N_1609);
or U2002 (N_2002,N_1235,N_1445);
or U2003 (N_2003,N_1157,N_1622);
or U2004 (N_2004,N_1467,N_1875);
nand U2005 (N_2005,N_1754,N_1575);
or U2006 (N_2006,N_1988,N_1471);
and U2007 (N_2007,N_1554,N_1099);
or U2008 (N_2008,N_1306,N_1000);
nor U2009 (N_2009,N_1008,N_1738);
and U2010 (N_2010,N_1568,N_1996);
nor U2011 (N_2011,N_1083,N_1185);
or U2012 (N_2012,N_1919,N_1274);
or U2013 (N_2013,N_1297,N_1705);
nand U2014 (N_2014,N_1014,N_1111);
nor U2015 (N_2015,N_1506,N_1123);
xnor U2016 (N_2016,N_1044,N_1736);
nand U2017 (N_2017,N_1908,N_1187);
and U2018 (N_2018,N_1419,N_1228);
nor U2019 (N_2019,N_1899,N_1366);
and U2020 (N_2020,N_1245,N_1217);
or U2021 (N_2021,N_1056,N_1567);
and U2022 (N_2022,N_1414,N_1986);
or U2023 (N_2023,N_1418,N_1147);
nor U2024 (N_2024,N_1329,N_1519);
or U2025 (N_2025,N_1588,N_1220);
nor U2026 (N_2026,N_1831,N_1317);
and U2027 (N_2027,N_1618,N_1648);
or U2028 (N_2028,N_1384,N_1474);
nor U2029 (N_2029,N_1520,N_1386);
and U2030 (N_2030,N_1508,N_1872);
and U2031 (N_2031,N_1053,N_1409);
or U2032 (N_2032,N_1625,N_1037);
and U2033 (N_2033,N_1624,N_1978);
nor U2034 (N_2034,N_1886,N_1861);
or U2035 (N_2035,N_1739,N_1021);
nor U2036 (N_2036,N_1019,N_1560);
and U2037 (N_2037,N_1006,N_1714);
and U2038 (N_2038,N_1837,N_1380);
or U2039 (N_2039,N_1027,N_1065);
nor U2040 (N_2040,N_1446,N_1548);
or U2041 (N_2041,N_1050,N_1197);
or U2042 (N_2042,N_1639,N_1940);
nor U2043 (N_2043,N_1815,N_1672);
and U2044 (N_2044,N_1853,N_1170);
nand U2045 (N_2045,N_1513,N_1054);
or U2046 (N_2046,N_1937,N_1312);
nor U2047 (N_2047,N_1393,N_1870);
nand U2048 (N_2048,N_1911,N_1320);
or U2049 (N_2049,N_1232,N_1289);
and U2050 (N_2050,N_1010,N_1694);
and U2051 (N_2051,N_1238,N_1135);
or U2052 (N_2052,N_1193,N_1348);
or U2053 (N_2053,N_1600,N_1150);
nand U2054 (N_2054,N_1025,N_1656);
xor U2055 (N_2055,N_1598,N_1133);
or U2056 (N_2056,N_1129,N_1449);
nand U2057 (N_2057,N_1051,N_1977);
and U2058 (N_2058,N_1401,N_1766);
and U2059 (N_2059,N_1810,N_1175);
nor U2060 (N_2060,N_1344,N_1230);
or U2061 (N_2061,N_1438,N_1042);
and U2062 (N_2062,N_1522,N_1069);
or U2063 (N_2063,N_1820,N_1173);
and U2064 (N_2064,N_1237,N_1594);
nor U2065 (N_2065,N_1347,N_1085);
nand U2066 (N_2066,N_1671,N_1106);
and U2067 (N_2067,N_1712,N_1194);
or U2068 (N_2068,N_1957,N_1140);
nor U2069 (N_2069,N_1071,N_1061);
nor U2070 (N_2070,N_1871,N_1285);
or U2071 (N_2071,N_1982,N_1523);
or U2072 (N_2072,N_1963,N_1502);
and U2073 (N_2073,N_1877,N_1336);
nor U2074 (N_2074,N_1112,N_1168);
nand U2075 (N_2075,N_1645,N_1439);
or U2076 (N_2076,N_1408,N_1234);
or U2077 (N_2077,N_1189,N_1064);
nand U2078 (N_2078,N_1435,N_1411);
or U2079 (N_2079,N_1190,N_1836);
nor U2080 (N_2080,N_1273,N_1256);
nor U2081 (N_2081,N_1587,N_1811);
and U2082 (N_2082,N_1891,N_1635);
nor U2083 (N_2083,N_1313,N_1878);
or U2084 (N_2084,N_1278,N_1149);
or U2085 (N_2085,N_1059,N_1565);
or U2086 (N_2086,N_1844,N_1751);
and U2087 (N_2087,N_1326,N_1559);
and U2088 (N_2088,N_1876,N_1487);
or U2089 (N_2089,N_1277,N_1660);
nor U2090 (N_2090,N_1678,N_1470);
nand U2091 (N_2091,N_1444,N_1379);
nor U2092 (N_2092,N_1733,N_1715);
and U2093 (N_2093,N_1492,N_1206);
nor U2094 (N_2094,N_1802,N_1131);
or U2095 (N_2095,N_1373,N_1975);
nand U2096 (N_2096,N_1698,N_1128);
or U2097 (N_2097,N_1651,N_1515);
nor U2098 (N_2098,N_1650,N_1242);
or U2099 (N_2099,N_1652,N_1001);
or U2100 (N_2100,N_1262,N_1310);
and U2101 (N_2101,N_1091,N_1400);
or U2102 (N_2102,N_1758,N_1556);
and U2103 (N_2103,N_1857,N_1130);
and U2104 (N_2104,N_1062,N_1668);
and U2105 (N_2105,N_1086,N_1354);
or U2106 (N_2106,N_1482,N_1874);
or U2107 (N_2107,N_1638,N_1774);
nor U2108 (N_2108,N_1574,N_1063);
nand U2109 (N_2109,N_1260,N_1316);
and U2110 (N_2110,N_1298,N_1103);
or U2111 (N_2111,N_1816,N_1564);
or U2112 (N_2112,N_1550,N_1785);
and U2113 (N_2113,N_1284,N_1208);
or U2114 (N_2114,N_1122,N_1304);
or U2115 (N_2115,N_1743,N_1158);
nor U2116 (N_2116,N_1395,N_1433);
nor U2117 (N_2117,N_1983,N_1180);
or U2118 (N_2118,N_1486,N_1126);
nand U2119 (N_2119,N_1015,N_1075);
and U2120 (N_2120,N_1707,N_1846);
or U2121 (N_2121,N_1729,N_1628);
and U2122 (N_2122,N_1356,N_1695);
nand U2123 (N_2123,N_1525,N_1191);
and U2124 (N_2124,N_1997,N_1457);
and U2125 (N_2125,N_1121,N_1763);
or U2126 (N_2126,N_1331,N_1361);
nor U2127 (N_2127,N_1020,N_1770);
or U2128 (N_2128,N_1301,N_1790);
and U2129 (N_2129,N_1787,N_1146);
nand U2130 (N_2130,N_1973,N_1473);
or U2131 (N_2131,N_1667,N_1167);
nand U2132 (N_2132,N_1749,N_1884);
nand U2133 (N_2133,N_1327,N_1780);
and U2134 (N_2134,N_1428,N_1458);
and U2135 (N_2135,N_1752,N_1362);
and U2136 (N_2136,N_1365,N_1782);
nor U2137 (N_2137,N_1999,N_1060);
nand U2138 (N_2138,N_1961,N_1530);
xnor U2139 (N_2139,N_1631,N_1632);
or U2140 (N_2140,N_1546,N_1499);
nor U2141 (N_2141,N_1640,N_1370);
nand U2142 (N_2142,N_1898,N_1357);
and U2143 (N_2143,N_1004,N_1082);
or U2144 (N_2144,N_1253,N_1209);
and U2145 (N_2145,N_1563,N_1935);
or U2146 (N_2146,N_1995,N_1478);
or U2147 (N_2147,N_1643,N_1674);
nor U2148 (N_2148,N_1677,N_1696);
or U2149 (N_2149,N_1324,N_1335);
nand U2150 (N_2150,N_1942,N_1906);
and U2151 (N_2151,N_1340,N_1318);
nand U2152 (N_2152,N_1547,N_1718);
or U2153 (N_2153,N_1965,N_1806);
nor U2154 (N_2154,N_1814,N_1462);
xnor U2155 (N_2155,N_1092,N_1711);
and U2156 (N_2156,N_1241,N_1646);
nand U2157 (N_2157,N_1850,N_1113);
nand U2158 (N_2158,N_1290,N_1679);
and U2159 (N_2159,N_1355,N_1504);
nor U2160 (N_2160,N_1294,N_1687);
or U2161 (N_2161,N_1440,N_1834);
and U2162 (N_2162,N_1442,N_1371);
or U2163 (N_2163,N_1862,N_1088);
or U2164 (N_2164,N_1219,N_1346);
xnor U2165 (N_2165,N_1953,N_1581);
nand U2166 (N_2166,N_1236,N_1293);
and U2167 (N_2167,N_1805,N_1102);
nand U2168 (N_2168,N_1394,N_1321);
and U2169 (N_2169,N_1453,N_1665);
nor U2170 (N_2170,N_1974,N_1521);
nand U2171 (N_2171,N_1755,N_1662);
or U2172 (N_2172,N_1532,N_1024);
and U2173 (N_2173,N_1590,N_1516);
or U2174 (N_2174,N_1697,N_1993);
nor U2175 (N_2175,N_1116,N_1583);
nor U2176 (N_2176,N_1926,N_1057);
and U2177 (N_2177,N_1510,N_1931);
nand U2178 (N_2178,N_1415,N_1930);
and U2179 (N_2179,N_1948,N_1918);
or U2180 (N_2180,N_1750,N_1726);
or U2181 (N_2181,N_1145,N_1949);
nor U2182 (N_2182,N_1903,N_1055);
nand U2183 (N_2183,N_1613,N_1552);
and U2184 (N_2184,N_1675,N_1873);
nand U2185 (N_2185,N_1566,N_1496);
nor U2186 (N_2186,N_1807,N_1270);
nand U2187 (N_2187,N_1352,N_1859);
or U2188 (N_2188,N_1860,N_1670);
and U2189 (N_2189,N_1518,N_1614);
nand U2190 (N_2190,N_1809,N_1448);
nand U2191 (N_2191,N_1136,N_1623);
nand U2192 (N_2192,N_1093,N_1866);
and U2193 (N_2193,N_1281,N_1251);
nor U2194 (N_2194,N_1704,N_1424);
or U2195 (N_2195,N_1827,N_1143);
and U2196 (N_2196,N_1562,N_1443);
nand U2197 (N_2197,N_1124,N_1781);
or U2198 (N_2198,N_1472,N_1735);
and U2199 (N_2199,N_1258,N_1954);
nand U2200 (N_2200,N_1779,N_1905);
or U2201 (N_2201,N_1881,N_1549);
nand U2202 (N_2202,N_1227,N_1275);
nand U2203 (N_2203,N_1405,N_1305);
nand U2204 (N_2204,N_1945,N_1322);
or U2205 (N_2205,N_1359,N_1046);
nand U2206 (N_2206,N_1368,N_1374);
or U2207 (N_2207,N_1529,N_1657);
nand U2208 (N_2208,N_1897,N_1654);
or U2209 (N_2209,N_1946,N_1720);
and U2210 (N_2210,N_1087,N_1267);
nor U2211 (N_2211,N_1231,N_1792);
or U2212 (N_2212,N_1390,N_1959);
and U2213 (N_2213,N_1034,N_1311);
nand U2214 (N_2214,N_1794,N_1325);
or U2215 (N_2215,N_1724,N_1161);
nand U2216 (N_2216,N_1803,N_1887);
or U2217 (N_2217,N_1314,N_1287);
nor U2218 (N_2218,N_1002,N_1821);
or U2219 (N_2219,N_1673,N_1682);
nand U2220 (N_2220,N_1915,N_1777);
nand U2221 (N_2221,N_1577,N_1734);
nor U2222 (N_2222,N_1603,N_1225);
nand U2223 (N_2223,N_1843,N_1215);
nand U2224 (N_2224,N_1360,N_1437);
or U2225 (N_2225,N_1647,N_1300);
nor U2226 (N_2226,N_1179,N_1107);
and U2227 (N_2227,N_1078,N_1702);
and U2228 (N_2228,N_1943,N_1163);
nor U2229 (N_2229,N_1153,N_1539);
nor U2230 (N_2230,N_1990,N_1271);
nand U2231 (N_2231,N_1538,N_1141);
or U2232 (N_2232,N_1421,N_1578);
nand U2233 (N_2233,N_1929,N_1456);
or U2234 (N_2234,N_1207,N_1385);
and U2235 (N_2235,N_1812,N_1964);
nand U2236 (N_2236,N_1484,N_1205);
and U2237 (N_2237,N_1350,N_1151);
or U2238 (N_2238,N_1389,N_1799);
or U2239 (N_2239,N_1617,N_1967);
and U2240 (N_2240,N_1100,N_1127);
nor U2241 (N_2241,N_1847,N_1801);
and U2242 (N_2242,N_1642,N_1741);
nor U2243 (N_2243,N_1171,N_1955);
nor U2244 (N_2244,N_1041,N_1254);
xnor U2245 (N_2245,N_1663,N_1376);
nor U2246 (N_2246,N_1725,N_1713);
and U2247 (N_2247,N_1722,N_1966);
or U2248 (N_2248,N_1265,N_1700);
or U2249 (N_2249,N_1488,N_1263);
or U2250 (N_2250,N_1485,N_1626);
and U2251 (N_2251,N_1011,N_1534);
and U2252 (N_2252,N_1589,N_1771);
and U2253 (N_2253,N_1381,N_1156);
and U2254 (N_2254,N_1970,N_1144);
nand U2255 (N_2255,N_1693,N_1172);
and U2256 (N_2256,N_1032,N_1721);
nand U2257 (N_2257,N_1531,N_1840);
nand U2258 (N_2258,N_1160,N_1018);
nand U2259 (N_2259,N_1772,N_1169);
nor U2260 (N_2260,N_1509,N_1343);
nor U2261 (N_2261,N_1507,N_1422);
or U2262 (N_2262,N_1892,N_1826);
nor U2263 (N_2263,N_1524,N_1543);
nor U2264 (N_2264,N_1944,N_1756);
and U2265 (N_2265,N_1201,N_1450);
and U2266 (N_2266,N_1923,N_1778);
or U2267 (N_2267,N_1382,N_1894);
and U2268 (N_2268,N_1653,N_1804);
nand U2269 (N_2269,N_1732,N_1035);
and U2270 (N_2270,N_1902,N_1952);
nor U2271 (N_2271,N_1012,N_1138);
nand U2272 (N_2272,N_1723,N_1030);
nand U2273 (N_2273,N_1701,N_1423);
nor U2274 (N_2274,N_1927,N_1447);
or U2275 (N_2275,N_1040,N_1685);
or U2276 (N_2276,N_1098,N_1214);
or U2277 (N_2277,N_1689,N_1845);
and U2278 (N_2278,N_1162,N_1555);
and U2279 (N_2279,N_1979,N_1584);
or U2280 (N_2280,N_1869,N_1296);
nand U2281 (N_2281,N_1601,N_1186);
nand U2282 (N_2282,N_1009,N_1412);
and U2283 (N_2283,N_1688,N_1375);
nor U2284 (N_2284,N_1045,N_1914);
nand U2285 (N_2285,N_1888,N_1659);
nor U2286 (N_2286,N_1669,N_1680);
or U2287 (N_2287,N_1341,N_1838);
and U2288 (N_2288,N_1760,N_1824);
xnor U2289 (N_2289,N_1833,N_1828);
or U2290 (N_2290,N_1031,N_1913);
nor U2291 (N_2291,N_1851,N_1364);
and U2292 (N_2292,N_1282,N_1429);
nand U2293 (N_2293,N_1315,N_1369);
nor U2294 (N_2294,N_1909,N_1514);
or U2295 (N_2295,N_1089,N_1561);
nand U2296 (N_2296,N_1746,N_1865);
nor U2297 (N_2297,N_1399,N_1292);
nand U2298 (N_2298,N_1683,N_1769);
nor U2299 (N_2299,N_1233,N_1250);
nor U2300 (N_2300,N_1468,N_1789);
nand U2301 (N_2301,N_1337,N_1924);
nand U2302 (N_2302,N_1269,N_1950);
xnor U2303 (N_2303,N_1863,N_1490);
and U2304 (N_2304,N_1330,N_1545);
or U2305 (N_2305,N_1586,N_1195);
nand U2306 (N_2306,N_1920,N_1731);
and U2307 (N_2307,N_1244,N_1922);
nor U2308 (N_2308,N_1615,N_1535);
or U2309 (N_2309,N_1434,N_1353);
nor U2310 (N_2310,N_1358,N_1323);
and U2311 (N_2311,N_1540,N_1666);
nor U2312 (N_2312,N_1896,N_1097);
nor U2313 (N_2313,N_1174,N_1068);
or U2314 (N_2314,N_1420,N_1791);
and U2315 (N_2315,N_1248,N_1066);
nand U2316 (N_2316,N_1585,N_1198);
nor U2317 (N_2317,N_1036,N_1120);
nand U2318 (N_2318,N_1607,N_1730);
or U2319 (N_2319,N_1139,N_1819);
nand U2320 (N_2320,N_1858,N_1798);
nor U2321 (N_2321,N_1115,N_1864);
and U2322 (N_2322,N_1925,N_1569);
nor U2323 (N_2323,N_1916,N_1299);
nand U2324 (N_2324,N_1039,N_1261);
or U2325 (N_2325,N_1676,N_1557);
nor U2326 (N_2326,N_1255,N_1432);
nand U2327 (N_2327,N_1229,N_1338);
nand U2328 (N_2328,N_1889,N_1753);
or U2329 (N_2329,N_1427,N_1655);
nand U2330 (N_2330,N_1007,N_1074);
nand U2331 (N_2331,N_1912,N_1934);
or U2332 (N_2332,N_1494,N_1101);
nand U2333 (N_2333,N_1416,N_1204);
or U2334 (N_2334,N_1775,N_1740);
or U2335 (N_2335,N_1339,N_1627);
and U2336 (N_2336,N_1043,N_1417);
and U2337 (N_2337,N_1681,N_1528);
nor U2338 (N_2338,N_1823,N_1483);
and U2339 (N_2339,N_1152,N_1709);
or U2340 (N_2340,N_1773,N_1383);
and U2341 (N_2341,N_1984,N_1223);
and U2342 (N_2342,N_1266,N_1570);
or U2343 (N_2343,N_1783,N_1413);
or U2344 (N_2344,N_1690,N_1398);
nor U2345 (N_2345,N_1291,N_1452);
or U2346 (N_2346,N_1363,N_1882);
nor U2347 (N_2347,N_1558,N_1989);
nor U2348 (N_2348,N_1795,N_1426);
and U2349 (N_2349,N_1822,N_1264);
or U2350 (N_2350,N_1511,N_1280);
or U2351 (N_2351,N_1747,N_1907);
or U2352 (N_2352,N_1620,N_1308);
and U2353 (N_2353,N_1932,N_1767);
or U2354 (N_2354,N_1868,N_1854);
nor U2355 (N_2355,N_1602,N_1246);
and U2356 (N_2356,N_1692,N_1855);
and U2357 (N_2357,N_1202,N_1178);
and U2358 (N_2358,N_1076,N_1058);
and U2359 (N_2359,N_1003,N_1764);
nand U2360 (N_2360,N_1571,N_1910);
or U2361 (N_2361,N_1226,N_1606);
or U2362 (N_2362,N_1155,N_1410);
or U2363 (N_2363,N_1904,N_1142);
or U2364 (N_2364,N_1272,N_1991);
nand U2365 (N_2365,N_1026,N_1016);
nand U2366 (N_2366,N_1883,N_1813);
or U2367 (N_2367,N_1388,N_1048);
and U2368 (N_2368,N_1307,N_1073);
or U2369 (N_2369,N_1023,N_1199);
nand U2370 (N_2370,N_1595,N_1593);
nand U2371 (N_2371,N_1372,N_1951);
or U2372 (N_2372,N_1431,N_1830);
or U2373 (N_2373,N_1402,N_1498);
nor U2374 (N_2374,N_1928,N_1599);
nand U2375 (N_2375,N_1958,N_1661);
and U2376 (N_2376,N_1212,N_1703);
and U2377 (N_2377,N_1118,N_1222);
or U2378 (N_2378,N_1176,N_1210);
or U2379 (N_2379,N_1829,N_1985);
or U2380 (N_2380,N_1503,N_1459);
nand U2381 (N_2381,N_1328,N_1481);
or U2382 (N_2382,N_1612,N_1096);
and U2383 (N_2383,N_1240,N_1334);
nand U2384 (N_2384,N_1611,N_1980);
nand U2385 (N_2385,N_1800,N_1070);
and U2386 (N_2386,N_1218,N_1029);
or U2387 (N_2387,N_1200,N_1211);
nor U2388 (N_2388,N_1987,N_1699);
nand U2389 (N_2389,N_1117,N_1079);
or U2390 (N_2390,N_1182,N_1033);
nor U2391 (N_2391,N_1464,N_1900);
or U2392 (N_2392,N_1765,N_1658);
nand U2393 (N_2393,N_1839,N_1786);
nor U2394 (N_2394,N_1960,N_1213);
or U2395 (N_2395,N_1466,N_1761);
nor U2396 (N_2396,N_1154,N_1166);
and U2397 (N_2397,N_1542,N_1493);
nand U2398 (N_2398,N_1745,N_1818);
nor U2399 (N_2399,N_1708,N_1936);
nand U2400 (N_2400,N_1971,N_1188);
or U2401 (N_2401,N_1252,N_1969);
nor U2402 (N_2402,N_1480,N_1797);
nand U2403 (N_2403,N_1268,N_1164);
nand U2404 (N_2404,N_1396,N_1533);
nor U2405 (N_2405,N_1748,N_1580);
or U2406 (N_2406,N_1491,N_1998);
and U2407 (N_2407,N_1596,N_1505);
and U2408 (N_2408,N_1633,N_1582);
nor U2409 (N_2409,N_1216,N_1664);
or U2410 (N_2410,N_1527,N_1407);
nor U2411 (N_2411,N_1972,N_1404);
nor U2412 (N_2412,N_1137,N_1183);
or U2413 (N_2413,N_1784,N_1114);
nor U2414 (N_2414,N_1049,N_1309);
or U2415 (N_2415,N_1776,N_1067);
nor U2416 (N_2416,N_1397,N_1387);
nor U2417 (N_2417,N_1108,N_1793);
nand U2418 (N_2418,N_1247,N_1392);
xnor U2419 (N_2419,N_1796,N_1104);
and U2420 (N_2420,N_1742,N_1842);
and U2421 (N_2421,N_1641,N_1895);
nor U2422 (N_2422,N_1028,N_1921);
and U2423 (N_2423,N_1080,N_1495);
nand U2424 (N_2424,N_1719,N_1684);
and U2425 (N_2425,N_1717,N_1196);
or U2426 (N_2426,N_1551,N_1541);
and U2427 (N_2427,N_1332,N_1022);
or U2428 (N_2428,N_1992,N_1500);
and U2429 (N_2429,N_1517,N_1159);
nand U2430 (N_2430,N_1095,N_1351);
nor U2431 (N_2431,N_1403,N_1848);
and U2432 (N_2432,N_1257,N_1081);
nor U2433 (N_2433,N_1109,N_1132);
nand U2434 (N_2434,N_1377,N_1345);
or U2435 (N_2435,N_1636,N_1038);
and U2436 (N_2436,N_1455,N_1573);
nand U2437 (N_2437,N_1295,N_1788);
nand U2438 (N_2438,N_1553,N_1497);
nand U2439 (N_2439,N_1544,N_1994);
or U2440 (N_2440,N_1630,N_1597);
nand U2441 (N_2441,N_1867,N_1879);
and U2442 (N_2442,N_1367,N_1105);
and U2443 (N_2443,N_1084,N_1832);
and U2444 (N_2444,N_1901,N_1072);
nor U2445 (N_2445,N_1716,N_1512);
nor U2446 (N_2446,N_1744,N_1706);
nand U2447 (N_2447,N_1460,N_1436);
or U2448 (N_2448,N_1184,N_1841);
or U2449 (N_2449,N_1825,N_1727);
nand U2450 (N_2450,N_1430,N_1005);
nor U2451 (N_2451,N_1333,N_1177);
and U2452 (N_2452,N_1454,N_1192);
nand U2453 (N_2453,N_1768,N_1479);
or U2454 (N_2454,N_1119,N_1013);
or U2455 (N_2455,N_1621,N_1221);
or U2456 (N_2456,N_1203,N_1283);
or U2457 (N_2457,N_1463,N_1469);
or U2458 (N_2458,N_1303,N_1477);
or U2459 (N_2459,N_1890,N_1425);
xor U2460 (N_2460,N_1090,N_1933);
nor U2461 (N_2461,N_1165,N_1441);
or U2462 (N_2462,N_1576,N_1134);
or U2463 (N_2463,N_1572,N_1757);
nand U2464 (N_2464,N_1579,N_1605);
xor U2465 (N_2465,N_1941,N_1835);
nor U2466 (N_2466,N_1239,N_1489);
and U2467 (N_2467,N_1052,N_1686);
nor U2468 (N_2468,N_1537,N_1017);
nor U2469 (N_2469,N_1604,N_1691);
nor U2470 (N_2470,N_1939,N_1461);
nor U2471 (N_2471,N_1947,N_1110);
and U2472 (N_2472,N_1759,N_1094);
or U2473 (N_2473,N_1616,N_1391);
or U2474 (N_2474,N_1856,N_1148);
and U2475 (N_2475,N_1634,N_1976);
or U2476 (N_2476,N_1536,N_1968);
and U2477 (N_2477,N_1808,N_1249);
and U2478 (N_2478,N_1181,N_1817);
nand U2479 (N_2479,N_1378,N_1762);
or U2480 (N_2480,N_1279,N_1644);
nand U2481 (N_2481,N_1276,N_1243);
and U2482 (N_2482,N_1286,N_1917);
nand U2483 (N_2483,N_1451,N_1880);
and U2484 (N_2484,N_1224,N_1077);
nor U2485 (N_2485,N_1938,N_1501);
or U2486 (N_2486,N_1125,N_1637);
nand U2487 (N_2487,N_1737,N_1728);
and U2488 (N_2488,N_1475,N_1885);
and U2489 (N_2489,N_1629,N_1047);
nand U2490 (N_2490,N_1302,N_1962);
and U2491 (N_2491,N_1610,N_1406);
or U2492 (N_2492,N_1608,N_1288);
and U2493 (N_2493,N_1476,N_1465);
or U2494 (N_2494,N_1956,N_1319);
or U2495 (N_2495,N_1349,N_1619);
nand U2496 (N_2496,N_1981,N_1852);
and U2497 (N_2497,N_1526,N_1592);
xor U2498 (N_2498,N_1342,N_1591);
and U2499 (N_2499,N_1893,N_1649);
nor U2500 (N_2500,N_1400,N_1818);
nand U2501 (N_2501,N_1489,N_1378);
or U2502 (N_2502,N_1121,N_1436);
xor U2503 (N_2503,N_1258,N_1643);
nor U2504 (N_2504,N_1272,N_1399);
or U2505 (N_2505,N_1080,N_1070);
or U2506 (N_2506,N_1984,N_1999);
or U2507 (N_2507,N_1356,N_1143);
and U2508 (N_2508,N_1557,N_1578);
nor U2509 (N_2509,N_1632,N_1400);
nor U2510 (N_2510,N_1774,N_1345);
or U2511 (N_2511,N_1112,N_1372);
nor U2512 (N_2512,N_1075,N_1907);
and U2513 (N_2513,N_1575,N_1632);
and U2514 (N_2514,N_1534,N_1874);
or U2515 (N_2515,N_1814,N_1305);
or U2516 (N_2516,N_1878,N_1560);
or U2517 (N_2517,N_1950,N_1466);
and U2518 (N_2518,N_1198,N_1946);
and U2519 (N_2519,N_1002,N_1661);
or U2520 (N_2520,N_1404,N_1993);
and U2521 (N_2521,N_1256,N_1899);
or U2522 (N_2522,N_1867,N_1458);
nand U2523 (N_2523,N_1499,N_1784);
or U2524 (N_2524,N_1803,N_1247);
nor U2525 (N_2525,N_1489,N_1510);
nor U2526 (N_2526,N_1209,N_1024);
nor U2527 (N_2527,N_1106,N_1462);
nor U2528 (N_2528,N_1038,N_1627);
nor U2529 (N_2529,N_1500,N_1580);
nand U2530 (N_2530,N_1781,N_1375);
or U2531 (N_2531,N_1765,N_1776);
or U2532 (N_2532,N_1727,N_1433);
and U2533 (N_2533,N_1253,N_1489);
nand U2534 (N_2534,N_1131,N_1856);
or U2535 (N_2535,N_1913,N_1277);
or U2536 (N_2536,N_1622,N_1186);
nor U2537 (N_2537,N_1170,N_1423);
or U2538 (N_2538,N_1547,N_1580);
or U2539 (N_2539,N_1865,N_1818);
or U2540 (N_2540,N_1381,N_1700);
nor U2541 (N_2541,N_1297,N_1339);
and U2542 (N_2542,N_1861,N_1157);
nand U2543 (N_2543,N_1486,N_1474);
nand U2544 (N_2544,N_1646,N_1763);
nor U2545 (N_2545,N_1162,N_1237);
or U2546 (N_2546,N_1689,N_1009);
nand U2547 (N_2547,N_1646,N_1123);
or U2548 (N_2548,N_1072,N_1306);
nand U2549 (N_2549,N_1686,N_1139);
nand U2550 (N_2550,N_1929,N_1527);
or U2551 (N_2551,N_1710,N_1897);
nand U2552 (N_2552,N_1457,N_1071);
or U2553 (N_2553,N_1337,N_1057);
and U2554 (N_2554,N_1961,N_1493);
or U2555 (N_2555,N_1974,N_1752);
and U2556 (N_2556,N_1901,N_1058);
or U2557 (N_2557,N_1092,N_1898);
nand U2558 (N_2558,N_1060,N_1965);
or U2559 (N_2559,N_1320,N_1715);
nor U2560 (N_2560,N_1031,N_1499);
nand U2561 (N_2561,N_1512,N_1923);
and U2562 (N_2562,N_1804,N_1932);
and U2563 (N_2563,N_1815,N_1221);
and U2564 (N_2564,N_1596,N_1614);
and U2565 (N_2565,N_1811,N_1945);
or U2566 (N_2566,N_1864,N_1867);
nand U2567 (N_2567,N_1894,N_1343);
and U2568 (N_2568,N_1374,N_1643);
or U2569 (N_2569,N_1081,N_1876);
and U2570 (N_2570,N_1988,N_1582);
nand U2571 (N_2571,N_1328,N_1870);
or U2572 (N_2572,N_1596,N_1996);
or U2573 (N_2573,N_1178,N_1088);
or U2574 (N_2574,N_1034,N_1915);
nor U2575 (N_2575,N_1494,N_1056);
nor U2576 (N_2576,N_1430,N_1832);
or U2577 (N_2577,N_1482,N_1122);
or U2578 (N_2578,N_1197,N_1976);
nor U2579 (N_2579,N_1468,N_1505);
and U2580 (N_2580,N_1861,N_1962);
nor U2581 (N_2581,N_1091,N_1008);
nand U2582 (N_2582,N_1527,N_1836);
nand U2583 (N_2583,N_1288,N_1390);
and U2584 (N_2584,N_1241,N_1948);
or U2585 (N_2585,N_1852,N_1058);
nor U2586 (N_2586,N_1873,N_1187);
or U2587 (N_2587,N_1647,N_1028);
nand U2588 (N_2588,N_1970,N_1700);
or U2589 (N_2589,N_1924,N_1173);
or U2590 (N_2590,N_1863,N_1528);
nor U2591 (N_2591,N_1073,N_1649);
nand U2592 (N_2592,N_1325,N_1404);
and U2593 (N_2593,N_1044,N_1901);
nor U2594 (N_2594,N_1039,N_1071);
or U2595 (N_2595,N_1573,N_1805);
and U2596 (N_2596,N_1278,N_1858);
and U2597 (N_2597,N_1989,N_1263);
nor U2598 (N_2598,N_1739,N_1366);
or U2599 (N_2599,N_1292,N_1030);
or U2600 (N_2600,N_1586,N_1855);
and U2601 (N_2601,N_1039,N_1537);
and U2602 (N_2602,N_1979,N_1479);
nand U2603 (N_2603,N_1634,N_1591);
nor U2604 (N_2604,N_1685,N_1122);
nor U2605 (N_2605,N_1281,N_1390);
nor U2606 (N_2606,N_1477,N_1849);
nor U2607 (N_2607,N_1252,N_1614);
nand U2608 (N_2608,N_1676,N_1923);
or U2609 (N_2609,N_1114,N_1584);
or U2610 (N_2610,N_1019,N_1780);
nand U2611 (N_2611,N_1347,N_1360);
nor U2612 (N_2612,N_1717,N_1983);
nand U2613 (N_2613,N_1352,N_1758);
or U2614 (N_2614,N_1390,N_1835);
and U2615 (N_2615,N_1351,N_1091);
nand U2616 (N_2616,N_1588,N_1438);
or U2617 (N_2617,N_1974,N_1869);
or U2618 (N_2618,N_1935,N_1006);
or U2619 (N_2619,N_1214,N_1945);
nand U2620 (N_2620,N_1690,N_1145);
nor U2621 (N_2621,N_1806,N_1252);
and U2622 (N_2622,N_1847,N_1085);
nand U2623 (N_2623,N_1862,N_1131);
or U2624 (N_2624,N_1817,N_1869);
nand U2625 (N_2625,N_1056,N_1511);
and U2626 (N_2626,N_1460,N_1959);
nand U2627 (N_2627,N_1695,N_1964);
and U2628 (N_2628,N_1037,N_1162);
nand U2629 (N_2629,N_1835,N_1664);
and U2630 (N_2630,N_1103,N_1131);
or U2631 (N_2631,N_1487,N_1379);
nor U2632 (N_2632,N_1111,N_1803);
nand U2633 (N_2633,N_1636,N_1676);
or U2634 (N_2634,N_1690,N_1860);
and U2635 (N_2635,N_1264,N_1515);
or U2636 (N_2636,N_1601,N_1977);
nand U2637 (N_2637,N_1124,N_1022);
nor U2638 (N_2638,N_1831,N_1721);
nor U2639 (N_2639,N_1069,N_1903);
nand U2640 (N_2640,N_1037,N_1514);
or U2641 (N_2641,N_1078,N_1500);
nand U2642 (N_2642,N_1260,N_1584);
nand U2643 (N_2643,N_1056,N_1766);
or U2644 (N_2644,N_1212,N_1612);
nand U2645 (N_2645,N_1652,N_1136);
or U2646 (N_2646,N_1728,N_1133);
nand U2647 (N_2647,N_1953,N_1981);
nand U2648 (N_2648,N_1380,N_1634);
and U2649 (N_2649,N_1612,N_1762);
nand U2650 (N_2650,N_1753,N_1818);
nand U2651 (N_2651,N_1828,N_1185);
or U2652 (N_2652,N_1233,N_1983);
and U2653 (N_2653,N_1235,N_1976);
nand U2654 (N_2654,N_1026,N_1765);
nand U2655 (N_2655,N_1206,N_1090);
or U2656 (N_2656,N_1786,N_1508);
and U2657 (N_2657,N_1304,N_1136);
nand U2658 (N_2658,N_1929,N_1010);
or U2659 (N_2659,N_1248,N_1445);
nor U2660 (N_2660,N_1427,N_1080);
or U2661 (N_2661,N_1976,N_1236);
nand U2662 (N_2662,N_1620,N_1528);
or U2663 (N_2663,N_1808,N_1374);
and U2664 (N_2664,N_1308,N_1542);
or U2665 (N_2665,N_1730,N_1235);
or U2666 (N_2666,N_1889,N_1555);
and U2667 (N_2667,N_1496,N_1839);
or U2668 (N_2668,N_1852,N_1874);
nor U2669 (N_2669,N_1025,N_1357);
and U2670 (N_2670,N_1888,N_1942);
nand U2671 (N_2671,N_1369,N_1879);
and U2672 (N_2672,N_1819,N_1822);
nand U2673 (N_2673,N_1703,N_1770);
or U2674 (N_2674,N_1030,N_1686);
or U2675 (N_2675,N_1664,N_1922);
or U2676 (N_2676,N_1760,N_1853);
or U2677 (N_2677,N_1988,N_1698);
nand U2678 (N_2678,N_1190,N_1332);
nand U2679 (N_2679,N_1489,N_1919);
nor U2680 (N_2680,N_1836,N_1764);
nor U2681 (N_2681,N_1359,N_1603);
nand U2682 (N_2682,N_1305,N_1050);
nor U2683 (N_2683,N_1682,N_1902);
nor U2684 (N_2684,N_1406,N_1697);
and U2685 (N_2685,N_1010,N_1540);
nand U2686 (N_2686,N_1434,N_1319);
or U2687 (N_2687,N_1243,N_1217);
and U2688 (N_2688,N_1849,N_1806);
and U2689 (N_2689,N_1771,N_1920);
or U2690 (N_2690,N_1202,N_1915);
nand U2691 (N_2691,N_1612,N_1533);
nor U2692 (N_2692,N_1654,N_1587);
xor U2693 (N_2693,N_1256,N_1896);
nand U2694 (N_2694,N_1936,N_1697);
or U2695 (N_2695,N_1204,N_1344);
xor U2696 (N_2696,N_1999,N_1742);
and U2697 (N_2697,N_1535,N_1015);
nor U2698 (N_2698,N_1391,N_1910);
nor U2699 (N_2699,N_1126,N_1654);
nor U2700 (N_2700,N_1649,N_1045);
or U2701 (N_2701,N_1765,N_1032);
nor U2702 (N_2702,N_1398,N_1624);
or U2703 (N_2703,N_1649,N_1837);
nand U2704 (N_2704,N_1896,N_1889);
and U2705 (N_2705,N_1437,N_1204);
nor U2706 (N_2706,N_1988,N_1061);
and U2707 (N_2707,N_1783,N_1139);
nor U2708 (N_2708,N_1950,N_1019);
nor U2709 (N_2709,N_1600,N_1966);
or U2710 (N_2710,N_1825,N_1410);
nor U2711 (N_2711,N_1432,N_1423);
and U2712 (N_2712,N_1021,N_1444);
or U2713 (N_2713,N_1505,N_1680);
or U2714 (N_2714,N_1093,N_1414);
nand U2715 (N_2715,N_1597,N_1785);
nand U2716 (N_2716,N_1055,N_1317);
xnor U2717 (N_2717,N_1551,N_1908);
nor U2718 (N_2718,N_1756,N_1028);
and U2719 (N_2719,N_1150,N_1697);
nor U2720 (N_2720,N_1226,N_1034);
and U2721 (N_2721,N_1176,N_1977);
nor U2722 (N_2722,N_1048,N_1306);
or U2723 (N_2723,N_1868,N_1981);
or U2724 (N_2724,N_1637,N_1240);
nand U2725 (N_2725,N_1311,N_1378);
nand U2726 (N_2726,N_1812,N_1493);
and U2727 (N_2727,N_1900,N_1372);
and U2728 (N_2728,N_1171,N_1172);
or U2729 (N_2729,N_1487,N_1650);
nand U2730 (N_2730,N_1127,N_1673);
nor U2731 (N_2731,N_1411,N_1167);
or U2732 (N_2732,N_1666,N_1773);
xnor U2733 (N_2733,N_1270,N_1133);
and U2734 (N_2734,N_1070,N_1495);
nor U2735 (N_2735,N_1046,N_1833);
and U2736 (N_2736,N_1003,N_1445);
nor U2737 (N_2737,N_1439,N_1404);
or U2738 (N_2738,N_1132,N_1566);
nand U2739 (N_2739,N_1962,N_1053);
nand U2740 (N_2740,N_1686,N_1391);
and U2741 (N_2741,N_1973,N_1101);
nand U2742 (N_2742,N_1528,N_1371);
and U2743 (N_2743,N_1708,N_1371);
nor U2744 (N_2744,N_1777,N_1098);
or U2745 (N_2745,N_1038,N_1653);
and U2746 (N_2746,N_1795,N_1340);
and U2747 (N_2747,N_1354,N_1328);
nor U2748 (N_2748,N_1517,N_1809);
and U2749 (N_2749,N_1990,N_1349);
or U2750 (N_2750,N_1934,N_1259);
or U2751 (N_2751,N_1180,N_1852);
and U2752 (N_2752,N_1110,N_1389);
nor U2753 (N_2753,N_1714,N_1880);
nor U2754 (N_2754,N_1919,N_1729);
and U2755 (N_2755,N_1716,N_1730);
and U2756 (N_2756,N_1268,N_1450);
and U2757 (N_2757,N_1206,N_1331);
or U2758 (N_2758,N_1590,N_1119);
and U2759 (N_2759,N_1659,N_1857);
nor U2760 (N_2760,N_1589,N_1475);
nor U2761 (N_2761,N_1524,N_1504);
nor U2762 (N_2762,N_1891,N_1275);
and U2763 (N_2763,N_1973,N_1501);
xnor U2764 (N_2764,N_1468,N_1415);
nand U2765 (N_2765,N_1697,N_1462);
or U2766 (N_2766,N_1090,N_1866);
nand U2767 (N_2767,N_1885,N_1271);
and U2768 (N_2768,N_1562,N_1278);
and U2769 (N_2769,N_1702,N_1669);
nand U2770 (N_2770,N_1921,N_1699);
or U2771 (N_2771,N_1646,N_1555);
nand U2772 (N_2772,N_1628,N_1583);
or U2773 (N_2773,N_1634,N_1073);
or U2774 (N_2774,N_1169,N_1275);
or U2775 (N_2775,N_1966,N_1347);
nor U2776 (N_2776,N_1356,N_1895);
nor U2777 (N_2777,N_1566,N_1954);
nand U2778 (N_2778,N_1013,N_1163);
nor U2779 (N_2779,N_1091,N_1612);
nand U2780 (N_2780,N_1294,N_1123);
nand U2781 (N_2781,N_1774,N_1979);
nand U2782 (N_2782,N_1805,N_1644);
nand U2783 (N_2783,N_1340,N_1784);
or U2784 (N_2784,N_1479,N_1729);
and U2785 (N_2785,N_1027,N_1670);
or U2786 (N_2786,N_1439,N_1136);
nand U2787 (N_2787,N_1725,N_1078);
nor U2788 (N_2788,N_1901,N_1650);
nand U2789 (N_2789,N_1314,N_1408);
and U2790 (N_2790,N_1652,N_1508);
and U2791 (N_2791,N_1719,N_1212);
and U2792 (N_2792,N_1670,N_1153);
nor U2793 (N_2793,N_1938,N_1482);
and U2794 (N_2794,N_1770,N_1782);
nor U2795 (N_2795,N_1600,N_1630);
or U2796 (N_2796,N_1331,N_1726);
nor U2797 (N_2797,N_1929,N_1758);
or U2798 (N_2798,N_1184,N_1362);
nand U2799 (N_2799,N_1137,N_1489);
nor U2800 (N_2800,N_1647,N_1566);
nand U2801 (N_2801,N_1181,N_1520);
nand U2802 (N_2802,N_1555,N_1254);
nor U2803 (N_2803,N_1126,N_1566);
nand U2804 (N_2804,N_1460,N_1973);
nand U2805 (N_2805,N_1524,N_1280);
or U2806 (N_2806,N_1495,N_1149);
and U2807 (N_2807,N_1496,N_1622);
or U2808 (N_2808,N_1081,N_1487);
nor U2809 (N_2809,N_1653,N_1163);
nand U2810 (N_2810,N_1560,N_1992);
nand U2811 (N_2811,N_1142,N_1778);
nand U2812 (N_2812,N_1671,N_1489);
or U2813 (N_2813,N_1182,N_1004);
nand U2814 (N_2814,N_1466,N_1255);
nor U2815 (N_2815,N_1439,N_1152);
and U2816 (N_2816,N_1994,N_1128);
or U2817 (N_2817,N_1053,N_1205);
nor U2818 (N_2818,N_1684,N_1190);
or U2819 (N_2819,N_1361,N_1532);
and U2820 (N_2820,N_1290,N_1841);
or U2821 (N_2821,N_1515,N_1972);
or U2822 (N_2822,N_1718,N_1015);
nor U2823 (N_2823,N_1951,N_1546);
or U2824 (N_2824,N_1839,N_1170);
nand U2825 (N_2825,N_1157,N_1510);
and U2826 (N_2826,N_1138,N_1777);
or U2827 (N_2827,N_1012,N_1238);
nand U2828 (N_2828,N_1130,N_1780);
or U2829 (N_2829,N_1177,N_1427);
nand U2830 (N_2830,N_1007,N_1172);
and U2831 (N_2831,N_1551,N_1685);
or U2832 (N_2832,N_1676,N_1453);
or U2833 (N_2833,N_1498,N_1652);
or U2834 (N_2834,N_1584,N_1699);
or U2835 (N_2835,N_1478,N_1414);
or U2836 (N_2836,N_1555,N_1777);
or U2837 (N_2837,N_1651,N_1381);
nor U2838 (N_2838,N_1070,N_1551);
nor U2839 (N_2839,N_1832,N_1867);
and U2840 (N_2840,N_1227,N_1855);
nand U2841 (N_2841,N_1504,N_1507);
nand U2842 (N_2842,N_1892,N_1415);
or U2843 (N_2843,N_1537,N_1805);
or U2844 (N_2844,N_1398,N_1332);
and U2845 (N_2845,N_1131,N_1820);
or U2846 (N_2846,N_1493,N_1631);
nand U2847 (N_2847,N_1560,N_1092);
nor U2848 (N_2848,N_1896,N_1682);
nand U2849 (N_2849,N_1505,N_1404);
nand U2850 (N_2850,N_1058,N_1445);
nand U2851 (N_2851,N_1086,N_1286);
xnor U2852 (N_2852,N_1592,N_1582);
and U2853 (N_2853,N_1433,N_1112);
and U2854 (N_2854,N_1554,N_1095);
and U2855 (N_2855,N_1202,N_1795);
and U2856 (N_2856,N_1429,N_1827);
nand U2857 (N_2857,N_1409,N_1065);
and U2858 (N_2858,N_1451,N_1784);
and U2859 (N_2859,N_1503,N_1413);
nand U2860 (N_2860,N_1650,N_1450);
nand U2861 (N_2861,N_1765,N_1197);
and U2862 (N_2862,N_1825,N_1892);
or U2863 (N_2863,N_1217,N_1180);
nand U2864 (N_2864,N_1532,N_1011);
nor U2865 (N_2865,N_1517,N_1769);
or U2866 (N_2866,N_1155,N_1209);
and U2867 (N_2867,N_1788,N_1984);
or U2868 (N_2868,N_1620,N_1432);
nor U2869 (N_2869,N_1717,N_1123);
nand U2870 (N_2870,N_1284,N_1278);
nor U2871 (N_2871,N_1535,N_1512);
nor U2872 (N_2872,N_1233,N_1692);
or U2873 (N_2873,N_1500,N_1791);
nand U2874 (N_2874,N_1578,N_1371);
nand U2875 (N_2875,N_1117,N_1191);
or U2876 (N_2876,N_1038,N_1643);
and U2877 (N_2877,N_1046,N_1158);
and U2878 (N_2878,N_1797,N_1757);
or U2879 (N_2879,N_1602,N_1505);
and U2880 (N_2880,N_1286,N_1609);
nor U2881 (N_2881,N_1486,N_1693);
nand U2882 (N_2882,N_1518,N_1154);
nor U2883 (N_2883,N_1693,N_1615);
nand U2884 (N_2884,N_1543,N_1414);
or U2885 (N_2885,N_1908,N_1666);
nor U2886 (N_2886,N_1907,N_1885);
nor U2887 (N_2887,N_1660,N_1104);
nand U2888 (N_2888,N_1676,N_1926);
nand U2889 (N_2889,N_1053,N_1960);
and U2890 (N_2890,N_1650,N_1267);
and U2891 (N_2891,N_1030,N_1572);
nor U2892 (N_2892,N_1053,N_1945);
or U2893 (N_2893,N_1912,N_1758);
nand U2894 (N_2894,N_1251,N_1289);
and U2895 (N_2895,N_1746,N_1353);
or U2896 (N_2896,N_1438,N_1596);
nor U2897 (N_2897,N_1753,N_1319);
nor U2898 (N_2898,N_1406,N_1189);
nor U2899 (N_2899,N_1023,N_1830);
or U2900 (N_2900,N_1389,N_1858);
nor U2901 (N_2901,N_1585,N_1117);
or U2902 (N_2902,N_1778,N_1019);
nor U2903 (N_2903,N_1771,N_1671);
or U2904 (N_2904,N_1287,N_1384);
nand U2905 (N_2905,N_1042,N_1029);
nand U2906 (N_2906,N_1275,N_1840);
nor U2907 (N_2907,N_1268,N_1558);
nor U2908 (N_2908,N_1432,N_1110);
and U2909 (N_2909,N_1771,N_1930);
nor U2910 (N_2910,N_1863,N_1649);
nor U2911 (N_2911,N_1073,N_1810);
nand U2912 (N_2912,N_1316,N_1711);
nand U2913 (N_2913,N_1598,N_1079);
nand U2914 (N_2914,N_1481,N_1299);
nor U2915 (N_2915,N_1590,N_1627);
and U2916 (N_2916,N_1515,N_1496);
and U2917 (N_2917,N_1578,N_1469);
nand U2918 (N_2918,N_1608,N_1791);
and U2919 (N_2919,N_1423,N_1481);
nand U2920 (N_2920,N_1040,N_1094);
and U2921 (N_2921,N_1363,N_1070);
or U2922 (N_2922,N_1616,N_1022);
nand U2923 (N_2923,N_1803,N_1285);
nor U2924 (N_2924,N_1891,N_1088);
nor U2925 (N_2925,N_1195,N_1464);
and U2926 (N_2926,N_1853,N_1886);
or U2927 (N_2927,N_1619,N_1691);
nor U2928 (N_2928,N_1298,N_1757);
or U2929 (N_2929,N_1758,N_1788);
nor U2930 (N_2930,N_1122,N_1362);
nand U2931 (N_2931,N_1621,N_1303);
and U2932 (N_2932,N_1371,N_1706);
nand U2933 (N_2933,N_1357,N_1790);
or U2934 (N_2934,N_1576,N_1899);
nor U2935 (N_2935,N_1515,N_1786);
nor U2936 (N_2936,N_1112,N_1295);
and U2937 (N_2937,N_1005,N_1121);
nand U2938 (N_2938,N_1721,N_1800);
and U2939 (N_2939,N_1632,N_1935);
nand U2940 (N_2940,N_1435,N_1841);
and U2941 (N_2941,N_1702,N_1993);
nand U2942 (N_2942,N_1415,N_1943);
nand U2943 (N_2943,N_1130,N_1257);
nor U2944 (N_2944,N_1837,N_1901);
and U2945 (N_2945,N_1091,N_1257);
or U2946 (N_2946,N_1848,N_1151);
or U2947 (N_2947,N_1721,N_1821);
and U2948 (N_2948,N_1709,N_1090);
nor U2949 (N_2949,N_1982,N_1782);
nand U2950 (N_2950,N_1753,N_1280);
nor U2951 (N_2951,N_1167,N_1775);
or U2952 (N_2952,N_1171,N_1865);
or U2953 (N_2953,N_1664,N_1465);
or U2954 (N_2954,N_1552,N_1246);
nor U2955 (N_2955,N_1059,N_1109);
nand U2956 (N_2956,N_1977,N_1740);
or U2957 (N_2957,N_1725,N_1527);
or U2958 (N_2958,N_1296,N_1918);
nand U2959 (N_2959,N_1102,N_1937);
nor U2960 (N_2960,N_1610,N_1428);
nand U2961 (N_2961,N_1018,N_1747);
nand U2962 (N_2962,N_1064,N_1670);
nand U2963 (N_2963,N_1563,N_1161);
or U2964 (N_2964,N_1439,N_1919);
nor U2965 (N_2965,N_1724,N_1971);
nor U2966 (N_2966,N_1831,N_1584);
nor U2967 (N_2967,N_1400,N_1765);
nor U2968 (N_2968,N_1097,N_1215);
nand U2969 (N_2969,N_1298,N_1045);
nor U2970 (N_2970,N_1850,N_1955);
or U2971 (N_2971,N_1006,N_1210);
or U2972 (N_2972,N_1912,N_1495);
or U2973 (N_2973,N_1234,N_1010);
and U2974 (N_2974,N_1781,N_1223);
nand U2975 (N_2975,N_1457,N_1688);
and U2976 (N_2976,N_1766,N_1579);
nand U2977 (N_2977,N_1942,N_1475);
nor U2978 (N_2978,N_1770,N_1368);
or U2979 (N_2979,N_1839,N_1107);
and U2980 (N_2980,N_1535,N_1646);
and U2981 (N_2981,N_1958,N_1899);
xor U2982 (N_2982,N_1296,N_1898);
nor U2983 (N_2983,N_1271,N_1629);
and U2984 (N_2984,N_1692,N_1056);
nand U2985 (N_2985,N_1786,N_1044);
and U2986 (N_2986,N_1066,N_1795);
nand U2987 (N_2987,N_1475,N_1862);
and U2988 (N_2988,N_1817,N_1039);
nand U2989 (N_2989,N_1656,N_1665);
and U2990 (N_2990,N_1565,N_1345);
nor U2991 (N_2991,N_1226,N_1299);
nand U2992 (N_2992,N_1677,N_1575);
nand U2993 (N_2993,N_1838,N_1245);
nor U2994 (N_2994,N_1951,N_1241);
nor U2995 (N_2995,N_1028,N_1817);
nor U2996 (N_2996,N_1680,N_1642);
and U2997 (N_2997,N_1326,N_1740);
nand U2998 (N_2998,N_1267,N_1597);
nor U2999 (N_2999,N_1186,N_1377);
or U3000 (N_3000,N_2806,N_2000);
nand U3001 (N_3001,N_2149,N_2599);
nand U3002 (N_3002,N_2694,N_2234);
nor U3003 (N_3003,N_2016,N_2221);
nor U3004 (N_3004,N_2103,N_2351);
nor U3005 (N_3005,N_2846,N_2436);
and U3006 (N_3006,N_2240,N_2706);
nor U3007 (N_3007,N_2156,N_2772);
or U3008 (N_3008,N_2708,N_2769);
nor U3009 (N_3009,N_2224,N_2515);
nor U3010 (N_3010,N_2774,N_2604);
nor U3011 (N_3011,N_2996,N_2329);
nor U3012 (N_3012,N_2181,N_2235);
and U3013 (N_3013,N_2114,N_2545);
nor U3014 (N_3014,N_2010,N_2294);
nand U3015 (N_3015,N_2736,N_2252);
or U3016 (N_3016,N_2731,N_2028);
nor U3017 (N_3017,N_2928,N_2402);
nor U3018 (N_3018,N_2423,N_2728);
nor U3019 (N_3019,N_2961,N_2897);
nand U3020 (N_3020,N_2442,N_2719);
nor U3021 (N_3021,N_2476,N_2607);
and U3022 (N_3022,N_2949,N_2984);
and U3023 (N_3023,N_2368,N_2095);
nor U3024 (N_3024,N_2723,N_2889);
or U3025 (N_3025,N_2173,N_2298);
and U3026 (N_3026,N_2781,N_2577);
xnor U3027 (N_3027,N_2504,N_2260);
nand U3028 (N_3028,N_2992,N_2033);
nand U3029 (N_3029,N_2524,N_2327);
nor U3030 (N_3030,N_2842,N_2051);
nand U3031 (N_3031,N_2013,N_2322);
nand U3032 (N_3032,N_2353,N_2315);
and U3033 (N_3033,N_2582,N_2486);
or U3034 (N_3034,N_2873,N_2112);
or U3035 (N_3035,N_2746,N_2779);
and U3036 (N_3036,N_2732,N_2912);
or U3037 (N_3037,N_2169,N_2118);
or U3038 (N_3038,N_2747,N_2784);
and U3039 (N_3039,N_2332,N_2501);
nor U3040 (N_3040,N_2271,N_2421);
nor U3041 (N_3041,N_2609,N_2280);
and U3042 (N_3042,N_2497,N_2080);
and U3043 (N_3043,N_2116,N_2291);
and U3044 (N_3044,N_2715,N_2552);
nand U3045 (N_3045,N_2935,N_2540);
and U3046 (N_3046,N_2324,N_2038);
nor U3047 (N_3047,N_2392,N_2069);
or U3048 (N_3048,N_2516,N_2771);
nor U3049 (N_3049,N_2496,N_2788);
nor U3050 (N_3050,N_2215,N_2418);
or U3051 (N_3051,N_2359,N_2020);
and U3052 (N_3052,N_2817,N_2677);
or U3053 (N_3053,N_2106,N_2342);
or U3054 (N_3054,N_2920,N_2239);
nand U3055 (N_3055,N_2693,N_2570);
and U3056 (N_3056,N_2888,N_2541);
nand U3057 (N_3057,N_2059,N_2440);
nand U3058 (N_3058,N_2659,N_2818);
or U3059 (N_3059,N_2441,N_2557);
nand U3060 (N_3060,N_2553,N_2437);
or U3061 (N_3061,N_2113,N_2244);
nand U3062 (N_3062,N_2823,N_2518);
or U3063 (N_3063,N_2575,N_2061);
or U3064 (N_3064,N_2339,N_2374);
nor U3065 (N_3065,N_2722,N_2197);
nand U3066 (N_3066,N_2633,N_2316);
nor U3067 (N_3067,N_2937,N_2132);
nor U3068 (N_3068,N_2355,N_2343);
nor U3069 (N_3069,N_2275,N_2981);
nand U3070 (N_3070,N_2473,N_2692);
or U3071 (N_3071,N_2201,N_2829);
nor U3072 (N_3072,N_2314,N_2675);
nor U3073 (N_3073,N_2001,N_2845);
and U3074 (N_3074,N_2308,N_2927);
and U3075 (N_3075,N_2695,N_2969);
and U3076 (N_3076,N_2810,N_2844);
nor U3077 (N_3077,N_2464,N_2670);
and U3078 (N_3078,N_2094,N_2566);
and U3079 (N_3079,N_2428,N_2972);
or U3080 (N_3080,N_2513,N_2931);
or U3081 (N_3081,N_2901,N_2556);
or U3082 (N_3082,N_2544,N_2596);
nand U3083 (N_3083,N_2372,N_2288);
nand U3084 (N_3084,N_2263,N_2373);
or U3085 (N_3085,N_2056,N_2024);
or U3086 (N_3086,N_2962,N_2292);
nand U3087 (N_3087,N_2579,N_2408);
nor U3088 (N_3088,N_2361,N_2131);
and U3089 (N_3089,N_2206,N_2711);
nor U3090 (N_3090,N_2395,N_2258);
or U3091 (N_3091,N_2347,N_2397);
and U3092 (N_3092,N_2537,N_2071);
and U3093 (N_3093,N_2470,N_2286);
or U3094 (N_3094,N_2958,N_2134);
nand U3095 (N_3095,N_2754,N_2145);
and U3096 (N_3096,N_2300,N_2519);
and U3097 (N_3097,N_2786,N_2750);
nor U3098 (N_3098,N_2186,N_2560);
nand U3099 (N_3099,N_2003,N_2220);
and U3100 (N_3100,N_2820,N_2008);
nand U3101 (N_3101,N_2041,N_2520);
nand U3102 (N_3102,N_2243,N_2539);
or U3103 (N_3103,N_2370,N_2994);
nand U3104 (N_3104,N_2768,N_2451);
or U3105 (N_3105,N_2232,N_2478);
and U3106 (N_3106,N_2611,N_2989);
nand U3107 (N_3107,N_2459,N_2574);
and U3108 (N_3108,N_2219,N_2046);
or U3109 (N_3109,N_2801,N_2336);
nand U3110 (N_3110,N_2667,N_2745);
nor U3111 (N_3111,N_2511,N_2642);
or U3112 (N_3112,N_2884,N_2109);
nand U3113 (N_3113,N_2689,N_2966);
nand U3114 (N_3114,N_2376,N_2320);
nand U3115 (N_3115,N_2489,N_2965);
nor U3116 (N_3116,N_2225,N_2724);
and U3117 (N_3117,N_2554,N_2123);
and U3118 (N_3118,N_2849,N_2763);
nor U3119 (N_3119,N_2696,N_2644);
and U3120 (N_3120,N_2472,N_2267);
and U3121 (N_3121,N_2254,N_2012);
nand U3122 (N_3122,N_2076,N_2507);
nor U3123 (N_3123,N_2494,N_2569);
and U3124 (N_3124,N_2455,N_2025);
nor U3125 (N_3125,N_2620,N_2680);
nor U3126 (N_3126,N_2624,N_2682);
and U3127 (N_3127,N_2616,N_2563);
or U3128 (N_3128,N_2142,N_2299);
nand U3129 (N_3129,N_2521,N_2727);
or U3130 (N_3130,N_2814,N_2301);
nand U3131 (N_3131,N_2531,N_2625);
nor U3132 (N_3132,N_2952,N_2629);
nand U3133 (N_3133,N_2483,N_2165);
and U3134 (N_3134,N_2793,N_2363);
and U3135 (N_3135,N_2617,N_2063);
or U3136 (N_3136,N_2757,N_2583);
and U3137 (N_3137,N_2939,N_2042);
nand U3138 (N_3138,N_2783,N_2111);
nand U3139 (N_3139,N_2861,N_2345);
and U3140 (N_3140,N_2088,N_2499);
or U3141 (N_3141,N_2229,N_2654);
and U3142 (N_3142,N_2782,N_2866);
and U3143 (N_3143,N_2333,N_2104);
nor U3144 (N_3144,N_2168,N_2307);
or U3145 (N_3145,N_2124,N_2641);
nand U3146 (N_3146,N_2188,N_2096);
nand U3147 (N_3147,N_2933,N_2050);
nand U3148 (N_3148,N_2990,N_2598);
nor U3149 (N_3149,N_2681,N_2434);
nand U3150 (N_3150,N_2973,N_2941);
nand U3151 (N_3151,N_2488,N_2004);
or U3152 (N_3152,N_2627,N_2205);
nor U3153 (N_3153,N_2837,N_2283);
nand U3154 (N_3154,N_2256,N_2527);
or U3155 (N_3155,N_2503,N_2075);
and U3156 (N_3156,N_2573,N_2883);
nor U3157 (N_3157,N_2491,N_2160);
or U3158 (N_3158,N_2601,N_2546);
nand U3159 (N_3159,N_2863,N_2517);
and U3160 (N_3160,N_2321,N_2404);
and U3161 (N_3161,N_2709,N_2018);
or U3162 (N_3162,N_2887,N_2212);
nand U3163 (N_3163,N_2506,N_2121);
or U3164 (N_3164,N_2652,N_2533);
or U3165 (N_3165,N_2279,N_2964);
nor U3166 (N_3166,N_2792,N_2128);
nand U3167 (N_3167,N_2637,N_2296);
nor U3168 (N_3168,N_2017,N_2306);
or U3169 (N_3169,N_2910,N_2335);
nand U3170 (N_3170,N_2334,N_2730);
or U3171 (N_3171,N_2185,N_2535);
nor U3172 (N_3172,N_2934,N_2362);
and U3173 (N_3173,N_2622,N_2276);
nor U3174 (N_3174,N_2151,N_2699);
or U3175 (N_3175,N_2077,N_2083);
and U3176 (N_3176,N_2740,N_2485);
or U3177 (N_3177,N_2490,N_2295);
nand U3178 (N_3178,N_2191,N_2893);
or U3179 (N_3179,N_2136,N_2751);
or U3180 (N_3180,N_2448,N_2936);
or U3181 (N_3181,N_2975,N_2636);
nand U3182 (N_3182,N_2761,N_2385);
nor U3183 (N_3183,N_2214,N_2991);
nor U3184 (N_3184,N_2146,N_2857);
nor U3185 (N_3185,N_2415,N_2281);
nor U3186 (N_3186,N_2364,N_2492);
or U3187 (N_3187,N_2119,N_2957);
or U3188 (N_3188,N_2498,N_2600);
nor U3189 (N_3189,N_2945,N_2053);
nand U3190 (N_3190,N_2237,N_2278);
nand U3191 (N_3191,N_2974,N_2311);
nand U3192 (N_3192,N_2477,N_2386);
or U3193 (N_3193,N_2407,N_2683);
or U3194 (N_3194,N_2564,N_2980);
and U3195 (N_3195,N_2812,N_2725);
nand U3196 (N_3196,N_2615,N_2797);
nand U3197 (N_3197,N_2815,N_2867);
nor U3198 (N_3198,N_2997,N_2389);
nand U3199 (N_3199,N_2838,N_2590);
nor U3200 (N_3200,N_2179,N_2729);
nand U3201 (N_3201,N_2847,N_2851);
or U3202 (N_3202,N_2836,N_2274);
or U3203 (N_3203,N_2377,N_2647);
or U3204 (N_3204,N_2799,N_2534);
and U3205 (N_3205,N_2460,N_2398);
nand U3206 (N_3206,N_2217,N_2192);
and U3207 (N_3207,N_2753,N_2326);
nand U3208 (N_3208,N_2900,N_2164);
and U3209 (N_3209,N_2828,N_2986);
and U3210 (N_3210,N_2850,N_2338);
nor U3211 (N_3211,N_2585,N_2551);
and U3212 (N_3212,N_2422,N_2198);
and U3213 (N_3213,N_2955,N_2942);
or U3214 (N_3214,N_2021,N_2303);
or U3215 (N_3215,N_2125,N_2657);
nor U3216 (N_3216,N_2171,N_2621);
nor U3217 (N_3217,N_2152,N_2686);
or U3218 (N_3218,N_2858,N_2035);
nand U3219 (N_3219,N_2227,N_2054);
or U3220 (N_3220,N_2938,N_2648);
or U3221 (N_3221,N_2147,N_2268);
or U3222 (N_3222,N_2576,N_2571);
nor U3223 (N_3223,N_2133,N_2098);
and U3224 (N_3224,N_2394,N_2525);
and U3225 (N_3225,N_2218,N_2161);
nor U3226 (N_3226,N_2758,N_2453);
and U3227 (N_3227,N_2302,N_2187);
or U3228 (N_3228,N_2045,N_2174);
or U3229 (N_3229,N_2650,N_2403);
or U3230 (N_3230,N_2505,N_2369);
or U3231 (N_3231,N_2452,N_2944);
and U3232 (N_3232,N_2854,N_2791);
or U3233 (N_3233,N_2108,N_2172);
or U3234 (N_3234,N_2047,N_2420);
nand U3235 (N_3235,N_2500,N_2284);
or U3236 (N_3236,N_2137,N_2262);
or U3237 (N_3237,N_2917,N_2919);
nor U3238 (N_3238,N_2406,N_2663);
or U3239 (N_3239,N_2091,N_2270);
or U3240 (N_3240,N_2795,N_2809);
and U3241 (N_3241,N_2638,N_2447);
nand U3242 (N_3242,N_2610,N_2261);
nor U3243 (N_3243,N_2899,N_2482);
or U3244 (N_3244,N_2862,N_2446);
nor U3245 (N_3245,N_2805,N_2387);
or U3246 (N_3246,N_2122,N_2821);
nor U3247 (N_3247,N_2684,N_2717);
nor U3248 (N_3248,N_2383,N_2926);
and U3249 (N_3249,N_2413,N_2399);
nor U3250 (N_3250,N_2932,N_2841);
or U3251 (N_3251,N_2568,N_2668);
xor U3252 (N_3252,N_2162,N_2129);
and U3253 (N_3253,N_2230,N_2705);
nand U3254 (N_3254,N_2742,N_2208);
and U3255 (N_3255,N_2767,N_2738);
or U3256 (N_3256,N_2330,N_2340);
or U3257 (N_3257,N_2360,N_2101);
and U3258 (N_3258,N_2060,N_2228);
or U3259 (N_3259,N_2643,N_2246);
and U3260 (N_3260,N_2860,N_2049);
nor U3261 (N_3261,N_2855,N_2840);
xnor U3262 (N_3262,N_2948,N_2803);
nor U3263 (N_3263,N_2796,N_2678);
or U3264 (N_3264,N_2744,N_2735);
or U3265 (N_3265,N_2921,N_2202);
nand U3266 (N_3266,N_2086,N_2209);
or U3267 (N_3267,N_2737,N_2529);
nand U3268 (N_3268,N_2318,N_2923);
or U3269 (N_3269,N_2027,N_2469);
nand U3270 (N_3270,N_2449,N_2640);
or U3271 (N_3271,N_2238,N_2143);
and U3272 (N_3272,N_2040,N_2593);
nor U3273 (N_3273,N_2223,N_2264);
or U3274 (N_3274,N_2183,N_2366);
and U3275 (N_3275,N_2831,N_2170);
and U3276 (N_3276,N_2586,N_2908);
or U3277 (N_3277,N_2210,N_2481);
nand U3278 (N_3278,N_2471,N_2733);
or U3279 (N_3279,N_2127,N_2073);
nor U3280 (N_3280,N_2430,N_2319);
and U3281 (N_3281,N_2072,N_2019);
or U3282 (N_3282,N_2358,N_2995);
and U3283 (N_3283,N_2068,N_2748);
nand U3284 (N_3284,N_2848,N_2178);
nand U3285 (N_3285,N_2512,N_2685);
and U3286 (N_3286,N_2026,N_2269);
and U3287 (N_3287,N_2594,N_2153);
nor U3288 (N_3288,N_2656,N_2247);
nor U3289 (N_3289,N_2508,N_2043);
nand U3290 (N_3290,N_2337,N_2480);
or U3291 (N_3291,N_2561,N_2804);
nor U3292 (N_3292,N_2463,N_2959);
nor U3293 (N_3293,N_2832,N_2597);
and U3294 (N_3294,N_2780,N_2743);
nor U3295 (N_3295,N_2005,N_2929);
or U3296 (N_3296,N_2734,N_2388);
and U3297 (N_3297,N_2493,N_2305);
nand U3298 (N_3298,N_2189,N_2802);
nand U3299 (N_3299,N_2628,N_2065);
and U3300 (N_3300,N_2658,N_2079);
and U3301 (N_3301,N_2431,N_2871);
or U3302 (N_3302,N_2349,N_2450);
and U3303 (N_3303,N_2317,N_2639);
nor U3304 (N_3304,N_2207,N_2352);
and U3305 (N_3305,N_2988,N_2902);
or U3306 (N_3306,N_2175,N_2196);
nor U3307 (N_3307,N_2752,N_2764);
and U3308 (N_3308,N_2588,N_2182);
nand U3309 (N_3309,N_2242,N_2954);
nor U3310 (N_3310,N_2584,N_2023);
nor U3311 (N_3311,N_2067,N_2869);
or U3312 (N_3312,N_2309,N_2562);
nor U3313 (N_3313,N_2265,N_2914);
nor U3314 (N_3314,N_2662,N_2213);
nand U3315 (N_3315,N_2474,N_2632);
nor U3316 (N_3316,N_2466,N_2089);
nand U3317 (N_3317,N_2378,N_2697);
nand U3318 (N_3318,N_2608,N_2924);
nand U3319 (N_3319,N_2688,N_2110);
or U3320 (N_3320,N_2475,N_2915);
nand U3321 (N_3321,N_2393,N_2798);
or U3322 (N_3322,N_2367,N_2282);
and U3323 (N_3323,N_2950,N_2141);
nor U3324 (N_3324,N_2726,N_2785);
xnor U3325 (N_3325,N_2911,N_2827);
or U3326 (N_3326,N_2140,N_2177);
nand U3327 (N_3327,N_2328,N_2755);
nor U3328 (N_3328,N_2167,N_2093);
and U3329 (N_3329,N_2396,N_2158);
or U3330 (N_3330,N_2536,N_2248);
or U3331 (N_3331,N_2789,N_2903);
nand U3332 (N_3332,N_2031,N_2864);
xor U3333 (N_3333,N_2435,N_2547);
nor U3334 (N_3334,N_2649,N_2672);
or U3335 (N_3335,N_2983,N_2424);
and U3336 (N_3336,N_2011,N_2679);
nor U3337 (N_3337,N_2700,N_2391);
and U3338 (N_3338,N_2555,N_2414);
nor U3339 (N_3339,N_2312,N_2843);
nand U3340 (N_3340,N_2707,N_2289);
nor U3341 (N_3341,N_2819,N_2985);
nand U3342 (N_3342,N_2532,N_2651);
nor U3343 (N_3343,N_2906,N_2787);
nor U3344 (N_3344,N_2691,N_2790);
or U3345 (N_3345,N_2885,N_2951);
nor U3346 (N_3346,N_2454,N_2226);
and U3347 (N_3347,N_2375,N_2412);
and U3348 (N_3348,N_2635,N_2890);
nand U3349 (N_3349,N_2417,N_2467);
nor U3350 (N_3350,N_2712,N_2749);
or U3351 (N_3351,N_2138,N_2419);
nand U3352 (N_3352,N_2390,N_2956);
nand U3353 (N_3353,N_2444,N_2022);
nand U3354 (N_3354,N_2613,N_2509);
or U3355 (N_3355,N_2405,N_2331);
or U3356 (N_3356,N_2007,N_2154);
or U3357 (N_3357,N_2578,N_2287);
nand U3358 (N_3358,N_2245,N_2999);
or U3359 (N_3359,N_2055,N_2826);
nor U3360 (N_3360,N_2909,N_2126);
nand U3361 (N_3361,N_2970,N_2427);
and U3362 (N_3362,N_2120,N_2105);
nand U3363 (N_3363,N_2117,N_2548);
or U3364 (N_3364,N_2665,N_2892);
nor U3365 (N_3365,N_2550,N_2203);
or U3366 (N_3366,N_2380,N_2543);
nand U3367 (N_3367,N_2631,N_2716);
and U3368 (N_3368,N_2993,N_2037);
and U3369 (N_3369,N_2510,N_2409);
or U3370 (N_3370,N_2479,N_2765);
nand U3371 (N_3371,N_2882,N_2874);
or U3372 (N_3372,N_2718,N_2704);
nand U3373 (N_3373,N_2382,N_2673);
or U3374 (N_3374,N_2411,N_2379);
nor U3375 (N_3375,N_2344,N_2676);
nor U3376 (N_3376,N_2350,N_2904);
nand U3377 (N_3377,N_2445,N_2487);
or U3378 (N_3378,N_2293,N_2356);
and U3379 (N_3379,N_2878,N_2484);
nor U3380 (N_3380,N_2222,N_2960);
nor U3381 (N_3381,N_2835,N_2630);
nand U3382 (N_3382,N_2664,N_2014);
or U3383 (N_3383,N_2090,N_2834);
or U3384 (N_3384,N_2528,N_2870);
nor U3385 (N_3385,N_2634,N_2432);
and U3386 (N_3386,N_2538,N_2253);
nor U3387 (N_3387,N_2830,N_2015);
or U3388 (N_3388,N_2940,N_2313);
nand U3389 (N_3389,N_2775,N_2297);
xor U3390 (N_3390,N_2304,N_2410);
xnor U3391 (N_3391,N_2916,N_2092);
or U3392 (N_3392,N_2323,N_2502);
and U3393 (N_3393,N_2868,N_2967);
or U3394 (N_3394,N_2953,N_2881);
xor U3395 (N_3395,N_2354,N_2925);
nand U3396 (N_3396,N_2907,N_2690);
nand U3397 (N_3397,N_2930,N_2074);
or U3398 (N_3398,N_2236,N_2852);
or U3399 (N_3399,N_2891,N_2211);
and U3400 (N_3400,N_2429,N_2619);
nand U3401 (N_3401,N_2439,N_2400);
or U3402 (N_3402,N_2759,N_2807);
nor U3403 (N_3403,N_2886,N_2381);
nand U3404 (N_3404,N_2070,N_2044);
nand U3405 (N_3405,N_2762,N_2655);
nor U3406 (N_3406,N_2872,N_2348);
or U3407 (N_3407,N_2800,N_2052);
and U3408 (N_3408,N_2987,N_2875);
nor U3409 (N_3409,N_2603,N_2231);
or U3410 (N_3410,N_2894,N_2272);
and U3411 (N_3411,N_2064,N_2710);
or U3412 (N_3412,N_2457,N_2002);
nor U3413 (N_3413,N_2963,N_2666);
or U3414 (N_3414,N_2241,N_2193);
and U3415 (N_3415,N_2346,N_2200);
or U3416 (N_3416,N_2032,N_2671);
and U3417 (N_3417,N_2426,N_2880);
or U3418 (N_3418,N_2739,N_2825);
nor U3419 (N_3419,N_2034,N_2465);
nand U3420 (N_3420,N_2943,N_2581);
or U3421 (N_3421,N_2559,N_2646);
and U3422 (N_3422,N_2078,N_2947);
and U3423 (N_3423,N_2039,N_2946);
or U3424 (N_3424,N_2194,N_2233);
xor U3425 (N_3425,N_2107,N_2898);
nor U3426 (N_3426,N_2130,N_2259);
and U3427 (N_3427,N_2567,N_2918);
and U3428 (N_3428,N_2922,N_2602);
or U3429 (N_3429,N_2565,N_2176);
or U3430 (N_3430,N_2580,N_2085);
or U3431 (N_3431,N_2687,N_2180);
and U3432 (N_3432,N_2251,N_2100);
nor U3433 (N_3433,N_2163,N_2057);
and U3434 (N_3434,N_2605,N_2285);
nand U3435 (N_3435,N_2905,N_2660);
nand U3436 (N_3436,N_2756,N_2614);
and U3437 (N_3437,N_2144,N_2066);
or U3438 (N_3438,N_2591,N_2184);
and U3439 (N_3439,N_2653,N_2526);
nor U3440 (N_3440,N_2458,N_2273);
or U3441 (N_3441,N_2084,N_2859);
nor U3442 (N_3442,N_2097,N_2514);
nand U3443 (N_3443,N_2009,N_2572);
and U3444 (N_3444,N_2876,N_2384);
or U3445 (N_3445,N_2778,N_2341);
or U3446 (N_3446,N_2062,N_2606);
nor U3447 (N_3447,N_2102,N_2618);
and U3448 (N_3448,N_2626,N_2853);
and U3449 (N_3449,N_2982,N_2865);
or U3450 (N_3450,N_2760,N_2674);
and U3451 (N_3451,N_2099,N_2416);
nor U3452 (N_3452,N_2816,N_2155);
or U3453 (N_3453,N_2773,N_2777);
or U3454 (N_3454,N_2468,N_2115);
nor U3455 (N_3455,N_2856,N_2813);
nand U3456 (N_3456,N_2462,N_2216);
and U3457 (N_3457,N_2461,N_2645);
nor U3458 (N_3458,N_2433,N_2794);
nor U3459 (N_3459,N_2166,N_2595);
nand U3460 (N_3460,N_2425,N_2082);
and U3461 (N_3461,N_2589,N_2978);
and U3462 (N_3462,N_2542,N_2776);
xnor U3463 (N_3463,N_2895,N_2592);
nor U3464 (N_3464,N_2839,N_2523);
nor U3465 (N_3465,N_2811,N_2150);
and U3466 (N_3466,N_2741,N_2702);
or U3467 (N_3467,N_2714,N_2558);
and U3468 (N_3468,N_2770,N_2877);
and U3469 (N_3469,N_2087,N_2979);
and U3470 (N_3470,N_2968,N_2721);
nand U3471 (N_3471,N_2157,N_2058);
nor U3472 (N_3472,N_2250,N_2443);
and U3473 (N_3473,N_2456,N_2204);
nand U3474 (N_3474,N_2896,N_2703);
and U3475 (N_3475,N_2824,N_2310);
nor U3476 (N_3476,N_2401,N_2255);
nor U3477 (N_3477,N_2290,N_2495);
nand U3478 (N_3478,N_2530,N_2998);
or U3479 (N_3479,N_2036,N_2522);
nand U3480 (N_3480,N_2195,N_2257);
or U3481 (N_3481,N_2159,N_2365);
nor U3482 (N_3482,N_2190,N_2371);
or U3483 (N_3483,N_2249,N_2612);
nor U3484 (N_3484,N_2913,N_2808);
and U3485 (N_3485,N_2135,N_2698);
xnor U3486 (N_3486,N_2669,N_2976);
nor U3487 (N_3487,N_2030,N_2587);
or U3488 (N_3488,N_2199,N_2879);
nand U3489 (N_3489,N_2822,N_2148);
and U3490 (N_3490,N_2048,N_2549);
nor U3491 (N_3491,N_2139,N_2833);
nand U3492 (N_3492,N_2720,N_2701);
and U3493 (N_3493,N_2661,N_2006);
nor U3494 (N_3494,N_2971,N_2266);
nor U3495 (N_3495,N_2357,N_2977);
and U3496 (N_3496,N_2277,N_2623);
nand U3497 (N_3497,N_2029,N_2325);
nand U3498 (N_3498,N_2081,N_2766);
xor U3499 (N_3499,N_2438,N_2713);
nor U3500 (N_3500,N_2406,N_2360);
xnor U3501 (N_3501,N_2804,N_2367);
or U3502 (N_3502,N_2572,N_2945);
and U3503 (N_3503,N_2433,N_2971);
or U3504 (N_3504,N_2075,N_2007);
nor U3505 (N_3505,N_2431,N_2425);
or U3506 (N_3506,N_2667,N_2174);
nand U3507 (N_3507,N_2702,N_2361);
and U3508 (N_3508,N_2910,N_2047);
nor U3509 (N_3509,N_2171,N_2821);
and U3510 (N_3510,N_2315,N_2751);
nand U3511 (N_3511,N_2222,N_2648);
nor U3512 (N_3512,N_2050,N_2876);
and U3513 (N_3513,N_2672,N_2429);
nand U3514 (N_3514,N_2706,N_2560);
nor U3515 (N_3515,N_2035,N_2925);
nand U3516 (N_3516,N_2049,N_2474);
and U3517 (N_3517,N_2650,N_2390);
and U3518 (N_3518,N_2360,N_2652);
nand U3519 (N_3519,N_2496,N_2660);
or U3520 (N_3520,N_2921,N_2370);
or U3521 (N_3521,N_2959,N_2865);
nor U3522 (N_3522,N_2204,N_2906);
nor U3523 (N_3523,N_2256,N_2964);
or U3524 (N_3524,N_2995,N_2712);
or U3525 (N_3525,N_2047,N_2273);
and U3526 (N_3526,N_2847,N_2899);
or U3527 (N_3527,N_2112,N_2870);
nand U3528 (N_3528,N_2437,N_2582);
nor U3529 (N_3529,N_2415,N_2429);
nor U3530 (N_3530,N_2071,N_2988);
or U3531 (N_3531,N_2830,N_2579);
nor U3532 (N_3532,N_2994,N_2738);
and U3533 (N_3533,N_2033,N_2014);
nand U3534 (N_3534,N_2851,N_2369);
and U3535 (N_3535,N_2333,N_2077);
or U3536 (N_3536,N_2172,N_2799);
nand U3537 (N_3537,N_2406,N_2299);
nand U3538 (N_3538,N_2155,N_2818);
and U3539 (N_3539,N_2627,N_2988);
nor U3540 (N_3540,N_2082,N_2139);
and U3541 (N_3541,N_2058,N_2269);
or U3542 (N_3542,N_2646,N_2442);
and U3543 (N_3543,N_2219,N_2302);
and U3544 (N_3544,N_2372,N_2052);
and U3545 (N_3545,N_2010,N_2179);
nor U3546 (N_3546,N_2188,N_2788);
nand U3547 (N_3547,N_2677,N_2453);
nor U3548 (N_3548,N_2186,N_2122);
nand U3549 (N_3549,N_2690,N_2694);
nor U3550 (N_3550,N_2059,N_2720);
and U3551 (N_3551,N_2473,N_2975);
or U3552 (N_3552,N_2718,N_2085);
nor U3553 (N_3553,N_2612,N_2232);
nor U3554 (N_3554,N_2458,N_2404);
and U3555 (N_3555,N_2332,N_2808);
and U3556 (N_3556,N_2411,N_2098);
and U3557 (N_3557,N_2376,N_2056);
nor U3558 (N_3558,N_2169,N_2481);
nor U3559 (N_3559,N_2766,N_2299);
nor U3560 (N_3560,N_2450,N_2681);
or U3561 (N_3561,N_2452,N_2039);
nor U3562 (N_3562,N_2103,N_2533);
nor U3563 (N_3563,N_2551,N_2708);
or U3564 (N_3564,N_2366,N_2333);
nand U3565 (N_3565,N_2882,N_2472);
or U3566 (N_3566,N_2145,N_2918);
nand U3567 (N_3567,N_2936,N_2861);
nand U3568 (N_3568,N_2336,N_2264);
or U3569 (N_3569,N_2058,N_2323);
or U3570 (N_3570,N_2987,N_2673);
nand U3571 (N_3571,N_2414,N_2610);
xor U3572 (N_3572,N_2359,N_2546);
and U3573 (N_3573,N_2657,N_2737);
nand U3574 (N_3574,N_2350,N_2554);
and U3575 (N_3575,N_2890,N_2716);
nand U3576 (N_3576,N_2319,N_2536);
nand U3577 (N_3577,N_2650,N_2988);
nor U3578 (N_3578,N_2263,N_2505);
nor U3579 (N_3579,N_2270,N_2059);
and U3580 (N_3580,N_2679,N_2377);
or U3581 (N_3581,N_2630,N_2958);
or U3582 (N_3582,N_2371,N_2855);
nor U3583 (N_3583,N_2640,N_2448);
nand U3584 (N_3584,N_2898,N_2191);
nor U3585 (N_3585,N_2778,N_2909);
or U3586 (N_3586,N_2349,N_2525);
nand U3587 (N_3587,N_2118,N_2381);
nand U3588 (N_3588,N_2746,N_2380);
nor U3589 (N_3589,N_2389,N_2951);
nor U3590 (N_3590,N_2634,N_2551);
and U3591 (N_3591,N_2134,N_2487);
nor U3592 (N_3592,N_2232,N_2635);
and U3593 (N_3593,N_2764,N_2183);
nand U3594 (N_3594,N_2310,N_2262);
and U3595 (N_3595,N_2021,N_2347);
nand U3596 (N_3596,N_2718,N_2368);
nor U3597 (N_3597,N_2644,N_2440);
or U3598 (N_3598,N_2723,N_2676);
or U3599 (N_3599,N_2167,N_2059);
or U3600 (N_3600,N_2458,N_2124);
nand U3601 (N_3601,N_2430,N_2582);
nor U3602 (N_3602,N_2961,N_2233);
nand U3603 (N_3603,N_2892,N_2315);
nor U3604 (N_3604,N_2921,N_2450);
nand U3605 (N_3605,N_2914,N_2603);
xnor U3606 (N_3606,N_2433,N_2282);
nor U3607 (N_3607,N_2966,N_2360);
or U3608 (N_3608,N_2097,N_2925);
nor U3609 (N_3609,N_2910,N_2065);
and U3610 (N_3610,N_2112,N_2723);
or U3611 (N_3611,N_2433,N_2071);
nand U3612 (N_3612,N_2115,N_2069);
nor U3613 (N_3613,N_2865,N_2067);
or U3614 (N_3614,N_2780,N_2990);
or U3615 (N_3615,N_2655,N_2951);
nor U3616 (N_3616,N_2012,N_2044);
nor U3617 (N_3617,N_2405,N_2458);
nor U3618 (N_3618,N_2108,N_2276);
nor U3619 (N_3619,N_2082,N_2954);
nor U3620 (N_3620,N_2868,N_2812);
and U3621 (N_3621,N_2245,N_2868);
nand U3622 (N_3622,N_2144,N_2593);
nand U3623 (N_3623,N_2750,N_2430);
or U3624 (N_3624,N_2503,N_2729);
nor U3625 (N_3625,N_2995,N_2167);
nand U3626 (N_3626,N_2612,N_2889);
nand U3627 (N_3627,N_2176,N_2148);
nor U3628 (N_3628,N_2510,N_2428);
and U3629 (N_3629,N_2130,N_2509);
nor U3630 (N_3630,N_2303,N_2367);
nand U3631 (N_3631,N_2095,N_2744);
nand U3632 (N_3632,N_2405,N_2697);
or U3633 (N_3633,N_2633,N_2025);
nor U3634 (N_3634,N_2035,N_2427);
and U3635 (N_3635,N_2409,N_2799);
and U3636 (N_3636,N_2036,N_2489);
and U3637 (N_3637,N_2375,N_2023);
and U3638 (N_3638,N_2579,N_2211);
and U3639 (N_3639,N_2055,N_2629);
or U3640 (N_3640,N_2752,N_2937);
and U3641 (N_3641,N_2743,N_2339);
and U3642 (N_3642,N_2603,N_2614);
and U3643 (N_3643,N_2405,N_2153);
nand U3644 (N_3644,N_2266,N_2486);
nand U3645 (N_3645,N_2597,N_2503);
nand U3646 (N_3646,N_2908,N_2729);
and U3647 (N_3647,N_2858,N_2250);
and U3648 (N_3648,N_2644,N_2505);
or U3649 (N_3649,N_2074,N_2083);
or U3650 (N_3650,N_2718,N_2273);
or U3651 (N_3651,N_2971,N_2959);
nand U3652 (N_3652,N_2888,N_2898);
and U3653 (N_3653,N_2883,N_2050);
nor U3654 (N_3654,N_2842,N_2430);
or U3655 (N_3655,N_2397,N_2654);
nand U3656 (N_3656,N_2242,N_2482);
nor U3657 (N_3657,N_2908,N_2336);
and U3658 (N_3658,N_2330,N_2546);
or U3659 (N_3659,N_2022,N_2493);
and U3660 (N_3660,N_2660,N_2255);
or U3661 (N_3661,N_2330,N_2920);
nand U3662 (N_3662,N_2834,N_2757);
and U3663 (N_3663,N_2848,N_2024);
or U3664 (N_3664,N_2038,N_2421);
nand U3665 (N_3665,N_2261,N_2908);
nand U3666 (N_3666,N_2817,N_2594);
or U3667 (N_3667,N_2607,N_2876);
nand U3668 (N_3668,N_2968,N_2630);
and U3669 (N_3669,N_2760,N_2713);
nand U3670 (N_3670,N_2423,N_2428);
nor U3671 (N_3671,N_2642,N_2652);
nor U3672 (N_3672,N_2007,N_2333);
or U3673 (N_3673,N_2235,N_2815);
or U3674 (N_3674,N_2650,N_2303);
nand U3675 (N_3675,N_2216,N_2388);
nor U3676 (N_3676,N_2032,N_2949);
and U3677 (N_3677,N_2351,N_2727);
and U3678 (N_3678,N_2218,N_2600);
nor U3679 (N_3679,N_2215,N_2250);
or U3680 (N_3680,N_2459,N_2861);
nor U3681 (N_3681,N_2038,N_2960);
and U3682 (N_3682,N_2918,N_2608);
and U3683 (N_3683,N_2806,N_2842);
and U3684 (N_3684,N_2811,N_2396);
nor U3685 (N_3685,N_2723,N_2067);
and U3686 (N_3686,N_2842,N_2998);
nor U3687 (N_3687,N_2950,N_2097);
and U3688 (N_3688,N_2250,N_2130);
and U3689 (N_3689,N_2129,N_2385);
nor U3690 (N_3690,N_2646,N_2768);
nand U3691 (N_3691,N_2583,N_2037);
and U3692 (N_3692,N_2766,N_2784);
and U3693 (N_3693,N_2681,N_2374);
nor U3694 (N_3694,N_2645,N_2871);
nor U3695 (N_3695,N_2837,N_2112);
and U3696 (N_3696,N_2539,N_2123);
nor U3697 (N_3697,N_2879,N_2035);
nand U3698 (N_3698,N_2621,N_2743);
nor U3699 (N_3699,N_2933,N_2201);
nand U3700 (N_3700,N_2682,N_2339);
or U3701 (N_3701,N_2711,N_2821);
or U3702 (N_3702,N_2865,N_2575);
nand U3703 (N_3703,N_2240,N_2484);
nand U3704 (N_3704,N_2198,N_2672);
nor U3705 (N_3705,N_2806,N_2794);
nand U3706 (N_3706,N_2137,N_2637);
nor U3707 (N_3707,N_2579,N_2606);
and U3708 (N_3708,N_2840,N_2500);
nand U3709 (N_3709,N_2650,N_2369);
or U3710 (N_3710,N_2847,N_2557);
nand U3711 (N_3711,N_2938,N_2039);
nor U3712 (N_3712,N_2977,N_2321);
nand U3713 (N_3713,N_2490,N_2170);
nand U3714 (N_3714,N_2966,N_2514);
or U3715 (N_3715,N_2851,N_2398);
nand U3716 (N_3716,N_2091,N_2613);
nand U3717 (N_3717,N_2882,N_2634);
and U3718 (N_3718,N_2430,N_2877);
nand U3719 (N_3719,N_2832,N_2272);
or U3720 (N_3720,N_2225,N_2380);
and U3721 (N_3721,N_2757,N_2362);
or U3722 (N_3722,N_2257,N_2128);
or U3723 (N_3723,N_2120,N_2020);
or U3724 (N_3724,N_2049,N_2064);
and U3725 (N_3725,N_2514,N_2515);
nor U3726 (N_3726,N_2784,N_2206);
or U3727 (N_3727,N_2781,N_2492);
or U3728 (N_3728,N_2883,N_2945);
or U3729 (N_3729,N_2654,N_2863);
or U3730 (N_3730,N_2968,N_2173);
nand U3731 (N_3731,N_2226,N_2591);
nand U3732 (N_3732,N_2284,N_2551);
nor U3733 (N_3733,N_2862,N_2949);
and U3734 (N_3734,N_2403,N_2250);
nand U3735 (N_3735,N_2660,N_2647);
and U3736 (N_3736,N_2944,N_2511);
nand U3737 (N_3737,N_2895,N_2827);
and U3738 (N_3738,N_2959,N_2222);
nand U3739 (N_3739,N_2388,N_2814);
and U3740 (N_3740,N_2758,N_2227);
or U3741 (N_3741,N_2351,N_2321);
nor U3742 (N_3742,N_2612,N_2983);
and U3743 (N_3743,N_2528,N_2915);
nor U3744 (N_3744,N_2024,N_2017);
nand U3745 (N_3745,N_2751,N_2062);
nand U3746 (N_3746,N_2391,N_2318);
or U3747 (N_3747,N_2087,N_2724);
nand U3748 (N_3748,N_2828,N_2021);
and U3749 (N_3749,N_2739,N_2481);
nand U3750 (N_3750,N_2121,N_2170);
and U3751 (N_3751,N_2123,N_2903);
nor U3752 (N_3752,N_2491,N_2275);
or U3753 (N_3753,N_2946,N_2664);
and U3754 (N_3754,N_2791,N_2247);
or U3755 (N_3755,N_2876,N_2109);
nand U3756 (N_3756,N_2168,N_2443);
or U3757 (N_3757,N_2965,N_2812);
and U3758 (N_3758,N_2314,N_2601);
or U3759 (N_3759,N_2608,N_2082);
nor U3760 (N_3760,N_2660,N_2475);
xnor U3761 (N_3761,N_2621,N_2495);
or U3762 (N_3762,N_2995,N_2883);
or U3763 (N_3763,N_2862,N_2193);
xnor U3764 (N_3764,N_2719,N_2220);
nor U3765 (N_3765,N_2907,N_2076);
nand U3766 (N_3766,N_2954,N_2120);
and U3767 (N_3767,N_2409,N_2685);
nor U3768 (N_3768,N_2110,N_2695);
and U3769 (N_3769,N_2126,N_2953);
and U3770 (N_3770,N_2210,N_2748);
nand U3771 (N_3771,N_2180,N_2311);
nor U3772 (N_3772,N_2007,N_2721);
and U3773 (N_3773,N_2679,N_2191);
nand U3774 (N_3774,N_2135,N_2546);
nand U3775 (N_3775,N_2888,N_2915);
nand U3776 (N_3776,N_2103,N_2225);
or U3777 (N_3777,N_2174,N_2685);
nor U3778 (N_3778,N_2936,N_2181);
and U3779 (N_3779,N_2117,N_2417);
xor U3780 (N_3780,N_2977,N_2244);
or U3781 (N_3781,N_2677,N_2615);
nor U3782 (N_3782,N_2640,N_2473);
and U3783 (N_3783,N_2366,N_2558);
nand U3784 (N_3784,N_2666,N_2168);
and U3785 (N_3785,N_2275,N_2273);
or U3786 (N_3786,N_2667,N_2851);
nand U3787 (N_3787,N_2622,N_2104);
and U3788 (N_3788,N_2929,N_2397);
nor U3789 (N_3789,N_2550,N_2072);
nor U3790 (N_3790,N_2695,N_2166);
and U3791 (N_3791,N_2146,N_2700);
nand U3792 (N_3792,N_2572,N_2085);
nor U3793 (N_3793,N_2560,N_2300);
nor U3794 (N_3794,N_2335,N_2065);
and U3795 (N_3795,N_2633,N_2739);
or U3796 (N_3796,N_2090,N_2537);
and U3797 (N_3797,N_2497,N_2948);
and U3798 (N_3798,N_2064,N_2823);
or U3799 (N_3799,N_2157,N_2717);
nor U3800 (N_3800,N_2651,N_2889);
nor U3801 (N_3801,N_2372,N_2677);
nand U3802 (N_3802,N_2622,N_2420);
and U3803 (N_3803,N_2509,N_2275);
nor U3804 (N_3804,N_2732,N_2123);
nand U3805 (N_3805,N_2771,N_2749);
nor U3806 (N_3806,N_2688,N_2708);
nor U3807 (N_3807,N_2430,N_2909);
and U3808 (N_3808,N_2530,N_2086);
or U3809 (N_3809,N_2410,N_2426);
xor U3810 (N_3810,N_2361,N_2264);
nor U3811 (N_3811,N_2381,N_2935);
or U3812 (N_3812,N_2639,N_2432);
or U3813 (N_3813,N_2643,N_2364);
and U3814 (N_3814,N_2477,N_2024);
or U3815 (N_3815,N_2119,N_2437);
nor U3816 (N_3816,N_2919,N_2463);
and U3817 (N_3817,N_2389,N_2102);
and U3818 (N_3818,N_2755,N_2788);
nand U3819 (N_3819,N_2167,N_2683);
nand U3820 (N_3820,N_2392,N_2403);
or U3821 (N_3821,N_2833,N_2249);
and U3822 (N_3822,N_2830,N_2602);
nand U3823 (N_3823,N_2960,N_2513);
nor U3824 (N_3824,N_2651,N_2841);
nand U3825 (N_3825,N_2818,N_2557);
nand U3826 (N_3826,N_2742,N_2924);
or U3827 (N_3827,N_2607,N_2934);
nand U3828 (N_3828,N_2875,N_2194);
nor U3829 (N_3829,N_2627,N_2080);
or U3830 (N_3830,N_2680,N_2584);
nand U3831 (N_3831,N_2315,N_2918);
nor U3832 (N_3832,N_2646,N_2124);
nor U3833 (N_3833,N_2566,N_2541);
nor U3834 (N_3834,N_2980,N_2204);
nand U3835 (N_3835,N_2468,N_2774);
and U3836 (N_3836,N_2749,N_2533);
or U3837 (N_3837,N_2733,N_2689);
nand U3838 (N_3838,N_2915,N_2376);
nor U3839 (N_3839,N_2108,N_2187);
or U3840 (N_3840,N_2657,N_2785);
or U3841 (N_3841,N_2226,N_2360);
nand U3842 (N_3842,N_2009,N_2211);
nor U3843 (N_3843,N_2582,N_2577);
nand U3844 (N_3844,N_2666,N_2789);
nor U3845 (N_3845,N_2028,N_2579);
and U3846 (N_3846,N_2894,N_2525);
or U3847 (N_3847,N_2851,N_2957);
and U3848 (N_3848,N_2417,N_2995);
nor U3849 (N_3849,N_2360,N_2215);
nand U3850 (N_3850,N_2084,N_2977);
nor U3851 (N_3851,N_2800,N_2138);
nor U3852 (N_3852,N_2289,N_2165);
nand U3853 (N_3853,N_2645,N_2685);
nand U3854 (N_3854,N_2572,N_2934);
and U3855 (N_3855,N_2538,N_2727);
nand U3856 (N_3856,N_2000,N_2993);
and U3857 (N_3857,N_2138,N_2964);
nor U3858 (N_3858,N_2689,N_2053);
or U3859 (N_3859,N_2808,N_2339);
nand U3860 (N_3860,N_2050,N_2662);
or U3861 (N_3861,N_2437,N_2512);
nor U3862 (N_3862,N_2027,N_2061);
and U3863 (N_3863,N_2186,N_2107);
or U3864 (N_3864,N_2003,N_2449);
nor U3865 (N_3865,N_2323,N_2721);
and U3866 (N_3866,N_2545,N_2696);
or U3867 (N_3867,N_2013,N_2893);
nand U3868 (N_3868,N_2889,N_2276);
and U3869 (N_3869,N_2926,N_2635);
and U3870 (N_3870,N_2138,N_2938);
or U3871 (N_3871,N_2272,N_2688);
nor U3872 (N_3872,N_2785,N_2035);
nor U3873 (N_3873,N_2487,N_2738);
nor U3874 (N_3874,N_2475,N_2351);
and U3875 (N_3875,N_2310,N_2289);
nor U3876 (N_3876,N_2527,N_2991);
nand U3877 (N_3877,N_2942,N_2497);
or U3878 (N_3878,N_2241,N_2149);
or U3879 (N_3879,N_2167,N_2620);
or U3880 (N_3880,N_2607,N_2790);
and U3881 (N_3881,N_2581,N_2168);
nand U3882 (N_3882,N_2459,N_2947);
or U3883 (N_3883,N_2572,N_2329);
nand U3884 (N_3884,N_2744,N_2925);
nor U3885 (N_3885,N_2624,N_2359);
nand U3886 (N_3886,N_2034,N_2573);
or U3887 (N_3887,N_2400,N_2819);
nand U3888 (N_3888,N_2108,N_2379);
and U3889 (N_3889,N_2522,N_2745);
nand U3890 (N_3890,N_2775,N_2351);
or U3891 (N_3891,N_2729,N_2110);
xnor U3892 (N_3892,N_2497,N_2388);
nor U3893 (N_3893,N_2713,N_2419);
nor U3894 (N_3894,N_2994,N_2514);
or U3895 (N_3895,N_2380,N_2329);
and U3896 (N_3896,N_2026,N_2280);
or U3897 (N_3897,N_2468,N_2286);
nand U3898 (N_3898,N_2265,N_2870);
and U3899 (N_3899,N_2803,N_2795);
and U3900 (N_3900,N_2963,N_2904);
and U3901 (N_3901,N_2670,N_2582);
and U3902 (N_3902,N_2826,N_2884);
or U3903 (N_3903,N_2940,N_2376);
and U3904 (N_3904,N_2457,N_2307);
nor U3905 (N_3905,N_2686,N_2877);
and U3906 (N_3906,N_2138,N_2394);
nand U3907 (N_3907,N_2282,N_2366);
and U3908 (N_3908,N_2398,N_2873);
nor U3909 (N_3909,N_2876,N_2371);
nor U3910 (N_3910,N_2992,N_2169);
nor U3911 (N_3911,N_2191,N_2903);
or U3912 (N_3912,N_2681,N_2778);
xnor U3913 (N_3913,N_2593,N_2351);
nor U3914 (N_3914,N_2193,N_2677);
nand U3915 (N_3915,N_2252,N_2387);
and U3916 (N_3916,N_2264,N_2166);
or U3917 (N_3917,N_2204,N_2426);
or U3918 (N_3918,N_2548,N_2858);
nor U3919 (N_3919,N_2235,N_2975);
or U3920 (N_3920,N_2944,N_2424);
nor U3921 (N_3921,N_2443,N_2160);
nor U3922 (N_3922,N_2180,N_2697);
nor U3923 (N_3923,N_2581,N_2513);
nand U3924 (N_3924,N_2172,N_2061);
and U3925 (N_3925,N_2790,N_2366);
nor U3926 (N_3926,N_2794,N_2108);
xnor U3927 (N_3927,N_2833,N_2611);
and U3928 (N_3928,N_2953,N_2161);
nand U3929 (N_3929,N_2604,N_2317);
or U3930 (N_3930,N_2041,N_2373);
nor U3931 (N_3931,N_2500,N_2787);
nand U3932 (N_3932,N_2277,N_2624);
nand U3933 (N_3933,N_2747,N_2654);
nand U3934 (N_3934,N_2708,N_2529);
or U3935 (N_3935,N_2724,N_2662);
and U3936 (N_3936,N_2087,N_2612);
or U3937 (N_3937,N_2367,N_2858);
nor U3938 (N_3938,N_2323,N_2189);
nor U3939 (N_3939,N_2238,N_2470);
and U3940 (N_3940,N_2024,N_2612);
nand U3941 (N_3941,N_2218,N_2126);
and U3942 (N_3942,N_2424,N_2069);
and U3943 (N_3943,N_2236,N_2338);
or U3944 (N_3944,N_2376,N_2502);
or U3945 (N_3945,N_2931,N_2345);
nand U3946 (N_3946,N_2936,N_2443);
or U3947 (N_3947,N_2201,N_2019);
nor U3948 (N_3948,N_2699,N_2833);
nand U3949 (N_3949,N_2948,N_2671);
and U3950 (N_3950,N_2726,N_2173);
nor U3951 (N_3951,N_2883,N_2098);
nor U3952 (N_3952,N_2378,N_2969);
or U3953 (N_3953,N_2090,N_2395);
or U3954 (N_3954,N_2169,N_2544);
or U3955 (N_3955,N_2213,N_2703);
and U3956 (N_3956,N_2420,N_2115);
nor U3957 (N_3957,N_2820,N_2367);
and U3958 (N_3958,N_2895,N_2168);
nor U3959 (N_3959,N_2260,N_2700);
nor U3960 (N_3960,N_2033,N_2107);
or U3961 (N_3961,N_2709,N_2391);
or U3962 (N_3962,N_2523,N_2836);
nor U3963 (N_3963,N_2771,N_2878);
or U3964 (N_3964,N_2994,N_2490);
and U3965 (N_3965,N_2588,N_2649);
nand U3966 (N_3966,N_2928,N_2001);
nand U3967 (N_3967,N_2114,N_2698);
and U3968 (N_3968,N_2592,N_2257);
nand U3969 (N_3969,N_2100,N_2469);
and U3970 (N_3970,N_2080,N_2106);
or U3971 (N_3971,N_2528,N_2259);
and U3972 (N_3972,N_2775,N_2813);
or U3973 (N_3973,N_2898,N_2881);
and U3974 (N_3974,N_2525,N_2344);
nand U3975 (N_3975,N_2986,N_2881);
and U3976 (N_3976,N_2384,N_2937);
and U3977 (N_3977,N_2745,N_2550);
and U3978 (N_3978,N_2593,N_2250);
or U3979 (N_3979,N_2721,N_2135);
nand U3980 (N_3980,N_2732,N_2922);
nor U3981 (N_3981,N_2514,N_2374);
or U3982 (N_3982,N_2710,N_2933);
and U3983 (N_3983,N_2443,N_2184);
nand U3984 (N_3984,N_2967,N_2813);
nor U3985 (N_3985,N_2064,N_2303);
or U3986 (N_3986,N_2415,N_2348);
nor U3987 (N_3987,N_2150,N_2483);
or U3988 (N_3988,N_2265,N_2362);
nor U3989 (N_3989,N_2312,N_2714);
or U3990 (N_3990,N_2316,N_2775);
nand U3991 (N_3991,N_2638,N_2114);
and U3992 (N_3992,N_2913,N_2571);
nor U3993 (N_3993,N_2430,N_2441);
or U3994 (N_3994,N_2769,N_2737);
and U3995 (N_3995,N_2679,N_2032);
or U3996 (N_3996,N_2442,N_2907);
or U3997 (N_3997,N_2882,N_2492);
nor U3998 (N_3998,N_2703,N_2781);
or U3999 (N_3999,N_2981,N_2756);
nor U4000 (N_4000,N_3300,N_3895);
nor U4001 (N_4001,N_3033,N_3835);
nand U4002 (N_4002,N_3212,N_3047);
or U4003 (N_4003,N_3875,N_3170);
xor U4004 (N_4004,N_3705,N_3818);
or U4005 (N_4005,N_3506,N_3099);
or U4006 (N_4006,N_3790,N_3620);
nor U4007 (N_4007,N_3772,N_3696);
nand U4008 (N_4008,N_3554,N_3352);
and U4009 (N_4009,N_3124,N_3956);
or U4010 (N_4010,N_3019,N_3912);
or U4011 (N_4011,N_3330,N_3163);
nand U4012 (N_4012,N_3510,N_3748);
and U4013 (N_4013,N_3396,N_3842);
and U4014 (N_4014,N_3967,N_3279);
or U4015 (N_4015,N_3935,N_3563);
and U4016 (N_4016,N_3976,N_3478);
nor U4017 (N_4017,N_3295,N_3940);
nand U4018 (N_4018,N_3246,N_3836);
nor U4019 (N_4019,N_3437,N_3118);
and U4020 (N_4020,N_3307,N_3407);
and U4021 (N_4021,N_3885,N_3222);
or U4022 (N_4022,N_3401,N_3302);
nor U4023 (N_4023,N_3397,N_3176);
nand U4024 (N_4024,N_3160,N_3077);
nand U4025 (N_4025,N_3061,N_3725);
and U4026 (N_4026,N_3674,N_3685);
and U4027 (N_4027,N_3410,N_3614);
nand U4028 (N_4028,N_3777,N_3482);
nand U4029 (N_4029,N_3970,N_3656);
nand U4030 (N_4030,N_3794,N_3332);
and U4031 (N_4031,N_3497,N_3792);
and U4032 (N_4032,N_3427,N_3783);
nor U4033 (N_4033,N_3334,N_3228);
nand U4034 (N_4034,N_3826,N_3162);
nor U4035 (N_4035,N_3564,N_3067);
or U4036 (N_4036,N_3272,N_3593);
nor U4037 (N_4037,N_3089,N_3120);
nand U4038 (N_4038,N_3440,N_3242);
nand U4039 (N_4039,N_3567,N_3652);
and U4040 (N_4040,N_3240,N_3661);
or U4041 (N_4041,N_3984,N_3207);
and U4042 (N_4042,N_3843,N_3608);
nor U4043 (N_4043,N_3541,N_3785);
or U4044 (N_4044,N_3886,N_3384);
nor U4045 (N_4045,N_3631,N_3179);
nand U4046 (N_4046,N_3721,N_3997);
or U4047 (N_4047,N_3199,N_3399);
or U4048 (N_4048,N_3788,N_3423);
and U4049 (N_4049,N_3736,N_3626);
nor U4050 (N_4050,N_3690,N_3741);
nand U4051 (N_4051,N_3110,N_3058);
nor U4052 (N_4052,N_3202,N_3994);
and U4053 (N_4053,N_3130,N_3582);
nor U4054 (N_4054,N_3195,N_3264);
and U4055 (N_4055,N_3566,N_3119);
nor U4056 (N_4056,N_3784,N_3000);
nor U4057 (N_4057,N_3171,N_3481);
or U4058 (N_4058,N_3244,N_3548);
and U4059 (N_4059,N_3284,N_3519);
nand U4060 (N_4060,N_3451,N_3596);
or U4061 (N_4061,N_3923,N_3346);
xnor U4062 (N_4062,N_3680,N_3666);
nor U4063 (N_4063,N_3357,N_3245);
nand U4064 (N_4064,N_3867,N_3525);
nor U4065 (N_4065,N_3756,N_3765);
or U4066 (N_4066,N_3734,N_3194);
nor U4067 (N_4067,N_3601,N_3393);
nor U4068 (N_4068,N_3846,N_3745);
nand U4069 (N_4069,N_3914,N_3776);
or U4070 (N_4070,N_3031,N_3670);
nor U4071 (N_4071,N_3965,N_3884);
and U4072 (N_4072,N_3688,N_3964);
and U4073 (N_4073,N_3356,N_3209);
and U4074 (N_4074,N_3966,N_3263);
and U4075 (N_4075,N_3100,N_3092);
nor U4076 (N_4076,N_3659,N_3646);
nor U4077 (N_4077,N_3801,N_3649);
nand U4078 (N_4078,N_3679,N_3798);
nand U4079 (N_4079,N_3412,N_3834);
and U4080 (N_4080,N_3502,N_3498);
or U4081 (N_4081,N_3852,N_3625);
and U4082 (N_4082,N_3739,N_3390);
nand U4083 (N_4083,N_3709,N_3858);
nor U4084 (N_4084,N_3671,N_3839);
or U4085 (N_4085,N_3675,N_3483);
or U4086 (N_4086,N_3268,N_3728);
nor U4087 (N_4087,N_3349,N_3773);
and U4088 (N_4088,N_3471,N_3667);
nand U4089 (N_4089,N_3365,N_3004);
or U4090 (N_4090,N_3897,N_3056);
and U4091 (N_4091,N_3030,N_3971);
nand U4092 (N_4092,N_3862,N_3612);
nand U4093 (N_4093,N_3947,N_3111);
and U4094 (N_4094,N_3753,N_3229);
nor U4095 (N_4095,N_3309,N_3445);
nor U4096 (N_4096,N_3304,N_3337);
nand U4097 (N_4097,N_3648,N_3761);
nor U4098 (N_4098,N_3426,N_3917);
nor U4099 (N_4099,N_3184,N_3723);
nor U4100 (N_4100,N_3764,N_3115);
and U4101 (N_4101,N_3770,N_3466);
nor U4102 (N_4102,N_3308,N_3186);
nand U4103 (N_4103,N_3879,N_3489);
nor U4104 (N_4104,N_3559,N_3145);
nand U4105 (N_4105,N_3320,N_3683);
and U4106 (N_4106,N_3987,N_3359);
and U4107 (N_4107,N_3012,N_3522);
or U4108 (N_4108,N_3322,N_3116);
nor U4109 (N_4109,N_3579,N_3493);
or U4110 (N_4110,N_3720,N_3021);
and U4111 (N_4111,N_3958,N_3135);
nor U4112 (N_4112,N_3805,N_3573);
and U4113 (N_4113,N_3899,N_3848);
or U4114 (N_4114,N_3473,N_3036);
nand U4115 (N_4115,N_3691,N_3260);
and U4116 (N_4116,N_3639,N_3323);
or U4117 (N_4117,N_3221,N_3664);
and U4118 (N_4118,N_3180,N_3206);
or U4119 (N_4119,N_3220,N_3062);
or U4120 (N_4120,N_3715,N_3536);
or U4121 (N_4121,N_3429,N_3371);
and U4122 (N_4122,N_3153,N_3029);
and U4123 (N_4123,N_3598,N_3041);
and U4124 (N_4124,N_3859,N_3324);
and U4125 (N_4125,N_3504,N_3619);
nand U4126 (N_4126,N_3795,N_3386);
nand U4127 (N_4127,N_3225,N_3565);
nor U4128 (N_4128,N_3192,N_3046);
or U4129 (N_4129,N_3475,N_3490);
nand U4130 (N_4130,N_3044,N_3640);
and U4131 (N_4131,N_3239,N_3543);
nor U4132 (N_4132,N_3876,N_3389);
and U4133 (N_4133,N_3151,N_3621);
nand U4134 (N_4134,N_3992,N_3286);
nor U4135 (N_4135,N_3941,N_3024);
nor U4136 (N_4136,N_3079,N_3779);
nand U4137 (N_4137,N_3963,N_3382);
nand U4138 (N_4138,N_3109,N_3530);
or U4139 (N_4139,N_3526,N_3901);
nor U4140 (N_4140,N_3296,N_3955);
nor U4141 (N_4141,N_3204,N_3518);
or U4142 (N_4142,N_3547,N_3977);
nand U4143 (N_4143,N_3040,N_3444);
nor U4144 (N_4144,N_3350,N_3432);
nand U4145 (N_4145,N_3319,N_3500);
or U4146 (N_4146,N_3453,N_3443);
and U4147 (N_4147,N_3628,N_3032);
nor U4148 (N_4148,N_3629,N_3896);
or U4149 (N_4149,N_3752,N_3123);
or U4150 (N_4150,N_3231,N_3226);
nor U4151 (N_4151,N_3161,N_3982);
nand U4152 (N_4152,N_3342,N_3078);
or U4153 (N_4153,N_3340,N_3817);
nor U4154 (N_4154,N_3767,N_3751);
nor U4155 (N_4155,N_3939,N_3368);
and U4156 (N_4156,N_3754,N_3749);
nor U4157 (N_4157,N_3157,N_3201);
nor U4158 (N_4158,N_3552,N_3665);
or U4159 (N_4159,N_3477,N_3121);
or U4160 (N_4160,N_3253,N_3146);
nand U4161 (N_4161,N_3789,N_3558);
or U4162 (N_4162,N_3388,N_3918);
or U4163 (N_4163,N_3400,N_3837);
and U4164 (N_4164,N_3583,N_3920);
and U4165 (N_4165,N_3529,N_3358);
nor U4166 (N_4166,N_3177,N_3537);
nor U4167 (N_4167,N_3611,N_3132);
nand U4168 (N_4168,N_3376,N_3452);
nand U4169 (N_4169,N_3066,N_3211);
and U4170 (N_4170,N_3002,N_3610);
or U4171 (N_4171,N_3823,N_3763);
or U4172 (N_4172,N_3880,N_3695);
and U4173 (N_4173,N_3613,N_3703);
nor U4174 (N_4174,N_3043,N_3136);
and U4175 (N_4175,N_3250,N_3542);
nor U4176 (N_4176,N_3081,N_3624);
and U4177 (N_4177,N_3810,N_3915);
nor U4178 (N_4178,N_3891,N_3187);
nand U4179 (N_4179,N_3329,N_3294);
or U4180 (N_4180,N_3570,N_3678);
nor U4181 (N_4181,N_3127,N_3603);
and U4182 (N_4182,N_3085,N_3236);
nor U4183 (N_4183,N_3314,N_3926);
nand U4184 (N_4184,N_3869,N_3532);
or U4185 (N_4185,N_3080,N_3589);
or U4186 (N_4186,N_3375,N_3045);
nand U4187 (N_4187,N_3280,N_3871);
or U4188 (N_4188,N_3414,N_3856);
or U4189 (N_4189,N_3945,N_3605);
or U4190 (N_4190,N_3636,N_3496);
or U4191 (N_4191,N_3105,N_3057);
nor U4192 (N_4192,N_3909,N_3405);
or U4193 (N_4193,N_3241,N_3052);
nand U4194 (N_4194,N_3069,N_3213);
or U4195 (N_4195,N_3824,N_3572);
and U4196 (N_4196,N_3035,N_3508);
or U4197 (N_4197,N_3011,N_3476);
nand U4198 (N_4198,N_3507,N_3232);
or U4199 (N_4199,N_3616,N_3948);
and U4200 (N_4200,N_3474,N_3906);
or U4201 (N_4201,N_3927,N_3463);
and U4202 (N_4202,N_3327,N_3025);
or U4203 (N_4203,N_3944,N_3172);
or U4204 (N_4204,N_3139,N_3424);
nor U4205 (N_4205,N_3505,N_3953);
and U4206 (N_4206,N_3581,N_3464);
nand U4207 (N_4207,N_3857,N_3088);
or U4208 (N_4208,N_3697,N_3439);
nand U4209 (N_4209,N_3459,N_3988);
nor U4210 (N_4210,N_3487,N_3039);
or U4211 (N_4211,N_3372,N_3845);
or U4212 (N_4212,N_3328,N_3149);
and U4213 (N_4213,N_3738,N_3617);
or U4214 (N_4214,N_3255,N_3718);
and U4215 (N_4215,N_3578,N_3273);
nor U4216 (N_4216,N_3657,N_3167);
and U4217 (N_4217,N_3627,N_3347);
nor U4218 (N_4218,N_3183,N_3339);
nor U4219 (N_4219,N_3299,N_3442);
nor U4220 (N_4220,N_3706,N_3872);
or U4221 (N_4221,N_3355,N_3458);
nand U4222 (N_4222,N_3422,N_3398);
and U4223 (N_4223,N_3998,N_3793);
or U4224 (N_4224,N_3147,N_3456);
nand U4225 (N_4225,N_3495,N_3306);
and U4226 (N_4226,N_3995,N_3866);
or U4227 (N_4227,N_3851,N_3083);
nor U4228 (N_4228,N_3148,N_3647);
and U4229 (N_4229,N_3301,N_3419);
or U4230 (N_4230,N_3873,N_3402);
or U4231 (N_4231,N_3711,N_3017);
or U4232 (N_4232,N_3185,N_3038);
and U4233 (N_4233,N_3902,N_3545);
nand U4234 (N_4234,N_3234,N_3802);
and U4235 (N_4235,N_3274,N_3870);
nand U4236 (N_4236,N_3618,N_3553);
or U4237 (N_4237,N_3560,N_3946);
nand U4238 (N_4238,N_3716,N_3978);
nand U4239 (N_4239,N_3684,N_3363);
nor U4240 (N_4240,N_3005,N_3406);
and U4241 (N_4241,N_3297,N_3847);
nor U4242 (N_4242,N_3114,N_3433);
and U4243 (N_4243,N_3203,N_3527);
or U4244 (N_4244,N_3403,N_3724);
and U4245 (N_4245,N_3571,N_3925);
nor U4246 (N_4246,N_3592,N_3107);
and U4247 (N_4247,N_3520,N_3181);
nand U4248 (N_4248,N_3740,N_3415);
nand U4249 (N_4249,N_3072,N_3993);
and U4250 (N_4250,N_3141,N_3877);
or U4251 (N_4251,N_3860,N_3854);
or U4252 (N_4252,N_3015,N_3849);
nor U4253 (N_4253,N_3972,N_3492);
nand U4254 (N_4254,N_3594,N_3395);
or U4255 (N_4255,N_3050,N_3354);
nand U4256 (N_4256,N_3026,N_3929);
and U4257 (N_4257,N_3137,N_3694);
or U4258 (N_4258,N_3832,N_3315);
or U4259 (N_4259,N_3800,N_3009);
or U4260 (N_4260,N_3076,N_3208);
and U4261 (N_4261,N_3808,N_3991);
xor U4262 (N_4262,N_3874,N_3028);
nand U4263 (N_4263,N_3367,N_3533);
nor U4264 (N_4264,N_3523,N_3103);
nand U4265 (N_4265,N_3434,N_3408);
nand U4266 (N_4266,N_3546,N_3362);
or U4267 (N_4267,N_3643,N_3766);
or U4268 (N_4268,N_3430,N_3774);
or U4269 (N_4269,N_3462,N_3893);
or U4270 (N_4270,N_3681,N_3797);
nor U4271 (N_4271,N_3075,N_3758);
or U4272 (N_4272,N_3922,N_3868);
or U4273 (N_4273,N_3677,N_3494);
nand U4274 (N_4274,N_3164,N_3635);
and U4275 (N_4275,N_3325,N_3786);
nor U4276 (N_4276,N_3934,N_3373);
or U4277 (N_4277,N_3864,N_3919);
and U4278 (N_4278,N_3383,N_3775);
and U4279 (N_4279,N_3737,N_3534);
or U4280 (N_4280,N_3961,N_3449);
or U4281 (N_4281,N_3150,N_3949);
and U4282 (N_4282,N_3238,N_3070);
and U4283 (N_4283,N_3305,N_3557);
nand U4284 (N_4284,N_3097,N_3930);
and U4285 (N_4285,N_3954,N_3133);
or U4286 (N_4286,N_3182,N_3606);
or U4287 (N_4287,N_3053,N_3962);
nor U4288 (N_4288,N_3531,N_3831);
nand U4289 (N_4289,N_3421,N_3913);
nor U4290 (N_4290,N_3457,N_3812);
and U4291 (N_4291,N_3054,N_3479);
nand U4292 (N_4292,N_3803,N_3676);
and U4293 (N_4293,N_3780,N_3750);
or U4294 (N_4294,N_3227,N_3517);
or U4295 (N_4295,N_3193,N_3265);
nor U4296 (N_4296,N_3951,N_3385);
or U4297 (N_4297,N_3568,N_3413);
nor U4298 (N_4298,N_3701,N_3189);
nor U4299 (N_4299,N_3576,N_3205);
xnor U4300 (N_4300,N_3950,N_3387);
and U4301 (N_4301,N_3258,N_3735);
nand U4302 (N_4302,N_3924,N_3822);
nand U4303 (N_4303,N_3460,N_3825);
and U4304 (N_4304,N_3173,N_3472);
and U4305 (N_4305,N_3027,N_3607);
nand U4306 (N_4306,N_3312,N_3259);
and U4307 (N_4307,N_3113,N_3760);
nand U4308 (N_4308,N_3428,N_3574);
nor U4309 (N_4309,N_3049,N_3855);
and U4310 (N_4310,N_3288,N_3343);
nor U4311 (N_4311,N_3480,N_3898);
nor U4312 (N_4312,N_3404,N_3344);
nor U4313 (N_4313,N_3037,N_3071);
or U4314 (N_4314,N_3001,N_3013);
nand U4315 (N_4315,N_3290,N_3746);
nor U4316 (N_4316,N_3095,N_3065);
nor U4317 (N_4317,N_3051,N_3807);
nand U4318 (N_4318,N_3455,N_3336);
nor U4319 (N_4319,N_3910,N_3602);
or U4320 (N_4320,N_3615,N_3318);
or U4321 (N_4321,N_3544,N_3285);
or U4322 (N_4322,N_3023,N_3599);
nand U4323 (N_4323,N_3178,N_3267);
nand U4324 (N_4324,N_3747,N_3587);
nand U4325 (N_4325,N_3214,N_3699);
and U4326 (N_4326,N_3197,N_3816);
and U4327 (N_4327,N_3999,N_3277);
nor U4328 (N_4328,N_3710,N_3377);
nand U4329 (N_4329,N_3435,N_3811);
or U4330 (N_4330,N_3952,N_3905);
nand U4331 (N_4331,N_3689,N_3708);
and U4332 (N_4332,N_3064,N_3799);
nor U4333 (N_4333,N_3217,N_3317);
nor U4334 (N_4334,N_3216,N_3486);
xor U4335 (N_4335,N_3727,N_3804);
or U4336 (N_4336,N_3539,N_3755);
nor U4337 (N_4337,N_3392,N_3303);
nand U4338 (N_4338,N_3907,N_3074);
or U4339 (N_4339,N_3438,N_3983);
nor U4340 (N_4340,N_3082,N_3682);
and U4341 (N_4341,N_3158,N_3420);
nand U4342 (N_4342,N_3714,N_3391);
or U4343 (N_4343,N_3622,N_3048);
and U4344 (N_4344,N_3278,N_3073);
nor U4345 (N_4345,N_3597,N_3704);
and U4346 (N_4346,N_3742,N_3590);
nor U4347 (N_4347,N_3448,N_3447);
and U4348 (N_4348,N_3292,N_3861);
nand U4349 (N_4349,N_3333,N_3271);
or U4350 (N_4350,N_3353,N_3693);
nand U4351 (N_4351,N_3112,N_3159);
and U4352 (N_4352,N_3129,N_3436);
nand U4353 (N_4353,N_3781,N_3974);
and U4354 (N_4354,N_3702,N_3722);
nand U4355 (N_4355,N_3577,N_3461);
nand U4356 (N_4356,N_3719,N_3882);
nand U4357 (N_4357,N_3311,N_3960);
nor U4358 (N_4358,N_3450,N_3936);
and U4359 (N_4359,N_3637,N_3819);
and U4360 (N_4360,N_3686,N_3561);
nor U4361 (N_4361,N_3655,N_3707);
nand U4362 (N_4362,N_3585,N_3374);
and U4363 (N_4363,N_3562,N_3446);
nand U4364 (N_4364,N_3890,N_3778);
or U4365 (N_4365,N_3806,N_3762);
and U4366 (N_4366,N_3730,N_3126);
and U4367 (N_4367,N_3521,N_3650);
and U4368 (N_4368,N_3516,N_3841);
nor U4369 (N_4369,N_3660,N_3465);
nand U4370 (N_4370,N_3068,N_3840);
nor U4371 (N_4371,N_3827,N_3535);
nand U4372 (N_4372,N_3441,N_3055);
nand U4373 (N_4373,N_3883,N_3633);
and U4374 (N_4374,N_3233,N_3022);
or U4375 (N_4375,N_3609,N_3512);
and U4376 (N_4376,N_3007,N_3484);
nand U4377 (N_4377,N_3369,N_3981);
nand U4378 (N_4378,N_3892,N_3975);
nor U4379 (N_4379,N_3980,N_3759);
nand U4380 (N_4380,N_3169,N_3266);
or U4381 (N_4381,N_3641,N_3200);
or U4382 (N_4382,N_3878,N_3379);
nand U4383 (N_4383,N_3468,N_3191);
nor U4384 (N_4384,N_3364,N_3488);
or U4385 (N_4385,N_3673,N_3509);
or U4386 (N_4386,N_3018,N_3293);
and U4387 (N_4387,N_3501,N_3888);
nor U4388 (N_4388,N_3887,N_3908);
nand U4389 (N_4389,N_3938,N_3165);
nor U4390 (N_4390,N_3782,N_3903);
nand U4391 (N_4391,N_3771,N_3224);
nor U4392 (N_4392,N_3351,N_3644);
and U4393 (N_4393,N_3973,N_3360);
and U4394 (N_4394,N_3128,N_3503);
and U4395 (N_4395,N_3152,N_3584);
and U4396 (N_4396,N_3672,N_3006);
or U4397 (N_4397,N_3555,N_3174);
nand U4398 (N_4398,N_3968,N_3580);
or U4399 (N_4399,N_3513,N_3916);
nor U4400 (N_4400,N_3485,N_3168);
nor U4401 (N_4401,N_3215,N_3687);
nand U4402 (N_4402,N_3247,N_3733);
and U4403 (N_4403,N_3251,N_3850);
nor U4404 (N_4404,N_3060,N_3904);
nand U4405 (N_4405,N_3932,N_3094);
nor U4406 (N_4406,N_3669,N_3863);
nand U4407 (N_4407,N_3630,N_3757);
and U4408 (N_4408,N_3198,N_3096);
nand U4409 (N_4409,N_3658,N_3090);
or U4410 (N_4410,N_3144,N_3087);
and U4411 (N_4411,N_3230,N_3218);
nor U4412 (N_4412,N_3237,N_3411);
nor U4413 (N_4413,N_3515,N_3287);
and U4414 (N_4414,N_3600,N_3042);
nand U4415 (N_4415,N_3166,N_3768);
or U4416 (N_4416,N_3814,N_3979);
and U4417 (N_4417,N_3829,N_3985);
and U4418 (N_4418,N_3809,N_3361);
xnor U4419 (N_4419,N_3623,N_3595);
or U4420 (N_4420,N_3791,N_3190);
nand U4421 (N_4421,N_3713,N_3154);
and U4422 (N_4422,N_3769,N_3138);
and U4423 (N_4423,N_3321,N_3270);
and U4424 (N_4424,N_3550,N_3499);
nand U4425 (N_4425,N_3010,N_3731);
or U4426 (N_4426,N_3059,N_3252);
and U4427 (N_4427,N_3249,N_3556);
nor U4428 (N_4428,N_3668,N_3175);
nand U4429 (N_4429,N_3140,N_3256);
or U4430 (N_4430,N_3491,N_3394);
nor U4431 (N_4431,N_3235,N_3634);
nand U4432 (N_4432,N_3524,N_3269);
nand U4433 (N_4433,N_3700,N_3853);
nor U4434 (N_4434,N_3335,N_3156);
xnor U4435 (N_4435,N_3514,N_3338);
nand U4436 (N_4436,N_3289,N_3131);
nor U4437 (N_4437,N_3538,N_3425);
or U4438 (N_4438,N_3881,N_3142);
xor U4439 (N_4439,N_3380,N_3418);
or U4440 (N_4440,N_3921,N_3416);
nand U4441 (N_4441,N_3986,N_3431);
and U4442 (N_4442,N_3223,N_3889);
and U4443 (N_4443,N_3063,N_3125);
nor U4444 (N_4444,N_3104,N_3101);
nand U4445 (N_4445,N_3108,N_3928);
or U4446 (N_4446,N_3370,N_3276);
nor U4447 (N_4447,N_3511,N_3102);
nand U4448 (N_4448,N_3830,N_3117);
and U4449 (N_4449,N_3787,N_3931);
and U4450 (N_4450,N_3942,N_3210);
nor U4451 (N_4451,N_3188,N_3698);
nor U4452 (N_4452,N_3865,N_3243);
and U4453 (N_4453,N_3016,N_3091);
or U4454 (N_4454,N_3743,N_3454);
or U4455 (N_4455,N_3262,N_3469);
or U4456 (N_4456,N_3959,N_3540);
or U4457 (N_4457,N_3020,N_3282);
or U4458 (N_4458,N_3575,N_3122);
or U4459 (N_4459,N_3933,N_3008);
nand U4460 (N_4460,N_3712,N_3143);
and U4461 (N_4461,N_3732,N_3381);
or U4462 (N_4462,N_3281,N_3313);
or U4463 (N_4463,N_3348,N_3894);
nand U4464 (N_4464,N_3591,N_3604);
nor U4465 (N_4465,N_3196,N_3833);
or U4466 (N_4466,N_3717,N_3989);
nand U4467 (N_4467,N_3417,N_3257);
nand U4468 (N_4468,N_3470,N_3937);
nand U4469 (N_4469,N_3326,N_3283);
and U4470 (N_4470,N_3549,N_3528);
and U4471 (N_4471,N_3331,N_3844);
nor U4472 (N_4472,N_3003,N_3645);
and U4473 (N_4473,N_3275,N_3796);
or U4474 (N_4474,N_3996,N_3651);
and U4475 (N_4475,N_3316,N_3990);
and U4476 (N_4476,N_3838,N_3345);
nand U4477 (N_4477,N_3957,N_3726);
or U4478 (N_4478,N_3943,N_3341);
or U4479 (N_4479,N_3744,N_3106);
nand U4480 (N_4480,N_3911,N_3084);
nor U4481 (N_4481,N_3663,N_3093);
and U4482 (N_4482,N_3310,N_3569);
or U4483 (N_4483,N_3261,N_3254);
and U4484 (N_4484,N_3821,N_3134);
nand U4485 (N_4485,N_3291,N_3588);
nand U4486 (N_4486,N_3662,N_3638);
and U4487 (N_4487,N_3366,N_3729);
nor U4488 (N_4488,N_3378,N_3900);
nand U4489 (N_4489,N_3632,N_3815);
and U4490 (N_4490,N_3820,N_3086);
nor U4491 (N_4491,N_3813,N_3692);
nor U4492 (N_4492,N_3642,N_3098);
and U4493 (N_4493,N_3219,N_3248);
or U4494 (N_4494,N_3298,N_3467);
and U4495 (N_4495,N_3654,N_3551);
and U4496 (N_4496,N_3014,N_3828);
nand U4497 (N_4497,N_3155,N_3653);
nand U4498 (N_4498,N_3409,N_3969);
nor U4499 (N_4499,N_3034,N_3586);
nand U4500 (N_4500,N_3342,N_3771);
nor U4501 (N_4501,N_3240,N_3794);
nand U4502 (N_4502,N_3767,N_3617);
nor U4503 (N_4503,N_3171,N_3797);
nor U4504 (N_4504,N_3658,N_3375);
nand U4505 (N_4505,N_3517,N_3923);
or U4506 (N_4506,N_3089,N_3602);
or U4507 (N_4507,N_3931,N_3261);
nor U4508 (N_4508,N_3677,N_3933);
and U4509 (N_4509,N_3937,N_3755);
or U4510 (N_4510,N_3835,N_3756);
nand U4511 (N_4511,N_3805,N_3918);
and U4512 (N_4512,N_3165,N_3360);
and U4513 (N_4513,N_3026,N_3148);
or U4514 (N_4514,N_3052,N_3783);
nand U4515 (N_4515,N_3861,N_3102);
nor U4516 (N_4516,N_3162,N_3974);
nor U4517 (N_4517,N_3157,N_3303);
or U4518 (N_4518,N_3683,N_3130);
or U4519 (N_4519,N_3720,N_3613);
nor U4520 (N_4520,N_3825,N_3676);
xor U4521 (N_4521,N_3526,N_3225);
nand U4522 (N_4522,N_3428,N_3852);
or U4523 (N_4523,N_3404,N_3252);
nand U4524 (N_4524,N_3776,N_3200);
or U4525 (N_4525,N_3437,N_3444);
and U4526 (N_4526,N_3842,N_3771);
and U4527 (N_4527,N_3746,N_3997);
or U4528 (N_4528,N_3709,N_3879);
or U4529 (N_4529,N_3722,N_3026);
nor U4530 (N_4530,N_3773,N_3581);
nand U4531 (N_4531,N_3884,N_3618);
and U4532 (N_4532,N_3491,N_3927);
nand U4533 (N_4533,N_3613,N_3890);
or U4534 (N_4534,N_3712,N_3285);
or U4535 (N_4535,N_3448,N_3675);
and U4536 (N_4536,N_3135,N_3992);
and U4537 (N_4537,N_3979,N_3362);
nor U4538 (N_4538,N_3650,N_3007);
nand U4539 (N_4539,N_3845,N_3947);
nor U4540 (N_4540,N_3672,N_3469);
nor U4541 (N_4541,N_3692,N_3340);
nand U4542 (N_4542,N_3467,N_3098);
nand U4543 (N_4543,N_3504,N_3163);
and U4544 (N_4544,N_3757,N_3579);
nor U4545 (N_4545,N_3377,N_3287);
nand U4546 (N_4546,N_3786,N_3795);
and U4547 (N_4547,N_3367,N_3390);
nor U4548 (N_4548,N_3951,N_3722);
and U4549 (N_4549,N_3977,N_3284);
and U4550 (N_4550,N_3672,N_3127);
or U4551 (N_4551,N_3436,N_3354);
xor U4552 (N_4552,N_3189,N_3654);
or U4553 (N_4553,N_3935,N_3881);
nand U4554 (N_4554,N_3932,N_3612);
nand U4555 (N_4555,N_3879,N_3200);
nand U4556 (N_4556,N_3091,N_3837);
or U4557 (N_4557,N_3689,N_3306);
nor U4558 (N_4558,N_3412,N_3117);
nor U4559 (N_4559,N_3493,N_3203);
or U4560 (N_4560,N_3493,N_3361);
nor U4561 (N_4561,N_3036,N_3864);
nor U4562 (N_4562,N_3411,N_3442);
or U4563 (N_4563,N_3741,N_3923);
and U4564 (N_4564,N_3195,N_3974);
nand U4565 (N_4565,N_3005,N_3583);
and U4566 (N_4566,N_3137,N_3644);
or U4567 (N_4567,N_3455,N_3168);
nor U4568 (N_4568,N_3690,N_3752);
nor U4569 (N_4569,N_3253,N_3438);
or U4570 (N_4570,N_3632,N_3017);
nor U4571 (N_4571,N_3162,N_3198);
and U4572 (N_4572,N_3033,N_3826);
and U4573 (N_4573,N_3511,N_3639);
or U4574 (N_4574,N_3042,N_3829);
nor U4575 (N_4575,N_3442,N_3425);
and U4576 (N_4576,N_3469,N_3762);
nor U4577 (N_4577,N_3556,N_3830);
nand U4578 (N_4578,N_3488,N_3321);
and U4579 (N_4579,N_3384,N_3905);
and U4580 (N_4580,N_3655,N_3229);
and U4581 (N_4581,N_3911,N_3377);
nand U4582 (N_4582,N_3306,N_3519);
or U4583 (N_4583,N_3814,N_3001);
or U4584 (N_4584,N_3828,N_3188);
or U4585 (N_4585,N_3375,N_3640);
or U4586 (N_4586,N_3140,N_3787);
and U4587 (N_4587,N_3223,N_3510);
nor U4588 (N_4588,N_3017,N_3205);
and U4589 (N_4589,N_3602,N_3395);
nand U4590 (N_4590,N_3188,N_3246);
and U4591 (N_4591,N_3502,N_3555);
nor U4592 (N_4592,N_3887,N_3676);
and U4593 (N_4593,N_3101,N_3366);
nand U4594 (N_4594,N_3666,N_3312);
or U4595 (N_4595,N_3057,N_3485);
nor U4596 (N_4596,N_3199,N_3987);
nor U4597 (N_4597,N_3927,N_3966);
or U4598 (N_4598,N_3800,N_3525);
and U4599 (N_4599,N_3799,N_3056);
nand U4600 (N_4600,N_3514,N_3043);
nand U4601 (N_4601,N_3329,N_3914);
and U4602 (N_4602,N_3668,N_3511);
nor U4603 (N_4603,N_3903,N_3401);
nand U4604 (N_4604,N_3806,N_3460);
nand U4605 (N_4605,N_3625,N_3472);
nor U4606 (N_4606,N_3773,N_3425);
and U4607 (N_4607,N_3956,N_3830);
and U4608 (N_4608,N_3135,N_3166);
nand U4609 (N_4609,N_3741,N_3065);
and U4610 (N_4610,N_3556,N_3248);
and U4611 (N_4611,N_3597,N_3451);
or U4612 (N_4612,N_3252,N_3226);
nor U4613 (N_4613,N_3056,N_3177);
and U4614 (N_4614,N_3543,N_3706);
nand U4615 (N_4615,N_3906,N_3020);
or U4616 (N_4616,N_3908,N_3464);
nand U4617 (N_4617,N_3159,N_3792);
or U4618 (N_4618,N_3524,N_3115);
or U4619 (N_4619,N_3188,N_3029);
nor U4620 (N_4620,N_3529,N_3845);
or U4621 (N_4621,N_3201,N_3143);
nor U4622 (N_4622,N_3688,N_3980);
and U4623 (N_4623,N_3267,N_3659);
nor U4624 (N_4624,N_3401,N_3609);
nor U4625 (N_4625,N_3705,N_3838);
nand U4626 (N_4626,N_3422,N_3574);
and U4627 (N_4627,N_3862,N_3195);
nor U4628 (N_4628,N_3178,N_3800);
nor U4629 (N_4629,N_3075,N_3080);
and U4630 (N_4630,N_3065,N_3094);
nand U4631 (N_4631,N_3722,N_3052);
nor U4632 (N_4632,N_3920,N_3447);
and U4633 (N_4633,N_3263,N_3862);
nor U4634 (N_4634,N_3821,N_3865);
nor U4635 (N_4635,N_3468,N_3483);
nand U4636 (N_4636,N_3355,N_3228);
and U4637 (N_4637,N_3257,N_3632);
xor U4638 (N_4638,N_3618,N_3685);
and U4639 (N_4639,N_3400,N_3614);
nor U4640 (N_4640,N_3117,N_3500);
or U4641 (N_4641,N_3385,N_3443);
and U4642 (N_4642,N_3507,N_3513);
or U4643 (N_4643,N_3797,N_3517);
and U4644 (N_4644,N_3133,N_3789);
and U4645 (N_4645,N_3762,N_3865);
nor U4646 (N_4646,N_3110,N_3088);
or U4647 (N_4647,N_3454,N_3531);
nand U4648 (N_4648,N_3794,N_3592);
or U4649 (N_4649,N_3773,N_3597);
and U4650 (N_4650,N_3775,N_3927);
nand U4651 (N_4651,N_3040,N_3507);
nor U4652 (N_4652,N_3174,N_3129);
or U4653 (N_4653,N_3147,N_3536);
nor U4654 (N_4654,N_3703,N_3596);
nor U4655 (N_4655,N_3862,N_3184);
and U4656 (N_4656,N_3155,N_3638);
or U4657 (N_4657,N_3601,N_3961);
and U4658 (N_4658,N_3957,N_3570);
and U4659 (N_4659,N_3896,N_3153);
and U4660 (N_4660,N_3321,N_3936);
or U4661 (N_4661,N_3563,N_3314);
or U4662 (N_4662,N_3327,N_3295);
xor U4663 (N_4663,N_3887,N_3229);
and U4664 (N_4664,N_3446,N_3841);
or U4665 (N_4665,N_3507,N_3757);
and U4666 (N_4666,N_3097,N_3894);
nand U4667 (N_4667,N_3916,N_3674);
or U4668 (N_4668,N_3707,N_3307);
or U4669 (N_4669,N_3478,N_3780);
or U4670 (N_4670,N_3954,N_3758);
and U4671 (N_4671,N_3509,N_3607);
and U4672 (N_4672,N_3845,N_3652);
nand U4673 (N_4673,N_3719,N_3794);
or U4674 (N_4674,N_3944,N_3064);
and U4675 (N_4675,N_3457,N_3950);
and U4676 (N_4676,N_3224,N_3117);
and U4677 (N_4677,N_3130,N_3613);
and U4678 (N_4678,N_3776,N_3423);
or U4679 (N_4679,N_3681,N_3942);
nand U4680 (N_4680,N_3512,N_3030);
nor U4681 (N_4681,N_3903,N_3136);
or U4682 (N_4682,N_3810,N_3359);
nor U4683 (N_4683,N_3927,N_3465);
nor U4684 (N_4684,N_3517,N_3165);
or U4685 (N_4685,N_3388,N_3545);
nor U4686 (N_4686,N_3255,N_3041);
or U4687 (N_4687,N_3851,N_3505);
and U4688 (N_4688,N_3177,N_3046);
and U4689 (N_4689,N_3705,N_3777);
nand U4690 (N_4690,N_3896,N_3370);
nand U4691 (N_4691,N_3866,N_3377);
nand U4692 (N_4692,N_3072,N_3699);
or U4693 (N_4693,N_3318,N_3473);
nand U4694 (N_4694,N_3045,N_3232);
nor U4695 (N_4695,N_3217,N_3965);
and U4696 (N_4696,N_3041,N_3525);
and U4697 (N_4697,N_3156,N_3601);
and U4698 (N_4698,N_3751,N_3907);
nor U4699 (N_4699,N_3284,N_3130);
nor U4700 (N_4700,N_3317,N_3046);
nand U4701 (N_4701,N_3752,N_3527);
nor U4702 (N_4702,N_3876,N_3871);
nand U4703 (N_4703,N_3318,N_3820);
nor U4704 (N_4704,N_3867,N_3037);
nor U4705 (N_4705,N_3431,N_3599);
or U4706 (N_4706,N_3416,N_3494);
nor U4707 (N_4707,N_3838,N_3435);
or U4708 (N_4708,N_3717,N_3943);
or U4709 (N_4709,N_3591,N_3123);
or U4710 (N_4710,N_3533,N_3553);
or U4711 (N_4711,N_3752,N_3145);
and U4712 (N_4712,N_3448,N_3551);
and U4713 (N_4713,N_3904,N_3480);
nand U4714 (N_4714,N_3181,N_3233);
and U4715 (N_4715,N_3232,N_3734);
nand U4716 (N_4716,N_3438,N_3395);
or U4717 (N_4717,N_3576,N_3466);
nand U4718 (N_4718,N_3036,N_3108);
nand U4719 (N_4719,N_3681,N_3277);
or U4720 (N_4720,N_3738,N_3234);
or U4721 (N_4721,N_3549,N_3349);
nand U4722 (N_4722,N_3062,N_3829);
and U4723 (N_4723,N_3063,N_3526);
or U4724 (N_4724,N_3977,N_3688);
and U4725 (N_4725,N_3587,N_3529);
and U4726 (N_4726,N_3995,N_3288);
nand U4727 (N_4727,N_3665,N_3565);
or U4728 (N_4728,N_3209,N_3883);
and U4729 (N_4729,N_3517,N_3794);
nand U4730 (N_4730,N_3324,N_3466);
nand U4731 (N_4731,N_3679,N_3599);
or U4732 (N_4732,N_3044,N_3749);
nor U4733 (N_4733,N_3476,N_3192);
or U4734 (N_4734,N_3122,N_3963);
or U4735 (N_4735,N_3531,N_3824);
and U4736 (N_4736,N_3973,N_3536);
and U4737 (N_4737,N_3424,N_3482);
nand U4738 (N_4738,N_3237,N_3620);
nand U4739 (N_4739,N_3348,N_3286);
nor U4740 (N_4740,N_3390,N_3240);
or U4741 (N_4741,N_3580,N_3053);
or U4742 (N_4742,N_3050,N_3984);
or U4743 (N_4743,N_3890,N_3117);
nor U4744 (N_4744,N_3213,N_3251);
or U4745 (N_4745,N_3564,N_3144);
and U4746 (N_4746,N_3766,N_3022);
or U4747 (N_4747,N_3109,N_3311);
nand U4748 (N_4748,N_3662,N_3944);
xor U4749 (N_4749,N_3334,N_3806);
nand U4750 (N_4750,N_3830,N_3060);
nor U4751 (N_4751,N_3510,N_3841);
or U4752 (N_4752,N_3794,N_3929);
or U4753 (N_4753,N_3874,N_3470);
nand U4754 (N_4754,N_3180,N_3123);
nand U4755 (N_4755,N_3378,N_3442);
or U4756 (N_4756,N_3100,N_3342);
or U4757 (N_4757,N_3492,N_3176);
or U4758 (N_4758,N_3650,N_3568);
or U4759 (N_4759,N_3037,N_3389);
and U4760 (N_4760,N_3725,N_3649);
nand U4761 (N_4761,N_3109,N_3965);
and U4762 (N_4762,N_3024,N_3594);
and U4763 (N_4763,N_3116,N_3345);
nor U4764 (N_4764,N_3601,N_3452);
nor U4765 (N_4765,N_3056,N_3399);
nand U4766 (N_4766,N_3387,N_3766);
or U4767 (N_4767,N_3995,N_3401);
and U4768 (N_4768,N_3032,N_3532);
nor U4769 (N_4769,N_3657,N_3002);
or U4770 (N_4770,N_3222,N_3996);
or U4771 (N_4771,N_3844,N_3470);
nand U4772 (N_4772,N_3311,N_3808);
and U4773 (N_4773,N_3108,N_3083);
nand U4774 (N_4774,N_3133,N_3014);
xnor U4775 (N_4775,N_3535,N_3370);
or U4776 (N_4776,N_3747,N_3855);
nand U4777 (N_4777,N_3926,N_3088);
or U4778 (N_4778,N_3421,N_3377);
or U4779 (N_4779,N_3880,N_3663);
nor U4780 (N_4780,N_3749,N_3389);
nor U4781 (N_4781,N_3939,N_3014);
nand U4782 (N_4782,N_3215,N_3010);
and U4783 (N_4783,N_3462,N_3210);
nor U4784 (N_4784,N_3380,N_3903);
nor U4785 (N_4785,N_3410,N_3643);
and U4786 (N_4786,N_3800,N_3310);
and U4787 (N_4787,N_3842,N_3600);
nor U4788 (N_4788,N_3268,N_3788);
and U4789 (N_4789,N_3223,N_3173);
and U4790 (N_4790,N_3981,N_3112);
nand U4791 (N_4791,N_3515,N_3266);
and U4792 (N_4792,N_3441,N_3110);
nor U4793 (N_4793,N_3962,N_3124);
nand U4794 (N_4794,N_3480,N_3009);
nor U4795 (N_4795,N_3932,N_3217);
nand U4796 (N_4796,N_3523,N_3486);
and U4797 (N_4797,N_3545,N_3316);
and U4798 (N_4798,N_3531,N_3154);
nand U4799 (N_4799,N_3830,N_3642);
nor U4800 (N_4800,N_3915,N_3661);
or U4801 (N_4801,N_3748,N_3142);
nand U4802 (N_4802,N_3685,N_3008);
nand U4803 (N_4803,N_3428,N_3361);
nor U4804 (N_4804,N_3861,N_3833);
nand U4805 (N_4805,N_3633,N_3208);
and U4806 (N_4806,N_3742,N_3875);
and U4807 (N_4807,N_3089,N_3961);
and U4808 (N_4808,N_3039,N_3120);
or U4809 (N_4809,N_3950,N_3354);
and U4810 (N_4810,N_3070,N_3544);
nor U4811 (N_4811,N_3354,N_3424);
nand U4812 (N_4812,N_3892,N_3349);
nor U4813 (N_4813,N_3395,N_3235);
nand U4814 (N_4814,N_3410,N_3877);
and U4815 (N_4815,N_3200,N_3817);
or U4816 (N_4816,N_3784,N_3729);
and U4817 (N_4817,N_3301,N_3954);
and U4818 (N_4818,N_3250,N_3411);
and U4819 (N_4819,N_3376,N_3404);
nand U4820 (N_4820,N_3236,N_3376);
nor U4821 (N_4821,N_3021,N_3085);
nor U4822 (N_4822,N_3116,N_3808);
nand U4823 (N_4823,N_3514,N_3794);
xor U4824 (N_4824,N_3471,N_3022);
nand U4825 (N_4825,N_3953,N_3621);
and U4826 (N_4826,N_3785,N_3535);
xnor U4827 (N_4827,N_3060,N_3601);
nand U4828 (N_4828,N_3445,N_3755);
and U4829 (N_4829,N_3386,N_3023);
nand U4830 (N_4830,N_3851,N_3005);
or U4831 (N_4831,N_3393,N_3790);
nand U4832 (N_4832,N_3381,N_3956);
or U4833 (N_4833,N_3816,N_3586);
nand U4834 (N_4834,N_3747,N_3730);
and U4835 (N_4835,N_3667,N_3365);
nand U4836 (N_4836,N_3012,N_3140);
and U4837 (N_4837,N_3934,N_3256);
nand U4838 (N_4838,N_3138,N_3548);
or U4839 (N_4839,N_3429,N_3274);
nand U4840 (N_4840,N_3345,N_3085);
and U4841 (N_4841,N_3232,N_3014);
nand U4842 (N_4842,N_3088,N_3685);
nand U4843 (N_4843,N_3311,N_3478);
nand U4844 (N_4844,N_3844,N_3224);
nand U4845 (N_4845,N_3015,N_3501);
nand U4846 (N_4846,N_3456,N_3142);
or U4847 (N_4847,N_3214,N_3968);
nand U4848 (N_4848,N_3478,N_3890);
nand U4849 (N_4849,N_3634,N_3805);
nand U4850 (N_4850,N_3897,N_3256);
and U4851 (N_4851,N_3203,N_3655);
nor U4852 (N_4852,N_3139,N_3378);
nand U4853 (N_4853,N_3815,N_3515);
and U4854 (N_4854,N_3542,N_3281);
nor U4855 (N_4855,N_3415,N_3804);
and U4856 (N_4856,N_3487,N_3296);
or U4857 (N_4857,N_3523,N_3753);
nand U4858 (N_4858,N_3161,N_3942);
and U4859 (N_4859,N_3272,N_3242);
or U4860 (N_4860,N_3463,N_3872);
and U4861 (N_4861,N_3047,N_3874);
nand U4862 (N_4862,N_3471,N_3184);
nor U4863 (N_4863,N_3024,N_3004);
nor U4864 (N_4864,N_3428,N_3614);
and U4865 (N_4865,N_3465,N_3289);
nor U4866 (N_4866,N_3100,N_3490);
and U4867 (N_4867,N_3562,N_3895);
or U4868 (N_4868,N_3646,N_3818);
and U4869 (N_4869,N_3283,N_3307);
nor U4870 (N_4870,N_3481,N_3335);
nor U4871 (N_4871,N_3316,N_3896);
and U4872 (N_4872,N_3603,N_3992);
or U4873 (N_4873,N_3796,N_3987);
nand U4874 (N_4874,N_3711,N_3244);
nand U4875 (N_4875,N_3468,N_3886);
nor U4876 (N_4876,N_3347,N_3228);
and U4877 (N_4877,N_3092,N_3921);
or U4878 (N_4878,N_3671,N_3350);
nor U4879 (N_4879,N_3919,N_3619);
or U4880 (N_4880,N_3855,N_3588);
or U4881 (N_4881,N_3893,N_3260);
nand U4882 (N_4882,N_3173,N_3036);
and U4883 (N_4883,N_3708,N_3864);
or U4884 (N_4884,N_3546,N_3276);
and U4885 (N_4885,N_3030,N_3853);
or U4886 (N_4886,N_3325,N_3473);
and U4887 (N_4887,N_3227,N_3432);
nor U4888 (N_4888,N_3463,N_3284);
nor U4889 (N_4889,N_3192,N_3822);
nand U4890 (N_4890,N_3398,N_3332);
nor U4891 (N_4891,N_3859,N_3822);
and U4892 (N_4892,N_3810,N_3135);
and U4893 (N_4893,N_3732,N_3247);
nor U4894 (N_4894,N_3147,N_3697);
nor U4895 (N_4895,N_3576,N_3368);
or U4896 (N_4896,N_3721,N_3815);
and U4897 (N_4897,N_3863,N_3102);
or U4898 (N_4898,N_3936,N_3437);
nand U4899 (N_4899,N_3412,N_3709);
or U4900 (N_4900,N_3757,N_3499);
nor U4901 (N_4901,N_3175,N_3016);
nand U4902 (N_4902,N_3848,N_3724);
nand U4903 (N_4903,N_3057,N_3411);
nor U4904 (N_4904,N_3032,N_3045);
and U4905 (N_4905,N_3550,N_3576);
and U4906 (N_4906,N_3663,N_3246);
nand U4907 (N_4907,N_3833,N_3266);
or U4908 (N_4908,N_3268,N_3819);
nor U4909 (N_4909,N_3079,N_3208);
nor U4910 (N_4910,N_3454,N_3314);
nor U4911 (N_4911,N_3316,N_3125);
or U4912 (N_4912,N_3629,N_3541);
or U4913 (N_4913,N_3330,N_3521);
nand U4914 (N_4914,N_3301,N_3696);
or U4915 (N_4915,N_3312,N_3964);
or U4916 (N_4916,N_3768,N_3616);
nand U4917 (N_4917,N_3311,N_3150);
nand U4918 (N_4918,N_3041,N_3149);
and U4919 (N_4919,N_3832,N_3383);
nand U4920 (N_4920,N_3436,N_3497);
or U4921 (N_4921,N_3223,N_3060);
nand U4922 (N_4922,N_3991,N_3511);
nand U4923 (N_4923,N_3928,N_3907);
and U4924 (N_4924,N_3216,N_3679);
nor U4925 (N_4925,N_3710,N_3406);
and U4926 (N_4926,N_3561,N_3452);
nand U4927 (N_4927,N_3857,N_3585);
nand U4928 (N_4928,N_3172,N_3521);
nand U4929 (N_4929,N_3618,N_3933);
nor U4930 (N_4930,N_3260,N_3967);
and U4931 (N_4931,N_3358,N_3606);
or U4932 (N_4932,N_3387,N_3992);
or U4933 (N_4933,N_3550,N_3108);
nor U4934 (N_4934,N_3502,N_3171);
or U4935 (N_4935,N_3725,N_3739);
nand U4936 (N_4936,N_3953,N_3103);
nor U4937 (N_4937,N_3443,N_3882);
and U4938 (N_4938,N_3391,N_3975);
nor U4939 (N_4939,N_3784,N_3534);
or U4940 (N_4940,N_3139,N_3815);
and U4941 (N_4941,N_3920,N_3733);
and U4942 (N_4942,N_3722,N_3808);
and U4943 (N_4943,N_3401,N_3940);
or U4944 (N_4944,N_3573,N_3402);
nor U4945 (N_4945,N_3314,N_3298);
nand U4946 (N_4946,N_3867,N_3336);
nand U4947 (N_4947,N_3817,N_3393);
or U4948 (N_4948,N_3189,N_3091);
or U4949 (N_4949,N_3330,N_3746);
nor U4950 (N_4950,N_3841,N_3545);
and U4951 (N_4951,N_3527,N_3552);
or U4952 (N_4952,N_3205,N_3280);
or U4953 (N_4953,N_3638,N_3161);
nand U4954 (N_4954,N_3441,N_3211);
and U4955 (N_4955,N_3822,N_3166);
nand U4956 (N_4956,N_3888,N_3515);
and U4957 (N_4957,N_3588,N_3676);
and U4958 (N_4958,N_3232,N_3081);
nand U4959 (N_4959,N_3906,N_3585);
nor U4960 (N_4960,N_3948,N_3048);
or U4961 (N_4961,N_3734,N_3431);
nor U4962 (N_4962,N_3170,N_3598);
or U4963 (N_4963,N_3598,N_3851);
nor U4964 (N_4964,N_3990,N_3318);
and U4965 (N_4965,N_3016,N_3094);
and U4966 (N_4966,N_3728,N_3976);
nor U4967 (N_4967,N_3811,N_3628);
or U4968 (N_4968,N_3918,N_3162);
and U4969 (N_4969,N_3092,N_3258);
and U4970 (N_4970,N_3829,N_3199);
nor U4971 (N_4971,N_3205,N_3632);
and U4972 (N_4972,N_3641,N_3779);
and U4973 (N_4973,N_3622,N_3257);
nand U4974 (N_4974,N_3980,N_3576);
or U4975 (N_4975,N_3272,N_3143);
nand U4976 (N_4976,N_3478,N_3151);
or U4977 (N_4977,N_3665,N_3766);
or U4978 (N_4978,N_3517,N_3380);
nand U4979 (N_4979,N_3170,N_3026);
and U4980 (N_4980,N_3280,N_3552);
nand U4981 (N_4981,N_3442,N_3046);
nor U4982 (N_4982,N_3248,N_3942);
and U4983 (N_4983,N_3600,N_3329);
nand U4984 (N_4984,N_3623,N_3703);
or U4985 (N_4985,N_3101,N_3586);
nor U4986 (N_4986,N_3282,N_3196);
nor U4987 (N_4987,N_3725,N_3054);
nand U4988 (N_4988,N_3712,N_3546);
nor U4989 (N_4989,N_3365,N_3171);
nand U4990 (N_4990,N_3889,N_3334);
nand U4991 (N_4991,N_3576,N_3339);
nand U4992 (N_4992,N_3310,N_3071);
and U4993 (N_4993,N_3759,N_3958);
nand U4994 (N_4994,N_3883,N_3505);
nor U4995 (N_4995,N_3840,N_3975);
xnor U4996 (N_4996,N_3973,N_3777);
and U4997 (N_4997,N_3893,N_3238);
nand U4998 (N_4998,N_3584,N_3512);
and U4999 (N_4999,N_3890,N_3941);
or UO_0 (O_0,N_4846,N_4227);
nor UO_1 (O_1,N_4475,N_4403);
nor UO_2 (O_2,N_4736,N_4716);
and UO_3 (O_3,N_4720,N_4079);
or UO_4 (O_4,N_4534,N_4580);
nor UO_5 (O_5,N_4663,N_4217);
nand UO_6 (O_6,N_4042,N_4059);
and UO_7 (O_7,N_4672,N_4583);
or UO_8 (O_8,N_4589,N_4255);
nor UO_9 (O_9,N_4935,N_4195);
and UO_10 (O_10,N_4727,N_4265);
and UO_11 (O_11,N_4587,N_4464);
nor UO_12 (O_12,N_4687,N_4825);
and UO_13 (O_13,N_4375,N_4602);
and UO_14 (O_14,N_4980,N_4168);
nor UO_15 (O_15,N_4396,N_4544);
or UO_16 (O_16,N_4940,N_4204);
or UO_17 (O_17,N_4837,N_4756);
nor UO_18 (O_18,N_4131,N_4325);
or UO_19 (O_19,N_4926,N_4271);
xnor UO_20 (O_20,N_4424,N_4369);
nand UO_21 (O_21,N_4680,N_4807);
nand UO_22 (O_22,N_4060,N_4330);
nand UO_23 (O_23,N_4921,N_4272);
and UO_24 (O_24,N_4978,N_4302);
and UO_25 (O_25,N_4838,N_4235);
or UO_26 (O_26,N_4642,N_4536);
or UO_27 (O_27,N_4684,N_4392);
or UO_28 (O_28,N_4713,N_4465);
nand UO_29 (O_29,N_4707,N_4327);
nand UO_30 (O_30,N_4755,N_4655);
and UO_31 (O_31,N_4632,N_4329);
nand UO_32 (O_32,N_4092,N_4076);
or UO_33 (O_33,N_4282,N_4426);
and UO_34 (O_34,N_4202,N_4947);
nand UO_35 (O_35,N_4192,N_4667);
nand UO_36 (O_36,N_4505,N_4117);
and UO_37 (O_37,N_4034,N_4022);
nor UO_38 (O_38,N_4001,N_4652);
and UO_39 (O_39,N_4733,N_4520);
nand UO_40 (O_40,N_4695,N_4798);
nand UO_41 (O_41,N_4146,N_4510);
or UO_42 (O_42,N_4898,N_4486);
and UO_43 (O_43,N_4135,N_4774);
or UO_44 (O_44,N_4409,N_4347);
nand UO_45 (O_45,N_4381,N_4547);
and UO_46 (O_46,N_4306,N_4918);
nor UO_47 (O_47,N_4213,N_4915);
or UO_48 (O_48,N_4961,N_4592);
nand UO_49 (O_49,N_4366,N_4887);
and UO_50 (O_50,N_4523,N_4710);
nor UO_51 (O_51,N_4087,N_4140);
or UO_52 (O_52,N_4964,N_4454);
nor UO_53 (O_53,N_4574,N_4145);
nor UO_54 (O_54,N_4990,N_4346);
or UO_55 (O_55,N_4788,N_4591);
nor UO_56 (O_56,N_4723,N_4354);
nor UO_57 (O_57,N_4223,N_4616);
and UO_58 (O_58,N_4842,N_4761);
nor UO_59 (O_59,N_4515,N_4112);
or UO_60 (O_60,N_4276,N_4446);
and UO_61 (O_61,N_4046,N_4634);
and UO_62 (O_62,N_4780,N_4872);
nand UO_63 (O_63,N_4316,N_4064);
nor UO_64 (O_64,N_4658,N_4670);
and UO_65 (O_65,N_4702,N_4814);
nand UO_66 (O_66,N_4850,N_4712);
or UO_67 (O_67,N_4675,N_4007);
and UO_68 (O_68,N_4199,N_4402);
nor UO_69 (O_69,N_4136,N_4167);
or UO_70 (O_70,N_4700,N_4533);
nand UO_71 (O_71,N_4002,N_4690);
nor UO_72 (O_72,N_4401,N_4953);
nand UO_73 (O_73,N_4806,N_4047);
nand UO_74 (O_74,N_4483,N_4252);
or UO_75 (O_75,N_4596,N_4019);
nor UO_76 (O_76,N_4422,N_4373);
nand UO_77 (O_77,N_4154,N_4037);
or UO_78 (O_78,N_4705,N_4758);
and UO_79 (O_79,N_4543,N_4304);
nor UO_80 (O_80,N_4012,N_4179);
or UO_81 (O_81,N_4169,N_4597);
nor UO_82 (O_82,N_4508,N_4086);
or UO_83 (O_83,N_4778,N_4718);
nor UO_84 (O_84,N_4811,N_4450);
or UO_85 (O_85,N_4228,N_4841);
and UO_86 (O_86,N_4506,N_4932);
nand UO_87 (O_87,N_4925,N_4423);
nor UO_88 (O_88,N_4539,N_4786);
nor UO_89 (O_89,N_4907,N_4490);
nand UO_90 (O_90,N_4879,N_4929);
nand UO_91 (O_91,N_4818,N_4630);
nor UO_92 (O_92,N_4903,N_4939);
nor UO_93 (O_93,N_4350,N_4560);
nor UO_94 (O_94,N_4793,N_4004);
nor UO_95 (O_95,N_4998,N_4966);
and UO_96 (O_96,N_4664,N_4683);
nand UO_97 (O_97,N_4671,N_4744);
nor UO_98 (O_98,N_4899,N_4686);
nand UO_99 (O_99,N_4342,N_4886);
nor UO_100 (O_100,N_4598,N_4126);
or UO_101 (O_101,N_4495,N_4882);
nor UO_102 (O_102,N_4181,N_4868);
nand UO_103 (O_103,N_4698,N_4288);
or UO_104 (O_104,N_4100,N_4021);
xor UO_105 (O_105,N_4751,N_4128);
and UO_106 (O_106,N_4413,N_4305);
and UO_107 (O_107,N_4732,N_4269);
nand UO_108 (O_108,N_4055,N_4258);
nand UO_109 (O_109,N_4447,N_4323);
nor UO_110 (O_110,N_4057,N_4906);
nor UO_111 (O_111,N_4562,N_4324);
nor UO_112 (O_112,N_4437,N_4032);
or UO_113 (O_113,N_4456,N_4063);
or UO_114 (O_114,N_4708,N_4922);
and UO_115 (O_115,N_4928,N_4586);
nor UO_116 (O_116,N_4296,N_4514);
or UO_117 (O_117,N_4322,N_4773);
nand UO_118 (O_118,N_4985,N_4274);
or UO_119 (O_119,N_4239,N_4127);
nor UO_120 (O_120,N_4895,N_4072);
and UO_121 (O_121,N_4476,N_4576);
nor UO_122 (O_122,N_4243,N_4648);
or UO_123 (O_123,N_4541,N_4949);
nand UO_124 (O_124,N_4266,N_4008);
nor UO_125 (O_125,N_4999,N_4113);
nand UO_126 (O_126,N_4451,N_4645);
or UO_127 (O_127,N_4384,N_4378);
nand UO_128 (O_128,N_4000,N_4083);
and UO_129 (O_129,N_4704,N_4196);
or UO_130 (O_130,N_4877,N_4362);
or UO_131 (O_131,N_4155,N_4283);
and UO_132 (O_132,N_4280,N_4784);
and UO_133 (O_133,N_4654,N_4003);
and UO_134 (O_134,N_4018,N_4105);
or UO_135 (O_135,N_4442,N_4689);
or UO_136 (O_136,N_4631,N_4443);
and UO_137 (O_137,N_4738,N_4946);
nand UO_138 (O_138,N_4184,N_4270);
and UO_139 (O_139,N_4029,N_4200);
nor UO_140 (O_140,N_4635,N_4153);
or UO_141 (O_141,N_4754,N_4367);
nor UO_142 (O_142,N_4555,N_4656);
nor UO_143 (O_143,N_4605,N_4688);
nand UO_144 (O_144,N_4933,N_4035);
xnor UO_145 (O_145,N_4352,N_4830);
nor UO_146 (O_146,N_4676,N_4649);
nor UO_147 (O_147,N_4237,N_4114);
and UO_148 (O_148,N_4344,N_4979);
nand UO_149 (O_149,N_4885,N_4130);
and UO_150 (O_150,N_4393,N_4318);
nor UO_151 (O_151,N_4441,N_4452);
nor UO_152 (O_152,N_4365,N_4682);
or UO_153 (O_153,N_4789,N_4428);
nor UO_154 (O_154,N_4870,N_4578);
or UO_155 (O_155,N_4822,N_4388);
or UO_156 (O_156,N_4833,N_4777);
or UO_157 (O_157,N_4829,N_4660);
nand UO_158 (O_158,N_4499,N_4397);
nand UO_159 (O_159,N_4124,N_4721);
and UO_160 (O_160,N_4760,N_4226);
or UO_161 (O_161,N_4799,N_4275);
nor UO_162 (O_162,N_4479,N_4488);
nor UO_163 (O_163,N_4024,N_4971);
nor UO_164 (O_164,N_4349,N_4896);
nor UO_165 (O_165,N_4033,N_4313);
nor UO_166 (O_166,N_4828,N_4414);
and UO_167 (O_167,N_4627,N_4026);
or UO_168 (O_168,N_4530,N_4876);
or UO_169 (O_169,N_4489,N_4449);
nor UO_170 (O_170,N_4015,N_4232);
nand UO_171 (O_171,N_4524,N_4636);
nand UO_172 (O_172,N_4501,N_4585);
nand UO_173 (O_173,N_4400,N_4206);
or UO_174 (O_174,N_4963,N_4750);
nor UO_175 (O_175,N_4041,N_4207);
nand UO_176 (O_176,N_4607,N_4208);
or UO_177 (O_177,N_4247,N_4201);
and UO_178 (O_178,N_4492,N_4725);
nand UO_179 (O_179,N_4189,N_4427);
and UO_180 (O_180,N_4817,N_4823);
and UO_181 (O_181,N_4281,N_4144);
nand UO_182 (O_182,N_4038,N_4930);
and UO_183 (O_183,N_4858,N_4336);
nor UO_184 (O_184,N_4808,N_4170);
nor UO_185 (O_185,N_4711,N_4372);
and UO_186 (O_186,N_4279,N_4941);
nand UO_187 (O_187,N_4741,N_4995);
nor UO_188 (O_188,N_4116,N_4078);
or UO_189 (O_189,N_4463,N_4093);
and UO_190 (O_190,N_4977,N_4861);
or UO_191 (O_191,N_4259,N_4225);
nor UO_192 (O_192,N_4053,N_4976);
or UO_193 (O_193,N_4440,N_4867);
nand UO_194 (O_194,N_4389,N_4640);
nand UO_195 (O_195,N_4728,N_4952);
nor UO_196 (O_196,N_4466,N_4852);
or UO_197 (O_197,N_4161,N_4783);
and UO_198 (O_198,N_4659,N_4923);
and UO_199 (O_199,N_4438,N_4950);
nand UO_200 (O_200,N_4968,N_4693);
nor UO_201 (O_201,N_4565,N_4415);
or UO_202 (O_202,N_4874,N_4070);
or UO_203 (O_203,N_4509,N_4717);
or UO_204 (O_204,N_4561,N_4795);
nand UO_205 (O_205,N_4782,N_4694);
nor UO_206 (O_206,N_4250,N_4892);
or UO_207 (O_207,N_4881,N_4317);
or UO_208 (O_208,N_4900,N_4832);
nand UO_209 (O_209,N_4519,N_4287);
and UO_210 (O_210,N_4066,N_4512);
or UO_211 (O_211,N_4101,N_4332);
and UO_212 (O_212,N_4956,N_4757);
nand UO_213 (O_213,N_4913,N_4297);
or UO_214 (O_214,N_4133,N_4821);
and UO_215 (O_215,N_4469,N_4831);
nand UO_216 (O_216,N_4851,N_4374);
and UO_217 (O_217,N_4395,N_4107);
nor UO_218 (O_218,N_4039,N_4550);
or UO_219 (O_219,N_4188,N_4238);
or UO_220 (O_220,N_4610,N_4657);
or UO_221 (O_221,N_4730,N_4859);
or UO_222 (O_222,N_4142,N_4612);
nand UO_223 (O_223,N_4827,N_4319);
nand UO_224 (O_224,N_4430,N_4884);
or UO_225 (O_225,N_4094,N_4575);
nand UO_226 (O_226,N_4767,N_4665);
or UO_227 (O_227,N_4531,N_4912);
nand UO_228 (O_228,N_4256,N_4084);
or UO_229 (O_229,N_4090,N_4701);
nand UO_230 (O_230,N_4944,N_4845);
nor UO_231 (O_231,N_4320,N_4740);
nor UO_232 (O_232,N_4425,N_4293);
nand UO_233 (O_233,N_4299,N_4068);
and UO_234 (O_234,N_4244,N_4061);
nor UO_235 (O_235,N_4706,N_4253);
or UO_236 (O_236,N_4205,N_4997);
nor UO_237 (O_237,N_4969,N_4198);
nor UO_238 (O_238,N_4099,N_4407);
nor UO_239 (O_239,N_4960,N_4633);
and UO_240 (O_240,N_4622,N_4163);
and UO_241 (O_241,N_4171,N_4159);
nor UO_242 (O_242,N_4219,N_4230);
nor UO_243 (O_243,N_4257,N_4538);
nand UO_244 (O_244,N_4996,N_4848);
or UO_245 (O_245,N_4781,N_4242);
nand UO_246 (O_246,N_4847,N_4310);
and UO_247 (O_247,N_4143,N_4584);
and UO_248 (O_248,N_4745,N_4518);
or UO_249 (O_249,N_4855,N_4759);
nand UO_250 (O_250,N_4156,N_4085);
and UO_251 (O_251,N_4044,N_4945);
or UO_252 (O_252,N_4618,N_4412);
nand UO_253 (O_253,N_4417,N_4619);
nor UO_254 (O_254,N_4890,N_4233);
or UO_255 (O_255,N_4766,N_4360);
nor UO_256 (O_256,N_4286,N_4569);
nor UO_257 (O_257,N_4908,N_4540);
nand UO_258 (O_258,N_4298,N_4069);
and UO_259 (O_259,N_4709,N_4992);
and UO_260 (O_260,N_4314,N_4074);
or UO_261 (O_261,N_4629,N_4160);
and UO_262 (O_262,N_4615,N_4762);
nor UO_263 (O_263,N_4497,N_4308);
and UO_264 (O_264,N_4394,N_4715);
and UO_265 (O_265,N_4726,N_4385);
and UO_266 (O_266,N_4662,N_4609);
nand UO_267 (O_267,N_4028,N_4182);
nand UO_268 (O_268,N_4871,N_4432);
nand UO_269 (O_269,N_4503,N_4975);
nand UO_270 (O_270,N_4771,N_4218);
and UO_271 (O_271,N_4348,N_4493);
nor UO_272 (O_272,N_4611,N_4548);
and UO_273 (O_273,N_4666,N_4284);
nand UO_274 (O_274,N_4473,N_4109);
and UO_275 (O_275,N_4909,N_4088);
and UO_276 (O_276,N_4797,N_4873);
and UO_277 (O_277,N_4644,N_4641);
nand UO_278 (O_278,N_4962,N_4563);
or UO_279 (O_279,N_4719,N_4516);
nor UO_280 (O_280,N_4535,N_4368);
or UO_281 (O_281,N_4058,N_4681);
xnor UO_282 (O_282,N_4125,N_4815);
nor UO_283 (O_283,N_4460,N_4957);
nor UO_284 (O_284,N_4056,N_4804);
or UO_285 (O_285,N_4231,N_4674);
nor UO_286 (O_286,N_4164,N_4307);
or UO_287 (O_287,N_4528,N_4785);
nand UO_288 (O_288,N_4857,N_4234);
or UO_289 (O_289,N_4986,N_4948);
xor UO_290 (O_290,N_4370,N_4052);
or UO_291 (O_291,N_4262,N_4601);
nor UO_292 (O_292,N_4186,N_4193);
nand UO_293 (O_293,N_4934,N_4025);
and UO_294 (O_294,N_4119,N_4180);
nand UO_295 (O_295,N_4120,N_4434);
nor UO_296 (O_296,N_4474,N_4418);
and UO_297 (O_297,N_4178,N_4731);
nand UO_298 (O_298,N_4608,N_4328);
or UO_299 (O_299,N_4746,N_4138);
nand UO_300 (O_300,N_4590,N_4445);
or UO_301 (O_301,N_4691,N_4606);
nand UO_302 (O_302,N_4439,N_4511);
or UO_303 (O_303,N_4914,N_4924);
and UO_304 (O_304,N_4151,N_4340);
nand UO_305 (O_305,N_4916,N_4987);
nor UO_306 (O_306,N_4954,N_4062);
or UO_307 (O_307,N_4739,N_4300);
and UO_308 (O_308,N_4507,N_4301);
or UO_309 (O_309,N_4653,N_4927);
or UO_310 (O_310,N_4840,N_4097);
and UO_311 (O_311,N_4826,N_4175);
nor UO_312 (O_312,N_4856,N_4537);
nor UO_313 (O_313,N_4498,N_4568);
nor UO_314 (O_314,N_4377,N_4137);
or UO_315 (O_315,N_4553,N_4714);
or UO_316 (O_316,N_4054,N_4936);
and UO_317 (O_317,N_4593,N_4787);
and UO_318 (O_318,N_4549,N_4617);
or UO_319 (O_319,N_4210,N_4311);
or UO_320 (O_320,N_4792,N_4991);
nand UO_321 (O_321,N_4546,N_4897);
or UO_322 (O_322,N_4812,N_4291);
nand UO_323 (O_323,N_4545,N_4770);
and UO_324 (O_324,N_4677,N_4165);
nor UO_325 (O_325,N_4118,N_4970);
and UO_326 (O_326,N_4485,N_4567);
nor UO_327 (O_327,N_4240,N_4212);
nor UO_328 (O_328,N_4431,N_4371);
or UO_329 (O_329,N_4095,N_4277);
and UO_330 (O_330,N_4579,N_4254);
and UO_331 (O_331,N_4863,N_4215);
or UO_332 (O_332,N_4875,N_4429);
nor UO_333 (O_333,N_4190,N_4955);
and UO_334 (O_334,N_4902,N_4920);
nor UO_335 (O_335,N_4480,N_4309);
and UO_336 (O_336,N_4264,N_4835);
or UO_337 (O_337,N_4108,N_4448);
and UO_338 (O_338,N_4468,N_4526);
or UO_339 (O_339,N_4843,N_4889);
and UO_340 (O_340,N_4355,N_4410);
nand UO_341 (O_341,N_4643,N_4292);
nand UO_342 (O_342,N_4134,N_4809);
nand UO_343 (O_343,N_4864,N_4260);
and UO_344 (O_344,N_4742,N_4484);
or UO_345 (O_345,N_4129,N_4571);
nand UO_346 (O_346,N_4819,N_4263);
and UO_347 (O_347,N_4361,N_4343);
or UO_348 (O_348,N_4158,N_4764);
and UO_349 (O_349,N_4749,N_4768);
or UO_350 (O_350,N_4236,N_4071);
or UO_351 (O_351,N_4974,N_4624);
and UO_352 (O_352,N_4457,N_4183);
nor UO_353 (O_353,N_4901,N_4075);
and UO_354 (O_354,N_4581,N_4836);
or UO_355 (O_355,N_4800,N_4339);
and UO_356 (O_356,N_4647,N_4982);
nand UO_357 (O_357,N_4883,N_4267);
nor UO_358 (O_358,N_4931,N_4839);
nor UO_359 (O_359,N_4132,N_4013);
and UO_360 (O_360,N_4203,N_4917);
nor UO_361 (O_361,N_4743,N_4172);
nor UO_362 (O_362,N_4104,N_4331);
nand UO_363 (O_363,N_4091,N_4650);
nor UO_364 (O_364,N_4081,N_4834);
or UO_365 (O_365,N_4734,N_4379);
nor UO_366 (O_366,N_4249,N_4905);
nor UO_367 (O_367,N_4628,N_4696);
nor UO_368 (O_368,N_4421,N_4794);
or UO_369 (O_369,N_4559,N_4157);
nor UO_370 (O_370,N_4775,N_4338);
nor UO_371 (O_371,N_4082,N_4853);
and UO_372 (O_372,N_4595,N_4220);
nand UO_373 (O_373,N_4865,N_4737);
nor UO_374 (O_374,N_4027,N_4194);
nor UO_375 (O_375,N_4994,N_4894);
and UO_376 (O_376,N_4214,N_4067);
and UO_377 (O_377,N_4639,N_4123);
nand UO_378 (O_378,N_4216,N_4405);
and UO_379 (O_379,N_4358,N_4176);
or UO_380 (O_380,N_4152,N_4011);
or UO_381 (O_381,N_4747,N_4573);
nor UO_382 (O_382,N_4345,N_4315);
nor UO_383 (O_383,N_4891,N_4461);
or UO_384 (O_384,N_4391,N_4139);
or UO_385 (O_385,N_4174,N_4014);
nor UO_386 (O_386,N_4937,N_4211);
nand UO_387 (O_387,N_4919,N_4522);
nand UO_388 (O_388,N_4722,N_4387);
nand UO_389 (O_389,N_4577,N_4462);
nand UO_390 (O_390,N_4436,N_4491);
and UO_391 (O_391,N_4763,N_4382);
nand UO_392 (O_392,N_4604,N_4525);
or UO_393 (O_393,N_4866,N_4010);
nand UO_394 (O_394,N_4110,N_4527);
nor UO_395 (O_395,N_4353,N_4496);
and UO_396 (O_396,N_4285,N_4599);
nor UO_397 (O_397,N_4162,N_4261);
nand UO_398 (O_398,N_4294,N_4951);
and UO_399 (O_399,N_4209,N_4096);
and UO_400 (O_400,N_4009,N_4564);
nor UO_401 (O_401,N_4295,N_4472);
or UO_402 (O_402,N_4661,N_4869);
nand UO_403 (O_403,N_4073,N_4433);
and UO_404 (O_404,N_4023,N_4542);
or UO_405 (O_405,N_4459,N_4359);
or UO_406 (O_406,N_4790,N_4552);
nor UO_407 (O_407,N_4036,N_4185);
nand UO_408 (O_408,N_4849,N_4411);
and UO_409 (O_409,N_4048,N_4844);
nand UO_410 (O_410,N_4582,N_4791);
nor UO_411 (O_411,N_4245,N_4748);
xnor UO_412 (O_412,N_4638,N_4221);
nor UO_413 (O_413,N_4416,N_4621);
nand UO_414 (O_414,N_4435,N_4697);
or UO_415 (O_415,N_4983,N_4685);
and UO_416 (O_416,N_4471,N_4769);
xor UO_417 (O_417,N_4121,N_4098);
and UO_418 (O_418,N_4993,N_4824);
and UO_419 (O_419,N_4248,N_4357);
and UO_420 (O_420,N_4419,N_4805);
or UO_421 (O_421,N_4625,N_4149);
nor UO_422 (O_422,N_4398,N_4984);
nand UO_423 (O_423,N_4802,N_4572);
nand UO_424 (O_424,N_4521,N_4187);
nor UO_425 (O_425,N_4326,N_4752);
nand UO_426 (O_426,N_4988,N_4958);
or UO_427 (O_427,N_4080,N_4888);
nand UO_428 (O_428,N_4973,N_4341);
and UO_429 (O_429,N_4753,N_4729);
or UO_430 (O_430,N_4532,N_4513);
nand UO_431 (O_431,N_4065,N_4017);
and UO_432 (O_432,N_4453,N_4494);
or UO_433 (O_433,N_4614,N_4333);
xnor UO_434 (O_434,N_4570,N_4620);
nand UO_435 (O_435,N_4289,N_4406);
nand UO_436 (O_436,N_4481,N_4989);
or UO_437 (O_437,N_4045,N_4278);
or UO_438 (O_438,N_4404,N_4651);
nor UO_439 (O_439,N_4363,N_4197);
nand UO_440 (O_440,N_4177,N_4600);
or UO_441 (O_441,N_4222,N_4478);
nor UO_442 (O_442,N_4273,N_4408);
and UO_443 (O_443,N_4102,N_4594);
or UO_444 (O_444,N_4303,N_4005);
nor UO_445 (O_445,N_4487,N_4673);
nor UO_446 (O_446,N_4588,N_4959);
nor UO_447 (O_447,N_4965,N_4904);
and UO_448 (O_448,N_4796,N_4376);
and UO_449 (O_449,N_4943,N_4334);
nand UO_450 (O_450,N_4699,N_4455);
nand UO_451 (O_451,N_4241,N_4312);
and UO_452 (O_452,N_4893,N_4938);
and UO_453 (O_453,N_4356,N_4030);
nand UO_454 (O_454,N_4810,N_4551);
and UO_455 (O_455,N_4290,N_4860);
or UO_456 (O_456,N_4477,N_4268);
nand UO_457 (O_457,N_4111,N_4517);
nor UO_458 (O_458,N_4386,N_4558);
nand UO_459 (O_459,N_4482,N_4504);
or UO_460 (O_460,N_4229,N_4967);
nor UO_461 (O_461,N_4458,N_4813);
or UO_462 (O_462,N_4779,N_4335);
nor UO_463 (O_463,N_4420,N_4972);
or UO_464 (O_464,N_4724,N_4051);
and UO_465 (O_465,N_4646,N_4089);
nor UO_466 (O_466,N_4141,N_4557);
nand UO_467 (O_467,N_4981,N_4820);
and UO_468 (O_468,N_4500,N_4173);
and UO_469 (O_469,N_4043,N_4390);
and UO_470 (O_470,N_4467,N_4880);
nor UO_471 (O_471,N_4016,N_4050);
nor UO_472 (O_472,N_4803,N_4364);
or UO_473 (O_473,N_4878,N_4668);
nor UO_474 (O_474,N_4031,N_4556);
nor UO_475 (O_475,N_4049,N_4251);
nor UO_476 (O_476,N_4103,N_4383);
nor UO_477 (O_477,N_4191,N_4246);
nand UO_478 (O_478,N_4765,N_4077);
and UO_479 (O_479,N_4862,N_4380);
or UO_480 (O_480,N_4776,N_4147);
and UO_481 (O_481,N_4623,N_4337);
nor UO_482 (O_482,N_4942,N_4735);
nor UO_483 (O_483,N_4224,N_4502);
and UO_484 (O_484,N_4566,N_4816);
and UO_485 (O_485,N_4801,N_4637);
nor UO_486 (O_486,N_4006,N_4603);
and UO_487 (O_487,N_4122,N_4772);
nor UO_488 (O_488,N_4613,N_4399);
nand UO_489 (O_489,N_4529,N_4321);
and UO_490 (O_490,N_4692,N_4669);
and UO_491 (O_491,N_4703,N_4115);
nor UO_492 (O_492,N_4444,N_4626);
and UO_493 (O_493,N_4040,N_4678);
and UO_494 (O_494,N_4166,N_4910);
nand UO_495 (O_495,N_4911,N_4470);
or UO_496 (O_496,N_4020,N_4150);
nor UO_497 (O_497,N_4679,N_4854);
nor UO_498 (O_498,N_4554,N_4351);
nor UO_499 (O_499,N_4148,N_4106);
xor UO_500 (O_500,N_4715,N_4080);
and UO_501 (O_501,N_4635,N_4754);
and UO_502 (O_502,N_4680,N_4911);
nor UO_503 (O_503,N_4232,N_4481);
or UO_504 (O_504,N_4509,N_4230);
nor UO_505 (O_505,N_4510,N_4226);
nor UO_506 (O_506,N_4429,N_4624);
and UO_507 (O_507,N_4088,N_4077);
nand UO_508 (O_508,N_4754,N_4342);
or UO_509 (O_509,N_4654,N_4984);
nor UO_510 (O_510,N_4832,N_4268);
and UO_511 (O_511,N_4131,N_4478);
nor UO_512 (O_512,N_4239,N_4874);
nand UO_513 (O_513,N_4241,N_4429);
nand UO_514 (O_514,N_4586,N_4843);
nor UO_515 (O_515,N_4906,N_4800);
nor UO_516 (O_516,N_4601,N_4246);
nand UO_517 (O_517,N_4646,N_4332);
and UO_518 (O_518,N_4801,N_4961);
nand UO_519 (O_519,N_4650,N_4613);
or UO_520 (O_520,N_4431,N_4023);
or UO_521 (O_521,N_4425,N_4866);
nor UO_522 (O_522,N_4857,N_4020);
or UO_523 (O_523,N_4692,N_4103);
xor UO_524 (O_524,N_4557,N_4285);
or UO_525 (O_525,N_4714,N_4319);
or UO_526 (O_526,N_4721,N_4967);
or UO_527 (O_527,N_4945,N_4931);
or UO_528 (O_528,N_4780,N_4259);
and UO_529 (O_529,N_4531,N_4921);
nand UO_530 (O_530,N_4249,N_4909);
and UO_531 (O_531,N_4177,N_4174);
and UO_532 (O_532,N_4147,N_4164);
and UO_533 (O_533,N_4288,N_4644);
nand UO_534 (O_534,N_4466,N_4174);
nand UO_535 (O_535,N_4868,N_4325);
nor UO_536 (O_536,N_4604,N_4522);
or UO_537 (O_537,N_4918,N_4647);
and UO_538 (O_538,N_4899,N_4087);
and UO_539 (O_539,N_4097,N_4685);
nand UO_540 (O_540,N_4922,N_4981);
and UO_541 (O_541,N_4507,N_4410);
and UO_542 (O_542,N_4557,N_4396);
nor UO_543 (O_543,N_4903,N_4518);
and UO_544 (O_544,N_4552,N_4742);
and UO_545 (O_545,N_4594,N_4873);
nand UO_546 (O_546,N_4565,N_4556);
nor UO_547 (O_547,N_4666,N_4022);
and UO_548 (O_548,N_4820,N_4141);
nor UO_549 (O_549,N_4880,N_4210);
nor UO_550 (O_550,N_4164,N_4163);
nand UO_551 (O_551,N_4719,N_4658);
and UO_552 (O_552,N_4211,N_4686);
nand UO_553 (O_553,N_4928,N_4550);
nor UO_554 (O_554,N_4131,N_4918);
or UO_555 (O_555,N_4287,N_4282);
nand UO_556 (O_556,N_4988,N_4511);
or UO_557 (O_557,N_4681,N_4622);
nor UO_558 (O_558,N_4459,N_4579);
or UO_559 (O_559,N_4591,N_4222);
nor UO_560 (O_560,N_4701,N_4923);
and UO_561 (O_561,N_4854,N_4115);
or UO_562 (O_562,N_4800,N_4719);
or UO_563 (O_563,N_4466,N_4776);
nand UO_564 (O_564,N_4212,N_4307);
and UO_565 (O_565,N_4220,N_4575);
or UO_566 (O_566,N_4692,N_4685);
xnor UO_567 (O_567,N_4447,N_4462);
and UO_568 (O_568,N_4343,N_4718);
nand UO_569 (O_569,N_4275,N_4099);
nand UO_570 (O_570,N_4414,N_4501);
and UO_571 (O_571,N_4354,N_4312);
and UO_572 (O_572,N_4106,N_4724);
and UO_573 (O_573,N_4081,N_4456);
or UO_574 (O_574,N_4447,N_4467);
or UO_575 (O_575,N_4622,N_4043);
or UO_576 (O_576,N_4669,N_4838);
nand UO_577 (O_577,N_4708,N_4202);
or UO_578 (O_578,N_4364,N_4275);
and UO_579 (O_579,N_4804,N_4133);
nand UO_580 (O_580,N_4535,N_4558);
or UO_581 (O_581,N_4391,N_4011);
nand UO_582 (O_582,N_4978,N_4982);
or UO_583 (O_583,N_4676,N_4437);
or UO_584 (O_584,N_4342,N_4494);
or UO_585 (O_585,N_4484,N_4122);
nand UO_586 (O_586,N_4542,N_4622);
and UO_587 (O_587,N_4884,N_4519);
nor UO_588 (O_588,N_4301,N_4156);
nor UO_589 (O_589,N_4571,N_4590);
nand UO_590 (O_590,N_4218,N_4908);
and UO_591 (O_591,N_4928,N_4923);
nand UO_592 (O_592,N_4871,N_4890);
and UO_593 (O_593,N_4806,N_4361);
nor UO_594 (O_594,N_4070,N_4807);
or UO_595 (O_595,N_4985,N_4689);
or UO_596 (O_596,N_4549,N_4443);
nand UO_597 (O_597,N_4796,N_4051);
nand UO_598 (O_598,N_4150,N_4181);
nor UO_599 (O_599,N_4040,N_4189);
or UO_600 (O_600,N_4519,N_4638);
nor UO_601 (O_601,N_4872,N_4864);
or UO_602 (O_602,N_4673,N_4516);
nor UO_603 (O_603,N_4057,N_4550);
or UO_604 (O_604,N_4953,N_4145);
nor UO_605 (O_605,N_4995,N_4213);
nor UO_606 (O_606,N_4755,N_4468);
nor UO_607 (O_607,N_4053,N_4717);
and UO_608 (O_608,N_4910,N_4841);
and UO_609 (O_609,N_4867,N_4542);
nand UO_610 (O_610,N_4861,N_4224);
nor UO_611 (O_611,N_4686,N_4702);
or UO_612 (O_612,N_4903,N_4984);
or UO_613 (O_613,N_4625,N_4800);
and UO_614 (O_614,N_4259,N_4736);
or UO_615 (O_615,N_4267,N_4415);
nand UO_616 (O_616,N_4691,N_4614);
nor UO_617 (O_617,N_4299,N_4146);
xor UO_618 (O_618,N_4967,N_4803);
and UO_619 (O_619,N_4736,N_4219);
and UO_620 (O_620,N_4669,N_4390);
or UO_621 (O_621,N_4371,N_4030);
nor UO_622 (O_622,N_4118,N_4081);
nor UO_623 (O_623,N_4908,N_4078);
nand UO_624 (O_624,N_4286,N_4076);
or UO_625 (O_625,N_4585,N_4098);
or UO_626 (O_626,N_4793,N_4296);
and UO_627 (O_627,N_4955,N_4105);
or UO_628 (O_628,N_4256,N_4228);
or UO_629 (O_629,N_4515,N_4974);
or UO_630 (O_630,N_4131,N_4208);
or UO_631 (O_631,N_4222,N_4273);
and UO_632 (O_632,N_4132,N_4261);
xnor UO_633 (O_633,N_4839,N_4296);
and UO_634 (O_634,N_4774,N_4694);
nand UO_635 (O_635,N_4228,N_4967);
or UO_636 (O_636,N_4511,N_4171);
nand UO_637 (O_637,N_4968,N_4301);
nor UO_638 (O_638,N_4008,N_4076);
or UO_639 (O_639,N_4255,N_4007);
and UO_640 (O_640,N_4521,N_4755);
and UO_641 (O_641,N_4736,N_4903);
nand UO_642 (O_642,N_4041,N_4028);
nor UO_643 (O_643,N_4732,N_4896);
and UO_644 (O_644,N_4468,N_4377);
nand UO_645 (O_645,N_4349,N_4103);
and UO_646 (O_646,N_4338,N_4586);
nand UO_647 (O_647,N_4313,N_4232);
and UO_648 (O_648,N_4195,N_4298);
and UO_649 (O_649,N_4910,N_4686);
nand UO_650 (O_650,N_4347,N_4179);
xnor UO_651 (O_651,N_4618,N_4023);
nor UO_652 (O_652,N_4264,N_4163);
or UO_653 (O_653,N_4661,N_4949);
nand UO_654 (O_654,N_4285,N_4244);
nor UO_655 (O_655,N_4696,N_4723);
nor UO_656 (O_656,N_4314,N_4717);
nand UO_657 (O_657,N_4285,N_4681);
nand UO_658 (O_658,N_4656,N_4951);
or UO_659 (O_659,N_4459,N_4358);
and UO_660 (O_660,N_4040,N_4205);
and UO_661 (O_661,N_4107,N_4005);
and UO_662 (O_662,N_4412,N_4756);
nor UO_663 (O_663,N_4926,N_4033);
nand UO_664 (O_664,N_4715,N_4524);
nand UO_665 (O_665,N_4633,N_4762);
or UO_666 (O_666,N_4535,N_4427);
nand UO_667 (O_667,N_4147,N_4121);
or UO_668 (O_668,N_4768,N_4111);
or UO_669 (O_669,N_4362,N_4514);
nand UO_670 (O_670,N_4848,N_4092);
nor UO_671 (O_671,N_4588,N_4632);
or UO_672 (O_672,N_4318,N_4413);
and UO_673 (O_673,N_4824,N_4600);
or UO_674 (O_674,N_4016,N_4222);
nand UO_675 (O_675,N_4566,N_4040);
or UO_676 (O_676,N_4963,N_4649);
or UO_677 (O_677,N_4181,N_4263);
or UO_678 (O_678,N_4859,N_4619);
and UO_679 (O_679,N_4890,N_4003);
and UO_680 (O_680,N_4562,N_4027);
nand UO_681 (O_681,N_4231,N_4383);
and UO_682 (O_682,N_4785,N_4096);
and UO_683 (O_683,N_4484,N_4971);
nor UO_684 (O_684,N_4099,N_4477);
nand UO_685 (O_685,N_4121,N_4778);
nand UO_686 (O_686,N_4920,N_4984);
and UO_687 (O_687,N_4977,N_4231);
nor UO_688 (O_688,N_4818,N_4386);
and UO_689 (O_689,N_4794,N_4383);
and UO_690 (O_690,N_4955,N_4887);
nand UO_691 (O_691,N_4261,N_4133);
or UO_692 (O_692,N_4483,N_4372);
nand UO_693 (O_693,N_4336,N_4166);
nor UO_694 (O_694,N_4090,N_4293);
nand UO_695 (O_695,N_4554,N_4597);
xor UO_696 (O_696,N_4962,N_4049);
or UO_697 (O_697,N_4327,N_4749);
nand UO_698 (O_698,N_4703,N_4446);
or UO_699 (O_699,N_4153,N_4697);
or UO_700 (O_700,N_4669,N_4165);
or UO_701 (O_701,N_4232,N_4638);
nor UO_702 (O_702,N_4031,N_4992);
and UO_703 (O_703,N_4135,N_4719);
or UO_704 (O_704,N_4972,N_4942);
and UO_705 (O_705,N_4333,N_4405);
nand UO_706 (O_706,N_4607,N_4973);
or UO_707 (O_707,N_4569,N_4219);
nand UO_708 (O_708,N_4612,N_4270);
nand UO_709 (O_709,N_4258,N_4409);
nor UO_710 (O_710,N_4069,N_4091);
nor UO_711 (O_711,N_4344,N_4593);
or UO_712 (O_712,N_4971,N_4202);
nor UO_713 (O_713,N_4877,N_4335);
or UO_714 (O_714,N_4904,N_4644);
or UO_715 (O_715,N_4857,N_4537);
nand UO_716 (O_716,N_4047,N_4716);
nand UO_717 (O_717,N_4012,N_4837);
nand UO_718 (O_718,N_4075,N_4846);
nor UO_719 (O_719,N_4660,N_4058);
nor UO_720 (O_720,N_4477,N_4676);
nor UO_721 (O_721,N_4462,N_4312);
or UO_722 (O_722,N_4392,N_4347);
nor UO_723 (O_723,N_4218,N_4940);
nand UO_724 (O_724,N_4672,N_4869);
or UO_725 (O_725,N_4982,N_4041);
and UO_726 (O_726,N_4166,N_4671);
or UO_727 (O_727,N_4913,N_4533);
nand UO_728 (O_728,N_4256,N_4486);
or UO_729 (O_729,N_4255,N_4368);
nor UO_730 (O_730,N_4405,N_4102);
and UO_731 (O_731,N_4317,N_4012);
xor UO_732 (O_732,N_4025,N_4581);
or UO_733 (O_733,N_4051,N_4683);
and UO_734 (O_734,N_4280,N_4654);
nand UO_735 (O_735,N_4008,N_4801);
and UO_736 (O_736,N_4154,N_4215);
nor UO_737 (O_737,N_4725,N_4373);
nand UO_738 (O_738,N_4316,N_4572);
or UO_739 (O_739,N_4149,N_4925);
or UO_740 (O_740,N_4741,N_4520);
nor UO_741 (O_741,N_4147,N_4680);
and UO_742 (O_742,N_4042,N_4851);
or UO_743 (O_743,N_4020,N_4751);
and UO_744 (O_744,N_4716,N_4952);
nor UO_745 (O_745,N_4582,N_4655);
or UO_746 (O_746,N_4953,N_4161);
and UO_747 (O_747,N_4100,N_4838);
nor UO_748 (O_748,N_4892,N_4647);
nand UO_749 (O_749,N_4786,N_4455);
and UO_750 (O_750,N_4174,N_4444);
nand UO_751 (O_751,N_4513,N_4279);
and UO_752 (O_752,N_4540,N_4323);
or UO_753 (O_753,N_4043,N_4912);
nor UO_754 (O_754,N_4292,N_4998);
and UO_755 (O_755,N_4233,N_4068);
nor UO_756 (O_756,N_4911,N_4280);
nor UO_757 (O_757,N_4995,N_4705);
nand UO_758 (O_758,N_4363,N_4565);
nand UO_759 (O_759,N_4698,N_4835);
or UO_760 (O_760,N_4508,N_4315);
nand UO_761 (O_761,N_4387,N_4432);
or UO_762 (O_762,N_4856,N_4387);
or UO_763 (O_763,N_4591,N_4135);
nor UO_764 (O_764,N_4493,N_4899);
or UO_765 (O_765,N_4570,N_4457);
and UO_766 (O_766,N_4927,N_4369);
nor UO_767 (O_767,N_4258,N_4066);
or UO_768 (O_768,N_4399,N_4496);
nor UO_769 (O_769,N_4839,N_4193);
nand UO_770 (O_770,N_4099,N_4507);
nor UO_771 (O_771,N_4525,N_4299);
nand UO_772 (O_772,N_4055,N_4722);
or UO_773 (O_773,N_4776,N_4920);
or UO_774 (O_774,N_4612,N_4345);
nor UO_775 (O_775,N_4246,N_4164);
nand UO_776 (O_776,N_4392,N_4057);
and UO_777 (O_777,N_4606,N_4372);
nor UO_778 (O_778,N_4096,N_4414);
nor UO_779 (O_779,N_4908,N_4227);
nor UO_780 (O_780,N_4696,N_4792);
or UO_781 (O_781,N_4161,N_4927);
nand UO_782 (O_782,N_4493,N_4465);
and UO_783 (O_783,N_4418,N_4236);
and UO_784 (O_784,N_4184,N_4543);
and UO_785 (O_785,N_4942,N_4632);
nor UO_786 (O_786,N_4300,N_4229);
nor UO_787 (O_787,N_4745,N_4189);
and UO_788 (O_788,N_4379,N_4219);
or UO_789 (O_789,N_4781,N_4288);
nor UO_790 (O_790,N_4200,N_4757);
or UO_791 (O_791,N_4702,N_4445);
nor UO_792 (O_792,N_4391,N_4847);
or UO_793 (O_793,N_4725,N_4321);
and UO_794 (O_794,N_4170,N_4215);
and UO_795 (O_795,N_4177,N_4157);
or UO_796 (O_796,N_4915,N_4225);
or UO_797 (O_797,N_4362,N_4361);
nand UO_798 (O_798,N_4400,N_4740);
nand UO_799 (O_799,N_4718,N_4519);
nand UO_800 (O_800,N_4517,N_4765);
nor UO_801 (O_801,N_4788,N_4122);
nand UO_802 (O_802,N_4676,N_4238);
nand UO_803 (O_803,N_4939,N_4828);
and UO_804 (O_804,N_4446,N_4077);
nand UO_805 (O_805,N_4012,N_4365);
and UO_806 (O_806,N_4410,N_4972);
and UO_807 (O_807,N_4049,N_4350);
or UO_808 (O_808,N_4380,N_4187);
or UO_809 (O_809,N_4146,N_4300);
nor UO_810 (O_810,N_4625,N_4319);
nor UO_811 (O_811,N_4806,N_4703);
and UO_812 (O_812,N_4466,N_4775);
nand UO_813 (O_813,N_4061,N_4632);
nor UO_814 (O_814,N_4347,N_4283);
nor UO_815 (O_815,N_4035,N_4530);
nor UO_816 (O_816,N_4430,N_4684);
or UO_817 (O_817,N_4601,N_4551);
nand UO_818 (O_818,N_4992,N_4900);
or UO_819 (O_819,N_4861,N_4849);
and UO_820 (O_820,N_4475,N_4169);
or UO_821 (O_821,N_4329,N_4474);
nand UO_822 (O_822,N_4806,N_4918);
nand UO_823 (O_823,N_4563,N_4888);
nand UO_824 (O_824,N_4063,N_4261);
nand UO_825 (O_825,N_4931,N_4703);
nor UO_826 (O_826,N_4157,N_4277);
nand UO_827 (O_827,N_4183,N_4169);
xnor UO_828 (O_828,N_4818,N_4861);
or UO_829 (O_829,N_4687,N_4593);
or UO_830 (O_830,N_4133,N_4203);
nor UO_831 (O_831,N_4168,N_4871);
and UO_832 (O_832,N_4619,N_4939);
or UO_833 (O_833,N_4601,N_4931);
and UO_834 (O_834,N_4689,N_4336);
nand UO_835 (O_835,N_4704,N_4153);
xor UO_836 (O_836,N_4391,N_4094);
or UO_837 (O_837,N_4070,N_4548);
and UO_838 (O_838,N_4777,N_4108);
or UO_839 (O_839,N_4541,N_4650);
or UO_840 (O_840,N_4322,N_4999);
and UO_841 (O_841,N_4242,N_4749);
or UO_842 (O_842,N_4732,N_4137);
nand UO_843 (O_843,N_4473,N_4276);
or UO_844 (O_844,N_4504,N_4683);
nand UO_845 (O_845,N_4573,N_4628);
nor UO_846 (O_846,N_4614,N_4310);
nand UO_847 (O_847,N_4077,N_4313);
or UO_848 (O_848,N_4451,N_4493);
nor UO_849 (O_849,N_4042,N_4271);
or UO_850 (O_850,N_4483,N_4349);
nand UO_851 (O_851,N_4970,N_4299);
nand UO_852 (O_852,N_4956,N_4032);
nor UO_853 (O_853,N_4456,N_4958);
nand UO_854 (O_854,N_4065,N_4974);
and UO_855 (O_855,N_4223,N_4650);
or UO_856 (O_856,N_4216,N_4969);
and UO_857 (O_857,N_4510,N_4582);
and UO_858 (O_858,N_4072,N_4493);
or UO_859 (O_859,N_4755,N_4678);
nor UO_860 (O_860,N_4169,N_4761);
nor UO_861 (O_861,N_4417,N_4937);
or UO_862 (O_862,N_4078,N_4325);
or UO_863 (O_863,N_4102,N_4840);
and UO_864 (O_864,N_4918,N_4629);
or UO_865 (O_865,N_4483,N_4700);
or UO_866 (O_866,N_4358,N_4222);
or UO_867 (O_867,N_4608,N_4315);
nand UO_868 (O_868,N_4059,N_4598);
or UO_869 (O_869,N_4714,N_4173);
or UO_870 (O_870,N_4530,N_4097);
nand UO_871 (O_871,N_4430,N_4947);
nor UO_872 (O_872,N_4373,N_4281);
or UO_873 (O_873,N_4171,N_4631);
nor UO_874 (O_874,N_4081,N_4165);
and UO_875 (O_875,N_4989,N_4799);
nor UO_876 (O_876,N_4056,N_4171);
nand UO_877 (O_877,N_4581,N_4295);
nor UO_878 (O_878,N_4755,N_4295);
nor UO_879 (O_879,N_4036,N_4276);
nand UO_880 (O_880,N_4234,N_4588);
nand UO_881 (O_881,N_4027,N_4302);
or UO_882 (O_882,N_4876,N_4851);
nor UO_883 (O_883,N_4888,N_4860);
and UO_884 (O_884,N_4823,N_4178);
or UO_885 (O_885,N_4118,N_4019);
or UO_886 (O_886,N_4949,N_4058);
nor UO_887 (O_887,N_4983,N_4324);
nand UO_888 (O_888,N_4566,N_4108);
and UO_889 (O_889,N_4049,N_4264);
and UO_890 (O_890,N_4164,N_4422);
and UO_891 (O_891,N_4378,N_4929);
nand UO_892 (O_892,N_4917,N_4852);
nand UO_893 (O_893,N_4868,N_4296);
or UO_894 (O_894,N_4350,N_4210);
and UO_895 (O_895,N_4075,N_4434);
nor UO_896 (O_896,N_4491,N_4185);
or UO_897 (O_897,N_4801,N_4835);
or UO_898 (O_898,N_4066,N_4024);
nand UO_899 (O_899,N_4380,N_4177);
nor UO_900 (O_900,N_4555,N_4091);
or UO_901 (O_901,N_4190,N_4331);
nor UO_902 (O_902,N_4895,N_4914);
nand UO_903 (O_903,N_4464,N_4084);
nand UO_904 (O_904,N_4992,N_4040);
nor UO_905 (O_905,N_4128,N_4992);
or UO_906 (O_906,N_4349,N_4695);
or UO_907 (O_907,N_4125,N_4048);
and UO_908 (O_908,N_4802,N_4826);
or UO_909 (O_909,N_4078,N_4600);
nor UO_910 (O_910,N_4207,N_4954);
or UO_911 (O_911,N_4543,N_4902);
and UO_912 (O_912,N_4272,N_4829);
or UO_913 (O_913,N_4945,N_4081);
nor UO_914 (O_914,N_4260,N_4575);
nand UO_915 (O_915,N_4128,N_4401);
xor UO_916 (O_916,N_4412,N_4696);
nand UO_917 (O_917,N_4136,N_4291);
nor UO_918 (O_918,N_4923,N_4732);
or UO_919 (O_919,N_4669,N_4014);
nand UO_920 (O_920,N_4991,N_4195);
nor UO_921 (O_921,N_4567,N_4405);
nand UO_922 (O_922,N_4433,N_4067);
nand UO_923 (O_923,N_4527,N_4382);
and UO_924 (O_924,N_4868,N_4171);
and UO_925 (O_925,N_4682,N_4899);
nor UO_926 (O_926,N_4845,N_4144);
nand UO_927 (O_927,N_4165,N_4740);
nand UO_928 (O_928,N_4346,N_4025);
nor UO_929 (O_929,N_4592,N_4758);
or UO_930 (O_930,N_4396,N_4081);
and UO_931 (O_931,N_4711,N_4929);
nand UO_932 (O_932,N_4894,N_4111);
or UO_933 (O_933,N_4298,N_4297);
nand UO_934 (O_934,N_4403,N_4110);
and UO_935 (O_935,N_4728,N_4561);
and UO_936 (O_936,N_4074,N_4825);
nand UO_937 (O_937,N_4427,N_4819);
or UO_938 (O_938,N_4346,N_4669);
or UO_939 (O_939,N_4062,N_4244);
or UO_940 (O_940,N_4750,N_4332);
and UO_941 (O_941,N_4355,N_4101);
nor UO_942 (O_942,N_4035,N_4794);
nand UO_943 (O_943,N_4285,N_4940);
and UO_944 (O_944,N_4649,N_4722);
or UO_945 (O_945,N_4543,N_4698);
or UO_946 (O_946,N_4225,N_4235);
or UO_947 (O_947,N_4471,N_4038);
or UO_948 (O_948,N_4919,N_4704);
and UO_949 (O_949,N_4344,N_4647);
or UO_950 (O_950,N_4810,N_4715);
nor UO_951 (O_951,N_4223,N_4959);
nor UO_952 (O_952,N_4438,N_4859);
nand UO_953 (O_953,N_4615,N_4888);
and UO_954 (O_954,N_4246,N_4241);
nand UO_955 (O_955,N_4822,N_4735);
or UO_956 (O_956,N_4563,N_4673);
nand UO_957 (O_957,N_4601,N_4051);
or UO_958 (O_958,N_4624,N_4591);
and UO_959 (O_959,N_4842,N_4527);
nor UO_960 (O_960,N_4964,N_4819);
and UO_961 (O_961,N_4940,N_4762);
or UO_962 (O_962,N_4574,N_4180);
nor UO_963 (O_963,N_4840,N_4576);
nand UO_964 (O_964,N_4334,N_4232);
nor UO_965 (O_965,N_4282,N_4393);
nor UO_966 (O_966,N_4249,N_4612);
nor UO_967 (O_967,N_4112,N_4883);
or UO_968 (O_968,N_4980,N_4239);
and UO_969 (O_969,N_4435,N_4536);
nor UO_970 (O_970,N_4438,N_4431);
or UO_971 (O_971,N_4415,N_4596);
and UO_972 (O_972,N_4799,N_4011);
nand UO_973 (O_973,N_4974,N_4750);
or UO_974 (O_974,N_4242,N_4957);
or UO_975 (O_975,N_4126,N_4420);
and UO_976 (O_976,N_4277,N_4391);
or UO_977 (O_977,N_4979,N_4548);
nor UO_978 (O_978,N_4889,N_4214);
or UO_979 (O_979,N_4576,N_4071);
or UO_980 (O_980,N_4745,N_4344);
nand UO_981 (O_981,N_4328,N_4561);
nor UO_982 (O_982,N_4664,N_4716);
and UO_983 (O_983,N_4450,N_4739);
nor UO_984 (O_984,N_4451,N_4098);
and UO_985 (O_985,N_4899,N_4869);
or UO_986 (O_986,N_4183,N_4194);
nand UO_987 (O_987,N_4044,N_4334);
nand UO_988 (O_988,N_4395,N_4059);
nand UO_989 (O_989,N_4356,N_4108);
nor UO_990 (O_990,N_4486,N_4858);
nand UO_991 (O_991,N_4159,N_4239);
nand UO_992 (O_992,N_4027,N_4610);
nor UO_993 (O_993,N_4280,N_4032);
and UO_994 (O_994,N_4955,N_4287);
and UO_995 (O_995,N_4422,N_4615);
nand UO_996 (O_996,N_4378,N_4293);
or UO_997 (O_997,N_4002,N_4410);
nor UO_998 (O_998,N_4159,N_4093);
nand UO_999 (O_999,N_4292,N_4725);
endmodule