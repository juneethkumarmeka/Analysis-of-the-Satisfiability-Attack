module basic_500_3000_500_50_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_384,In_176);
or U1 (N_1,In_434,In_157);
nor U2 (N_2,In_105,In_149);
nand U3 (N_3,In_293,In_302);
or U4 (N_4,In_50,In_440);
and U5 (N_5,In_306,In_197);
nand U6 (N_6,In_270,In_163);
nand U7 (N_7,In_261,In_195);
or U8 (N_8,In_295,In_439);
nand U9 (N_9,In_36,In_57);
nand U10 (N_10,In_314,In_449);
nand U11 (N_11,In_121,In_482);
nor U12 (N_12,In_430,In_154);
nand U13 (N_13,In_249,In_405);
or U14 (N_14,In_259,In_130);
nand U15 (N_15,In_235,In_373);
nor U16 (N_16,In_414,In_488);
nor U17 (N_17,In_422,In_43);
nor U18 (N_18,In_180,In_364);
nand U19 (N_19,In_355,In_55);
or U20 (N_20,In_416,In_174);
and U21 (N_21,In_369,In_64);
or U22 (N_22,In_146,In_320);
nor U23 (N_23,In_85,In_400);
or U24 (N_24,In_44,In_327);
or U25 (N_25,In_374,In_98);
nor U26 (N_26,In_183,In_429);
or U27 (N_27,In_478,In_11);
nand U28 (N_28,In_466,In_172);
and U29 (N_29,In_47,In_428);
nand U30 (N_30,In_204,In_145);
nand U31 (N_31,In_419,In_442);
xnor U32 (N_32,In_375,In_73);
nand U33 (N_33,In_14,In_467);
or U34 (N_34,In_95,In_451);
nor U35 (N_35,In_15,In_288);
nand U36 (N_36,In_240,In_18);
nor U37 (N_37,In_424,In_492);
and U38 (N_38,In_486,In_331);
nand U39 (N_39,In_378,In_371);
nor U40 (N_40,In_388,In_390);
nor U41 (N_41,In_443,In_99);
or U42 (N_42,In_418,In_411);
nand U43 (N_43,In_103,In_316);
or U44 (N_44,In_338,In_318);
and U45 (N_45,In_309,In_7);
nand U46 (N_46,In_382,In_412);
nor U47 (N_47,In_311,In_35);
nand U48 (N_48,In_462,In_269);
and U49 (N_49,In_305,In_361);
and U50 (N_50,In_366,In_358);
nand U51 (N_51,In_193,In_106);
nor U52 (N_52,In_243,In_395);
or U53 (N_53,In_170,In_403);
or U54 (N_54,In_137,In_83);
and U55 (N_55,In_3,In_209);
nor U56 (N_56,In_232,In_112);
nand U57 (N_57,In_100,In_75);
nand U58 (N_58,In_194,In_463);
and U59 (N_59,In_92,In_168);
and U60 (N_60,In_426,In_201);
nand U61 (N_61,In_188,In_237);
and U62 (N_62,In_228,In_433);
nor U63 (N_63,In_359,In_25);
and U64 (N_64,In_281,In_367);
nor U65 (N_65,In_167,N_10);
xor U66 (N_66,In_377,In_16);
or U67 (N_67,In_475,In_271);
xnor U68 (N_68,In_333,In_141);
nor U69 (N_69,In_284,In_315);
nor U70 (N_70,In_385,In_186);
and U71 (N_71,In_33,N_55);
nor U72 (N_72,In_253,In_287);
nand U73 (N_73,In_241,In_152);
nand U74 (N_74,In_88,In_54);
and U75 (N_75,N_58,N_2);
nor U76 (N_76,N_26,In_238);
or U77 (N_77,In_150,In_122);
and U78 (N_78,In_415,In_89);
or U79 (N_79,In_187,In_289);
xor U80 (N_80,N_12,In_109);
or U81 (N_81,In_234,N_34);
nand U82 (N_82,N_15,In_436);
or U83 (N_83,In_67,In_323);
xor U84 (N_84,In_211,In_431);
and U85 (N_85,In_53,In_410);
or U86 (N_86,In_450,In_252);
nand U87 (N_87,In_372,In_79);
nor U88 (N_88,In_370,In_340);
nand U89 (N_89,In_404,In_493);
nor U90 (N_90,In_86,In_386);
nor U91 (N_91,In_296,N_56);
nor U92 (N_92,N_27,In_107);
or U93 (N_93,In_23,In_266);
nand U94 (N_94,In_126,In_401);
or U95 (N_95,In_68,N_21);
or U96 (N_96,N_39,In_90);
nor U97 (N_97,In_267,In_205);
or U98 (N_98,In_13,In_184);
and U99 (N_99,In_268,In_94);
and U100 (N_100,In_448,In_460);
or U101 (N_101,In_217,In_59);
nand U102 (N_102,In_353,In_477);
xnor U103 (N_103,In_37,In_185);
xnor U104 (N_104,In_138,In_265);
nor U105 (N_105,In_343,In_39);
or U106 (N_106,In_147,In_165);
nand U107 (N_107,In_402,N_24);
or U108 (N_108,N_29,In_489);
nand U109 (N_109,In_227,In_461);
nand U110 (N_110,In_274,N_32);
nor U111 (N_111,N_52,N_40);
and U112 (N_112,In_283,In_84);
and U113 (N_113,N_49,In_273);
nand U114 (N_114,N_16,In_61);
and U115 (N_115,In_58,In_104);
nand U116 (N_116,In_496,In_4);
or U117 (N_117,In_423,In_111);
and U118 (N_118,In_465,In_41);
and U119 (N_119,In_81,In_455);
and U120 (N_120,In_459,In_363);
xnor U121 (N_121,N_114,In_304);
and U122 (N_122,In_71,In_139);
nor U123 (N_123,N_37,In_135);
or U124 (N_124,In_479,In_297);
and U125 (N_125,In_480,In_239);
nand U126 (N_126,In_116,In_263);
or U127 (N_127,In_198,N_50);
nor U128 (N_128,In_159,N_117);
xnor U129 (N_129,In_226,In_381);
and U130 (N_130,In_133,N_76);
and U131 (N_131,In_409,In_328);
or U132 (N_132,N_47,N_73);
xor U133 (N_133,N_66,In_65);
nor U134 (N_134,In_233,In_387);
or U135 (N_135,In_317,In_12);
nand U136 (N_136,In_245,N_81);
or U137 (N_137,N_18,In_421);
nand U138 (N_138,In_352,In_24);
nand U139 (N_139,N_51,In_5);
nand U140 (N_140,In_335,In_291);
nor U141 (N_141,N_23,In_120);
nor U142 (N_142,In_148,In_321);
nand U143 (N_143,In_202,In_34);
xnor U144 (N_144,In_380,N_100);
or U145 (N_145,In_322,N_89);
nand U146 (N_146,N_86,In_66);
nand U147 (N_147,In_319,In_360);
and U148 (N_148,In_379,N_80);
or U149 (N_149,N_68,In_128);
and U150 (N_150,N_99,In_212);
and U151 (N_151,In_332,N_91);
nand U152 (N_152,In_21,In_230);
nand U153 (N_153,In_119,In_491);
and U154 (N_154,N_35,In_307);
and U155 (N_155,In_236,N_118);
or U156 (N_156,N_43,In_22);
nand U157 (N_157,In_203,In_495);
or U158 (N_158,In_487,In_474);
or U159 (N_159,In_101,In_312);
nand U160 (N_160,N_103,In_300);
nor U161 (N_161,In_27,In_473);
or U162 (N_162,In_215,N_110);
nor U163 (N_163,N_70,In_278);
nand U164 (N_164,In_470,In_216);
nor U165 (N_165,In_69,N_42);
nor U166 (N_166,In_52,N_61);
nor U167 (N_167,N_92,In_394);
xnor U168 (N_168,In_51,In_324);
nand U169 (N_169,In_452,N_106);
or U170 (N_170,In_30,N_77);
nor U171 (N_171,N_22,In_357);
and U172 (N_172,In_399,N_9);
or U173 (N_173,N_5,In_191);
and U174 (N_174,In_80,In_339);
xor U175 (N_175,In_337,N_116);
nor U176 (N_176,In_348,In_303);
xnor U177 (N_177,N_14,In_254);
nand U178 (N_178,N_104,In_264);
nand U179 (N_179,N_1,In_351);
nor U180 (N_180,In_77,In_349);
and U181 (N_181,In_161,In_8);
and U182 (N_182,N_149,In_93);
and U183 (N_183,In_250,N_126);
nand U184 (N_184,N_48,In_444);
nor U185 (N_185,In_142,In_389);
nand U186 (N_186,In_26,In_483);
or U187 (N_187,In_279,In_498);
or U188 (N_188,In_290,N_101);
or U189 (N_189,N_65,N_83);
nand U190 (N_190,In_272,In_169);
xnor U191 (N_191,N_107,In_2);
or U192 (N_192,In_464,In_155);
and U193 (N_193,N_0,In_118);
nand U194 (N_194,In_256,In_425);
or U195 (N_195,N_125,In_334);
or U196 (N_196,N_148,N_123);
or U197 (N_197,In_115,N_168);
nor U198 (N_198,In_74,In_246);
nor U199 (N_199,N_45,N_62);
nor U200 (N_200,In_49,In_143);
and U201 (N_201,In_456,N_129);
nand U202 (N_202,N_140,In_432);
and U203 (N_203,N_7,In_407);
nand U204 (N_204,N_28,In_255);
nand U205 (N_205,In_481,N_130);
xnor U206 (N_206,In_28,In_91);
nor U207 (N_207,In_247,N_115);
or U208 (N_208,In_9,N_108);
nor U209 (N_209,N_175,In_285);
xor U210 (N_210,In_244,In_454);
and U211 (N_211,In_63,N_36);
nor U212 (N_212,N_138,In_262);
and U213 (N_213,N_142,In_383);
nand U214 (N_214,N_84,N_147);
nand U215 (N_215,N_128,In_397);
nand U216 (N_216,In_189,In_179);
or U217 (N_217,N_6,N_44);
or U218 (N_218,In_392,N_78);
and U219 (N_219,In_354,In_220);
nand U220 (N_220,In_110,In_6);
nor U221 (N_221,N_85,In_218);
or U222 (N_222,In_10,N_173);
and U223 (N_223,In_391,N_137);
and U224 (N_224,In_362,N_141);
and U225 (N_225,N_167,N_174);
nand U226 (N_226,In_131,In_132);
or U227 (N_227,In_282,In_207);
or U228 (N_228,In_175,In_260);
and U229 (N_229,In_472,N_53);
nand U230 (N_230,In_102,N_46);
and U231 (N_231,N_8,In_485);
nor U232 (N_232,In_347,N_67);
and U233 (N_233,In_484,In_341);
or U234 (N_234,In_342,In_457);
nor U235 (N_235,In_1,N_60);
and U236 (N_236,In_231,In_277);
xnor U237 (N_237,In_129,In_82);
nand U238 (N_238,In_376,In_393);
or U239 (N_239,N_166,N_169);
xnor U240 (N_240,N_127,In_219);
nor U241 (N_241,N_231,In_144);
nand U242 (N_242,N_192,N_178);
nor U243 (N_243,In_301,N_162);
nor U244 (N_244,N_233,In_329);
nand U245 (N_245,In_298,N_201);
nor U246 (N_246,N_79,In_427);
nor U247 (N_247,In_286,N_145);
nor U248 (N_248,In_458,N_194);
nand U249 (N_249,In_221,In_294);
nor U250 (N_250,In_471,In_206);
nand U251 (N_251,In_114,In_313);
and U252 (N_252,In_134,In_446);
or U253 (N_253,In_40,In_224);
nand U254 (N_254,N_236,In_97);
nand U255 (N_255,N_11,N_163);
xnor U256 (N_256,N_144,In_42);
and U257 (N_257,N_181,N_202);
nand U258 (N_258,In_345,In_417);
xnor U259 (N_259,In_257,In_45);
or U260 (N_260,N_209,In_166);
nor U261 (N_261,N_139,N_218);
xnor U262 (N_262,N_204,In_160);
nand U263 (N_263,In_72,N_120);
nand U264 (N_264,In_17,In_76);
and U265 (N_265,In_70,N_30);
xnor U266 (N_266,N_184,In_31);
or U267 (N_267,In_60,N_186);
or U268 (N_268,In_229,N_97);
and U269 (N_269,N_211,N_13);
or U270 (N_270,N_25,In_453);
nor U271 (N_271,N_221,N_112);
or U272 (N_272,N_87,N_180);
and U273 (N_273,In_136,In_182);
xor U274 (N_274,N_220,In_248);
nor U275 (N_275,In_213,N_216);
and U276 (N_276,N_237,N_226);
nand U277 (N_277,N_111,N_224);
nor U278 (N_278,N_96,N_219);
or U279 (N_279,N_74,In_164);
nand U280 (N_280,In_398,N_187);
and U281 (N_281,N_239,N_195);
nor U282 (N_282,N_205,In_29);
xor U283 (N_283,In_275,N_132);
or U284 (N_284,N_227,N_33);
or U285 (N_285,In_435,In_96);
nand U286 (N_286,In_336,In_325);
nor U287 (N_287,In_344,N_172);
nor U288 (N_288,N_94,N_71);
nor U289 (N_289,N_238,N_88);
nor U290 (N_290,In_396,N_152);
nand U291 (N_291,In_210,N_133);
or U292 (N_292,N_232,In_140);
and U293 (N_293,In_192,N_157);
nand U294 (N_294,N_213,In_171);
and U295 (N_295,In_78,In_199);
or U296 (N_296,N_161,In_153);
and U297 (N_297,In_124,In_308);
nor U298 (N_298,In_178,In_330);
nor U299 (N_299,N_191,N_164);
or U300 (N_300,N_82,N_292);
or U301 (N_301,N_159,In_127);
and U302 (N_302,In_20,N_93);
nor U303 (N_303,N_280,In_32);
xnor U304 (N_304,N_284,N_296);
and U305 (N_305,N_196,In_38);
or U306 (N_306,N_252,In_469);
and U307 (N_307,N_295,N_143);
and U308 (N_308,N_247,N_261);
nand U309 (N_309,N_158,N_54);
nor U310 (N_310,N_135,N_156);
nand U311 (N_311,In_490,N_95);
nor U312 (N_312,N_283,N_241);
xnor U313 (N_313,In_225,In_177);
or U314 (N_314,N_153,N_64);
nand U315 (N_315,N_256,N_240);
nor U316 (N_316,In_497,N_249);
nor U317 (N_317,N_207,In_299);
and U318 (N_318,N_257,N_229);
and U319 (N_319,In_468,In_356);
or U320 (N_320,N_20,In_222);
xnor U321 (N_321,N_271,N_206);
nor U322 (N_322,N_113,In_413);
xnor U323 (N_323,N_259,N_151);
nand U324 (N_324,In_46,In_350);
nand U325 (N_325,N_75,N_109);
nor U326 (N_326,N_299,N_246);
and U327 (N_327,N_260,N_131);
or U328 (N_328,N_146,N_189);
nor U329 (N_329,N_276,N_136);
xnor U330 (N_330,In_445,N_182);
and U331 (N_331,N_179,In_406);
or U332 (N_332,N_263,N_177);
or U333 (N_333,N_171,N_274);
or U334 (N_334,N_121,N_254);
xnor U335 (N_335,In_365,N_217);
nand U336 (N_336,N_98,N_294);
nor U337 (N_337,N_160,N_275);
nor U338 (N_338,N_31,In_113);
or U339 (N_339,In_156,N_230);
nand U340 (N_340,N_264,N_199);
xnor U341 (N_341,N_228,N_63);
nand U342 (N_342,N_102,N_253);
or U343 (N_343,In_420,In_173);
nand U344 (N_344,In_208,In_158);
or U345 (N_345,N_203,In_196);
or U346 (N_346,In_499,N_208);
or U347 (N_347,In_242,N_223);
and U348 (N_348,In_190,N_270);
nor U349 (N_349,N_290,N_287);
nor U350 (N_350,In_441,N_278);
or U351 (N_351,N_277,N_289);
nand U352 (N_352,In_223,In_62);
nand U353 (N_353,In_258,N_105);
nand U354 (N_354,In_214,N_212);
or U355 (N_355,N_248,N_69);
and U356 (N_356,N_124,N_197);
nand U357 (N_357,In_276,In_476);
or U358 (N_358,In_125,N_183);
nor U359 (N_359,In_108,N_210);
nor U360 (N_360,N_335,In_200);
and U361 (N_361,N_341,N_258);
and U362 (N_362,N_293,N_298);
xor U363 (N_363,N_269,N_332);
nand U364 (N_364,In_438,N_337);
nand U365 (N_365,N_349,N_119);
and U366 (N_366,N_286,N_265);
nand U367 (N_367,N_321,N_198);
nor U368 (N_368,N_155,N_3);
or U369 (N_369,N_327,In_151);
nand U370 (N_370,N_57,In_56);
or U371 (N_371,N_329,N_312);
nor U372 (N_372,N_328,N_316);
nor U373 (N_373,N_326,N_225);
nand U374 (N_374,In_19,N_324);
or U375 (N_375,N_242,In_494);
nor U376 (N_376,N_185,N_268);
or U377 (N_377,N_250,N_193);
nand U378 (N_378,N_317,N_338);
and U379 (N_379,N_303,In_326);
nand U380 (N_380,N_354,N_334);
and U381 (N_381,N_336,N_262);
or U382 (N_382,In_87,N_4);
nor U383 (N_383,N_319,N_214);
nand U384 (N_384,In_408,N_188);
nand U385 (N_385,N_281,N_251);
and U386 (N_386,N_320,N_314);
nand U387 (N_387,N_355,N_304);
or U388 (N_388,In_310,N_134);
xor U389 (N_389,N_285,N_235);
and U390 (N_390,N_346,N_342);
or U391 (N_391,N_200,N_351);
and U392 (N_392,N_308,N_288);
or U393 (N_393,N_345,N_301);
nor U394 (N_394,N_356,In_0);
or U395 (N_395,In_346,N_17);
nand U396 (N_396,N_300,In_251);
or U397 (N_397,N_273,N_234);
and U398 (N_398,N_309,In_162);
or U399 (N_399,N_176,N_72);
and U400 (N_400,N_302,N_306);
nand U401 (N_401,N_244,In_447);
nand U402 (N_402,N_313,N_297);
nand U403 (N_403,N_311,N_344);
and U404 (N_404,N_330,N_272);
or U405 (N_405,N_291,N_267);
nor U406 (N_406,N_245,N_307);
nor U407 (N_407,In_117,N_279);
nor U408 (N_408,N_190,In_368);
nor U409 (N_409,In_48,N_310);
nor U410 (N_410,N_357,N_215);
or U411 (N_411,N_266,N_150);
nand U412 (N_412,N_325,N_170);
nor U413 (N_413,N_315,N_122);
or U414 (N_414,N_348,N_19);
and U415 (N_415,In_280,N_243);
and U416 (N_416,N_154,In_181);
and U417 (N_417,N_305,In_292);
nand U418 (N_418,In_123,N_340);
nand U419 (N_419,N_255,N_322);
nor U420 (N_420,N_412,N_418);
and U421 (N_421,N_379,N_391);
nor U422 (N_422,N_374,N_395);
xnor U423 (N_423,N_339,N_366);
nor U424 (N_424,N_403,N_397);
or U425 (N_425,N_387,N_407);
and U426 (N_426,N_333,N_390);
nor U427 (N_427,N_361,N_222);
nand U428 (N_428,N_417,N_392);
or U429 (N_429,N_409,N_377);
nor U430 (N_430,N_415,N_370);
or U431 (N_431,N_389,N_347);
or U432 (N_432,N_380,N_358);
nor U433 (N_433,N_410,N_394);
or U434 (N_434,N_419,N_401);
and U435 (N_435,N_352,In_437);
and U436 (N_436,N_38,N_386);
and U437 (N_437,N_388,N_406);
nor U438 (N_438,N_383,N_331);
nor U439 (N_439,N_402,N_398);
nor U440 (N_440,N_375,N_371);
nand U441 (N_441,N_384,N_59);
and U442 (N_442,N_343,N_90);
or U443 (N_443,N_396,N_360);
nor U444 (N_444,N_365,N_414);
nor U445 (N_445,N_359,N_363);
or U446 (N_446,N_385,N_350);
nor U447 (N_447,N_368,N_41);
nor U448 (N_448,N_405,N_282);
and U449 (N_449,N_378,N_373);
nand U450 (N_450,N_165,N_408);
or U451 (N_451,N_416,N_393);
nor U452 (N_452,N_411,N_382);
nor U453 (N_453,N_364,N_400);
nor U454 (N_454,N_362,N_353);
and U455 (N_455,N_372,N_381);
or U456 (N_456,N_413,N_323);
nand U457 (N_457,N_376,N_369);
nor U458 (N_458,N_318,N_404);
and U459 (N_459,N_399,N_367);
and U460 (N_460,N_411,N_401);
nand U461 (N_461,N_282,N_372);
and U462 (N_462,N_382,N_417);
or U463 (N_463,N_333,N_405);
nand U464 (N_464,N_371,N_410);
or U465 (N_465,N_365,N_390);
or U466 (N_466,N_347,N_413);
nand U467 (N_467,N_59,N_392);
nand U468 (N_468,N_384,N_343);
nor U469 (N_469,N_391,N_41);
nor U470 (N_470,N_415,N_360);
nor U471 (N_471,N_382,N_363);
or U472 (N_472,N_367,N_318);
or U473 (N_473,N_399,N_403);
nor U474 (N_474,N_379,N_396);
and U475 (N_475,N_372,N_382);
and U476 (N_476,N_380,N_365);
xor U477 (N_477,N_396,N_419);
nor U478 (N_478,N_407,N_404);
nor U479 (N_479,N_395,N_381);
nand U480 (N_480,N_443,N_435);
nor U481 (N_481,N_444,N_437);
nor U482 (N_482,N_427,N_454);
nor U483 (N_483,N_434,N_457);
nor U484 (N_484,N_425,N_421);
nor U485 (N_485,N_440,N_433);
and U486 (N_486,N_459,N_448);
and U487 (N_487,N_447,N_436);
or U488 (N_488,N_450,N_478);
or U489 (N_489,N_471,N_423);
nand U490 (N_490,N_474,N_476);
nand U491 (N_491,N_479,N_467);
and U492 (N_492,N_432,N_461);
nor U493 (N_493,N_422,N_446);
xor U494 (N_494,N_473,N_428);
and U495 (N_495,N_477,N_426);
nor U496 (N_496,N_441,N_468);
and U497 (N_497,N_438,N_460);
and U498 (N_498,N_470,N_464);
xnor U499 (N_499,N_451,N_456);
nor U500 (N_500,N_431,N_469);
nor U501 (N_501,N_462,N_458);
and U502 (N_502,N_430,N_465);
and U503 (N_503,N_472,N_424);
or U504 (N_504,N_466,N_452);
or U505 (N_505,N_453,N_455);
xnor U506 (N_506,N_442,N_449);
and U507 (N_507,N_463,N_475);
nand U508 (N_508,N_420,N_445);
xor U509 (N_509,N_439,N_429);
nor U510 (N_510,N_456,N_467);
or U511 (N_511,N_424,N_441);
nand U512 (N_512,N_445,N_431);
and U513 (N_513,N_420,N_429);
nand U514 (N_514,N_442,N_471);
nand U515 (N_515,N_430,N_474);
nor U516 (N_516,N_450,N_427);
nor U517 (N_517,N_432,N_440);
nand U518 (N_518,N_476,N_460);
nor U519 (N_519,N_450,N_430);
nand U520 (N_520,N_475,N_443);
nor U521 (N_521,N_426,N_475);
nand U522 (N_522,N_423,N_450);
or U523 (N_523,N_423,N_420);
and U524 (N_524,N_479,N_451);
or U525 (N_525,N_433,N_458);
nand U526 (N_526,N_473,N_449);
nand U527 (N_527,N_446,N_437);
or U528 (N_528,N_437,N_467);
and U529 (N_529,N_472,N_452);
and U530 (N_530,N_479,N_429);
nor U531 (N_531,N_434,N_459);
nor U532 (N_532,N_466,N_451);
nand U533 (N_533,N_424,N_430);
nand U534 (N_534,N_463,N_467);
or U535 (N_535,N_446,N_477);
or U536 (N_536,N_459,N_479);
and U537 (N_537,N_472,N_440);
nand U538 (N_538,N_453,N_461);
and U539 (N_539,N_427,N_477);
xor U540 (N_540,N_489,N_534);
or U541 (N_541,N_508,N_536);
nand U542 (N_542,N_529,N_491);
nand U543 (N_543,N_490,N_496);
or U544 (N_544,N_525,N_537);
nor U545 (N_545,N_500,N_486);
nand U546 (N_546,N_485,N_521);
nor U547 (N_547,N_480,N_502);
nor U548 (N_548,N_524,N_519);
nand U549 (N_549,N_531,N_511);
xnor U550 (N_550,N_481,N_518);
nor U551 (N_551,N_495,N_539);
or U552 (N_552,N_522,N_513);
nor U553 (N_553,N_527,N_497);
nand U554 (N_554,N_493,N_492);
or U555 (N_555,N_505,N_499);
xnor U556 (N_556,N_516,N_520);
and U557 (N_557,N_510,N_498);
and U558 (N_558,N_530,N_514);
nand U559 (N_559,N_517,N_512);
xor U560 (N_560,N_506,N_528);
nand U561 (N_561,N_535,N_504);
or U562 (N_562,N_532,N_482);
or U563 (N_563,N_487,N_509);
nor U564 (N_564,N_507,N_538);
and U565 (N_565,N_501,N_483);
nor U566 (N_566,N_523,N_488);
and U567 (N_567,N_526,N_503);
or U568 (N_568,N_484,N_494);
nand U569 (N_569,N_515,N_533);
xor U570 (N_570,N_518,N_520);
or U571 (N_571,N_504,N_526);
nand U572 (N_572,N_498,N_504);
or U573 (N_573,N_512,N_534);
or U574 (N_574,N_499,N_487);
xnor U575 (N_575,N_536,N_539);
xnor U576 (N_576,N_539,N_490);
nor U577 (N_577,N_517,N_494);
xnor U578 (N_578,N_499,N_535);
nor U579 (N_579,N_516,N_501);
nand U580 (N_580,N_533,N_531);
or U581 (N_581,N_515,N_502);
nor U582 (N_582,N_538,N_509);
nor U583 (N_583,N_529,N_503);
or U584 (N_584,N_504,N_488);
nor U585 (N_585,N_489,N_506);
and U586 (N_586,N_506,N_521);
or U587 (N_587,N_514,N_499);
xnor U588 (N_588,N_480,N_535);
or U589 (N_589,N_508,N_487);
or U590 (N_590,N_535,N_505);
xnor U591 (N_591,N_539,N_513);
nor U592 (N_592,N_482,N_517);
nor U593 (N_593,N_480,N_506);
and U594 (N_594,N_529,N_486);
nor U595 (N_595,N_493,N_519);
nand U596 (N_596,N_516,N_534);
or U597 (N_597,N_510,N_526);
nor U598 (N_598,N_513,N_530);
or U599 (N_599,N_531,N_485);
nor U600 (N_600,N_548,N_592);
or U601 (N_601,N_562,N_566);
nor U602 (N_602,N_578,N_541);
nand U603 (N_603,N_586,N_550);
nor U604 (N_604,N_554,N_549);
nor U605 (N_605,N_573,N_588);
nand U606 (N_606,N_553,N_579);
nor U607 (N_607,N_564,N_552);
or U608 (N_608,N_572,N_565);
nor U609 (N_609,N_546,N_577);
nor U610 (N_610,N_580,N_598);
nand U611 (N_611,N_574,N_567);
nand U612 (N_612,N_563,N_593);
or U613 (N_613,N_583,N_571);
or U614 (N_614,N_575,N_544);
nand U615 (N_615,N_587,N_540);
nand U616 (N_616,N_596,N_590);
and U617 (N_617,N_556,N_594);
or U618 (N_618,N_595,N_576);
and U619 (N_619,N_584,N_561);
nand U620 (N_620,N_560,N_545);
or U621 (N_621,N_597,N_557);
or U622 (N_622,N_589,N_599);
and U623 (N_623,N_570,N_558);
nand U624 (N_624,N_542,N_582);
nor U625 (N_625,N_585,N_547);
nand U626 (N_626,N_591,N_551);
or U627 (N_627,N_555,N_559);
nor U628 (N_628,N_569,N_543);
nor U629 (N_629,N_581,N_568);
and U630 (N_630,N_562,N_580);
nor U631 (N_631,N_557,N_547);
or U632 (N_632,N_554,N_589);
xnor U633 (N_633,N_565,N_568);
nor U634 (N_634,N_591,N_569);
nand U635 (N_635,N_555,N_551);
or U636 (N_636,N_588,N_592);
nor U637 (N_637,N_550,N_592);
or U638 (N_638,N_591,N_552);
and U639 (N_639,N_564,N_568);
and U640 (N_640,N_574,N_571);
nand U641 (N_641,N_571,N_560);
or U642 (N_642,N_577,N_579);
xor U643 (N_643,N_583,N_575);
nor U644 (N_644,N_575,N_540);
nand U645 (N_645,N_575,N_560);
or U646 (N_646,N_558,N_589);
nor U647 (N_647,N_585,N_574);
nand U648 (N_648,N_597,N_542);
xnor U649 (N_649,N_579,N_559);
nand U650 (N_650,N_544,N_565);
nand U651 (N_651,N_554,N_551);
and U652 (N_652,N_582,N_552);
nor U653 (N_653,N_588,N_549);
nor U654 (N_654,N_545,N_590);
nor U655 (N_655,N_582,N_595);
xnor U656 (N_656,N_585,N_586);
xor U657 (N_657,N_568,N_544);
or U658 (N_658,N_555,N_552);
or U659 (N_659,N_599,N_581);
nor U660 (N_660,N_621,N_610);
nor U661 (N_661,N_607,N_613);
xor U662 (N_662,N_641,N_653);
xnor U663 (N_663,N_604,N_616);
nor U664 (N_664,N_626,N_654);
nand U665 (N_665,N_609,N_634);
or U666 (N_666,N_605,N_622);
or U667 (N_667,N_656,N_658);
nor U668 (N_668,N_617,N_643);
nand U669 (N_669,N_648,N_618);
nor U670 (N_670,N_600,N_639);
or U671 (N_671,N_611,N_633);
nand U672 (N_672,N_614,N_603);
xor U673 (N_673,N_608,N_637);
nand U674 (N_674,N_612,N_652);
or U675 (N_675,N_647,N_650);
nand U676 (N_676,N_624,N_635);
or U677 (N_677,N_651,N_620);
or U678 (N_678,N_628,N_644);
nor U679 (N_679,N_645,N_623);
and U680 (N_680,N_627,N_629);
and U681 (N_681,N_642,N_625);
or U682 (N_682,N_640,N_632);
nand U683 (N_683,N_638,N_615);
nand U684 (N_684,N_606,N_636);
and U685 (N_685,N_602,N_601);
and U686 (N_686,N_619,N_657);
nor U687 (N_687,N_655,N_631);
and U688 (N_688,N_646,N_630);
and U689 (N_689,N_659,N_649);
nand U690 (N_690,N_627,N_602);
nand U691 (N_691,N_635,N_620);
nand U692 (N_692,N_615,N_647);
nand U693 (N_693,N_607,N_657);
nand U694 (N_694,N_651,N_609);
xnor U695 (N_695,N_649,N_607);
nor U696 (N_696,N_612,N_637);
or U697 (N_697,N_635,N_605);
xor U698 (N_698,N_637,N_629);
nor U699 (N_699,N_627,N_649);
nand U700 (N_700,N_656,N_603);
nor U701 (N_701,N_610,N_604);
nor U702 (N_702,N_645,N_616);
nor U703 (N_703,N_609,N_631);
xor U704 (N_704,N_645,N_624);
and U705 (N_705,N_613,N_614);
and U706 (N_706,N_649,N_639);
nor U707 (N_707,N_650,N_637);
nand U708 (N_708,N_657,N_646);
or U709 (N_709,N_649,N_646);
nand U710 (N_710,N_631,N_658);
nor U711 (N_711,N_634,N_644);
and U712 (N_712,N_649,N_624);
nor U713 (N_713,N_630,N_612);
nor U714 (N_714,N_653,N_645);
nor U715 (N_715,N_657,N_649);
nor U716 (N_716,N_658,N_657);
nor U717 (N_717,N_623,N_636);
and U718 (N_718,N_644,N_615);
and U719 (N_719,N_620,N_608);
or U720 (N_720,N_668,N_718);
and U721 (N_721,N_688,N_673);
and U722 (N_722,N_686,N_666);
and U723 (N_723,N_667,N_710);
or U724 (N_724,N_696,N_700);
and U725 (N_725,N_712,N_682);
nor U726 (N_726,N_683,N_691);
xor U727 (N_727,N_664,N_672);
or U728 (N_728,N_661,N_678);
and U729 (N_729,N_684,N_717);
nand U730 (N_730,N_714,N_709);
and U731 (N_731,N_670,N_719);
and U732 (N_732,N_705,N_677);
nand U733 (N_733,N_690,N_698);
nor U734 (N_734,N_697,N_703);
xnor U735 (N_735,N_675,N_704);
and U736 (N_736,N_687,N_701);
or U737 (N_737,N_663,N_695);
nor U738 (N_738,N_676,N_660);
nor U739 (N_739,N_711,N_685);
nand U740 (N_740,N_716,N_713);
and U741 (N_741,N_707,N_694);
and U742 (N_742,N_665,N_671);
and U743 (N_743,N_706,N_715);
xnor U744 (N_744,N_662,N_708);
nand U745 (N_745,N_693,N_680);
nor U746 (N_746,N_674,N_669);
xor U747 (N_747,N_689,N_699);
and U748 (N_748,N_692,N_679);
or U749 (N_749,N_681,N_702);
or U750 (N_750,N_661,N_679);
nand U751 (N_751,N_682,N_660);
xor U752 (N_752,N_695,N_708);
xor U753 (N_753,N_670,N_693);
and U754 (N_754,N_673,N_718);
or U755 (N_755,N_689,N_668);
and U756 (N_756,N_692,N_663);
nand U757 (N_757,N_661,N_677);
xor U758 (N_758,N_670,N_678);
or U759 (N_759,N_701,N_700);
and U760 (N_760,N_706,N_688);
nand U761 (N_761,N_670,N_666);
or U762 (N_762,N_708,N_699);
nand U763 (N_763,N_660,N_714);
or U764 (N_764,N_661,N_660);
nor U765 (N_765,N_682,N_695);
nand U766 (N_766,N_688,N_709);
or U767 (N_767,N_678,N_702);
nor U768 (N_768,N_700,N_681);
nor U769 (N_769,N_676,N_692);
xnor U770 (N_770,N_680,N_701);
nor U771 (N_771,N_696,N_690);
nand U772 (N_772,N_694,N_712);
or U773 (N_773,N_700,N_679);
nand U774 (N_774,N_716,N_699);
nor U775 (N_775,N_699,N_707);
nor U776 (N_776,N_694,N_710);
and U777 (N_777,N_678,N_684);
and U778 (N_778,N_714,N_710);
nor U779 (N_779,N_705,N_666);
or U780 (N_780,N_722,N_755);
xnor U781 (N_781,N_749,N_739);
nand U782 (N_782,N_775,N_753);
and U783 (N_783,N_730,N_774);
or U784 (N_784,N_738,N_769);
or U785 (N_785,N_724,N_732);
and U786 (N_786,N_761,N_766);
nor U787 (N_787,N_728,N_771);
nor U788 (N_788,N_751,N_733);
xor U789 (N_789,N_744,N_748);
nor U790 (N_790,N_721,N_762);
nor U791 (N_791,N_745,N_760);
nand U792 (N_792,N_768,N_747);
xnor U793 (N_793,N_756,N_742);
nand U794 (N_794,N_723,N_776);
and U795 (N_795,N_737,N_754);
xor U796 (N_796,N_736,N_779);
and U797 (N_797,N_720,N_759);
nor U798 (N_798,N_767,N_726);
xor U799 (N_799,N_725,N_778);
nand U800 (N_800,N_750,N_757);
nand U801 (N_801,N_777,N_743);
nand U802 (N_802,N_752,N_740);
nand U803 (N_803,N_731,N_763);
nor U804 (N_804,N_741,N_770);
and U805 (N_805,N_764,N_734);
nand U806 (N_806,N_735,N_772);
nand U807 (N_807,N_746,N_729);
and U808 (N_808,N_727,N_773);
and U809 (N_809,N_765,N_758);
xor U810 (N_810,N_727,N_742);
nor U811 (N_811,N_745,N_764);
xnor U812 (N_812,N_738,N_749);
and U813 (N_813,N_724,N_761);
xnor U814 (N_814,N_750,N_772);
and U815 (N_815,N_748,N_727);
or U816 (N_816,N_751,N_727);
and U817 (N_817,N_761,N_725);
nand U818 (N_818,N_779,N_757);
or U819 (N_819,N_762,N_739);
nor U820 (N_820,N_772,N_770);
or U821 (N_821,N_775,N_727);
or U822 (N_822,N_755,N_758);
or U823 (N_823,N_772,N_747);
or U824 (N_824,N_752,N_753);
or U825 (N_825,N_726,N_723);
nand U826 (N_826,N_757,N_758);
or U827 (N_827,N_773,N_723);
and U828 (N_828,N_745,N_742);
nand U829 (N_829,N_720,N_771);
and U830 (N_830,N_746,N_759);
nor U831 (N_831,N_770,N_747);
nand U832 (N_832,N_762,N_753);
nand U833 (N_833,N_744,N_723);
and U834 (N_834,N_768,N_741);
and U835 (N_835,N_774,N_763);
and U836 (N_836,N_746,N_755);
and U837 (N_837,N_747,N_762);
nor U838 (N_838,N_759,N_762);
or U839 (N_839,N_746,N_734);
xor U840 (N_840,N_809,N_790);
and U841 (N_841,N_831,N_818);
nand U842 (N_842,N_791,N_792);
nand U843 (N_843,N_795,N_814);
and U844 (N_844,N_794,N_796);
or U845 (N_845,N_789,N_788);
or U846 (N_846,N_830,N_808);
or U847 (N_847,N_804,N_803);
nor U848 (N_848,N_800,N_829);
or U849 (N_849,N_838,N_780);
nand U850 (N_850,N_834,N_817);
or U851 (N_851,N_823,N_793);
xnor U852 (N_852,N_824,N_787);
nor U853 (N_853,N_781,N_785);
or U854 (N_854,N_797,N_822);
or U855 (N_855,N_836,N_819);
nor U856 (N_856,N_784,N_833);
and U857 (N_857,N_806,N_813);
and U858 (N_858,N_835,N_828);
nor U859 (N_859,N_812,N_811);
and U860 (N_860,N_820,N_798);
nor U861 (N_861,N_832,N_837);
and U862 (N_862,N_805,N_825);
xnor U863 (N_863,N_807,N_782);
nor U864 (N_864,N_799,N_783);
nor U865 (N_865,N_827,N_839);
nor U866 (N_866,N_815,N_802);
xnor U867 (N_867,N_801,N_816);
and U868 (N_868,N_821,N_810);
or U869 (N_869,N_826,N_786);
and U870 (N_870,N_835,N_799);
nor U871 (N_871,N_786,N_822);
xor U872 (N_872,N_824,N_802);
nand U873 (N_873,N_827,N_801);
or U874 (N_874,N_790,N_811);
nor U875 (N_875,N_794,N_800);
nor U876 (N_876,N_810,N_811);
and U877 (N_877,N_814,N_819);
nand U878 (N_878,N_829,N_793);
nand U879 (N_879,N_794,N_808);
nand U880 (N_880,N_784,N_832);
nor U881 (N_881,N_824,N_825);
nor U882 (N_882,N_821,N_799);
nand U883 (N_883,N_805,N_837);
and U884 (N_884,N_791,N_831);
and U885 (N_885,N_811,N_838);
or U886 (N_886,N_813,N_815);
or U887 (N_887,N_788,N_800);
nand U888 (N_888,N_839,N_834);
or U889 (N_889,N_780,N_814);
xor U890 (N_890,N_830,N_781);
or U891 (N_891,N_839,N_830);
nand U892 (N_892,N_803,N_786);
nor U893 (N_893,N_810,N_808);
or U894 (N_894,N_786,N_828);
or U895 (N_895,N_792,N_830);
or U896 (N_896,N_838,N_784);
nor U897 (N_897,N_810,N_826);
nand U898 (N_898,N_836,N_784);
nor U899 (N_899,N_829,N_811);
or U900 (N_900,N_874,N_854);
nand U901 (N_901,N_869,N_887);
nor U902 (N_902,N_856,N_883);
nor U903 (N_903,N_871,N_843);
xor U904 (N_904,N_852,N_847);
nor U905 (N_905,N_881,N_876);
and U906 (N_906,N_858,N_855);
xnor U907 (N_907,N_897,N_853);
nand U908 (N_908,N_888,N_899);
nor U909 (N_909,N_877,N_898);
or U910 (N_910,N_865,N_867);
nor U911 (N_911,N_875,N_849);
nand U912 (N_912,N_859,N_882);
or U913 (N_913,N_862,N_894);
xor U914 (N_914,N_850,N_879);
nor U915 (N_915,N_889,N_842);
nor U916 (N_916,N_864,N_845);
and U917 (N_917,N_896,N_886);
and U918 (N_918,N_895,N_866);
nor U919 (N_919,N_846,N_878);
and U920 (N_920,N_873,N_884);
nand U921 (N_921,N_893,N_890);
nand U922 (N_922,N_861,N_840);
and U923 (N_923,N_880,N_872);
or U924 (N_924,N_851,N_860);
nor U925 (N_925,N_844,N_870);
and U926 (N_926,N_841,N_891);
xor U927 (N_927,N_863,N_868);
and U928 (N_928,N_892,N_885);
nor U929 (N_929,N_848,N_857);
or U930 (N_930,N_850,N_842);
nand U931 (N_931,N_859,N_872);
or U932 (N_932,N_851,N_868);
and U933 (N_933,N_854,N_840);
nand U934 (N_934,N_847,N_896);
nand U935 (N_935,N_845,N_879);
or U936 (N_936,N_865,N_846);
xnor U937 (N_937,N_866,N_869);
nand U938 (N_938,N_886,N_885);
nor U939 (N_939,N_845,N_866);
or U940 (N_940,N_880,N_896);
xor U941 (N_941,N_845,N_893);
and U942 (N_942,N_893,N_881);
or U943 (N_943,N_886,N_888);
xnor U944 (N_944,N_894,N_879);
or U945 (N_945,N_894,N_886);
nor U946 (N_946,N_877,N_884);
nand U947 (N_947,N_891,N_880);
or U948 (N_948,N_856,N_896);
nand U949 (N_949,N_879,N_877);
and U950 (N_950,N_896,N_863);
and U951 (N_951,N_868,N_873);
and U952 (N_952,N_859,N_845);
nand U953 (N_953,N_845,N_888);
nor U954 (N_954,N_841,N_853);
nor U955 (N_955,N_850,N_856);
nand U956 (N_956,N_881,N_847);
and U957 (N_957,N_854,N_869);
or U958 (N_958,N_866,N_880);
and U959 (N_959,N_887,N_860);
nand U960 (N_960,N_943,N_923);
nor U961 (N_961,N_947,N_941);
xor U962 (N_962,N_910,N_914);
and U963 (N_963,N_921,N_945);
xor U964 (N_964,N_902,N_934);
xnor U965 (N_965,N_959,N_939);
and U966 (N_966,N_957,N_950);
nor U967 (N_967,N_901,N_911);
nand U968 (N_968,N_958,N_908);
and U969 (N_969,N_904,N_903);
xnor U970 (N_970,N_942,N_930);
xnor U971 (N_971,N_917,N_933);
nor U972 (N_972,N_949,N_940);
and U973 (N_973,N_954,N_913);
nand U974 (N_974,N_905,N_952);
xnor U975 (N_975,N_927,N_928);
nand U976 (N_976,N_956,N_948);
nand U977 (N_977,N_918,N_931);
nor U978 (N_978,N_951,N_955);
and U979 (N_979,N_906,N_929);
or U980 (N_980,N_909,N_919);
nor U981 (N_981,N_915,N_932);
nor U982 (N_982,N_936,N_907);
nor U983 (N_983,N_925,N_922);
or U984 (N_984,N_924,N_920);
nor U985 (N_985,N_944,N_900);
or U986 (N_986,N_935,N_926);
and U987 (N_987,N_946,N_938);
and U988 (N_988,N_953,N_916);
nand U989 (N_989,N_937,N_912);
nor U990 (N_990,N_915,N_947);
nand U991 (N_991,N_955,N_944);
xnor U992 (N_992,N_935,N_946);
or U993 (N_993,N_910,N_959);
or U994 (N_994,N_931,N_920);
nor U995 (N_995,N_939,N_915);
or U996 (N_996,N_916,N_926);
and U997 (N_997,N_952,N_932);
nand U998 (N_998,N_940,N_950);
and U999 (N_999,N_902,N_923);
or U1000 (N_1000,N_906,N_939);
xor U1001 (N_1001,N_901,N_958);
and U1002 (N_1002,N_950,N_954);
nor U1003 (N_1003,N_903,N_906);
nand U1004 (N_1004,N_923,N_959);
or U1005 (N_1005,N_946,N_941);
nand U1006 (N_1006,N_909,N_901);
and U1007 (N_1007,N_900,N_923);
and U1008 (N_1008,N_952,N_948);
or U1009 (N_1009,N_928,N_953);
and U1010 (N_1010,N_952,N_933);
and U1011 (N_1011,N_937,N_942);
xor U1012 (N_1012,N_917,N_955);
nor U1013 (N_1013,N_938,N_936);
nand U1014 (N_1014,N_907,N_927);
nor U1015 (N_1015,N_924,N_916);
xnor U1016 (N_1016,N_919,N_941);
nand U1017 (N_1017,N_931,N_915);
or U1018 (N_1018,N_913,N_958);
and U1019 (N_1019,N_905,N_915);
nor U1020 (N_1020,N_998,N_1011);
nand U1021 (N_1021,N_1010,N_971);
nor U1022 (N_1022,N_994,N_995);
or U1023 (N_1023,N_1019,N_966);
and U1024 (N_1024,N_986,N_992);
nand U1025 (N_1025,N_988,N_976);
nand U1026 (N_1026,N_975,N_978);
nand U1027 (N_1027,N_969,N_987);
nand U1028 (N_1028,N_982,N_983);
nand U1029 (N_1029,N_993,N_1002);
xor U1030 (N_1030,N_1009,N_964);
nor U1031 (N_1031,N_970,N_1018);
or U1032 (N_1032,N_984,N_960);
nor U1033 (N_1033,N_1006,N_996);
nor U1034 (N_1034,N_1004,N_1015);
nand U1035 (N_1035,N_973,N_967);
and U1036 (N_1036,N_1008,N_1001);
and U1037 (N_1037,N_979,N_990);
nand U1038 (N_1038,N_985,N_1012);
xnor U1039 (N_1039,N_1003,N_997);
nor U1040 (N_1040,N_961,N_968);
xor U1041 (N_1041,N_1016,N_963);
nand U1042 (N_1042,N_962,N_1007);
xor U1043 (N_1043,N_980,N_1013);
and U1044 (N_1044,N_989,N_1014);
and U1045 (N_1045,N_977,N_981);
xnor U1046 (N_1046,N_1000,N_991);
nor U1047 (N_1047,N_999,N_972);
nor U1048 (N_1048,N_974,N_1017);
nor U1049 (N_1049,N_965,N_1005);
xor U1050 (N_1050,N_1003,N_1017);
and U1051 (N_1051,N_979,N_971);
nand U1052 (N_1052,N_1017,N_1013);
nand U1053 (N_1053,N_999,N_978);
and U1054 (N_1054,N_978,N_1015);
nor U1055 (N_1055,N_1016,N_1001);
nor U1056 (N_1056,N_974,N_982);
or U1057 (N_1057,N_1004,N_976);
and U1058 (N_1058,N_997,N_975);
nand U1059 (N_1059,N_963,N_995);
and U1060 (N_1060,N_961,N_963);
or U1061 (N_1061,N_1007,N_985);
and U1062 (N_1062,N_1012,N_960);
nor U1063 (N_1063,N_998,N_992);
xor U1064 (N_1064,N_1015,N_960);
nor U1065 (N_1065,N_991,N_975);
nor U1066 (N_1066,N_1002,N_1015);
nand U1067 (N_1067,N_967,N_1018);
or U1068 (N_1068,N_963,N_984);
nor U1069 (N_1069,N_1007,N_975);
nor U1070 (N_1070,N_969,N_1016);
nor U1071 (N_1071,N_1014,N_1016);
nor U1072 (N_1072,N_985,N_1011);
nand U1073 (N_1073,N_992,N_973);
nor U1074 (N_1074,N_965,N_973);
or U1075 (N_1075,N_960,N_997);
nand U1076 (N_1076,N_980,N_1003);
nand U1077 (N_1077,N_1018,N_982);
nor U1078 (N_1078,N_966,N_970);
nor U1079 (N_1079,N_971,N_987);
or U1080 (N_1080,N_1069,N_1063);
or U1081 (N_1081,N_1023,N_1043);
or U1082 (N_1082,N_1051,N_1068);
and U1083 (N_1083,N_1039,N_1050);
nand U1084 (N_1084,N_1027,N_1077);
nand U1085 (N_1085,N_1052,N_1079);
nand U1086 (N_1086,N_1044,N_1047);
nand U1087 (N_1087,N_1049,N_1076);
and U1088 (N_1088,N_1037,N_1061);
nor U1089 (N_1089,N_1056,N_1067);
and U1090 (N_1090,N_1073,N_1078);
nor U1091 (N_1091,N_1072,N_1057);
nor U1092 (N_1092,N_1062,N_1035);
nor U1093 (N_1093,N_1033,N_1022);
xor U1094 (N_1094,N_1074,N_1038);
xor U1095 (N_1095,N_1075,N_1045);
and U1096 (N_1096,N_1021,N_1071);
or U1097 (N_1097,N_1024,N_1020);
nor U1098 (N_1098,N_1040,N_1054);
nor U1099 (N_1099,N_1025,N_1031);
nor U1100 (N_1100,N_1070,N_1060);
nand U1101 (N_1101,N_1032,N_1028);
nand U1102 (N_1102,N_1034,N_1046);
nor U1103 (N_1103,N_1029,N_1048);
or U1104 (N_1104,N_1059,N_1041);
and U1105 (N_1105,N_1065,N_1055);
nand U1106 (N_1106,N_1058,N_1030);
nor U1107 (N_1107,N_1026,N_1036);
or U1108 (N_1108,N_1066,N_1042);
nor U1109 (N_1109,N_1053,N_1064);
nor U1110 (N_1110,N_1051,N_1039);
nor U1111 (N_1111,N_1064,N_1063);
and U1112 (N_1112,N_1031,N_1020);
and U1113 (N_1113,N_1031,N_1069);
and U1114 (N_1114,N_1022,N_1059);
or U1115 (N_1115,N_1053,N_1071);
or U1116 (N_1116,N_1031,N_1037);
xor U1117 (N_1117,N_1023,N_1069);
nand U1118 (N_1118,N_1042,N_1058);
or U1119 (N_1119,N_1076,N_1074);
or U1120 (N_1120,N_1026,N_1063);
and U1121 (N_1121,N_1056,N_1040);
nor U1122 (N_1122,N_1042,N_1039);
xor U1123 (N_1123,N_1052,N_1042);
nor U1124 (N_1124,N_1046,N_1022);
and U1125 (N_1125,N_1071,N_1063);
nor U1126 (N_1126,N_1040,N_1074);
nand U1127 (N_1127,N_1065,N_1033);
xnor U1128 (N_1128,N_1022,N_1067);
nand U1129 (N_1129,N_1078,N_1079);
nand U1130 (N_1130,N_1033,N_1038);
and U1131 (N_1131,N_1055,N_1061);
nand U1132 (N_1132,N_1046,N_1037);
nand U1133 (N_1133,N_1041,N_1049);
nor U1134 (N_1134,N_1079,N_1056);
nor U1135 (N_1135,N_1060,N_1065);
and U1136 (N_1136,N_1043,N_1075);
or U1137 (N_1137,N_1045,N_1051);
and U1138 (N_1138,N_1051,N_1049);
nand U1139 (N_1139,N_1075,N_1044);
nand U1140 (N_1140,N_1087,N_1122);
nor U1141 (N_1141,N_1121,N_1091);
nor U1142 (N_1142,N_1098,N_1086);
nand U1143 (N_1143,N_1083,N_1126);
nand U1144 (N_1144,N_1102,N_1101);
nor U1145 (N_1145,N_1090,N_1137);
or U1146 (N_1146,N_1124,N_1134);
nor U1147 (N_1147,N_1112,N_1136);
nand U1148 (N_1148,N_1133,N_1113);
nand U1149 (N_1149,N_1095,N_1123);
nor U1150 (N_1150,N_1104,N_1115);
or U1151 (N_1151,N_1088,N_1080);
nor U1152 (N_1152,N_1096,N_1116);
nor U1153 (N_1153,N_1081,N_1110);
nor U1154 (N_1154,N_1111,N_1094);
and U1155 (N_1155,N_1119,N_1109);
or U1156 (N_1156,N_1132,N_1127);
or U1157 (N_1157,N_1139,N_1138);
nor U1158 (N_1158,N_1089,N_1129);
and U1159 (N_1159,N_1135,N_1130);
nor U1160 (N_1160,N_1114,N_1103);
and U1161 (N_1161,N_1084,N_1082);
or U1162 (N_1162,N_1117,N_1131);
xor U1163 (N_1163,N_1125,N_1106);
nor U1164 (N_1164,N_1092,N_1093);
or U1165 (N_1165,N_1118,N_1100);
nand U1166 (N_1166,N_1107,N_1108);
nand U1167 (N_1167,N_1097,N_1085);
nor U1168 (N_1168,N_1105,N_1099);
xnor U1169 (N_1169,N_1120,N_1128);
nor U1170 (N_1170,N_1100,N_1093);
nor U1171 (N_1171,N_1086,N_1121);
and U1172 (N_1172,N_1085,N_1093);
nor U1173 (N_1173,N_1106,N_1088);
and U1174 (N_1174,N_1135,N_1129);
or U1175 (N_1175,N_1085,N_1096);
and U1176 (N_1176,N_1097,N_1105);
nor U1177 (N_1177,N_1136,N_1080);
or U1178 (N_1178,N_1135,N_1125);
nand U1179 (N_1179,N_1129,N_1107);
and U1180 (N_1180,N_1111,N_1095);
xnor U1181 (N_1181,N_1104,N_1139);
nor U1182 (N_1182,N_1124,N_1083);
nand U1183 (N_1183,N_1118,N_1087);
nand U1184 (N_1184,N_1103,N_1090);
or U1185 (N_1185,N_1084,N_1106);
nand U1186 (N_1186,N_1122,N_1091);
nand U1187 (N_1187,N_1083,N_1110);
and U1188 (N_1188,N_1111,N_1107);
nor U1189 (N_1189,N_1112,N_1115);
nand U1190 (N_1190,N_1102,N_1109);
nor U1191 (N_1191,N_1109,N_1135);
nor U1192 (N_1192,N_1132,N_1086);
xnor U1193 (N_1193,N_1121,N_1139);
or U1194 (N_1194,N_1132,N_1080);
or U1195 (N_1195,N_1124,N_1094);
or U1196 (N_1196,N_1115,N_1099);
and U1197 (N_1197,N_1123,N_1089);
nand U1198 (N_1198,N_1103,N_1121);
or U1199 (N_1199,N_1113,N_1112);
or U1200 (N_1200,N_1176,N_1177);
nor U1201 (N_1201,N_1196,N_1149);
nand U1202 (N_1202,N_1145,N_1193);
nor U1203 (N_1203,N_1199,N_1173);
or U1204 (N_1204,N_1184,N_1190);
and U1205 (N_1205,N_1161,N_1178);
nand U1206 (N_1206,N_1197,N_1162);
or U1207 (N_1207,N_1167,N_1166);
xnor U1208 (N_1208,N_1153,N_1181);
nor U1209 (N_1209,N_1163,N_1164);
nor U1210 (N_1210,N_1179,N_1147);
nor U1211 (N_1211,N_1156,N_1160);
nand U1212 (N_1212,N_1183,N_1159);
and U1213 (N_1213,N_1185,N_1148);
and U1214 (N_1214,N_1165,N_1175);
nor U1215 (N_1215,N_1144,N_1151);
nand U1216 (N_1216,N_1143,N_1140);
nor U1217 (N_1217,N_1146,N_1172);
nor U1218 (N_1218,N_1182,N_1141);
or U1219 (N_1219,N_1154,N_1192);
nor U1220 (N_1220,N_1142,N_1188);
xor U1221 (N_1221,N_1155,N_1187);
and U1222 (N_1222,N_1194,N_1168);
nor U1223 (N_1223,N_1189,N_1198);
nand U1224 (N_1224,N_1174,N_1158);
nor U1225 (N_1225,N_1169,N_1180);
or U1226 (N_1226,N_1170,N_1191);
or U1227 (N_1227,N_1186,N_1171);
xor U1228 (N_1228,N_1152,N_1150);
or U1229 (N_1229,N_1195,N_1157);
nor U1230 (N_1230,N_1174,N_1178);
and U1231 (N_1231,N_1171,N_1177);
or U1232 (N_1232,N_1173,N_1195);
or U1233 (N_1233,N_1162,N_1196);
nor U1234 (N_1234,N_1146,N_1181);
and U1235 (N_1235,N_1191,N_1142);
nand U1236 (N_1236,N_1175,N_1164);
and U1237 (N_1237,N_1189,N_1168);
and U1238 (N_1238,N_1174,N_1196);
nand U1239 (N_1239,N_1199,N_1165);
or U1240 (N_1240,N_1180,N_1148);
or U1241 (N_1241,N_1164,N_1198);
nand U1242 (N_1242,N_1163,N_1147);
or U1243 (N_1243,N_1175,N_1148);
nand U1244 (N_1244,N_1189,N_1148);
or U1245 (N_1245,N_1160,N_1164);
xnor U1246 (N_1246,N_1166,N_1148);
nor U1247 (N_1247,N_1145,N_1156);
xor U1248 (N_1248,N_1173,N_1164);
nor U1249 (N_1249,N_1146,N_1154);
or U1250 (N_1250,N_1155,N_1178);
or U1251 (N_1251,N_1141,N_1145);
and U1252 (N_1252,N_1145,N_1151);
nand U1253 (N_1253,N_1142,N_1186);
and U1254 (N_1254,N_1177,N_1194);
nand U1255 (N_1255,N_1198,N_1183);
nand U1256 (N_1256,N_1184,N_1167);
and U1257 (N_1257,N_1194,N_1166);
and U1258 (N_1258,N_1159,N_1177);
nand U1259 (N_1259,N_1145,N_1196);
nor U1260 (N_1260,N_1227,N_1252);
and U1261 (N_1261,N_1249,N_1215);
nor U1262 (N_1262,N_1254,N_1207);
nor U1263 (N_1263,N_1209,N_1253);
nor U1264 (N_1264,N_1214,N_1235);
xnor U1265 (N_1265,N_1246,N_1229);
nor U1266 (N_1266,N_1201,N_1219);
or U1267 (N_1267,N_1248,N_1233);
and U1268 (N_1268,N_1251,N_1226);
and U1269 (N_1269,N_1228,N_1225);
or U1270 (N_1270,N_1241,N_1243);
nand U1271 (N_1271,N_1245,N_1213);
nand U1272 (N_1272,N_1221,N_1240);
or U1273 (N_1273,N_1224,N_1223);
or U1274 (N_1274,N_1250,N_1211);
nor U1275 (N_1275,N_1238,N_1230);
nand U1276 (N_1276,N_1257,N_1218);
or U1277 (N_1277,N_1234,N_1205);
and U1278 (N_1278,N_1247,N_1217);
nand U1279 (N_1279,N_1255,N_1237);
nand U1280 (N_1280,N_1202,N_1242);
nand U1281 (N_1281,N_1232,N_1259);
and U1282 (N_1282,N_1208,N_1258);
nor U1283 (N_1283,N_1239,N_1216);
and U1284 (N_1284,N_1220,N_1236);
and U1285 (N_1285,N_1212,N_1200);
and U1286 (N_1286,N_1203,N_1210);
and U1287 (N_1287,N_1244,N_1256);
nand U1288 (N_1288,N_1222,N_1231);
nand U1289 (N_1289,N_1204,N_1206);
xor U1290 (N_1290,N_1255,N_1204);
and U1291 (N_1291,N_1228,N_1247);
and U1292 (N_1292,N_1237,N_1239);
and U1293 (N_1293,N_1209,N_1227);
or U1294 (N_1294,N_1236,N_1221);
nand U1295 (N_1295,N_1242,N_1249);
or U1296 (N_1296,N_1234,N_1252);
or U1297 (N_1297,N_1249,N_1253);
nor U1298 (N_1298,N_1247,N_1224);
or U1299 (N_1299,N_1245,N_1219);
and U1300 (N_1300,N_1208,N_1225);
and U1301 (N_1301,N_1204,N_1202);
xor U1302 (N_1302,N_1234,N_1220);
or U1303 (N_1303,N_1248,N_1257);
nor U1304 (N_1304,N_1221,N_1211);
or U1305 (N_1305,N_1201,N_1208);
nor U1306 (N_1306,N_1241,N_1238);
and U1307 (N_1307,N_1233,N_1224);
nand U1308 (N_1308,N_1235,N_1225);
or U1309 (N_1309,N_1246,N_1251);
nor U1310 (N_1310,N_1212,N_1257);
xnor U1311 (N_1311,N_1256,N_1208);
nand U1312 (N_1312,N_1231,N_1226);
and U1313 (N_1313,N_1220,N_1244);
or U1314 (N_1314,N_1216,N_1205);
and U1315 (N_1315,N_1229,N_1256);
or U1316 (N_1316,N_1202,N_1219);
xnor U1317 (N_1317,N_1236,N_1239);
nor U1318 (N_1318,N_1257,N_1236);
nor U1319 (N_1319,N_1208,N_1226);
and U1320 (N_1320,N_1315,N_1272);
nand U1321 (N_1321,N_1305,N_1267);
and U1322 (N_1322,N_1260,N_1285);
or U1323 (N_1323,N_1303,N_1261);
nand U1324 (N_1324,N_1283,N_1306);
or U1325 (N_1325,N_1314,N_1308);
nor U1326 (N_1326,N_1276,N_1286);
nand U1327 (N_1327,N_1284,N_1291);
xor U1328 (N_1328,N_1313,N_1273);
or U1329 (N_1329,N_1297,N_1279);
or U1330 (N_1330,N_1296,N_1265);
and U1331 (N_1331,N_1301,N_1310);
or U1332 (N_1332,N_1312,N_1311);
and U1333 (N_1333,N_1318,N_1292);
nor U1334 (N_1334,N_1300,N_1282);
nand U1335 (N_1335,N_1299,N_1309);
or U1336 (N_1336,N_1294,N_1281);
or U1337 (N_1337,N_1316,N_1295);
or U1338 (N_1338,N_1289,N_1304);
nor U1339 (N_1339,N_1319,N_1280);
or U1340 (N_1340,N_1274,N_1302);
nand U1341 (N_1341,N_1268,N_1277);
and U1342 (N_1342,N_1290,N_1307);
nand U1343 (N_1343,N_1288,N_1262);
or U1344 (N_1344,N_1298,N_1266);
or U1345 (N_1345,N_1270,N_1317);
or U1346 (N_1346,N_1271,N_1293);
or U1347 (N_1347,N_1264,N_1287);
nor U1348 (N_1348,N_1275,N_1269);
or U1349 (N_1349,N_1278,N_1263);
nand U1350 (N_1350,N_1289,N_1287);
nor U1351 (N_1351,N_1292,N_1312);
nand U1352 (N_1352,N_1265,N_1286);
nand U1353 (N_1353,N_1304,N_1272);
nand U1354 (N_1354,N_1271,N_1286);
and U1355 (N_1355,N_1272,N_1277);
or U1356 (N_1356,N_1269,N_1296);
nand U1357 (N_1357,N_1271,N_1274);
and U1358 (N_1358,N_1283,N_1305);
or U1359 (N_1359,N_1288,N_1280);
nor U1360 (N_1360,N_1303,N_1265);
nand U1361 (N_1361,N_1273,N_1291);
xnor U1362 (N_1362,N_1291,N_1317);
and U1363 (N_1363,N_1311,N_1283);
xnor U1364 (N_1364,N_1312,N_1273);
nor U1365 (N_1365,N_1315,N_1276);
nand U1366 (N_1366,N_1278,N_1309);
or U1367 (N_1367,N_1295,N_1307);
xnor U1368 (N_1368,N_1270,N_1299);
nor U1369 (N_1369,N_1313,N_1276);
and U1370 (N_1370,N_1277,N_1300);
and U1371 (N_1371,N_1271,N_1295);
nand U1372 (N_1372,N_1268,N_1293);
nand U1373 (N_1373,N_1315,N_1263);
xnor U1374 (N_1374,N_1273,N_1302);
and U1375 (N_1375,N_1284,N_1274);
and U1376 (N_1376,N_1310,N_1278);
or U1377 (N_1377,N_1292,N_1311);
or U1378 (N_1378,N_1292,N_1293);
and U1379 (N_1379,N_1315,N_1271);
or U1380 (N_1380,N_1349,N_1322);
nand U1381 (N_1381,N_1328,N_1355);
or U1382 (N_1382,N_1373,N_1360);
nor U1383 (N_1383,N_1343,N_1340);
nor U1384 (N_1384,N_1354,N_1326);
nor U1385 (N_1385,N_1367,N_1353);
xor U1386 (N_1386,N_1369,N_1337);
or U1387 (N_1387,N_1361,N_1350);
nand U1388 (N_1388,N_1368,N_1325);
or U1389 (N_1389,N_1324,N_1348);
or U1390 (N_1390,N_1345,N_1334);
or U1391 (N_1391,N_1372,N_1356);
nand U1392 (N_1392,N_1338,N_1376);
nand U1393 (N_1393,N_1364,N_1359);
nor U1394 (N_1394,N_1358,N_1332);
or U1395 (N_1395,N_1329,N_1330);
nor U1396 (N_1396,N_1370,N_1363);
nor U1397 (N_1397,N_1327,N_1339);
nand U1398 (N_1398,N_1365,N_1366);
nor U1399 (N_1399,N_1362,N_1341);
nor U1400 (N_1400,N_1352,N_1321);
or U1401 (N_1401,N_1377,N_1371);
or U1402 (N_1402,N_1378,N_1336);
nor U1403 (N_1403,N_1357,N_1347);
nor U1404 (N_1404,N_1342,N_1344);
or U1405 (N_1405,N_1379,N_1323);
nor U1406 (N_1406,N_1351,N_1335);
xnor U1407 (N_1407,N_1375,N_1333);
nand U1408 (N_1408,N_1331,N_1320);
nand U1409 (N_1409,N_1346,N_1374);
or U1410 (N_1410,N_1377,N_1355);
or U1411 (N_1411,N_1344,N_1347);
or U1412 (N_1412,N_1354,N_1324);
nand U1413 (N_1413,N_1343,N_1368);
or U1414 (N_1414,N_1364,N_1370);
nand U1415 (N_1415,N_1326,N_1376);
and U1416 (N_1416,N_1370,N_1350);
and U1417 (N_1417,N_1348,N_1375);
nand U1418 (N_1418,N_1348,N_1351);
and U1419 (N_1419,N_1370,N_1351);
and U1420 (N_1420,N_1363,N_1367);
or U1421 (N_1421,N_1339,N_1351);
or U1422 (N_1422,N_1320,N_1374);
nor U1423 (N_1423,N_1360,N_1374);
nand U1424 (N_1424,N_1339,N_1325);
and U1425 (N_1425,N_1363,N_1344);
nor U1426 (N_1426,N_1367,N_1368);
and U1427 (N_1427,N_1324,N_1353);
or U1428 (N_1428,N_1328,N_1337);
nor U1429 (N_1429,N_1345,N_1376);
xnor U1430 (N_1430,N_1339,N_1366);
nand U1431 (N_1431,N_1327,N_1346);
xor U1432 (N_1432,N_1324,N_1327);
nand U1433 (N_1433,N_1358,N_1341);
and U1434 (N_1434,N_1340,N_1335);
nor U1435 (N_1435,N_1333,N_1351);
and U1436 (N_1436,N_1337,N_1322);
or U1437 (N_1437,N_1338,N_1369);
nand U1438 (N_1438,N_1341,N_1347);
nand U1439 (N_1439,N_1351,N_1342);
and U1440 (N_1440,N_1437,N_1439);
nor U1441 (N_1441,N_1404,N_1423);
or U1442 (N_1442,N_1430,N_1384);
nand U1443 (N_1443,N_1396,N_1388);
nand U1444 (N_1444,N_1395,N_1422);
or U1445 (N_1445,N_1411,N_1429);
and U1446 (N_1446,N_1417,N_1381);
xor U1447 (N_1447,N_1431,N_1383);
nand U1448 (N_1448,N_1391,N_1406);
or U1449 (N_1449,N_1407,N_1402);
nand U1450 (N_1450,N_1393,N_1392);
nand U1451 (N_1451,N_1425,N_1409);
nand U1452 (N_1452,N_1380,N_1415);
nand U1453 (N_1453,N_1420,N_1394);
nand U1454 (N_1454,N_1427,N_1397);
and U1455 (N_1455,N_1419,N_1390);
nor U1456 (N_1456,N_1424,N_1413);
or U1457 (N_1457,N_1416,N_1389);
or U1458 (N_1458,N_1426,N_1418);
nor U1459 (N_1459,N_1412,N_1434);
or U1460 (N_1460,N_1410,N_1408);
and U1461 (N_1461,N_1436,N_1403);
or U1462 (N_1462,N_1398,N_1400);
or U1463 (N_1463,N_1387,N_1435);
and U1464 (N_1464,N_1438,N_1433);
and U1465 (N_1465,N_1414,N_1405);
nor U1466 (N_1466,N_1385,N_1401);
xor U1467 (N_1467,N_1432,N_1428);
and U1468 (N_1468,N_1399,N_1421);
nand U1469 (N_1469,N_1386,N_1382);
or U1470 (N_1470,N_1431,N_1410);
nand U1471 (N_1471,N_1428,N_1381);
nor U1472 (N_1472,N_1431,N_1422);
or U1473 (N_1473,N_1400,N_1391);
and U1474 (N_1474,N_1391,N_1383);
nor U1475 (N_1475,N_1425,N_1395);
or U1476 (N_1476,N_1381,N_1438);
nor U1477 (N_1477,N_1414,N_1398);
nand U1478 (N_1478,N_1388,N_1387);
and U1479 (N_1479,N_1418,N_1429);
and U1480 (N_1480,N_1406,N_1409);
nand U1481 (N_1481,N_1390,N_1434);
nand U1482 (N_1482,N_1385,N_1384);
or U1483 (N_1483,N_1391,N_1381);
or U1484 (N_1484,N_1394,N_1433);
nand U1485 (N_1485,N_1381,N_1429);
and U1486 (N_1486,N_1394,N_1386);
nand U1487 (N_1487,N_1436,N_1434);
nand U1488 (N_1488,N_1421,N_1396);
nor U1489 (N_1489,N_1422,N_1392);
nor U1490 (N_1490,N_1380,N_1399);
xnor U1491 (N_1491,N_1416,N_1386);
nor U1492 (N_1492,N_1387,N_1400);
or U1493 (N_1493,N_1431,N_1406);
nor U1494 (N_1494,N_1427,N_1400);
nor U1495 (N_1495,N_1382,N_1416);
xor U1496 (N_1496,N_1411,N_1410);
and U1497 (N_1497,N_1386,N_1434);
nor U1498 (N_1498,N_1422,N_1412);
nor U1499 (N_1499,N_1428,N_1389);
and U1500 (N_1500,N_1492,N_1473);
and U1501 (N_1501,N_1499,N_1488);
nand U1502 (N_1502,N_1479,N_1478);
nand U1503 (N_1503,N_1469,N_1493);
nand U1504 (N_1504,N_1449,N_1447);
nor U1505 (N_1505,N_1475,N_1485);
nor U1506 (N_1506,N_1482,N_1466);
or U1507 (N_1507,N_1464,N_1465);
nor U1508 (N_1508,N_1495,N_1463);
or U1509 (N_1509,N_1454,N_1491);
xor U1510 (N_1510,N_1443,N_1448);
or U1511 (N_1511,N_1462,N_1490);
and U1512 (N_1512,N_1440,N_1472);
nor U1513 (N_1513,N_1455,N_1451);
or U1514 (N_1514,N_1456,N_1471);
or U1515 (N_1515,N_1477,N_1480);
and U1516 (N_1516,N_1476,N_1453);
or U1517 (N_1517,N_1496,N_1483);
and U1518 (N_1518,N_1441,N_1442);
nand U1519 (N_1519,N_1481,N_1468);
or U1520 (N_1520,N_1450,N_1487);
nor U1521 (N_1521,N_1498,N_1489);
and U1522 (N_1522,N_1445,N_1470);
nor U1523 (N_1523,N_1458,N_1460);
xnor U1524 (N_1524,N_1497,N_1484);
or U1525 (N_1525,N_1459,N_1457);
or U1526 (N_1526,N_1486,N_1467);
nor U1527 (N_1527,N_1474,N_1446);
or U1528 (N_1528,N_1452,N_1494);
nor U1529 (N_1529,N_1461,N_1444);
nor U1530 (N_1530,N_1474,N_1441);
or U1531 (N_1531,N_1498,N_1477);
and U1532 (N_1532,N_1483,N_1455);
or U1533 (N_1533,N_1486,N_1470);
nand U1534 (N_1534,N_1496,N_1470);
and U1535 (N_1535,N_1441,N_1463);
xnor U1536 (N_1536,N_1475,N_1447);
nor U1537 (N_1537,N_1499,N_1498);
nor U1538 (N_1538,N_1460,N_1498);
and U1539 (N_1539,N_1471,N_1489);
or U1540 (N_1540,N_1476,N_1473);
nor U1541 (N_1541,N_1450,N_1489);
or U1542 (N_1542,N_1446,N_1493);
or U1543 (N_1543,N_1483,N_1484);
nand U1544 (N_1544,N_1455,N_1450);
or U1545 (N_1545,N_1451,N_1450);
nor U1546 (N_1546,N_1488,N_1448);
or U1547 (N_1547,N_1441,N_1462);
or U1548 (N_1548,N_1446,N_1459);
and U1549 (N_1549,N_1482,N_1473);
and U1550 (N_1550,N_1461,N_1479);
nand U1551 (N_1551,N_1443,N_1471);
nor U1552 (N_1552,N_1474,N_1442);
and U1553 (N_1553,N_1493,N_1472);
nand U1554 (N_1554,N_1484,N_1470);
xor U1555 (N_1555,N_1451,N_1473);
or U1556 (N_1556,N_1461,N_1441);
or U1557 (N_1557,N_1462,N_1456);
or U1558 (N_1558,N_1477,N_1493);
and U1559 (N_1559,N_1499,N_1486);
and U1560 (N_1560,N_1527,N_1550);
nor U1561 (N_1561,N_1514,N_1512);
nor U1562 (N_1562,N_1555,N_1541);
and U1563 (N_1563,N_1548,N_1526);
and U1564 (N_1564,N_1538,N_1536);
nor U1565 (N_1565,N_1530,N_1513);
or U1566 (N_1566,N_1542,N_1502);
and U1567 (N_1567,N_1523,N_1511);
nor U1568 (N_1568,N_1539,N_1544);
and U1569 (N_1569,N_1510,N_1528);
nor U1570 (N_1570,N_1519,N_1503);
nor U1571 (N_1571,N_1524,N_1517);
or U1572 (N_1572,N_1553,N_1557);
nand U1573 (N_1573,N_1532,N_1543);
or U1574 (N_1574,N_1507,N_1549);
xor U1575 (N_1575,N_1551,N_1521);
or U1576 (N_1576,N_1509,N_1547);
and U1577 (N_1577,N_1515,N_1508);
nor U1578 (N_1578,N_1500,N_1505);
nand U1579 (N_1579,N_1534,N_1556);
nor U1580 (N_1580,N_1559,N_1540);
or U1581 (N_1581,N_1529,N_1554);
and U1582 (N_1582,N_1522,N_1516);
nor U1583 (N_1583,N_1546,N_1518);
and U1584 (N_1584,N_1501,N_1525);
and U1585 (N_1585,N_1537,N_1504);
xnor U1586 (N_1586,N_1531,N_1535);
xnor U1587 (N_1587,N_1533,N_1552);
and U1588 (N_1588,N_1558,N_1545);
nor U1589 (N_1589,N_1520,N_1506);
and U1590 (N_1590,N_1538,N_1518);
or U1591 (N_1591,N_1548,N_1540);
nor U1592 (N_1592,N_1540,N_1518);
and U1593 (N_1593,N_1558,N_1527);
and U1594 (N_1594,N_1547,N_1530);
and U1595 (N_1595,N_1517,N_1513);
nor U1596 (N_1596,N_1504,N_1535);
nor U1597 (N_1597,N_1507,N_1541);
or U1598 (N_1598,N_1531,N_1551);
nor U1599 (N_1599,N_1550,N_1520);
or U1600 (N_1600,N_1522,N_1553);
or U1601 (N_1601,N_1505,N_1544);
nor U1602 (N_1602,N_1508,N_1540);
nand U1603 (N_1603,N_1536,N_1501);
or U1604 (N_1604,N_1525,N_1507);
xnor U1605 (N_1605,N_1554,N_1536);
or U1606 (N_1606,N_1526,N_1528);
nand U1607 (N_1607,N_1536,N_1529);
xor U1608 (N_1608,N_1552,N_1551);
nand U1609 (N_1609,N_1501,N_1552);
nand U1610 (N_1610,N_1547,N_1517);
or U1611 (N_1611,N_1513,N_1552);
and U1612 (N_1612,N_1542,N_1504);
and U1613 (N_1613,N_1557,N_1549);
or U1614 (N_1614,N_1550,N_1518);
or U1615 (N_1615,N_1512,N_1506);
xnor U1616 (N_1616,N_1525,N_1511);
nor U1617 (N_1617,N_1528,N_1501);
nor U1618 (N_1618,N_1513,N_1512);
and U1619 (N_1619,N_1559,N_1500);
nand U1620 (N_1620,N_1604,N_1562);
nor U1621 (N_1621,N_1561,N_1610);
nor U1622 (N_1622,N_1591,N_1619);
or U1623 (N_1623,N_1593,N_1602);
xnor U1624 (N_1624,N_1581,N_1609);
nor U1625 (N_1625,N_1596,N_1566);
nand U1626 (N_1626,N_1590,N_1613);
nor U1627 (N_1627,N_1607,N_1594);
and U1628 (N_1628,N_1589,N_1588);
and U1629 (N_1629,N_1580,N_1584);
or U1630 (N_1630,N_1560,N_1614);
nor U1631 (N_1631,N_1618,N_1606);
nor U1632 (N_1632,N_1615,N_1585);
and U1633 (N_1633,N_1569,N_1617);
xnor U1634 (N_1634,N_1582,N_1570);
or U1635 (N_1635,N_1587,N_1579);
nor U1636 (N_1636,N_1599,N_1592);
or U1637 (N_1637,N_1576,N_1567);
xor U1638 (N_1638,N_1571,N_1598);
and U1639 (N_1639,N_1568,N_1575);
nand U1640 (N_1640,N_1608,N_1586);
nor U1641 (N_1641,N_1603,N_1605);
or U1642 (N_1642,N_1572,N_1616);
or U1643 (N_1643,N_1601,N_1578);
nand U1644 (N_1644,N_1563,N_1611);
and U1645 (N_1645,N_1595,N_1565);
nor U1646 (N_1646,N_1612,N_1583);
or U1647 (N_1647,N_1577,N_1573);
nor U1648 (N_1648,N_1597,N_1574);
nor U1649 (N_1649,N_1564,N_1600);
or U1650 (N_1650,N_1579,N_1562);
nand U1651 (N_1651,N_1585,N_1598);
or U1652 (N_1652,N_1609,N_1568);
and U1653 (N_1653,N_1577,N_1562);
or U1654 (N_1654,N_1603,N_1571);
or U1655 (N_1655,N_1560,N_1578);
nor U1656 (N_1656,N_1563,N_1617);
and U1657 (N_1657,N_1584,N_1578);
xor U1658 (N_1658,N_1602,N_1600);
nor U1659 (N_1659,N_1614,N_1568);
nand U1660 (N_1660,N_1566,N_1603);
or U1661 (N_1661,N_1594,N_1595);
and U1662 (N_1662,N_1608,N_1579);
and U1663 (N_1663,N_1572,N_1601);
xor U1664 (N_1664,N_1567,N_1561);
and U1665 (N_1665,N_1593,N_1596);
and U1666 (N_1666,N_1573,N_1611);
and U1667 (N_1667,N_1580,N_1599);
nand U1668 (N_1668,N_1567,N_1594);
nand U1669 (N_1669,N_1571,N_1609);
or U1670 (N_1670,N_1569,N_1564);
and U1671 (N_1671,N_1573,N_1581);
nor U1672 (N_1672,N_1575,N_1589);
or U1673 (N_1673,N_1568,N_1617);
or U1674 (N_1674,N_1604,N_1602);
and U1675 (N_1675,N_1587,N_1589);
and U1676 (N_1676,N_1619,N_1599);
nor U1677 (N_1677,N_1567,N_1579);
or U1678 (N_1678,N_1602,N_1599);
nor U1679 (N_1679,N_1560,N_1615);
nor U1680 (N_1680,N_1642,N_1659);
or U1681 (N_1681,N_1675,N_1641);
nand U1682 (N_1682,N_1635,N_1627);
and U1683 (N_1683,N_1637,N_1624);
and U1684 (N_1684,N_1633,N_1677);
and U1685 (N_1685,N_1660,N_1674);
and U1686 (N_1686,N_1667,N_1646);
nor U1687 (N_1687,N_1636,N_1666);
nor U1688 (N_1688,N_1621,N_1676);
nor U1689 (N_1689,N_1645,N_1671);
nor U1690 (N_1690,N_1670,N_1630);
and U1691 (N_1691,N_1669,N_1672);
nand U1692 (N_1692,N_1665,N_1663);
nand U1693 (N_1693,N_1678,N_1644);
or U1694 (N_1694,N_1640,N_1634);
nor U1695 (N_1695,N_1631,N_1626);
nand U1696 (N_1696,N_1628,N_1656);
xor U1697 (N_1697,N_1629,N_1662);
nand U1698 (N_1698,N_1623,N_1647);
nand U1699 (N_1699,N_1679,N_1654);
or U1700 (N_1700,N_1650,N_1652);
or U1701 (N_1701,N_1673,N_1657);
and U1702 (N_1702,N_1649,N_1622);
nor U1703 (N_1703,N_1648,N_1661);
nand U1704 (N_1704,N_1639,N_1668);
or U1705 (N_1705,N_1651,N_1655);
nor U1706 (N_1706,N_1643,N_1632);
or U1707 (N_1707,N_1620,N_1625);
xnor U1708 (N_1708,N_1638,N_1653);
and U1709 (N_1709,N_1664,N_1658);
and U1710 (N_1710,N_1643,N_1678);
or U1711 (N_1711,N_1674,N_1658);
or U1712 (N_1712,N_1675,N_1643);
and U1713 (N_1713,N_1655,N_1673);
or U1714 (N_1714,N_1668,N_1621);
or U1715 (N_1715,N_1678,N_1675);
nand U1716 (N_1716,N_1665,N_1679);
or U1717 (N_1717,N_1625,N_1657);
nand U1718 (N_1718,N_1626,N_1676);
or U1719 (N_1719,N_1637,N_1626);
and U1720 (N_1720,N_1651,N_1637);
or U1721 (N_1721,N_1661,N_1659);
xor U1722 (N_1722,N_1646,N_1671);
and U1723 (N_1723,N_1661,N_1657);
xnor U1724 (N_1724,N_1636,N_1654);
and U1725 (N_1725,N_1637,N_1620);
or U1726 (N_1726,N_1651,N_1624);
nor U1727 (N_1727,N_1658,N_1652);
or U1728 (N_1728,N_1631,N_1641);
nand U1729 (N_1729,N_1677,N_1631);
xnor U1730 (N_1730,N_1635,N_1668);
nor U1731 (N_1731,N_1634,N_1633);
nor U1732 (N_1732,N_1650,N_1649);
nor U1733 (N_1733,N_1644,N_1651);
xor U1734 (N_1734,N_1657,N_1664);
xnor U1735 (N_1735,N_1669,N_1658);
and U1736 (N_1736,N_1672,N_1623);
or U1737 (N_1737,N_1637,N_1674);
nand U1738 (N_1738,N_1635,N_1672);
nor U1739 (N_1739,N_1648,N_1634);
nor U1740 (N_1740,N_1696,N_1714);
nand U1741 (N_1741,N_1706,N_1727);
nand U1742 (N_1742,N_1720,N_1702);
nand U1743 (N_1743,N_1710,N_1734);
and U1744 (N_1744,N_1731,N_1717);
and U1745 (N_1745,N_1695,N_1704);
and U1746 (N_1746,N_1692,N_1713);
nand U1747 (N_1747,N_1680,N_1687);
xor U1748 (N_1748,N_1684,N_1705);
nand U1749 (N_1749,N_1712,N_1729);
and U1750 (N_1750,N_1736,N_1711);
nand U1751 (N_1751,N_1719,N_1722);
nand U1752 (N_1752,N_1685,N_1688);
nor U1753 (N_1753,N_1699,N_1716);
xor U1754 (N_1754,N_1700,N_1709);
or U1755 (N_1755,N_1698,N_1707);
nor U1756 (N_1756,N_1726,N_1721);
nor U1757 (N_1757,N_1724,N_1694);
and U1758 (N_1758,N_1690,N_1733);
nor U1759 (N_1759,N_1737,N_1703);
nor U1760 (N_1760,N_1701,N_1730);
and U1761 (N_1761,N_1723,N_1725);
nor U1762 (N_1762,N_1697,N_1691);
or U1763 (N_1763,N_1715,N_1683);
nor U1764 (N_1764,N_1735,N_1693);
and U1765 (N_1765,N_1686,N_1738);
nor U1766 (N_1766,N_1732,N_1718);
or U1767 (N_1767,N_1739,N_1682);
xnor U1768 (N_1768,N_1708,N_1728);
or U1769 (N_1769,N_1689,N_1681);
nand U1770 (N_1770,N_1702,N_1713);
nor U1771 (N_1771,N_1702,N_1704);
nor U1772 (N_1772,N_1701,N_1733);
nor U1773 (N_1773,N_1723,N_1686);
and U1774 (N_1774,N_1710,N_1683);
nand U1775 (N_1775,N_1700,N_1712);
or U1776 (N_1776,N_1733,N_1722);
nand U1777 (N_1777,N_1710,N_1726);
or U1778 (N_1778,N_1697,N_1716);
nand U1779 (N_1779,N_1686,N_1682);
and U1780 (N_1780,N_1710,N_1711);
or U1781 (N_1781,N_1703,N_1705);
or U1782 (N_1782,N_1696,N_1734);
nor U1783 (N_1783,N_1699,N_1732);
nor U1784 (N_1784,N_1701,N_1736);
or U1785 (N_1785,N_1691,N_1721);
xnor U1786 (N_1786,N_1722,N_1728);
nor U1787 (N_1787,N_1710,N_1714);
or U1788 (N_1788,N_1724,N_1697);
nor U1789 (N_1789,N_1695,N_1684);
or U1790 (N_1790,N_1695,N_1694);
or U1791 (N_1791,N_1687,N_1682);
nand U1792 (N_1792,N_1702,N_1724);
nand U1793 (N_1793,N_1732,N_1703);
nor U1794 (N_1794,N_1734,N_1695);
and U1795 (N_1795,N_1716,N_1696);
nor U1796 (N_1796,N_1699,N_1718);
nor U1797 (N_1797,N_1708,N_1739);
xnor U1798 (N_1798,N_1684,N_1689);
nor U1799 (N_1799,N_1691,N_1703);
nand U1800 (N_1800,N_1741,N_1748);
nor U1801 (N_1801,N_1797,N_1740);
and U1802 (N_1802,N_1795,N_1773);
nor U1803 (N_1803,N_1777,N_1780);
xor U1804 (N_1804,N_1778,N_1774);
nor U1805 (N_1805,N_1758,N_1744);
nand U1806 (N_1806,N_1743,N_1787);
nand U1807 (N_1807,N_1749,N_1766);
nand U1808 (N_1808,N_1757,N_1786);
nand U1809 (N_1809,N_1746,N_1785);
nand U1810 (N_1810,N_1779,N_1798);
and U1811 (N_1811,N_1753,N_1784);
nor U1812 (N_1812,N_1792,N_1756);
xor U1813 (N_1813,N_1755,N_1772);
nand U1814 (N_1814,N_1745,N_1770);
and U1815 (N_1815,N_1776,N_1769);
and U1816 (N_1816,N_1771,N_1760);
nand U1817 (N_1817,N_1747,N_1791);
nand U1818 (N_1818,N_1799,N_1775);
or U1819 (N_1819,N_1751,N_1793);
and U1820 (N_1820,N_1742,N_1759);
nor U1821 (N_1821,N_1754,N_1783);
xor U1822 (N_1822,N_1794,N_1764);
nor U1823 (N_1823,N_1789,N_1796);
nor U1824 (N_1824,N_1788,N_1750);
nand U1825 (N_1825,N_1761,N_1752);
and U1826 (N_1826,N_1790,N_1781);
nor U1827 (N_1827,N_1763,N_1762);
nor U1828 (N_1828,N_1768,N_1767);
or U1829 (N_1829,N_1765,N_1782);
and U1830 (N_1830,N_1763,N_1748);
and U1831 (N_1831,N_1758,N_1774);
nor U1832 (N_1832,N_1764,N_1746);
or U1833 (N_1833,N_1753,N_1766);
and U1834 (N_1834,N_1791,N_1773);
and U1835 (N_1835,N_1793,N_1762);
nand U1836 (N_1836,N_1772,N_1752);
or U1837 (N_1837,N_1797,N_1756);
and U1838 (N_1838,N_1793,N_1741);
nand U1839 (N_1839,N_1795,N_1761);
xor U1840 (N_1840,N_1796,N_1797);
and U1841 (N_1841,N_1793,N_1790);
or U1842 (N_1842,N_1781,N_1762);
xor U1843 (N_1843,N_1743,N_1745);
nor U1844 (N_1844,N_1770,N_1742);
nand U1845 (N_1845,N_1779,N_1785);
and U1846 (N_1846,N_1772,N_1767);
and U1847 (N_1847,N_1761,N_1758);
and U1848 (N_1848,N_1742,N_1768);
and U1849 (N_1849,N_1795,N_1780);
and U1850 (N_1850,N_1786,N_1774);
and U1851 (N_1851,N_1779,N_1796);
nor U1852 (N_1852,N_1790,N_1780);
and U1853 (N_1853,N_1740,N_1744);
nand U1854 (N_1854,N_1740,N_1769);
nand U1855 (N_1855,N_1769,N_1747);
nand U1856 (N_1856,N_1799,N_1787);
and U1857 (N_1857,N_1768,N_1743);
nand U1858 (N_1858,N_1765,N_1791);
or U1859 (N_1859,N_1754,N_1787);
nor U1860 (N_1860,N_1830,N_1836);
nand U1861 (N_1861,N_1812,N_1814);
nor U1862 (N_1862,N_1847,N_1832);
nor U1863 (N_1863,N_1842,N_1831);
or U1864 (N_1864,N_1829,N_1840);
nor U1865 (N_1865,N_1854,N_1834);
xor U1866 (N_1866,N_1824,N_1811);
nor U1867 (N_1867,N_1806,N_1835);
and U1868 (N_1868,N_1856,N_1817);
xnor U1869 (N_1869,N_1821,N_1841);
xor U1870 (N_1870,N_1827,N_1849);
or U1871 (N_1871,N_1838,N_1837);
and U1872 (N_1872,N_1851,N_1828);
nor U1873 (N_1873,N_1822,N_1804);
nand U1874 (N_1874,N_1807,N_1853);
nor U1875 (N_1875,N_1848,N_1819);
nand U1876 (N_1876,N_1823,N_1859);
xnor U1877 (N_1877,N_1833,N_1852);
and U1878 (N_1878,N_1813,N_1818);
xor U1879 (N_1879,N_1810,N_1805);
nor U1880 (N_1880,N_1858,N_1802);
nor U1881 (N_1881,N_1839,N_1809);
or U1882 (N_1882,N_1845,N_1800);
nor U1883 (N_1883,N_1826,N_1815);
nand U1884 (N_1884,N_1825,N_1850);
nand U1885 (N_1885,N_1843,N_1846);
nor U1886 (N_1886,N_1816,N_1803);
nand U1887 (N_1887,N_1857,N_1820);
nand U1888 (N_1888,N_1855,N_1808);
nor U1889 (N_1889,N_1844,N_1801);
and U1890 (N_1890,N_1845,N_1855);
or U1891 (N_1891,N_1820,N_1843);
nand U1892 (N_1892,N_1807,N_1847);
and U1893 (N_1893,N_1801,N_1859);
or U1894 (N_1894,N_1806,N_1844);
and U1895 (N_1895,N_1803,N_1827);
and U1896 (N_1896,N_1846,N_1852);
xor U1897 (N_1897,N_1822,N_1844);
nand U1898 (N_1898,N_1818,N_1823);
and U1899 (N_1899,N_1815,N_1823);
nor U1900 (N_1900,N_1806,N_1852);
xor U1901 (N_1901,N_1844,N_1831);
nand U1902 (N_1902,N_1800,N_1833);
nand U1903 (N_1903,N_1811,N_1845);
nor U1904 (N_1904,N_1856,N_1804);
xor U1905 (N_1905,N_1834,N_1803);
and U1906 (N_1906,N_1813,N_1811);
nor U1907 (N_1907,N_1853,N_1802);
and U1908 (N_1908,N_1828,N_1801);
xor U1909 (N_1909,N_1812,N_1831);
or U1910 (N_1910,N_1801,N_1852);
or U1911 (N_1911,N_1820,N_1805);
and U1912 (N_1912,N_1826,N_1802);
xor U1913 (N_1913,N_1841,N_1856);
and U1914 (N_1914,N_1816,N_1824);
and U1915 (N_1915,N_1857,N_1817);
nand U1916 (N_1916,N_1829,N_1808);
or U1917 (N_1917,N_1822,N_1832);
nor U1918 (N_1918,N_1835,N_1821);
nand U1919 (N_1919,N_1857,N_1821);
nor U1920 (N_1920,N_1891,N_1865);
nand U1921 (N_1921,N_1872,N_1864);
or U1922 (N_1922,N_1876,N_1901);
or U1923 (N_1923,N_1875,N_1917);
nor U1924 (N_1924,N_1916,N_1874);
and U1925 (N_1925,N_1861,N_1894);
nor U1926 (N_1926,N_1882,N_1897);
nor U1927 (N_1927,N_1887,N_1886);
nand U1928 (N_1928,N_1910,N_1905);
or U1929 (N_1929,N_1878,N_1896);
or U1930 (N_1930,N_1903,N_1869);
nor U1931 (N_1931,N_1866,N_1873);
nand U1932 (N_1932,N_1881,N_1915);
nor U1933 (N_1933,N_1885,N_1880);
nor U1934 (N_1934,N_1899,N_1893);
and U1935 (N_1935,N_1862,N_1909);
and U1936 (N_1936,N_1877,N_1904);
nor U1937 (N_1937,N_1868,N_1900);
and U1938 (N_1938,N_1898,N_1884);
and U1939 (N_1939,N_1890,N_1911);
or U1940 (N_1940,N_1883,N_1907);
and U1941 (N_1941,N_1902,N_1906);
or U1942 (N_1942,N_1892,N_1888);
and U1943 (N_1943,N_1870,N_1879);
xnor U1944 (N_1944,N_1871,N_1863);
or U1945 (N_1945,N_1908,N_1860);
or U1946 (N_1946,N_1918,N_1912);
nand U1947 (N_1947,N_1867,N_1919);
nor U1948 (N_1948,N_1913,N_1914);
and U1949 (N_1949,N_1895,N_1889);
and U1950 (N_1950,N_1867,N_1868);
nor U1951 (N_1951,N_1894,N_1867);
and U1952 (N_1952,N_1909,N_1899);
or U1953 (N_1953,N_1874,N_1863);
xnor U1954 (N_1954,N_1867,N_1902);
nor U1955 (N_1955,N_1897,N_1877);
xor U1956 (N_1956,N_1864,N_1869);
and U1957 (N_1957,N_1875,N_1874);
nand U1958 (N_1958,N_1873,N_1907);
or U1959 (N_1959,N_1919,N_1895);
nand U1960 (N_1960,N_1880,N_1860);
nor U1961 (N_1961,N_1909,N_1868);
nor U1962 (N_1962,N_1919,N_1883);
nor U1963 (N_1963,N_1907,N_1879);
or U1964 (N_1964,N_1917,N_1900);
and U1965 (N_1965,N_1881,N_1883);
nor U1966 (N_1966,N_1890,N_1876);
and U1967 (N_1967,N_1872,N_1868);
and U1968 (N_1968,N_1885,N_1890);
or U1969 (N_1969,N_1907,N_1864);
nor U1970 (N_1970,N_1880,N_1882);
or U1971 (N_1971,N_1883,N_1880);
or U1972 (N_1972,N_1902,N_1884);
and U1973 (N_1973,N_1902,N_1883);
xnor U1974 (N_1974,N_1879,N_1880);
or U1975 (N_1975,N_1863,N_1866);
and U1976 (N_1976,N_1918,N_1886);
and U1977 (N_1977,N_1867,N_1907);
or U1978 (N_1978,N_1894,N_1876);
nand U1979 (N_1979,N_1881,N_1896);
and U1980 (N_1980,N_1954,N_1957);
nand U1981 (N_1981,N_1931,N_1922);
nand U1982 (N_1982,N_1958,N_1970);
and U1983 (N_1983,N_1937,N_1972);
nor U1984 (N_1984,N_1924,N_1952);
nor U1985 (N_1985,N_1962,N_1941);
and U1986 (N_1986,N_1977,N_1939);
and U1987 (N_1987,N_1934,N_1973);
and U1988 (N_1988,N_1965,N_1921);
or U1989 (N_1989,N_1946,N_1951);
and U1990 (N_1990,N_1926,N_1932);
nor U1991 (N_1991,N_1930,N_1953);
nand U1992 (N_1992,N_1925,N_1920);
nor U1993 (N_1993,N_1947,N_1942);
or U1994 (N_1994,N_1966,N_1955);
and U1995 (N_1995,N_1964,N_1945);
nor U1996 (N_1996,N_1976,N_1936);
nor U1997 (N_1997,N_1975,N_1956);
and U1998 (N_1998,N_1971,N_1950);
nand U1999 (N_1999,N_1944,N_1923);
nor U2000 (N_2000,N_1968,N_1961);
and U2001 (N_2001,N_1929,N_1935);
nand U2002 (N_2002,N_1928,N_1959);
or U2003 (N_2003,N_1949,N_1969);
or U2004 (N_2004,N_1948,N_1974);
nor U2005 (N_2005,N_1943,N_1940);
or U2006 (N_2006,N_1927,N_1933);
nor U2007 (N_2007,N_1960,N_1963);
nor U2008 (N_2008,N_1967,N_1978);
and U2009 (N_2009,N_1979,N_1938);
nand U2010 (N_2010,N_1941,N_1932);
nor U2011 (N_2011,N_1942,N_1943);
or U2012 (N_2012,N_1924,N_1948);
xnor U2013 (N_2013,N_1971,N_1959);
or U2014 (N_2014,N_1940,N_1970);
nand U2015 (N_2015,N_1958,N_1972);
nand U2016 (N_2016,N_1953,N_1920);
nor U2017 (N_2017,N_1973,N_1942);
or U2018 (N_2018,N_1937,N_1978);
and U2019 (N_2019,N_1954,N_1936);
or U2020 (N_2020,N_1951,N_1944);
nand U2021 (N_2021,N_1957,N_1978);
nor U2022 (N_2022,N_1951,N_1957);
nor U2023 (N_2023,N_1955,N_1958);
nor U2024 (N_2024,N_1968,N_1943);
xnor U2025 (N_2025,N_1972,N_1930);
nand U2026 (N_2026,N_1927,N_1974);
and U2027 (N_2027,N_1942,N_1956);
and U2028 (N_2028,N_1960,N_1923);
nand U2029 (N_2029,N_1966,N_1921);
nand U2030 (N_2030,N_1937,N_1967);
nand U2031 (N_2031,N_1949,N_1936);
nor U2032 (N_2032,N_1976,N_1958);
or U2033 (N_2033,N_1963,N_1958);
nor U2034 (N_2034,N_1959,N_1927);
and U2035 (N_2035,N_1947,N_1959);
and U2036 (N_2036,N_1927,N_1957);
nor U2037 (N_2037,N_1948,N_1960);
nand U2038 (N_2038,N_1954,N_1931);
or U2039 (N_2039,N_1929,N_1933);
nand U2040 (N_2040,N_2012,N_2030);
nor U2041 (N_2041,N_2004,N_2005);
nand U2042 (N_2042,N_2011,N_2001);
nor U2043 (N_2043,N_1997,N_1993);
nand U2044 (N_2044,N_2035,N_2002);
or U2045 (N_2045,N_1983,N_2010);
and U2046 (N_2046,N_1986,N_1991);
and U2047 (N_2047,N_2020,N_2022);
xor U2048 (N_2048,N_2016,N_2033);
and U2049 (N_2049,N_2032,N_2037);
and U2050 (N_2050,N_1999,N_2014);
and U2051 (N_2051,N_2025,N_1994);
and U2052 (N_2052,N_1984,N_2027);
xor U2053 (N_2053,N_2038,N_2008);
or U2054 (N_2054,N_2018,N_1982);
xnor U2055 (N_2055,N_1981,N_2009);
and U2056 (N_2056,N_2039,N_1996);
and U2057 (N_2057,N_1990,N_2034);
or U2058 (N_2058,N_2028,N_1992);
nor U2059 (N_2059,N_2015,N_2036);
xnor U2060 (N_2060,N_2024,N_2000);
nand U2061 (N_2061,N_2003,N_2026);
nor U2062 (N_2062,N_1989,N_2019);
or U2063 (N_2063,N_2021,N_2023);
or U2064 (N_2064,N_1985,N_2031);
nand U2065 (N_2065,N_2007,N_2006);
and U2066 (N_2066,N_1980,N_2017);
and U2067 (N_2067,N_2013,N_1988);
or U2068 (N_2068,N_1995,N_1987);
or U2069 (N_2069,N_2029,N_1998);
nand U2070 (N_2070,N_2033,N_2014);
nor U2071 (N_2071,N_1987,N_1998);
nand U2072 (N_2072,N_1981,N_1992);
nor U2073 (N_2073,N_2036,N_1995);
nor U2074 (N_2074,N_2030,N_2028);
nand U2075 (N_2075,N_1988,N_2004);
xor U2076 (N_2076,N_1992,N_2034);
and U2077 (N_2077,N_2039,N_2012);
nand U2078 (N_2078,N_2007,N_1981);
nor U2079 (N_2079,N_2017,N_2037);
nor U2080 (N_2080,N_1989,N_2034);
or U2081 (N_2081,N_2021,N_1991);
and U2082 (N_2082,N_1989,N_2006);
and U2083 (N_2083,N_1999,N_2024);
or U2084 (N_2084,N_2026,N_2015);
nor U2085 (N_2085,N_2037,N_1989);
nor U2086 (N_2086,N_1984,N_2037);
nor U2087 (N_2087,N_2010,N_1987);
and U2088 (N_2088,N_1989,N_2004);
or U2089 (N_2089,N_2016,N_1980);
or U2090 (N_2090,N_2006,N_2038);
nor U2091 (N_2091,N_1991,N_1996);
xnor U2092 (N_2092,N_2005,N_2035);
and U2093 (N_2093,N_2006,N_2020);
or U2094 (N_2094,N_2000,N_1992);
and U2095 (N_2095,N_2004,N_1994);
nor U2096 (N_2096,N_2033,N_2005);
and U2097 (N_2097,N_1999,N_1980);
or U2098 (N_2098,N_2010,N_2027);
nor U2099 (N_2099,N_2031,N_2021);
and U2100 (N_2100,N_2099,N_2075);
nor U2101 (N_2101,N_2041,N_2092);
or U2102 (N_2102,N_2063,N_2079);
xnor U2103 (N_2103,N_2070,N_2094);
nor U2104 (N_2104,N_2093,N_2097);
xor U2105 (N_2105,N_2091,N_2089);
xnor U2106 (N_2106,N_2049,N_2060);
nand U2107 (N_2107,N_2053,N_2040);
nor U2108 (N_2108,N_2059,N_2074);
or U2109 (N_2109,N_2042,N_2064);
xor U2110 (N_2110,N_2058,N_2069);
nand U2111 (N_2111,N_2095,N_2088);
and U2112 (N_2112,N_2055,N_2083);
xor U2113 (N_2113,N_2084,N_2052);
and U2114 (N_2114,N_2090,N_2062);
and U2115 (N_2115,N_2082,N_2073);
xor U2116 (N_2116,N_2087,N_2047);
or U2117 (N_2117,N_2081,N_2066);
or U2118 (N_2118,N_2051,N_2046);
nand U2119 (N_2119,N_2072,N_2068);
or U2120 (N_2120,N_2085,N_2080);
nor U2121 (N_2121,N_2054,N_2077);
nand U2122 (N_2122,N_2050,N_2076);
nor U2123 (N_2123,N_2067,N_2096);
nand U2124 (N_2124,N_2065,N_2071);
nand U2125 (N_2125,N_2057,N_2045);
or U2126 (N_2126,N_2044,N_2048);
or U2127 (N_2127,N_2056,N_2098);
nor U2128 (N_2128,N_2061,N_2043);
nor U2129 (N_2129,N_2086,N_2078);
xnor U2130 (N_2130,N_2061,N_2088);
or U2131 (N_2131,N_2099,N_2093);
nand U2132 (N_2132,N_2044,N_2068);
nand U2133 (N_2133,N_2054,N_2071);
nand U2134 (N_2134,N_2059,N_2069);
xnor U2135 (N_2135,N_2056,N_2073);
xor U2136 (N_2136,N_2091,N_2046);
or U2137 (N_2137,N_2074,N_2070);
nor U2138 (N_2138,N_2096,N_2060);
and U2139 (N_2139,N_2076,N_2059);
and U2140 (N_2140,N_2043,N_2082);
or U2141 (N_2141,N_2081,N_2095);
or U2142 (N_2142,N_2048,N_2097);
xor U2143 (N_2143,N_2088,N_2051);
nor U2144 (N_2144,N_2072,N_2059);
or U2145 (N_2145,N_2080,N_2093);
nor U2146 (N_2146,N_2075,N_2051);
xor U2147 (N_2147,N_2079,N_2089);
nand U2148 (N_2148,N_2092,N_2050);
nor U2149 (N_2149,N_2071,N_2070);
nor U2150 (N_2150,N_2069,N_2087);
nand U2151 (N_2151,N_2071,N_2074);
or U2152 (N_2152,N_2084,N_2096);
and U2153 (N_2153,N_2089,N_2060);
or U2154 (N_2154,N_2052,N_2090);
or U2155 (N_2155,N_2042,N_2067);
nor U2156 (N_2156,N_2086,N_2089);
nand U2157 (N_2157,N_2058,N_2073);
nor U2158 (N_2158,N_2072,N_2077);
or U2159 (N_2159,N_2087,N_2092);
nand U2160 (N_2160,N_2110,N_2107);
nand U2161 (N_2161,N_2112,N_2109);
nand U2162 (N_2162,N_2104,N_2122);
nand U2163 (N_2163,N_2115,N_2123);
xor U2164 (N_2164,N_2101,N_2140);
nor U2165 (N_2165,N_2119,N_2149);
or U2166 (N_2166,N_2138,N_2129);
nor U2167 (N_2167,N_2134,N_2150);
xor U2168 (N_2168,N_2120,N_2139);
or U2169 (N_2169,N_2118,N_2106);
or U2170 (N_2170,N_2141,N_2113);
nand U2171 (N_2171,N_2108,N_2147);
nor U2172 (N_2172,N_2146,N_2127);
nor U2173 (N_2173,N_2116,N_2132);
nor U2174 (N_2174,N_2126,N_2153);
nor U2175 (N_2175,N_2103,N_2133);
or U2176 (N_2176,N_2155,N_2158);
and U2177 (N_2177,N_2142,N_2145);
nor U2178 (N_2178,N_2125,N_2148);
nor U2179 (N_2179,N_2143,N_2137);
nand U2180 (N_2180,N_2156,N_2102);
and U2181 (N_2181,N_2157,N_2130);
or U2182 (N_2182,N_2105,N_2111);
and U2183 (N_2183,N_2100,N_2159);
and U2184 (N_2184,N_2124,N_2151);
nand U2185 (N_2185,N_2136,N_2131);
or U2186 (N_2186,N_2144,N_2117);
nor U2187 (N_2187,N_2154,N_2114);
and U2188 (N_2188,N_2121,N_2135);
and U2189 (N_2189,N_2152,N_2128);
or U2190 (N_2190,N_2128,N_2104);
and U2191 (N_2191,N_2131,N_2116);
and U2192 (N_2192,N_2102,N_2145);
and U2193 (N_2193,N_2116,N_2140);
or U2194 (N_2194,N_2157,N_2139);
nand U2195 (N_2195,N_2108,N_2111);
or U2196 (N_2196,N_2141,N_2147);
nor U2197 (N_2197,N_2150,N_2109);
or U2198 (N_2198,N_2118,N_2136);
nor U2199 (N_2199,N_2134,N_2103);
and U2200 (N_2200,N_2110,N_2121);
or U2201 (N_2201,N_2155,N_2137);
xnor U2202 (N_2202,N_2112,N_2147);
and U2203 (N_2203,N_2101,N_2123);
nand U2204 (N_2204,N_2151,N_2125);
or U2205 (N_2205,N_2129,N_2134);
nor U2206 (N_2206,N_2104,N_2152);
and U2207 (N_2207,N_2128,N_2101);
and U2208 (N_2208,N_2120,N_2147);
and U2209 (N_2209,N_2111,N_2156);
or U2210 (N_2210,N_2159,N_2134);
and U2211 (N_2211,N_2148,N_2105);
nand U2212 (N_2212,N_2153,N_2110);
nor U2213 (N_2213,N_2116,N_2143);
nand U2214 (N_2214,N_2146,N_2102);
nor U2215 (N_2215,N_2108,N_2124);
nor U2216 (N_2216,N_2115,N_2119);
nor U2217 (N_2217,N_2143,N_2159);
or U2218 (N_2218,N_2155,N_2150);
or U2219 (N_2219,N_2138,N_2147);
and U2220 (N_2220,N_2195,N_2178);
or U2221 (N_2221,N_2213,N_2191);
or U2222 (N_2222,N_2211,N_2165);
xnor U2223 (N_2223,N_2200,N_2169);
nand U2224 (N_2224,N_2163,N_2201);
or U2225 (N_2225,N_2188,N_2181);
nor U2226 (N_2226,N_2192,N_2189);
or U2227 (N_2227,N_2167,N_2168);
and U2228 (N_2228,N_2217,N_2197);
nor U2229 (N_2229,N_2205,N_2160);
nand U2230 (N_2230,N_2196,N_2203);
or U2231 (N_2231,N_2198,N_2161);
xor U2232 (N_2232,N_2182,N_2199);
nor U2233 (N_2233,N_2204,N_2206);
nand U2234 (N_2234,N_2194,N_2190);
and U2235 (N_2235,N_2193,N_2184);
and U2236 (N_2236,N_2164,N_2171);
nand U2237 (N_2237,N_2172,N_2219);
or U2238 (N_2238,N_2183,N_2186);
and U2239 (N_2239,N_2214,N_2185);
xnor U2240 (N_2240,N_2166,N_2210);
nor U2241 (N_2241,N_2208,N_2176);
nand U2242 (N_2242,N_2174,N_2218);
nand U2243 (N_2243,N_2179,N_2212);
nand U2244 (N_2244,N_2202,N_2170);
and U2245 (N_2245,N_2180,N_2175);
nand U2246 (N_2246,N_2207,N_2216);
or U2247 (N_2247,N_2215,N_2173);
nand U2248 (N_2248,N_2177,N_2209);
and U2249 (N_2249,N_2187,N_2162);
or U2250 (N_2250,N_2190,N_2213);
and U2251 (N_2251,N_2217,N_2186);
and U2252 (N_2252,N_2194,N_2202);
nand U2253 (N_2253,N_2203,N_2163);
and U2254 (N_2254,N_2201,N_2186);
nand U2255 (N_2255,N_2188,N_2211);
and U2256 (N_2256,N_2164,N_2209);
nand U2257 (N_2257,N_2161,N_2182);
or U2258 (N_2258,N_2161,N_2205);
and U2259 (N_2259,N_2210,N_2197);
nand U2260 (N_2260,N_2180,N_2211);
and U2261 (N_2261,N_2208,N_2192);
or U2262 (N_2262,N_2182,N_2188);
or U2263 (N_2263,N_2211,N_2204);
and U2264 (N_2264,N_2209,N_2165);
nor U2265 (N_2265,N_2161,N_2171);
xor U2266 (N_2266,N_2167,N_2183);
or U2267 (N_2267,N_2165,N_2208);
nor U2268 (N_2268,N_2212,N_2193);
nor U2269 (N_2269,N_2170,N_2209);
and U2270 (N_2270,N_2164,N_2219);
or U2271 (N_2271,N_2184,N_2175);
and U2272 (N_2272,N_2160,N_2184);
nand U2273 (N_2273,N_2209,N_2202);
or U2274 (N_2274,N_2208,N_2204);
nor U2275 (N_2275,N_2163,N_2160);
and U2276 (N_2276,N_2192,N_2206);
nor U2277 (N_2277,N_2206,N_2197);
xnor U2278 (N_2278,N_2215,N_2184);
or U2279 (N_2279,N_2205,N_2212);
and U2280 (N_2280,N_2240,N_2237);
nor U2281 (N_2281,N_2272,N_2257);
xnor U2282 (N_2282,N_2250,N_2260);
and U2283 (N_2283,N_2224,N_2267);
or U2284 (N_2284,N_2222,N_2228);
or U2285 (N_2285,N_2236,N_2238);
or U2286 (N_2286,N_2234,N_2261);
xor U2287 (N_2287,N_2239,N_2230);
and U2288 (N_2288,N_2259,N_2226);
or U2289 (N_2289,N_2276,N_2232);
and U2290 (N_2290,N_2268,N_2273);
nor U2291 (N_2291,N_2277,N_2275);
nand U2292 (N_2292,N_2229,N_2278);
nand U2293 (N_2293,N_2274,N_2264);
nand U2294 (N_2294,N_2263,N_2252);
nand U2295 (N_2295,N_2247,N_2262);
nor U2296 (N_2296,N_2246,N_2245);
xor U2297 (N_2297,N_2279,N_2248);
nor U2298 (N_2298,N_2255,N_2258);
nand U2299 (N_2299,N_2243,N_2265);
and U2300 (N_2300,N_2253,N_2233);
nand U2301 (N_2301,N_2231,N_2266);
nor U2302 (N_2302,N_2249,N_2225);
and U2303 (N_2303,N_2256,N_2270);
and U2304 (N_2304,N_2221,N_2242);
nor U2305 (N_2305,N_2223,N_2241);
and U2306 (N_2306,N_2269,N_2254);
and U2307 (N_2307,N_2220,N_2235);
nor U2308 (N_2308,N_2227,N_2251);
or U2309 (N_2309,N_2271,N_2244);
xnor U2310 (N_2310,N_2241,N_2233);
or U2311 (N_2311,N_2274,N_2241);
nor U2312 (N_2312,N_2263,N_2269);
and U2313 (N_2313,N_2272,N_2270);
and U2314 (N_2314,N_2221,N_2274);
xor U2315 (N_2315,N_2260,N_2279);
or U2316 (N_2316,N_2231,N_2273);
nand U2317 (N_2317,N_2278,N_2238);
nor U2318 (N_2318,N_2228,N_2250);
nand U2319 (N_2319,N_2249,N_2267);
xor U2320 (N_2320,N_2246,N_2242);
nand U2321 (N_2321,N_2242,N_2233);
nor U2322 (N_2322,N_2224,N_2260);
or U2323 (N_2323,N_2257,N_2239);
nand U2324 (N_2324,N_2221,N_2249);
nor U2325 (N_2325,N_2254,N_2229);
xnor U2326 (N_2326,N_2236,N_2260);
xor U2327 (N_2327,N_2247,N_2266);
nor U2328 (N_2328,N_2269,N_2229);
and U2329 (N_2329,N_2263,N_2222);
and U2330 (N_2330,N_2231,N_2258);
or U2331 (N_2331,N_2271,N_2263);
and U2332 (N_2332,N_2261,N_2271);
nand U2333 (N_2333,N_2246,N_2277);
xor U2334 (N_2334,N_2253,N_2273);
nand U2335 (N_2335,N_2238,N_2245);
nor U2336 (N_2336,N_2253,N_2240);
nand U2337 (N_2337,N_2268,N_2252);
nand U2338 (N_2338,N_2239,N_2244);
nand U2339 (N_2339,N_2246,N_2224);
and U2340 (N_2340,N_2319,N_2330);
xnor U2341 (N_2341,N_2335,N_2291);
and U2342 (N_2342,N_2302,N_2333);
and U2343 (N_2343,N_2314,N_2337);
and U2344 (N_2344,N_2283,N_2290);
nor U2345 (N_2345,N_2334,N_2311);
or U2346 (N_2346,N_2295,N_2318);
nand U2347 (N_2347,N_2285,N_2317);
nor U2348 (N_2348,N_2320,N_2312);
or U2349 (N_2349,N_2322,N_2323);
and U2350 (N_2350,N_2321,N_2313);
nor U2351 (N_2351,N_2310,N_2339);
nor U2352 (N_2352,N_2306,N_2289);
or U2353 (N_2353,N_2286,N_2316);
nor U2354 (N_2354,N_2298,N_2328);
or U2355 (N_2355,N_2336,N_2307);
xor U2356 (N_2356,N_2299,N_2296);
and U2357 (N_2357,N_2292,N_2325);
and U2358 (N_2358,N_2332,N_2300);
xnor U2359 (N_2359,N_2282,N_2288);
nand U2360 (N_2360,N_2287,N_2280);
or U2361 (N_2361,N_2301,N_2281);
xor U2362 (N_2362,N_2297,N_2303);
nor U2363 (N_2363,N_2331,N_2326);
xnor U2364 (N_2364,N_2327,N_2305);
nand U2365 (N_2365,N_2329,N_2309);
nor U2366 (N_2366,N_2324,N_2294);
and U2367 (N_2367,N_2308,N_2293);
nand U2368 (N_2368,N_2315,N_2304);
or U2369 (N_2369,N_2338,N_2284);
and U2370 (N_2370,N_2323,N_2300);
xnor U2371 (N_2371,N_2319,N_2323);
nor U2372 (N_2372,N_2328,N_2293);
nand U2373 (N_2373,N_2281,N_2336);
xnor U2374 (N_2374,N_2289,N_2303);
and U2375 (N_2375,N_2316,N_2338);
nand U2376 (N_2376,N_2312,N_2305);
or U2377 (N_2377,N_2301,N_2323);
nor U2378 (N_2378,N_2284,N_2282);
nor U2379 (N_2379,N_2325,N_2294);
or U2380 (N_2380,N_2333,N_2311);
and U2381 (N_2381,N_2336,N_2335);
and U2382 (N_2382,N_2338,N_2294);
nand U2383 (N_2383,N_2323,N_2327);
nand U2384 (N_2384,N_2308,N_2312);
nand U2385 (N_2385,N_2323,N_2283);
or U2386 (N_2386,N_2327,N_2315);
or U2387 (N_2387,N_2291,N_2327);
and U2388 (N_2388,N_2297,N_2296);
and U2389 (N_2389,N_2293,N_2290);
nor U2390 (N_2390,N_2327,N_2338);
xnor U2391 (N_2391,N_2330,N_2318);
and U2392 (N_2392,N_2309,N_2307);
nor U2393 (N_2393,N_2313,N_2300);
or U2394 (N_2394,N_2310,N_2322);
and U2395 (N_2395,N_2298,N_2300);
nand U2396 (N_2396,N_2306,N_2339);
nand U2397 (N_2397,N_2303,N_2287);
xor U2398 (N_2398,N_2319,N_2334);
or U2399 (N_2399,N_2295,N_2310);
and U2400 (N_2400,N_2351,N_2370);
nor U2401 (N_2401,N_2377,N_2379);
nor U2402 (N_2402,N_2381,N_2366);
nand U2403 (N_2403,N_2387,N_2345);
xor U2404 (N_2404,N_2346,N_2347);
and U2405 (N_2405,N_2349,N_2367);
and U2406 (N_2406,N_2382,N_2375);
nor U2407 (N_2407,N_2342,N_2390);
nor U2408 (N_2408,N_2392,N_2356);
or U2409 (N_2409,N_2341,N_2380);
nand U2410 (N_2410,N_2350,N_2355);
nor U2411 (N_2411,N_2386,N_2357);
nor U2412 (N_2412,N_2359,N_2398);
nand U2413 (N_2413,N_2372,N_2396);
nand U2414 (N_2414,N_2376,N_2393);
nor U2415 (N_2415,N_2395,N_2360);
or U2416 (N_2416,N_2394,N_2378);
nand U2417 (N_2417,N_2399,N_2389);
or U2418 (N_2418,N_2363,N_2353);
nor U2419 (N_2419,N_2385,N_2361);
xor U2420 (N_2420,N_2354,N_2368);
and U2421 (N_2421,N_2384,N_2371);
or U2422 (N_2422,N_2374,N_2352);
or U2423 (N_2423,N_2358,N_2383);
and U2424 (N_2424,N_2348,N_2362);
xor U2425 (N_2425,N_2344,N_2365);
and U2426 (N_2426,N_2391,N_2340);
or U2427 (N_2427,N_2364,N_2388);
nor U2428 (N_2428,N_2373,N_2369);
and U2429 (N_2429,N_2343,N_2397);
nor U2430 (N_2430,N_2378,N_2393);
or U2431 (N_2431,N_2354,N_2389);
nor U2432 (N_2432,N_2359,N_2396);
nor U2433 (N_2433,N_2389,N_2387);
or U2434 (N_2434,N_2359,N_2387);
and U2435 (N_2435,N_2395,N_2372);
nor U2436 (N_2436,N_2341,N_2398);
and U2437 (N_2437,N_2363,N_2364);
and U2438 (N_2438,N_2365,N_2359);
and U2439 (N_2439,N_2342,N_2348);
nand U2440 (N_2440,N_2370,N_2348);
or U2441 (N_2441,N_2394,N_2365);
nand U2442 (N_2442,N_2364,N_2389);
nand U2443 (N_2443,N_2385,N_2386);
nand U2444 (N_2444,N_2390,N_2366);
and U2445 (N_2445,N_2383,N_2359);
nand U2446 (N_2446,N_2357,N_2369);
nor U2447 (N_2447,N_2359,N_2395);
nand U2448 (N_2448,N_2356,N_2375);
or U2449 (N_2449,N_2390,N_2350);
or U2450 (N_2450,N_2376,N_2367);
nand U2451 (N_2451,N_2357,N_2380);
and U2452 (N_2452,N_2367,N_2377);
nor U2453 (N_2453,N_2371,N_2344);
xnor U2454 (N_2454,N_2363,N_2395);
xor U2455 (N_2455,N_2393,N_2360);
and U2456 (N_2456,N_2373,N_2380);
nand U2457 (N_2457,N_2389,N_2343);
and U2458 (N_2458,N_2345,N_2347);
or U2459 (N_2459,N_2344,N_2398);
nor U2460 (N_2460,N_2456,N_2409);
and U2461 (N_2461,N_2430,N_2446);
or U2462 (N_2462,N_2437,N_2458);
nand U2463 (N_2463,N_2427,N_2423);
nor U2464 (N_2464,N_2452,N_2404);
or U2465 (N_2465,N_2453,N_2420);
nor U2466 (N_2466,N_2411,N_2444);
nor U2467 (N_2467,N_2421,N_2450);
or U2468 (N_2468,N_2401,N_2432);
and U2469 (N_2469,N_2433,N_2414);
nor U2470 (N_2470,N_2410,N_2429);
nand U2471 (N_2471,N_2407,N_2406);
nor U2472 (N_2472,N_2403,N_2455);
and U2473 (N_2473,N_2457,N_2408);
nor U2474 (N_2474,N_2424,N_2440);
or U2475 (N_2475,N_2451,N_2426);
xor U2476 (N_2476,N_2417,N_2447);
nand U2477 (N_2477,N_2428,N_2416);
nand U2478 (N_2478,N_2412,N_2439);
or U2479 (N_2479,N_2413,N_2459);
and U2480 (N_2480,N_2441,N_2400);
and U2481 (N_2481,N_2438,N_2402);
nor U2482 (N_2482,N_2405,N_2449);
nor U2483 (N_2483,N_2422,N_2448);
or U2484 (N_2484,N_2436,N_2435);
nor U2485 (N_2485,N_2454,N_2415);
xnor U2486 (N_2486,N_2431,N_2445);
or U2487 (N_2487,N_2425,N_2442);
and U2488 (N_2488,N_2418,N_2434);
or U2489 (N_2489,N_2419,N_2443);
nand U2490 (N_2490,N_2424,N_2445);
and U2491 (N_2491,N_2419,N_2411);
and U2492 (N_2492,N_2453,N_2433);
and U2493 (N_2493,N_2430,N_2423);
nor U2494 (N_2494,N_2430,N_2447);
or U2495 (N_2495,N_2403,N_2432);
or U2496 (N_2496,N_2456,N_2433);
nor U2497 (N_2497,N_2458,N_2422);
or U2498 (N_2498,N_2425,N_2409);
and U2499 (N_2499,N_2428,N_2442);
or U2500 (N_2500,N_2430,N_2425);
or U2501 (N_2501,N_2457,N_2450);
and U2502 (N_2502,N_2412,N_2405);
xor U2503 (N_2503,N_2451,N_2422);
and U2504 (N_2504,N_2420,N_2444);
nor U2505 (N_2505,N_2410,N_2437);
and U2506 (N_2506,N_2454,N_2444);
nand U2507 (N_2507,N_2401,N_2440);
xor U2508 (N_2508,N_2454,N_2437);
or U2509 (N_2509,N_2435,N_2456);
nor U2510 (N_2510,N_2448,N_2450);
nor U2511 (N_2511,N_2443,N_2437);
nand U2512 (N_2512,N_2409,N_2423);
and U2513 (N_2513,N_2411,N_2436);
xnor U2514 (N_2514,N_2413,N_2448);
nor U2515 (N_2515,N_2437,N_2400);
nand U2516 (N_2516,N_2419,N_2427);
and U2517 (N_2517,N_2435,N_2418);
and U2518 (N_2518,N_2412,N_2432);
nor U2519 (N_2519,N_2401,N_2416);
xor U2520 (N_2520,N_2513,N_2514);
nor U2521 (N_2521,N_2506,N_2467);
or U2522 (N_2522,N_2491,N_2476);
nand U2523 (N_2523,N_2499,N_2502);
nor U2524 (N_2524,N_2495,N_2484);
or U2525 (N_2525,N_2477,N_2483);
or U2526 (N_2526,N_2475,N_2516);
and U2527 (N_2527,N_2519,N_2482);
and U2528 (N_2528,N_2490,N_2472);
or U2529 (N_2529,N_2481,N_2461);
nor U2530 (N_2530,N_2487,N_2508);
and U2531 (N_2531,N_2515,N_2466);
nand U2532 (N_2532,N_2473,N_2494);
or U2533 (N_2533,N_2480,N_2503);
xnor U2534 (N_2534,N_2511,N_2507);
nor U2535 (N_2535,N_2470,N_2504);
nor U2536 (N_2536,N_2493,N_2469);
nor U2537 (N_2537,N_2463,N_2474);
or U2538 (N_2538,N_2488,N_2486);
nand U2539 (N_2539,N_2492,N_2501);
or U2540 (N_2540,N_2478,N_2464);
or U2541 (N_2541,N_2518,N_2496);
or U2542 (N_2542,N_2505,N_2471);
nor U2543 (N_2543,N_2517,N_2512);
nor U2544 (N_2544,N_2489,N_2509);
nand U2545 (N_2545,N_2468,N_2479);
nand U2546 (N_2546,N_2462,N_2500);
nor U2547 (N_2547,N_2460,N_2510);
nor U2548 (N_2548,N_2498,N_2465);
nor U2549 (N_2549,N_2497,N_2485);
or U2550 (N_2550,N_2511,N_2512);
nor U2551 (N_2551,N_2480,N_2507);
nand U2552 (N_2552,N_2483,N_2479);
nor U2553 (N_2553,N_2467,N_2485);
and U2554 (N_2554,N_2503,N_2498);
nor U2555 (N_2555,N_2465,N_2466);
nor U2556 (N_2556,N_2508,N_2498);
xor U2557 (N_2557,N_2486,N_2469);
nor U2558 (N_2558,N_2514,N_2507);
and U2559 (N_2559,N_2518,N_2512);
and U2560 (N_2560,N_2482,N_2484);
or U2561 (N_2561,N_2518,N_2480);
and U2562 (N_2562,N_2475,N_2496);
and U2563 (N_2563,N_2493,N_2490);
nor U2564 (N_2564,N_2505,N_2475);
and U2565 (N_2565,N_2511,N_2462);
or U2566 (N_2566,N_2486,N_2514);
and U2567 (N_2567,N_2465,N_2516);
nand U2568 (N_2568,N_2519,N_2512);
nand U2569 (N_2569,N_2511,N_2499);
and U2570 (N_2570,N_2508,N_2507);
and U2571 (N_2571,N_2501,N_2496);
nand U2572 (N_2572,N_2470,N_2462);
and U2573 (N_2573,N_2473,N_2516);
or U2574 (N_2574,N_2507,N_2469);
nand U2575 (N_2575,N_2511,N_2505);
nor U2576 (N_2576,N_2479,N_2508);
or U2577 (N_2577,N_2502,N_2501);
xnor U2578 (N_2578,N_2468,N_2484);
or U2579 (N_2579,N_2519,N_2497);
or U2580 (N_2580,N_2538,N_2531);
nor U2581 (N_2581,N_2535,N_2522);
xor U2582 (N_2582,N_2575,N_2558);
or U2583 (N_2583,N_2566,N_2523);
xnor U2584 (N_2584,N_2525,N_2559);
nand U2585 (N_2585,N_2556,N_2555);
nor U2586 (N_2586,N_2530,N_2551);
nor U2587 (N_2587,N_2564,N_2569);
or U2588 (N_2588,N_2528,N_2553);
or U2589 (N_2589,N_2560,N_2579);
and U2590 (N_2590,N_2529,N_2554);
xnor U2591 (N_2591,N_2561,N_2521);
xor U2592 (N_2592,N_2526,N_2536);
nor U2593 (N_2593,N_2550,N_2541);
nor U2594 (N_2594,N_2543,N_2563);
nand U2595 (N_2595,N_2576,N_2533);
nand U2596 (N_2596,N_2547,N_2545);
xnor U2597 (N_2597,N_2573,N_2578);
xnor U2598 (N_2598,N_2532,N_2552);
and U2599 (N_2599,N_2537,N_2549);
and U2600 (N_2600,N_2570,N_2574);
and U2601 (N_2601,N_2542,N_2548);
nor U2602 (N_2602,N_2577,N_2562);
nand U2603 (N_2603,N_2524,N_2557);
or U2604 (N_2604,N_2534,N_2565);
and U2605 (N_2605,N_2540,N_2544);
nand U2606 (N_2606,N_2572,N_2568);
nand U2607 (N_2607,N_2567,N_2571);
and U2608 (N_2608,N_2539,N_2520);
nor U2609 (N_2609,N_2546,N_2527);
xor U2610 (N_2610,N_2526,N_2547);
or U2611 (N_2611,N_2522,N_2549);
nor U2612 (N_2612,N_2552,N_2548);
nand U2613 (N_2613,N_2524,N_2546);
and U2614 (N_2614,N_2537,N_2536);
nand U2615 (N_2615,N_2560,N_2536);
nand U2616 (N_2616,N_2561,N_2545);
and U2617 (N_2617,N_2575,N_2536);
or U2618 (N_2618,N_2579,N_2552);
xnor U2619 (N_2619,N_2530,N_2555);
nor U2620 (N_2620,N_2575,N_2533);
nor U2621 (N_2621,N_2540,N_2576);
and U2622 (N_2622,N_2546,N_2547);
and U2623 (N_2623,N_2576,N_2553);
nor U2624 (N_2624,N_2562,N_2551);
nand U2625 (N_2625,N_2571,N_2561);
or U2626 (N_2626,N_2541,N_2552);
nor U2627 (N_2627,N_2562,N_2535);
or U2628 (N_2628,N_2559,N_2561);
nor U2629 (N_2629,N_2554,N_2558);
or U2630 (N_2630,N_2576,N_2527);
nand U2631 (N_2631,N_2527,N_2547);
xor U2632 (N_2632,N_2562,N_2566);
or U2633 (N_2633,N_2558,N_2563);
or U2634 (N_2634,N_2541,N_2560);
or U2635 (N_2635,N_2544,N_2554);
nor U2636 (N_2636,N_2538,N_2551);
or U2637 (N_2637,N_2564,N_2546);
xor U2638 (N_2638,N_2531,N_2525);
nand U2639 (N_2639,N_2545,N_2579);
nor U2640 (N_2640,N_2627,N_2582);
xor U2641 (N_2641,N_2606,N_2603);
nor U2642 (N_2642,N_2580,N_2589);
and U2643 (N_2643,N_2610,N_2605);
xor U2644 (N_2644,N_2602,N_2633);
xor U2645 (N_2645,N_2609,N_2612);
or U2646 (N_2646,N_2621,N_2599);
nand U2647 (N_2647,N_2629,N_2588);
or U2648 (N_2648,N_2597,N_2592);
nand U2649 (N_2649,N_2637,N_2586);
or U2650 (N_2650,N_2593,N_2581);
and U2651 (N_2651,N_2616,N_2587);
and U2652 (N_2652,N_2594,N_2584);
and U2653 (N_2653,N_2631,N_2639);
and U2654 (N_2654,N_2618,N_2628);
and U2655 (N_2655,N_2617,N_2626);
xnor U2656 (N_2656,N_2632,N_2619);
nand U2657 (N_2657,N_2636,N_2614);
and U2658 (N_2658,N_2611,N_2634);
or U2659 (N_2659,N_2585,N_2638);
nand U2660 (N_2660,N_2604,N_2620);
and U2661 (N_2661,N_2625,N_2598);
or U2662 (N_2662,N_2630,N_2590);
and U2663 (N_2663,N_2591,N_2607);
and U2664 (N_2664,N_2601,N_2635);
and U2665 (N_2665,N_2622,N_2615);
nor U2666 (N_2666,N_2596,N_2624);
and U2667 (N_2667,N_2608,N_2613);
or U2668 (N_2668,N_2583,N_2595);
nor U2669 (N_2669,N_2623,N_2600);
nor U2670 (N_2670,N_2613,N_2601);
and U2671 (N_2671,N_2607,N_2625);
nand U2672 (N_2672,N_2604,N_2586);
and U2673 (N_2673,N_2615,N_2614);
nor U2674 (N_2674,N_2634,N_2615);
and U2675 (N_2675,N_2636,N_2623);
nor U2676 (N_2676,N_2607,N_2604);
nor U2677 (N_2677,N_2630,N_2602);
and U2678 (N_2678,N_2638,N_2611);
and U2679 (N_2679,N_2631,N_2621);
nor U2680 (N_2680,N_2599,N_2600);
and U2681 (N_2681,N_2582,N_2588);
nor U2682 (N_2682,N_2626,N_2622);
nor U2683 (N_2683,N_2587,N_2637);
or U2684 (N_2684,N_2614,N_2620);
or U2685 (N_2685,N_2606,N_2626);
and U2686 (N_2686,N_2580,N_2626);
nand U2687 (N_2687,N_2609,N_2607);
or U2688 (N_2688,N_2591,N_2590);
and U2689 (N_2689,N_2631,N_2584);
or U2690 (N_2690,N_2638,N_2601);
or U2691 (N_2691,N_2612,N_2638);
nand U2692 (N_2692,N_2631,N_2609);
nand U2693 (N_2693,N_2582,N_2629);
nor U2694 (N_2694,N_2606,N_2631);
xor U2695 (N_2695,N_2611,N_2637);
nand U2696 (N_2696,N_2627,N_2630);
nor U2697 (N_2697,N_2634,N_2585);
or U2698 (N_2698,N_2603,N_2586);
nor U2699 (N_2699,N_2620,N_2595);
or U2700 (N_2700,N_2692,N_2662);
or U2701 (N_2701,N_2664,N_2660);
xor U2702 (N_2702,N_2667,N_2681);
and U2703 (N_2703,N_2696,N_2655);
xor U2704 (N_2704,N_2685,N_2641);
and U2705 (N_2705,N_2697,N_2647);
or U2706 (N_2706,N_2679,N_2657);
nor U2707 (N_2707,N_2666,N_2680);
nor U2708 (N_2708,N_2693,N_2674);
nand U2709 (N_2709,N_2695,N_2675);
or U2710 (N_2710,N_2659,N_2670);
nor U2711 (N_2711,N_2646,N_2658);
or U2712 (N_2712,N_2690,N_2640);
nand U2713 (N_2713,N_2688,N_2653);
or U2714 (N_2714,N_2652,N_2698);
nand U2715 (N_2715,N_2661,N_2691);
and U2716 (N_2716,N_2672,N_2665);
or U2717 (N_2717,N_2678,N_2682);
or U2718 (N_2718,N_2644,N_2687);
and U2719 (N_2719,N_2654,N_2684);
nand U2720 (N_2720,N_2649,N_2650);
nor U2721 (N_2721,N_2699,N_2668);
or U2722 (N_2722,N_2643,N_2694);
nand U2723 (N_2723,N_2645,N_2642);
and U2724 (N_2724,N_2686,N_2676);
nand U2725 (N_2725,N_2677,N_2669);
xor U2726 (N_2726,N_2689,N_2683);
xor U2727 (N_2727,N_2656,N_2648);
nand U2728 (N_2728,N_2673,N_2671);
or U2729 (N_2729,N_2663,N_2651);
xor U2730 (N_2730,N_2664,N_2679);
nor U2731 (N_2731,N_2682,N_2669);
or U2732 (N_2732,N_2676,N_2691);
or U2733 (N_2733,N_2646,N_2678);
or U2734 (N_2734,N_2696,N_2678);
and U2735 (N_2735,N_2674,N_2691);
nor U2736 (N_2736,N_2692,N_2650);
nor U2737 (N_2737,N_2665,N_2699);
and U2738 (N_2738,N_2697,N_2648);
or U2739 (N_2739,N_2640,N_2665);
nand U2740 (N_2740,N_2662,N_2666);
nand U2741 (N_2741,N_2674,N_2694);
or U2742 (N_2742,N_2664,N_2689);
and U2743 (N_2743,N_2679,N_2647);
nand U2744 (N_2744,N_2657,N_2673);
or U2745 (N_2745,N_2656,N_2672);
nor U2746 (N_2746,N_2647,N_2672);
xor U2747 (N_2747,N_2641,N_2658);
or U2748 (N_2748,N_2686,N_2696);
or U2749 (N_2749,N_2663,N_2643);
and U2750 (N_2750,N_2695,N_2677);
or U2751 (N_2751,N_2663,N_2640);
nand U2752 (N_2752,N_2689,N_2651);
and U2753 (N_2753,N_2668,N_2648);
and U2754 (N_2754,N_2646,N_2681);
and U2755 (N_2755,N_2665,N_2692);
nand U2756 (N_2756,N_2687,N_2648);
and U2757 (N_2757,N_2669,N_2681);
or U2758 (N_2758,N_2640,N_2678);
and U2759 (N_2759,N_2648,N_2676);
xor U2760 (N_2760,N_2715,N_2709);
xnor U2761 (N_2761,N_2755,N_2706);
nand U2762 (N_2762,N_2744,N_2724);
nand U2763 (N_2763,N_2729,N_2743);
or U2764 (N_2764,N_2725,N_2702);
nand U2765 (N_2765,N_2708,N_2736);
and U2766 (N_2766,N_2719,N_2734);
nand U2767 (N_2767,N_2759,N_2738);
nor U2768 (N_2768,N_2748,N_2717);
and U2769 (N_2769,N_2716,N_2726);
nor U2770 (N_2770,N_2723,N_2735);
and U2771 (N_2771,N_2728,N_2746);
and U2772 (N_2772,N_2751,N_2756);
nor U2773 (N_2773,N_2710,N_2737);
nor U2774 (N_2774,N_2745,N_2742);
xnor U2775 (N_2775,N_2754,N_2733);
nand U2776 (N_2776,N_2732,N_2730);
or U2777 (N_2777,N_2700,N_2701);
nor U2778 (N_2778,N_2749,N_2739);
and U2779 (N_2779,N_2757,N_2705);
and U2780 (N_2780,N_2727,N_2714);
nor U2781 (N_2781,N_2704,N_2731);
or U2782 (N_2782,N_2753,N_2712);
nor U2783 (N_2783,N_2720,N_2741);
and U2784 (N_2784,N_2707,N_2740);
nand U2785 (N_2785,N_2718,N_2752);
and U2786 (N_2786,N_2722,N_2711);
nand U2787 (N_2787,N_2747,N_2750);
nand U2788 (N_2788,N_2703,N_2713);
nor U2789 (N_2789,N_2721,N_2758);
nand U2790 (N_2790,N_2701,N_2748);
and U2791 (N_2791,N_2734,N_2755);
nor U2792 (N_2792,N_2712,N_2736);
and U2793 (N_2793,N_2732,N_2757);
nand U2794 (N_2794,N_2759,N_2727);
and U2795 (N_2795,N_2746,N_2756);
nand U2796 (N_2796,N_2722,N_2738);
nor U2797 (N_2797,N_2744,N_2746);
nand U2798 (N_2798,N_2709,N_2735);
and U2799 (N_2799,N_2713,N_2727);
and U2800 (N_2800,N_2748,N_2758);
nand U2801 (N_2801,N_2716,N_2722);
nand U2802 (N_2802,N_2751,N_2729);
and U2803 (N_2803,N_2724,N_2745);
nand U2804 (N_2804,N_2741,N_2721);
or U2805 (N_2805,N_2741,N_2710);
nand U2806 (N_2806,N_2730,N_2725);
and U2807 (N_2807,N_2757,N_2734);
or U2808 (N_2808,N_2705,N_2744);
xor U2809 (N_2809,N_2715,N_2716);
nor U2810 (N_2810,N_2717,N_2734);
nand U2811 (N_2811,N_2751,N_2719);
nor U2812 (N_2812,N_2731,N_2742);
nand U2813 (N_2813,N_2734,N_2742);
or U2814 (N_2814,N_2748,N_2703);
nand U2815 (N_2815,N_2715,N_2740);
and U2816 (N_2816,N_2755,N_2701);
nand U2817 (N_2817,N_2724,N_2716);
xnor U2818 (N_2818,N_2701,N_2702);
nor U2819 (N_2819,N_2714,N_2720);
nand U2820 (N_2820,N_2784,N_2766);
nor U2821 (N_2821,N_2791,N_2760);
and U2822 (N_2822,N_2783,N_2802);
xor U2823 (N_2823,N_2776,N_2800);
nor U2824 (N_2824,N_2806,N_2818);
nand U2825 (N_2825,N_2798,N_2770);
nor U2826 (N_2826,N_2761,N_2797);
xnor U2827 (N_2827,N_2777,N_2792);
xnor U2828 (N_2828,N_2793,N_2765);
and U2829 (N_2829,N_2786,N_2772);
or U2830 (N_2830,N_2812,N_2808);
nor U2831 (N_2831,N_2795,N_2788);
or U2832 (N_2832,N_2767,N_2778);
xor U2833 (N_2833,N_2787,N_2811);
nand U2834 (N_2834,N_2807,N_2815);
and U2835 (N_2835,N_2763,N_2764);
or U2836 (N_2836,N_2779,N_2780);
and U2837 (N_2837,N_2817,N_2774);
or U2838 (N_2838,N_2768,N_2773);
nand U2839 (N_2839,N_2803,N_2785);
nor U2840 (N_2840,N_2769,N_2782);
and U2841 (N_2841,N_2781,N_2790);
nor U2842 (N_2842,N_2810,N_2775);
xnor U2843 (N_2843,N_2789,N_2819);
xnor U2844 (N_2844,N_2771,N_2814);
nand U2845 (N_2845,N_2801,N_2813);
and U2846 (N_2846,N_2805,N_2762);
nand U2847 (N_2847,N_2816,N_2809);
nor U2848 (N_2848,N_2796,N_2804);
nand U2849 (N_2849,N_2794,N_2799);
nor U2850 (N_2850,N_2816,N_2767);
or U2851 (N_2851,N_2764,N_2786);
or U2852 (N_2852,N_2804,N_2760);
nand U2853 (N_2853,N_2783,N_2781);
or U2854 (N_2854,N_2809,N_2808);
nand U2855 (N_2855,N_2819,N_2760);
nor U2856 (N_2856,N_2797,N_2807);
and U2857 (N_2857,N_2786,N_2805);
nand U2858 (N_2858,N_2805,N_2780);
nor U2859 (N_2859,N_2813,N_2818);
nand U2860 (N_2860,N_2786,N_2809);
or U2861 (N_2861,N_2775,N_2771);
nor U2862 (N_2862,N_2791,N_2799);
and U2863 (N_2863,N_2796,N_2765);
and U2864 (N_2864,N_2769,N_2803);
nand U2865 (N_2865,N_2772,N_2782);
and U2866 (N_2866,N_2815,N_2808);
and U2867 (N_2867,N_2796,N_2786);
nor U2868 (N_2868,N_2778,N_2773);
nor U2869 (N_2869,N_2781,N_2761);
nand U2870 (N_2870,N_2817,N_2791);
and U2871 (N_2871,N_2786,N_2813);
nor U2872 (N_2872,N_2781,N_2765);
and U2873 (N_2873,N_2790,N_2774);
nor U2874 (N_2874,N_2806,N_2789);
and U2875 (N_2875,N_2782,N_2792);
nand U2876 (N_2876,N_2798,N_2787);
nor U2877 (N_2877,N_2774,N_2787);
nor U2878 (N_2878,N_2799,N_2777);
nor U2879 (N_2879,N_2809,N_2790);
and U2880 (N_2880,N_2848,N_2843);
and U2881 (N_2881,N_2863,N_2850);
and U2882 (N_2882,N_2876,N_2856);
nand U2883 (N_2883,N_2872,N_2827);
nand U2884 (N_2884,N_2825,N_2854);
nand U2885 (N_2885,N_2851,N_2874);
nor U2886 (N_2886,N_2832,N_2878);
and U2887 (N_2887,N_2824,N_2870);
nand U2888 (N_2888,N_2820,N_2867);
nand U2889 (N_2889,N_2841,N_2861);
and U2890 (N_2890,N_2837,N_2866);
or U2891 (N_2891,N_2849,N_2871);
or U2892 (N_2892,N_2838,N_2862);
xnor U2893 (N_2893,N_2846,N_2845);
nand U2894 (N_2894,N_2853,N_2833);
or U2895 (N_2895,N_2836,N_2859);
nor U2896 (N_2896,N_2830,N_2847);
nand U2897 (N_2897,N_2826,N_2831);
xnor U2898 (N_2898,N_2835,N_2821);
xor U2899 (N_2899,N_2842,N_2834);
xor U2900 (N_2900,N_2864,N_2828);
nand U2901 (N_2901,N_2869,N_2829);
nor U2902 (N_2902,N_2877,N_2823);
xnor U2903 (N_2903,N_2857,N_2844);
xor U2904 (N_2904,N_2860,N_2840);
or U2905 (N_2905,N_2852,N_2873);
or U2906 (N_2906,N_2839,N_2865);
and U2907 (N_2907,N_2822,N_2855);
or U2908 (N_2908,N_2868,N_2858);
xnor U2909 (N_2909,N_2879,N_2875);
nand U2910 (N_2910,N_2842,N_2821);
and U2911 (N_2911,N_2829,N_2853);
nand U2912 (N_2912,N_2827,N_2857);
or U2913 (N_2913,N_2858,N_2822);
nor U2914 (N_2914,N_2841,N_2828);
nand U2915 (N_2915,N_2824,N_2839);
or U2916 (N_2916,N_2878,N_2856);
nor U2917 (N_2917,N_2873,N_2835);
and U2918 (N_2918,N_2832,N_2865);
and U2919 (N_2919,N_2837,N_2865);
nor U2920 (N_2920,N_2839,N_2866);
xnor U2921 (N_2921,N_2855,N_2875);
nor U2922 (N_2922,N_2833,N_2840);
nor U2923 (N_2923,N_2825,N_2828);
xnor U2924 (N_2924,N_2846,N_2875);
and U2925 (N_2925,N_2840,N_2851);
nand U2926 (N_2926,N_2827,N_2835);
or U2927 (N_2927,N_2868,N_2855);
and U2928 (N_2928,N_2867,N_2849);
nand U2929 (N_2929,N_2878,N_2860);
nor U2930 (N_2930,N_2879,N_2834);
and U2931 (N_2931,N_2868,N_2842);
nand U2932 (N_2932,N_2851,N_2824);
xnor U2933 (N_2933,N_2831,N_2852);
nand U2934 (N_2934,N_2828,N_2839);
nor U2935 (N_2935,N_2825,N_2877);
or U2936 (N_2936,N_2844,N_2867);
and U2937 (N_2937,N_2878,N_2833);
nand U2938 (N_2938,N_2845,N_2875);
nand U2939 (N_2939,N_2841,N_2864);
and U2940 (N_2940,N_2934,N_2937);
and U2941 (N_2941,N_2887,N_2895);
nor U2942 (N_2942,N_2908,N_2893);
and U2943 (N_2943,N_2932,N_2916);
and U2944 (N_2944,N_2905,N_2909);
or U2945 (N_2945,N_2894,N_2891);
nor U2946 (N_2946,N_2892,N_2914);
nor U2947 (N_2947,N_2936,N_2933);
or U2948 (N_2948,N_2915,N_2917);
xnor U2949 (N_2949,N_2900,N_2913);
nand U2950 (N_2950,N_2920,N_2903);
or U2951 (N_2951,N_2939,N_2912);
and U2952 (N_2952,N_2931,N_2896);
nor U2953 (N_2953,N_2884,N_2885);
nand U2954 (N_2954,N_2899,N_2935);
and U2955 (N_2955,N_2881,N_2923);
and U2956 (N_2956,N_2910,N_2888);
and U2957 (N_2957,N_2880,N_2907);
or U2958 (N_2958,N_2902,N_2901);
nor U2959 (N_2959,N_2925,N_2924);
nand U2960 (N_2960,N_2930,N_2938);
and U2961 (N_2961,N_2882,N_2890);
nor U2962 (N_2962,N_2921,N_2927);
nor U2963 (N_2963,N_2906,N_2889);
xor U2964 (N_2964,N_2926,N_2886);
and U2965 (N_2965,N_2922,N_2918);
nor U2966 (N_2966,N_2898,N_2929);
and U2967 (N_2967,N_2919,N_2897);
nand U2968 (N_2968,N_2911,N_2883);
nand U2969 (N_2969,N_2904,N_2928);
and U2970 (N_2970,N_2928,N_2890);
nand U2971 (N_2971,N_2920,N_2890);
nand U2972 (N_2972,N_2912,N_2924);
nand U2973 (N_2973,N_2912,N_2880);
or U2974 (N_2974,N_2927,N_2920);
and U2975 (N_2975,N_2920,N_2900);
and U2976 (N_2976,N_2922,N_2904);
nand U2977 (N_2977,N_2925,N_2920);
nand U2978 (N_2978,N_2905,N_2910);
nand U2979 (N_2979,N_2880,N_2911);
nand U2980 (N_2980,N_2913,N_2918);
xor U2981 (N_2981,N_2900,N_2919);
and U2982 (N_2982,N_2919,N_2895);
nand U2983 (N_2983,N_2884,N_2902);
and U2984 (N_2984,N_2927,N_2883);
or U2985 (N_2985,N_2920,N_2887);
nand U2986 (N_2986,N_2899,N_2884);
or U2987 (N_2987,N_2907,N_2917);
xnor U2988 (N_2988,N_2917,N_2934);
or U2989 (N_2989,N_2920,N_2922);
and U2990 (N_2990,N_2923,N_2896);
and U2991 (N_2991,N_2907,N_2929);
or U2992 (N_2992,N_2927,N_2926);
or U2993 (N_2993,N_2935,N_2905);
or U2994 (N_2994,N_2923,N_2888);
or U2995 (N_2995,N_2896,N_2891);
nor U2996 (N_2996,N_2929,N_2896);
and U2997 (N_2997,N_2932,N_2912);
and U2998 (N_2998,N_2939,N_2903);
or U2999 (N_2999,N_2889,N_2891);
nor UO_0 (O_0,N_2952,N_2940);
and UO_1 (O_1,N_2976,N_2941);
nand UO_2 (O_2,N_2950,N_2996);
nor UO_3 (O_3,N_2972,N_2964);
nand UO_4 (O_4,N_2960,N_2967);
or UO_5 (O_5,N_2981,N_2977);
nand UO_6 (O_6,N_2962,N_2954);
nand UO_7 (O_7,N_2970,N_2994);
nor UO_8 (O_8,N_2942,N_2990);
nand UO_9 (O_9,N_2988,N_2997);
and UO_10 (O_10,N_2953,N_2995);
or UO_11 (O_11,N_2999,N_2969);
xor UO_12 (O_12,N_2945,N_2968);
or UO_13 (O_13,N_2979,N_2978);
nand UO_14 (O_14,N_2986,N_2966);
nor UO_15 (O_15,N_2959,N_2992);
or UO_16 (O_16,N_2985,N_2974);
nand UO_17 (O_17,N_2944,N_2971);
xnor UO_18 (O_18,N_2947,N_2989);
nor UO_19 (O_19,N_2963,N_2984);
nor UO_20 (O_20,N_2993,N_2983);
xnor UO_21 (O_21,N_2980,N_2958);
and UO_22 (O_22,N_2951,N_2965);
or UO_23 (O_23,N_2961,N_2943);
xor UO_24 (O_24,N_2973,N_2975);
or UO_25 (O_25,N_2982,N_2955);
nand UO_26 (O_26,N_2987,N_2998);
or UO_27 (O_27,N_2946,N_2991);
nor UO_28 (O_28,N_2957,N_2949);
or UO_29 (O_29,N_2956,N_2948);
and UO_30 (O_30,N_2969,N_2981);
or UO_31 (O_31,N_2964,N_2995);
or UO_32 (O_32,N_2983,N_2963);
xor UO_33 (O_33,N_2976,N_2995);
and UO_34 (O_34,N_2973,N_2993);
nor UO_35 (O_35,N_2998,N_2985);
nand UO_36 (O_36,N_2968,N_2960);
or UO_37 (O_37,N_2980,N_2994);
or UO_38 (O_38,N_2978,N_2968);
xnor UO_39 (O_39,N_2992,N_2952);
nand UO_40 (O_40,N_2966,N_2975);
nor UO_41 (O_41,N_2979,N_2946);
xnor UO_42 (O_42,N_2974,N_2990);
nor UO_43 (O_43,N_2990,N_2983);
and UO_44 (O_44,N_2959,N_2946);
and UO_45 (O_45,N_2984,N_2944);
or UO_46 (O_46,N_2963,N_2965);
nor UO_47 (O_47,N_2957,N_2966);
or UO_48 (O_48,N_2964,N_2949);
and UO_49 (O_49,N_2966,N_2962);
nand UO_50 (O_50,N_2955,N_2970);
or UO_51 (O_51,N_2979,N_2999);
and UO_52 (O_52,N_2963,N_2993);
nand UO_53 (O_53,N_2991,N_2992);
nand UO_54 (O_54,N_2981,N_2950);
xnor UO_55 (O_55,N_2959,N_2949);
nand UO_56 (O_56,N_2960,N_2951);
or UO_57 (O_57,N_2957,N_2972);
or UO_58 (O_58,N_2978,N_2986);
or UO_59 (O_59,N_2961,N_2998);
or UO_60 (O_60,N_2996,N_2976);
or UO_61 (O_61,N_2990,N_2985);
and UO_62 (O_62,N_2993,N_2945);
and UO_63 (O_63,N_2993,N_2964);
or UO_64 (O_64,N_2998,N_2963);
nor UO_65 (O_65,N_2942,N_2954);
and UO_66 (O_66,N_2991,N_2950);
xnor UO_67 (O_67,N_2991,N_2965);
nor UO_68 (O_68,N_2950,N_2970);
nand UO_69 (O_69,N_2966,N_2984);
nand UO_70 (O_70,N_2962,N_2945);
and UO_71 (O_71,N_2986,N_2956);
and UO_72 (O_72,N_2945,N_2996);
or UO_73 (O_73,N_2960,N_2959);
nor UO_74 (O_74,N_2947,N_2978);
or UO_75 (O_75,N_2960,N_2999);
nor UO_76 (O_76,N_2960,N_2996);
or UO_77 (O_77,N_2992,N_2957);
nand UO_78 (O_78,N_2980,N_2983);
nor UO_79 (O_79,N_2959,N_2954);
nand UO_80 (O_80,N_2980,N_2948);
or UO_81 (O_81,N_2980,N_2975);
or UO_82 (O_82,N_2983,N_2986);
xor UO_83 (O_83,N_2969,N_2972);
and UO_84 (O_84,N_2952,N_2953);
nor UO_85 (O_85,N_2947,N_2969);
xnor UO_86 (O_86,N_2949,N_2989);
xnor UO_87 (O_87,N_2975,N_2957);
and UO_88 (O_88,N_2967,N_2991);
nor UO_89 (O_89,N_2969,N_2970);
or UO_90 (O_90,N_2996,N_2956);
and UO_91 (O_91,N_2964,N_2942);
nor UO_92 (O_92,N_2994,N_2952);
or UO_93 (O_93,N_2986,N_2990);
and UO_94 (O_94,N_2968,N_2999);
nand UO_95 (O_95,N_2993,N_2989);
and UO_96 (O_96,N_2952,N_2947);
nand UO_97 (O_97,N_2996,N_2989);
nor UO_98 (O_98,N_2950,N_2956);
nor UO_99 (O_99,N_2942,N_2962);
or UO_100 (O_100,N_2973,N_2978);
or UO_101 (O_101,N_2985,N_2976);
xnor UO_102 (O_102,N_2952,N_2963);
nand UO_103 (O_103,N_2999,N_2985);
nor UO_104 (O_104,N_2956,N_2990);
or UO_105 (O_105,N_2985,N_2943);
and UO_106 (O_106,N_2972,N_2978);
and UO_107 (O_107,N_2953,N_2992);
nand UO_108 (O_108,N_2958,N_2955);
nand UO_109 (O_109,N_2978,N_2956);
nand UO_110 (O_110,N_2990,N_2950);
and UO_111 (O_111,N_2987,N_2976);
xor UO_112 (O_112,N_2963,N_2975);
and UO_113 (O_113,N_2951,N_2983);
nand UO_114 (O_114,N_2986,N_2947);
and UO_115 (O_115,N_2980,N_2987);
nand UO_116 (O_116,N_2949,N_2976);
and UO_117 (O_117,N_2985,N_2959);
nor UO_118 (O_118,N_2988,N_2980);
xnor UO_119 (O_119,N_2961,N_2969);
nor UO_120 (O_120,N_2968,N_2965);
or UO_121 (O_121,N_2970,N_2971);
nor UO_122 (O_122,N_2969,N_2949);
nand UO_123 (O_123,N_2963,N_2940);
nand UO_124 (O_124,N_2992,N_2954);
and UO_125 (O_125,N_2989,N_2971);
nand UO_126 (O_126,N_2953,N_2983);
nor UO_127 (O_127,N_2963,N_2962);
or UO_128 (O_128,N_2946,N_2982);
nor UO_129 (O_129,N_2994,N_2996);
or UO_130 (O_130,N_2959,N_2963);
nand UO_131 (O_131,N_2941,N_2994);
and UO_132 (O_132,N_2958,N_2952);
or UO_133 (O_133,N_2947,N_2987);
or UO_134 (O_134,N_2967,N_2971);
nor UO_135 (O_135,N_2949,N_2981);
nand UO_136 (O_136,N_2948,N_2966);
nor UO_137 (O_137,N_2973,N_2962);
nand UO_138 (O_138,N_2955,N_2981);
nand UO_139 (O_139,N_2961,N_2955);
or UO_140 (O_140,N_2993,N_2959);
nor UO_141 (O_141,N_2940,N_2996);
nor UO_142 (O_142,N_2953,N_2986);
or UO_143 (O_143,N_2986,N_2954);
nor UO_144 (O_144,N_2948,N_2951);
nor UO_145 (O_145,N_2974,N_2950);
xnor UO_146 (O_146,N_2971,N_2984);
nor UO_147 (O_147,N_2982,N_2995);
nand UO_148 (O_148,N_2980,N_2953);
or UO_149 (O_149,N_2956,N_2987);
and UO_150 (O_150,N_2997,N_2991);
or UO_151 (O_151,N_2961,N_2962);
nand UO_152 (O_152,N_2953,N_2964);
xnor UO_153 (O_153,N_2976,N_2962);
nand UO_154 (O_154,N_2999,N_2955);
or UO_155 (O_155,N_2987,N_2990);
xnor UO_156 (O_156,N_2950,N_2986);
or UO_157 (O_157,N_2991,N_2994);
and UO_158 (O_158,N_2940,N_2946);
nor UO_159 (O_159,N_2962,N_2968);
and UO_160 (O_160,N_2990,N_2992);
nand UO_161 (O_161,N_2949,N_2942);
nand UO_162 (O_162,N_2985,N_2995);
nor UO_163 (O_163,N_2975,N_2956);
nand UO_164 (O_164,N_2971,N_2955);
or UO_165 (O_165,N_2964,N_2965);
and UO_166 (O_166,N_2943,N_2956);
nand UO_167 (O_167,N_2965,N_2941);
nand UO_168 (O_168,N_2957,N_2993);
and UO_169 (O_169,N_2972,N_2968);
or UO_170 (O_170,N_2953,N_2944);
or UO_171 (O_171,N_2955,N_2977);
nor UO_172 (O_172,N_2957,N_2985);
nor UO_173 (O_173,N_2963,N_2979);
or UO_174 (O_174,N_2951,N_2966);
or UO_175 (O_175,N_2974,N_2966);
nor UO_176 (O_176,N_2989,N_2965);
xor UO_177 (O_177,N_2965,N_2974);
nor UO_178 (O_178,N_2952,N_2982);
xor UO_179 (O_179,N_2962,N_2977);
nand UO_180 (O_180,N_2997,N_2993);
and UO_181 (O_181,N_2944,N_2955);
xor UO_182 (O_182,N_2998,N_2954);
nand UO_183 (O_183,N_2945,N_2975);
and UO_184 (O_184,N_2967,N_2943);
nand UO_185 (O_185,N_2981,N_2958);
nor UO_186 (O_186,N_2993,N_2992);
nand UO_187 (O_187,N_2963,N_2992);
xor UO_188 (O_188,N_2997,N_2994);
or UO_189 (O_189,N_2993,N_2978);
nand UO_190 (O_190,N_2947,N_2951);
nor UO_191 (O_191,N_2956,N_2957);
nand UO_192 (O_192,N_2983,N_2985);
or UO_193 (O_193,N_2965,N_2979);
nand UO_194 (O_194,N_2964,N_2966);
or UO_195 (O_195,N_2994,N_2976);
or UO_196 (O_196,N_2949,N_2993);
and UO_197 (O_197,N_2941,N_2946);
or UO_198 (O_198,N_2998,N_2975);
and UO_199 (O_199,N_2998,N_2948);
or UO_200 (O_200,N_2982,N_2970);
and UO_201 (O_201,N_2951,N_2943);
xnor UO_202 (O_202,N_2965,N_2981);
nand UO_203 (O_203,N_2946,N_2973);
xor UO_204 (O_204,N_2953,N_2945);
nand UO_205 (O_205,N_2962,N_2948);
and UO_206 (O_206,N_2989,N_2973);
nor UO_207 (O_207,N_2971,N_2950);
and UO_208 (O_208,N_2956,N_2962);
nor UO_209 (O_209,N_2961,N_2997);
nand UO_210 (O_210,N_2944,N_2992);
or UO_211 (O_211,N_2951,N_2987);
or UO_212 (O_212,N_2951,N_2986);
xor UO_213 (O_213,N_2944,N_2978);
nand UO_214 (O_214,N_2955,N_2996);
and UO_215 (O_215,N_2995,N_2973);
nor UO_216 (O_216,N_2992,N_2987);
nand UO_217 (O_217,N_2974,N_2944);
or UO_218 (O_218,N_2979,N_2976);
xnor UO_219 (O_219,N_2949,N_2988);
or UO_220 (O_220,N_2989,N_2987);
nor UO_221 (O_221,N_2959,N_2962);
and UO_222 (O_222,N_2959,N_2998);
and UO_223 (O_223,N_2951,N_2995);
and UO_224 (O_224,N_2986,N_2946);
and UO_225 (O_225,N_2944,N_2973);
nand UO_226 (O_226,N_2956,N_2966);
or UO_227 (O_227,N_2970,N_2985);
or UO_228 (O_228,N_2998,N_2967);
nor UO_229 (O_229,N_2940,N_2956);
or UO_230 (O_230,N_2978,N_2962);
or UO_231 (O_231,N_2970,N_2961);
and UO_232 (O_232,N_2948,N_2974);
nor UO_233 (O_233,N_2965,N_2957);
and UO_234 (O_234,N_2952,N_2945);
and UO_235 (O_235,N_2978,N_2964);
nor UO_236 (O_236,N_2989,N_2978);
nor UO_237 (O_237,N_2976,N_2952);
nand UO_238 (O_238,N_2960,N_2984);
nor UO_239 (O_239,N_2953,N_2967);
or UO_240 (O_240,N_2959,N_2964);
nand UO_241 (O_241,N_2995,N_2978);
nor UO_242 (O_242,N_2995,N_2996);
and UO_243 (O_243,N_2957,N_2976);
nor UO_244 (O_244,N_2996,N_2961);
nor UO_245 (O_245,N_2956,N_2976);
and UO_246 (O_246,N_2994,N_2965);
or UO_247 (O_247,N_2975,N_2968);
and UO_248 (O_248,N_2941,N_2978);
or UO_249 (O_249,N_2995,N_2942);
and UO_250 (O_250,N_2948,N_2983);
nor UO_251 (O_251,N_2945,N_2947);
xnor UO_252 (O_252,N_2951,N_2984);
xnor UO_253 (O_253,N_2979,N_2970);
xor UO_254 (O_254,N_2962,N_2983);
xor UO_255 (O_255,N_2943,N_2944);
and UO_256 (O_256,N_2970,N_2940);
or UO_257 (O_257,N_2948,N_2986);
or UO_258 (O_258,N_2987,N_2983);
nor UO_259 (O_259,N_2969,N_2959);
or UO_260 (O_260,N_2977,N_2959);
nand UO_261 (O_261,N_2974,N_2968);
and UO_262 (O_262,N_2971,N_2986);
or UO_263 (O_263,N_2944,N_2956);
nor UO_264 (O_264,N_2986,N_2976);
xnor UO_265 (O_265,N_2940,N_2944);
nor UO_266 (O_266,N_2943,N_2942);
nand UO_267 (O_267,N_2971,N_2992);
and UO_268 (O_268,N_2968,N_2970);
nor UO_269 (O_269,N_2971,N_2966);
and UO_270 (O_270,N_2993,N_2962);
nand UO_271 (O_271,N_2988,N_2960);
nor UO_272 (O_272,N_2949,N_2977);
nand UO_273 (O_273,N_2961,N_2994);
and UO_274 (O_274,N_2983,N_2952);
and UO_275 (O_275,N_2991,N_2958);
nor UO_276 (O_276,N_2993,N_2987);
nor UO_277 (O_277,N_2941,N_2986);
nand UO_278 (O_278,N_2965,N_2978);
xor UO_279 (O_279,N_2999,N_2981);
nor UO_280 (O_280,N_2962,N_2965);
or UO_281 (O_281,N_2940,N_2967);
or UO_282 (O_282,N_2946,N_2953);
or UO_283 (O_283,N_2973,N_2981);
nor UO_284 (O_284,N_2967,N_2997);
or UO_285 (O_285,N_2982,N_2981);
and UO_286 (O_286,N_2953,N_2961);
nor UO_287 (O_287,N_2960,N_2964);
nand UO_288 (O_288,N_2999,N_2982);
xnor UO_289 (O_289,N_2954,N_2973);
or UO_290 (O_290,N_2968,N_2941);
and UO_291 (O_291,N_2996,N_2953);
nand UO_292 (O_292,N_2986,N_2940);
or UO_293 (O_293,N_2996,N_2975);
and UO_294 (O_294,N_2975,N_2985);
or UO_295 (O_295,N_2949,N_2965);
nor UO_296 (O_296,N_2957,N_2970);
and UO_297 (O_297,N_2993,N_2961);
or UO_298 (O_298,N_2981,N_2974);
nor UO_299 (O_299,N_2972,N_2960);
nor UO_300 (O_300,N_2985,N_2946);
and UO_301 (O_301,N_2985,N_2993);
nor UO_302 (O_302,N_2950,N_2964);
nand UO_303 (O_303,N_2992,N_2973);
nand UO_304 (O_304,N_2964,N_2943);
and UO_305 (O_305,N_2997,N_2976);
nor UO_306 (O_306,N_2941,N_2990);
nand UO_307 (O_307,N_2968,N_2940);
xnor UO_308 (O_308,N_2947,N_2984);
xnor UO_309 (O_309,N_2978,N_2961);
nor UO_310 (O_310,N_2990,N_2960);
or UO_311 (O_311,N_2951,N_2981);
or UO_312 (O_312,N_2968,N_2984);
and UO_313 (O_313,N_2940,N_2954);
or UO_314 (O_314,N_2995,N_2962);
and UO_315 (O_315,N_2972,N_2941);
or UO_316 (O_316,N_2993,N_2990);
nor UO_317 (O_317,N_2999,N_2978);
nor UO_318 (O_318,N_2995,N_2969);
or UO_319 (O_319,N_2967,N_2963);
and UO_320 (O_320,N_2970,N_2958);
or UO_321 (O_321,N_2946,N_2954);
nand UO_322 (O_322,N_2967,N_2976);
nand UO_323 (O_323,N_2997,N_2958);
and UO_324 (O_324,N_2954,N_2947);
nand UO_325 (O_325,N_2996,N_2942);
nor UO_326 (O_326,N_2996,N_2944);
nor UO_327 (O_327,N_2944,N_2958);
or UO_328 (O_328,N_2954,N_2968);
and UO_329 (O_329,N_2940,N_2982);
and UO_330 (O_330,N_2958,N_2962);
nand UO_331 (O_331,N_2990,N_2970);
and UO_332 (O_332,N_2953,N_2970);
or UO_333 (O_333,N_2975,N_2941);
and UO_334 (O_334,N_2980,N_2950);
and UO_335 (O_335,N_2944,N_2951);
nor UO_336 (O_336,N_2943,N_2971);
or UO_337 (O_337,N_2986,N_2988);
xor UO_338 (O_338,N_2962,N_2988);
nand UO_339 (O_339,N_2959,N_2955);
xor UO_340 (O_340,N_2991,N_2987);
nor UO_341 (O_341,N_2944,N_2970);
nand UO_342 (O_342,N_2985,N_2987);
or UO_343 (O_343,N_2947,N_2962);
or UO_344 (O_344,N_2959,N_2995);
and UO_345 (O_345,N_2964,N_2985);
nor UO_346 (O_346,N_2966,N_2968);
nand UO_347 (O_347,N_2989,N_2982);
and UO_348 (O_348,N_2949,N_2995);
and UO_349 (O_349,N_2948,N_2975);
nor UO_350 (O_350,N_2999,N_2945);
and UO_351 (O_351,N_2978,N_2982);
or UO_352 (O_352,N_2969,N_2948);
xnor UO_353 (O_353,N_2988,N_2981);
nor UO_354 (O_354,N_2999,N_2958);
nor UO_355 (O_355,N_2969,N_2946);
xor UO_356 (O_356,N_2986,N_2960);
nand UO_357 (O_357,N_2985,N_2948);
nor UO_358 (O_358,N_2985,N_2968);
nand UO_359 (O_359,N_2948,N_2955);
xnor UO_360 (O_360,N_2955,N_2985);
nand UO_361 (O_361,N_2982,N_2993);
or UO_362 (O_362,N_2956,N_2979);
nor UO_363 (O_363,N_2958,N_2988);
and UO_364 (O_364,N_2983,N_2969);
and UO_365 (O_365,N_2947,N_2960);
nand UO_366 (O_366,N_2991,N_2986);
nand UO_367 (O_367,N_2979,N_2958);
nor UO_368 (O_368,N_2969,N_2996);
or UO_369 (O_369,N_2964,N_2956);
nor UO_370 (O_370,N_2960,N_2956);
nor UO_371 (O_371,N_2975,N_2976);
or UO_372 (O_372,N_2942,N_2968);
and UO_373 (O_373,N_2944,N_2963);
xnor UO_374 (O_374,N_2958,N_2964);
and UO_375 (O_375,N_2993,N_2974);
nand UO_376 (O_376,N_2994,N_2948);
and UO_377 (O_377,N_2983,N_2943);
or UO_378 (O_378,N_2944,N_2957);
nor UO_379 (O_379,N_2968,N_2996);
or UO_380 (O_380,N_2944,N_2950);
nor UO_381 (O_381,N_2952,N_2957);
nor UO_382 (O_382,N_2989,N_2966);
and UO_383 (O_383,N_2994,N_2990);
or UO_384 (O_384,N_2954,N_2966);
or UO_385 (O_385,N_2976,N_2946);
and UO_386 (O_386,N_2990,N_2976);
and UO_387 (O_387,N_2968,N_2947);
nor UO_388 (O_388,N_2962,N_2980);
and UO_389 (O_389,N_2959,N_2979);
and UO_390 (O_390,N_2971,N_2990);
nor UO_391 (O_391,N_2980,N_2954);
nor UO_392 (O_392,N_2997,N_2955);
or UO_393 (O_393,N_2941,N_2983);
or UO_394 (O_394,N_2970,N_2992);
or UO_395 (O_395,N_2966,N_2993);
nand UO_396 (O_396,N_2995,N_2956);
xnor UO_397 (O_397,N_2941,N_2959);
or UO_398 (O_398,N_2965,N_2943);
nand UO_399 (O_399,N_2966,N_2970);
nand UO_400 (O_400,N_2990,N_2967);
nor UO_401 (O_401,N_2991,N_2978);
nor UO_402 (O_402,N_2953,N_2998);
nor UO_403 (O_403,N_2981,N_2972);
nor UO_404 (O_404,N_2947,N_2959);
and UO_405 (O_405,N_2955,N_2990);
and UO_406 (O_406,N_2943,N_2997);
or UO_407 (O_407,N_2987,N_2962);
nand UO_408 (O_408,N_2976,N_2972);
nor UO_409 (O_409,N_2980,N_2968);
or UO_410 (O_410,N_2970,N_2952);
and UO_411 (O_411,N_2969,N_2962);
nand UO_412 (O_412,N_2980,N_2976);
nor UO_413 (O_413,N_2978,N_2940);
or UO_414 (O_414,N_2974,N_2975);
nor UO_415 (O_415,N_2961,N_2950);
or UO_416 (O_416,N_2973,N_2949);
nor UO_417 (O_417,N_2975,N_2961);
and UO_418 (O_418,N_2946,N_2950);
nor UO_419 (O_419,N_2971,N_2951);
nand UO_420 (O_420,N_2940,N_2988);
or UO_421 (O_421,N_2944,N_2983);
xnor UO_422 (O_422,N_2953,N_2993);
nand UO_423 (O_423,N_2999,N_2986);
and UO_424 (O_424,N_2974,N_2988);
nor UO_425 (O_425,N_2995,N_2986);
or UO_426 (O_426,N_2974,N_2962);
and UO_427 (O_427,N_2994,N_2944);
and UO_428 (O_428,N_2977,N_2945);
nor UO_429 (O_429,N_2984,N_2996);
and UO_430 (O_430,N_2955,N_2952);
nor UO_431 (O_431,N_2964,N_2963);
or UO_432 (O_432,N_2992,N_2977);
nand UO_433 (O_433,N_2973,N_2985);
and UO_434 (O_434,N_2996,N_2985);
and UO_435 (O_435,N_2960,N_2977);
nand UO_436 (O_436,N_2940,N_2959);
nor UO_437 (O_437,N_2951,N_2967);
nand UO_438 (O_438,N_2956,N_2963);
nor UO_439 (O_439,N_2998,N_2972);
or UO_440 (O_440,N_2994,N_2973);
and UO_441 (O_441,N_2994,N_2950);
nor UO_442 (O_442,N_2997,N_2963);
nor UO_443 (O_443,N_2982,N_2980);
nor UO_444 (O_444,N_2984,N_2993);
nor UO_445 (O_445,N_2970,N_2984);
and UO_446 (O_446,N_2952,N_2959);
or UO_447 (O_447,N_2998,N_2992);
or UO_448 (O_448,N_2981,N_2971);
nand UO_449 (O_449,N_2976,N_2988);
or UO_450 (O_450,N_2985,N_2986);
nor UO_451 (O_451,N_2998,N_2978);
nor UO_452 (O_452,N_2971,N_2997);
and UO_453 (O_453,N_2942,N_2979);
nor UO_454 (O_454,N_2946,N_2955);
and UO_455 (O_455,N_2995,N_2967);
nand UO_456 (O_456,N_2988,N_2991);
and UO_457 (O_457,N_2951,N_2958);
nor UO_458 (O_458,N_2979,N_2945);
nor UO_459 (O_459,N_2965,N_2983);
nor UO_460 (O_460,N_2995,N_2957);
nand UO_461 (O_461,N_2972,N_2944);
nor UO_462 (O_462,N_2988,N_2950);
and UO_463 (O_463,N_2982,N_2941);
or UO_464 (O_464,N_2974,N_2957);
nand UO_465 (O_465,N_2998,N_2982);
nor UO_466 (O_466,N_2993,N_2958);
or UO_467 (O_467,N_2979,N_2982);
nor UO_468 (O_468,N_2943,N_2958);
and UO_469 (O_469,N_2959,N_2971);
nand UO_470 (O_470,N_2972,N_2946);
or UO_471 (O_471,N_2953,N_2988);
nand UO_472 (O_472,N_2975,N_2951);
xnor UO_473 (O_473,N_2992,N_2968);
nand UO_474 (O_474,N_2973,N_2948);
and UO_475 (O_475,N_2948,N_2941);
nand UO_476 (O_476,N_2972,N_2977);
and UO_477 (O_477,N_2999,N_2998);
nand UO_478 (O_478,N_2955,N_2989);
nor UO_479 (O_479,N_2954,N_2960);
and UO_480 (O_480,N_2987,N_2961);
and UO_481 (O_481,N_2997,N_2951);
or UO_482 (O_482,N_2987,N_2968);
and UO_483 (O_483,N_2986,N_2963);
nand UO_484 (O_484,N_2947,N_2993);
nand UO_485 (O_485,N_2960,N_2943);
nand UO_486 (O_486,N_2957,N_2973);
nand UO_487 (O_487,N_2974,N_2996);
nand UO_488 (O_488,N_2989,N_2992);
xor UO_489 (O_489,N_2956,N_2953);
and UO_490 (O_490,N_2977,N_2991);
and UO_491 (O_491,N_2961,N_2995);
nand UO_492 (O_492,N_2975,N_2983);
nand UO_493 (O_493,N_2949,N_2940);
and UO_494 (O_494,N_2983,N_2957);
xnor UO_495 (O_495,N_2947,N_2958);
nand UO_496 (O_496,N_2983,N_2989);
and UO_497 (O_497,N_2944,N_2987);
nand UO_498 (O_498,N_2944,N_2947);
and UO_499 (O_499,N_2970,N_2995);
endmodule